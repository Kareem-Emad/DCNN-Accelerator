
-- 
-- Definition of  Controller
-- 
--      Sat May 11 13:08:15 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Queue_5 is
   port (
      d : IN std_logic_vector (15 DOWNTO 0) ;
      q_0_15 : OUT std_logic ;
      q_0_14 : OUT std_logic ;
      q_0_13 : OUT std_logic ;
      q_0_12 : OUT std_logic ;
      q_0_11 : OUT std_logic ;
      q_0_10 : OUT std_logic ;
      q_0_9 : OUT std_logic ;
      q_0_8 : OUT std_logic ;
      q_0_7 : OUT std_logic ;
      q_0_6 : OUT std_logic ;
      q_0_5 : OUT std_logic ;
      q_0_4 : OUT std_logic ;
      q_0_3 : OUT std_logic ;
      q_0_2 : OUT std_logic ;
      q_0_1 : OUT std_logic ;
      q_0_0 : OUT std_logic ;
      q_1_15 : OUT std_logic ;
      q_1_14 : OUT std_logic ;
      q_1_13 : OUT std_logic ;
      q_1_12 : OUT std_logic ;
      q_1_11 : OUT std_logic ;
      q_1_10 : OUT std_logic ;
      q_1_9 : OUT std_logic ;
      q_1_8 : OUT std_logic ;
      q_1_7 : OUT std_logic ;
      q_1_6 : OUT std_logic ;
      q_1_5 : OUT std_logic ;
      q_1_4 : OUT std_logic ;
      q_1_3 : OUT std_logic ;
      q_1_2 : OUT std_logic ;
      q_1_1 : OUT std_logic ;
      q_1_0 : OUT std_logic ;
      q_2_15 : OUT std_logic ;
      q_2_14 : OUT std_logic ;
      q_2_13 : OUT std_logic ;
      q_2_12 : OUT std_logic ;
      q_2_11 : OUT std_logic ;
      q_2_10 : OUT std_logic ;
      q_2_9 : OUT std_logic ;
      q_2_8 : OUT std_logic ;
      q_2_7 : OUT std_logic ;
      q_2_6 : OUT std_logic ;
      q_2_5 : OUT std_logic ;
      q_2_4 : OUT std_logic ;
      q_2_3 : OUT std_logic ;
      q_2_2 : OUT std_logic ;
      q_2_1 : OUT std_logic ;
      q_2_0 : OUT std_logic ;
      q_3_15 : OUT std_logic ;
      q_3_14 : OUT std_logic ;
      q_3_13 : OUT std_logic ;
      q_3_12 : OUT std_logic ;
      q_3_11 : OUT std_logic ;
      q_3_10 : OUT std_logic ;
      q_3_9 : OUT std_logic ;
      q_3_8 : OUT std_logic ;
      q_3_7 : OUT std_logic ;
      q_3_6 : OUT std_logic ;
      q_3_5 : OUT std_logic ;
      q_3_4 : OUT std_logic ;
      q_3_3 : OUT std_logic ;
      q_3_2 : OUT std_logic ;
      q_3_1 : OUT std_logic ;
      q_3_0 : OUT std_logic ;
      q_4_15 : OUT std_logic ;
      q_4_14 : OUT std_logic ;
      q_4_13 : OUT std_logic ;
      q_4_12 : OUT std_logic ;
      q_4_11 : OUT std_logic ;
      q_4_10 : OUT std_logic ;
      q_4_9 : OUT std_logic ;
      q_4_8 : OUT std_logic ;
      q_4_7 : OUT std_logic ;
      q_4_6 : OUT std_logic ;
      q_4_5 : OUT std_logic ;
      q_4_4 : OUT std_logic ;
      q_4_3 : OUT std_logic ;
      q_4_2 : OUT std_logic ;
      q_4_1 : OUT std_logic ;
      q_4_0 : OUT std_logic ;
      clk : IN std_logic ;
      load : IN std_logic ;
      reset : IN std_logic) ;
end Queue_5 ;

architecture Dataflow of Queue_5 is
   signal q_0_15_EXMPLR, q_0_14_EXMPLR, q_0_13_EXMPLR, q_0_12_EXMPLR, 
      q_0_11_EXMPLR, q_0_10_EXMPLR, q_0_9_EXMPLR, q_0_8_EXMPLR, q_0_7_EXMPLR, 
      q_0_6_EXMPLR, q_0_5_EXMPLR, q_0_4_EXMPLR, q_0_3_EXMPLR, q_0_2_EXMPLR, 
      q_0_1_EXMPLR, q_0_0_EXMPLR, q_1_15_EXMPLR, q_1_14_EXMPLR, 
      q_1_13_EXMPLR, q_1_12_EXMPLR, q_1_11_EXMPLR, q_1_10_EXMPLR, 
      q_1_9_EXMPLR, q_1_8_EXMPLR, q_1_7_EXMPLR, q_1_6_EXMPLR, q_1_5_EXMPLR, 
      q_1_4_EXMPLR, q_1_3_EXMPLR, q_1_2_EXMPLR, q_1_1_EXMPLR, q_1_0_EXMPLR, 
      q_2_15_EXMPLR, q_2_14_EXMPLR, q_2_13_EXMPLR, q_2_12_EXMPLR, 
      q_2_11_EXMPLR, q_2_10_EXMPLR, q_2_9_EXMPLR, q_2_8_EXMPLR, q_2_7_EXMPLR, 
      q_2_6_EXMPLR, q_2_5_EXMPLR, q_2_4_EXMPLR, q_2_3_EXMPLR, q_2_2_EXMPLR, 
      q_2_1_EXMPLR, q_2_0_EXMPLR, q_3_15_EXMPLR, q_3_14_EXMPLR, 
      q_3_13_EXMPLR, q_3_12_EXMPLR, q_3_11_EXMPLR, q_3_10_EXMPLR, 
      q_3_9_EXMPLR, q_3_8_EXMPLR, q_3_7_EXMPLR, q_3_6_EXMPLR, q_3_5_EXMPLR, 
      q_3_4_EXMPLR, q_3_3_EXMPLR, q_3_2_EXMPLR, q_3_1_EXMPLR, q_3_0_EXMPLR, 
      q_4_15_EXMPLR, q_4_14_EXMPLR, q_4_13_EXMPLR, q_4_12_EXMPLR, 
      q_4_11_EXMPLR, q_4_10_EXMPLR, q_4_9_EXMPLR, q_4_8_EXMPLR, q_4_7_EXMPLR, 
      q_4_6_EXMPLR, q_4_5_EXMPLR, q_4_4_EXMPLR, q_4_3_EXMPLR, q_4_2_EXMPLR, 
      q_4_1_EXMPLR, q_4_0_EXMPLR, nx393, nx403, nx413, nx423, nx433, nx443, 
      nx453, nx463, nx473, nx483, nx493, nx503, nx513, nx523, nx533, nx543, 
      nx553, nx563, nx573, nx583, nx593, nx603, nx613, nx623, nx633, nx643, 
      nx653, nx663, nx673, nx683, nx693, nx703, nx713, nx723, nx733, nx743, 
      nx753, nx763, nx773, nx783, nx793, nx803, nx813, nx823, nx833, nx843, 
      nx853, nx863, nx873, nx883, nx893, nx903, nx913, nx923, nx933, nx943, 
      nx953, nx963, nx973, nx983, nx993, nx1003, nx1013, nx1023, nx1033, 
      nx1043, nx1053, nx1063, nx1073, nx1083, nx1093, nx1103, nx1113, nx1123, 
      nx1133, nx1143, nx1153, nx1163, nx1173, nx1183, nx1440, nx1442, nx1444, 
      nx1446, nx1448, nx1450, nx1452, nx1454, nx1456, nx1458, nx1460, nx1462, 
      nx1466, nx1468, nx1470, nx1472, nx1474, nx1476, nx1478, nx1480, nx1482, 
      nx1484, nx1486, nx1488, nx1492, nx1494, nx1496, nx1498, nx1500, nx1502, 
      nx1504, nx1506, nx1508, nx1510, nx1512, nx1514, nx1516, nx1518, nx1520, 
      nx1522, nx1524, nx1526: std_logic ;

begin
   q_0_15 <= q_0_15_EXMPLR ;
   q_0_14 <= q_0_14_EXMPLR ;
   q_0_13 <= q_0_13_EXMPLR ;
   q_0_12 <= q_0_12_EXMPLR ;
   q_0_11 <= q_0_11_EXMPLR ;
   q_0_10 <= q_0_10_EXMPLR ;
   q_0_9 <= q_0_9_EXMPLR ;
   q_0_8 <= q_0_8_EXMPLR ;
   q_0_7 <= q_0_7_EXMPLR ;
   q_0_6 <= q_0_6_EXMPLR ;
   q_0_5 <= q_0_5_EXMPLR ;
   q_0_4 <= q_0_4_EXMPLR ;
   q_0_3 <= q_0_3_EXMPLR ;
   q_0_2 <= q_0_2_EXMPLR ;
   q_0_1 <= q_0_1_EXMPLR ;
   q_0_0 <= q_0_0_EXMPLR ;
   q_1_15 <= q_1_15_EXMPLR ;
   q_1_14 <= q_1_14_EXMPLR ;
   q_1_13 <= q_1_13_EXMPLR ;
   q_1_12 <= q_1_12_EXMPLR ;
   q_1_11 <= q_1_11_EXMPLR ;
   q_1_10 <= q_1_10_EXMPLR ;
   q_1_9 <= q_1_9_EXMPLR ;
   q_1_8 <= q_1_8_EXMPLR ;
   q_1_7 <= q_1_7_EXMPLR ;
   q_1_6 <= q_1_6_EXMPLR ;
   q_1_5 <= q_1_5_EXMPLR ;
   q_1_4 <= q_1_4_EXMPLR ;
   q_1_3 <= q_1_3_EXMPLR ;
   q_1_2 <= q_1_2_EXMPLR ;
   q_1_1 <= q_1_1_EXMPLR ;
   q_1_0 <= q_1_0_EXMPLR ;
   q_2_15 <= q_2_15_EXMPLR ;
   q_2_14 <= q_2_14_EXMPLR ;
   q_2_13 <= q_2_13_EXMPLR ;
   q_2_12 <= q_2_12_EXMPLR ;
   q_2_11 <= q_2_11_EXMPLR ;
   q_2_10 <= q_2_10_EXMPLR ;
   q_2_9 <= q_2_9_EXMPLR ;
   q_2_8 <= q_2_8_EXMPLR ;
   q_2_7 <= q_2_7_EXMPLR ;
   q_2_6 <= q_2_6_EXMPLR ;
   q_2_5 <= q_2_5_EXMPLR ;
   q_2_4 <= q_2_4_EXMPLR ;
   q_2_3 <= q_2_3_EXMPLR ;
   q_2_2 <= q_2_2_EXMPLR ;
   q_2_1 <= q_2_1_EXMPLR ;
   q_2_0 <= q_2_0_EXMPLR ;
   q_3_15 <= q_3_15_EXMPLR ;
   q_3_14 <= q_3_14_EXMPLR ;
   q_3_13 <= q_3_13_EXMPLR ;
   q_3_12 <= q_3_12_EXMPLR ;
   q_3_11 <= q_3_11_EXMPLR ;
   q_3_10 <= q_3_10_EXMPLR ;
   q_3_9 <= q_3_9_EXMPLR ;
   q_3_8 <= q_3_8_EXMPLR ;
   q_3_7 <= q_3_7_EXMPLR ;
   q_3_6 <= q_3_6_EXMPLR ;
   q_3_5 <= q_3_5_EXMPLR ;
   q_3_4 <= q_3_4_EXMPLR ;
   q_3_3 <= q_3_3_EXMPLR ;
   q_3_2 <= q_3_2_EXMPLR ;
   q_3_1 <= q_3_1_EXMPLR ;
   q_3_0 <= q_3_0_EXMPLR ;
   q_4_15 <= q_4_15_EXMPLR ;
   q_4_14 <= q_4_14_EXMPLR ;
   q_4_13 <= q_4_13_EXMPLR ;
   q_4_12 <= q_4_12_EXMPLR ;
   q_4_11 <= q_4_11_EXMPLR ;
   q_4_10 <= q_4_10_EXMPLR ;
   q_4_9 <= q_4_9_EXMPLR ;
   q_4_8 <= q_4_8_EXMPLR ;
   q_4_7 <= q_4_7_EXMPLR ;
   q_4_6 <= q_4_6_EXMPLR ;
   q_4_5 <= q_4_5_EXMPLR ;
   q_4_4 <= q_4_4_EXMPLR ;
   q_4_3 <= q_4_3_EXMPLR ;
   q_4_2 <= q_4_2_EXMPLR ;
   q_4_1 <= q_4_1_EXMPLR ;
   q_4_0 <= q_4_0_EXMPLR ;
   gen_regs_4_regi_reg_q_0 : dffr port map ( Q=>q_4_0_EXMPLR, QB=>OPEN, D=>
      nx433, CLK=>nx1492, R=>nx1466);
   ix434 : mux21_ni port map ( Y=>nx433, A0=>q_4_0_EXMPLR, A1=>q_3_0_EXMPLR, 
      S0=>nx1440);
   gen_regs_3_regi_reg_q_0 : dffr port map ( Q=>q_3_0_EXMPLR, QB=>OPEN, D=>
      nx423, CLK=>nx1492, R=>nx1466);
   ix424 : mux21_ni port map ( Y=>nx423, A0=>q_3_0_EXMPLR, A1=>q_2_0_EXMPLR, 
      S0=>nx1440);
   gen_regs_2_regi_reg_q_0 : dffr port map ( Q=>q_2_0_EXMPLR, QB=>OPEN, D=>
      nx413, CLK=>nx1492, R=>nx1466);
   ix414 : mux21_ni port map ( Y=>nx413, A0=>q_2_0_EXMPLR, A1=>q_1_0_EXMPLR, 
      S0=>nx1440);
   gen_regs_1_regi_reg_q_0 : dffr port map ( Q=>q_1_0_EXMPLR, QB=>OPEN, D=>
      nx403, CLK=>nx1492, R=>nx1466);
   ix404 : mux21_ni port map ( Y=>nx403, A0=>q_1_0_EXMPLR, A1=>q_0_0_EXMPLR, 
      S0=>nx1440);
   reg0_reg_q_0 : dffr port map ( Q=>q_0_0_EXMPLR, QB=>OPEN, D=>nx393, CLK=>
      nx1492, R=>nx1466);
   ix394 : mux21_ni port map ( Y=>nx393, A0=>q_0_0_EXMPLR, A1=>d(0), S0=>
      nx1440);
   gen_regs_4_regi_reg_q_1 : dffr port map ( Q=>q_4_1_EXMPLR, QB=>OPEN, D=>
      nx483, CLK=>nx1494, R=>nx1468);
   ix484 : mux21_ni port map ( Y=>nx483, A0=>q_4_1_EXMPLR, A1=>q_3_1_EXMPLR, 
      S0=>nx1442);
   gen_regs_3_regi_reg_q_1 : dffr port map ( Q=>q_3_1_EXMPLR, QB=>OPEN, D=>
      nx473, CLK=>nx1494, R=>nx1468);
   ix474 : mux21_ni port map ( Y=>nx473, A0=>q_3_1_EXMPLR, A1=>q_2_1_EXMPLR, 
      S0=>nx1442);
   gen_regs_2_regi_reg_q_1 : dffr port map ( Q=>q_2_1_EXMPLR, QB=>OPEN, D=>
      nx463, CLK=>nx1494, R=>nx1468);
   ix464 : mux21_ni port map ( Y=>nx463, A0=>q_2_1_EXMPLR, A1=>q_1_1_EXMPLR, 
      S0=>nx1442);
   gen_regs_1_regi_reg_q_1 : dffr port map ( Q=>q_1_1_EXMPLR, QB=>OPEN, D=>
      nx453, CLK=>nx1492, R=>nx1466);
   ix454 : mux21_ni port map ( Y=>nx453, A0=>q_1_1_EXMPLR, A1=>q_0_1_EXMPLR, 
      S0=>nx1440);
   reg0_reg_q_1 : dffr port map ( Q=>q_0_1_EXMPLR, QB=>OPEN, D=>nx443, CLK=>
      nx1492, R=>nx1466);
   ix444 : mux21_ni port map ( Y=>nx443, A0=>q_0_1_EXMPLR, A1=>d(1), S0=>
      nx1440);
   gen_regs_4_regi_reg_q_2 : dffr port map ( Q=>q_4_2_EXMPLR, QB=>OPEN, D=>
      nx533, CLK=>nx1496, R=>nx1470);
   ix534 : mux21_ni port map ( Y=>nx533, A0=>q_4_2_EXMPLR, A1=>q_3_2_EXMPLR, 
      S0=>nx1444);
   gen_regs_3_regi_reg_q_2 : dffr port map ( Q=>q_3_2_EXMPLR, QB=>OPEN, D=>
      nx523, CLK=>nx1494, R=>nx1468);
   ix524 : mux21_ni port map ( Y=>nx523, A0=>q_3_2_EXMPLR, A1=>q_2_2_EXMPLR, 
      S0=>nx1442);
   gen_regs_2_regi_reg_q_2 : dffr port map ( Q=>q_2_2_EXMPLR, QB=>OPEN, D=>
      nx513, CLK=>nx1494, R=>nx1468);
   ix514 : mux21_ni port map ( Y=>nx513, A0=>q_2_2_EXMPLR, A1=>q_1_2_EXMPLR, 
      S0=>nx1442);
   gen_regs_1_regi_reg_q_2 : dffr port map ( Q=>q_1_2_EXMPLR, QB=>OPEN, D=>
      nx503, CLK=>nx1494, R=>nx1468);
   ix504 : mux21_ni port map ( Y=>nx503, A0=>q_1_2_EXMPLR, A1=>q_0_2_EXMPLR, 
      S0=>nx1442);
   reg0_reg_q_2 : dffr port map ( Q=>q_0_2_EXMPLR, QB=>OPEN, D=>nx493, CLK=>
      nx1494, R=>nx1468);
   ix494 : mux21_ni port map ( Y=>nx493, A0=>q_0_2_EXMPLR, A1=>d(2), S0=>
      nx1442);
   gen_regs_4_regi_reg_q_3 : dffr port map ( Q=>q_4_3_EXMPLR, QB=>OPEN, D=>
      nx583, CLK=>nx1496, R=>nx1470);
   ix584 : mux21_ni port map ( Y=>nx583, A0=>q_4_3_EXMPLR, A1=>q_3_3_EXMPLR, 
      S0=>nx1444);
   gen_regs_3_regi_reg_q_3 : dffr port map ( Q=>q_3_3_EXMPLR, QB=>OPEN, D=>
      nx573, CLK=>nx1496, R=>nx1470);
   ix574 : mux21_ni port map ( Y=>nx573, A0=>q_3_3_EXMPLR, A1=>q_2_3_EXMPLR, 
      S0=>nx1444);
   gen_regs_2_regi_reg_q_3 : dffr port map ( Q=>q_2_3_EXMPLR, QB=>OPEN, D=>
      nx563, CLK=>nx1496, R=>nx1470);
   ix564 : mux21_ni port map ( Y=>nx563, A0=>q_2_3_EXMPLR, A1=>q_1_3_EXMPLR, 
      S0=>nx1444);
   gen_regs_1_regi_reg_q_3 : dffr port map ( Q=>q_1_3_EXMPLR, QB=>OPEN, D=>
      nx553, CLK=>nx1496, R=>nx1470);
   ix554 : mux21_ni port map ( Y=>nx553, A0=>q_1_3_EXMPLR, A1=>q_0_3_EXMPLR, 
      S0=>nx1444);
   reg0_reg_q_3 : dffr port map ( Q=>q_0_3_EXMPLR, QB=>OPEN, D=>nx543, CLK=>
      nx1496, R=>nx1470);
   ix544 : mux21_ni port map ( Y=>nx543, A0=>q_0_3_EXMPLR, A1=>d(3), S0=>
      nx1444);
   gen_regs_4_regi_reg_q_4 : dffr port map ( Q=>q_4_4_EXMPLR, QB=>OPEN, D=>
      nx633, CLK=>nx1498, R=>nx1472);
   ix634 : mux21_ni port map ( Y=>nx633, A0=>q_4_4_EXMPLR, A1=>q_3_4_EXMPLR, 
      S0=>nx1446);
   gen_regs_3_regi_reg_q_4 : dffr port map ( Q=>q_3_4_EXMPLR, QB=>OPEN, D=>
      nx623, CLK=>nx1498, R=>nx1472);
   ix624 : mux21_ni port map ( Y=>nx623, A0=>q_3_4_EXMPLR, A1=>q_2_4_EXMPLR, 
      S0=>nx1446);
   gen_regs_2_regi_reg_q_4 : dffr port map ( Q=>q_2_4_EXMPLR, QB=>OPEN, D=>
      nx613, CLK=>nx1498, R=>nx1472);
   ix614 : mux21_ni port map ( Y=>nx613, A0=>q_2_4_EXMPLR, A1=>q_1_4_EXMPLR, 
      S0=>nx1446);
   gen_regs_1_regi_reg_q_4 : dffr port map ( Q=>q_1_4_EXMPLR, QB=>OPEN, D=>
      nx603, CLK=>nx1498, R=>nx1472);
   ix604 : mux21_ni port map ( Y=>nx603, A0=>q_1_4_EXMPLR, A1=>q_0_4_EXMPLR, 
      S0=>nx1446);
   reg0_reg_q_4 : dffr port map ( Q=>q_0_4_EXMPLR, QB=>OPEN, D=>nx593, CLK=>
      nx1496, R=>nx1470);
   ix594 : mux21_ni port map ( Y=>nx593, A0=>q_0_4_EXMPLR, A1=>d(4), S0=>
      nx1444);
   gen_regs_4_regi_reg_q_5 : dffr port map ( Q=>q_4_5_EXMPLR, QB=>OPEN, D=>
      nx683, CLK=>nx1500, R=>nx1474);
   ix684 : mux21_ni port map ( Y=>nx683, A0=>q_4_5_EXMPLR, A1=>q_3_5_EXMPLR, 
      S0=>nx1448);
   gen_regs_3_regi_reg_q_5 : dffr port map ( Q=>q_3_5_EXMPLR, QB=>OPEN, D=>
      nx673, CLK=>nx1500, R=>nx1474);
   ix674 : mux21_ni port map ( Y=>nx673, A0=>q_3_5_EXMPLR, A1=>q_2_5_EXMPLR, 
      S0=>nx1448);
   gen_regs_2_regi_reg_q_5 : dffr port map ( Q=>q_2_5_EXMPLR, QB=>OPEN, D=>
      nx663, CLK=>nx1498, R=>nx1472);
   ix664 : mux21_ni port map ( Y=>nx663, A0=>q_2_5_EXMPLR, A1=>q_1_5_EXMPLR, 
      S0=>nx1446);
   gen_regs_1_regi_reg_q_5 : dffr port map ( Q=>q_1_5_EXMPLR, QB=>OPEN, D=>
      nx653, CLK=>nx1498, R=>nx1472);
   ix654 : mux21_ni port map ( Y=>nx653, A0=>q_1_5_EXMPLR, A1=>q_0_5_EXMPLR, 
      S0=>nx1446);
   reg0_reg_q_5 : dffr port map ( Q=>q_0_5_EXMPLR, QB=>OPEN, D=>nx643, CLK=>
      nx1498, R=>nx1472);
   ix644 : mux21_ni port map ( Y=>nx643, A0=>q_0_5_EXMPLR, A1=>d(5), S0=>
      nx1446);
   gen_regs_4_regi_reg_q_6 : dffr port map ( Q=>q_4_6_EXMPLR, QB=>OPEN, D=>
      nx733, CLK=>nx1500, R=>nx1474);
   ix734 : mux21_ni port map ( Y=>nx733, A0=>q_4_6_EXMPLR, A1=>q_3_6_EXMPLR, 
      S0=>nx1448);
   gen_regs_3_regi_reg_q_6 : dffr port map ( Q=>q_3_6_EXMPLR, QB=>OPEN, D=>
      nx723, CLK=>nx1500, R=>nx1474);
   ix724 : mux21_ni port map ( Y=>nx723, A0=>q_3_6_EXMPLR, A1=>q_2_6_EXMPLR, 
      S0=>nx1448);
   gen_regs_2_regi_reg_q_6 : dffr port map ( Q=>q_2_6_EXMPLR, QB=>OPEN, D=>
      nx713, CLK=>nx1500, R=>nx1474);
   ix714 : mux21_ni port map ( Y=>nx713, A0=>q_2_6_EXMPLR, A1=>q_1_6_EXMPLR, 
      S0=>nx1448);
   gen_regs_1_regi_reg_q_6 : dffr port map ( Q=>q_1_6_EXMPLR, QB=>OPEN, D=>
      nx703, CLK=>nx1500, R=>nx1474);
   ix704 : mux21_ni port map ( Y=>nx703, A0=>q_1_6_EXMPLR, A1=>q_0_6_EXMPLR, 
      S0=>nx1448);
   reg0_reg_q_6 : dffr port map ( Q=>q_0_6_EXMPLR, QB=>OPEN, D=>nx693, CLK=>
      nx1500, R=>nx1474);
   ix694 : mux21_ni port map ( Y=>nx693, A0=>q_0_6_EXMPLR, A1=>d(6), S0=>
      nx1448);
   gen_regs_4_regi_reg_q_7 : dffr port map ( Q=>q_4_7_EXMPLR, QB=>OPEN, D=>
      nx783, CLK=>nx1502, R=>nx1476);
   ix784 : mux21_ni port map ( Y=>nx783, A0=>q_4_7_EXMPLR, A1=>q_3_7_EXMPLR, 
      S0=>nx1450);
   gen_regs_3_regi_reg_q_7 : dffr port map ( Q=>q_3_7_EXMPLR, QB=>OPEN, D=>
      nx773, CLK=>nx1502, R=>nx1476);
   ix774 : mux21_ni port map ( Y=>nx773, A0=>q_3_7_EXMPLR, A1=>q_2_7_EXMPLR, 
      S0=>nx1450);
   gen_regs_2_regi_reg_q_7 : dffr port map ( Q=>q_2_7_EXMPLR, QB=>OPEN, D=>
      nx763, CLK=>nx1502, R=>nx1476);
   ix764 : mux21_ni port map ( Y=>nx763, A0=>q_2_7_EXMPLR, A1=>q_1_7_EXMPLR, 
      S0=>nx1450);
   gen_regs_1_regi_reg_q_7 : dffr port map ( Q=>q_1_7_EXMPLR, QB=>OPEN, D=>
      nx753, CLK=>nx1502, R=>nx1476);
   ix754 : mux21_ni port map ( Y=>nx753, A0=>q_1_7_EXMPLR, A1=>q_0_7_EXMPLR, 
      S0=>nx1450);
   reg0_reg_q_7 : dffr port map ( Q=>q_0_7_EXMPLR, QB=>OPEN, D=>nx743, CLK=>
      nx1502, R=>nx1476);
   ix744 : mux21_ni port map ( Y=>nx743, A0=>q_0_7_EXMPLR, A1=>d(7), S0=>
      nx1450);
   gen_regs_4_regi_reg_q_8 : dffr port map ( Q=>q_4_8_EXMPLR, QB=>OPEN, D=>
      nx833, CLK=>nx1504, R=>nx1478);
   ix834 : mux21_ni port map ( Y=>nx833, A0=>q_4_8_EXMPLR, A1=>q_3_8_EXMPLR, 
      S0=>nx1452);
   gen_regs_3_regi_reg_q_8 : dffr port map ( Q=>q_3_8_EXMPLR, QB=>OPEN, D=>
      nx823, CLK=>nx1504, R=>nx1478);
   ix824 : mux21_ni port map ( Y=>nx823, A0=>q_3_8_EXMPLR, A1=>q_2_8_EXMPLR, 
      S0=>nx1452);
   gen_regs_2_regi_reg_q_8 : dffr port map ( Q=>q_2_8_EXMPLR, QB=>OPEN, D=>
      nx813, CLK=>nx1504, R=>nx1478);
   ix814 : mux21_ni port map ( Y=>nx813, A0=>q_2_8_EXMPLR, A1=>q_1_8_EXMPLR, 
      S0=>nx1452);
   gen_regs_1_regi_reg_q_8 : dffr port map ( Q=>q_1_8_EXMPLR, QB=>OPEN, D=>
      nx803, CLK=>nx1502, R=>nx1476);
   ix804 : mux21_ni port map ( Y=>nx803, A0=>q_1_8_EXMPLR, A1=>q_0_8_EXMPLR, 
      S0=>nx1450);
   reg0_reg_q_8 : dffr port map ( Q=>q_0_8_EXMPLR, QB=>OPEN, D=>nx793, CLK=>
      nx1502, R=>nx1476);
   ix794 : mux21_ni port map ( Y=>nx793, A0=>q_0_8_EXMPLR, A1=>d(8), S0=>
      nx1450);
   gen_regs_4_regi_reg_q_9 : dffr port map ( Q=>q_4_9_EXMPLR, QB=>OPEN, D=>
      nx883, CLK=>nx1506, R=>nx1480);
   ix884 : mux21_ni port map ( Y=>nx883, A0=>q_4_9_EXMPLR, A1=>q_3_9_EXMPLR, 
      S0=>nx1454);
   gen_regs_3_regi_reg_q_9 : dffr port map ( Q=>q_3_9_EXMPLR, QB=>OPEN, D=>
      nx873, CLK=>nx1504, R=>nx1478);
   ix874 : mux21_ni port map ( Y=>nx873, A0=>q_3_9_EXMPLR, A1=>q_2_9_EXMPLR, 
      S0=>nx1452);
   gen_regs_2_regi_reg_q_9 : dffr port map ( Q=>q_2_9_EXMPLR, QB=>OPEN, D=>
      nx863, CLK=>nx1504, R=>nx1478);
   ix864 : mux21_ni port map ( Y=>nx863, A0=>q_2_9_EXMPLR, A1=>q_1_9_EXMPLR, 
      S0=>nx1452);
   gen_regs_1_regi_reg_q_9 : dffr port map ( Q=>q_1_9_EXMPLR, QB=>OPEN, D=>
      nx853, CLK=>nx1504, R=>nx1478);
   ix854 : mux21_ni port map ( Y=>nx853, A0=>q_1_9_EXMPLR, A1=>q_0_9_EXMPLR, 
      S0=>nx1452);
   reg0_reg_q_9 : dffr port map ( Q=>q_0_9_EXMPLR, QB=>OPEN, D=>nx843, CLK=>
      nx1504, R=>nx1478);
   ix844 : mux21_ni port map ( Y=>nx843, A0=>q_0_9_EXMPLR, A1=>d(9), S0=>
      nx1452);
   gen_regs_4_regi_reg_q_10 : dffr port map ( Q=>q_4_10_EXMPLR, QB=>OPEN, D
      =>nx933, CLK=>nx1506, R=>nx1480);
   ix934 : mux21_ni port map ( Y=>nx933, A0=>q_4_10_EXMPLR, A1=>
      q_3_10_EXMPLR, S0=>nx1454);
   gen_regs_3_regi_reg_q_10 : dffr port map ( Q=>q_3_10_EXMPLR, QB=>OPEN, D
      =>nx923, CLK=>nx1506, R=>nx1480);
   ix924 : mux21_ni port map ( Y=>nx923, A0=>q_3_10_EXMPLR, A1=>
      q_2_10_EXMPLR, S0=>nx1454);
   gen_regs_2_regi_reg_q_10 : dffr port map ( Q=>q_2_10_EXMPLR, QB=>OPEN, D
      =>nx913, CLK=>nx1506, R=>nx1480);
   ix914 : mux21_ni port map ( Y=>nx913, A0=>q_2_10_EXMPLR, A1=>
      q_1_10_EXMPLR, S0=>nx1454);
   gen_regs_1_regi_reg_q_10 : dffr port map ( Q=>q_1_10_EXMPLR, QB=>OPEN, D
      =>nx903, CLK=>nx1506, R=>nx1480);
   ix904 : mux21_ni port map ( Y=>nx903, A0=>q_1_10_EXMPLR, A1=>
      q_0_10_EXMPLR, S0=>nx1454);
   reg0_reg_q_10 : dffr port map ( Q=>q_0_10_EXMPLR, QB=>OPEN, D=>nx893, CLK
      =>nx1506, R=>nx1480);
   ix894 : mux21_ni port map ( Y=>nx893, A0=>q_0_10_EXMPLR, A1=>d(10), S0=>
      nx1454);
   gen_regs_4_regi_reg_q_11 : dffr port map ( Q=>q_4_11_EXMPLR, QB=>OPEN, D
      =>nx983, CLK=>nx1508, R=>nx1482);
   ix984 : mux21_ni port map ( Y=>nx983, A0=>q_4_11_EXMPLR, A1=>
      q_3_11_EXMPLR, S0=>nx1456);
   gen_regs_3_regi_reg_q_11 : dffr port map ( Q=>q_3_11_EXMPLR, QB=>OPEN, D
      =>nx973, CLK=>nx1508, R=>nx1482);
   ix974 : mux21_ni port map ( Y=>nx973, A0=>q_3_11_EXMPLR, A1=>
      q_2_11_EXMPLR, S0=>nx1456);
   gen_regs_2_regi_reg_q_11 : dffr port map ( Q=>q_2_11_EXMPLR, QB=>OPEN, D
      =>nx963, CLK=>nx1508, R=>nx1482);
   ix964 : mux21_ni port map ( Y=>nx963, A0=>q_2_11_EXMPLR, A1=>
      q_1_11_EXMPLR, S0=>nx1456);
   gen_regs_1_regi_reg_q_11 : dffr port map ( Q=>q_1_11_EXMPLR, QB=>OPEN, D
      =>nx953, CLK=>nx1508, R=>nx1482);
   ix954 : mux21_ni port map ( Y=>nx953, A0=>q_1_11_EXMPLR, A1=>
      q_0_11_EXMPLR, S0=>nx1456);
   reg0_reg_q_11 : dffr port map ( Q=>q_0_11_EXMPLR, QB=>OPEN, D=>nx943, CLK
      =>nx1506, R=>nx1480);
   ix944 : mux21_ni port map ( Y=>nx943, A0=>q_0_11_EXMPLR, A1=>d(11), S0=>
      nx1454);
   gen_regs_4_regi_reg_q_12 : dffr port map ( Q=>q_4_12_EXMPLR, QB=>OPEN, D
      =>nx1033, CLK=>nx1510, R=>nx1484);
   ix1034 : mux21_ni port map ( Y=>nx1033, A0=>q_4_12_EXMPLR, A1=>
      q_3_12_EXMPLR, S0=>nx1458);
   gen_regs_3_regi_reg_q_12 : dffr port map ( Q=>q_3_12_EXMPLR, QB=>OPEN, D
      =>nx1023, CLK=>nx1510, R=>nx1484);
   ix1024 : mux21_ni port map ( Y=>nx1023, A0=>q_3_12_EXMPLR, A1=>
      q_2_12_EXMPLR, S0=>nx1458);
   gen_regs_2_regi_reg_q_12 : dffr port map ( Q=>q_2_12_EXMPLR, QB=>OPEN, D
      =>nx1013, CLK=>nx1508, R=>nx1482);
   ix1014 : mux21_ni port map ( Y=>nx1013, A0=>q_2_12_EXMPLR, A1=>
      q_1_12_EXMPLR, S0=>nx1456);
   gen_regs_1_regi_reg_q_12 : dffr port map ( Q=>q_1_12_EXMPLR, QB=>OPEN, D
      =>nx1003, CLK=>nx1508, R=>nx1482);
   ix1004 : mux21_ni port map ( Y=>nx1003, A0=>q_1_12_EXMPLR, A1=>
      q_0_12_EXMPLR, S0=>nx1456);
   reg0_reg_q_12 : dffr port map ( Q=>q_0_12_EXMPLR, QB=>OPEN, D=>nx993, CLK
      =>nx1508, R=>nx1482);
   ix994 : mux21_ni port map ( Y=>nx993, A0=>q_0_12_EXMPLR, A1=>d(12), S0=>
      nx1456);
   gen_regs_4_regi_reg_q_13 : dffr port map ( Q=>q_4_13_EXMPLR, QB=>OPEN, D
      =>nx1083, CLK=>nx1510, R=>nx1484);
   ix1084 : mux21_ni port map ( Y=>nx1083, A0=>q_4_13_EXMPLR, A1=>
      q_3_13_EXMPLR, S0=>nx1458);
   gen_regs_3_regi_reg_q_13 : dffr port map ( Q=>q_3_13_EXMPLR, QB=>OPEN, D
      =>nx1073, CLK=>nx1510, R=>nx1484);
   ix1074 : mux21_ni port map ( Y=>nx1073, A0=>q_3_13_EXMPLR, A1=>
      q_2_13_EXMPLR, S0=>nx1458);
   gen_regs_2_regi_reg_q_13 : dffr port map ( Q=>q_2_13_EXMPLR, QB=>OPEN, D
      =>nx1063, CLK=>nx1510, R=>nx1484);
   ix1064 : mux21_ni port map ( Y=>nx1063, A0=>q_2_13_EXMPLR, A1=>
      q_1_13_EXMPLR, S0=>nx1458);
   gen_regs_1_regi_reg_q_13 : dffr port map ( Q=>q_1_13_EXMPLR, QB=>OPEN, D
      =>nx1053, CLK=>nx1510, R=>nx1484);
   ix1054 : mux21_ni port map ( Y=>nx1053, A0=>q_1_13_EXMPLR, A1=>
      q_0_13_EXMPLR, S0=>nx1458);
   reg0_reg_q_13 : dffr port map ( Q=>q_0_13_EXMPLR, QB=>OPEN, D=>nx1043, 
      CLK=>nx1510, R=>nx1484);
   ix1044 : mux21_ni port map ( Y=>nx1043, A0=>q_0_13_EXMPLR, A1=>d(13), S0
      =>nx1458);
   gen_regs_4_regi_reg_q_14 : dffr port map ( Q=>q_4_14_EXMPLR, QB=>OPEN, D
      =>nx1133, CLK=>nx1512, R=>nx1486);
   ix1134 : mux21_ni port map ( Y=>nx1133, A0=>q_4_14_EXMPLR, A1=>
      q_3_14_EXMPLR, S0=>nx1460);
   gen_regs_3_regi_reg_q_14 : dffr port map ( Q=>q_3_14_EXMPLR, QB=>OPEN, D
      =>nx1123, CLK=>nx1512, R=>nx1486);
   ix1124 : mux21_ni port map ( Y=>nx1123, A0=>q_3_14_EXMPLR, A1=>
      q_2_14_EXMPLR, S0=>nx1460);
   gen_regs_2_regi_reg_q_14 : dffr port map ( Q=>q_2_14_EXMPLR, QB=>OPEN, D
      =>nx1113, CLK=>nx1512, R=>nx1486);
   ix1114 : mux21_ni port map ( Y=>nx1113, A0=>q_2_14_EXMPLR, A1=>
      q_1_14_EXMPLR, S0=>nx1460);
   gen_regs_1_regi_reg_q_14 : dffr port map ( Q=>q_1_14_EXMPLR, QB=>OPEN, D
      =>nx1103, CLK=>nx1512, R=>nx1486);
   ix1104 : mux21_ni port map ( Y=>nx1103, A0=>q_1_14_EXMPLR, A1=>
      q_0_14_EXMPLR, S0=>nx1460);
   reg0_reg_q_14 : dffr port map ( Q=>q_0_14_EXMPLR, QB=>OPEN, D=>nx1093, 
      CLK=>nx1512, R=>nx1486);
   ix1094 : mux21_ni port map ( Y=>nx1093, A0=>q_0_14_EXMPLR, A1=>d(14), S0
      =>nx1460);
   gen_regs_4_regi_reg_q_15 : dffr port map ( Q=>q_4_15_EXMPLR, QB=>OPEN, D
      =>nx1183, CLK=>nx1514, R=>nx1488);
   ix1184 : mux21_ni port map ( Y=>nx1183, A0=>q_4_15_EXMPLR, A1=>
      q_3_15_EXMPLR, S0=>nx1462);
   gen_regs_3_regi_reg_q_15 : dffr port map ( Q=>q_3_15_EXMPLR, QB=>OPEN, D
      =>nx1173, CLK=>nx1514, R=>nx1488);
   ix1174 : mux21_ni port map ( Y=>nx1173, A0=>q_3_15_EXMPLR, A1=>
      q_2_15_EXMPLR, S0=>nx1462);
   gen_regs_2_regi_reg_q_15 : dffr port map ( Q=>q_2_15_EXMPLR, QB=>OPEN, D
      =>nx1163, CLK=>nx1514, R=>nx1488);
   ix1164 : mux21_ni port map ( Y=>nx1163, A0=>q_2_15_EXMPLR, A1=>
      q_1_15_EXMPLR, S0=>nx1462);
   gen_regs_1_regi_reg_q_15 : dffr port map ( Q=>q_1_15_EXMPLR, QB=>OPEN, D
      =>nx1153, CLK=>nx1512, R=>nx1486);
   ix1154 : mux21_ni port map ( Y=>nx1153, A0=>q_1_15_EXMPLR, A1=>
      q_0_15_EXMPLR, S0=>nx1460);
   reg0_reg_q_15 : dffr port map ( Q=>q_0_15_EXMPLR, QB=>OPEN, D=>nx1143, 
      CLK=>nx1512, R=>nx1486);
   ix1144 : mux21_ni port map ( Y=>nx1143, A0=>q_0_15_EXMPLR, A1=>d(15), S0
      =>nx1460);
   ix1439 : inv02 port map ( Y=>nx1440, A=>nx1516);
   ix1441 : inv02 port map ( Y=>nx1442, A=>nx1516);
   ix1443 : inv02 port map ( Y=>nx1444, A=>nx1516);
   ix1445 : inv02 port map ( Y=>nx1446, A=>nx1516);
   ix1447 : inv02 port map ( Y=>nx1448, A=>nx1516);
   ix1449 : inv02 port map ( Y=>nx1450, A=>nx1516);
   ix1451 : inv02 port map ( Y=>nx1452, A=>nx1516);
   ix1453 : inv02 port map ( Y=>nx1454, A=>nx1518);
   ix1455 : inv02 port map ( Y=>nx1456, A=>nx1518);
   ix1457 : inv02 port map ( Y=>nx1458, A=>nx1518);
   ix1459 : inv02 port map ( Y=>nx1460, A=>nx1518);
   ix1461 : inv02 port map ( Y=>nx1462, A=>nx1518);
   ix1465 : inv02 port map ( Y=>nx1466, A=>nx1520);
   ix1467 : inv02 port map ( Y=>nx1468, A=>nx1520);
   ix1469 : inv02 port map ( Y=>nx1470, A=>nx1520);
   ix1471 : inv02 port map ( Y=>nx1472, A=>nx1520);
   ix1473 : inv02 port map ( Y=>nx1474, A=>nx1520);
   ix1475 : inv02 port map ( Y=>nx1476, A=>nx1520);
   ix1477 : inv02 port map ( Y=>nx1478, A=>nx1520);
   ix1479 : inv02 port map ( Y=>nx1480, A=>nx1522);
   ix1481 : inv02 port map ( Y=>nx1482, A=>nx1522);
   ix1483 : inv02 port map ( Y=>nx1484, A=>nx1522);
   ix1485 : inv02 port map ( Y=>nx1486, A=>nx1522);
   ix1487 : inv02 port map ( Y=>nx1488, A=>nx1522);
   ix1491 : inv02 port map ( Y=>nx1492, A=>nx1524);
   ix1493 : inv02 port map ( Y=>nx1494, A=>nx1524);
   ix1495 : inv02 port map ( Y=>nx1496, A=>nx1524);
   ix1497 : inv02 port map ( Y=>nx1498, A=>nx1524);
   ix1499 : inv02 port map ( Y=>nx1500, A=>nx1524);
   ix1501 : inv02 port map ( Y=>nx1502, A=>nx1524);
   ix1503 : inv02 port map ( Y=>nx1504, A=>nx1524);
   ix1505 : inv02 port map ( Y=>nx1506, A=>nx1526);
   ix1507 : inv02 port map ( Y=>nx1508, A=>nx1526);
   ix1509 : inv02 port map ( Y=>nx1510, A=>nx1526);
   ix1511 : inv02 port map ( Y=>nx1512, A=>nx1526);
   ix1513 : inv02 port map ( Y=>nx1514, A=>nx1526);
   ix1515 : inv02 port map ( Y=>nx1516, A=>load);
   ix1517 : inv02 port map ( Y=>nx1518, A=>load);
   ix1519 : inv02 port map ( Y=>nx1520, A=>reset);
   ix1521 : inv02 port map ( Y=>nx1522, A=>reset);
   ix1523 : inv02 port map ( Y=>nx1524, A=>clk);
   ix1525 : inv02 port map ( Y=>nx1526, A=>clk);
end Dataflow ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Cache_5_16_28_5 is
   port (
      in_word : IN std_logic_vector (15 DOWNTO 0) ;
      cache_in_sel : IN std_logic_vector (4 DOWNTO 0) ;
      cache_out_sel : IN std_logic_vector (4 DOWNTO 0) ;
      decoder_enable : IN std_logic ;
      out_column_0_15 : OUT std_logic ;
      out_column_0_14 : OUT std_logic ;
      out_column_0_13 : OUT std_logic ;
      out_column_0_12 : OUT std_logic ;
      out_column_0_11 : OUT std_logic ;
      out_column_0_10 : OUT std_logic ;
      out_column_0_9 : OUT std_logic ;
      out_column_0_8 : OUT std_logic ;
      out_column_0_7 : OUT std_logic ;
      out_column_0_6 : OUT std_logic ;
      out_column_0_5 : OUT std_logic ;
      out_column_0_4 : OUT std_logic ;
      out_column_0_3 : OUT std_logic ;
      out_column_0_2 : OUT std_logic ;
      out_column_0_1 : OUT std_logic ;
      out_column_0_0 : OUT std_logic ;
      out_column_1_15 : OUT std_logic ;
      out_column_1_14 : OUT std_logic ;
      out_column_1_13 : OUT std_logic ;
      out_column_1_12 : OUT std_logic ;
      out_column_1_11 : OUT std_logic ;
      out_column_1_10 : OUT std_logic ;
      out_column_1_9 : OUT std_logic ;
      out_column_1_8 : OUT std_logic ;
      out_column_1_7 : OUT std_logic ;
      out_column_1_6 : OUT std_logic ;
      out_column_1_5 : OUT std_logic ;
      out_column_1_4 : OUT std_logic ;
      out_column_1_3 : OUT std_logic ;
      out_column_1_2 : OUT std_logic ;
      out_column_1_1 : OUT std_logic ;
      out_column_1_0 : OUT std_logic ;
      out_column_2_15 : OUT std_logic ;
      out_column_2_14 : OUT std_logic ;
      out_column_2_13 : OUT std_logic ;
      out_column_2_12 : OUT std_logic ;
      out_column_2_11 : OUT std_logic ;
      out_column_2_10 : OUT std_logic ;
      out_column_2_9 : OUT std_logic ;
      out_column_2_8 : OUT std_logic ;
      out_column_2_7 : OUT std_logic ;
      out_column_2_6 : OUT std_logic ;
      out_column_2_5 : OUT std_logic ;
      out_column_2_4 : OUT std_logic ;
      out_column_2_3 : OUT std_logic ;
      out_column_2_2 : OUT std_logic ;
      out_column_2_1 : OUT std_logic ;
      out_column_2_0 : OUT std_logic ;
      out_column_3_15 : OUT std_logic ;
      out_column_3_14 : OUT std_logic ;
      out_column_3_13 : OUT std_logic ;
      out_column_3_12 : OUT std_logic ;
      out_column_3_11 : OUT std_logic ;
      out_column_3_10 : OUT std_logic ;
      out_column_3_9 : OUT std_logic ;
      out_column_3_8 : OUT std_logic ;
      out_column_3_7 : OUT std_logic ;
      out_column_3_6 : OUT std_logic ;
      out_column_3_5 : OUT std_logic ;
      out_column_3_4 : OUT std_logic ;
      out_column_3_3 : OUT std_logic ;
      out_column_3_2 : OUT std_logic ;
      out_column_3_1 : OUT std_logic ;
      out_column_3_0 : OUT std_logic ;
      out_column_4_15 : OUT std_logic ;
      out_column_4_14 : OUT std_logic ;
      out_column_4_13 : OUT std_logic ;
      out_column_4_12 : OUT std_logic ;
      out_column_4_11 : OUT std_logic ;
      out_column_4_10 : OUT std_logic ;
      out_column_4_9 : OUT std_logic ;
      out_column_4_8 : OUT std_logic ;
      out_column_4_7 : OUT std_logic ;
      out_column_4_6 : OUT std_logic ;
      out_column_4_5 : OUT std_logic ;
      out_column_4_4 : OUT std_logic ;
      out_column_4_3 : OUT std_logic ;
      out_column_4_2 : OUT std_logic ;
      out_column_4_1 : OUT std_logic ;
      out_column_4_0 : OUT std_logic ;
      clk : IN std_logic ;
      reset : IN std_logic) ;
end Cache_5_16_28_5 ;

architecture Dataflow of Cache_5_16_28_5 is
   component Queue_5
      port (
         d : IN std_logic_vector (15 DOWNTO 0) ;
         q_0_15 : OUT std_logic ;
         q_0_14 : OUT std_logic ;
         q_0_13 : OUT std_logic ;
         q_0_12 : OUT std_logic ;
         q_0_11 : OUT std_logic ;
         q_0_10 : OUT std_logic ;
         q_0_9 : OUT std_logic ;
         q_0_8 : OUT std_logic ;
         q_0_7 : OUT std_logic ;
         q_0_6 : OUT std_logic ;
         q_0_5 : OUT std_logic ;
         q_0_4 : OUT std_logic ;
         q_0_3 : OUT std_logic ;
         q_0_2 : OUT std_logic ;
         q_0_1 : OUT std_logic ;
         q_0_0 : OUT std_logic ;
         q_1_15 : OUT std_logic ;
         q_1_14 : OUT std_logic ;
         q_1_13 : OUT std_logic ;
         q_1_12 : OUT std_logic ;
         q_1_11 : OUT std_logic ;
         q_1_10 : OUT std_logic ;
         q_1_9 : OUT std_logic ;
         q_1_8 : OUT std_logic ;
         q_1_7 : OUT std_logic ;
         q_1_6 : OUT std_logic ;
         q_1_5 : OUT std_logic ;
         q_1_4 : OUT std_logic ;
         q_1_3 : OUT std_logic ;
         q_1_2 : OUT std_logic ;
         q_1_1 : OUT std_logic ;
         q_1_0 : OUT std_logic ;
         q_2_15 : OUT std_logic ;
         q_2_14 : OUT std_logic ;
         q_2_13 : OUT std_logic ;
         q_2_12 : OUT std_logic ;
         q_2_11 : OUT std_logic ;
         q_2_10 : OUT std_logic ;
         q_2_9 : OUT std_logic ;
         q_2_8 : OUT std_logic ;
         q_2_7 : OUT std_logic ;
         q_2_6 : OUT std_logic ;
         q_2_5 : OUT std_logic ;
         q_2_4 : OUT std_logic ;
         q_2_3 : OUT std_logic ;
         q_2_2 : OUT std_logic ;
         q_2_1 : OUT std_logic ;
         q_2_0 : OUT std_logic ;
         q_3_15 : OUT std_logic ;
         q_3_14 : OUT std_logic ;
         q_3_13 : OUT std_logic ;
         q_3_12 : OUT std_logic ;
         q_3_11 : OUT std_logic ;
         q_3_10 : OUT std_logic ;
         q_3_9 : OUT std_logic ;
         q_3_8 : OUT std_logic ;
         q_3_7 : OUT std_logic ;
         q_3_6 : OUT std_logic ;
         q_3_5 : OUT std_logic ;
         q_3_4 : OUT std_logic ;
         q_3_3 : OUT std_logic ;
         q_3_2 : OUT std_logic ;
         q_3_1 : OUT std_logic ;
         q_3_0 : OUT std_logic ;
         q_4_15 : OUT std_logic ;
         q_4_14 : OUT std_logic ;
         q_4_13 : OUT std_logic ;
         q_4_12 : OUT std_logic ;
         q_4_11 : OUT std_logic ;
         q_4_10 : OUT std_logic ;
         q_4_9 : OUT std_logic ;
         q_4_8 : OUT std_logic ;
         q_4_7 : OUT std_logic ;
         q_4_6 : OUT std_logic ;
         q_4_5 : OUT std_logic ;
         q_4_4 : OUT std_logic ;
         q_4_3 : OUT std_logic ;
         q_4_2 : OUT std_logic ;
         q_4_1 : OUT std_logic ;
         q_4_0 : OUT std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         reset : IN std_logic) ;
   end component ;
   signal que_out_0_0_15, que_out_0_0_14, que_out_0_0_13, que_out_0_0_12, 
      que_out_0_0_11, que_out_0_0_10, que_out_0_0_9, que_out_0_0_8, 
      que_out_0_0_7, que_out_0_0_6, que_out_0_0_5, que_out_0_0_4, 
      que_out_0_0_3, que_out_0_0_2, que_out_0_0_1, que_out_0_0_0, 
      que_out_0_1_15, que_out_0_1_14, que_out_0_1_13, que_out_0_1_12, 
      que_out_0_1_11, que_out_0_1_10, que_out_0_1_9, que_out_0_1_8, 
      que_out_0_1_7, que_out_0_1_6, que_out_0_1_5, que_out_0_1_4, 
      que_out_0_1_3, que_out_0_1_2, que_out_0_1_1, que_out_0_1_0, 
      que_out_0_2_15, que_out_0_2_14, que_out_0_2_13, que_out_0_2_12, 
      que_out_0_2_11, que_out_0_2_10, que_out_0_2_9, que_out_0_2_8, 
      que_out_0_2_7, que_out_0_2_6, que_out_0_2_5, que_out_0_2_4, 
      que_out_0_2_3, que_out_0_2_2, que_out_0_2_1, que_out_0_2_0, 
      que_out_0_3_15, que_out_0_3_14, que_out_0_3_13, que_out_0_3_12, 
      que_out_0_3_11, que_out_0_3_10, que_out_0_3_9, que_out_0_3_8, 
      que_out_0_3_7, que_out_0_3_6, que_out_0_3_5, que_out_0_3_4, 
      que_out_0_3_3, que_out_0_3_2, que_out_0_3_1, que_out_0_3_0, 
      que_out_0_4_15, que_out_0_4_14, que_out_0_4_13, que_out_0_4_12, 
      que_out_0_4_11, que_out_0_4_10, que_out_0_4_9, que_out_0_4_8, 
      que_out_0_4_7, que_out_0_4_6, que_out_0_4_5, que_out_0_4_4, 
      que_out_0_4_3, que_out_0_4_2, que_out_0_4_1, que_out_0_4_0, 
      que_out_1_0_15, que_out_1_0_14, que_out_1_0_13, que_out_1_0_12, 
      que_out_1_0_11, que_out_1_0_10, que_out_1_0_9, que_out_1_0_8, 
      que_out_1_0_7, que_out_1_0_6, que_out_1_0_5, que_out_1_0_4, 
      que_out_1_0_3, que_out_1_0_2, que_out_1_0_1, que_out_1_0_0, 
      que_out_1_1_15, que_out_1_1_14, que_out_1_1_13, que_out_1_1_12, 
      que_out_1_1_11, que_out_1_1_10, que_out_1_1_9, que_out_1_1_8, 
      que_out_1_1_7, que_out_1_1_6, que_out_1_1_5, que_out_1_1_4, 
      que_out_1_1_3, que_out_1_1_2, que_out_1_1_1, que_out_1_1_0, 
      que_out_1_2_15, que_out_1_2_14, que_out_1_2_13, que_out_1_2_12, 
      que_out_1_2_11, que_out_1_2_10, que_out_1_2_9, que_out_1_2_8, 
      que_out_1_2_7, que_out_1_2_6, que_out_1_2_5, que_out_1_2_4, 
      que_out_1_2_3, que_out_1_2_2, que_out_1_2_1, que_out_1_2_0, 
      que_out_1_3_15, que_out_1_3_14, que_out_1_3_13, que_out_1_3_12, 
      que_out_1_3_11, que_out_1_3_10, que_out_1_3_9, que_out_1_3_8, 
      que_out_1_3_7, que_out_1_3_6, que_out_1_3_5, que_out_1_3_4, 
      que_out_1_3_3, que_out_1_3_2, que_out_1_3_1, que_out_1_3_0, 
      que_out_1_4_15, que_out_1_4_14, que_out_1_4_13, que_out_1_4_12, 
      que_out_1_4_11, que_out_1_4_10, que_out_1_4_9, que_out_1_4_8, 
      que_out_1_4_7, que_out_1_4_6, que_out_1_4_5, que_out_1_4_4, 
      que_out_1_4_3, que_out_1_4_2, que_out_1_4_1, que_out_1_4_0, 
      que_out_2_0_15, que_out_2_0_14, que_out_2_0_13, que_out_2_0_12, 
      que_out_2_0_11, que_out_2_0_10, que_out_2_0_9, que_out_2_0_8, 
      que_out_2_0_7, que_out_2_0_6, que_out_2_0_5, que_out_2_0_4, 
      que_out_2_0_3, que_out_2_0_2, que_out_2_0_1, que_out_2_0_0, 
      que_out_2_1_15, que_out_2_1_14, que_out_2_1_13, que_out_2_1_12, 
      que_out_2_1_11, que_out_2_1_10, que_out_2_1_9, que_out_2_1_8, 
      que_out_2_1_7, que_out_2_1_6, que_out_2_1_5, que_out_2_1_4, 
      que_out_2_1_3, que_out_2_1_2, que_out_2_1_1, que_out_2_1_0, 
      que_out_2_2_15, que_out_2_2_14, que_out_2_2_13, que_out_2_2_12, 
      que_out_2_2_11, que_out_2_2_10, que_out_2_2_9, que_out_2_2_8, 
      que_out_2_2_7, que_out_2_2_6, que_out_2_2_5, que_out_2_2_4, 
      que_out_2_2_3, que_out_2_2_2, que_out_2_2_1, que_out_2_2_0, 
      que_out_2_3_15, que_out_2_3_14, que_out_2_3_13, que_out_2_3_12, 
      que_out_2_3_11, que_out_2_3_10, que_out_2_3_9, que_out_2_3_8, 
      que_out_2_3_7, que_out_2_3_6, que_out_2_3_5, que_out_2_3_4, 
      que_out_2_3_3, que_out_2_3_2, que_out_2_3_1, que_out_2_3_0, 
      que_out_2_4_15, que_out_2_4_14, que_out_2_4_13, que_out_2_4_12, 
      que_out_2_4_11, que_out_2_4_10, que_out_2_4_9, que_out_2_4_8, 
      que_out_2_4_7, que_out_2_4_6, que_out_2_4_5, que_out_2_4_4, 
      que_out_2_4_3, que_out_2_4_2, que_out_2_4_1, que_out_2_4_0, 
      que_out_3_0_15, que_out_3_0_14, que_out_3_0_13, que_out_3_0_12, 
      que_out_3_0_11, que_out_3_0_10, que_out_3_0_9, que_out_3_0_8, 
      que_out_3_0_7, que_out_3_0_6, que_out_3_0_5, que_out_3_0_4, 
      que_out_3_0_3, que_out_3_0_2, que_out_3_0_1, que_out_3_0_0, 
      que_out_3_1_15, que_out_3_1_14, que_out_3_1_13, que_out_3_1_12, 
      que_out_3_1_11, que_out_3_1_10, que_out_3_1_9, que_out_3_1_8, 
      que_out_3_1_7, que_out_3_1_6, que_out_3_1_5, que_out_3_1_4, 
      que_out_3_1_3, que_out_3_1_2, que_out_3_1_1, que_out_3_1_0, 
      que_out_3_2_15, que_out_3_2_14, que_out_3_2_13, que_out_3_2_12, 
      que_out_3_2_11, que_out_3_2_10, que_out_3_2_9, que_out_3_2_8, 
      que_out_3_2_7, que_out_3_2_6, que_out_3_2_5, que_out_3_2_4, 
      que_out_3_2_3, que_out_3_2_2, que_out_3_2_1, que_out_3_2_0, 
      que_out_3_3_15, que_out_3_3_14, que_out_3_3_13, que_out_3_3_12, 
      que_out_3_3_11, que_out_3_3_10, que_out_3_3_9, que_out_3_3_8, 
      que_out_3_3_7, que_out_3_3_6, que_out_3_3_5, que_out_3_3_4, 
      que_out_3_3_3, que_out_3_3_2, que_out_3_3_1, que_out_3_3_0, 
      que_out_3_4_15, que_out_3_4_14, que_out_3_4_13, que_out_3_4_12, 
      que_out_3_4_11, que_out_3_4_10, que_out_3_4_9, que_out_3_4_8, 
      que_out_3_4_7, que_out_3_4_6, que_out_3_4_5, que_out_3_4_4, 
      que_out_3_4_3, que_out_3_4_2, que_out_3_4_1, que_out_3_4_0, 
      que_out_4_0_15, que_out_4_0_14, que_out_4_0_13, que_out_4_0_12, 
      que_out_4_0_11, que_out_4_0_10, que_out_4_0_9, que_out_4_0_8, 
      que_out_4_0_7, que_out_4_0_6, que_out_4_0_5, que_out_4_0_4, 
      que_out_4_0_3, que_out_4_0_2, que_out_4_0_1, que_out_4_0_0, 
      que_out_4_1_15, que_out_4_1_14, que_out_4_1_13, que_out_4_1_12, 
      que_out_4_1_11, que_out_4_1_10, que_out_4_1_9, que_out_4_1_8, 
      que_out_4_1_7, que_out_4_1_6, que_out_4_1_5, que_out_4_1_4, 
      que_out_4_1_3, que_out_4_1_2, que_out_4_1_1, que_out_4_1_0, 
      que_out_4_2_15, que_out_4_2_14, que_out_4_2_13, que_out_4_2_12, 
      que_out_4_2_11, que_out_4_2_10, que_out_4_2_9, que_out_4_2_8, 
      que_out_4_2_7, que_out_4_2_6, que_out_4_2_5, que_out_4_2_4, 
      que_out_4_2_3, que_out_4_2_2, que_out_4_2_1, que_out_4_2_0, 
      que_out_4_3_15, que_out_4_3_14, que_out_4_3_13, que_out_4_3_12, 
      que_out_4_3_11, que_out_4_3_10, que_out_4_3_9, que_out_4_3_8, 
      que_out_4_3_7, que_out_4_3_6, que_out_4_3_5, que_out_4_3_4, 
      que_out_4_3_3, que_out_4_3_2, que_out_4_3_1, que_out_4_3_0, 
      que_out_4_4_15, que_out_4_4_14, que_out_4_4_13, que_out_4_4_12, 
      que_out_4_4_11, que_out_4_4_10, que_out_4_4_9, que_out_4_4_8, 
      que_out_4_4_7, que_out_4_4_6, que_out_4_4_5, que_out_4_4_4, 
      que_out_4_4_3, que_out_4_4_2, que_out_4_4_1, que_out_4_4_0, 
      que_out_5_0_15, que_out_5_0_14, que_out_5_0_13, que_out_5_0_12, 
      que_out_5_0_11, que_out_5_0_10, que_out_5_0_9, que_out_5_0_8, 
      que_out_5_0_7, que_out_5_0_6, que_out_5_0_5, que_out_5_0_4, 
      que_out_5_0_3, que_out_5_0_2, que_out_5_0_1, que_out_5_0_0, 
      que_out_5_1_15, que_out_5_1_14, que_out_5_1_13, que_out_5_1_12, 
      que_out_5_1_11, que_out_5_1_10, que_out_5_1_9, que_out_5_1_8, 
      que_out_5_1_7, que_out_5_1_6, que_out_5_1_5, que_out_5_1_4, 
      que_out_5_1_3, que_out_5_1_2, que_out_5_1_1, que_out_5_1_0, 
      que_out_5_2_15, que_out_5_2_14, que_out_5_2_13, que_out_5_2_12, 
      que_out_5_2_11, que_out_5_2_10, que_out_5_2_9, que_out_5_2_8, 
      que_out_5_2_7, que_out_5_2_6, que_out_5_2_5, que_out_5_2_4, 
      que_out_5_2_3, que_out_5_2_2, que_out_5_2_1, que_out_5_2_0, 
      que_out_5_3_15, que_out_5_3_14, que_out_5_3_13, que_out_5_3_12, 
      que_out_5_3_11, que_out_5_3_10, que_out_5_3_9, que_out_5_3_8, 
      que_out_5_3_7, que_out_5_3_6, que_out_5_3_5, que_out_5_3_4, 
      que_out_5_3_3, que_out_5_3_2, que_out_5_3_1, que_out_5_3_0, 
      que_out_5_4_15, que_out_5_4_14, que_out_5_4_13, que_out_5_4_12, 
      que_out_5_4_11, que_out_5_4_10, que_out_5_4_9, que_out_5_4_8, 
      que_out_5_4_7, que_out_5_4_6, que_out_5_4_5, que_out_5_4_4, 
      que_out_5_4_3, que_out_5_4_2, que_out_5_4_1, que_out_5_4_0, 
      que_out_6_0_15, que_out_6_0_14, que_out_6_0_13, que_out_6_0_12, 
      que_out_6_0_11, que_out_6_0_10, que_out_6_0_9, que_out_6_0_8, 
      que_out_6_0_7, que_out_6_0_6, que_out_6_0_5, que_out_6_0_4, 
      que_out_6_0_3, que_out_6_0_2, que_out_6_0_1, que_out_6_0_0, 
      que_out_6_1_15, que_out_6_1_14, que_out_6_1_13, que_out_6_1_12, 
      que_out_6_1_11, que_out_6_1_10, que_out_6_1_9, que_out_6_1_8, 
      que_out_6_1_7, que_out_6_1_6, que_out_6_1_5, que_out_6_1_4, 
      que_out_6_1_3, que_out_6_1_2, que_out_6_1_1, que_out_6_1_0, 
      que_out_6_2_15, que_out_6_2_14, que_out_6_2_13, que_out_6_2_12, 
      que_out_6_2_11, que_out_6_2_10, que_out_6_2_9, que_out_6_2_8, 
      que_out_6_2_7, que_out_6_2_6, que_out_6_2_5, que_out_6_2_4, 
      que_out_6_2_3, que_out_6_2_2, que_out_6_2_1, que_out_6_2_0, 
      que_out_6_3_15, que_out_6_3_14, que_out_6_3_13, que_out_6_3_12, 
      que_out_6_3_11, que_out_6_3_10, que_out_6_3_9, que_out_6_3_8, 
      que_out_6_3_7, que_out_6_3_6, que_out_6_3_5, que_out_6_3_4, 
      que_out_6_3_3, que_out_6_3_2, que_out_6_3_1, que_out_6_3_0, 
      que_out_6_4_15, que_out_6_4_14, que_out_6_4_13, que_out_6_4_12, 
      que_out_6_4_11, que_out_6_4_10, que_out_6_4_9, que_out_6_4_8, 
      que_out_6_4_7, que_out_6_4_6, que_out_6_4_5, que_out_6_4_4, 
      que_out_6_4_3, que_out_6_4_2, que_out_6_4_1, que_out_6_4_0, 
      que_out_7_0_15, que_out_7_0_14, que_out_7_0_13, que_out_7_0_12, 
      que_out_7_0_11, que_out_7_0_10, que_out_7_0_9, que_out_7_0_8, 
      que_out_7_0_7, que_out_7_0_6, que_out_7_0_5, que_out_7_0_4, 
      que_out_7_0_3, que_out_7_0_2, que_out_7_0_1, que_out_7_0_0, 
      que_out_7_1_15, que_out_7_1_14, que_out_7_1_13, que_out_7_1_12, 
      que_out_7_1_11, que_out_7_1_10, que_out_7_1_9, que_out_7_1_8, 
      que_out_7_1_7, que_out_7_1_6, que_out_7_1_5, que_out_7_1_4, 
      que_out_7_1_3, que_out_7_1_2, que_out_7_1_1, que_out_7_1_0, 
      que_out_7_2_15, que_out_7_2_14, que_out_7_2_13, que_out_7_2_12, 
      que_out_7_2_11, que_out_7_2_10, que_out_7_2_9, que_out_7_2_8, 
      que_out_7_2_7, que_out_7_2_6, que_out_7_2_5, que_out_7_2_4, 
      que_out_7_2_3, que_out_7_2_2, que_out_7_2_1, que_out_7_2_0, 
      que_out_7_3_15, que_out_7_3_14, que_out_7_3_13, que_out_7_3_12, 
      que_out_7_3_11, que_out_7_3_10, que_out_7_3_9, que_out_7_3_8, 
      que_out_7_3_7, que_out_7_3_6, que_out_7_3_5, que_out_7_3_4, 
      que_out_7_3_3, que_out_7_3_2, que_out_7_3_1, que_out_7_3_0, 
      que_out_7_4_15, que_out_7_4_14, que_out_7_4_13, que_out_7_4_12, 
      que_out_7_4_11, que_out_7_4_10, que_out_7_4_9, que_out_7_4_8, 
      que_out_7_4_7, que_out_7_4_6, que_out_7_4_5, que_out_7_4_4, 
      que_out_7_4_3, que_out_7_4_2, que_out_7_4_1, que_out_7_4_0, 
      que_out_8_0_15, que_out_8_0_14, que_out_8_0_13, que_out_8_0_12, 
      que_out_8_0_11, que_out_8_0_10, que_out_8_0_9, que_out_8_0_8, 
      que_out_8_0_7, que_out_8_0_6, que_out_8_0_5, que_out_8_0_4, 
      que_out_8_0_3, que_out_8_0_2, que_out_8_0_1, que_out_8_0_0, 
      que_out_8_1_15, que_out_8_1_14, que_out_8_1_13, que_out_8_1_12, 
      que_out_8_1_11, que_out_8_1_10, que_out_8_1_9, que_out_8_1_8, 
      que_out_8_1_7, que_out_8_1_6, que_out_8_1_5, que_out_8_1_4, 
      que_out_8_1_3, que_out_8_1_2, que_out_8_1_1, que_out_8_1_0, 
      que_out_8_2_15, que_out_8_2_14, que_out_8_2_13, que_out_8_2_12, 
      que_out_8_2_11, que_out_8_2_10, que_out_8_2_9, que_out_8_2_8, 
      que_out_8_2_7, que_out_8_2_6, que_out_8_2_5, que_out_8_2_4, 
      que_out_8_2_3, que_out_8_2_2, que_out_8_2_1, que_out_8_2_0, 
      que_out_8_3_15, que_out_8_3_14, que_out_8_3_13, que_out_8_3_12, 
      que_out_8_3_11, que_out_8_3_10, que_out_8_3_9, que_out_8_3_8, 
      que_out_8_3_7, que_out_8_3_6, que_out_8_3_5, que_out_8_3_4, 
      que_out_8_3_3, que_out_8_3_2, que_out_8_3_1, que_out_8_3_0, 
      que_out_8_4_15, que_out_8_4_14, que_out_8_4_13, que_out_8_4_12, 
      que_out_8_4_11, que_out_8_4_10, que_out_8_4_9, que_out_8_4_8, 
      que_out_8_4_7, que_out_8_4_6, que_out_8_4_5, que_out_8_4_4, 
      que_out_8_4_3, que_out_8_4_2, que_out_8_4_1, que_out_8_4_0, 
      que_out_9_0_15, que_out_9_0_14, que_out_9_0_13, que_out_9_0_12, 
      que_out_9_0_11, que_out_9_0_10, que_out_9_0_9, que_out_9_0_8, 
      que_out_9_0_7, que_out_9_0_6, que_out_9_0_5, que_out_9_0_4, 
      que_out_9_0_3, que_out_9_0_2, que_out_9_0_1, que_out_9_0_0, 
      que_out_9_1_15, que_out_9_1_14, que_out_9_1_13, que_out_9_1_12, 
      que_out_9_1_11, que_out_9_1_10, que_out_9_1_9, que_out_9_1_8, 
      que_out_9_1_7, que_out_9_1_6, que_out_9_1_5, que_out_9_1_4, 
      que_out_9_1_3, que_out_9_1_2, que_out_9_1_1, que_out_9_1_0, 
      que_out_9_2_15, que_out_9_2_14, que_out_9_2_13, que_out_9_2_12, 
      que_out_9_2_11, que_out_9_2_10, que_out_9_2_9, que_out_9_2_8, 
      que_out_9_2_7, que_out_9_2_6, que_out_9_2_5, que_out_9_2_4, 
      que_out_9_2_3, que_out_9_2_2, que_out_9_2_1, que_out_9_2_0, 
      que_out_9_3_15, que_out_9_3_14, que_out_9_3_13, que_out_9_3_12, 
      que_out_9_3_11, que_out_9_3_10, que_out_9_3_9, que_out_9_3_8, 
      que_out_9_3_7, que_out_9_3_6, que_out_9_3_5, que_out_9_3_4, 
      que_out_9_3_3, que_out_9_3_2, que_out_9_3_1, que_out_9_3_0, 
      que_out_9_4_15, que_out_9_4_14, que_out_9_4_13, que_out_9_4_12, 
      que_out_9_4_11, que_out_9_4_10, que_out_9_4_9, que_out_9_4_8, 
      que_out_9_4_7, que_out_9_4_6, que_out_9_4_5, que_out_9_4_4, 
      que_out_9_4_3, que_out_9_4_2, que_out_9_4_1, que_out_9_4_0, 
      que_out_10_0_15, que_out_10_0_14, que_out_10_0_13, que_out_10_0_12, 
      que_out_10_0_11, que_out_10_0_10, que_out_10_0_9, que_out_10_0_8, 
      que_out_10_0_7, que_out_10_0_6, que_out_10_0_5, que_out_10_0_4, 
      que_out_10_0_3, que_out_10_0_2, que_out_10_0_1, que_out_10_0_0, 
      que_out_10_1_15, que_out_10_1_14, que_out_10_1_13, que_out_10_1_12, 
      que_out_10_1_11, que_out_10_1_10, que_out_10_1_9, que_out_10_1_8, 
      que_out_10_1_7, que_out_10_1_6, que_out_10_1_5, que_out_10_1_4, 
      que_out_10_1_3, que_out_10_1_2, que_out_10_1_1, que_out_10_1_0, 
      que_out_10_2_15, que_out_10_2_14, que_out_10_2_13, que_out_10_2_12, 
      que_out_10_2_11, que_out_10_2_10, que_out_10_2_9, que_out_10_2_8, 
      que_out_10_2_7, que_out_10_2_6, que_out_10_2_5, que_out_10_2_4, 
      que_out_10_2_3, que_out_10_2_2, que_out_10_2_1, que_out_10_2_0, 
      que_out_10_3_15, que_out_10_3_14, que_out_10_3_13, que_out_10_3_12, 
      que_out_10_3_11, que_out_10_3_10, que_out_10_3_9, que_out_10_3_8, 
      que_out_10_3_7, que_out_10_3_6, que_out_10_3_5, que_out_10_3_4, 
      que_out_10_3_3, que_out_10_3_2, que_out_10_3_1, que_out_10_3_0, 
      que_out_10_4_15, que_out_10_4_14, que_out_10_4_13, que_out_10_4_12, 
      que_out_10_4_11, que_out_10_4_10, que_out_10_4_9, que_out_10_4_8, 
      que_out_10_4_7, que_out_10_4_6, que_out_10_4_5, que_out_10_4_4, 
      que_out_10_4_3, que_out_10_4_2, que_out_10_4_1, que_out_10_4_0, 
      que_out_11_0_15, que_out_11_0_14, que_out_11_0_13, que_out_11_0_12, 
      que_out_11_0_11, que_out_11_0_10, que_out_11_0_9, que_out_11_0_8, 
      que_out_11_0_7, que_out_11_0_6, que_out_11_0_5, que_out_11_0_4, 
      que_out_11_0_3, que_out_11_0_2, que_out_11_0_1, que_out_11_0_0, 
      que_out_11_1_15, que_out_11_1_14, que_out_11_1_13, que_out_11_1_12, 
      que_out_11_1_11, que_out_11_1_10, que_out_11_1_9, que_out_11_1_8, 
      que_out_11_1_7, que_out_11_1_6, que_out_11_1_5, que_out_11_1_4, 
      que_out_11_1_3, que_out_11_1_2, que_out_11_1_1, que_out_11_1_0, 
      que_out_11_2_15, que_out_11_2_14, que_out_11_2_13, que_out_11_2_12, 
      que_out_11_2_11, que_out_11_2_10, que_out_11_2_9, que_out_11_2_8, 
      que_out_11_2_7, que_out_11_2_6, que_out_11_2_5, que_out_11_2_4, 
      que_out_11_2_3, que_out_11_2_2, que_out_11_2_1, que_out_11_2_0, 
      que_out_11_3_15, que_out_11_3_14, que_out_11_3_13, que_out_11_3_12, 
      que_out_11_3_11, que_out_11_3_10, que_out_11_3_9, que_out_11_3_8, 
      que_out_11_3_7, que_out_11_3_6, que_out_11_3_5, que_out_11_3_4, 
      que_out_11_3_3, que_out_11_3_2, que_out_11_3_1, que_out_11_3_0, 
      que_out_11_4_15, que_out_11_4_14, que_out_11_4_13, que_out_11_4_12, 
      que_out_11_4_11, que_out_11_4_10, que_out_11_4_9, que_out_11_4_8, 
      que_out_11_4_7, que_out_11_4_6, que_out_11_4_5, que_out_11_4_4, 
      que_out_11_4_3, que_out_11_4_2, que_out_11_4_1, que_out_11_4_0, 
      que_out_12_0_15, que_out_12_0_14, que_out_12_0_13, que_out_12_0_12, 
      que_out_12_0_11, que_out_12_0_10, que_out_12_0_9, que_out_12_0_8, 
      que_out_12_0_7, que_out_12_0_6, que_out_12_0_5, que_out_12_0_4, 
      que_out_12_0_3, que_out_12_0_2, que_out_12_0_1, que_out_12_0_0, 
      que_out_12_1_15, que_out_12_1_14, que_out_12_1_13, que_out_12_1_12, 
      que_out_12_1_11, que_out_12_1_10, que_out_12_1_9, que_out_12_1_8, 
      que_out_12_1_7, que_out_12_1_6, que_out_12_1_5, que_out_12_1_4, 
      que_out_12_1_3, que_out_12_1_2, que_out_12_1_1, que_out_12_1_0, 
      que_out_12_2_15, que_out_12_2_14, que_out_12_2_13, que_out_12_2_12, 
      que_out_12_2_11, que_out_12_2_10, que_out_12_2_9, que_out_12_2_8, 
      que_out_12_2_7, que_out_12_2_6, que_out_12_2_5, que_out_12_2_4, 
      que_out_12_2_3, que_out_12_2_2, que_out_12_2_1, que_out_12_2_0, 
      que_out_12_3_15, que_out_12_3_14, que_out_12_3_13, que_out_12_3_12, 
      que_out_12_3_11, que_out_12_3_10, que_out_12_3_9, que_out_12_3_8, 
      que_out_12_3_7, que_out_12_3_6, que_out_12_3_5, que_out_12_3_4, 
      que_out_12_3_3, que_out_12_3_2, que_out_12_3_1, que_out_12_3_0, 
      que_out_12_4_15, que_out_12_4_14, que_out_12_4_13, que_out_12_4_12, 
      que_out_12_4_11, que_out_12_4_10, que_out_12_4_9, que_out_12_4_8, 
      que_out_12_4_7, que_out_12_4_6, que_out_12_4_5, que_out_12_4_4, 
      que_out_12_4_3, que_out_12_4_2, que_out_12_4_1, que_out_12_4_0, 
      que_out_13_0_15, que_out_13_0_14, que_out_13_0_13, que_out_13_0_12, 
      que_out_13_0_11, que_out_13_0_10, que_out_13_0_9, que_out_13_0_8, 
      que_out_13_0_7, que_out_13_0_6, que_out_13_0_5, que_out_13_0_4, 
      que_out_13_0_3, que_out_13_0_2, que_out_13_0_1, que_out_13_0_0, 
      que_out_13_1_15, que_out_13_1_14, que_out_13_1_13, que_out_13_1_12, 
      que_out_13_1_11, que_out_13_1_10, que_out_13_1_9, que_out_13_1_8, 
      que_out_13_1_7, que_out_13_1_6, que_out_13_1_5, que_out_13_1_4, 
      que_out_13_1_3, que_out_13_1_2, que_out_13_1_1, que_out_13_1_0, 
      que_out_13_2_15, que_out_13_2_14, que_out_13_2_13, que_out_13_2_12, 
      que_out_13_2_11, que_out_13_2_10, que_out_13_2_9, que_out_13_2_8, 
      que_out_13_2_7, que_out_13_2_6, que_out_13_2_5, que_out_13_2_4, 
      que_out_13_2_3, que_out_13_2_2, que_out_13_2_1, que_out_13_2_0, 
      que_out_13_3_15, que_out_13_3_14, que_out_13_3_13, que_out_13_3_12, 
      que_out_13_3_11, que_out_13_3_10, que_out_13_3_9, que_out_13_3_8, 
      que_out_13_3_7, que_out_13_3_6, que_out_13_3_5, que_out_13_3_4, 
      que_out_13_3_3, que_out_13_3_2, que_out_13_3_1, que_out_13_3_0, 
      que_out_13_4_15, que_out_13_4_14, que_out_13_4_13, que_out_13_4_12, 
      que_out_13_4_11, que_out_13_4_10, que_out_13_4_9, que_out_13_4_8, 
      que_out_13_4_7, que_out_13_4_6, que_out_13_4_5, que_out_13_4_4, 
      que_out_13_4_3, que_out_13_4_2, que_out_13_4_1, que_out_13_4_0, 
      que_out_14_0_15, que_out_14_0_14, que_out_14_0_13, que_out_14_0_12, 
      que_out_14_0_11, que_out_14_0_10, que_out_14_0_9, que_out_14_0_8, 
      que_out_14_0_7, que_out_14_0_6, que_out_14_0_5, que_out_14_0_4, 
      que_out_14_0_3, que_out_14_0_2, que_out_14_0_1, que_out_14_0_0, 
      que_out_14_1_15, que_out_14_1_14, que_out_14_1_13, que_out_14_1_12, 
      que_out_14_1_11, que_out_14_1_10, que_out_14_1_9, que_out_14_1_8, 
      que_out_14_1_7, que_out_14_1_6, que_out_14_1_5, que_out_14_1_4, 
      que_out_14_1_3, que_out_14_1_2, que_out_14_1_1, que_out_14_1_0, 
      que_out_14_2_15, que_out_14_2_14, que_out_14_2_13, que_out_14_2_12, 
      que_out_14_2_11, que_out_14_2_10, que_out_14_2_9, que_out_14_2_8, 
      que_out_14_2_7, que_out_14_2_6, que_out_14_2_5, que_out_14_2_4, 
      que_out_14_2_3, que_out_14_2_2, que_out_14_2_1, que_out_14_2_0, 
      que_out_14_3_15, que_out_14_3_14, que_out_14_3_13, que_out_14_3_12, 
      que_out_14_3_11, que_out_14_3_10, que_out_14_3_9, que_out_14_3_8, 
      que_out_14_3_7, que_out_14_3_6, que_out_14_3_5, que_out_14_3_4, 
      que_out_14_3_3, que_out_14_3_2, que_out_14_3_1, que_out_14_3_0, 
      que_out_14_4_15, que_out_14_4_14, que_out_14_4_13, que_out_14_4_12, 
      que_out_14_4_11, que_out_14_4_10, que_out_14_4_9, que_out_14_4_8, 
      que_out_14_4_7, que_out_14_4_6, que_out_14_4_5, que_out_14_4_4, 
      que_out_14_4_3, que_out_14_4_2, que_out_14_4_1, que_out_14_4_0, 
      que_out_15_0_15, que_out_15_0_14, que_out_15_0_13, que_out_15_0_12, 
      que_out_15_0_11, que_out_15_0_10, que_out_15_0_9, que_out_15_0_8, 
      que_out_15_0_7, que_out_15_0_6, que_out_15_0_5, que_out_15_0_4, 
      que_out_15_0_3, que_out_15_0_2, que_out_15_0_1, que_out_15_0_0, 
      que_out_15_1_15, que_out_15_1_14, que_out_15_1_13, que_out_15_1_12, 
      que_out_15_1_11, que_out_15_1_10, que_out_15_1_9, que_out_15_1_8, 
      que_out_15_1_7, que_out_15_1_6, que_out_15_1_5, que_out_15_1_4, 
      que_out_15_1_3, que_out_15_1_2, que_out_15_1_1, que_out_15_1_0, 
      que_out_15_2_15, que_out_15_2_14, que_out_15_2_13, que_out_15_2_12, 
      que_out_15_2_11, que_out_15_2_10, que_out_15_2_9, que_out_15_2_8, 
      que_out_15_2_7, que_out_15_2_6, que_out_15_2_5, que_out_15_2_4, 
      que_out_15_2_3, que_out_15_2_2, que_out_15_2_1, que_out_15_2_0, 
      que_out_15_3_15, que_out_15_3_14, que_out_15_3_13, que_out_15_3_12, 
      que_out_15_3_11, que_out_15_3_10, que_out_15_3_9, que_out_15_3_8, 
      que_out_15_3_7, que_out_15_3_6, que_out_15_3_5, que_out_15_3_4, 
      que_out_15_3_3, que_out_15_3_2, que_out_15_3_1, que_out_15_3_0, 
      que_out_15_4_15, que_out_15_4_14, que_out_15_4_13, que_out_15_4_12, 
      que_out_15_4_11, que_out_15_4_10, que_out_15_4_9, que_out_15_4_8, 
      que_out_15_4_7, que_out_15_4_6, que_out_15_4_5, que_out_15_4_4, 
      que_out_15_4_3, que_out_15_4_2, que_out_15_4_1, que_out_15_4_0, 
      que_out_16_0_15, que_out_16_0_14, que_out_16_0_13, que_out_16_0_12, 
      que_out_16_0_11, que_out_16_0_10, que_out_16_0_9, que_out_16_0_8, 
      que_out_16_0_7, que_out_16_0_6, que_out_16_0_5, que_out_16_0_4, 
      que_out_16_0_3, que_out_16_0_2, que_out_16_0_1, que_out_16_0_0, 
      que_out_16_1_15, que_out_16_1_14, que_out_16_1_13, que_out_16_1_12, 
      que_out_16_1_11, que_out_16_1_10, que_out_16_1_9, que_out_16_1_8, 
      que_out_16_1_7, que_out_16_1_6, que_out_16_1_5, que_out_16_1_4, 
      que_out_16_1_3, que_out_16_1_2, que_out_16_1_1, que_out_16_1_0, 
      que_out_16_2_15, que_out_16_2_14, que_out_16_2_13, que_out_16_2_12, 
      que_out_16_2_11, que_out_16_2_10, que_out_16_2_9, que_out_16_2_8, 
      que_out_16_2_7, que_out_16_2_6, que_out_16_2_5, que_out_16_2_4, 
      que_out_16_2_3, que_out_16_2_2, que_out_16_2_1, que_out_16_2_0, 
      que_out_16_3_15, que_out_16_3_14, que_out_16_3_13, que_out_16_3_12, 
      que_out_16_3_11, que_out_16_3_10, que_out_16_3_9, que_out_16_3_8, 
      que_out_16_3_7, que_out_16_3_6, que_out_16_3_5, que_out_16_3_4, 
      que_out_16_3_3, que_out_16_3_2, que_out_16_3_1, que_out_16_3_0, 
      que_out_16_4_15, que_out_16_4_14, que_out_16_4_13, que_out_16_4_12, 
      que_out_16_4_11, que_out_16_4_10, que_out_16_4_9, que_out_16_4_8, 
      que_out_16_4_7, que_out_16_4_6, que_out_16_4_5, que_out_16_4_4, 
      que_out_16_4_3, que_out_16_4_2, que_out_16_4_1, que_out_16_4_0, 
      que_out_17_0_15, que_out_17_0_14, que_out_17_0_13, que_out_17_0_12, 
      que_out_17_0_11, que_out_17_0_10, que_out_17_0_9, que_out_17_0_8, 
      que_out_17_0_7, que_out_17_0_6, que_out_17_0_5, que_out_17_0_4, 
      que_out_17_0_3, que_out_17_0_2, que_out_17_0_1, que_out_17_0_0, 
      que_out_17_1_15, que_out_17_1_14, que_out_17_1_13, que_out_17_1_12, 
      que_out_17_1_11, que_out_17_1_10, que_out_17_1_9, que_out_17_1_8, 
      que_out_17_1_7, que_out_17_1_6, que_out_17_1_5, que_out_17_1_4, 
      que_out_17_1_3, que_out_17_1_2, que_out_17_1_1, que_out_17_1_0, 
      que_out_17_2_15, que_out_17_2_14, que_out_17_2_13, que_out_17_2_12, 
      que_out_17_2_11, que_out_17_2_10, que_out_17_2_9, que_out_17_2_8, 
      que_out_17_2_7, que_out_17_2_6, que_out_17_2_5, que_out_17_2_4, 
      que_out_17_2_3, que_out_17_2_2, que_out_17_2_1, que_out_17_2_0, 
      que_out_17_3_15, que_out_17_3_14, que_out_17_3_13, que_out_17_3_12, 
      que_out_17_3_11, que_out_17_3_10, que_out_17_3_9, que_out_17_3_8, 
      que_out_17_3_7, que_out_17_3_6, que_out_17_3_5, que_out_17_3_4, 
      que_out_17_3_3, que_out_17_3_2, que_out_17_3_1, que_out_17_3_0, 
      que_out_17_4_15, que_out_17_4_14, que_out_17_4_13, que_out_17_4_12, 
      que_out_17_4_11, que_out_17_4_10, que_out_17_4_9, que_out_17_4_8, 
      que_out_17_4_7, que_out_17_4_6, que_out_17_4_5, que_out_17_4_4, 
      que_out_17_4_3, que_out_17_4_2, que_out_17_4_1, que_out_17_4_0, 
      que_out_18_0_15, que_out_18_0_14, que_out_18_0_13, que_out_18_0_12, 
      que_out_18_0_11, que_out_18_0_10, que_out_18_0_9, que_out_18_0_8, 
      que_out_18_0_7, que_out_18_0_6, que_out_18_0_5, que_out_18_0_4, 
      que_out_18_0_3, que_out_18_0_2, que_out_18_0_1, que_out_18_0_0, 
      que_out_18_1_15, que_out_18_1_14, que_out_18_1_13, que_out_18_1_12, 
      que_out_18_1_11, que_out_18_1_10, que_out_18_1_9, que_out_18_1_8, 
      que_out_18_1_7, que_out_18_1_6, que_out_18_1_5, que_out_18_1_4, 
      que_out_18_1_3, que_out_18_1_2, que_out_18_1_1, que_out_18_1_0, 
      que_out_18_2_15, que_out_18_2_14, que_out_18_2_13, que_out_18_2_12, 
      que_out_18_2_11, que_out_18_2_10, que_out_18_2_9, que_out_18_2_8, 
      que_out_18_2_7, que_out_18_2_6, que_out_18_2_5, que_out_18_2_4, 
      que_out_18_2_3, que_out_18_2_2, que_out_18_2_1, que_out_18_2_0, 
      que_out_18_3_15, que_out_18_3_14, que_out_18_3_13, que_out_18_3_12, 
      que_out_18_3_11, que_out_18_3_10, que_out_18_3_9, que_out_18_3_8, 
      que_out_18_3_7, que_out_18_3_6, que_out_18_3_5, que_out_18_3_4, 
      que_out_18_3_3, que_out_18_3_2, que_out_18_3_1, que_out_18_3_0, 
      que_out_18_4_15, que_out_18_4_14, que_out_18_4_13, que_out_18_4_12, 
      que_out_18_4_11, que_out_18_4_10, que_out_18_4_9, que_out_18_4_8, 
      que_out_18_4_7, que_out_18_4_6, que_out_18_4_5, que_out_18_4_4, 
      que_out_18_4_3, que_out_18_4_2, que_out_18_4_1, que_out_18_4_0, 
      que_out_19_0_15, que_out_19_0_14, que_out_19_0_13, que_out_19_0_12, 
      que_out_19_0_11, que_out_19_0_10, que_out_19_0_9, que_out_19_0_8, 
      que_out_19_0_7, que_out_19_0_6, que_out_19_0_5, que_out_19_0_4, 
      que_out_19_0_3, que_out_19_0_2, que_out_19_0_1, que_out_19_0_0, 
      que_out_19_1_15, que_out_19_1_14, que_out_19_1_13, que_out_19_1_12, 
      que_out_19_1_11, que_out_19_1_10, que_out_19_1_9, que_out_19_1_8, 
      que_out_19_1_7, que_out_19_1_6, que_out_19_1_5, que_out_19_1_4, 
      que_out_19_1_3, que_out_19_1_2, que_out_19_1_1, que_out_19_1_0, 
      que_out_19_2_15, que_out_19_2_14, que_out_19_2_13, que_out_19_2_12, 
      que_out_19_2_11, que_out_19_2_10, que_out_19_2_9, que_out_19_2_8, 
      que_out_19_2_7, que_out_19_2_6, que_out_19_2_5, que_out_19_2_4, 
      que_out_19_2_3, que_out_19_2_2, que_out_19_2_1, que_out_19_2_0, 
      que_out_19_3_15, que_out_19_3_14, que_out_19_3_13, que_out_19_3_12, 
      que_out_19_3_11, que_out_19_3_10, que_out_19_3_9, que_out_19_3_8, 
      que_out_19_3_7, que_out_19_3_6, que_out_19_3_5, que_out_19_3_4, 
      que_out_19_3_3, que_out_19_3_2, que_out_19_3_1, que_out_19_3_0, 
      que_out_19_4_15, que_out_19_4_14, que_out_19_4_13, que_out_19_4_12, 
      que_out_19_4_11, que_out_19_4_10, que_out_19_4_9, que_out_19_4_8, 
      que_out_19_4_7, que_out_19_4_6, que_out_19_4_5, que_out_19_4_4, 
      que_out_19_4_3, que_out_19_4_2, que_out_19_4_1, que_out_19_4_0, 
      que_out_20_0_15, que_out_20_0_14, que_out_20_0_13, que_out_20_0_12, 
      que_out_20_0_11, que_out_20_0_10, que_out_20_0_9, que_out_20_0_8, 
      que_out_20_0_7, que_out_20_0_6, que_out_20_0_5, que_out_20_0_4, 
      que_out_20_0_3, que_out_20_0_2, que_out_20_0_1, que_out_20_0_0, 
      que_out_20_1_15, que_out_20_1_14, que_out_20_1_13, que_out_20_1_12, 
      que_out_20_1_11, que_out_20_1_10, que_out_20_1_9, que_out_20_1_8, 
      que_out_20_1_7, que_out_20_1_6, que_out_20_1_5, que_out_20_1_4, 
      que_out_20_1_3, que_out_20_1_2, que_out_20_1_1, que_out_20_1_0, 
      que_out_20_2_15, que_out_20_2_14, que_out_20_2_13, que_out_20_2_12, 
      que_out_20_2_11, que_out_20_2_10, que_out_20_2_9, que_out_20_2_8, 
      que_out_20_2_7, que_out_20_2_6, que_out_20_2_5, que_out_20_2_4, 
      que_out_20_2_3, que_out_20_2_2, que_out_20_2_1, que_out_20_2_0, 
      que_out_20_3_15, que_out_20_3_14, que_out_20_3_13, que_out_20_3_12, 
      que_out_20_3_11, que_out_20_3_10, que_out_20_3_9, que_out_20_3_8, 
      que_out_20_3_7, que_out_20_3_6, que_out_20_3_5, que_out_20_3_4, 
      que_out_20_3_3, que_out_20_3_2, que_out_20_3_1, que_out_20_3_0, 
      que_out_20_4_15, que_out_20_4_14, que_out_20_4_13, que_out_20_4_12, 
      que_out_20_4_11, que_out_20_4_10, que_out_20_4_9, que_out_20_4_8, 
      que_out_20_4_7, que_out_20_4_6, que_out_20_4_5, que_out_20_4_4, 
      que_out_20_4_3, que_out_20_4_2, que_out_20_4_1, que_out_20_4_0, 
      que_out_21_0_15, que_out_21_0_14, que_out_21_0_13, que_out_21_0_12, 
      que_out_21_0_11, que_out_21_0_10, que_out_21_0_9, que_out_21_0_8, 
      que_out_21_0_7, que_out_21_0_6, que_out_21_0_5, que_out_21_0_4, 
      que_out_21_0_3, que_out_21_0_2, que_out_21_0_1, que_out_21_0_0, 
      que_out_21_1_15, que_out_21_1_14, que_out_21_1_13, que_out_21_1_12, 
      que_out_21_1_11, que_out_21_1_10, que_out_21_1_9, que_out_21_1_8, 
      que_out_21_1_7, que_out_21_1_6, que_out_21_1_5, que_out_21_1_4, 
      que_out_21_1_3, que_out_21_1_2, que_out_21_1_1, que_out_21_1_0, 
      que_out_21_2_15, que_out_21_2_14, que_out_21_2_13, que_out_21_2_12, 
      que_out_21_2_11, que_out_21_2_10, que_out_21_2_9, que_out_21_2_8, 
      que_out_21_2_7, que_out_21_2_6, que_out_21_2_5, que_out_21_2_4, 
      que_out_21_2_3, que_out_21_2_2, que_out_21_2_1, que_out_21_2_0, 
      que_out_21_3_15, que_out_21_3_14, que_out_21_3_13, que_out_21_3_12, 
      que_out_21_3_11, que_out_21_3_10, que_out_21_3_9, que_out_21_3_8, 
      que_out_21_3_7, que_out_21_3_6, que_out_21_3_5, que_out_21_3_4, 
      que_out_21_3_3, que_out_21_3_2, que_out_21_3_1, que_out_21_3_0, 
      que_out_21_4_15, que_out_21_4_14, que_out_21_4_13, que_out_21_4_12, 
      que_out_21_4_11, que_out_21_4_10, que_out_21_4_9, que_out_21_4_8, 
      que_out_21_4_7, que_out_21_4_6, que_out_21_4_5, que_out_21_4_4, 
      que_out_21_4_3, que_out_21_4_2, que_out_21_4_1, que_out_21_4_0, 
      que_out_22_0_15, que_out_22_0_14, que_out_22_0_13, que_out_22_0_12, 
      que_out_22_0_11, que_out_22_0_10, que_out_22_0_9, que_out_22_0_8, 
      que_out_22_0_7, que_out_22_0_6, que_out_22_0_5, que_out_22_0_4, 
      que_out_22_0_3, que_out_22_0_2, que_out_22_0_1, que_out_22_0_0, 
      que_out_22_1_15, que_out_22_1_14, que_out_22_1_13, que_out_22_1_12, 
      que_out_22_1_11, que_out_22_1_10, que_out_22_1_9, que_out_22_1_8, 
      que_out_22_1_7, que_out_22_1_6, que_out_22_1_5, que_out_22_1_4, 
      que_out_22_1_3, que_out_22_1_2, que_out_22_1_1, que_out_22_1_0, 
      que_out_22_2_15, que_out_22_2_14, que_out_22_2_13, que_out_22_2_12, 
      que_out_22_2_11, que_out_22_2_10, que_out_22_2_9, que_out_22_2_8, 
      que_out_22_2_7, que_out_22_2_6, que_out_22_2_5, que_out_22_2_4, 
      que_out_22_2_3, que_out_22_2_2, que_out_22_2_1, que_out_22_2_0, 
      que_out_22_3_15, que_out_22_3_14, que_out_22_3_13, que_out_22_3_12, 
      que_out_22_3_11, que_out_22_3_10, que_out_22_3_9, que_out_22_3_8, 
      que_out_22_3_7, que_out_22_3_6, que_out_22_3_5, que_out_22_3_4, 
      que_out_22_3_3, que_out_22_3_2, que_out_22_3_1, que_out_22_3_0, 
      que_out_22_4_15, que_out_22_4_14, que_out_22_4_13, que_out_22_4_12, 
      que_out_22_4_11, que_out_22_4_10, que_out_22_4_9, que_out_22_4_8, 
      que_out_22_4_7, que_out_22_4_6, que_out_22_4_5, que_out_22_4_4, 
      que_out_22_4_3, que_out_22_4_2, que_out_22_4_1, que_out_22_4_0, 
      que_out_23_0_15, que_out_23_0_14, que_out_23_0_13, que_out_23_0_12, 
      que_out_23_0_11, que_out_23_0_10, que_out_23_0_9, que_out_23_0_8, 
      que_out_23_0_7, que_out_23_0_6, que_out_23_0_5, que_out_23_0_4, 
      que_out_23_0_3, que_out_23_0_2, que_out_23_0_1, que_out_23_0_0, 
      que_out_23_1_15, que_out_23_1_14, que_out_23_1_13, que_out_23_1_12, 
      que_out_23_1_11, que_out_23_1_10, que_out_23_1_9, que_out_23_1_8, 
      que_out_23_1_7, que_out_23_1_6, que_out_23_1_5, que_out_23_1_4, 
      que_out_23_1_3, que_out_23_1_2, que_out_23_1_1, que_out_23_1_0, 
      que_out_23_2_15, que_out_23_2_14, que_out_23_2_13, que_out_23_2_12, 
      que_out_23_2_11, que_out_23_2_10, que_out_23_2_9, que_out_23_2_8, 
      que_out_23_2_7, que_out_23_2_6, que_out_23_2_5, que_out_23_2_4, 
      que_out_23_2_3, que_out_23_2_2, que_out_23_2_1, que_out_23_2_0, 
      que_out_23_3_15, que_out_23_3_14, que_out_23_3_13, que_out_23_3_12, 
      que_out_23_3_11, que_out_23_3_10, que_out_23_3_9, que_out_23_3_8, 
      que_out_23_3_7, que_out_23_3_6, que_out_23_3_5, que_out_23_3_4, 
      que_out_23_3_3, que_out_23_3_2, que_out_23_3_1, que_out_23_3_0, 
      que_out_23_4_15, que_out_23_4_14, que_out_23_4_13, que_out_23_4_12, 
      que_out_23_4_11, que_out_23_4_10, que_out_23_4_9, que_out_23_4_8, 
      que_out_23_4_7, que_out_23_4_6, que_out_23_4_5, que_out_23_4_4, 
      que_out_23_4_3, que_out_23_4_2, que_out_23_4_1, que_out_23_4_0, 
      que_out_24_0_15, que_out_24_0_14, que_out_24_0_13, que_out_24_0_12, 
      que_out_24_0_11, que_out_24_0_10, que_out_24_0_9, que_out_24_0_8, 
      que_out_24_0_7, que_out_24_0_6, que_out_24_0_5, que_out_24_0_4, 
      que_out_24_0_3, que_out_24_0_2, que_out_24_0_1, que_out_24_0_0, 
      que_out_24_1_15, que_out_24_1_14, que_out_24_1_13, que_out_24_1_12, 
      que_out_24_1_11, que_out_24_1_10, que_out_24_1_9, que_out_24_1_8, 
      que_out_24_1_7, que_out_24_1_6, que_out_24_1_5, que_out_24_1_4, 
      que_out_24_1_3, que_out_24_1_2, que_out_24_1_1, que_out_24_1_0, 
      que_out_24_2_15, que_out_24_2_14, que_out_24_2_13, que_out_24_2_12, 
      que_out_24_2_11, que_out_24_2_10, que_out_24_2_9, que_out_24_2_8, 
      que_out_24_2_7, que_out_24_2_6, que_out_24_2_5, que_out_24_2_4, 
      que_out_24_2_3, que_out_24_2_2, que_out_24_2_1, que_out_24_2_0, 
      que_out_24_3_15, que_out_24_3_14, que_out_24_3_13, que_out_24_3_12, 
      que_out_24_3_11, que_out_24_3_10, que_out_24_3_9, que_out_24_3_8, 
      que_out_24_3_7, que_out_24_3_6, que_out_24_3_5, que_out_24_3_4, 
      que_out_24_3_3, que_out_24_3_2, que_out_24_3_1, que_out_24_3_0, 
      que_out_24_4_15, que_out_24_4_14, que_out_24_4_13, que_out_24_4_12, 
      que_out_24_4_11, que_out_24_4_10, que_out_24_4_9, que_out_24_4_8, 
      que_out_24_4_7, que_out_24_4_6, que_out_24_4_5, que_out_24_4_4, 
      que_out_24_4_3, que_out_24_4_2, que_out_24_4_1, que_out_24_4_0, 
      que_out_25_0_15, que_out_25_0_14, que_out_25_0_13, que_out_25_0_12, 
      que_out_25_0_11, que_out_25_0_10, que_out_25_0_9, que_out_25_0_8, 
      que_out_25_0_7, que_out_25_0_6, que_out_25_0_5, que_out_25_0_4, 
      que_out_25_0_3, que_out_25_0_2, que_out_25_0_1, que_out_25_0_0, 
      que_out_25_1_15, que_out_25_1_14, que_out_25_1_13, que_out_25_1_12, 
      que_out_25_1_11, que_out_25_1_10, que_out_25_1_9, que_out_25_1_8, 
      que_out_25_1_7, que_out_25_1_6, que_out_25_1_5, que_out_25_1_4, 
      que_out_25_1_3, que_out_25_1_2, que_out_25_1_1, que_out_25_1_0, 
      que_out_25_2_15, que_out_25_2_14, que_out_25_2_13, que_out_25_2_12, 
      que_out_25_2_11, que_out_25_2_10, que_out_25_2_9, que_out_25_2_8, 
      que_out_25_2_7, que_out_25_2_6, que_out_25_2_5, que_out_25_2_4, 
      que_out_25_2_3, que_out_25_2_2, que_out_25_2_1, que_out_25_2_0, 
      que_out_25_3_15, que_out_25_3_14, que_out_25_3_13, que_out_25_3_12, 
      que_out_25_3_11, que_out_25_3_10, que_out_25_3_9, que_out_25_3_8, 
      que_out_25_3_7, que_out_25_3_6, que_out_25_3_5, que_out_25_3_4, 
      que_out_25_3_3, que_out_25_3_2, que_out_25_3_1, que_out_25_3_0, 
      que_out_25_4_15, que_out_25_4_14, que_out_25_4_13, que_out_25_4_12, 
      que_out_25_4_11, que_out_25_4_10, que_out_25_4_9, que_out_25_4_8, 
      que_out_25_4_7, que_out_25_4_6, que_out_25_4_5, que_out_25_4_4, 
      que_out_25_4_3, que_out_25_4_2, que_out_25_4_1, que_out_25_4_0, 
      que_out_26_0_15, que_out_26_0_14, que_out_26_0_13, que_out_26_0_12, 
      que_out_26_0_11, que_out_26_0_10, que_out_26_0_9, que_out_26_0_8, 
      que_out_26_0_7, que_out_26_0_6, que_out_26_0_5, que_out_26_0_4, 
      que_out_26_0_3, que_out_26_0_2, que_out_26_0_1, que_out_26_0_0, 
      que_out_26_1_15, que_out_26_1_14, que_out_26_1_13, que_out_26_1_12, 
      que_out_26_1_11, que_out_26_1_10, que_out_26_1_9, que_out_26_1_8, 
      que_out_26_1_7, que_out_26_1_6, que_out_26_1_5, que_out_26_1_4, 
      que_out_26_1_3, que_out_26_1_2, que_out_26_1_1, que_out_26_1_0, 
      que_out_26_2_15, que_out_26_2_14, que_out_26_2_13, que_out_26_2_12, 
      que_out_26_2_11, que_out_26_2_10, que_out_26_2_9, que_out_26_2_8, 
      que_out_26_2_7, que_out_26_2_6, que_out_26_2_5, que_out_26_2_4, 
      que_out_26_2_3, que_out_26_2_2, que_out_26_2_1, que_out_26_2_0, 
      que_out_26_3_15, que_out_26_3_14, que_out_26_3_13, que_out_26_3_12, 
      que_out_26_3_11, que_out_26_3_10, que_out_26_3_9, que_out_26_3_8, 
      que_out_26_3_7, que_out_26_3_6, que_out_26_3_5, que_out_26_3_4, 
      que_out_26_3_3, que_out_26_3_2, que_out_26_3_1, que_out_26_3_0, 
      que_out_26_4_15, que_out_26_4_14, que_out_26_4_13, que_out_26_4_12, 
      que_out_26_4_11, que_out_26_4_10, que_out_26_4_9, que_out_26_4_8, 
      que_out_26_4_7, que_out_26_4_6, que_out_26_4_5, que_out_26_4_4, 
      que_out_26_4_3, que_out_26_4_2, que_out_26_4_1, que_out_26_4_0, 
      que_out_27_0_15, que_out_27_0_14, que_out_27_0_13, que_out_27_0_12, 
      que_out_27_0_11, que_out_27_0_10, que_out_27_0_9, que_out_27_0_8, 
      que_out_27_0_7, que_out_27_0_6, que_out_27_0_5, que_out_27_0_4, 
      que_out_27_0_3, que_out_27_0_2, que_out_27_0_1, que_out_27_0_0, 
      que_out_27_1_15, que_out_27_1_14, que_out_27_1_13, que_out_27_1_12, 
      que_out_27_1_11, que_out_27_1_10, que_out_27_1_9, que_out_27_1_8, 
      que_out_27_1_7, que_out_27_1_6, que_out_27_1_5, que_out_27_1_4, 
      que_out_27_1_3, que_out_27_1_2, que_out_27_1_1, que_out_27_1_0, 
      que_out_27_2_15, que_out_27_2_14, que_out_27_2_13, que_out_27_2_12, 
      que_out_27_2_11, que_out_27_2_10, que_out_27_2_9, que_out_27_2_8, 
      que_out_27_2_7, que_out_27_2_6, que_out_27_2_5, que_out_27_2_4, 
      que_out_27_2_3, que_out_27_2_2, que_out_27_2_1, que_out_27_2_0, 
      que_out_27_3_15, que_out_27_3_14, que_out_27_3_13, que_out_27_3_12, 
      que_out_27_3_11, que_out_27_3_10, que_out_27_3_9, que_out_27_3_8, 
      que_out_27_3_7, que_out_27_3_6, que_out_27_3_5, que_out_27_3_4, 
      que_out_27_3_3, que_out_27_3_2, que_out_27_3_1, que_out_27_3_0, 
      que_out_27_4_15, que_out_27_4_14, que_out_27_4_13, que_out_27_4_12, 
      que_out_27_4_11, que_out_27_4_10, que_out_27_4_9, que_out_27_4_8, 
      que_out_27_4_7, que_out_27_4_6, que_out_27_4_5, que_out_27_4_4, 
      que_out_27_4_3, que_out_27_4_2, que_out_27_4_1, que_out_27_4_0, 
      sel_que_27, sel_que_26, sel_que_25, sel_que_24, sel_que_23, sel_que_22, 
      sel_que_21, sel_que_20, sel_que_19, sel_que_18, sel_que_17, sel_que_16, 
      sel_que_15, sel_que_14, sel_que_13, sel_que_12, sel_que_11, sel_que_10, 
      sel_que_9, sel_que_8, sel_que_7, sel_que_6, sel_que_5, sel_que_4, 
      sel_que_3, sel_que_2, sel_que_1, sel_que_0, nx12, nx14, nx28, nx30, 
      nx42, nx48, nx62, nx64, nx68, nx74, nx82, nx88, nx90, nx94, nx100, 
      nx104, nx114, nx118, nx122, nx130, nx136, nx144, nx150, nx158, nx166, 
      nx172, nx180, nx188, nx192, nx200, nx206, nx214, nx222, nx226, nx230, 
      nx238, nx268, nx294, nx322, nx348, nx378, nx404, nx432, nx458, nx488, 
      nx514, nx542, nx568, nx598, nx624, nx652, nx678, nx708, nx734, nx762, 
      nx788, nx818, nx844, nx872, nx898, nx928, nx954, nx982, nx1008, nx1038, 
      nx1064, nx1092, nx1118, nx1148, nx1174, nx1202, nx1228, nx1258, nx1284, 
      nx1312, nx1338, nx1368, nx1394, nx1422, nx1448, nx1478, nx1504, nx1532, 
      nx1558, nx1588, nx1614, nx1642, nx1668, nx1698, nx1724, nx1752, nx1778, 
      nx1808, nx1834, nx1862, nx1888, nx1918, nx1944, nx1972, nx1998, nx2028, 
      nx2054, nx2082, nx2108, nx2138, nx2164, nx2192, nx2218, nx2248, nx2274, 
      nx2302, nx2328, nx2358, nx2384, nx2412, nx2438, nx2468, nx2494, nx2522, 
      nx2548, nx2578, nx2604, nx2632, nx2658, nx2688, nx2714, nx2742, nx2768, 
      nx2798, nx2824, nx2852, nx2878, nx2908, nx2934, nx2962, nx2988, nx3018, 
      nx3044, nx3072, nx3098, nx3128, nx3154, nx3182, nx3208, nx3238, nx3264, 
      nx3292, nx3318, nx3348, nx3374, nx3402, nx3428, nx3458, nx3484, nx3512, 
      nx3538, nx3568, nx3594, nx3622, nx3648, nx3678, nx3704, nx3732, nx3758, 
      nx3788, nx3814, nx3842, nx3868, nx3898, nx3924, nx3952, nx3978, nx4008, 
      nx4034, nx4062, nx4088, nx4118, nx4144, nx4172, nx4198, nx4228, nx4254, 
      nx4282, nx4308, nx4338, nx4364, nx4392, nx4418, nx4448, nx4474, nx4502, 
      nx4528, nx4558, nx4584, nx4612, nx4638, nx4668, nx4694, nx4722, nx4748, 
      nx4778, nx4804, nx4832, nx4858, nx4888, nx4914, nx4942, nx4968, nx4998, 
      nx5024, nx5052, nx5078, nx5108, nx5134, nx5162, nx5188, nx5218, nx5244, 
      nx5272, nx5298, nx5328, nx5354, nx5382, nx5408, nx5438, nx5464, nx5492, 
      nx5518, nx5548, nx5574, nx5602, nx5628, nx5658, nx5684, nx5712, nx5738, 
      nx5768, nx5794, nx5822, nx5848, nx5878, nx5904, nx5932, nx5958, nx5988, 
      nx6014, nx6042, nx6068, nx6098, nx6124, nx6152, nx6178, nx6208, nx6234, 
      nx6262, nx6288, nx6318, nx6344, nx6372, nx6398, nx6428, nx6454, nx6482, 
      nx6508, nx6538, nx6564, nx6592, nx6618, nx6648, nx6674, nx6702, nx6728, 
      nx6758, nx6784, nx6812, nx6838, nx6868, nx6894, nx6922, nx6948, nx6978, 
      nx7004, nx7032, nx7058, nx7088, nx7114, nx7142, nx7168, nx7198, nx7224, 
      nx7252, nx7278, nx7308, nx7334, nx7362, nx7388, nx7418, nx7444, nx7472, 
      nx7498, nx7528, nx7554, nx7582, nx7608, nx7638, nx7664, nx7692, nx7718, 
      nx7748, nx7774, nx7802, nx7828, nx7858, nx7884, nx7912, nx7938, nx7968, 
      nx7994, nx8022, nx8048, nx8078, nx8104, nx8132, nx8158, nx8188, nx8214, 
      nx8242, nx8268, nx8298, nx8324, nx8352, nx8378, nx8408, nx8434, nx8462, 
      nx8488, nx8518, nx8544, nx8572, nx8598, nx8628, nx8654, nx8682, nx8708, 
      nx8738, nx8764, nx8792, nx8818, nx8848, nx8874, nx8902, nx8928, nx8938, 
      nx9038, nx6829, nx6833, nx6835, nx6839, nx6843, nx6847, nx6875, nx6885, 
      nx6889, nx6893, nx6897, nx6901, nx6905, nx6915, nx6927, nx6931, nx6933, 
      nx6937, nx6939, nx6943, nx6945, nx6949, nx6951, nx6955, nx6957, nx6961, 
      nx6965, nx6967, nx6971, nx6977, nx6985, nx6991, nx6999, nx7007, nx7017, 
      nx7029, nx7037, nx7043, nx7053, nx7055, nx7057, nx7061, nx7063, nx7065, 
      nx7069, nx7071, nx7073, nx7077, nx7079, nx7081, nx7087, nx7089, nx7091, 
      nx7095, nx7097, nx7099, nx7103, nx7105, nx7107, nx7111, nx7113, nx7115, 
      nx7121, nx7123, nx7125, nx7129, nx7131, nx7133, nx7137, nx7139, nx7141, 
      nx7145, nx7147, nx7149, nx7155, nx7157, nx7159, nx7163, nx7165, nx7167, 
      nx7171, nx7173, nx7175, nx7179, nx7181, nx7183, nx7189, nx7191, nx7193, 
      nx7197, nx7199, nx7201, nx7205, nx7207, nx7209, nx7213, nx7215, nx7217, 
      nx7223, nx7225, nx7227, nx7231, nx7233, nx7235, nx7239, nx7241, nx7243, 
      nx7247, nx7249, nx7251, nx7257, nx7259, nx7261, nx7265, nx7267, nx7269, 
      nx7273, nx7275, nx7277, nx7281, nx7283, nx7285, nx7291, nx7293, nx7295, 
      nx7299, nx7301, nx7303, nx7307, nx7309, nx7311, nx7315, nx7317, nx7319, 
      nx7325, nx7327, nx7329, nx7333, nx7335, nx7337, nx7341, nx7343, nx7345, 
      nx7349, nx7351, nx7353, nx7359, nx7361, nx7363, nx7367, nx7369, nx7371, 
      nx7375, nx7377, nx7379, nx7383, nx7385, nx7387, nx7393, nx7395, nx7397, 
      nx7401, nx7403, nx7405, nx7409, nx7411, nx7413, nx7417, nx7419, nx7421, 
      nx7427, nx7429, nx7431, nx7435, nx7437, nx7439, nx7443, nx7445, nx7447, 
      nx7451, nx7453, nx7455, nx7461, nx7463, nx7465, nx7469, nx7471, nx7473, 
      nx7477, nx7479, nx7481, nx7485, nx7487, nx7489, nx7495, nx7497, nx7499, 
      nx7503, nx7505, nx7507, nx7511, nx7513, nx7515, nx7519, nx7521, nx7523, 
      nx7529, nx7531, nx7533, nx7537, nx7539, nx7541, nx7545, nx7547, nx7549, 
      nx7553, nx7555, nx7557, nx7563, nx7565, nx7567, nx7571, nx7573, nx7575, 
      nx7579, nx7581, nx7583, nx7587, nx7589, nx7591, nx7597, nx7599, nx7601, 
      nx7605, nx7607, nx7609, nx7613, nx7615, nx7617, nx7621, nx7623, nx7625, 
      nx7631, nx7633, nx7635, nx7639, nx7641, nx7643, nx7647, nx7649, nx7651, 
      nx7655, nx7657, nx7659, nx7665, nx7667, nx7669, nx7673, nx7675, nx7677, 
      nx7681, nx7683, nx7685, nx7689, nx7691, nx7693, nx7699, nx7701, nx7703, 
      nx7707, nx7709, nx7711, nx7715, nx7717, nx7719, nx7723, nx7725, nx7727, 
      nx7733, nx7735, nx7737, nx7741, nx7743, nx7745, nx7749, nx7751, nx7753, 
      nx7757, nx7759, nx7761, nx7767, nx7769, nx7771, nx7775, nx7777, nx7779, 
      nx7783, nx7785, nx7787, nx7791, nx7793, nx7795, nx7801, nx7803, nx7805, 
      nx7809, nx7811, nx7813, nx7817, nx7819, nx7821, nx7825, nx7827, nx7829, 
      nx7835, nx7837, nx7839, nx7843, nx7845, nx7847, nx7851, nx7853, nx7855, 
      nx7859, nx7861, nx7863, nx7869, nx7871, nx7873, nx7877, nx7879, nx7881, 
      nx7885, nx7887, nx7889, nx7893, nx7895, nx7897, nx7903, nx7905, nx7907, 
      nx7911, nx7913, nx7915, nx7919, nx7921, nx7923, nx7927, nx7929, nx7931, 
      nx7937, nx7939, nx7941, nx7945, nx7947, nx7949, nx7953, nx7955, nx7957, 
      nx7961, nx7963, nx7965, nx7971, nx7973, nx7975, nx7979, nx7981, nx7983, 
      nx7987, nx7989, nx7991, nx7995, nx7997, nx7999, nx8005, nx8007, nx8009, 
      nx8013, nx8015, nx8017, nx8021, nx8023, nx8025, nx8029, nx8031, nx8033, 
      nx8039, nx8041, nx8043, nx8047, nx8049, nx8051, nx8055, nx8057, nx8059, 
      nx8063, nx8065, nx8067, nx8073, nx8075, nx8077, nx8081, nx8083, nx8085, 
      nx8089, nx8091, nx8093, nx8097, nx8099, nx8101, nx8107, nx8109, nx8111, 
      nx8115, nx8117, nx8119, nx8123, nx8125, nx8127, nx8131, nx8133, nx8135, 
      nx8141, nx8143, nx8145, nx8149, nx8151, nx8153, nx8157, nx8159, nx8161, 
      nx8165, nx8167, nx8169, nx8175, nx8177, nx8179, nx8183, nx8185, nx8187, 
      nx8191, nx8193, nx8195, nx8199, nx8201, nx8203, nx8209, nx8211, nx8213, 
      nx8217, nx8219, nx8221, nx8225, nx8227, nx8229, nx8233, nx8235, nx8237, 
      nx8243, nx8245, nx8247, nx8251, nx8253, nx8255, nx8259, nx8261, nx8263, 
      nx8267, nx8269, nx8271, nx8277, nx8279, nx8281, nx8285, nx8287, nx8289, 
      nx8293, nx8295, nx8297, nx8301, nx8303, nx8305, nx8311, nx8313, nx8315, 
      nx8319, nx8321, nx8323, nx8327, nx8329, nx8331, nx8335, nx8337, nx8339, 
      nx8345, nx8347, nx8349, nx8353, nx8355, nx8357, nx8361, nx8363, nx8365, 
      nx8369, nx8371, nx8373, nx8379, nx8381, nx8383, nx8387, nx8389, nx8391, 
      nx8395, nx8397, nx8399, nx8403, nx8405, nx8407, nx8413, nx8415, nx8417, 
      nx8421, nx8423, nx8425, nx8429, nx8431, nx8433, nx8437, nx8439, nx8441, 
      nx8447, nx8449, nx8451, nx8455, nx8457, nx8459, nx8463, nx8465, nx8467, 
      nx8471, nx8473, nx8475, nx8481, nx8483, nx8485, nx8489, nx8491, nx8493, 
      nx8497, nx8499, nx8501, nx8505, nx8507, nx8509, nx8515, nx8517, nx8519, 
      nx8523, nx8525, nx8527, nx8531, nx8533, nx8535, nx8539, nx8541, nx8543, 
      nx8549, nx8551, nx8553, nx8557, nx8559, nx8561, nx8565, nx8567, nx8569, 
      nx8573, nx8575, nx8577, nx8583, nx8585, nx8587, nx8591, nx8593, nx8595, 
      nx8599, nx8601, nx8603, nx8607, nx8609, nx8611, nx8617, nx8619, nx8621, 
      nx8625, nx8627, nx8629, nx8633, nx8635, nx8637, nx8641, nx8643, nx8645, 
      nx8651, nx8653, nx8655, nx8659, nx8661, nx8663, nx8667, nx8669, nx8671, 
      nx8675, nx8677, nx8679, nx8685, nx8687, nx8689, nx8693, nx8695, nx8697, 
      nx8701, nx8703, nx8705, nx8709, nx8711, nx8713, nx8719, nx8721, nx8723, 
      nx8727, nx8729, nx8731, nx8735, nx8737, nx8739, nx8743, nx8745, nx8747, 
      nx8753, nx8755, nx8757, nx8761, nx8763, nx8765, nx8769, nx8771, nx8773, 
      nx8777, nx8779, nx8781, nx8787, nx8789, nx8791, nx8795, nx8797, nx8799, 
      nx8803, nx8805, nx8807, nx8811, nx8813, nx8815, nx8821, nx8823, nx8825, 
      nx8829, nx8831, nx8833, nx8837, nx8839, nx8841, nx8845, nx8847, nx8849, 
      nx8855, nx8857, nx8859, nx8863, nx8865, nx8867, nx8871, nx8873, nx8875, 
      nx8879, nx8881, nx8883, nx8889, nx8891, nx8893, nx8897, nx8899, nx8901, 
      nx8905, nx8907, nx8909, nx8913, nx8915, nx8917, nx8923, nx8925, nx8927, 
      nx8931, nx8933, nx8935, nx8939, nx8941, nx8943, nx8947, nx8949, nx8951, 
      nx8955, nx8957, nx8959, nx8963, nx8965, nx8967, nx8970, nx8973, nx8975, 
      nx8978, nx8981, nx8983, nx8989, nx8991, nx8993, nx8997, nx8999, nx9001, 
      nx9005, nx9007, nx9009, nx9013, nx9015, nx9017, nx9023, nx9025, nx9027, 
      nx9031, nx9033, nx9035, nx9039, nx9041, nx9043, nx9047, nx9049, nx9051, 
      nx9057, nx9059, nx9061, nx9065, nx9067, nx9069, nx9073, nx9075, nx9077, 
      nx9081, nx9083, nx9085, nx9090, nx9093, nx9095, nx9098, nx9101, nx9103, 
      nx9106, nx9108, nx9110, nx9113, nx9115, nx9117, nx9121, nx9123, nx9125, 
      nx9128, nx9130, nx9132, nx9135, nx9137, nx9139, nx9142, nx9144, nx9146, 
      nx9150, nx9152, nx9154, nx9157, nx9159, nx9161, nx9164, nx9166, nx9168, 
      nx9171, nx9173, nx9175, nx9179, nx9181, nx9183, nx9186, nx9188, nx9190, 
      nx9193, nx9195, nx9197, nx9200, nx9202, nx9204, nx9208, nx9210, nx9212, 
      nx9215, nx9217, nx9219, nx9222, nx9224, nx9226, nx9229, nx9231, nx9233, 
      nx9237, nx9239, nx9241, nx9244, nx9246, nx9248, nx9251, nx9253, nx9255, 
      nx9258, nx9260, nx9262, nx9266, nx9268, nx9270, nx9273, nx9275, nx9277, 
      nx9280, nx9282, nx9284, nx9287, nx9289, nx9291, nx9295, nx9297, nx9299, 
      nx9302, nx9304, nx9306, nx9309, nx9311, nx9313, nx9316, nx9318, nx9320, 
      nx9324, nx9326, nx9328, nx9331, nx9333, nx9335, nx9338, nx9340, nx9342, 
      nx9345, nx9347, nx9349, nx9353, nx9355, nx9357, nx9360, nx9362, nx9364, 
      nx9367, nx9369, nx9371, nx9374, nx9376, nx9378, nx9382, nx9384, nx9386, 
      nx9389, nx9391, nx9393, nx9396, nx9398, nx9400, nx9403, nx9405, nx9407, 
      nx9411, nx9413, nx9415, nx9418, nx9420, nx9422, nx9425, nx9427, nx9429, 
      nx9432, nx9434, nx9436, nx9440, nx9442, nx9444, nx9447, nx9449, nx9451, 
      nx9454, nx9456, nx9458, nx9461, nx9463, nx9465, nx9469, nx9471, nx9473, 
      nx9476, nx9478, nx9480, nx9483, nx9485, nx9487, nx9490, nx9492, nx9494, 
      nx9498, nx9500, nx9502, nx9505, nx9507, nx9509, nx9512, nx9514, nx9516, 
      nx9519, nx9521, nx9523, nx9527, nx9529, nx9531, nx9534, nx9536, nx9538, 
      nx9541, nx9543, nx9545, nx9548, nx9550, nx9552, nx9556, nx9558, nx9560, 
      nx9563, nx9565, nx9567, nx9570, nx9572, nx9574, nx9577, nx9579, nx9581, 
      nx9585, nx9587, nx9589, nx9592, nx9594, nx9596, nx9599, nx9601, nx9603, 
      nx9606, nx9608, nx9610, nx9614, nx9616, nx9618, nx9621, nx9623, nx9625, 
      nx9628, nx9630, nx9632, nx9635, nx9637, nx9639, nx9648, nx9650, nx9652, 
      nx9654, nx9656, nx9658, nx9660, nx9662, nx9664, nx9666, nx9668, nx9670, 
      nx9674, nx9676, nx9678, nx9680, nx9682, nx9684, nx9686, nx9688, nx9690, 
      nx9692, nx9694, nx9696, nx9700, nx9702, nx9704, nx9706, nx9708, nx9710, 
      nx9712, nx9714, nx9716, nx9718, nx9720, nx9722, nx9726, nx9728, nx9730, 
      nx9732, nx9734, nx9736, nx9738, nx9740, nx9742, nx9744, nx9746, nx9748, 
      nx9752, nx9754, nx9756, nx9758, nx9760, nx9762, nx9764, nx9766, nx9768, 
      nx9770, nx9772, nx9774, nx9778, nx9780, nx9782, nx9784, nx9786, nx9788, 
      nx9790, nx9792, nx9794, nx9796, nx9798, nx9800, nx9804, nx9806, nx9808, 
      nx9810, nx9812, nx9814, nx9816, nx9818, nx9820, nx9822, nx9824, nx9826, 
      nx9830, nx9832, nx9834, nx9836, nx9838, nx9840, nx9842, nx9844, nx9846, 
      nx9848, nx9850, nx9852, nx9856, nx9858, nx9860, nx9862, nx9864, nx9866, 
      nx9868, nx9870, nx9872, nx9874, nx9876, nx9878, nx9882, nx9884, nx9886, 
      nx9888, nx9890, nx9892, nx9894, nx9896, nx9898, nx9900, nx9902, nx9904, 
      nx9908, nx9910, nx9912, nx9914, nx9916, nx9918, nx9920, nx9922, nx9924, 
      nx9926, nx9928, nx9930, nx9934, nx9936, nx9938, nx9940, nx9942, nx9944, 
      nx9946, nx9948, nx9950, nx9952, nx9954, nx9956, nx9960, nx9962, nx9964, 
      nx9966, nx9968, nx9970, nx9972, nx9974, nx9976, nx9978, nx9980, nx9982, 
      nx9986, nx9988, nx9990, nx9992, nx9994, nx9996, nx9998, nx10000, 
      nx10002, nx10004, nx10006, nx10008, nx10012, nx10014, nx10016, nx10018, 
      nx10020, nx10022, nx10024, nx10026, nx10028, nx10030, nx10032, nx10034, 
      nx10038, nx10040, nx10042, nx10044, nx10046, nx10048, nx10050, nx10052, 
      nx10054, nx10056, nx10058, nx10060, nx10064, nx10066, nx10068, nx10070, 
      nx10072, nx10074, nx10076, nx10078, nx10080, nx10082, nx10084, nx10086, 
      nx10090, nx10092, nx10094, nx10096, nx10098, nx10100, nx10102, nx10104, 
      nx10106, nx10108, nx10110, nx10112, nx10116, nx10118, nx10120, nx10122, 
      nx10124, nx10126, nx10128, nx10130, nx10132, nx10134, nx10136, nx10138, 
      nx10142, nx10144, nx10146, nx10148, nx10150, nx10152, nx10154, nx10156, 
      nx10158, nx10160, nx10162, nx10164, nx10168, nx10170, nx10172, nx10174, 
      nx10176, nx10178, nx10180, nx10182, nx10184, nx10186, nx10188, nx10190, 
      nx10194, nx10196, nx10198, nx10200, nx10202, nx10204, nx10206, nx10208, 
      nx10210, nx10212, nx10214, nx10216, nx10220, nx10222, nx10224, nx10226, 
      nx10228, nx10230, nx10232, nx10234, nx10236, nx10238, nx10240, nx10242, 
      nx10246, nx10248, nx10250, nx10252, nx10254, nx10256, nx10258, nx10260, 
      nx10262, nx10264, nx10266, nx10268, nx10272, nx10274, nx10276, nx10278, 
      nx10280, nx10282, nx10284, nx10286, nx10288, nx10290, nx10292, nx10294, 
      nx10298, nx10300, nx10302, nx10304, nx10306, nx10308, nx10310, nx10312, 
      nx10314, nx10316, nx10318, nx10320, nx10324, nx10326, nx10328, nx10330, 
      nx10332, nx10334, nx10336, nx10338, nx10340, nx10342, nx10344, nx10346, 
      nx10350, nx10352, nx10354, nx10356, nx10358, nx10360, nx10362, nx10364, 
      nx10366, nx10368, nx10370, nx10372, nx10374, nx10376, nx10378, nx10380, 
      nx10382, nx10384, nx10386, nx10388, nx10390, nx10392, nx10394, nx10396, 
      nx10398, nx10400, nx10402, nx10404, nx10406, nx10408, nx10410, nx10412, 
      nx10414, nx10416, nx10418, nx10420, nx10422, nx10424, nx10426, nx10428, 
      nx10430, nx10432, nx10434, nx10436, nx10438, nx10440, nx10442, nx10444, 
      nx10446, nx10448, nx10450, nx10452, nx10454, nx10456, nx10458, nx10460, 
      nx10462, nx10464, nx10466, nx10468, nx10470, nx10472, nx10474, nx10476, 
      nx10478, nx10480, nx10482, nx10484, nx10486, nx10488, nx10494, nx10496, 
      nx10498, nx10500, nx10502, nx10504, nx10506, nx10508, nx10510, nx10512, 
      nx10514, nx10516, nx10518, nx10520, nx10522, nx10524, nx10526, nx10528, 
      nx10530, nx10532, nx10534, nx10536, nx10538, nx10540, nx10542, nx10544, 
      nx10546, nx10548, nx10550, nx10552, nx10554, nx10556, nx10558, nx10560, 
      nx10562, nx10564, nx10566, nx10568, nx10570, nx10572, nx10574, nx10576, 
      nx10578, nx10580, nx10582, nx10584, nx10586, nx10588, nx10590, nx10592, 
      nx10594, nx10596, nx10598, nx10600, nx10602, nx10604, nx10606, nx10608, 
      nx10610, nx10612, nx10614, nx10616, nx10618, nx10620, nx10622, nx10624, 
      nx10626, nx10628, nx10630, nx10632, nx10634, nx10636, nx10638, nx10640, 
      nx10642, nx10644, nx10646, nx10648, nx10650, nx10652, nx10654, nx10656, 
      nx10658, nx10660, nx10662, nx10664, nx10666, nx10668, nx10690, nx10692, 
      nx10694, nx10696, nx10698, nx10700, nx10702, nx10704, nx10706, nx10708, 
      nx10710, nx10712, nx10714, nx10716, nx10718, nx10720, nx10722, nx10724, 
      nx10726, nx10728, nx10730, nx10732, nx10734, nx10736, nx10742, nx10744, 
      nx10746, nx10748: std_logic ;

begin
   gen_queues_0_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_0_0_15, q_0_14=>que_out_0_0_14, q_0_13=>
      que_out_0_0_13, q_0_12=>que_out_0_0_12, q_0_11=>que_out_0_0_11, q_0_10
      =>que_out_0_0_10, q_0_9=>que_out_0_0_9, q_0_8=>que_out_0_0_8, q_0_7=>
      que_out_0_0_7, q_0_6=>que_out_0_0_6, q_0_5=>que_out_0_0_5, q_0_4=>
      que_out_0_0_4, q_0_3=>que_out_0_0_3, q_0_2=>que_out_0_0_2, q_0_1=>
      que_out_0_0_1, q_0_0=>que_out_0_0_0, q_1_15=>que_out_0_1_15, q_1_14=>
      que_out_0_1_14, q_1_13=>que_out_0_1_13, q_1_12=>que_out_0_1_12, q_1_11
      =>que_out_0_1_11, q_1_10=>que_out_0_1_10, q_1_9=>que_out_0_1_9, q_1_8
      =>que_out_0_1_8, q_1_7=>que_out_0_1_7, q_1_6=>que_out_0_1_6, q_1_5=>
      que_out_0_1_5, q_1_4=>que_out_0_1_4, q_1_3=>que_out_0_1_3, q_1_2=>
      que_out_0_1_2, q_1_1=>que_out_0_1_1, q_1_0=>que_out_0_1_0, q_2_15=>
      que_out_0_2_15, q_2_14=>que_out_0_2_14, q_2_13=>que_out_0_2_13, q_2_12
      =>que_out_0_2_12, q_2_11=>que_out_0_2_11, q_2_10=>que_out_0_2_10, 
      q_2_9=>que_out_0_2_9, q_2_8=>que_out_0_2_8, q_2_7=>que_out_0_2_7, 
      q_2_6=>que_out_0_2_6, q_2_5=>que_out_0_2_5, q_2_4=>que_out_0_2_4, 
      q_2_3=>que_out_0_2_3, q_2_2=>que_out_0_2_2, q_2_1=>que_out_0_2_1, 
      q_2_0=>que_out_0_2_0, q_3_15=>que_out_0_3_15, q_3_14=>que_out_0_3_14, 
      q_3_13=>que_out_0_3_13, q_3_12=>que_out_0_3_12, q_3_11=>que_out_0_3_11, 
      q_3_10=>que_out_0_3_10, q_3_9=>que_out_0_3_9, q_3_8=>que_out_0_3_8, 
      q_3_7=>que_out_0_3_7, q_3_6=>que_out_0_3_6, q_3_5=>que_out_0_3_5, 
      q_3_4=>que_out_0_3_4, q_3_3=>que_out_0_3_3, q_3_2=>que_out_0_3_2, 
      q_3_1=>que_out_0_3_1, q_3_0=>que_out_0_3_0, q_4_15=>que_out_0_4_15, 
      q_4_14=>que_out_0_4_14, q_4_13=>que_out_0_4_13, q_4_12=>que_out_0_4_12, 
      q_4_11=>que_out_0_4_11, q_4_10=>que_out_0_4_10, q_4_9=>que_out_0_4_9, 
      q_4_8=>que_out_0_4_8, q_4_7=>que_out_0_4_7, q_4_6=>que_out_0_4_6, 
      q_4_5=>que_out_0_4_5, q_4_4=>que_out_0_4_4, q_4_3=>que_out_0_4_3, 
      q_4_2=>que_out_0_4_2, q_4_1=>que_out_0_4_1, q_4_0=>que_out_0_4_0, clk
      =>nx10714, load=>sel_que_0, reset=>nx10690);
   gen_queues_1_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_1_0_15, q_0_14=>que_out_1_0_14, q_0_13=>
      que_out_1_0_13, q_0_12=>que_out_1_0_12, q_0_11=>que_out_1_0_11, q_0_10
      =>que_out_1_0_10, q_0_9=>que_out_1_0_9, q_0_8=>que_out_1_0_8, q_0_7=>
      que_out_1_0_7, q_0_6=>que_out_1_0_6, q_0_5=>que_out_1_0_5, q_0_4=>
      que_out_1_0_4, q_0_3=>que_out_1_0_3, q_0_2=>que_out_1_0_2, q_0_1=>
      que_out_1_0_1, q_0_0=>que_out_1_0_0, q_1_15=>que_out_1_1_15, q_1_14=>
      que_out_1_1_14, q_1_13=>que_out_1_1_13, q_1_12=>que_out_1_1_12, q_1_11
      =>que_out_1_1_11, q_1_10=>que_out_1_1_10, q_1_9=>que_out_1_1_9, q_1_8
      =>que_out_1_1_8, q_1_7=>que_out_1_1_7, q_1_6=>que_out_1_1_6, q_1_5=>
      que_out_1_1_5, q_1_4=>que_out_1_1_4, q_1_3=>que_out_1_1_3, q_1_2=>
      que_out_1_1_2, q_1_1=>que_out_1_1_1, q_1_0=>que_out_1_1_0, q_2_15=>
      que_out_1_2_15, q_2_14=>que_out_1_2_14, q_2_13=>que_out_1_2_13, q_2_12
      =>que_out_1_2_12, q_2_11=>que_out_1_2_11, q_2_10=>que_out_1_2_10, 
      q_2_9=>que_out_1_2_9, q_2_8=>que_out_1_2_8, q_2_7=>que_out_1_2_7, 
      q_2_6=>que_out_1_2_6, q_2_5=>que_out_1_2_5, q_2_4=>que_out_1_2_4, 
      q_2_3=>que_out_1_2_3, q_2_2=>que_out_1_2_2, q_2_1=>que_out_1_2_1, 
      q_2_0=>que_out_1_2_0, q_3_15=>que_out_1_3_15, q_3_14=>que_out_1_3_14, 
      q_3_13=>que_out_1_3_13, q_3_12=>que_out_1_3_12, q_3_11=>que_out_1_3_11, 
      q_3_10=>que_out_1_3_10, q_3_9=>que_out_1_3_9, q_3_8=>que_out_1_3_8, 
      q_3_7=>que_out_1_3_7, q_3_6=>que_out_1_3_6, q_3_5=>que_out_1_3_5, 
      q_3_4=>que_out_1_3_4, q_3_3=>que_out_1_3_3, q_3_2=>que_out_1_3_2, 
      q_3_1=>que_out_1_3_1, q_3_0=>que_out_1_3_0, q_4_15=>que_out_1_4_15, 
      q_4_14=>que_out_1_4_14, q_4_13=>que_out_1_4_13, q_4_12=>que_out_1_4_12, 
      q_4_11=>que_out_1_4_11, q_4_10=>que_out_1_4_10, q_4_9=>que_out_1_4_9, 
      q_4_8=>que_out_1_4_8, q_4_7=>que_out_1_4_7, q_4_6=>que_out_1_4_6, 
      q_4_5=>que_out_1_4_5, q_4_4=>que_out_1_4_4, q_4_3=>que_out_1_4_3, 
      q_4_2=>que_out_1_4_2, q_4_1=>que_out_1_4_1, q_4_0=>que_out_1_4_0, clk
      =>nx10714, load=>sel_que_1, reset=>nx10690);
   gen_queues_2_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_2_0_15, q_0_14=>que_out_2_0_14, q_0_13=>
      que_out_2_0_13, q_0_12=>que_out_2_0_12, q_0_11=>que_out_2_0_11, q_0_10
      =>que_out_2_0_10, q_0_9=>que_out_2_0_9, q_0_8=>que_out_2_0_8, q_0_7=>
      que_out_2_0_7, q_0_6=>que_out_2_0_6, q_0_5=>que_out_2_0_5, q_0_4=>
      que_out_2_0_4, q_0_3=>que_out_2_0_3, q_0_2=>que_out_2_0_2, q_0_1=>
      que_out_2_0_1, q_0_0=>que_out_2_0_0, q_1_15=>que_out_2_1_15, q_1_14=>
      que_out_2_1_14, q_1_13=>que_out_2_1_13, q_1_12=>que_out_2_1_12, q_1_11
      =>que_out_2_1_11, q_1_10=>que_out_2_1_10, q_1_9=>que_out_2_1_9, q_1_8
      =>que_out_2_1_8, q_1_7=>que_out_2_1_7, q_1_6=>que_out_2_1_6, q_1_5=>
      que_out_2_1_5, q_1_4=>que_out_2_1_4, q_1_3=>que_out_2_1_3, q_1_2=>
      que_out_2_1_2, q_1_1=>que_out_2_1_1, q_1_0=>que_out_2_1_0, q_2_15=>
      que_out_2_2_15, q_2_14=>que_out_2_2_14, q_2_13=>que_out_2_2_13, q_2_12
      =>que_out_2_2_12, q_2_11=>que_out_2_2_11, q_2_10=>que_out_2_2_10, 
      q_2_9=>que_out_2_2_9, q_2_8=>que_out_2_2_8, q_2_7=>que_out_2_2_7, 
      q_2_6=>que_out_2_2_6, q_2_5=>que_out_2_2_5, q_2_4=>que_out_2_2_4, 
      q_2_3=>que_out_2_2_3, q_2_2=>que_out_2_2_2, q_2_1=>que_out_2_2_1, 
      q_2_0=>que_out_2_2_0, q_3_15=>que_out_2_3_15, q_3_14=>que_out_2_3_14, 
      q_3_13=>que_out_2_3_13, q_3_12=>que_out_2_3_12, q_3_11=>que_out_2_3_11, 
      q_3_10=>que_out_2_3_10, q_3_9=>que_out_2_3_9, q_3_8=>que_out_2_3_8, 
      q_3_7=>que_out_2_3_7, q_3_6=>que_out_2_3_6, q_3_5=>que_out_2_3_5, 
      q_3_4=>que_out_2_3_4, q_3_3=>que_out_2_3_3, q_3_2=>que_out_2_3_2, 
      q_3_1=>que_out_2_3_1, q_3_0=>que_out_2_3_0, q_4_15=>que_out_2_4_15, 
      q_4_14=>que_out_2_4_14, q_4_13=>que_out_2_4_13, q_4_12=>que_out_2_4_12, 
      q_4_11=>que_out_2_4_11, q_4_10=>que_out_2_4_10, q_4_9=>que_out_2_4_9, 
      q_4_8=>que_out_2_4_8, q_4_7=>que_out_2_4_7, q_4_6=>que_out_2_4_6, 
      q_4_5=>que_out_2_4_5, q_4_4=>que_out_2_4_4, q_4_3=>que_out_2_4_3, 
      q_4_2=>que_out_2_4_2, q_4_1=>que_out_2_4_1, q_4_0=>que_out_2_4_0, clk
      =>nx10714, load=>sel_que_2, reset=>nx10690);
   gen_queues_3_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_3_0_15, q_0_14=>que_out_3_0_14, q_0_13=>
      que_out_3_0_13, q_0_12=>que_out_3_0_12, q_0_11=>que_out_3_0_11, q_0_10
      =>que_out_3_0_10, q_0_9=>que_out_3_0_9, q_0_8=>que_out_3_0_8, q_0_7=>
      que_out_3_0_7, q_0_6=>que_out_3_0_6, q_0_5=>que_out_3_0_5, q_0_4=>
      que_out_3_0_4, q_0_3=>que_out_3_0_3, q_0_2=>que_out_3_0_2, q_0_1=>
      que_out_3_0_1, q_0_0=>que_out_3_0_0, q_1_15=>que_out_3_1_15, q_1_14=>
      que_out_3_1_14, q_1_13=>que_out_3_1_13, q_1_12=>que_out_3_1_12, q_1_11
      =>que_out_3_1_11, q_1_10=>que_out_3_1_10, q_1_9=>que_out_3_1_9, q_1_8
      =>que_out_3_1_8, q_1_7=>que_out_3_1_7, q_1_6=>que_out_3_1_6, q_1_5=>
      que_out_3_1_5, q_1_4=>que_out_3_1_4, q_1_3=>que_out_3_1_3, q_1_2=>
      que_out_3_1_2, q_1_1=>que_out_3_1_1, q_1_0=>que_out_3_1_0, q_2_15=>
      que_out_3_2_15, q_2_14=>que_out_3_2_14, q_2_13=>que_out_3_2_13, q_2_12
      =>que_out_3_2_12, q_2_11=>que_out_3_2_11, q_2_10=>que_out_3_2_10, 
      q_2_9=>que_out_3_2_9, q_2_8=>que_out_3_2_8, q_2_7=>que_out_3_2_7, 
      q_2_6=>que_out_3_2_6, q_2_5=>que_out_3_2_5, q_2_4=>que_out_3_2_4, 
      q_2_3=>que_out_3_2_3, q_2_2=>que_out_3_2_2, q_2_1=>que_out_3_2_1, 
      q_2_0=>que_out_3_2_0, q_3_15=>que_out_3_3_15, q_3_14=>que_out_3_3_14, 
      q_3_13=>que_out_3_3_13, q_3_12=>que_out_3_3_12, q_3_11=>que_out_3_3_11, 
      q_3_10=>que_out_3_3_10, q_3_9=>que_out_3_3_9, q_3_8=>que_out_3_3_8, 
      q_3_7=>que_out_3_3_7, q_3_6=>que_out_3_3_6, q_3_5=>que_out_3_3_5, 
      q_3_4=>que_out_3_3_4, q_3_3=>que_out_3_3_3, q_3_2=>que_out_3_3_2, 
      q_3_1=>que_out_3_3_1, q_3_0=>que_out_3_3_0, q_4_15=>que_out_3_4_15, 
      q_4_14=>que_out_3_4_14, q_4_13=>que_out_3_4_13, q_4_12=>que_out_3_4_12, 
      q_4_11=>que_out_3_4_11, q_4_10=>que_out_3_4_10, q_4_9=>que_out_3_4_9, 
      q_4_8=>que_out_3_4_8, q_4_7=>que_out_3_4_7, q_4_6=>que_out_3_4_6, 
      q_4_5=>que_out_3_4_5, q_4_4=>que_out_3_4_4, q_4_3=>que_out_3_4_3, 
      q_4_2=>que_out_3_4_2, q_4_1=>que_out_3_4_1, q_4_0=>que_out_3_4_0, clk
      =>nx10716, load=>sel_que_3, reset=>nx10692);
   gen_queues_4_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_4_0_15, q_0_14=>que_out_4_0_14, q_0_13=>
      que_out_4_0_13, q_0_12=>que_out_4_0_12, q_0_11=>que_out_4_0_11, q_0_10
      =>que_out_4_0_10, q_0_9=>que_out_4_0_9, q_0_8=>que_out_4_0_8, q_0_7=>
      que_out_4_0_7, q_0_6=>que_out_4_0_6, q_0_5=>que_out_4_0_5, q_0_4=>
      que_out_4_0_4, q_0_3=>que_out_4_0_3, q_0_2=>que_out_4_0_2, q_0_1=>
      que_out_4_0_1, q_0_0=>que_out_4_0_0, q_1_15=>que_out_4_1_15, q_1_14=>
      que_out_4_1_14, q_1_13=>que_out_4_1_13, q_1_12=>que_out_4_1_12, q_1_11
      =>que_out_4_1_11, q_1_10=>que_out_4_1_10, q_1_9=>que_out_4_1_9, q_1_8
      =>que_out_4_1_8, q_1_7=>que_out_4_1_7, q_1_6=>que_out_4_1_6, q_1_5=>
      que_out_4_1_5, q_1_4=>que_out_4_1_4, q_1_3=>que_out_4_1_3, q_1_2=>
      que_out_4_1_2, q_1_1=>que_out_4_1_1, q_1_0=>que_out_4_1_0, q_2_15=>
      que_out_4_2_15, q_2_14=>que_out_4_2_14, q_2_13=>que_out_4_2_13, q_2_12
      =>que_out_4_2_12, q_2_11=>que_out_4_2_11, q_2_10=>que_out_4_2_10, 
      q_2_9=>que_out_4_2_9, q_2_8=>que_out_4_2_8, q_2_7=>que_out_4_2_7, 
      q_2_6=>que_out_4_2_6, q_2_5=>que_out_4_2_5, q_2_4=>que_out_4_2_4, 
      q_2_3=>que_out_4_2_3, q_2_2=>que_out_4_2_2, q_2_1=>que_out_4_2_1, 
      q_2_0=>que_out_4_2_0, q_3_15=>que_out_4_3_15, q_3_14=>que_out_4_3_14, 
      q_3_13=>que_out_4_3_13, q_3_12=>que_out_4_3_12, q_3_11=>que_out_4_3_11, 
      q_3_10=>que_out_4_3_10, q_3_9=>que_out_4_3_9, q_3_8=>que_out_4_3_8, 
      q_3_7=>que_out_4_3_7, q_3_6=>que_out_4_3_6, q_3_5=>que_out_4_3_5, 
      q_3_4=>que_out_4_3_4, q_3_3=>que_out_4_3_3, q_3_2=>que_out_4_3_2, 
      q_3_1=>que_out_4_3_1, q_3_0=>que_out_4_3_0, q_4_15=>que_out_4_4_15, 
      q_4_14=>que_out_4_4_14, q_4_13=>que_out_4_4_13, q_4_12=>que_out_4_4_12, 
      q_4_11=>que_out_4_4_11, q_4_10=>que_out_4_4_10, q_4_9=>que_out_4_4_9, 
      q_4_8=>que_out_4_4_8, q_4_7=>que_out_4_4_7, q_4_6=>que_out_4_4_6, 
      q_4_5=>que_out_4_4_5, q_4_4=>que_out_4_4_4, q_4_3=>que_out_4_4_3, 
      q_4_2=>que_out_4_4_2, q_4_1=>que_out_4_4_1, q_4_0=>que_out_4_4_0, clk
      =>nx10716, load=>sel_que_4, reset=>nx10692);
   gen_queues_5_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_5_0_15, q_0_14=>que_out_5_0_14, q_0_13=>
      que_out_5_0_13, q_0_12=>que_out_5_0_12, q_0_11=>que_out_5_0_11, q_0_10
      =>que_out_5_0_10, q_0_9=>que_out_5_0_9, q_0_8=>que_out_5_0_8, q_0_7=>
      que_out_5_0_7, q_0_6=>que_out_5_0_6, q_0_5=>que_out_5_0_5, q_0_4=>
      que_out_5_0_4, q_0_3=>que_out_5_0_3, q_0_2=>que_out_5_0_2, q_0_1=>
      que_out_5_0_1, q_0_0=>que_out_5_0_0, q_1_15=>que_out_5_1_15, q_1_14=>
      que_out_5_1_14, q_1_13=>que_out_5_1_13, q_1_12=>que_out_5_1_12, q_1_11
      =>que_out_5_1_11, q_1_10=>que_out_5_1_10, q_1_9=>que_out_5_1_9, q_1_8
      =>que_out_5_1_8, q_1_7=>que_out_5_1_7, q_1_6=>que_out_5_1_6, q_1_5=>
      que_out_5_1_5, q_1_4=>que_out_5_1_4, q_1_3=>que_out_5_1_3, q_1_2=>
      que_out_5_1_2, q_1_1=>que_out_5_1_1, q_1_0=>que_out_5_1_0, q_2_15=>
      que_out_5_2_15, q_2_14=>que_out_5_2_14, q_2_13=>que_out_5_2_13, q_2_12
      =>que_out_5_2_12, q_2_11=>que_out_5_2_11, q_2_10=>que_out_5_2_10, 
      q_2_9=>que_out_5_2_9, q_2_8=>que_out_5_2_8, q_2_7=>que_out_5_2_7, 
      q_2_6=>que_out_5_2_6, q_2_5=>que_out_5_2_5, q_2_4=>que_out_5_2_4, 
      q_2_3=>que_out_5_2_3, q_2_2=>que_out_5_2_2, q_2_1=>que_out_5_2_1, 
      q_2_0=>que_out_5_2_0, q_3_15=>que_out_5_3_15, q_3_14=>que_out_5_3_14, 
      q_3_13=>que_out_5_3_13, q_3_12=>que_out_5_3_12, q_3_11=>que_out_5_3_11, 
      q_3_10=>que_out_5_3_10, q_3_9=>que_out_5_3_9, q_3_8=>que_out_5_3_8, 
      q_3_7=>que_out_5_3_7, q_3_6=>que_out_5_3_6, q_3_5=>que_out_5_3_5, 
      q_3_4=>que_out_5_3_4, q_3_3=>que_out_5_3_3, q_3_2=>que_out_5_3_2, 
      q_3_1=>que_out_5_3_1, q_3_0=>que_out_5_3_0, q_4_15=>que_out_5_4_15, 
      q_4_14=>que_out_5_4_14, q_4_13=>que_out_5_4_13, q_4_12=>que_out_5_4_12, 
      q_4_11=>que_out_5_4_11, q_4_10=>que_out_5_4_10, q_4_9=>que_out_5_4_9, 
      q_4_8=>que_out_5_4_8, q_4_7=>que_out_5_4_7, q_4_6=>que_out_5_4_6, 
      q_4_5=>que_out_5_4_5, q_4_4=>que_out_5_4_4, q_4_3=>que_out_5_4_3, 
      q_4_2=>que_out_5_4_2, q_4_1=>que_out_5_4_1, q_4_0=>que_out_5_4_0, clk
      =>nx10716, load=>sel_que_5, reset=>nx10692);
   gen_queues_6_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_6_0_15, q_0_14=>que_out_6_0_14, q_0_13=>
      que_out_6_0_13, q_0_12=>que_out_6_0_12, q_0_11=>que_out_6_0_11, q_0_10
      =>que_out_6_0_10, q_0_9=>que_out_6_0_9, q_0_8=>que_out_6_0_8, q_0_7=>
      que_out_6_0_7, q_0_6=>que_out_6_0_6, q_0_5=>que_out_6_0_5, q_0_4=>
      que_out_6_0_4, q_0_3=>que_out_6_0_3, q_0_2=>que_out_6_0_2, q_0_1=>
      que_out_6_0_1, q_0_0=>que_out_6_0_0, q_1_15=>que_out_6_1_15, q_1_14=>
      que_out_6_1_14, q_1_13=>que_out_6_1_13, q_1_12=>que_out_6_1_12, q_1_11
      =>que_out_6_1_11, q_1_10=>que_out_6_1_10, q_1_9=>que_out_6_1_9, q_1_8
      =>que_out_6_1_8, q_1_7=>que_out_6_1_7, q_1_6=>que_out_6_1_6, q_1_5=>
      que_out_6_1_5, q_1_4=>que_out_6_1_4, q_1_3=>que_out_6_1_3, q_1_2=>
      que_out_6_1_2, q_1_1=>que_out_6_1_1, q_1_0=>que_out_6_1_0, q_2_15=>
      que_out_6_2_15, q_2_14=>que_out_6_2_14, q_2_13=>que_out_6_2_13, q_2_12
      =>que_out_6_2_12, q_2_11=>que_out_6_2_11, q_2_10=>que_out_6_2_10, 
      q_2_9=>que_out_6_2_9, q_2_8=>que_out_6_2_8, q_2_7=>que_out_6_2_7, 
      q_2_6=>que_out_6_2_6, q_2_5=>que_out_6_2_5, q_2_4=>que_out_6_2_4, 
      q_2_3=>que_out_6_2_3, q_2_2=>que_out_6_2_2, q_2_1=>que_out_6_2_1, 
      q_2_0=>que_out_6_2_0, q_3_15=>que_out_6_3_15, q_3_14=>que_out_6_3_14, 
      q_3_13=>que_out_6_3_13, q_3_12=>que_out_6_3_12, q_3_11=>que_out_6_3_11, 
      q_3_10=>que_out_6_3_10, q_3_9=>que_out_6_3_9, q_3_8=>que_out_6_3_8, 
      q_3_7=>que_out_6_3_7, q_3_6=>que_out_6_3_6, q_3_5=>que_out_6_3_5, 
      q_3_4=>que_out_6_3_4, q_3_3=>que_out_6_3_3, q_3_2=>que_out_6_3_2, 
      q_3_1=>que_out_6_3_1, q_3_0=>que_out_6_3_0, q_4_15=>que_out_6_4_15, 
      q_4_14=>que_out_6_4_14, q_4_13=>que_out_6_4_13, q_4_12=>que_out_6_4_12, 
      q_4_11=>que_out_6_4_11, q_4_10=>que_out_6_4_10, q_4_9=>que_out_6_4_9, 
      q_4_8=>que_out_6_4_8, q_4_7=>que_out_6_4_7, q_4_6=>que_out_6_4_6, 
      q_4_5=>que_out_6_4_5, q_4_4=>que_out_6_4_4, q_4_3=>que_out_6_4_3, 
      q_4_2=>que_out_6_4_2, q_4_1=>que_out_6_4_1, q_4_0=>que_out_6_4_0, clk
      =>nx10718, load=>sel_que_6, reset=>nx10694);
   gen_queues_7_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_7_0_15, q_0_14=>que_out_7_0_14, q_0_13=>
      que_out_7_0_13, q_0_12=>que_out_7_0_12, q_0_11=>que_out_7_0_11, q_0_10
      =>que_out_7_0_10, q_0_9=>que_out_7_0_9, q_0_8=>que_out_7_0_8, q_0_7=>
      que_out_7_0_7, q_0_6=>que_out_7_0_6, q_0_5=>que_out_7_0_5, q_0_4=>
      que_out_7_0_4, q_0_3=>que_out_7_0_3, q_0_2=>que_out_7_0_2, q_0_1=>
      que_out_7_0_1, q_0_0=>que_out_7_0_0, q_1_15=>que_out_7_1_15, q_1_14=>
      que_out_7_1_14, q_1_13=>que_out_7_1_13, q_1_12=>que_out_7_1_12, q_1_11
      =>que_out_7_1_11, q_1_10=>que_out_7_1_10, q_1_9=>que_out_7_1_9, q_1_8
      =>que_out_7_1_8, q_1_7=>que_out_7_1_7, q_1_6=>que_out_7_1_6, q_1_5=>
      que_out_7_1_5, q_1_4=>que_out_7_1_4, q_1_3=>que_out_7_1_3, q_1_2=>
      que_out_7_1_2, q_1_1=>que_out_7_1_1, q_1_0=>que_out_7_1_0, q_2_15=>
      que_out_7_2_15, q_2_14=>que_out_7_2_14, q_2_13=>que_out_7_2_13, q_2_12
      =>que_out_7_2_12, q_2_11=>que_out_7_2_11, q_2_10=>que_out_7_2_10, 
      q_2_9=>que_out_7_2_9, q_2_8=>que_out_7_2_8, q_2_7=>que_out_7_2_7, 
      q_2_6=>que_out_7_2_6, q_2_5=>que_out_7_2_5, q_2_4=>que_out_7_2_4, 
      q_2_3=>que_out_7_2_3, q_2_2=>que_out_7_2_2, q_2_1=>que_out_7_2_1, 
      q_2_0=>que_out_7_2_0, q_3_15=>que_out_7_3_15, q_3_14=>que_out_7_3_14, 
      q_3_13=>que_out_7_3_13, q_3_12=>que_out_7_3_12, q_3_11=>que_out_7_3_11, 
      q_3_10=>que_out_7_3_10, q_3_9=>que_out_7_3_9, q_3_8=>que_out_7_3_8, 
      q_3_7=>que_out_7_3_7, q_3_6=>que_out_7_3_6, q_3_5=>que_out_7_3_5, 
      q_3_4=>que_out_7_3_4, q_3_3=>que_out_7_3_3, q_3_2=>que_out_7_3_2, 
      q_3_1=>que_out_7_3_1, q_3_0=>que_out_7_3_0, q_4_15=>que_out_7_4_15, 
      q_4_14=>que_out_7_4_14, q_4_13=>que_out_7_4_13, q_4_12=>que_out_7_4_12, 
      q_4_11=>que_out_7_4_11, q_4_10=>que_out_7_4_10, q_4_9=>que_out_7_4_9, 
      q_4_8=>que_out_7_4_8, q_4_7=>que_out_7_4_7, q_4_6=>que_out_7_4_6, 
      q_4_5=>que_out_7_4_5, q_4_4=>que_out_7_4_4, q_4_3=>que_out_7_4_3, 
      q_4_2=>que_out_7_4_2, q_4_1=>que_out_7_4_1, q_4_0=>que_out_7_4_0, clk
      =>nx10720, load=>sel_que_7, reset=>nx10696);
   gen_queues_8_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_8_0_15, q_0_14=>que_out_8_0_14, q_0_13=>
      que_out_8_0_13, q_0_12=>que_out_8_0_12, q_0_11=>que_out_8_0_11, q_0_10
      =>que_out_8_0_10, q_0_9=>que_out_8_0_9, q_0_8=>que_out_8_0_8, q_0_7=>
      que_out_8_0_7, q_0_6=>que_out_8_0_6, q_0_5=>que_out_8_0_5, q_0_4=>
      que_out_8_0_4, q_0_3=>que_out_8_0_3, q_0_2=>que_out_8_0_2, q_0_1=>
      que_out_8_0_1, q_0_0=>que_out_8_0_0, q_1_15=>que_out_8_1_15, q_1_14=>
      que_out_8_1_14, q_1_13=>que_out_8_1_13, q_1_12=>que_out_8_1_12, q_1_11
      =>que_out_8_1_11, q_1_10=>que_out_8_1_10, q_1_9=>que_out_8_1_9, q_1_8
      =>que_out_8_1_8, q_1_7=>que_out_8_1_7, q_1_6=>que_out_8_1_6, q_1_5=>
      que_out_8_1_5, q_1_4=>que_out_8_1_4, q_1_3=>que_out_8_1_3, q_1_2=>
      que_out_8_1_2, q_1_1=>que_out_8_1_1, q_1_0=>que_out_8_1_0, q_2_15=>
      que_out_8_2_15, q_2_14=>que_out_8_2_14, q_2_13=>que_out_8_2_13, q_2_12
      =>que_out_8_2_12, q_2_11=>que_out_8_2_11, q_2_10=>que_out_8_2_10, 
      q_2_9=>que_out_8_2_9, q_2_8=>que_out_8_2_8, q_2_7=>que_out_8_2_7, 
      q_2_6=>que_out_8_2_6, q_2_5=>que_out_8_2_5, q_2_4=>que_out_8_2_4, 
      q_2_3=>que_out_8_2_3, q_2_2=>que_out_8_2_2, q_2_1=>que_out_8_2_1, 
      q_2_0=>que_out_8_2_0, q_3_15=>que_out_8_3_15, q_3_14=>que_out_8_3_14, 
      q_3_13=>que_out_8_3_13, q_3_12=>que_out_8_3_12, q_3_11=>que_out_8_3_11, 
      q_3_10=>que_out_8_3_10, q_3_9=>que_out_8_3_9, q_3_8=>que_out_8_3_8, 
      q_3_7=>que_out_8_3_7, q_3_6=>que_out_8_3_6, q_3_5=>que_out_8_3_5, 
      q_3_4=>que_out_8_3_4, q_3_3=>que_out_8_3_3, q_3_2=>que_out_8_3_2, 
      q_3_1=>que_out_8_3_1, q_3_0=>que_out_8_3_0, q_4_15=>que_out_8_4_15, 
      q_4_14=>que_out_8_4_14, q_4_13=>que_out_8_4_13, q_4_12=>que_out_8_4_12, 
      q_4_11=>que_out_8_4_11, q_4_10=>que_out_8_4_10, q_4_9=>que_out_8_4_9, 
      q_4_8=>que_out_8_4_8, q_4_7=>que_out_8_4_7, q_4_6=>que_out_8_4_6, 
      q_4_5=>que_out_8_4_5, q_4_4=>que_out_8_4_4, q_4_3=>que_out_8_4_3, 
      q_4_2=>que_out_8_4_2, q_4_1=>que_out_8_4_1, q_4_0=>que_out_8_4_0, clk
      =>nx10720, load=>sel_que_8, reset=>nx10696);
   gen_queues_9_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_9_0_15, q_0_14=>que_out_9_0_14, q_0_13=>
      que_out_9_0_13, q_0_12=>que_out_9_0_12, q_0_11=>que_out_9_0_11, q_0_10
      =>que_out_9_0_10, q_0_9=>que_out_9_0_9, q_0_8=>que_out_9_0_8, q_0_7=>
      que_out_9_0_7, q_0_6=>que_out_9_0_6, q_0_5=>que_out_9_0_5, q_0_4=>
      que_out_9_0_4, q_0_3=>que_out_9_0_3, q_0_2=>que_out_9_0_2, q_0_1=>
      que_out_9_0_1, q_0_0=>que_out_9_0_0, q_1_15=>que_out_9_1_15, q_1_14=>
      que_out_9_1_14, q_1_13=>que_out_9_1_13, q_1_12=>que_out_9_1_12, q_1_11
      =>que_out_9_1_11, q_1_10=>que_out_9_1_10, q_1_9=>que_out_9_1_9, q_1_8
      =>que_out_9_1_8, q_1_7=>que_out_9_1_7, q_1_6=>que_out_9_1_6, q_1_5=>
      que_out_9_1_5, q_1_4=>que_out_9_1_4, q_1_3=>que_out_9_1_3, q_1_2=>
      que_out_9_1_2, q_1_1=>que_out_9_1_1, q_1_0=>que_out_9_1_0, q_2_15=>
      que_out_9_2_15, q_2_14=>que_out_9_2_14, q_2_13=>que_out_9_2_13, q_2_12
      =>que_out_9_2_12, q_2_11=>que_out_9_2_11, q_2_10=>que_out_9_2_10, 
      q_2_9=>que_out_9_2_9, q_2_8=>que_out_9_2_8, q_2_7=>que_out_9_2_7, 
      q_2_6=>que_out_9_2_6, q_2_5=>que_out_9_2_5, q_2_4=>que_out_9_2_4, 
      q_2_3=>que_out_9_2_3, q_2_2=>que_out_9_2_2, q_2_1=>que_out_9_2_1, 
      q_2_0=>que_out_9_2_0, q_3_15=>que_out_9_3_15, q_3_14=>que_out_9_3_14, 
      q_3_13=>que_out_9_3_13, q_3_12=>que_out_9_3_12, q_3_11=>que_out_9_3_11, 
      q_3_10=>que_out_9_3_10, q_3_9=>que_out_9_3_9, q_3_8=>que_out_9_3_8, 
      q_3_7=>que_out_9_3_7, q_3_6=>que_out_9_3_6, q_3_5=>que_out_9_3_5, 
      q_3_4=>que_out_9_3_4, q_3_3=>que_out_9_3_3, q_3_2=>que_out_9_3_2, 
      q_3_1=>que_out_9_3_1, q_3_0=>que_out_9_3_0, q_4_15=>que_out_9_4_15, 
      q_4_14=>que_out_9_4_14, q_4_13=>que_out_9_4_13, q_4_12=>que_out_9_4_12, 
      q_4_11=>que_out_9_4_11, q_4_10=>que_out_9_4_10, q_4_9=>que_out_9_4_9, 
      q_4_8=>que_out_9_4_8, q_4_7=>que_out_9_4_7, q_4_6=>que_out_9_4_6, 
      q_4_5=>que_out_9_4_5, q_4_4=>que_out_9_4_4, q_4_3=>que_out_9_4_3, 
      q_4_2=>que_out_9_4_2, q_4_1=>que_out_9_4_1, q_4_0=>que_out_9_4_0, clk
      =>nx10720, load=>sel_que_9, reset=>nx10696);
   gen_queues_10_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_10_0_15, q_0_14=>que_out_10_0_14, q_0_13=>
      que_out_10_0_13, q_0_12=>que_out_10_0_12, q_0_11=>que_out_10_0_11, 
      q_0_10=>que_out_10_0_10, q_0_9=>que_out_10_0_9, q_0_8=>que_out_10_0_8, 
      q_0_7=>que_out_10_0_7, q_0_6=>que_out_10_0_6, q_0_5=>que_out_10_0_5, 
      q_0_4=>que_out_10_0_4, q_0_3=>que_out_10_0_3, q_0_2=>que_out_10_0_2, 
      q_0_1=>que_out_10_0_1, q_0_0=>que_out_10_0_0, q_1_15=>que_out_10_1_15, 
      q_1_14=>que_out_10_1_14, q_1_13=>que_out_10_1_13, q_1_12=>
      que_out_10_1_12, q_1_11=>que_out_10_1_11, q_1_10=>que_out_10_1_10, 
      q_1_9=>que_out_10_1_9, q_1_8=>que_out_10_1_8, q_1_7=>que_out_10_1_7, 
      q_1_6=>que_out_10_1_6, q_1_5=>que_out_10_1_5, q_1_4=>que_out_10_1_4, 
      q_1_3=>que_out_10_1_3, q_1_2=>que_out_10_1_2, q_1_1=>que_out_10_1_1, 
      q_1_0=>que_out_10_1_0, q_2_15=>que_out_10_2_15, q_2_14=>
      que_out_10_2_14, q_2_13=>que_out_10_2_13, q_2_12=>que_out_10_2_12, 
      q_2_11=>que_out_10_2_11, q_2_10=>que_out_10_2_10, q_2_9=>
      que_out_10_2_9, q_2_8=>que_out_10_2_8, q_2_7=>que_out_10_2_7, q_2_6=>
      que_out_10_2_6, q_2_5=>que_out_10_2_5, q_2_4=>que_out_10_2_4, q_2_3=>
      que_out_10_2_3, q_2_2=>que_out_10_2_2, q_2_1=>que_out_10_2_1, q_2_0=>
      que_out_10_2_0, q_3_15=>que_out_10_3_15, q_3_14=>que_out_10_3_14, 
      q_3_13=>que_out_10_3_13, q_3_12=>que_out_10_3_12, q_3_11=>
      que_out_10_3_11, q_3_10=>que_out_10_3_10, q_3_9=>que_out_10_3_9, q_3_8
      =>que_out_10_3_8, q_3_7=>que_out_10_3_7, q_3_6=>que_out_10_3_6, q_3_5
      =>que_out_10_3_5, q_3_4=>que_out_10_3_4, q_3_3=>que_out_10_3_3, q_3_2
      =>que_out_10_3_2, q_3_1=>que_out_10_3_1, q_3_0=>que_out_10_3_0, q_4_15
      =>que_out_10_4_15, q_4_14=>que_out_10_4_14, q_4_13=>que_out_10_4_13, 
      q_4_12=>que_out_10_4_12, q_4_11=>que_out_10_4_11, q_4_10=>
      que_out_10_4_10, q_4_9=>que_out_10_4_9, q_4_8=>que_out_10_4_8, q_4_7=>
      que_out_10_4_7, q_4_6=>que_out_10_4_6, q_4_5=>que_out_10_4_5, q_4_4=>
      que_out_10_4_4, q_4_3=>que_out_10_4_3, q_4_2=>que_out_10_4_2, q_4_1=>
      que_out_10_4_1, q_4_0=>que_out_10_4_0, clk=>nx10722, load=>sel_que_10, 
      reset=>nx10698);
   gen_queues_11_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_11_0_15, q_0_14=>que_out_11_0_14, q_0_13=>
      que_out_11_0_13, q_0_12=>que_out_11_0_12, q_0_11=>que_out_11_0_11, 
      q_0_10=>que_out_11_0_10, q_0_9=>que_out_11_0_9, q_0_8=>que_out_11_0_8, 
      q_0_7=>que_out_11_0_7, q_0_6=>que_out_11_0_6, q_0_5=>que_out_11_0_5, 
      q_0_4=>que_out_11_0_4, q_0_3=>que_out_11_0_3, q_0_2=>que_out_11_0_2, 
      q_0_1=>que_out_11_0_1, q_0_0=>que_out_11_0_0, q_1_15=>que_out_11_1_15, 
      q_1_14=>que_out_11_1_14, q_1_13=>que_out_11_1_13, q_1_12=>
      que_out_11_1_12, q_1_11=>que_out_11_1_11, q_1_10=>que_out_11_1_10, 
      q_1_9=>que_out_11_1_9, q_1_8=>que_out_11_1_8, q_1_7=>que_out_11_1_7, 
      q_1_6=>que_out_11_1_6, q_1_5=>que_out_11_1_5, q_1_4=>que_out_11_1_4, 
      q_1_3=>que_out_11_1_3, q_1_2=>que_out_11_1_2, q_1_1=>que_out_11_1_1, 
      q_1_0=>que_out_11_1_0, q_2_15=>que_out_11_2_15, q_2_14=>
      que_out_11_2_14, q_2_13=>que_out_11_2_13, q_2_12=>que_out_11_2_12, 
      q_2_11=>que_out_11_2_11, q_2_10=>que_out_11_2_10, q_2_9=>
      que_out_11_2_9, q_2_8=>que_out_11_2_8, q_2_7=>que_out_11_2_7, q_2_6=>
      que_out_11_2_6, q_2_5=>que_out_11_2_5, q_2_4=>que_out_11_2_4, q_2_3=>
      que_out_11_2_3, q_2_2=>que_out_11_2_2, q_2_1=>que_out_11_2_1, q_2_0=>
      que_out_11_2_0, q_3_15=>que_out_11_3_15, q_3_14=>que_out_11_3_14, 
      q_3_13=>que_out_11_3_13, q_3_12=>que_out_11_3_12, q_3_11=>
      que_out_11_3_11, q_3_10=>que_out_11_3_10, q_3_9=>que_out_11_3_9, q_3_8
      =>que_out_11_3_8, q_3_7=>que_out_11_3_7, q_3_6=>que_out_11_3_6, q_3_5
      =>que_out_11_3_5, q_3_4=>que_out_11_3_4, q_3_3=>que_out_11_3_3, q_3_2
      =>que_out_11_3_2, q_3_1=>que_out_11_3_1, q_3_0=>que_out_11_3_0, q_4_15
      =>que_out_11_4_15, q_4_14=>que_out_11_4_14, q_4_13=>que_out_11_4_13, 
      q_4_12=>que_out_11_4_12, q_4_11=>que_out_11_4_11, q_4_10=>
      que_out_11_4_10, q_4_9=>que_out_11_4_9, q_4_8=>que_out_11_4_8, q_4_7=>
      que_out_11_4_7, q_4_6=>que_out_11_4_6, q_4_5=>que_out_11_4_5, q_4_4=>
      que_out_11_4_4, q_4_3=>que_out_11_4_3, q_4_2=>que_out_11_4_2, q_4_1=>
      que_out_11_4_1, q_4_0=>que_out_11_4_0, clk=>nx10722, load=>sel_que_11, 
      reset=>nx10698);
   gen_queues_12_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_12_0_15, q_0_14=>que_out_12_0_14, q_0_13=>
      que_out_12_0_13, q_0_12=>que_out_12_0_12, q_0_11=>que_out_12_0_11, 
      q_0_10=>que_out_12_0_10, q_0_9=>que_out_12_0_9, q_0_8=>que_out_12_0_8, 
      q_0_7=>que_out_12_0_7, q_0_6=>que_out_12_0_6, q_0_5=>que_out_12_0_5, 
      q_0_4=>que_out_12_0_4, q_0_3=>que_out_12_0_3, q_0_2=>que_out_12_0_2, 
      q_0_1=>que_out_12_0_1, q_0_0=>que_out_12_0_0, q_1_15=>que_out_12_1_15, 
      q_1_14=>que_out_12_1_14, q_1_13=>que_out_12_1_13, q_1_12=>
      que_out_12_1_12, q_1_11=>que_out_12_1_11, q_1_10=>que_out_12_1_10, 
      q_1_9=>que_out_12_1_9, q_1_8=>que_out_12_1_8, q_1_7=>que_out_12_1_7, 
      q_1_6=>que_out_12_1_6, q_1_5=>que_out_12_1_5, q_1_4=>que_out_12_1_4, 
      q_1_3=>que_out_12_1_3, q_1_2=>que_out_12_1_2, q_1_1=>que_out_12_1_1, 
      q_1_0=>que_out_12_1_0, q_2_15=>que_out_12_2_15, q_2_14=>
      que_out_12_2_14, q_2_13=>que_out_12_2_13, q_2_12=>que_out_12_2_12, 
      q_2_11=>que_out_12_2_11, q_2_10=>que_out_12_2_10, q_2_9=>
      que_out_12_2_9, q_2_8=>que_out_12_2_8, q_2_7=>que_out_12_2_7, q_2_6=>
      que_out_12_2_6, q_2_5=>que_out_12_2_5, q_2_4=>que_out_12_2_4, q_2_3=>
      que_out_12_2_3, q_2_2=>que_out_12_2_2, q_2_1=>que_out_12_2_1, q_2_0=>
      que_out_12_2_0, q_3_15=>que_out_12_3_15, q_3_14=>que_out_12_3_14, 
      q_3_13=>que_out_12_3_13, q_3_12=>que_out_12_3_12, q_3_11=>
      que_out_12_3_11, q_3_10=>que_out_12_3_10, q_3_9=>que_out_12_3_9, q_3_8
      =>que_out_12_3_8, q_3_7=>que_out_12_3_7, q_3_6=>que_out_12_3_6, q_3_5
      =>que_out_12_3_5, q_3_4=>que_out_12_3_4, q_3_3=>que_out_12_3_3, q_3_2
      =>que_out_12_3_2, q_3_1=>que_out_12_3_1, q_3_0=>que_out_12_3_0, q_4_15
      =>que_out_12_4_15, q_4_14=>que_out_12_4_14, q_4_13=>que_out_12_4_13, 
      q_4_12=>que_out_12_4_12, q_4_11=>que_out_12_4_11, q_4_10=>
      que_out_12_4_10, q_4_9=>que_out_12_4_9, q_4_8=>que_out_12_4_8, q_4_7=>
      que_out_12_4_7, q_4_6=>que_out_12_4_6, q_4_5=>que_out_12_4_5, q_4_4=>
      que_out_12_4_4, q_4_3=>que_out_12_4_3, q_4_2=>que_out_12_4_2, q_4_1=>
      que_out_12_4_1, q_4_0=>que_out_12_4_0, clk=>nx10722, load=>sel_que_12, 
      reset=>nx10698);
   gen_queues_13_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_13_0_15, q_0_14=>que_out_13_0_14, q_0_13=>
      que_out_13_0_13, q_0_12=>que_out_13_0_12, q_0_11=>que_out_13_0_11, 
      q_0_10=>que_out_13_0_10, q_0_9=>que_out_13_0_9, q_0_8=>que_out_13_0_8, 
      q_0_7=>que_out_13_0_7, q_0_6=>que_out_13_0_6, q_0_5=>que_out_13_0_5, 
      q_0_4=>que_out_13_0_4, q_0_3=>que_out_13_0_3, q_0_2=>que_out_13_0_2, 
      q_0_1=>que_out_13_0_1, q_0_0=>que_out_13_0_0, q_1_15=>que_out_13_1_15, 
      q_1_14=>que_out_13_1_14, q_1_13=>que_out_13_1_13, q_1_12=>
      que_out_13_1_12, q_1_11=>que_out_13_1_11, q_1_10=>que_out_13_1_10, 
      q_1_9=>que_out_13_1_9, q_1_8=>que_out_13_1_8, q_1_7=>que_out_13_1_7, 
      q_1_6=>que_out_13_1_6, q_1_5=>que_out_13_1_5, q_1_4=>que_out_13_1_4, 
      q_1_3=>que_out_13_1_3, q_1_2=>que_out_13_1_2, q_1_1=>que_out_13_1_1, 
      q_1_0=>que_out_13_1_0, q_2_15=>que_out_13_2_15, q_2_14=>
      que_out_13_2_14, q_2_13=>que_out_13_2_13, q_2_12=>que_out_13_2_12, 
      q_2_11=>que_out_13_2_11, q_2_10=>que_out_13_2_10, q_2_9=>
      que_out_13_2_9, q_2_8=>que_out_13_2_8, q_2_7=>que_out_13_2_7, q_2_6=>
      que_out_13_2_6, q_2_5=>que_out_13_2_5, q_2_4=>que_out_13_2_4, q_2_3=>
      que_out_13_2_3, q_2_2=>que_out_13_2_2, q_2_1=>que_out_13_2_1, q_2_0=>
      que_out_13_2_0, q_3_15=>que_out_13_3_15, q_3_14=>que_out_13_3_14, 
      q_3_13=>que_out_13_3_13, q_3_12=>que_out_13_3_12, q_3_11=>
      que_out_13_3_11, q_3_10=>que_out_13_3_10, q_3_9=>que_out_13_3_9, q_3_8
      =>que_out_13_3_8, q_3_7=>que_out_13_3_7, q_3_6=>que_out_13_3_6, q_3_5
      =>que_out_13_3_5, q_3_4=>que_out_13_3_4, q_3_3=>que_out_13_3_3, q_3_2
      =>que_out_13_3_2, q_3_1=>que_out_13_3_1, q_3_0=>que_out_13_3_0, q_4_15
      =>que_out_13_4_15, q_4_14=>que_out_13_4_14, q_4_13=>que_out_13_4_13, 
      q_4_12=>que_out_13_4_12, q_4_11=>que_out_13_4_11, q_4_10=>
      que_out_13_4_10, q_4_9=>que_out_13_4_9, q_4_8=>que_out_13_4_8, q_4_7=>
      que_out_13_4_7, q_4_6=>que_out_13_4_6, q_4_5=>que_out_13_4_5, q_4_4=>
      que_out_13_4_4, q_4_3=>que_out_13_4_3, q_4_2=>que_out_13_4_2, q_4_1=>
      que_out_13_4_1, q_4_0=>que_out_13_4_0, clk=>nx10724, load=>sel_que_13, 
      reset=>nx10700);
   gen_queues_14_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_14_0_15, q_0_14=>que_out_14_0_14, q_0_13=>
      que_out_14_0_13, q_0_12=>que_out_14_0_12, q_0_11=>que_out_14_0_11, 
      q_0_10=>que_out_14_0_10, q_0_9=>que_out_14_0_9, q_0_8=>que_out_14_0_8, 
      q_0_7=>que_out_14_0_7, q_0_6=>que_out_14_0_6, q_0_5=>que_out_14_0_5, 
      q_0_4=>que_out_14_0_4, q_0_3=>que_out_14_0_3, q_0_2=>que_out_14_0_2, 
      q_0_1=>que_out_14_0_1, q_0_0=>que_out_14_0_0, q_1_15=>que_out_14_1_15, 
      q_1_14=>que_out_14_1_14, q_1_13=>que_out_14_1_13, q_1_12=>
      que_out_14_1_12, q_1_11=>que_out_14_1_11, q_1_10=>que_out_14_1_10, 
      q_1_9=>que_out_14_1_9, q_1_8=>que_out_14_1_8, q_1_7=>que_out_14_1_7, 
      q_1_6=>que_out_14_1_6, q_1_5=>que_out_14_1_5, q_1_4=>que_out_14_1_4, 
      q_1_3=>que_out_14_1_3, q_1_2=>que_out_14_1_2, q_1_1=>que_out_14_1_1, 
      q_1_0=>que_out_14_1_0, q_2_15=>que_out_14_2_15, q_2_14=>
      que_out_14_2_14, q_2_13=>que_out_14_2_13, q_2_12=>que_out_14_2_12, 
      q_2_11=>que_out_14_2_11, q_2_10=>que_out_14_2_10, q_2_9=>
      que_out_14_2_9, q_2_8=>que_out_14_2_8, q_2_7=>que_out_14_2_7, q_2_6=>
      que_out_14_2_6, q_2_5=>que_out_14_2_5, q_2_4=>que_out_14_2_4, q_2_3=>
      que_out_14_2_3, q_2_2=>que_out_14_2_2, q_2_1=>que_out_14_2_1, q_2_0=>
      que_out_14_2_0, q_3_15=>que_out_14_3_15, q_3_14=>que_out_14_3_14, 
      q_3_13=>que_out_14_3_13, q_3_12=>que_out_14_3_12, q_3_11=>
      que_out_14_3_11, q_3_10=>que_out_14_3_10, q_3_9=>que_out_14_3_9, q_3_8
      =>que_out_14_3_8, q_3_7=>que_out_14_3_7, q_3_6=>que_out_14_3_6, q_3_5
      =>que_out_14_3_5, q_3_4=>que_out_14_3_4, q_3_3=>que_out_14_3_3, q_3_2
      =>que_out_14_3_2, q_3_1=>que_out_14_3_1, q_3_0=>que_out_14_3_0, q_4_15
      =>que_out_14_4_15, q_4_14=>que_out_14_4_14, q_4_13=>que_out_14_4_13, 
      q_4_12=>que_out_14_4_12, q_4_11=>que_out_14_4_11, q_4_10=>
      que_out_14_4_10, q_4_9=>que_out_14_4_9, q_4_8=>que_out_14_4_8, q_4_7=>
      que_out_14_4_7, q_4_6=>que_out_14_4_6, q_4_5=>que_out_14_4_5, q_4_4=>
      que_out_14_4_4, q_4_3=>que_out_14_4_3, q_4_2=>que_out_14_4_2, q_4_1=>
      que_out_14_4_1, q_4_0=>que_out_14_4_0, clk=>nx10726, load=>sel_que_14, 
      reset=>nx10702);
   gen_queues_15_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_15_0_15, q_0_14=>que_out_15_0_14, q_0_13=>
      que_out_15_0_13, q_0_12=>que_out_15_0_12, q_0_11=>que_out_15_0_11, 
      q_0_10=>que_out_15_0_10, q_0_9=>que_out_15_0_9, q_0_8=>que_out_15_0_8, 
      q_0_7=>que_out_15_0_7, q_0_6=>que_out_15_0_6, q_0_5=>que_out_15_0_5, 
      q_0_4=>que_out_15_0_4, q_0_3=>que_out_15_0_3, q_0_2=>que_out_15_0_2, 
      q_0_1=>que_out_15_0_1, q_0_0=>que_out_15_0_0, q_1_15=>que_out_15_1_15, 
      q_1_14=>que_out_15_1_14, q_1_13=>que_out_15_1_13, q_1_12=>
      que_out_15_1_12, q_1_11=>que_out_15_1_11, q_1_10=>que_out_15_1_10, 
      q_1_9=>que_out_15_1_9, q_1_8=>que_out_15_1_8, q_1_7=>que_out_15_1_7, 
      q_1_6=>que_out_15_1_6, q_1_5=>que_out_15_1_5, q_1_4=>que_out_15_1_4, 
      q_1_3=>que_out_15_1_3, q_1_2=>que_out_15_1_2, q_1_1=>que_out_15_1_1, 
      q_1_0=>que_out_15_1_0, q_2_15=>que_out_15_2_15, q_2_14=>
      que_out_15_2_14, q_2_13=>que_out_15_2_13, q_2_12=>que_out_15_2_12, 
      q_2_11=>que_out_15_2_11, q_2_10=>que_out_15_2_10, q_2_9=>
      que_out_15_2_9, q_2_8=>que_out_15_2_8, q_2_7=>que_out_15_2_7, q_2_6=>
      que_out_15_2_6, q_2_5=>que_out_15_2_5, q_2_4=>que_out_15_2_4, q_2_3=>
      que_out_15_2_3, q_2_2=>que_out_15_2_2, q_2_1=>que_out_15_2_1, q_2_0=>
      que_out_15_2_0, q_3_15=>que_out_15_3_15, q_3_14=>que_out_15_3_14, 
      q_3_13=>que_out_15_3_13, q_3_12=>que_out_15_3_12, q_3_11=>
      que_out_15_3_11, q_3_10=>que_out_15_3_10, q_3_9=>que_out_15_3_9, q_3_8
      =>que_out_15_3_8, q_3_7=>que_out_15_3_7, q_3_6=>que_out_15_3_6, q_3_5
      =>que_out_15_3_5, q_3_4=>que_out_15_3_4, q_3_3=>que_out_15_3_3, q_3_2
      =>que_out_15_3_2, q_3_1=>que_out_15_3_1, q_3_0=>que_out_15_3_0, q_4_15
      =>que_out_15_4_15, q_4_14=>que_out_15_4_14, q_4_13=>que_out_15_4_13, 
      q_4_12=>que_out_15_4_12, q_4_11=>que_out_15_4_11, q_4_10=>
      que_out_15_4_10, q_4_9=>que_out_15_4_9, q_4_8=>que_out_15_4_8, q_4_7=>
      que_out_15_4_7, q_4_6=>que_out_15_4_6, q_4_5=>que_out_15_4_5, q_4_4=>
      que_out_15_4_4, q_4_3=>que_out_15_4_3, q_4_2=>que_out_15_4_2, q_4_1=>
      que_out_15_4_1, q_4_0=>que_out_15_4_0, clk=>nx10726, load=>sel_que_15, 
      reset=>nx10702);
   gen_queues_16_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_16_0_15, q_0_14=>que_out_16_0_14, q_0_13=>
      que_out_16_0_13, q_0_12=>que_out_16_0_12, q_0_11=>que_out_16_0_11, 
      q_0_10=>que_out_16_0_10, q_0_9=>que_out_16_0_9, q_0_8=>que_out_16_0_8, 
      q_0_7=>que_out_16_0_7, q_0_6=>que_out_16_0_6, q_0_5=>que_out_16_0_5, 
      q_0_4=>que_out_16_0_4, q_0_3=>que_out_16_0_3, q_0_2=>que_out_16_0_2, 
      q_0_1=>que_out_16_0_1, q_0_0=>que_out_16_0_0, q_1_15=>que_out_16_1_15, 
      q_1_14=>que_out_16_1_14, q_1_13=>que_out_16_1_13, q_1_12=>
      que_out_16_1_12, q_1_11=>que_out_16_1_11, q_1_10=>que_out_16_1_10, 
      q_1_9=>que_out_16_1_9, q_1_8=>que_out_16_1_8, q_1_7=>que_out_16_1_7, 
      q_1_6=>que_out_16_1_6, q_1_5=>que_out_16_1_5, q_1_4=>que_out_16_1_4, 
      q_1_3=>que_out_16_1_3, q_1_2=>que_out_16_1_2, q_1_1=>que_out_16_1_1, 
      q_1_0=>que_out_16_1_0, q_2_15=>que_out_16_2_15, q_2_14=>
      que_out_16_2_14, q_2_13=>que_out_16_2_13, q_2_12=>que_out_16_2_12, 
      q_2_11=>que_out_16_2_11, q_2_10=>que_out_16_2_10, q_2_9=>
      que_out_16_2_9, q_2_8=>que_out_16_2_8, q_2_7=>que_out_16_2_7, q_2_6=>
      que_out_16_2_6, q_2_5=>que_out_16_2_5, q_2_4=>que_out_16_2_4, q_2_3=>
      que_out_16_2_3, q_2_2=>que_out_16_2_2, q_2_1=>que_out_16_2_1, q_2_0=>
      que_out_16_2_0, q_3_15=>que_out_16_3_15, q_3_14=>que_out_16_3_14, 
      q_3_13=>que_out_16_3_13, q_3_12=>que_out_16_3_12, q_3_11=>
      que_out_16_3_11, q_3_10=>que_out_16_3_10, q_3_9=>que_out_16_3_9, q_3_8
      =>que_out_16_3_8, q_3_7=>que_out_16_3_7, q_3_6=>que_out_16_3_6, q_3_5
      =>que_out_16_3_5, q_3_4=>que_out_16_3_4, q_3_3=>que_out_16_3_3, q_3_2
      =>que_out_16_3_2, q_3_1=>que_out_16_3_1, q_3_0=>que_out_16_3_0, q_4_15
      =>que_out_16_4_15, q_4_14=>que_out_16_4_14, q_4_13=>que_out_16_4_13, 
      q_4_12=>que_out_16_4_12, q_4_11=>que_out_16_4_11, q_4_10=>
      que_out_16_4_10, q_4_9=>que_out_16_4_9, q_4_8=>que_out_16_4_8, q_4_7=>
      que_out_16_4_7, q_4_6=>que_out_16_4_6, q_4_5=>que_out_16_4_5, q_4_4=>
      que_out_16_4_4, q_4_3=>que_out_16_4_3, q_4_2=>que_out_16_4_2, q_4_1=>
      que_out_16_4_1, q_4_0=>que_out_16_4_0, clk=>nx10726, load=>sel_que_16, 
      reset=>nx10702);
   gen_queues_17_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_17_0_15, q_0_14=>que_out_17_0_14, q_0_13=>
      que_out_17_0_13, q_0_12=>que_out_17_0_12, q_0_11=>que_out_17_0_11, 
      q_0_10=>que_out_17_0_10, q_0_9=>que_out_17_0_9, q_0_8=>que_out_17_0_8, 
      q_0_7=>que_out_17_0_7, q_0_6=>que_out_17_0_6, q_0_5=>que_out_17_0_5, 
      q_0_4=>que_out_17_0_4, q_0_3=>que_out_17_0_3, q_0_2=>que_out_17_0_2, 
      q_0_1=>que_out_17_0_1, q_0_0=>que_out_17_0_0, q_1_15=>que_out_17_1_15, 
      q_1_14=>que_out_17_1_14, q_1_13=>que_out_17_1_13, q_1_12=>
      que_out_17_1_12, q_1_11=>que_out_17_1_11, q_1_10=>que_out_17_1_10, 
      q_1_9=>que_out_17_1_9, q_1_8=>que_out_17_1_8, q_1_7=>que_out_17_1_7, 
      q_1_6=>que_out_17_1_6, q_1_5=>que_out_17_1_5, q_1_4=>que_out_17_1_4, 
      q_1_3=>que_out_17_1_3, q_1_2=>que_out_17_1_2, q_1_1=>que_out_17_1_1, 
      q_1_0=>que_out_17_1_0, q_2_15=>que_out_17_2_15, q_2_14=>
      que_out_17_2_14, q_2_13=>que_out_17_2_13, q_2_12=>que_out_17_2_12, 
      q_2_11=>que_out_17_2_11, q_2_10=>que_out_17_2_10, q_2_9=>
      que_out_17_2_9, q_2_8=>que_out_17_2_8, q_2_7=>que_out_17_2_7, q_2_6=>
      que_out_17_2_6, q_2_5=>que_out_17_2_5, q_2_4=>que_out_17_2_4, q_2_3=>
      que_out_17_2_3, q_2_2=>que_out_17_2_2, q_2_1=>que_out_17_2_1, q_2_0=>
      que_out_17_2_0, q_3_15=>que_out_17_3_15, q_3_14=>que_out_17_3_14, 
      q_3_13=>que_out_17_3_13, q_3_12=>que_out_17_3_12, q_3_11=>
      que_out_17_3_11, q_3_10=>que_out_17_3_10, q_3_9=>que_out_17_3_9, q_3_8
      =>que_out_17_3_8, q_3_7=>que_out_17_3_7, q_3_6=>que_out_17_3_6, q_3_5
      =>que_out_17_3_5, q_3_4=>que_out_17_3_4, q_3_3=>que_out_17_3_3, q_3_2
      =>que_out_17_3_2, q_3_1=>que_out_17_3_1, q_3_0=>que_out_17_3_0, q_4_15
      =>que_out_17_4_15, q_4_14=>que_out_17_4_14, q_4_13=>que_out_17_4_13, 
      q_4_12=>que_out_17_4_12, q_4_11=>que_out_17_4_11, q_4_10=>
      que_out_17_4_10, q_4_9=>que_out_17_4_9, q_4_8=>que_out_17_4_8, q_4_7=>
      que_out_17_4_7, q_4_6=>que_out_17_4_6, q_4_5=>que_out_17_4_5, q_4_4=>
      que_out_17_4_4, q_4_3=>que_out_17_4_3, q_4_2=>que_out_17_4_2, q_4_1=>
      que_out_17_4_1, q_4_0=>que_out_17_4_0, clk=>nx10728, load=>sel_que_17, 
      reset=>nx10704);
   gen_queues_18_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_18_0_15, q_0_14=>que_out_18_0_14, q_0_13=>
      que_out_18_0_13, q_0_12=>que_out_18_0_12, q_0_11=>que_out_18_0_11, 
      q_0_10=>que_out_18_0_10, q_0_9=>que_out_18_0_9, q_0_8=>que_out_18_0_8, 
      q_0_7=>que_out_18_0_7, q_0_6=>que_out_18_0_6, q_0_5=>que_out_18_0_5, 
      q_0_4=>que_out_18_0_4, q_0_3=>que_out_18_0_3, q_0_2=>que_out_18_0_2, 
      q_0_1=>que_out_18_0_1, q_0_0=>que_out_18_0_0, q_1_15=>que_out_18_1_15, 
      q_1_14=>que_out_18_1_14, q_1_13=>que_out_18_1_13, q_1_12=>
      que_out_18_1_12, q_1_11=>que_out_18_1_11, q_1_10=>que_out_18_1_10, 
      q_1_9=>que_out_18_1_9, q_1_8=>que_out_18_1_8, q_1_7=>que_out_18_1_7, 
      q_1_6=>que_out_18_1_6, q_1_5=>que_out_18_1_5, q_1_4=>que_out_18_1_4, 
      q_1_3=>que_out_18_1_3, q_1_2=>que_out_18_1_2, q_1_1=>que_out_18_1_1, 
      q_1_0=>que_out_18_1_0, q_2_15=>que_out_18_2_15, q_2_14=>
      que_out_18_2_14, q_2_13=>que_out_18_2_13, q_2_12=>que_out_18_2_12, 
      q_2_11=>que_out_18_2_11, q_2_10=>que_out_18_2_10, q_2_9=>
      que_out_18_2_9, q_2_8=>que_out_18_2_8, q_2_7=>que_out_18_2_7, q_2_6=>
      que_out_18_2_6, q_2_5=>que_out_18_2_5, q_2_4=>que_out_18_2_4, q_2_3=>
      que_out_18_2_3, q_2_2=>que_out_18_2_2, q_2_1=>que_out_18_2_1, q_2_0=>
      que_out_18_2_0, q_3_15=>que_out_18_3_15, q_3_14=>que_out_18_3_14, 
      q_3_13=>que_out_18_3_13, q_3_12=>que_out_18_3_12, q_3_11=>
      que_out_18_3_11, q_3_10=>que_out_18_3_10, q_3_9=>que_out_18_3_9, q_3_8
      =>que_out_18_3_8, q_3_7=>que_out_18_3_7, q_3_6=>que_out_18_3_6, q_3_5
      =>que_out_18_3_5, q_3_4=>que_out_18_3_4, q_3_3=>que_out_18_3_3, q_3_2
      =>que_out_18_3_2, q_3_1=>que_out_18_3_1, q_3_0=>que_out_18_3_0, q_4_15
      =>que_out_18_4_15, q_4_14=>que_out_18_4_14, q_4_13=>que_out_18_4_13, 
      q_4_12=>que_out_18_4_12, q_4_11=>que_out_18_4_11, q_4_10=>
      que_out_18_4_10, q_4_9=>que_out_18_4_9, q_4_8=>que_out_18_4_8, q_4_7=>
      que_out_18_4_7, q_4_6=>que_out_18_4_6, q_4_5=>que_out_18_4_5, q_4_4=>
      que_out_18_4_4, q_4_3=>que_out_18_4_3, q_4_2=>que_out_18_4_2, q_4_1=>
      que_out_18_4_1, q_4_0=>que_out_18_4_0, clk=>nx10728, load=>sel_que_18, 
      reset=>nx10704);
   gen_queues_19_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_19_0_15, q_0_14=>que_out_19_0_14, q_0_13=>
      que_out_19_0_13, q_0_12=>que_out_19_0_12, q_0_11=>que_out_19_0_11, 
      q_0_10=>que_out_19_0_10, q_0_9=>que_out_19_0_9, q_0_8=>que_out_19_0_8, 
      q_0_7=>que_out_19_0_7, q_0_6=>que_out_19_0_6, q_0_5=>que_out_19_0_5, 
      q_0_4=>que_out_19_0_4, q_0_3=>que_out_19_0_3, q_0_2=>que_out_19_0_2, 
      q_0_1=>que_out_19_0_1, q_0_0=>que_out_19_0_0, q_1_15=>que_out_19_1_15, 
      q_1_14=>que_out_19_1_14, q_1_13=>que_out_19_1_13, q_1_12=>
      que_out_19_1_12, q_1_11=>que_out_19_1_11, q_1_10=>que_out_19_1_10, 
      q_1_9=>que_out_19_1_9, q_1_8=>que_out_19_1_8, q_1_7=>que_out_19_1_7, 
      q_1_6=>que_out_19_1_6, q_1_5=>que_out_19_1_5, q_1_4=>que_out_19_1_4, 
      q_1_3=>que_out_19_1_3, q_1_2=>que_out_19_1_2, q_1_1=>que_out_19_1_1, 
      q_1_0=>que_out_19_1_0, q_2_15=>que_out_19_2_15, q_2_14=>
      que_out_19_2_14, q_2_13=>que_out_19_2_13, q_2_12=>que_out_19_2_12, 
      q_2_11=>que_out_19_2_11, q_2_10=>que_out_19_2_10, q_2_9=>
      que_out_19_2_9, q_2_8=>que_out_19_2_8, q_2_7=>que_out_19_2_7, q_2_6=>
      que_out_19_2_6, q_2_5=>que_out_19_2_5, q_2_4=>que_out_19_2_4, q_2_3=>
      que_out_19_2_3, q_2_2=>que_out_19_2_2, q_2_1=>que_out_19_2_1, q_2_0=>
      que_out_19_2_0, q_3_15=>que_out_19_3_15, q_3_14=>que_out_19_3_14, 
      q_3_13=>que_out_19_3_13, q_3_12=>que_out_19_3_12, q_3_11=>
      que_out_19_3_11, q_3_10=>que_out_19_3_10, q_3_9=>que_out_19_3_9, q_3_8
      =>que_out_19_3_8, q_3_7=>que_out_19_3_7, q_3_6=>que_out_19_3_6, q_3_5
      =>que_out_19_3_5, q_3_4=>que_out_19_3_4, q_3_3=>que_out_19_3_3, q_3_2
      =>que_out_19_3_2, q_3_1=>que_out_19_3_1, q_3_0=>que_out_19_3_0, q_4_15
      =>que_out_19_4_15, q_4_14=>que_out_19_4_14, q_4_13=>que_out_19_4_13, 
      q_4_12=>que_out_19_4_12, q_4_11=>que_out_19_4_11, q_4_10=>
      que_out_19_4_10, q_4_9=>que_out_19_4_9, q_4_8=>que_out_19_4_8, q_4_7=>
      que_out_19_4_7, q_4_6=>que_out_19_4_6, q_4_5=>que_out_19_4_5, q_4_4=>
      que_out_19_4_4, q_4_3=>que_out_19_4_3, q_4_2=>que_out_19_4_2, q_4_1=>
      que_out_19_4_1, q_4_0=>que_out_19_4_0, clk=>nx10728, load=>sel_que_19, 
      reset=>nx10704);
   gen_queues_20_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_20_0_15, q_0_14=>que_out_20_0_14, q_0_13=>
      que_out_20_0_13, q_0_12=>que_out_20_0_12, q_0_11=>que_out_20_0_11, 
      q_0_10=>que_out_20_0_10, q_0_9=>que_out_20_0_9, q_0_8=>que_out_20_0_8, 
      q_0_7=>que_out_20_0_7, q_0_6=>que_out_20_0_6, q_0_5=>que_out_20_0_5, 
      q_0_4=>que_out_20_0_4, q_0_3=>que_out_20_0_3, q_0_2=>que_out_20_0_2, 
      q_0_1=>que_out_20_0_1, q_0_0=>que_out_20_0_0, q_1_15=>que_out_20_1_15, 
      q_1_14=>que_out_20_1_14, q_1_13=>que_out_20_1_13, q_1_12=>
      que_out_20_1_12, q_1_11=>que_out_20_1_11, q_1_10=>que_out_20_1_10, 
      q_1_9=>que_out_20_1_9, q_1_8=>que_out_20_1_8, q_1_7=>que_out_20_1_7, 
      q_1_6=>que_out_20_1_6, q_1_5=>que_out_20_1_5, q_1_4=>que_out_20_1_4, 
      q_1_3=>que_out_20_1_3, q_1_2=>que_out_20_1_2, q_1_1=>que_out_20_1_1, 
      q_1_0=>que_out_20_1_0, q_2_15=>que_out_20_2_15, q_2_14=>
      que_out_20_2_14, q_2_13=>que_out_20_2_13, q_2_12=>que_out_20_2_12, 
      q_2_11=>que_out_20_2_11, q_2_10=>que_out_20_2_10, q_2_9=>
      que_out_20_2_9, q_2_8=>que_out_20_2_8, q_2_7=>que_out_20_2_7, q_2_6=>
      que_out_20_2_6, q_2_5=>que_out_20_2_5, q_2_4=>que_out_20_2_4, q_2_3=>
      que_out_20_2_3, q_2_2=>que_out_20_2_2, q_2_1=>que_out_20_2_1, q_2_0=>
      que_out_20_2_0, q_3_15=>que_out_20_3_15, q_3_14=>que_out_20_3_14, 
      q_3_13=>que_out_20_3_13, q_3_12=>que_out_20_3_12, q_3_11=>
      que_out_20_3_11, q_3_10=>que_out_20_3_10, q_3_9=>que_out_20_3_9, q_3_8
      =>que_out_20_3_8, q_3_7=>que_out_20_3_7, q_3_6=>que_out_20_3_6, q_3_5
      =>que_out_20_3_5, q_3_4=>que_out_20_3_4, q_3_3=>que_out_20_3_3, q_3_2
      =>que_out_20_3_2, q_3_1=>que_out_20_3_1, q_3_0=>que_out_20_3_0, q_4_15
      =>que_out_20_4_15, q_4_14=>que_out_20_4_14, q_4_13=>que_out_20_4_13, 
      q_4_12=>que_out_20_4_12, q_4_11=>que_out_20_4_11, q_4_10=>
      que_out_20_4_10, q_4_9=>que_out_20_4_9, q_4_8=>que_out_20_4_8, q_4_7=>
      que_out_20_4_7, q_4_6=>que_out_20_4_6, q_4_5=>que_out_20_4_5, q_4_4=>
      que_out_20_4_4, q_4_3=>que_out_20_4_3, q_4_2=>que_out_20_4_2, q_4_1=>
      que_out_20_4_1, q_4_0=>que_out_20_4_0, clk=>nx10730, load=>sel_que_20, 
      reset=>nx10706);
   gen_queues_21_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_21_0_15, q_0_14=>que_out_21_0_14, q_0_13=>
      que_out_21_0_13, q_0_12=>que_out_21_0_12, q_0_11=>que_out_21_0_11, 
      q_0_10=>que_out_21_0_10, q_0_9=>que_out_21_0_9, q_0_8=>que_out_21_0_8, 
      q_0_7=>que_out_21_0_7, q_0_6=>que_out_21_0_6, q_0_5=>que_out_21_0_5, 
      q_0_4=>que_out_21_0_4, q_0_3=>que_out_21_0_3, q_0_2=>que_out_21_0_2, 
      q_0_1=>que_out_21_0_1, q_0_0=>que_out_21_0_0, q_1_15=>que_out_21_1_15, 
      q_1_14=>que_out_21_1_14, q_1_13=>que_out_21_1_13, q_1_12=>
      que_out_21_1_12, q_1_11=>que_out_21_1_11, q_1_10=>que_out_21_1_10, 
      q_1_9=>que_out_21_1_9, q_1_8=>que_out_21_1_8, q_1_7=>que_out_21_1_7, 
      q_1_6=>que_out_21_1_6, q_1_5=>que_out_21_1_5, q_1_4=>que_out_21_1_4, 
      q_1_3=>que_out_21_1_3, q_1_2=>que_out_21_1_2, q_1_1=>que_out_21_1_1, 
      q_1_0=>que_out_21_1_0, q_2_15=>que_out_21_2_15, q_2_14=>
      que_out_21_2_14, q_2_13=>que_out_21_2_13, q_2_12=>que_out_21_2_12, 
      q_2_11=>que_out_21_2_11, q_2_10=>que_out_21_2_10, q_2_9=>
      que_out_21_2_9, q_2_8=>que_out_21_2_8, q_2_7=>que_out_21_2_7, q_2_6=>
      que_out_21_2_6, q_2_5=>que_out_21_2_5, q_2_4=>que_out_21_2_4, q_2_3=>
      que_out_21_2_3, q_2_2=>que_out_21_2_2, q_2_1=>que_out_21_2_1, q_2_0=>
      que_out_21_2_0, q_3_15=>que_out_21_3_15, q_3_14=>que_out_21_3_14, 
      q_3_13=>que_out_21_3_13, q_3_12=>que_out_21_3_12, q_3_11=>
      que_out_21_3_11, q_3_10=>que_out_21_3_10, q_3_9=>que_out_21_3_9, q_3_8
      =>que_out_21_3_8, q_3_7=>que_out_21_3_7, q_3_6=>que_out_21_3_6, q_3_5
      =>que_out_21_3_5, q_3_4=>que_out_21_3_4, q_3_3=>que_out_21_3_3, q_3_2
      =>que_out_21_3_2, q_3_1=>que_out_21_3_1, q_3_0=>que_out_21_3_0, q_4_15
      =>que_out_21_4_15, q_4_14=>que_out_21_4_14, q_4_13=>que_out_21_4_13, 
      q_4_12=>que_out_21_4_12, q_4_11=>que_out_21_4_11, q_4_10=>
      que_out_21_4_10, q_4_9=>que_out_21_4_9, q_4_8=>que_out_21_4_8, q_4_7=>
      que_out_21_4_7, q_4_6=>que_out_21_4_6, q_4_5=>que_out_21_4_5, q_4_4=>
      que_out_21_4_4, q_4_3=>que_out_21_4_3, q_4_2=>que_out_21_4_2, q_4_1=>
      que_out_21_4_1, q_4_0=>que_out_21_4_0, clk=>nx10732, load=>sel_que_21, 
      reset=>nx10708);
   gen_queues_22_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_22_0_15, q_0_14=>que_out_22_0_14, q_0_13=>
      que_out_22_0_13, q_0_12=>que_out_22_0_12, q_0_11=>que_out_22_0_11, 
      q_0_10=>que_out_22_0_10, q_0_9=>que_out_22_0_9, q_0_8=>que_out_22_0_8, 
      q_0_7=>que_out_22_0_7, q_0_6=>que_out_22_0_6, q_0_5=>que_out_22_0_5, 
      q_0_4=>que_out_22_0_4, q_0_3=>que_out_22_0_3, q_0_2=>que_out_22_0_2, 
      q_0_1=>que_out_22_0_1, q_0_0=>que_out_22_0_0, q_1_15=>que_out_22_1_15, 
      q_1_14=>que_out_22_1_14, q_1_13=>que_out_22_1_13, q_1_12=>
      que_out_22_1_12, q_1_11=>que_out_22_1_11, q_1_10=>que_out_22_1_10, 
      q_1_9=>que_out_22_1_9, q_1_8=>que_out_22_1_8, q_1_7=>que_out_22_1_7, 
      q_1_6=>que_out_22_1_6, q_1_5=>que_out_22_1_5, q_1_4=>que_out_22_1_4, 
      q_1_3=>que_out_22_1_3, q_1_2=>que_out_22_1_2, q_1_1=>que_out_22_1_1, 
      q_1_0=>que_out_22_1_0, q_2_15=>que_out_22_2_15, q_2_14=>
      que_out_22_2_14, q_2_13=>que_out_22_2_13, q_2_12=>que_out_22_2_12, 
      q_2_11=>que_out_22_2_11, q_2_10=>que_out_22_2_10, q_2_9=>
      que_out_22_2_9, q_2_8=>que_out_22_2_8, q_2_7=>que_out_22_2_7, q_2_6=>
      que_out_22_2_6, q_2_5=>que_out_22_2_5, q_2_4=>que_out_22_2_4, q_2_3=>
      que_out_22_2_3, q_2_2=>que_out_22_2_2, q_2_1=>que_out_22_2_1, q_2_0=>
      que_out_22_2_0, q_3_15=>que_out_22_3_15, q_3_14=>que_out_22_3_14, 
      q_3_13=>que_out_22_3_13, q_3_12=>que_out_22_3_12, q_3_11=>
      que_out_22_3_11, q_3_10=>que_out_22_3_10, q_3_9=>que_out_22_3_9, q_3_8
      =>que_out_22_3_8, q_3_7=>que_out_22_3_7, q_3_6=>que_out_22_3_6, q_3_5
      =>que_out_22_3_5, q_3_4=>que_out_22_3_4, q_3_3=>que_out_22_3_3, q_3_2
      =>que_out_22_3_2, q_3_1=>que_out_22_3_1, q_3_0=>que_out_22_3_0, q_4_15
      =>que_out_22_4_15, q_4_14=>que_out_22_4_14, q_4_13=>que_out_22_4_13, 
      q_4_12=>que_out_22_4_12, q_4_11=>que_out_22_4_11, q_4_10=>
      que_out_22_4_10, q_4_9=>que_out_22_4_9, q_4_8=>que_out_22_4_8, q_4_7=>
      que_out_22_4_7, q_4_6=>que_out_22_4_6, q_4_5=>que_out_22_4_5, q_4_4=>
      que_out_22_4_4, q_4_3=>que_out_22_4_3, q_4_2=>que_out_22_4_2, q_4_1=>
      que_out_22_4_1, q_4_0=>que_out_22_4_0, clk=>nx10732, load=>sel_que_22, 
      reset=>nx10708);
   gen_queues_23_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_23_0_15, q_0_14=>que_out_23_0_14, q_0_13=>
      que_out_23_0_13, q_0_12=>que_out_23_0_12, q_0_11=>que_out_23_0_11, 
      q_0_10=>que_out_23_0_10, q_0_9=>que_out_23_0_9, q_0_8=>que_out_23_0_8, 
      q_0_7=>que_out_23_0_7, q_0_6=>que_out_23_0_6, q_0_5=>que_out_23_0_5, 
      q_0_4=>que_out_23_0_4, q_0_3=>que_out_23_0_3, q_0_2=>que_out_23_0_2, 
      q_0_1=>que_out_23_0_1, q_0_0=>que_out_23_0_0, q_1_15=>que_out_23_1_15, 
      q_1_14=>que_out_23_1_14, q_1_13=>que_out_23_1_13, q_1_12=>
      que_out_23_1_12, q_1_11=>que_out_23_1_11, q_1_10=>que_out_23_1_10, 
      q_1_9=>que_out_23_1_9, q_1_8=>que_out_23_1_8, q_1_7=>que_out_23_1_7, 
      q_1_6=>que_out_23_1_6, q_1_5=>que_out_23_1_5, q_1_4=>que_out_23_1_4, 
      q_1_3=>que_out_23_1_3, q_1_2=>que_out_23_1_2, q_1_1=>que_out_23_1_1, 
      q_1_0=>que_out_23_1_0, q_2_15=>que_out_23_2_15, q_2_14=>
      que_out_23_2_14, q_2_13=>que_out_23_2_13, q_2_12=>que_out_23_2_12, 
      q_2_11=>que_out_23_2_11, q_2_10=>que_out_23_2_10, q_2_9=>
      que_out_23_2_9, q_2_8=>que_out_23_2_8, q_2_7=>que_out_23_2_7, q_2_6=>
      que_out_23_2_6, q_2_5=>que_out_23_2_5, q_2_4=>que_out_23_2_4, q_2_3=>
      que_out_23_2_3, q_2_2=>que_out_23_2_2, q_2_1=>que_out_23_2_1, q_2_0=>
      que_out_23_2_0, q_3_15=>que_out_23_3_15, q_3_14=>que_out_23_3_14, 
      q_3_13=>que_out_23_3_13, q_3_12=>que_out_23_3_12, q_3_11=>
      que_out_23_3_11, q_3_10=>que_out_23_3_10, q_3_9=>que_out_23_3_9, q_3_8
      =>que_out_23_3_8, q_3_7=>que_out_23_3_7, q_3_6=>que_out_23_3_6, q_3_5
      =>que_out_23_3_5, q_3_4=>que_out_23_3_4, q_3_3=>que_out_23_3_3, q_3_2
      =>que_out_23_3_2, q_3_1=>que_out_23_3_1, q_3_0=>que_out_23_3_0, q_4_15
      =>que_out_23_4_15, q_4_14=>que_out_23_4_14, q_4_13=>que_out_23_4_13, 
      q_4_12=>que_out_23_4_12, q_4_11=>que_out_23_4_11, q_4_10=>
      que_out_23_4_10, q_4_9=>que_out_23_4_9, q_4_8=>que_out_23_4_8, q_4_7=>
      que_out_23_4_7, q_4_6=>que_out_23_4_6, q_4_5=>que_out_23_4_5, q_4_4=>
      que_out_23_4_4, q_4_3=>que_out_23_4_3, q_4_2=>que_out_23_4_2, q_4_1=>
      que_out_23_4_1, q_4_0=>que_out_23_4_0, clk=>nx10732, load=>sel_que_23, 
      reset=>nx10708);
   gen_queues_24_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_24_0_15, q_0_14=>que_out_24_0_14, q_0_13=>
      que_out_24_0_13, q_0_12=>que_out_24_0_12, q_0_11=>que_out_24_0_11, 
      q_0_10=>que_out_24_0_10, q_0_9=>que_out_24_0_9, q_0_8=>que_out_24_0_8, 
      q_0_7=>que_out_24_0_7, q_0_6=>que_out_24_0_6, q_0_5=>que_out_24_0_5, 
      q_0_4=>que_out_24_0_4, q_0_3=>que_out_24_0_3, q_0_2=>que_out_24_0_2, 
      q_0_1=>que_out_24_0_1, q_0_0=>que_out_24_0_0, q_1_15=>que_out_24_1_15, 
      q_1_14=>que_out_24_1_14, q_1_13=>que_out_24_1_13, q_1_12=>
      que_out_24_1_12, q_1_11=>que_out_24_1_11, q_1_10=>que_out_24_1_10, 
      q_1_9=>que_out_24_1_9, q_1_8=>que_out_24_1_8, q_1_7=>que_out_24_1_7, 
      q_1_6=>que_out_24_1_6, q_1_5=>que_out_24_1_5, q_1_4=>que_out_24_1_4, 
      q_1_3=>que_out_24_1_3, q_1_2=>que_out_24_1_2, q_1_1=>que_out_24_1_1, 
      q_1_0=>que_out_24_1_0, q_2_15=>que_out_24_2_15, q_2_14=>
      que_out_24_2_14, q_2_13=>que_out_24_2_13, q_2_12=>que_out_24_2_12, 
      q_2_11=>que_out_24_2_11, q_2_10=>que_out_24_2_10, q_2_9=>
      que_out_24_2_9, q_2_8=>que_out_24_2_8, q_2_7=>que_out_24_2_7, q_2_6=>
      que_out_24_2_6, q_2_5=>que_out_24_2_5, q_2_4=>que_out_24_2_4, q_2_3=>
      que_out_24_2_3, q_2_2=>que_out_24_2_2, q_2_1=>que_out_24_2_1, q_2_0=>
      que_out_24_2_0, q_3_15=>que_out_24_3_15, q_3_14=>que_out_24_3_14, 
      q_3_13=>que_out_24_3_13, q_3_12=>que_out_24_3_12, q_3_11=>
      que_out_24_3_11, q_3_10=>que_out_24_3_10, q_3_9=>que_out_24_3_9, q_3_8
      =>que_out_24_3_8, q_3_7=>que_out_24_3_7, q_3_6=>que_out_24_3_6, q_3_5
      =>que_out_24_3_5, q_3_4=>que_out_24_3_4, q_3_3=>que_out_24_3_3, q_3_2
      =>que_out_24_3_2, q_3_1=>que_out_24_3_1, q_3_0=>que_out_24_3_0, q_4_15
      =>que_out_24_4_15, q_4_14=>que_out_24_4_14, q_4_13=>que_out_24_4_13, 
      q_4_12=>que_out_24_4_12, q_4_11=>que_out_24_4_11, q_4_10=>
      que_out_24_4_10, q_4_9=>que_out_24_4_9, q_4_8=>que_out_24_4_8, q_4_7=>
      que_out_24_4_7, q_4_6=>que_out_24_4_6, q_4_5=>que_out_24_4_5, q_4_4=>
      que_out_24_4_4, q_4_3=>que_out_24_4_3, q_4_2=>que_out_24_4_2, q_4_1=>
      que_out_24_4_1, q_4_0=>que_out_24_4_0, clk=>nx10734, load=>sel_que_24, 
      reset=>nx10710);
   gen_queues_25_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_25_0_15, q_0_14=>que_out_25_0_14, q_0_13=>
      que_out_25_0_13, q_0_12=>que_out_25_0_12, q_0_11=>que_out_25_0_11, 
      q_0_10=>que_out_25_0_10, q_0_9=>que_out_25_0_9, q_0_8=>que_out_25_0_8, 
      q_0_7=>que_out_25_0_7, q_0_6=>que_out_25_0_6, q_0_5=>que_out_25_0_5, 
      q_0_4=>que_out_25_0_4, q_0_3=>que_out_25_0_3, q_0_2=>que_out_25_0_2, 
      q_0_1=>que_out_25_0_1, q_0_0=>que_out_25_0_0, q_1_15=>que_out_25_1_15, 
      q_1_14=>que_out_25_1_14, q_1_13=>que_out_25_1_13, q_1_12=>
      que_out_25_1_12, q_1_11=>que_out_25_1_11, q_1_10=>que_out_25_1_10, 
      q_1_9=>que_out_25_1_9, q_1_8=>que_out_25_1_8, q_1_7=>que_out_25_1_7, 
      q_1_6=>que_out_25_1_6, q_1_5=>que_out_25_1_5, q_1_4=>que_out_25_1_4, 
      q_1_3=>que_out_25_1_3, q_1_2=>que_out_25_1_2, q_1_1=>que_out_25_1_1, 
      q_1_0=>que_out_25_1_0, q_2_15=>que_out_25_2_15, q_2_14=>
      que_out_25_2_14, q_2_13=>que_out_25_2_13, q_2_12=>que_out_25_2_12, 
      q_2_11=>que_out_25_2_11, q_2_10=>que_out_25_2_10, q_2_9=>
      que_out_25_2_9, q_2_8=>que_out_25_2_8, q_2_7=>que_out_25_2_7, q_2_6=>
      que_out_25_2_6, q_2_5=>que_out_25_2_5, q_2_4=>que_out_25_2_4, q_2_3=>
      que_out_25_2_3, q_2_2=>que_out_25_2_2, q_2_1=>que_out_25_2_1, q_2_0=>
      que_out_25_2_0, q_3_15=>que_out_25_3_15, q_3_14=>que_out_25_3_14, 
      q_3_13=>que_out_25_3_13, q_3_12=>que_out_25_3_12, q_3_11=>
      que_out_25_3_11, q_3_10=>que_out_25_3_10, q_3_9=>que_out_25_3_9, q_3_8
      =>que_out_25_3_8, q_3_7=>que_out_25_3_7, q_3_6=>que_out_25_3_6, q_3_5
      =>que_out_25_3_5, q_3_4=>que_out_25_3_4, q_3_3=>que_out_25_3_3, q_3_2
      =>que_out_25_3_2, q_3_1=>que_out_25_3_1, q_3_0=>que_out_25_3_0, q_4_15
      =>que_out_25_4_15, q_4_14=>que_out_25_4_14, q_4_13=>que_out_25_4_13, 
      q_4_12=>que_out_25_4_12, q_4_11=>que_out_25_4_11, q_4_10=>
      que_out_25_4_10, q_4_9=>que_out_25_4_9, q_4_8=>que_out_25_4_8, q_4_7=>
      que_out_25_4_7, q_4_6=>que_out_25_4_6, q_4_5=>que_out_25_4_5, q_4_4=>
      que_out_25_4_4, q_4_3=>que_out_25_4_3, q_4_2=>que_out_25_4_2, q_4_1=>
      que_out_25_4_1, q_4_0=>que_out_25_4_0, clk=>nx10734, load=>sel_que_25, 
      reset=>nx10710);
   gen_queues_26_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_26_0_15, q_0_14=>que_out_26_0_14, q_0_13=>
      que_out_26_0_13, q_0_12=>que_out_26_0_12, q_0_11=>que_out_26_0_11, 
      q_0_10=>que_out_26_0_10, q_0_9=>que_out_26_0_9, q_0_8=>que_out_26_0_8, 
      q_0_7=>que_out_26_0_7, q_0_6=>que_out_26_0_6, q_0_5=>que_out_26_0_5, 
      q_0_4=>que_out_26_0_4, q_0_3=>que_out_26_0_3, q_0_2=>que_out_26_0_2, 
      q_0_1=>que_out_26_0_1, q_0_0=>que_out_26_0_0, q_1_15=>que_out_26_1_15, 
      q_1_14=>que_out_26_1_14, q_1_13=>que_out_26_1_13, q_1_12=>
      que_out_26_1_12, q_1_11=>que_out_26_1_11, q_1_10=>que_out_26_1_10, 
      q_1_9=>que_out_26_1_9, q_1_8=>que_out_26_1_8, q_1_7=>que_out_26_1_7, 
      q_1_6=>que_out_26_1_6, q_1_5=>que_out_26_1_5, q_1_4=>que_out_26_1_4, 
      q_1_3=>que_out_26_1_3, q_1_2=>que_out_26_1_2, q_1_1=>que_out_26_1_1, 
      q_1_0=>que_out_26_1_0, q_2_15=>que_out_26_2_15, q_2_14=>
      que_out_26_2_14, q_2_13=>que_out_26_2_13, q_2_12=>que_out_26_2_12, 
      q_2_11=>que_out_26_2_11, q_2_10=>que_out_26_2_10, q_2_9=>
      que_out_26_2_9, q_2_8=>que_out_26_2_8, q_2_7=>que_out_26_2_7, q_2_6=>
      que_out_26_2_6, q_2_5=>que_out_26_2_5, q_2_4=>que_out_26_2_4, q_2_3=>
      que_out_26_2_3, q_2_2=>que_out_26_2_2, q_2_1=>que_out_26_2_1, q_2_0=>
      que_out_26_2_0, q_3_15=>que_out_26_3_15, q_3_14=>que_out_26_3_14, 
      q_3_13=>que_out_26_3_13, q_3_12=>que_out_26_3_12, q_3_11=>
      que_out_26_3_11, q_3_10=>que_out_26_3_10, q_3_9=>que_out_26_3_9, q_3_8
      =>que_out_26_3_8, q_3_7=>que_out_26_3_7, q_3_6=>que_out_26_3_6, q_3_5
      =>que_out_26_3_5, q_3_4=>que_out_26_3_4, q_3_3=>que_out_26_3_3, q_3_2
      =>que_out_26_3_2, q_3_1=>que_out_26_3_1, q_3_0=>que_out_26_3_0, q_4_15
      =>que_out_26_4_15, q_4_14=>que_out_26_4_14, q_4_13=>que_out_26_4_13, 
      q_4_12=>que_out_26_4_12, q_4_11=>que_out_26_4_11, q_4_10=>
      que_out_26_4_10, q_4_9=>que_out_26_4_9, q_4_8=>que_out_26_4_8, q_4_7=>
      que_out_26_4_7, q_4_6=>que_out_26_4_6, q_4_5=>que_out_26_4_5, q_4_4=>
      que_out_26_4_4, q_4_3=>que_out_26_4_3, q_4_2=>que_out_26_4_2, q_4_1=>
      que_out_26_4_1, q_4_0=>que_out_26_4_0, clk=>nx10734, load=>sel_que_26, 
      reset=>nx10710);
   gen_queues_27_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_27_0_15, q_0_14=>que_out_27_0_14, q_0_13=>
      que_out_27_0_13, q_0_12=>que_out_27_0_12, q_0_11=>que_out_27_0_11, 
      q_0_10=>que_out_27_0_10, q_0_9=>que_out_27_0_9, q_0_8=>que_out_27_0_8, 
      q_0_7=>que_out_27_0_7, q_0_6=>que_out_27_0_6, q_0_5=>que_out_27_0_5, 
      q_0_4=>que_out_27_0_4, q_0_3=>que_out_27_0_3, q_0_2=>que_out_27_0_2, 
      q_0_1=>que_out_27_0_1, q_0_0=>que_out_27_0_0, q_1_15=>que_out_27_1_15, 
      q_1_14=>que_out_27_1_14, q_1_13=>que_out_27_1_13, q_1_12=>
      que_out_27_1_12, q_1_11=>que_out_27_1_11, q_1_10=>que_out_27_1_10, 
      q_1_9=>que_out_27_1_9, q_1_8=>que_out_27_1_8, q_1_7=>que_out_27_1_7, 
      q_1_6=>que_out_27_1_6, q_1_5=>que_out_27_1_5, q_1_4=>que_out_27_1_4, 
      q_1_3=>que_out_27_1_3, q_1_2=>que_out_27_1_2, q_1_1=>que_out_27_1_1, 
      q_1_0=>que_out_27_1_0, q_2_15=>que_out_27_2_15, q_2_14=>
      que_out_27_2_14, q_2_13=>que_out_27_2_13, q_2_12=>que_out_27_2_12, 
      q_2_11=>que_out_27_2_11, q_2_10=>que_out_27_2_10, q_2_9=>
      que_out_27_2_9, q_2_8=>que_out_27_2_8, q_2_7=>que_out_27_2_7, q_2_6=>
      que_out_27_2_6, q_2_5=>que_out_27_2_5, q_2_4=>que_out_27_2_4, q_2_3=>
      que_out_27_2_3, q_2_2=>que_out_27_2_2, q_2_1=>que_out_27_2_1, q_2_0=>
      que_out_27_2_0, q_3_15=>que_out_27_3_15, q_3_14=>que_out_27_3_14, 
      q_3_13=>que_out_27_3_13, q_3_12=>que_out_27_3_12, q_3_11=>
      que_out_27_3_11, q_3_10=>que_out_27_3_10, q_3_9=>que_out_27_3_9, q_3_8
      =>que_out_27_3_8, q_3_7=>que_out_27_3_7, q_3_6=>que_out_27_3_6, q_3_5
      =>que_out_27_3_5, q_3_4=>que_out_27_3_4, q_3_3=>que_out_27_3_3, q_3_2
      =>que_out_27_3_2, q_3_1=>que_out_27_3_1, q_3_0=>que_out_27_3_0, q_4_15
      =>que_out_27_4_15, q_4_14=>que_out_27_4_14, q_4_13=>que_out_27_4_13, 
      q_4_12=>que_out_27_4_12, q_4_11=>que_out_27_4_11, q_4_10=>
      que_out_27_4_10, q_4_9=>que_out_27_4_9, q_4_8=>que_out_27_4_8, q_4_7=>
      que_out_27_4_7, q_4_6=>que_out_27_4_6, q_4_5=>que_out_27_4_5, q_4_4=>
      que_out_27_4_4, q_4_3=>que_out_27_4_3, q_4_2=>que_out_27_4_2, q_4_1=>
      que_out_27_4_1, q_4_0=>que_out_27_4_0, clk=>nx10736, load=>sel_que_27, 
      reset=>nx10712);
   ix6830 : nand03 port map ( Y=>nx6829, A0=>nx8938, A1=>nx6833, A2=>nx6835
   );
   ix8939 : nor02ii port map ( Y=>nx8938, A0=>cache_in_sel(4), A1=>
      decoder_enable);
   ix6834 : inv01 port map ( Y=>nx6833, A=>cache_in_sel(1));
   ix6836 : inv01 port map ( Y=>nx6835, A=>cache_in_sel(0));
   ix6840 : nand03 port map ( Y=>nx6839, A0=>nx8938, A1=>nx6833, A2=>nx10508
   );
   ix6844 : nand03 port map ( Y=>nx6843, A0=>nx8938, A1=>nx10506, A2=>nx6835
   );
   ix6848 : nand03 port map ( Y=>nx6847, A0=>nx8938, A1=>nx10506, A2=>
      nx10508);
   ix9023 : nor02_2x port map ( Y=>sel_que_12, A0=>nx6875, A1=>nx6829);
   ix6876 : nand02 port map ( Y=>nx6875, A0=>cache_in_sel(3), A1=>
      cache_in_sel(2));
   ix9025 : nor02_2x port map ( Y=>sel_que_13, A0=>nx6875, A1=>nx6839);
   ix9027 : nor02_2x port map ( Y=>sel_que_14, A0=>nx6843, A1=>nx6875);
   ix9029 : nor02_2x port map ( Y=>sel_que_15, A0=>nx6875, A1=>nx6847);
   ix9043 : and02 port map ( Y=>sel_que_16, A0=>nx6885, A1=>nx9038);
   ix6886 : nor02_2x port map ( Y=>nx6885, A0=>cache_in_sel(2), A1=>
      cache_in_sel(3));
   ix9039 : nor03_2x port map ( Y=>nx9038, A0=>nx6889, A1=>nx10506, A2=>
      nx10508);
   ix6890 : nand02 port map ( Y=>nx6889, A0=>cache_in_sel(4), A1=>
      decoder_enable);
   ix6894 : nand04 port map ( Y=>nx6893, A0=>cache_in_sel(4), A1=>
      decoder_enable, A2=>nx6833, A3=>nx10508);
   ix6898 : nand04 port map ( Y=>nx6897, A0=>cache_in_sel(4), A1=>
      decoder_enable, A2=>nx10506, A3=>nx6835);
   ix6902 : nand04 port map ( Y=>nx6901, A0=>cache_in_sel(4), A1=>
      decoder_enable, A2=>nx10506, A3=>nx10508);
   ix9075 : and02 port map ( Y=>sel_que_20, A0=>nx6905, A1=>nx9038);
   ix9091 : and02 port map ( Y=>sel_que_24, A0=>nx6915, A1=>nx9038);
   ix243 : or04 port map ( Y=>out_column_4_0, A0=>nx238, A1=>nx188, A2=>
      nx130, A3=>nx82);
   ix239 : nand03 port map ( Y=>nx238, A0=>nx6927, A1=>nx6951, A2=>nx6967);
   ix6928 : aoi222 port map ( Y=>nx6927, A0=>que_out_10_4_0, A1=>nx10298, B0
      =>que_out_6_4_0, B1=>nx10350, C0=>que_out_9_4_0, C1=>nx10324);
   ix6932 : nand02_2x port map ( Y=>nx6931, A0=>cache_out_sel(3), A1=>nx6933
   );
   ix6934 : inv01 port map ( Y=>nx6933, A=>cache_out_sel(0));
   ix6938 : inv01 port map ( Y=>nx6937, A=>cache_out_sel(4));
   ix6940 : inv02 port map ( Y=>nx6939, A=>cache_out_sel(2));
   ix6946 : nand03 port map ( Y=>nx6945, A0=>nx10502, A1=>nx6937, A2=>
      nx10498);
   ix227 : nor04 port map ( Y=>nx226, A0=>nx6949, A1=>nx10502, A2=>nx10494, 
      A3=>nx10498);
   ix6950 : nand02_2x port map ( Y=>nx6949, A0=>cache_out_sel(3), A1=>
      cache_out_sel(0));
   ix6952 : aoi22 port map ( Y=>nx6951, A0=>que_out_5_4_0, A1=>nx10246, B0=>
      que_out_18_4_0, B1=>nx10272);
   ix6956 : nand02 port map ( Y=>nx6955, A0=>nx6957, A1=>cache_out_sel(0));
   ix6958 : inv01 port map ( Y=>nx6957, A=>cache_out_sel(3));
   ix6962 : inv01 port map ( Y=>nx6961, A=>cache_out_sel(1));
   ix215 : nor03_2x port map ( Y=>nx214, A0=>nx6965, A1=>nx10498, A2=>nx6943
   );
   ix6966 : nand02_2x port map ( Y=>nx6965, A0=>nx10494, A1=>nx10504);
   ix6968 : aoi22 port map ( Y=>nx6967, A0=>que_out_17_4_0, A1=>nx10220, B0
      =>que_out_20_4_0, B1=>nx10194);
   ix201 : nor03_2x port map ( Y=>nx200, A0=>nx6971, A1=>nx10498, A2=>
      nx10374);
   ix6972 : nand02_2x port map ( Y=>nx6971, A0=>nx10496, A1=>nx6961);
   ix193 : nor03_2x port map ( Y=>nx192, A0=>nx6971, A1=>nx6939, A2=>nx6943
   );
   ix189 : nand03 port map ( Y=>nx188, A0=>nx6977, A1=>nx6985, A2=>nx6991);
   ix6978 : aoi222 port map ( Y=>nx6977, A0=>que_out_19_4_0, A1=>nx10168, B0
      =>que_out_21_4_0, B1=>nx10142, C0=>que_out_8_4_0, C1=>nx10116);
   ix181 : nor03_2x port map ( Y=>nx180, A0=>nx6965, A1=>nx10498, A2=>
      nx10374);
   ix173 : nor03_2x port map ( Y=>nx172, A0=>nx6971, A1=>nx6939, A2=>nx10374
   );
   ix167 : nor04 port map ( Y=>nx166, A0=>nx6931, A1=>nx10502, A2=>nx10494, 
      A3=>nx10498);
   ix6986 : aoi22 port map ( Y=>nx6985, A0=>que_out_25_4_0, A1=>nx10064, B0
      =>que_out_16_4_0, B1=>nx10090);
   ix151 : nor02_2x port map ( Y=>nx150, A0=>nx6949, A1=>nx6971);
   ix159 : nor03_2x port map ( Y=>nx158, A0=>nx6971, A1=>nx10498, A2=>nx6943
   );
   ix6992 : aoi22 port map ( Y=>nx6991, A0=>que_out_24_4_0, A1=>nx10038, B0
      =>que_out_22_4_0, B1=>nx10012);
   ix145 : nor02_2x port map ( Y=>nx144, A0=>nx6971, A1=>nx6931);
   ix137 : nor03_2x port map ( Y=>nx136, A0=>nx6965, A1=>nx6939, A2=>nx6943
   );
   ix131 : nand03 port map ( Y=>nx130, A0=>nx6999, A1=>nx7007, A2=>nx7017);
   ix7000 : aoi222 port map ( Y=>nx6999, A0=>que_out_15_4_0, A1=>nx9960, B0
      =>que_out_3_4_0, B1=>nx9986, C0=>que_out_23_4_0, C1=>nx9934);
   ix119 : nor02_2x port map ( Y=>nx118, A0=>nx6949, A1=>nx6945);
   ix115 : nor03_2x port map ( Y=>nx114, A0=>nx6965, A1=>nx6939, A2=>nx10374
   );
   ix7008 : aoi22 port map ( Y=>nx7007, A0=>que_out_27_4_0, A1=>nx9908, B0=>
      que_out_4_4_0, B1=>nx9882);
   ix105 : nor02_2x port map ( Y=>nx104, A0=>nx6949, A1=>nx6965);
   ix101 : and02 port map ( Y=>nx100, A0=>nx88, A1=>nx28);
   ix89 : nor02_2x port map ( Y=>nx88, A0=>cache_out_sel(3), A1=>
      cache_out_sel(0));
   ix29 : nor03_2x port map ( Y=>nx28, A0=>nx10502, A1=>nx10494, A2=>nx6939
   );
   ix7018 : aoi22 port map ( Y=>nx7017, A0=>que_out_0_4_0, A1=>nx9830, B0=>
      que_out_2_4_0, B1=>nx9856);
   ix91 : and02 port map ( Y=>nx90, A0=>nx88, A1=>nx12);
   ix13 : nor03_2x port map ( Y=>nx12, A0=>nx10504, A1=>nx10494, A2=>nx10500
   );
   ix95 : and02 port map ( Y=>nx94, A0=>nx88, A1=>nx62);
   ix63 : nor03_2x port map ( Y=>nx62, A0=>nx6961, A1=>nx10494, A2=>nx10500
   );
   ix83 : nand03 port map ( Y=>nx82, A0=>nx7029, A1=>nx7037, A2=>nx7043);
   ix7030 : aoi222 port map ( Y=>nx7029, A0=>que_out_26_4_0, A1=>nx9804, B0
      =>que_out_14_4_0, B1=>nx9778, C0=>que_out_11_4_0, C1=>nx9752);
   ix75 : nor02_2x port map ( Y=>nx74, A0=>nx6965, A1=>nx6931);
   ix69 : nor02_2x port map ( Y=>nx68, A0=>nx6931, A1=>nx6945);
   ix7038 : aoi22 port map ( Y=>nx7037, A0=>que_out_13_4_0, A1=>nx9726, B0=>
      que_out_7_4_0, B1=>nx9700);
   ix43 : nor02_2x port map ( Y=>nx42, A0=>nx10374, A1=>nx6945);
   ix7044 : aoi22 port map ( Y=>nx7043, A0=>que_out_12_4_0, A1=>nx9674, B0=>
      que_out_1_4_0, B1=>nx9648);
   ix15 : nor04 port map ( Y=>nx14, A0=>nx10376, A1=>nx10504, A2=>nx10494, 
      A3=>nx10500);
   ix353 : or04 port map ( Y=>out_column_4_1, A0=>nx348, A1=>nx322, A2=>
      nx294, A3=>nx268);
   ix349 : nand03 port map ( Y=>nx348, A0=>nx7053, A1=>nx7055, A2=>nx7057);
   ix7054 : aoi222 port map ( Y=>nx7053, A0=>que_out_10_4_1, A1=>nx10298, B0
      =>que_out_6_4_1, B1=>nx10350, C0=>que_out_9_4_1, C1=>nx10324);
   ix7056 : aoi22 port map ( Y=>nx7055, A0=>que_out_5_4_1, A1=>nx10246, B0=>
      que_out_18_4_1, B1=>nx10272);
   ix7058 : aoi22 port map ( Y=>nx7057, A0=>que_out_17_4_1, A1=>nx10220, B0
      =>que_out_20_4_1, B1=>nx10194);
   ix323 : nand03 port map ( Y=>nx322, A0=>nx7061, A1=>nx7063, A2=>nx7065);
   ix7062 : aoi222 port map ( Y=>nx7061, A0=>que_out_19_4_1, A1=>nx10168, B0
      =>que_out_21_4_1, B1=>nx10142, C0=>que_out_8_4_1, C1=>nx10116);
   ix7064 : aoi22 port map ( Y=>nx7063, A0=>que_out_25_4_1, A1=>nx10064, B0
      =>que_out_16_4_1, B1=>nx10090);
   ix7066 : aoi22 port map ( Y=>nx7065, A0=>que_out_24_4_1, A1=>nx10038, B0
      =>que_out_22_4_1, B1=>nx10012);
   ix295 : nand03 port map ( Y=>nx294, A0=>nx7069, A1=>nx7071, A2=>nx7073);
   ix7070 : aoi222 port map ( Y=>nx7069, A0=>que_out_15_4_1, A1=>nx9960, B0
      =>que_out_3_4_1, B1=>nx9986, C0=>que_out_23_4_1, C1=>nx9934);
   ix7072 : aoi22 port map ( Y=>nx7071, A0=>que_out_27_4_1, A1=>nx9908, B0=>
      que_out_4_4_1, B1=>nx9882);
   ix7074 : aoi22 port map ( Y=>nx7073, A0=>que_out_0_4_1, A1=>nx9830, B0=>
      que_out_2_4_1, B1=>nx9856);
   ix269 : nand03 port map ( Y=>nx268, A0=>nx7077, A1=>nx7079, A2=>nx7081);
   ix7078 : aoi222 port map ( Y=>nx7077, A0=>que_out_26_4_1, A1=>nx9804, B0
      =>que_out_14_4_1, B1=>nx9778, C0=>que_out_11_4_1, C1=>nx9752);
   ix7080 : aoi22 port map ( Y=>nx7079, A0=>que_out_13_4_1, A1=>nx9726, B0=>
      que_out_7_4_1, B1=>nx9700);
   ix7082 : aoi22 port map ( Y=>nx7081, A0=>que_out_12_4_1, A1=>nx9674, B0=>
      que_out_1_4_1, B1=>nx9648);
   ix463 : or04 port map ( Y=>out_column_4_2, A0=>nx458, A1=>nx432, A2=>
      nx404, A3=>nx378);
   ix459 : nand03 port map ( Y=>nx458, A0=>nx7087, A1=>nx7089, A2=>nx7091);
   ix7088 : aoi222 port map ( Y=>nx7087, A0=>que_out_10_4_2, A1=>nx10298, B0
      =>que_out_6_4_2, B1=>nx10350, C0=>que_out_9_4_2, C1=>nx10324);
   ix7090 : aoi22 port map ( Y=>nx7089, A0=>que_out_5_4_2, A1=>nx10246, B0=>
      que_out_18_4_2, B1=>nx10272);
   ix7092 : aoi22 port map ( Y=>nx7091, A0=>que_out_17_4_2, A1=>nx10220, B0
      =>que_out_20_4_2, B1=>nx10194);
   ix433 : nand03 port map ( Y=>nx432, A0=>nx7095, A1=>nx7097, A2=>nx7099);
   ix7096 : aoi222 port map ( Y=>nx7095, A0=>que_out_19_4_2, A1=>nx10168, B0
      =>que_out_21_4_2, B1=>nx10142, C0=>que_out_8_4_2, C1=>nx10116);
   ix7098 : aoi22 port map ( Y=>nx7097, A0=>que_out_25_4_2, A1=>nx10064, B0
      =>que_out_16_4_2, B1=>nx10090);
   ix7100 : aoi22 port map ( Y=>nx7099, A0=>que_out_24_4_2, A1=>nx10038, B0
      =>que_out_22_4_2, B1=>nx10012);
   ix405 : nand03 port map ( Y=>nx404, A0=>nx7103, A1=>nx7105, A2=>nx7107);
   ix7104 : aoi222 port map ( Y=>nx7103, A0=>que_out_15_4_2, A1=>nx9960, B0
      =>que_out_3_4_2, B1=>nx9986, C0=>que_out_23_4_2, C1=>nx9934);
   ix7106 : aoi22 port map ( Y=>nx7105, A0=>que_out_27_4_2, A1=>nx9908, B0=>
      que_out_4_4_2, B1=>nx9882);
   ix7108 : aoi22 port map ( Y=>nx7107, A0=>que_out_0_4_2, A1=>nx9830, B0=>
      que_out_2_4_2, B1=>nx9856);
   ix379 : nand03 port map ( Y=>nx378, A0=>nx7111, A1=>nx7113, A2=>nx7115);
   ix7112 : aoi222 port map ( Y=>nx7111, A0=>que_out_26_4_2, A1=>nx9804, B0
      =>que_out_14_4_2, B1=>nx9778, C0=>que_out_11_4_2, C1=>nx9752);
   ix7114 : aoi22 port map ( Y=>nx7113, A0=>que_out_13_4_2, A1=>nx9726, B0=>
      que_out_7_4_2, B1=>nx9700);
   ix7116 : aoi22 port map ( Y=>nx7115, A0=>que_out_12_4_2, A1=>nx9674, B0=>
      que_out_1_4_2, B1=>nx9648);
   ix573 : or04 port map ( Y=>out_column_4_3, A0=>nx568, A1=>nx542, A2=>
      nx514, A3=>nx488);
   ix569 : nand03 port map ( Y=>nx568, A0=>nx7121, A1=>nx7123, A2=>nx7125);
   ix7122 : aoi222 port map ( Y=>nx7121, A0=>que_out_10_4_3, A1=>nx10298, B0
      =>que_out_6_4_3, B1=>nx10350, C0=>que_out_9_4_3, C1=>nx10324);
   ix7124 : aoi22 port map ( Y=>nx7123, A0=>que_out_5_4_3, A1=>nx10246, B0=>
      que_out_18_4_3, B1=>nx10272);
   ix7126 : aoi22 port map ( Y=>nx7125, A0=>que_out_17_4_3, A1=>nx10220, B0
      =>que_out_20_4_3, B1=>nx10194);
   ix543 : nand03 port map ( Y=>nx542, A0=>nx7129, A1=>nx7131, A2=>nx7133);
   ix7130 : aoi222 port map ( Y=>nx7129, A0=>que_out_19_4_3, A1=>nx10168, B0
      =>que_out_21_4_3, B1=>nx10142, C0=>que_out_8_4_3, C1=>nx10116);
   ix7132 : aoi22 port map ( Y=>nx7131, A0=>que_out_25_4_3, A1=>nx10064, B0
      =>que_out_16_4_3, B1=>nx10090);
   ix7134 : aoi22 port map ( Y=>nx7133, A0=>que_out_24_4_3, A1=>nx10038, B0
      =>que_out_22_4_3, B1=>nx10012);
   ix515 : nand03 port map ( Y=>nx514, A0=>nx7137, A1=>nx7139, A2=>nx7141);
   ix7138 : aoi222 port map ( Y=>nx7137, A0=>que_out_15_4_3, A1=>nx9960, B0
      =>que_out_3_4_3, B1=>nx9986, C0=>que_out_23_4_3, C1=>nx9934);
   ix7140 : aoi22 port map ( Y=>nx7139, A0=>que_out_27_4_3, A1=>nx9908, B0=>
      que_out_4_4_3, B1=>nx9882);
   ix7142 : aoi22 port map ( Y=>nx7141, A0=>que_out_0_4_3, A1=>nx9830, B0=>
      que_out_2_4_3, B1=>nx9856);
   ix489 : nand03 port map ( Y=>nx488, A0=>nx7145, A1=>nx7147, A2=>nx7149);
   ix7146 : aoi222 port map ( Y=>nx7145, A0=>que_out_26_4_3, A1=>nx9804, B0
      =>que_out_14_4_3, B1=>nx9778, C0=>que_out_11_4_3, C1=>nx9752);
   ix7148 : aoi22 port map ( Y=>nx7147, A0=>que_out_13_4_3, A1=>nx9726, B0=>
      que_out_7_4_3, B1=>nx9700);
   ix7150 : aoi22 port map ( Y=>nx7149, A0=>que_out_12_4_3, A1=>nx9674, B0=>
      que_out_1_4_3, B1=>nx9648);
   ix683 : or04 port map ( Y=>out_column_4_4, A0=>nx678, A1=>nx652, A2=>
      nx624, A3=>nx598);
   ix679 : nand03 port map ( Y=>nx678, A0=>nx7155, A1=>nx7157, A2=>nx7159);
   ix7156 : aoi222 port map ( Y=>nx7155, A0=>que_out_10_4_4, A1=>nx10298, B0
      =>que_out_6_4_4, B1=>nx10350, C0=>que_out_9_4_4, C1=>nx10324);
   ix7158 : aoi22 port map ( Y=>nx7157, A0=>que_out_5_4_4, A1=>nx10246, B0=>
      que_out_18_4_4, B1=>nx10272);
   ix7160 : aoi22 port map ( Y=>nx7159, A0=>que_out_17_4_4, A1=>nx10220, B0
      =>que_out_20_4_4, B1=>nx10194);
   ix653 : nand03 port map ( Y=>nx652, A0=>nx7163, A1=>nx7165, A2=>nx7167);
   ix7164 : aoi222 port map ( Y=>nx7163, A0=>que_out_19_4_4, A1=>nx10168, B0
      =>que_out_21_4_4, B1=>nx10142, C0=>que_out_8_4_4, C1=>nx10116);
   ix7166 : aoi22 port map ( Y=>nx7165, A0=>que_out_25_4_4, A1=>nx10064, B0
      =>que_out_16_4_4, B1=>nx10090);
   ix7168 : aoi22 port map ( Y=>nx7167, A0=>que_out_24_4_4, A1=>nx10038, B0
      =>que_out_22_4_4, B1=>nx10012);
   ix625 : nand03 port map ( Y=>nx624, A0=>nx7171, A1=>nx7173, A2=>nx7175);
   ix7172 : aoi222 port map ( Y=>nx7171, A0=>que_out_15_4_4, A1=>nx9960, B0
      =>que_out_3_4_4, B1=>nx9986, C0=>que_out_23_4_4, C1=>nx9934);
   ix7174 : aoi22 port map ( Y=>nx7173, A0=>que_out_27_4_4, A1=>nx9908, B0=>
      que_out_4_4_4, B1=>nx9882);
   ix7176 : aoi22 port map ( Y=>nx7175, A0=>que_out_0_4_4, A1=>nx9830, B0=>
      que_out_2_4_4, B1=>nx9856);
   ix599 : nand03 port map ( Y=>nx598, A0=>nx7179, A1=>nx7181, A2=>nx7183);
   ix7180 : aoi222 port map ( Y=>nx7179, A0=>que_out_26_4_4, A1=>nx9804, B0
      =>que_out_14_4_4, B1=>nx9778, C0=>que_out_11_4_4, C1=>nx9752);
   ix7182 : aoi22 port map ( Y=>nx7181, A0=>que_out_13_4_4, A1=>nx9726, B0=>
      que_out_7_4_4, B1=>nx9700);
   ix7184 : aoi22 port map ( Y=>nx7183, A0=>que_out_12_4_4, A1=>nx9674, B0=>
      que_out_1_4_4, B1=>nx9648);
   ix793 : or04 port map ( Y=>out_column_4_5, A0=>nx788, A1=>nx762, A2=>
      nx734, A3=>nx708);
   ix789 : nand03 port map ( Y=>nx788, A0=>nx7189, A1=>nx7191, A2=>nx7193);
   ix7190 : aoi222 port map ( Y=>nx7189, A0=>que_out_10_4_5, A1=>nx10298, B0
      =>que_out_6_4_5, B1=>nx10350, C0=>que_out_9_4_5, C1=>nx10324);
   ix7192 : aoi22 port map ( Y=>nx7191, A0=>que_out_5_4_5, A1=>nx10246, B0=>
      que_out_18_4_5, B1=>nx10272);
   ix7194 : aoi22 port map ( Y=>nx7193, A0=>que_out_17_4_5, A1=>nx10220, B0
      =>que_out_20_4_5, B1=>nx10194);
   ix763 : nand03 port map ( Y=>nx762, A0=>nx7197, A1=>nx7199, A2=>nx7201);
   ix7198 : aoi222 port map ( Y=>nx7197, A0=>que_out_19_4_5, A1=>nx10168, B0
      =>que_out_21_4_5, B1=>nx10142, C0=>que_out_8_4_5, C1=>nx10116);
   ix7200 : aoi22 port map ( Y=>nx7199, A0=>que_out_25_4_5, A1=>nx10064, B0
      =>que_out_16_4_5, B1=>nx10090);
   ix7202 : aoi22 port map ( Y=>nx7201, A0=>que_out_24_4_5, A1=>nx10038, B0
      =>que_out_22_4_5, B1=>nx10012);
   ix735 : nand03 port map ( Y=>nx734, A0=>nx7205, A1=>nx7207, A2=>nx7209);
   ix7206 : aoi222 port map ( Y=>nx7205, A0=>que_out_15_4_5, A1=>nx9960, B0
      =>que_out_3_4_5, B1=>nx9986, C0=>que_out_23_4_5, C1=>nx9934);
   ix7208 : aoi22 port map ( Y=>nx7207, A0=>que_out_27_4_5, A1=>nx9908, B0=>
      que_out_4_4_5, B1=>nx9882);
   ix7210 : aoi22 port map ( Y=>nx7209, A0=>que_out_0_4_5, A1=>nx9830, B0=>
      que_out_2_4_5, B1=>nx9856);
   ix709 : nand03 port map ( Y=>nx708, A0=>nx7213, A1=>nx7215, A2=>nx7217);
   ix7214 : aoi222 port map ( Y=>nx7213, A0=>que_out_26_4_5, A1=>nx9804, B0
      =>que_out_14_4_5, B1=>nx9778, C0=>que_out_11_4_5, C1=>nx9752);
   ix7216 : aoi22 port map ( Y=>nx7215, A0=>que_out_13_4_5, A1=>nx9726, B0=>
      que_out_7_4_5, B1=>nx9700);
   ix7218 : aoi22 port map ( Y=>nx7217, A0=>que_out_12_4_5, A1=>nx9674, B0=>
      que_out_1_4_5, B1=>nx9648);
   ix903 : or04 port map ( Y=>out_column_4_6, A0=>nx898, A1=>nx872, A2=>
      nx844, A3=>nx818);
   ix899 : nand03 port map ( Y=>nx898, A0=>nx7223, A1=>nx7225, A2=>nx7227);
   ix7224 : aoi222 port map ( Y=>nx7223, A0=>que_out_10_4_6, A1=>nx10298, B0
      =>que_out_6_4_6, B1=>nx10350, C0=>que_out_9_4_6, C1=>nx10324);
   ix7226 : aoi22 port map ( Y=>nx7225, A0=>que_out_5_4_6, A1=>nx10246, B0=>
      que_out_18_4_6, B1=>nx10272);
   ix7228 : aoi22 port map ( Y=>nx7227, A0=>que_out_17_4_6, A1=>nx10220, B0
      =>que_out_20_4_6, B1=>nx10194);
   ix873 : nand03 port map ( Y=>nx872, A0=>nx7231, A1=>nx7233, A2=>nx7235);
   ix7232 : aoi222 port map ( Y=>nx7231, A0=>que_out_19_4_6, A1=>nx10168, B0
      =>que_out_21_4_6, B1=>nx10142, C0=>que_out_8_4_6, C1=>nx10116);
   ix7234 : aoi22 port map ( Y=>nx7233, A0=>que_out_25_4_6, A1=>nx10064, B0
      =>que_out_16_4_6, B1=>nx10090);
   ix7236 : aoi22 port map ( Y=>nx7235, A0=>que_out_24_4_6, A1=>nx10038, B0
      =>que_out_22_4_6, B1=>nx10012);
   ix845 : nand03 port map ( Y=>nx844, A0=>nx7239, A1=>nx7241, A2=>nx7243);
   ix7240 : aoi222 port map ( Y=>nx7239, A0=>que_out_15_4_6, A1=>nx9960, B0
      =>que_out_3_4_6, B1=>nx9986, C0=>que_out_23_4_6, C1=>nx9934);
   ix7242 : aoi22 port map ( Y=>nx7241, A0=>que_out_27_4_6, A1=>nx9908, B0=>
      que_out_4_4_6, B1=>nx9882);
   ix7244 : aoi22 port map ( Y=>nx7243, A0=>que_out_0_4_6, A1=>nx9830, B0=>
      que_out_2_4_6, B1=>nx9856);
   ix819 : nand03 port map ( Y=>nx818, A0=>nx7247, A1=>nx7249, A2=>nx7251);
   ix7248 : aoi222 port map ( Y=>nx7247, A0=>que_out_26_4_6, A1=>nx9804, B0
      =>que_out_14_4_6, B1=>nx9778, C0=>que_out_11_4_6, C1=>nx9752);
   ix7250 : aoi22 port map ( Y=>nx7249, A0=>que_out_13_4_6, A1=>nx9726, B0=>
      que_out_7_4_6, B1=>nx9700);
   ix7252 : aoi22 port map ( Y=>nx7251, A0=>que_out_12_4_6, A1=>nx9674, B0=>
      que_out_1_4_6, B1=>nx9648);
   ix1013 : or04 port map ( Y=>out_column_4_7, A0=>nx1008, A1=>nx982, A2=>
      nx954, A3=>nx928);
   ix1009 : nand03 port map ( Y=>nx1008, A0=>nx7257, A1=>nx7259, A2=>nx7261
   );
   ix7258 : aoi222 port map ( Y=>nx7257, A0=>que_out_10_4_7, A1=>nx10300, B0
      =>que_out_6_4_7, B1=>nx10352, C0=>que_out_9_4_7, C1=>nx10326);
   ix7260 : aoi22 port map ( Y=>nx7259, A0=>que_out_5_4_7, A1=>nx10248, B0=>
      que_out_18_4_7, B1=>nx10274);
   ix7262 : aoi22 port map ( Y=>nx7261, A0=>que_out_17_4_7, A1=>nx10222, B0
      =>que_out_20_4_7, B1=>nx10196);
   ix983 : nand03 port map ( Y=>nx982, A0=>nx7265, A1=>nx7267, A2=>nx7269);
   ix7266 : aoi222 port map ( Y=>nx7265, A0=>que_out_19_4_7, A1=>nx10170, B0
      =>que_out_21_4_7, B1=>nx10144, C0=>que_out_8_4_7, C1=>nx10118);
   ix7268 : aoi22 port map ( Y=>nx7267, A0=>que_out_25_4_7, A1=>nx10066, B0
      =>que_out_16_4_7, B1=>nx10092);
   ix7270 : aoi22 port map ( Y=>nx7269, A0=>que_out_24_4_7, A1=>nx10040, B0
      =>que_out_22_4_7, B1=>nx10014);
   ix955 : nand03 port map ( Y=>nx954, A0=>nx7273, A1=>nx7275, A2=>nx7277);
   ix7274 : aoi222 port map ( Y=>nx7273, A0=>que_out_15_4_7, A1=>nx9962, B0
      =>que_out_3_4_7, B1=>nx9988, C0=>que_out_23_4_7, C1=>nx9936);
   ix7276 : aoi22 port map ( Y=>nx7275, A0=>que_out_27_4_7, A1=>nx9910, B0=>
      que_out_4_4_7, B1=>nx9884);
   ix7278 : aoi22 port map ( Y=>nx7277, A0=>que_out_0_4_7, A1=>nx9832, B0=>
      que_out_2_4_7, B1=>nx9858);
   ix929 : nand03 port map ( Y=>nx928, A0=>nx7281, A1=>nx7283, A2=>nx7285);
   ix7282 : aoi222 port map ( Y=>nx7281, A0=>que_out_26_4_7, A1=>nx9806, B0
      =>que_out_14_4_7, B1=>nx9780, C0=>que_out_11_4_7, C1=>nx9754);
   ix7284 : aoi22 port map ( Y=>nx7283, A0=>que_out_13_4_7, A1=>nx9728, B0=>
      que_out_7_4_7, B1=>nx9702);
   ix7286 : aoi22 port map ( Y=>nx7285, A0=>que_out_12_4_7, A1=>nx9676, B0=>
      que_out_1_4_7, B1=>nx9650);
   ix1123 : or04 port map ( Y=>out_column_4_8, A0=>nx1118, A1=>nx1092, A2=>
      nx1064, A3=>nx1038);
   ix1119 : nand03 port map ( Y=>nx1118, A0=>nx7291, A1=>nx7293, A2=>nx7295
   );
   ix7292 : aoi222 port map ( Y=>nx7291, A0=>que_out_10_4_8, A1=>nx10300, B0
      =>que_out_6_4_8, B1=>nx10352, C0=>que_out_9_4_8, C1=>nx10326);
   ix7294 : aoi22 port map ( Y=>nx7293, A0=>que_out_5_4_8, A1=>nx10248, B0=>
      que_out_18_4_8, B1=>nx10274);
   ix7296 : aoi22 port map ( Y=>nx7295, A0=>que_out_17_4_8, A1=>nx10222, B0
      =>que_out_20_4_8, B1=>nx10196);
   ix1093 : nand03 port map ( Y=>nx1092, A0=>nx7299, A1=>nx7301, A2=>nx7303
   );
   ix7300 : aoi222 port map ( Y=>nx7299, A0=>que_out_19_4_8, A1=>nx10170, B0
      =>que_out_21_4_8, B1=>nx10144, C0=>que_out_8_4_8, C1=>nx10118);
   ix7302 : aoi22 port map ( Y=>nx7301, A0=>que_out_25_4_8, A1=>nx10066, B0
      =>que_out_16_4_8, B1=>nx10092);
   ix7304 : aoi22 port map ( Y=>nx7303, A0=>que_out_24_4_8, A1=>nx10040, B0
      =>que_out_22_4_8, B1=>nx10014);
   ix1065 : nand03 port map ( Y=>nx1064, A0=>nx7307, A1=>nx7309, A2=>nx7311
   );
   ix7308 : aoi222 port map ( Y=>nx7307, A0=>que_out_15_4_8, A1=>nx9962, B0
      =>que_out_3_4_8, B1=>nx9988, C0=>que_out_23_4_8, C1=>nx9936);
   ix7310 : aoi22 port map ( Y=>nx7309, A0=>que_out_27_4_8, A1=>nx9910, B0=>
      que_out_4_4_8, B1=>nx9884);
   ix7312 : aoi22 port map ( Y=>nx7311, A0=>que_out_0_4_8, A1=>nx9832, B0=>
      que_out_2_4_8, B1=>nx9858);
   ix1039 : nand03 port map ( Y=>nx1038, A0=>nx7315, A1=>nx7317, A2=>nx7319
   );
   ix7316 : aoi222 port map ( Y=>nx7315, A0=>que_out_26_4_8, A1=>nx9806, B0
      =>que_out_14_4_8, B1=>nx9780, C0=>que_out_11_4_8, C1=>nx9754);
   ix7318 : aoi22 port map ( Y=>nx7317, A0=>que_out_13_4_8, A1=>nx9728, B0=>
      que_out_7_4_8, B1=>nx9702);
   ix7320 : aoi22 port map ( Y=>nx7319, A0=>que_out_12_4_8, A1=>nx9676, B0=>
      que_out_1_4_8, B1=>nx9650);
   ix1233 : or04 port map ( Y=>out_column_4_9, A0=>nx1228, A1=>nx1202, A2=>
      nx1174, A3=>nx1148);
   ix1229 : nand03 port map ( Y=>nx1228, A0=>nx7325, A1=>nx7327, A2=>nx7329
   );
   ix7326 : aoi222 port map ( Y=>nx7325, A0=>que_out_10_4_9, A1=>nx10300, B0
      =>que_out_6_4_9, B1=>nx10352, C0=>que_out_9_4_9, C1=>nx10326);
   ix7328 : aoi22 port map ( Y=>nx7327, A0=>que_out_5_4_9, A1=>nx10248, B0=>
      que_out_18_4_9, B1=>nx10274);
   ix7330 : aoi22 port map ( Y=>nx7329, A0=>que_out_17_4_9, A1=>nx10222, B0
      =>que_out_20_4_9, B1=>nx10196);
   ix1203 : nand03 port map ( Y=>nx1202, A0=>nx7333, A1=>nx7335, A2=>nx7337
   );
   ix7334 : aoi222 port map ( Y=>nx7333, A0=>que_out_19_4_9, A1=>nx10170, B0
      =>que_out_21_4_9, B1=>nx10144, C0=>que_out_8_4_9, C1=>nx10118);
   ix7336 : aoi22 port map ( Y=>nx7335, A0=>que_out_25_4_9, A1=>nx10066, B0
      =>que_out_16_4_9, B1=>nx10092);
   ix7338 : aoi22 port map ( Y=>nx7337, A0=>que_out_24_4_9, A1=>nx10040, B0
      =>que_out_22_4_9, B1=>nx10014);
   ix1175 : nand03 port map ( Y=>nx1174, A0=>nx7341, A1=>nx7343, A2=>nx7345
   );
   ix7342 : aoi222 port map ( Y=>nx7341, A0=>que_out_15_4_9, A1=>nx9962, B0
      =>que_out_3_4_9, B1=>nx9988, C0=>que_out_23_4_9, C1=>nx9936);
   ix7344 : aoi22 port map ( Y=>nx7343, A0=>que_out_27_4_9, A1=>nx9910, B0=>
      que_out_4_4_9, B1=>nx9884);
   ix7346 : aoi22 port map ( Y=>nx7345, A0=>que_out_0_4_9, A1=>nx9832, B0=>
      que_out_2_4_9, B1=>nx9858);
   ix1149 : nand03 port map ( Y=>nx1148, A0=>nx7349, A1=>nx7351, A2=>nx7353
   );
   ix7350 : aoi222 port map ( Y=>nx7349, A0=>que_out_26_4_9, A1=>nx9806, B0
      =>que_out_14_4_9, B1=>nx9780, C0=>que_out_11_4_9, C1=>nx9754);
   ix7352 : aoi22 port map ( Y=>nx7351, A0=>que_out_13_4_9, A1=>nx9728, B0=>
      que_out_7_4_9, B1=>nx9702);
   ix7354 : aoi22 port map ( Y=>nx7353, A0=>que_out_12_4_9, A1=>nx9676, B0=>
      que_out_1_4_9, B1=>nx9650);
   ix1343 : or04 port map ( Y=>out_column_4_10, A0=>nx1338, A1=>nx1312, A2=>
      nx1284, A3=>nx1258);
   ix1339 : nand03 port map ( Y=>nx1338, A0=>nx7359, A1=>nx7361, A2=>nx7363
   );
   ix7360 : aoi222 port map ( Y=>nx7359, A0=>que_out_10_4_10, A1=>nx10300, 
      B0=>que_out_6_4_10, B1=>nx10352, C0=>que_out_9_4_10, C1=>nx10326);
   ix7362 : aoi22 port map ( Y=>nx7361, A0=>que_out_5_4_10, A1=>nx10248, B0
      =>que_out_18_4_10, B1=>nx10274);
   ix7364 : aoi22 port map ( Y=>nx7363, A0=>que_out_17_4_10, A1=>nx10222, B0
      =>que_out_20_4_10, B1=>nx10196);
   ix1313 : nand03 port map ( Y=>nx1312, A0=>nx7367, A1=>nx7369, A2=>nx7371
   );
   ix7368 : aoi222 port map ( Y=>nx7367, A0=>que_out_19_4_10, A1=>nx10170, 
      B0=>que_out_21_4_10, B1=>nx10144, C0=>que_out_8_4_10, C1=>nx10118);
   ix7370 : aoi22 port map ( Y=>nx7369, A0=>que_out_25_4_10, A1=>nx10066, B0
      =>que_out_16_4_10, B1=>nx10092);
   ix7372 : aoi22 port map ( Y=>nx7371, A0=>que_out_24_4_10, A1=>nx10040, B0
      =>que_out_22_4_10, B1=>nx10014);
   ix1285 : nand03 port map ( Y=>nx1284, A0=>nx7375, A1=>nx7377, A2=>nx7379
   );
   ix7376 : aoi222 port map ( Y=>nx7375, A0=>que_out_15_4_10, A1=>nx9962, B0
      =>que_out_3_4_10, B1=>nx9988, C0=>que_out_23_4_10, C1=>nx9936);
   ix7378 : aoi22 port map ( Y=>nx7377, A0=>que_out_27_4_10, A1=>nx9910, B0
      =>que_out_4_4_10, B1=>nx9884);
   ix7380 : aoi22 port map ( Y=>nx7379, A0=>que_out_0_4_10, A1=>nx9832, B0=>
      que_out_2_4_10, B1=>nx9858);
   ix1259 : nand03 port map ( Y=>nx1258, A0=>nx7383, A1=>nx7385, A2=>nx7387
   );
   ix7384 : aoi222 port map ( Y=>nx7383, A0=>que_out_26_4_10, A1=>nx9806, B0
      =>que_out_14_4_10, B1=>nx9780, C0=>que_out_11_4_10, C1=>nx9754);
   ix7386 : aoi22 port map ( Y=>nx7385, A0=>que_out_13_4_10, A1=>nx9728, B0
      =>que_out_7_4_10, B1=>nx9702);
   ix7388 : aoi22 port map ( Y=>nx7387, A0=>que_out_12_4_10, A1=>nx9676, B0
      =>que_out_1_4_10, B1=>nx9650);
   ix1453 : or04 port map ( Y=>out_column_4_11, A0=>nx1448, A1=>nx1422, A2=>
      nx1394, A3=>nx1368);
   ix1449 : nand03 port map ( Y=>nx1448, A0=>nx7393, A1=>nx7395, A2=>nx7397
   );
   ix7394 : aoi222 port map ( Y=>nx7393, A0=>que_out_10_4_11, A1=>nx10300, 
      B0=>que_out_6_4_11, B1=>nx10352, C0=>que_out_9_4_11, C1=>nx10326);
   ix7396 : aoi22 port map ( Y=>nx7395, A0=>que_out_5_4_11, A1=>nx10248, B0
      =>que_out_18_4_11, B1=>nx10274);
   ix7398 : aoi22 port map ( Y=>nx7397, A0=>que_out_17_4_11, A1=>nx10222, B0
      =>que_out_20_4_11, B1=>nx10196);
   ix1423 : nand03 port map ( Y=>nx1422, A0=>nx7401, A1=>nx7403, A2=>nx7405
   );
   ix7402 : aoi222 port map ( Y=>nx7401, A0=>que_out_19_4_11, A1=>nx10170, 
      B0=>que_out_21_4_11, B1=>nx10144, C0=>que_out_8_4_11, C1=>nx10118);
   ix7404 : aoi22 port map ( Y=>nx7403, A0=>que_out_25_4_11, A1=>nx10066, B0
      =>que_out_16_4_11, B1=>nx10092);
   ix7406 : aoi22 port map ( Y=>nx7405, A0=>que_out_24_4_11, A1=>nx10040, B0
      =>que_out_22_4_11, B1=>nx10014);
   ix1395 : nand03 port map ( Y=>nx1394, A0=>nx7409, A1=>nx7411, A2=>nx7413
   );
   ix7410 : aoi222 port map ( Y=>nx7409, A0=>que_out_15_4_11, A1=>nx9962, B0
      =>que_out_3_4_11, B1=>nx9988, C0=>que_out_23_4_11, C1=>nx9936);
   ix7412 : aoi22 port map ( Y=>nx7411, A0=>que_out_27_4_11, A1=>nx9910, B0
      =>que_out_4_4_11, B1=>nx9884);
   ix7414 : aoi22 port map ( Y=>nx7413, A0=>que_out_0_4_11, A1=>nx9832, B0=>
      que_out_2_4_11, B1=>nx9858);
   ix1369 : nand03 port map ( Y=>nx1368, A0=>nx7417, A1=>nx7419, A2=>nx7421
   );
   ix7418 : aoi222 port map ( Y=>nx7417, A0=>que_out_26_4_11, A1=>nx9806, B0
      =>que_out_14_4_11, B1=>nx9780, C0=>que_out_11_4_11, C1=>nx9754);
   ix7420 : aoi22 port map ( Y=>nx7419, A0=>que_out_13_4_11, A1=>nx9728, B0
      =>que_out_7_4_11, B1=>nx9702);
   ix7422 : aoi22 port map ( Y=>nx7421, A0=>que_out_12_4_11, A1=>nx9676, B0
      =>que_out_1_4_11, B1=>nx9650);
   ix1563 : or04 port map ( Y=>out_column_4_12, A0=>nx1558, A1=>nx1532, A2=>
      nx1504, A3=>nx1478);
   ix1559 : nand03 port map ( Y=>nx1558, A0=>nx7427, A1=>nx7429, A2=>nx7431
   );
   ix7428 : aoi222 port map ( Y=>nx7427, A0=>que_out_10_4_12, A1=>nx10300, 
      B0=>que_out_6_4_12, B1=>nx10352, C0=>que_out_9_4_12, C1=>nx10326);
   ix7430 : aoi22 port map ( Y=>nx7429, A0=>que_out_5_4_12, A1=>nx10248, B0
      =>que_out_18_4_12, B1=>nx10274);
   ix7432 : aoi22 port map ( Y=>nx7431, A0=>que_out_17_4_12, A1=>nx10222, B0
      =>que_out_20_4_12, B1=>nx10196);
   ix1533 : nand03 port map ( Y=>nx1532, A0=>nx7435, A1=>nx7437, A2=>nx7439
   );
   ix7436 : aoi222 port map ( Y=>nx7435, A0=>que_out_19_4_12, A1=>nx10170, 
      B0=>que_out_21_4_12, B1=>nx10144, C0=>que_out_8_4_12, C1=>nx10118);
   ix7438 : aoi22 port map ( Y=>nx7437, A0=>que_out_25_4_12, A1=>nx10066, B0
      =>que_out_16_4_12, B1=>nx10092);
   ix7440 : aoi22 port map ( Y=>nx7439, A0=>que_out_24_4_12, A1=>nx10040, B0
      =>que_out_22_4_12, B1=>nx10014);
   ix1505 : nand03 port map ( Y=>nx1504, A0=>nx7443, A1=>nx7445, A2=>nx7447
   );
   ix7444 : aoi222 port map ( Y=>nx7443, A0=>que_out_15_4_12, A1=>nx9962, B0
      =>que_out_3_4_12, B1=>nx9988, C0=>que_out_23_4_12, C1=>nx9936);
   ix7446 : aoi22 port map ( Y=>nx7445, A0=>que_out_27_4_12, A1=>nx9910, B0
      =>que_out_4_4_12, B1=>nx9884);
   ix7448 : aoi22 port map ( Y=>nx7447, A0=>que_out_0_4_12, A1=>nx9832, B0=>
      que_out_2_4_12, B1=>nx9858);
   ix1479 : nand03 port map ( Y=>nx1478, A0=>nx7451, A1=>nx7453, A2=>nx7455
   );
   ix7452 : aoi222 port map ( Y=>nx7451, A0=>que_out_26_4_12, A1=>nx9806, B0
      =>que_out_14_4_12, B1=>nx9780, C0=>que_out_11_4_12, C1=>nx9754);
   ix7454 : aoi22 port map ( Y=>nx7453, A0=>que_out_13_4_12, A1=>nx9728, B0
      =>que_out_7_4_12, B1=>nx9702);
   ix7456 : aoi22 port map ( Y=>nx7455, A0=>que_out_12_4_12, A1=>nx9676, B0
      =>que_out_1_4_12, B1=>nx9650);
   ix1673 : or04 port map ( Y=>out_column_4_13, A0=>nx1668, A1=>nx1642, A2=>
      nx1614, A3=>nx1588);
   ix1669 : nand03 port map ( Y=>nx1668, A0=>nx7461, A1=>nx7463, A2=>nx7465
   );
   ix7462 : aoi222 port map ( Y=>nx7461, A0=>que_out_10_4_13, A1=>nx10300, 
      B0=>que_out_6_4_13, B1=>nx10352, C0=>que_out_9_4_13, C1=>nx10326);
   ix7464 : aoi22 port map ( Y=>nx7463, A0=>que_out_5_4_13, A1=>nx10248, B0
      =>que_out_18_4_13, B1=>nx10274);
   ix7466 : aoi22 port map ( Y=>nx7465, A0=>que_out_17_4_13, A1=>nx10222, B0
      =>que_out_20_4_13, B1=>nx10196);
   ix1643 : nand03 port map ( Y=>nx1642, A0=>nx7469, A1=>nx7471, A2=>nx7473
   );
   ix7470 : aoi222 port map ( Y=>nx7469, A0=>que_out_19_4_13, A1=>nx10170, 
      B0=>que_out_21_4_13, B1=>nx10144, C0=>que_out_8_4_13, C1=>nx10118);
   ix7472 : aoi22 port map ( Y=>nx7471, A0=>que_out_25_4_13, A1=>nx10066, B0
      =>que_out_16_4_13, B1=>nx10092);
   ix7474 : aoi22 port map ( Y=>nx7473, A0=>que_out_24_4_13, A1=>nx10040, B0
      =>que_out_22_4_13, B1=>nx10014);
   ix1615 : nand03 port map ( Y=>nx1614, A0=>nx7477, A1=>nx7479, A2=>nx7481
   );
   ix7478 : aoi222 port map ( Y=>nx7477, A0=>que_out_15_4_13, A1=>nx9962, B0
      =>que_out_3_4_13, B1=>nx9988, C0=>que_out_23_4_13, C1=>nx9936);
   ix7480 : aoi22 port map ( Y=>nx7479, A0=>que_out_27_4_13, A1=>nx9910, B0
      =>que_out_4_4_13, B1=>nx9884);
   ix7482 : aoi22 port map ( Y=>nx7481, A0=>que_out_0_4_13, A1=>nx9832, B0=>
      que_out_2_4_13, B1=>nx9858);
   ix1589 : nand03 port map ( Y=>nx1588, A0=>nx7485, A1=>nx7487, A2=>nx7489
   );
   ix7486 : aoi222 port map ( Y=>nx7485, A0=>que_out_26_4_13, A1=>nx9806, B0
      =>que_out_14_4_13, B1=>nx9780, C0=>que_out_11_4_13, C1=>nx9754);
   ix7488 : aoi22 port map ( Y=>nx7487, A0=>que_out_13_4_13, A1=>nx9728, B0
      =>que_out_7_4_13, B1=>nx9702);
   ix7490 : aoi22 port map ( Y=>nx7489, A0=>que_out_12_4_13, A1=>nx9676, B0
      =>que_out_1_4_13, B1=>nx9650);
   ix1783 : or04 port map ( Y=>out_column_4_14, A0=>nx1778, A1=>nx1752, A2=>
      nx1724, A3=>nx1698);
   ix1779 : nand03 port map ( Y=>nx1778, A0=>nx7495, A1=>nx7497, A2=>nx7499
   );
   ix7496 : aoi222 port map ( Y=>nx7495, A0=>que_out_10_4_14, A1=>nx10302, 
      B0=>que_out_6_4_14, B1=>nx10354, C0=>que_out_9_4_14, C1=>nx10328);
   ix7498 : aoi22 port map ( Y=>nx7497, A0=>que_out_5_4_14, A1=>nx10250, B0
      =>que_out_18_4_14, B1=>nx10276);
   ix7500 : aoi22 port map ( Y=>nx7499, A0=>que_out_17_4_14, A1=>nx10224, B0
      =>que_out_20_4_14, B1=>nx10198);
   ix1753 : nand03 port map ( Y=>nx1752, A0=>nx7503, A1=>nx7505, A2=>nx7507
   );
   ix7504 : aoi222 port map ( Y=>nx7503, A0=>que_out_19_4_14, A1=>nx10172, 
      B0=>que_out_21_4_14, B1=>nx10146, C0=>que_out_8_4_14, C1=>nx10120);
   ix7506 : aoi22 port map ( Y=>nx7505, A0=>que_out_25_4_14, A1=>nx10068, B0
      =>que_out_16_4_14, B1=>nx10094);
   ix7508 : aoi22 port map ( Y=>nx7507, A0=>que_out_24_4_14, A1=>nx10042, B0
      =>que_out_22_4_14, B1=>nx10016);
   ix1725 : nand03 port map ( Y=>nx1724, A0=>nx7511, A1=>nx7513, A2=>nx7515
   );
   ix7512 : aoi222 port map ( Y=>nx7511, A0=>que_out_15_4_14, A1=>nx9964, B0
      =>que_out_3_4_14, B1=>nx9990, C0=>que_out_23_4_14, C1=>nx9938);
   ix7514 : aoi22 port map ( Y=>nx7513, A0=>que_out_27_4_14, A1=>nx9912, B0
      =>que_out_4_4_14, B1=>nx9886);
   ix7516 : aoi22 port map ( Y=>nx7515, A0=>que_out_0_4_14, A1=>nx9834, B0=>
      que_out_2_4_14, B1=>nx9860);
   ix1699 : nand03 port map ( Y=>nx1698, A0=>nx7519, A1=>nx7521, A2=>nx7523
   );
   ix7520 : aoi222 port map ( Y=>nx7519, A0=>que_out_26_4_14, A1=>nx9808, B0
      =>que_out_14_4_14, B1=>nx9782, C0=>que_out_11_4_14, C1=>nx9756);
   ix7522 : aoi22 port map ( Y=>nx7521, A0=>que_out_13_4_14, A1=>nx9730, B0
      =>que_out_7_4_14, B1=>nx9704);
   ix7524 : aoi22 port map ( Y=>nx7523, A0=>que_out_12_4_14, A1=>nx9678, B0
      =>que_out_1_4_14, B1=>nx9652);
   ix1893 : or04 port map ( Y=>out_column_4_15, A0=>nx1888, A1=>nx1862, A2=>
      nx1834, A3=>nx1808);
   ix1889 : nand03 port map ( Y=>nx1888, A0=>nx7529, A1=>nx7531, A2=>nx7533
   );
   ix7530 : aoi222 port map ( Y=>nx7529, A0=>que_out_10_4_15, A1=>nx10302, 
      B0=>que_out_6_4_15, B1=>nx10354, C0=>que_out_9_4_15, C1=>nx10328);
   ix7532 : aoi22 port map ( Y=>nx7531, A0=>que_out_5_4_15, A1=>nx10250, B0
      =>que_out_18_4_15, B1=>nx10276);
   ix7534 : aoi22 port map ( Y=>nx7533, A0=>que_out_17_4_15, A1=>nx10224, B0
      =>que_out_20_4_15, B1=>nx10198);
   ix1863 : nand03 port map ( Y=>nx1862, A0=>nx7537, A1=>nx7539, A2=>nx7541
   );
   ix7538 : aoi222 port map ( Y=>nx7537, A0=>que_out_19_4_15, A1=>nx10172, 
      B0=>que_out_21_4_15, B1=>nx10146, C0=>que_out_8_4_15, C1=>nx10120);
   ix7540 : aoi22 port map ( Y=>nx7539, A0=>que_out_25_4_15, A1=>nx10068, B0
      =>que_out_16_4_15, B1=>nx10094);
   ix7542 : aoi22 port map ( Y=>nx7541, A0=>que_out_24_4_15, A1=>nx10042, B0
      =>que_out_22_4_15, B1=>nx10016);
   ix1835 : nand03 port map ( Y=>nx1834, A0=>nx7545, A1=>nx7547, A2=>nx7549
   );
   ix7546 : aoi222 port map ( Y=>nx7545, A0=>que_out_15_4_15, A1=>nx9964, B0
      =>que_out_3_4_15, B1=>nx9990, C0=>que_out_23_4_15, C1=>nx9938);
   ix7548 : aoi22 port map ( Y=>nx7547, A0=>que_out_27_4_15, A1=>nx9912, B0
      =>que_out_4_4_15, B1=>nx9886);
   ix7550 : aoi22 port map ( Y=>nx7549, A0=>que_out_0_4_15, A1=>nx9834, B0=>
      que_out_2_4_15, B1=>nx9860);
   ix1809 : nand03 port map ( Y=>nx1808, A0=>nx7553, A1=>nx7555, A2=>nx7557
   );
   ix7554 : aoi222 port map ( Y=>nx7553, A0=>que_out_26_4_15, A1=>nx9808, B0
      =>que_out_14_4_15, B1=>nx9782, C0=>que_out_11_4_15, C1=>nx9756);
   ix7556 : aoi22 port map ( Y=>nx7555, A0=>que_out_13_4_15, A1=>nx9730, B0
      =>que_out_7_4_15, B1=>nx9704);
   ix7558 : aoi22 port map ( Y=>nx7557, A0=>que_out_12_4_15, A1=>nx9678, B0
      =>que_out_1_4_15, B1=>nx9652);
   ix2003 : or04 port map ( Y=>out_column_3_0, A0=>nx1998, A1=>nx1972, A2=>
      nx1944, A3=>nx1918);
   ix1999 : nand03 port map ( Y=>nx1998, A0=>nx7563, A1=>nx7565, A2=>nx7567
   );
   ix7564 : aoi222 port map ( Y=>nx7563, A0=>que_out_10_3_0, A1=>nx10302, B0
      =>que_out_6_3_0, B1=>nx10354, C0=>que_out_9_3_0, C1=>nx10328);
   ix7566 : aoi22 port map ( Y=>nx7565, A0=>que_out_5_3_0, A1=>nx10250, B0=>
      que_out_18_3_0, B1=>nx10276);
   ix7568 : aoi22 port map ( Y=>nx7567, A0=>que_out_17_3_0, A1=>nx10224, B0
      =>que_out_20_3_0, B1=>nx10198);
   ix1973 : nand03 port map ( Y=>nx1972, A0=>nx7571, A1=>nx7573, A2=>nx7575
   );
   ix7572 : aoi222 port map ( Y=>nx7571, A0=>que_out_19_3_0, A1=>nx10172, B0
      =>que_out_21_3_0, B1=>nx10146, C0=>que_out_8_3_0, C1=>nx10120);
   ix7574 : aoi22 port map ( Y=>nx7573, A0=>que_out_25_3_0, A1=>nx10068, B0
      =>que_out_16_3_0, B1=>nx10094);
   ix7576 : aoi22 port map ( Y=>nx7575, A0=>que_out_24_3_0, A1=>nx10042, B0
      =>que_out_22_3_0, B1=>nx10016);
   ix1945 : nand03 port map ( Y=>nx1944, A0=>nx7579, A1=>nx7581, A2=>nx7583
   );
   ix7580 : aoi222 port map ( Y=>nx7579, A0=>que_out_15_3_0, A1=>nx9964, B0
      =>que_out_3_3_0, B1=>nx9990, C0=>que_out_23_3_0, C1=>nx9938);
   ix7582 : aoi22 port map ( Y=>nx7581, A0=>que_out_27_3_0, A1=>nx9912, B0=>
      que_out_4_3_0, B1=>nx9886);
   ix7584 : aoi22 port map ( Y=>nx7583, A0=>que_out_0_3_0, A1=>nx9834, B0=>
      que_out_2_3_0, B1=>nx9860);
   ix1919 : nand03 port map ( Y=>nx1918, A0=>nx7587, A1=>nx7589, A2=>nx7591
   );
   ix7588 : aoi222 port map ( Y=>nx7587, A0=>que_out_26_3_0, A1=>nx9808, B0
      =>que_out_14_3_0, B1=>nx9782, C0=>que_out_11_3_0, C1=>nx9756);
   ix7590 : aoi22 port map ( Y=>nx7589, A0=>que_out_13_3_0, A1=>nx9730, B0=>
      que_out_7_3_0, B1=>nx9704);
   ix7592 : aoi22 port map ( Y=>nx7591, A0=>que_out_12_3_0, A1=>nx9678, B0=>
      que_out_1_3_0, B1=>nx9652);
   ix2113 : or04 port map ( Y=>out_column_3_1, A0=>nx2108, A1=>nx2082, A2=>
      nx2054, A3=>nx2028);
   ix2109 : nand03 port map ( Y=>nx2108, A0=>nx7597, A1=>nx7599, A2=>nx7601
   );
   ix7598 : aoi222 port map ( Y=>nx7597, A0=>que_out_10_3_1, A1=>nx10302, B0
      =>que_out_6_3_1, B1=>nx10354, C0=>que_out_9_3_1, C1=>nx10328);
   ix7600 : aoi22 port map ( Y=>nx7599, A0=>que_out_5_3_1, A1=>nx10250, B0=>
      que_out_18_3_1, B1=>nx10276);
   ix7602 : aoi22 port map ( Y=>nx7601, A0=>que_out_17_3_1, A1=>nx10224, B0
      =>que_out_20_3_1, B1=>nx10198);
   ix2083 : nand03 port map ( Y=>nx2082, A0=>nx7605, A1=>nx7607, A2=>nx7609
   );
   ix7606 : aoi222 port map ( Y=>nx7605, A0=>que_out_19_3_1, A1=>nx10172, B0
      =>que_out_21_3_1, B1=>nx10146, C0=>que_out_8_3_1, C1=>nx10120);
   ix7608 : aoi22 port map ( Y=>nx7607, A0=>que_out_25_3_1, A1=>nx10068, B0
      =>que_out_16_3_1, B1=>nx10094);
   ix7610 : aoi22 port map ( Y=>nx7609, A0=>que_out_24_3_1, A1=>nx10042, B0
      =>que_out_22_3_1, B1=>nx10016);
   ix2055 : nand03 port map ( Y=>nx2054, A0=>nx7613, A1=>nx7615, A2=>nx7617
   );
   ix7614 : aoi222 port map ( Y=>nx7613, A0=>que_out_15_3_1, A1=>nx9964, B0
      =>que_out_3_3_1, B1=>nx9990, C0=>que_out_23_3_1, C1=>nx9938);
   ix7616 : aoi22 port map ( Y=>nx7615, A0=>que_out_27_3_1, A1=>nx9912, B0=>
      que_out_4_3_1, B1=>nx9886);
   ix7618 : aoi22 port map ( Y=>nx7617, A0=>que_out_0_3_1, A1=>nx9834, B0=>
      que_out_2_3_1, B1=>nx9860);
   ix2029 : nand03 port map ( Y=>nx2028, A0=>nx7621, A1=>nx7623, A2=>nx7625
   );
   ix7622 : aoi222 port map ( Y=>nx7621, A0=>que_out_26_3_1, A1=>nx9808, B0
      =>que_out_14_3_1, B1=>nx9782, C0=>que_out_11_3_1, C1=>nx9756);
   ix7624 : aoi22 port map ( Y=>nx7623, A0=>que_out_13_3_1, A1=>nx9730, B0=>
      que_out_7_3_1, B1=>nx9704);
   ix7626 : aoi22 port map ( Y=>nx7625, A0=>que_out_12_3_1, A1=>nx9678, B0=>
      que_out_1_3_1, B1=>nx9652);
   ix2223 : or04 port map ( Y=>out_column_3_2, A0=>nx2218, A1=>nx2192, A2=>
      nx2164, A3=>nx2138);
   ix2219 : nand03 port map ( Y=>nx2218, A0=>nx7631, A1=>nx7633, A2=>nx7635
   );
   ix7632 : aoi222 port map ( Y=>nx7631, A0=>que_out_10_3_2, A1=>nx10302, B0
      =>que_out_6_3_2, B1=>nx10354, C0=>que_out_9_3_2, C1=>nx10328);
   ix7634 : aoi22 port map ( Y=>nx7633, A0=>que_out_5_3_2, A1=>nx10250, B0=>
      que_out_18_3_2, B1=>nx10276);
   ix7636 : aoi22 port map ( Y=>nx7635, A0=>que_out_17_3_2, A1=>nx10224, B0
      =>que_out_20_3_2, B1=>nx10198);
   ix2193 : nand03 port map ( Y=>nx2192, A0=>nx7639, A1=>nx7641, A2=>nx7643
   );
   ix7640 : aoi222 port map ( Y=>nx7639, A0=>que_out_19_3_2, A1=>nx10172, B0
      =>que_out_21_3_2, B1=>nx10146, C0=>que_out_8_3_2, C1=>nx10120);
   ix7642 : aoi22 port map ( Y=>nx7641, A0=>que_out_25_3_2, A1=>nx10068, B0
      =>que_out_16_3_2, B1=>nx10094);
   ix7644 : aoi22 port map ( Y=>nx7643, A0=>que_out_24_3_2, A1=>nx10042, B0
      =>que_out_22_3_2, B1=>nx10016);
   ix2165 : nand03 port map ( Y=>nx2164, A0=>nx7647, A1=>nx7649, A2=>nx7651
   );
   ix7648 : aoi222 port map ( Y=>nx7647, A0=>que_out_15_3_2, A1=>nx9964, B0
      =>que_out_3_3_2, B1=>nx9990, C0=>que_out_23_3_2, C1=>nx9938);
   ix7650 : aoi22 port map ( Y=>nx7649, A0=>que_out_27_3_2, A1=>nx9912, B0=>
      que_out_4_3_2, B1=>nx9886);
   ix7652 : aoi22 port map ( Y=>nx7651, A0=>que_out_0_3_2, A1=>nx9834, B0=>
      que_out_2_3_2, B1=>nx9860);
   ix2139 : nand03 port map ( Y=>nx2138, A0=>nx7655, A1=>nx7657, A2=>nx7659
   );
   ix7656 : aoi222 port map ( Y=>nx7655, A0=>que_out_26_3_2, A1=>nx9808, B0
      =>que_out_14_3_2, B1=>nx9782, C0=>que_out_11_3_2, C1=>nx9756);
   ix7658 : aoi22 port map ( Y=>nx7657, A0=>que_out_13_3_2, A1=>nx9730, B0=>
      que_out_7_3_2, B1=>nx9704);
   ix7660 : aoi22 port map ( Y=>nx7659, A0=>que_out_12_3_2, A1=>nx9678, B0=>
      que_out_1_3_2, B1=>nx9652);
   ix2333 : or04 port map ( Y=>out_column_3_3, A0=>nx2328, A1=>nx2302, A2=>
      nx2274, A3=>nx2248);
   ix2329 : nand03 port map ( Y=>nx2328, A0=>nx7665, A1=>nx7667, A2=>nx7669
   );
   ix7666 : aoi222 port map ( Y=>nx7665, A0=>que_out_10_3_3, A1=>nx10302, B0
      =>que_out_6_3_3, B1=>nx10354, C0=>que_out_9_3_3, C1=>nx10328);
   ix7668 : aoi22 port map ( Y=>nx7667, A0=>que_out_5_3_3, A1=>nx10250, B0=>
      que_out_18_3_3, B1=>nx10276);
   ix7670 : aoi22 port map ( Y=>nx7669, A0=>que_out_17_3_3, A1=>nx10224, B0
      =>que_out_20_3_3, B1=>nx10198);
   ix2303 : nand03 port map ( Y=>nx2302, A0=>nx7673, A1=>nx7675, A2=>nx7677
   );
   ix7674 : aoi222 port map ( Y=>nx7673, A0=>que_out_19_3_3, A1=>nx10172, B0
      =>que_out_21_3_3, B1=>nx10146, C0=>que_out_8_3_3, C1=>nx10120);
   ix7676 : aoi22 port map ( Y=>nx7675, A0=>que_out_25_3_3, A1=>nx10068, B0
      =>que_out_16_3_3, B1=>nx10094);
   ix7678 : aoi22 port map ( Y=>nx7677, A0=>que_out_24_3_3, A1=>nx10042, B0
      =>que_out_22_3_3, B1=>nx10016);
   ix2275 : nand03 port map ( Y=>nx2274, A0=>nx7681, A1=>nx7683, A2=>nx7685
   );
   ix7682 : aoi222 port map ( Y=>nx7681, A0=>que_out_15_3_3, A1=>nx9964, B0
      =>que_out_3_3_3, B1=>nx9990, C0=>que_out_23_3_3, C1=>nx9938);
   ix7684 : aoi22 port map ( Y=>nx7683, A0=>que_out_27_3_3, A1=>nx9912, B0=>
      que_out_4_3_3, B1=>nx9886);
   ix7686 : aoi22 port map ( Y=>nx7685, A0=>que_out_0_3_3, A1=>nx9834, B0=>
      que_out_2_3_3, B1=>nx9860);
   ix2249 : nand03 port map ( Y=>nx2248, A0=>nx7689, A1=>nx7691, A2=>nx7693
   );
   ix7690 : aoi222 port map ( Y=>nx7689, A0=>que_out_26_3_3, A1=>nx9808, B0
      =>que_out_14_3_3, B1=>nx9782, C0=>que_out_11_3_3, C1=>nx9756);
   ix7692 : aoi22 port map ( Y=>nx7691, A0=>que_out_13_3_3, A1=>nx9730, B0=>
      que_out_7_3_3, B1=>nx9704);
   ix7694 : aoi22 port map ( Y=>nx7693, A0=>que_out_12_3_3, A1=>nx9678, B0=>
      que_out_1_3_3, B1=>nx9652);
   ix2443 : or04 port map ( Y=>out_column_3_4, A0=>nx2438, A1=>nx2412, A2=>
      nx2384, A3=>nx2358);
   ix2439 : nand03 port map ( Y=>nx2438, A0=>nx7699, A1=>nx7701, A2=>nx7703
   );
   ix7700 : aoi222 port map ( Y=>nx7699, A0=>que_out_10_3_4, A1=>nx10302, B0
      =>que_out_6_3_4, B1=>nx10354, C0=>que_out_9_3_4, C1=>nx10328);
   ix7702 : aoi22 port map ( Y=>nx7701, A0=>que_out_5_3_4, A1=>nx10250, B0=>
      que_out_18_3_4, B1=>nx10276);
   ix7704 : aoi22 port map ( Y=>nx7703, A0=>que_out_17_3_4, A1=>nx10224, B0
      =>que_out_20_3_4, B1=>nx10198);
   ix2413 : nand03 port map ( Y=>nx2412, A0=>nx7707, A1=>nx7709, A2=>nx7711
   );
   ix7708 : aoi222 port map ( Y=>nx7707, A0=>que_out_19_3_4, A1=>nx10172, B0
      =>que_out_21_3_4, B1=>nx10146, C0=>que_out_8_3_4, C1=>nx10120);
   ix7710 : aoi22 port map ( Y=>nx7709, A0=>que_out_25_3_4, A1=>nx10068, B0
      =>que_out_16_3_4, B1=>nx10094);
   ix7712 : aoi22 port map ( Y=>nx7711, A0=>que_out_24_3_4, A1=>nx10042, B0
      =>que_out_22_3_4, B1=>nx10016);
   ix2385 : nand03 port map ( Y=>nx2384, A0=>nx7715, A1=>nx7717, A2=>nx7719
   );
   ix7716 : aoi222 port map ( Y=>nx7715, A0=>que_out_15_3_4, A1=>nx9964, B0
      =>que_out_3_3_4, B1=>nx9990, C0=>que_out_23_3_4, C1=>nx9938);
   ix7718 : aoi22 port map ( Y=>nx7717, A0=>que_out_27_3_4, A1=>nx9912, B0=>
      que_out_4_3_4, B1=>nx9886);
   ix7720 : aoi22 port map ( Y=>nx7719, A0=>que_out_0_3_4, A1=>nx9834, B0=>
      que_out_2_3_4, B1=>nx9860);
   ix2359 : nand03 port map ( Y=>nx2358, A0=>nx7723, A1=>nx7725, A2=>nx7727
   );
   ix7724 : aoi222 port map ( Y=>nx7723, A0=>que_out_26_3_4, A1=>nx9808, B0
      =>que_out_14_3_4, B1=>nx9782, C0=>que_out_11_3_4, C1=>nx9756);
   ix7726 : aoi22 port map ( Y=>nx7725, A0=>que_out_13_3_4, A1=>nx9730, B0=>
      que_out_7_3_4, B1=>nx9704);
   ix7728 : aoi22 port map ( Y=>nx7727, A0=>que_out_12_3_4, A1=>nx9678, B0=>
      que_out_1_3_4, B1=>nx9652);
   ix2553 : or04 port map ( Y=>out_column_3_5, A0=>nx2548, A1=>nx2522, A2=>
      nx2494, A3=>nx2468);
   ix2549 : nand03 port map ( Y=>nx2548, A0=>nx7733, A1=>nx7735, A2=>nx7737
   );
   ix7734 : aoi222 port map ( Y=>nx7733, A0=>que_out_10_3_5, A1=>nx10304, B0
      =>que_out_6_3_5, B1=>nx10356, C0=>que_out_9_3_5, C1=>nx10330);
   ix7736 : aoi22 port map ( Y=>nx7735, A0=>que_out_5_3_5, A1=>nx10252, B0=>
      que_out_18_3_5, B1=>nx10278);
   ix7738 : aoi22 port map ( Y=>nx7737, A0=>que_out_17_3_5, A1=>nx10226, B0
      =>que_out_20_3_5, B1=>nx10200);
   ix2523 : nand03 port map ( Y=>nx2522, A0=>nx7741, A1=>nx7743, A2=>nx7745
   );
   ix7742 : aoi222 port map ( Y=>nx7741, A0=>que_out_19_3_5, A1=>nx10174, B0
      =>que_out_21_3_5, B1=>nx10148, C0=>que_out_8_3_5, C1=>nx10122);
   ix7744 : aoi22 port map ( Y=>nx7743, A0=>que_out_25_3_5, A1=>nx10070, B0
      =>que_out_16_3_5, B1=>nx10096);
   ix7746 : aoi22 port map ( Y=>nx7745, A0=>que_out_24_3_5, A1=>nx10044, B0
      =>que_out_22_3_5, B1=>nx10018);
   ix2495 : nand03 port map ( Y=>nx2494, A0=>nx7749, A1=>nx7751, A2=>nx7753
   );
   ix7750 : aoi222 port map ( Y=>nx7749, A0=>que_out_15_3_5, A1=>nx9966, B0
      =>que_out_3_3_5, B1=>nx9992, C0=>que_out_23_3_5, C1=>nx9940);
   ix7752 : aoi22 port map ( Y=>nx7751, A0=>que_out_27_3_5, A1=>nx9914, B0=>
      que_out_4_3_5, B1=>nx9888);
   ix7754 : aoi22 port map ( Y=>nx7753, A0=>que_out_0_3_5, A1=>nx9836, B0=>
      que_out_2_3_5, B1=>nx9862);
   ix2469 : nand03 port map ( Y=>nx2468, A0=>nx7757, A1=>nx7759, A2=>nx7761
   );
   ix7758 : aoi222 port map ( Y=>nx7757, A0=>que_out_26_3_5, A1=>nx9810, B0
      =>que_out_14_3_5, B1=>nx9784, C0=>que_out_11_3_5, C1=>nx9758);
   ix7760 : aoi22 port map ( Y=>nx7759, A0=>que_out_13_3_5, A1=>nx9732, B0=>
      que_out_7_3_5, B1=>nx9706);
   ix7762 : aoi22 port map ( Y=>nx7761, A0=>que_out_12_3_5, A1=>nx9680, B0=>
      que_out_1_3_5, B1=>nx9654);
   ix2663 : or04 port map ( Y=>out_column_3_6, A0=>nx2658, A1=>nx2632, A2=>
      nx2604, A3=>nx2578);
   ix2659 : nand03 port map ( Y=>nx2658, A0=>nx7767, A1=>nx7769, A2=>nx7771
   );
   ix7768 : aoi222 port map ( Y=>nx7767, A0=>que_out_10_3_6, A1=>nx10304, B0
      =>que_out_6_3_6, B1=>nx10356, C0=>que_out_9_3_6, C1=>nx10330);
   ix7770 : aoi22 port map ( Y=>nx7769, A0=>que_out_5_3_6, A1=>nx10252, B0=>
      que_out_18_3_6, B1=>nx10278);
   ix7772 : aoi22 port map ( Y=>nx7771, A0=>que_out_17_3_6, A1=>nx10226, B0
      =>que_out_20_3_6, B1=>nx10200);
   ix2633 : nand03 port map ( Y=>nx2632, A0=>nx7775, A1=>nx7777, A2=>nx7779
   );
   ix7776 : aoi222 port map ( Y=>nx7775, A0=>que_out_19_3_6, A1=>nx10174, B0
      =>que_out_21_3_6, B1=>nx10148, C0=>que_out_8_3_6, C1=>nx10122);
   ix7778 : aoi22 port map ( Y=>nx7777, A0=>que_out_25_3_6, A1=>nx10070, B0
      =>que_out_16_3_6, B1=>nx10096);
   ix7780 : aoi22 port map ( Y=>nx7779, A0=>que_out_24_3_6, A1=>nx10044, B0
      =>que_out_22_3_6, B1=>nx10018);
   ix2605 : nand03 port map ( Y=>nx2604, A0=>nx7783, A1=>nx7785, A2=>nx7787
   );
   ix7784 : aoi222 port map ( Y=>nx7783, A0=>que_out_15_3_6, A1=>nx9966, B0
      =>que_out_3_3_6, B1=>nx9992, C0=>que_out_23_3_6, C1=>nx9940);
   ix7786 : aoi22 port map ( Y=>nx7785, A0=>que_out_27_3_6, A1=>nx9914, B0=>
      que_out_4_3_6, B1=>nx9888);
   ix7788 : aoi22 port map ( Y=>nx7787, A0=>que_out_0_3_6, A1=>nx9836, B0=>
      que_out_2_3_6, B1=>nx9862);
   ix2579 : nand03 port map ( Y=>nx2578, A0=>nx7791, A1=>nx7793, A2=>nx7795
   );
   ix7792 : aoi222 port map ( Y=>nx7791, A0=>que_out_26_3_6, A1=>nx9810, B0
      =>que_out_14_3_6, B1=>nx9784, C0=>que_out_11_3_6, C1=>nx9758);
   ix7794 : aoi22 port map ( Y=>nx7793, A0=>que_out_13_3_6, A1=>nx9732, B0=>
      que_out_7_3_6, B1=>nx9706);
   ix7796 : aoi22 port map ( Y=>nx7795, A0=>que_out_12_3_6, A1=>nx9680, B0=>
      que_out_1_3_6, B1=>nx9654);
   ix2773 : or04 port map ( Y=>out_column_3_7, A0=>nx2768, A1=>nx2742, A2=>
      nx2714, A3=>nx2688);
   ix2769 : nand03 port map ( Y=>nx2768, A0=>nx7801, A1=>nx7803, A2=>nx7805
   );
   ix7802 : aoi222 port map ( Y=>nx7801, A0=>que_out_10_3_7, A1=>nx10304, B0
      =>que_out_6_3_7, B1=>nx10356, C0=>que_out_9_3_7, C1=>nx10330);
   ix7804 : aoi22 port map ( Y=>nx7803, A0=>que_out_5_3_7, A1=>nx10252, B0=>
      que_out_18_3_7, B1=>nx10278);
   ix7806 : aoi22 port map ( Y=>nx7805, A0=>que_out_17_3_7, A1=>nx10226, B0
      =>que_out_20_3_7, B1=>nx10200);
   ix2743 : nand03 port map ( Y=>nx2742, A0=>nx7809, A1=>nx7811, A2=>nx7813
   );
   ix7810 : aoi222 port map ( Y=>nx7809, A0=>que_out_19_3_7, A1=>nx10174, B0
      =>que_out_21_3_7, B1=>nx10148, C0=>que_out_8_3_7, C1=>nx10122);
   ix7812 : aoi22 port map ( Y=>nx7811, A0=>que_out_25_3_7, A1=>nx10070, B0
      =>que_out_16_3_7, B1=>nx10096);
   ix7814 : aoi22 port map ( Y=>nx7813, A0=>que_out_24_3_7, A1=>nx10044, B0
      =>que_out_22_3_7, B1=>nx10018);
   ix2715 : nand03 port map ( Y=>nx2714, A0=>nx7817, A1=>nx7819, A2=>nx7821
   );
   ix7818 : aoi222 port map ( Y=>nx7817, A0=>que_out_15_3_7, A1=>nx9966, B0
      =>que_out_3_3_7, B1=>nx9992, C0=>que_out_23_3_7, C1=>nx9940);
   ix7820 : aoi22 port map ( Y=>nx7819, A0=>que_out_27_3_7, A1=>nx9914, B0=>
      que_out_4_3_7, B1=>nx9888);
   ix7822 : aoi22 port map ( Y=>nx7821, A0=>que_out_0_3_7, A1=>nx9836, B0=>
      que_out_2_3_7, B1=>nx9862);
   ix2689 : nand03 port map ( Y=>nx2688, A0=>nx7825, A1=>nx7827, A2=>nx7829
   );
   ix7826 : aoi222 port map ( Y=>nx7825, A0=>que_out_26_3_7, A1=>nx9810, B0
      =>que_out_14_3_7, B1=>nx9784, C0=>que_out_11_3_7, C1=>nx9758);
   ix7828 : aoi22 port map ( Y=>nx7827, A0=>que_out_13_3_7, A1=>nx9732, B0=>
      que_out_7_3_7, B1=>nx9706);
   ix7830 : aoi22 port map ( Y=>nx7829, A0=>que_out_12_3_7, A1=>nx9680, B0=>
      que_out_1_3_7, B1=>nx9654);
   ix2883 : or04 port map ( Y=>out_column_3_8, A0=>nx2878, A1=>nx2852, A2=>
      nx2824, A3=>nx2798);
   ix2879 : nand03 port map ( Y=>nx2878, A0=>nx7835, A1=>nx7837, A2=>nx7839
   );
   ix7836 : aoi222 port map ( Y=>nx7835, A0=>que_out_10_3_8, A1=>nx10304, B0
      =>que_out_6_3_8, B1=>nx10356, C0=>que_out_9_3_8, C1=>nx10330);
   ix7838 : aoi22 port map ( Y=>nx7837, A0=>que_out_5_3_8, A1=>nx10252, B0=>
      que_out_18_3_8, B1=>nx10278);
   ix7840 : aoi22 port map ( Y=>nx7839, A0=>que_out_17_3_8, A1=>nx10226, B0
      =>que_out_20_3_8, B1=>nx10200);
   ix2853 : nand03 port map ( Y=>nx2852, A0=>nx7843, A1=>nx7845, A2=>nx7847
   );
   ix7844 : aoi222 port map ( Y=>nx7843, A0=>que_out_19_3_8, A1=>nx10174, B0
      =>que_out_21_3_8, B1=>nx10148, C0=>que_out_8_3_8, C1=>nx10122);
   ix7846 : aoi22 port map ( Y=>nx7845, A0=>que_out_25_3_8, A1=>nx10070, B0
      =>que_out_16_3_8, B1=>nx10096);
   ix7848 : aoi22 port map ( Y=>nx7847, A0=>que_out_24_3_8, A1=>nx10044, B0
      =>que_out_22_3_8, B1=>nx10018);
   ix2825 : nand03 port map ( Y=>nx2824, A0=>nx7851, A1=>nx7853, A2=>nx7855
   );
   ix7852 : aoi222 port map ( Y=>nx7851, A0=>que_out_15_3_8, A1=>nx9966, B0
      =>que_out_3_3_8, B1=>nx9992, C0=>que_out_23_3_8, C1=>nx9940);
   ix7854 : aoi22 port map ( Y=>nx7853, A0=>que_out_27_3_8, A1=>nx9914, B0=>
      que_out_4_3_8, B1=>nx9888);
   ix7856 : aoi22 port map ( Y=>nx7855, A0=>que_out_0_3_8, A1=>nx9836, B0=>
      que_out_2_3_8, B1=>nx9862);
   ix2799 : nand03 port map ( Y=>nx2798, A0=>nx7859, A1=>nx7861, A2=>nx7863
   );
   ix7860 : aoi222 port map ( Y=>nx7859, A0=>que_out_26_3_8, A1=>nx9810, B0
      =>que_out_14_3_8, B1=>nx9784, C0=>que_out_11_3_8, C1=>nx9758);
   ix7862 : aoi22 port map ( Y=>nx7861, A0=>que_out_13_3_8, A1=>nx9732, B0=>
      que_out_7_3_8, B1=>nx9706);
   ix7864 : aoi22 port map ( Y=>nx7863, A0=>que_out_12_3_8, A1=>nx9680, B0=>
      que_out_1_3_8, B1=>nx9654);
   ix2993 : or04 port map ( Y=>out_column_3_9, A0=>nx2988, A1=>nx2962, A2=>
      nx2934, A3=>nx2908);
   ix2989 : nand03 port map ( Y=>nx2988, A0=>nx7869, A1=>nx7871, A2=>nx7873
   );
   ix7870 : aoi222 port map ( Y=>nx7869, A0=>que_out_10_3_9, A1=>nx10304, B0
      =>que_out_6_3_9, B1=>nx10356, C0=>que_out_9_3_9, C1=>nx10330);
   ix7872 : aoi22 port map ( Y=>nx7871, A0=>que_out_5_3_9, A1=>nx10252, B0=>
      que_out_18_3_9, B1=>nx10278);
   ix7874 : aoi22 port map ( Y=>nx7873, A0=>que_out_17_3_9, A1=>nx10226, B0
      =>que_out_20_3_9, B1=>nx10200);
   ix2963 : nand03 port map ( Y=>nx2962, A0=>nx7877, A1=>nx7879, A2=>nx7881
   );
   ix7878 : aoi222 port map ( Y=>nx7877, A0=>que_out_19_3_9, A1=>nx10174, B0
      =>que_out_21_3_9, B1=>nx10148, C0=>que_out_8_3_9, C1=>nx10122);
   ix7880 : aoi22 port map ( Y=>nx7879, A0=>que_out_25_3_9, A1=>nx10070, B0
      =>que_out_16_3_9, B1=>nx10096);
   ix7882 : aoi22 port map ( Y=>nx7881, A0=>que_out_24_3_9, A1=>nx10044, B0
      =>que_out_22_3_9, B1=>nx10018);
   ix2935 : nand03 port map ( Y=>nx2934, A0=>nx7885, A1=>nx7887, A2=>nx7889
   );
   ix7886 : aoi222 port map ( Y=>nx7885, A0=>que_out_15_3_9, A1=>nx9966, B0
      =>que_out_3_3_9, B1=>nx9992, C0=>que_out_23_3_9, C1=>nx9940);
   ix7888 : aoi22 port map ( Y=>nx7887, A0=>que_out_27_3_9, A1=>nx9914, B0=>
      que_out_4_3_9, B1=>nx9888);
   ix7890 : aoi22 port map ( Y=>nx7889, A0=>que_out_0_3_9, A1=>nx9836, B0=>
      que_out_2_3_9, B1=>nx9862);
   ix2909 : nand03 port map ( Y=>nx2908, A0=>nx7893, A1=>nx7895, A2=>nx7897
   );
   ix7894 : aoi222 port map ( Y=>nx7893, A0=>que_out_26_3_9, A1=>nx9810, B0
      =>que_out_14_3_9, B1=>nx9784, C0=>que_out_11_3_9, C1=>nx9758);
   ix7896 : aoi22 port map ( Y=>nx7895, A0=>que_out_13_3_9, A1=>nx9732, B0=>
      que_out_7_3_9, B1=>nx9706);
   ix7898 : aoi22 port map ( Y=>nx7897, A0=>que_out_12_3_9, A1=>nx9680, B0=>
      que_out_1_3_9, B1=>nx9654);
   ix3103 : or04 port map ( Y=>out_column_3_10, A0=>nx3098, A1=>nx3072, A2=>
      nx3044, A3=>nx3018);
   ix3099 : nand03 port map ( Y=>nx3098, A0=>nx7903, A1=>nx7905, A2=>nx7907
   );
   ix7904 : aoi222 port map ( Y=>nx7903, A0=>que_out_10_3_10, A1=>nx10304, 
      B0=>que_out_6_3_10, B1=>nx10356, C0=>que_out_9_3_10, C1=>nx10330);
   ix7906 : aoi22 port map ( Y=>nx7905, A0=>que_out_5_3_10, A1=>nx10252, B0
      =>que_out_18_3_10, B1=>nx10278);
   ix7908 : aoi22 port map ( Y=>nx7907, A0=>que_out_17_3_10, A1=>nx10226, B0
      =>que_out_20_3_10, B1=>nx10200);
   ix3073 : nand03 port map ( Y=>nx3072, A0=>nx7911, A1=>nx7913, A2=>nx7915
   );
   ix7912 : aoi222 port map ( Y=>nx7911, A0=>que_out_19_3_10, A1=>nx10174, 
      B0=>que_out_21_3_10, B1=>nx10148, C0=>que_out_8_3_10, C1=>nx10122);
   ix7914 : aoi22 port map ( Y=>nx7913, A0=>que_out_25_3_10, A1=>nx10070, B0
      =>que_out_16_3_10, B1=>nx10096);
   ix7916 : aoi22 port map ( Y=>nx7915, A0=>que_out_24_3_10, A1=>nx10044, B0
      =>que_out_22_3_10, B1=>nx10018);
   ix3045 : nand03 port map ( Y=>nx3044, A0=>nx7919, A1=>nx7921, A2=>nx7923
   );
   ix7920 : aoi222 port map ( Y=>nx7919, A0=>que_out_15_3_10, A1=>nx9966, B0
      =>que_out_3_3_10, B1=>nx9992, C0=>que_out_23_3_10, C1=>nx9940);
   ix7922 : aoi22 port map ( Y=>nx7921, A0=>que_out_27_3_10, A1=>nx9914, B0
      =>que_out_4_3_10, B1=>nx9888);
   ix7924 : aoi22 port map ( Y=>nx7923, A0=>que_out_0_3_10, A1=>nx9836, B0=>
      que_out_2_3_10, B1=>nx9862);
   ix3019 : nand03 port map ( Y=>nx3018, A0=>nx7927, A1=>nx7929, A2=>nx7931
   );
   ix7928 : aoi222 port map ( Y=>nx7927, A0=>que_out_26_3_10, A1=>nx9810, B0
      =>que_out_14_3_10, B1=>nx9784, C0=>que_out_11_3_10, C1=>nx9758);
   ix7930 : aoi22 port map ( Y=>nx7929, A0=>que_out_13_3_10, A1=>nx9732, B0
      =>que_out_7_3_10, B1=>nx9706);
   ix7932 : aoi22 port map ( Y=>nx7931, A0=>que_out_12_3_10, A1=>nx9680, B0
      =>que_out_1_3_10, B1=>nx9654);
   ix3213 : or04 port map ( Y=>out_column_3_11, A0=>nx3208, A1=>nx3182, A2=>
      nx3154, A3=>nx3128);
   ix3209 : nand03 port map ( Y=>nx3208, A0=>nx7937, A1=>nx7939, A2=>nx7941
   );
   ix7938 : aoi222 port map ( Y=>nx7937, A0=>que_out_10_3_11, A1=>nx10304, 
      B0=>que_out_6_3_11, B1=>nx10356, C0=>que_out_9_3_11, C1=>nx10330);
   ix7940 : aoi22 port map ( Y=>nx7939, A0=>que_out_5_3_11, A1=>nx10252, B0
      =>que_out_18_3_11, B1=>nx10278);
   ix7942 : aoi22 port map ( Y=>nx7941, A0=>que_out_17_3_11, A1=>nx10226, B0
      =>que_out_20_3_11, B1=>nx10200);
   ix3183 : nand03 port map ( Y=>nx3182, A0=>nx7945, A1=>nx7947, A2=>nx7949
   );
   ix7946 : aoi222 port map ( Y=>nx7945, A0=>que_out_19_3_11, A1=>nx10174, 
      B0=>que_out_21_3_11, B1=>nx10148, C0=>que_out_8_3_11, C1=>nx10122);
   ix7948 : aoi22 port map ( Y=>nx7947, A0=>que_out_25_3_11, A1=>nx10070, B0
      =>que_out_16_3_11, B1=>nx10096);
   ix7950 : aoi22 port map ( Y=>nx7949, A0=>que_out_24_3_11, A1=>nx10044, B0
      =>que_out_22_3_11, B1=>nx10018);
   ix3155 : nand03 port map ( Y=>nx3154, A0=>nx7953, A1=>nx7955, A2=>nx7957
   );
   ix7954 : aoi222 port map ( Y=>nx7953, A0=>que_out_15_3_11, A1=>nx9966, B0
      =>que_out_3_3_11, B1=>nx9992, C0=>que_out_23_3_11, C1=>nx9940);
   ix7956 : aoi22 port map ( Y=>nx7955, A0=>que_out_27_3_11, A1=>nx9914, B0
      =>que_out_4_3_11, B1=>nx9888);
   ix7958 : aoi22 port map ( Y=>nx7957, A0=>que_out_0_3_11, A1=>nx9836, B0=>
      que_out_2_3_11, B1=>nx9862);
   ix3129 : nand03 port map ( Y=>nx3128, A0=>nx7961, A1=>nx7963, A2=>nx7965
   );
   ix7962 : aoi222 port map ( Y=>nx7961, A0=>que_out_26_3_11, A1=>nx9810, B0
      =>que_out_14_3_11, B1=>nx9784, C0=>que_out_11_3_11, C1=>nx9758);
   ix7964 : aoi22 port map ( Y=>nx7963, A0=>que_out_13_3_11, A1=>nx9732, B0
      =>que_out_7_3_11, B1=>nx9706);
   ix7966 : aoi22 port map ( Y=>nx7965, A0=>que_out_12_3_11, A1=>nx9680, B0
      =>que_out_1_3_11, B1=>nx9654);
   ix3323 : or04 port map ( Y=>out_column_3_12, A0=>nx3318, A1=>nx3292, A2=>
      nx3264, A3=>nx3238);
   ix3319 : nand03 port map ( Y=>nx3318, A0=>nx7971, A1=>nx7973, A2=>nx7975
   );
   ix7972 : aoi222 port map ( Y=>nx7971, A0=>que_out_10_3_12, A1=>nx10306, 
      B0=>que_out_6_3_12, B1=>nx10358, C0=>que_out_9_3_12, C1=>nx10332);
   ix7974 : aoi22 port map ( Y=>nx7973, A0=>que_out_5_3_12, A1=>nx10254, B0
      =>que_out_18_3_12, B1=>nx10280);
   ix7976 : aoi22 port map ( Y=>nx7975, A0=>que_out_17_3_12, A1=>nx10228, B0
      =>que_out_20_3_12, B1=>nx10202);
   ix3293 : nand03 port map ( Y=>nx3292, A0=>nx7979, A1=>nx7981, A2=>nx7983
   );
   ix7980 : aoi222 port map ( Y=>nx7979, A0=>que_out_19_3_12, A1=>nx10176, 
      B0=>que_out_21_3_12, B1=>nx10150, C0=>que_out_8_3_12, C1=>nx10124);
   ix7982 : aoi22 port map ( Y=>nx7981, A0=>que_out_25_3_12, A1=>nx10072, B0
      =>que_out_16_3_12, B1=>nx10098);
   ix7984 : aoi22 port map ( Y=>nx7983, A0=>que_out_24_3_12, A1=>nx10046, B0
      =>que_out_22_3_12, B1=>nx10020);
   ix3265 : nand03 port map ( Y=>nx3264, A0=>nx7987, A1=>nx7989, A2=>nx7991
   );
   ix7988 : aoi222 port map ( Y=>nx7987, A0=>que_out_15_3_12, A1=>nx9968, B0
      =>que_out_3_3_12, B1=>nx9994, C0=>que_out_23_3_12, C1=>nx9942);
   ix7990 : aoi22 port map ( Y=>nx7989, A0=>que_out_27_3_12, A1=>nx9916, B0
      =>que_out_4_3_12, B1=>nx9890);
   ix7992 : aoi22 port map ( Y=>nx7991, A0=>que_out_0_3_12, A1=>nx9838, B0=>
      que_out_2_3_12, B1=>nx9864);
   ix3239 : nand03 port map ( Y=>nx3238, A0=>nx7995, A1=>nx7997, A2=>nx7999
   );
   ix7996 : aoi222 port map ( Y=>nx7995, A0=>que_out_26_3_12, A1=>nx9812, B0
      =>que_out_14_3_12, B1=>nx9786, C0=>que_out_11_3_12, C1=>nx9760);
   ix7998 : aoi22 port map ( Y=>nx7997, A0=>que_out_13_3_12, A1=>nx9734, B0
      =>que_out_7_3_12, B1=>nx9708);
   ix8000 : aoi22 port map ( Y=>nx7999, A0=>que_out_12_3_12, A1=>nx9682, B0
      =>que_out_1_3_12, B1=>nx9656);
   ix3433 : or04 port map ( Y=>out_column_3_13, A0=>nx3428, A1=>nx3402, A2=>
      nx3374, A3=>nx3348);
   ix3429 : nand03 port map ( Y=>nx3428, A0=>nx8005, A1=>nx8007, A2=>nx8009
   );
   ix8006 : aoi222 port map ( Y=>nx8005, A0=>que_out_10_3_13, A1=>nx10306, 
      B0=>que_out_6_3_13, B1=>nx10358, C0=>que_out_9_3_13, C1=>nx10332);
   ix8008 : aoi22 port map ( Y=>nx8007, A0=>que_out_5_3_13, A1=>nx10254, B0
      =>que_out_18_3_13, B1=>nx10280);
   ix8010 : aoi22 port map ( Y=>nx8009, A0=>que_out_17_3_13, A1=>nx10228, B0
      =>que_out_20_3_13, B1=>nx10202);
   ix3403 : nand03 port map ( Y=>nx3402, A0=>nx8013, A1=>nx8015, A2=>nx8017
   );
   ix8014 : aoi222 port map ( Y=>nx8013, A0=>que_out_19_3_13, A1=>nx10176, 
      B0=>que_out_21_3_13, B1=>nx10150, C0=>que_out_8_3_13, C1=>nx10124);
   ix8016 : aoi22 port map ( Y=>nx8015, A0=>que_out_25_3_13, A1=>nx10072, B0
      =>que_out_16_3_13, B1=>nx10098);
   ix8018 : aoi22 port map ( Y=>nx8017, A0=>que_out_24_3_13, A1=>nx10046, B0
      =>que_out_22_3_13, B1=>nx10020);
   ix3375 : nand03 port map ( Y=>nx3374, A0=>nx8021, A1=>nx8023, A2=>nx8025
   );
   ix8022 : aoi222 port map ( Y=>nx8021, A0=>que_out_15_3_13, A1=>nx9968, B0
      =>que_out_3_3_13, B1=>nx9994, C0=>que_out_23_3_13, C1=>nx9942);
   ix8024 : aoi22 port map ( Y=>nx8023, A0=>que_out_27_3_13, A1=>nx9916, B0
      =>que_out_4_3_13, B1=>nx9890);
   ix8026 : aoi22 port map ( Y=>nx8025, A0=>que_out_0_3_13, A1=>nx9838, B0=>
      que_out_2_3_13, B1=>nx9864);
   ix3349 : nand03 port map ( Y=>nx3348, A0=>nx8029, A1=>nx8031, A2=>nx8033
   );
   ix8030 : aoi222 port map ( Y=>nx8029, A0=>que_out_26_3_13, A1=>nx9812, B0
      =>que_out_14_3_13, B1=>nx9786, C0=>que_out_11_3_13, C1=>nx9760);
   ix8032 : aoi22 port map ( Y=>nx8031, A0=>que_out_13_3_13, A1=>nx9734, B0
      =>que_out_7_3_13, B1=>nx9708);
   ix8034 : aoi22 port map ( Y=>nx8033, A0=>que_out_12_3_13, A1=>nx9682, B0
      =>que_out_1_3_13, B1=>nx9656);
   ix3543 : or04 port map ( Y=>out_column_3_14, A0=>nx3538, A1=>nx3512, A2=>
      nx3484, A3=>nx3458);
   ix3539 : nand03 port map ( Y=>nx3538, A0=>nx8039, A1=>nx8041, A2=>nx8043
   );
   ix8040 : aoi222 port map ( Y=>nx8039, A0=>que_out_10_3_14, A1=>nx10306, 
      B0=>que_out_6_3_14, B1=>nx10358, C0=>que_out_9_3_14, C1=>nx10332);
   ix8042 : aoi22 port map ( Y=>nx8041, A0=>que_out_5_3_14, A1=>nx10254, B0
      =>que_out_18_3_14, B1=>nx10280);
   ix8044 : aoi22 port map ( Y=>nx8043, A0=>que_out_17_3_14, A1=>nx10228, B0
      =>que_out_20_3_14, B1=>nx10202);
   ix3513 : nand03 port map ( Y=>nx3512, A0=>nx8047, A1=>nx8049, A2=>nx8051
   );
   ix8048 : aoi222 port map ( Y=>nx8047, A0=>que_out_19_3_14, A1=>nx10176, 
      B0=>que_out_21_3_14, B1=>nx10150, C0=>que_out_8_3_14, C1=>nx10124);
   ix8050 : aoi22 port map ( Y=>nx8049, A0=>que_out_25_3_14, A1=>nx10072, B0
      =>que_out_16_3_14, B1=>nx10098);
   ix8052 : aoi22 port map ( Y=>nx8051, A0=>que_out_24_3_14, A1=>nx10046, B0
      =>que_out_22_3_14, B1=>nx10020);
   ix3485 : nand03 port map ( Y=>nx3484, A0=>nx8055, A1=>nx8057, A2=>nx8059
   );
   ix8056 : aoi222 port map ( Y=>nx8055, A0=>que_out_15_3_14, A1=>nx9968, B0
      =>que_out_3_3_14, B1=>nx9994, C0=>que_out_23_3_14, C1=>nx9942);
   ix8058 : aoi22 port map ( Y=>nx8057, A0=>que_out_27_3_14, A1=>nx9916, B0
      =>que_out_4_3_14, B1=>nx9890);
   ix8060 : aoi22 port map ( Y=>nx8059, A0=>que_out_0_3_14, A1=>nx9838, B0=>
      que_out_2_3_14, B1=>nx9864);
   ix3459 : nand03 port map ( Y=>nx3458, A0=>nx8063, A1=>nx8065, A2=>nx8067
   );
   ix8064 : aoi222 port map ( Y=>nx8063, A0=>que_out_26_3_14, A1=>nx9812, B0
      =>que_out_14_3_14, B1=>nx9786, C0=>que_out_11_3_14, C1=>nx9760);
   ix8066 : aoi22 port map ( Y=>nx8065, A0=>que_out_13_3_14, A1=>nx9734, B0
      =>que_out_7_3_14, B1=>nx9708);
   ix8068 : aoi22 port map ( Y=>nx8067, A0=>que_out_12_3_14, A1=>nx9682, B0
      =>que_out_1_3_14, B1=>nx9656);
   ix3653 : or04 port map ( Y=>out_column_3_15, A0=>nx3648, A1=>nx3622, A2=>
      nx3594, A3=>nx3568);
   ix3649 : nand03 port map ( Y=>nx3648, A0=>nx8073, A1=>nx8075, A2=>nx8077
   );
   ix8074 : aoi222 port map ( Y=>nx8073, A0=>que_out_10_3_15, A1=>nx10306, 
      B0=>que_out_6_3_15, B1=>nx10358, C0=>que_out_9_3_15, C1=>nx10332);
   ix8076 : aoi22 port map ( Y=>nx8075, A0=>que_out_5_3_15, A1=>nx10254, B0
      =>que_out_18_3_15, B1=>nx10280);
   ix8078 : aoi22 port map ( Y=>nx8077, A0=>que_out_17_3_15, A1=>nx10228, B0
      =>que_out_20_3_15, B1=>nx10202);
   ix3623 : nand03 port map ( Y=>nx3622, A0=>nx8081, A1=>nx8083, A2=>nx8085
   );
   ix8082 : aoi222 port map ( Y=>nx8081, A0=>que_out_19_3_15, A1=>nx10176, 
      B0=>que_out_21_3_15, B1=>nx10150, C0=>que_out_8_3_15, C1=>nx10124);
   ix8084 : aoi22 port map ( Y=>nx8083, A0=>que_out_25_3_15, A1=>nx10072, B0
      =>que_out_16_3_15, B1=>nx10098);
   ix8086 : aoi22 port map ( Y=>nx8085, A0=>que_out_24_3_15, A1=>nx10046, B0
      =>que_out_22_3_15, B1=>nx10020);
   ix3595 : nand03 port map ( Y=>nx3594, A0=>nx8089, A1=>nx8091, A2=>nx8093
   );
   ix8090 : aoi222 port map ( Y=>nx8089, A0=>que_out_15_3_15, A1=>nx9968, B0
      =>que_out_3_3_15, B1=>nx9994, C0=>que_out_23_3_15, C1=>nx9942);
   ix8092 : aoi22 port map ( Y=>nx8091, A0=>que_out_27_3_15, A1=>nx9916, B0
      =>que_out_4_3_15, B1=>nx9890);
   ix8094 : aoi22 port map ( Y=>nx8093, A0=>que_out_0_3_15, A1=>nx9838, B0=>
      que_out_2_3_15, B1=>nx9864);
   ix3569 : nand03 port map ( Y=>nx3568, A0=>nx8097, A1=>nx8099, A2=>nx8101
   );
   ix8098 : aoi222 port map ( Y=>nx8097, A0=>que_out_26_3_15, A1=>nx9812, B0
      =>que_out_14_3_15, B1=>nx9786, C0=>que_out_11_3_15, C1=>nx9760);
   ix8100 : aoi22 port map ( Y=>nx8099, A0=>que_out_13_3_15, A1=>nx9734, B0
      =>que_out_7_3_15, B1=>nx9708);
   ix8102 : aoi22 port map ( Y=>nx8101, A0=>que_out_12_3_15, A1=>nx9682, B0
      =>que_out_1_3_15, B1=>nx9656);
   ix3763 : or04 port map ( Y=>out_column_2_0, A0=>nx3758, A1=>nx3732, A2=>
      nx3704, A3=>nx3678);
   ix3759 : nand03 port map ( Y=>nx3758, A0=>nx8107, A1=>nx8109, A2=>nx8111
   );
   ix8108 : aoi222 port map ( Y=>nx8107, A0=>que_out_10_2_0, A1=>nx10306, B0
      =>que_out_6_2_0, B1=>nx10358, C0=>que_out_9_2_0, C1=>nx10332);
   ix8110 : aoi22 port map ( Y=>nx8109, A0=>que_out_5_2_0, A1=>nx10254, B0=>
      que_out_18_2_0, B1=>nx10280);
   ix8112 : aoi22 port map ( Y=>nx8111, A0=>que_out_17_2_0, A1=>nx10228, B0
      =>que_out_20_2_0, B1=>nx10202);
   ix3733 : nand03 port map ( Y=>nx3732, A0=>nx8115, A1=>nx8117, A2=>nx8119
   );
   ix8116 : aoi222 port map ( Y=>nx8115, A0=>que_out_19_2_0, A1=>nx10176, B0
      =>que_out_21_2_0, B1=>nx10150, C0=>que_out_8_2_0, C1=>nx10124);
   ix8118 : aoi22 port map ( Y=>nx8117, A0=>que_out_25_2_0, A1=>nx10072, B0
      =>que_out_16_2_0, B1=>nx10098);
   ix8120 : aoi22 port map ( Y=>nx8119, A0=>que_out_24_2_0, A1=>nx10046, B0
      =>que_out_22_2_0, B1=>nx10020);
   ix3705 : nand03 port map ( Y=>nx3704, A0=>nx8123, A1=>nx8125, A2=>nx8127
   );
   ix8124 : aoi222 port map ( Y=>nx8123, A0=>que_out_15_2_0, A1=>nx9968, B0
      =>que_out_3_2_0, B1=>nx9994, C0=>que_out_23_2_0, C1=>nx9942);
   ix8126 : aoi22 port map ( Y=>nx8125, A0=>que_out_27_2_0, A1=>nx9916, B0=>
      que_out_4_2_0, B1=>nx9890);
   ix8128 : aoi22 port map ( Y=>nx8127, A0=>que_out_0_2_0, A1=>nx9838, B0=>
      que_out_2_2_0, B1=>nx9864);
   ix3679 : nand03 port map ( Y=>nx3678, A0=>nx8131, A1=>nx8133, A2=>nx8135
   );
   ix8132 : aoi222 port map ( Y=>nx8131, A0=>que_out_26_2_0, A1=>nx9812, B0
      =>que_out_14_2_0, B1=>nx9786, C0=>que_out_11_2_0, C1=>nx9760);
   ix8134 : aoi22 port map ( Y=>nx8133, A0=>que_out_13_2_0, A1=>nx9734, B0=>
      que_out_7_2_0, B1=>nx9708);
   ix8136 : aoi22 port map ( Y=>nx8135, A0=>que_out_12_2_0, A1=>nx9682, B0=>
      que_out_1_2_0, B1=>nx9656);
   ix3873 : or04 port map ( Y=>out_column_2_1, A0=>nx3868, A1=>nx3842, A2=>
      nx3814, A3=>nx3788);
   ix3869 : nand03 port map ( Y=>nx3868, A0=>nx8141, A1=>nx8143, A2=>nx8145
   );
   ix8142 : aoi222 port map ( Y=>nx8141, A0=>que_out_10_2_1, A1=>nx10306, B0
      =>que_out_6_2_1, B1=>nx10358, C0=>que_out_9_2_1, C1=>nx10332);
   ix8144 : aoi22 port map ( Y=>nx8143, A0=>que_out_5_2_1, A1=>nx10254, B0=>
      que_out_18_2_1, B1=>nx10280);
   ix8146 : aoi22 port map ( Y=>nx8145, A0=>que_out_17_2_1, A1=>nx10228, B0
      =>que_out_20_2_1, B1=>nx10202);
   ix3843 : nand03 port map ( Y=>nx3842, A0=>nx8149, A1=>nx8151, A2=>nx8153
   );
   ix8150 : aoi222 port map ( Y=>nx8149, A0=>que_out_19_2_1, A1=>nx10176, B0
      =>que_out_21_2_1, B1=>nx10150, C0=>que_out_8_2_1, C1=>nx10124);
   ix8152 : aoi22 port map ( Y=>nx8151, A0=>que_out_25_2_1, A1=>nx10072, B0
      =>que_out_16_2_1, B1=>nx10098);
   ix8154 : aoi22 port map ( Y=>nx8153, A0=>que_out_24_2_1, A1=>nx10046, B0
      =>que_out_22_2_1, B1=>nx10020);
   ix3815 : nand03 port map ( Y=>nx3814, A0=>nx8157, A1=>nx8159, A2=>nx8161
   );
   ix8158 : aoi222 port map ( Y=>nx8157, A0=>que_out_15_2_1, A1=>nx9968, B0
      =>que_out_3_2_1, B1=>nx9994, C0=>que_out_23_2_1, C1=>nx9942);
   ix8160 : aoi22 port map ( Y=>nx8159, A0=>que_out_27_2_1, A1=>nx9916, B0=>
      que_out_4_2_1, B1=>nx9890);
   ix8162 : aoi22 port map ( Y=>nx8161, A0=>que_out_0_2_1, A1=>nx9838, B0=>
      que_out_2_2_1, B1=>nx9864);
   ix3789 : nand03 port map ( Y=>nx3788, A0=>nx8165, A1=>nx8167, A2=>nx8169
   );
   ix8166 : aoi222 port map ( Y=>nx8165, A0=>que_out_26_2_1, A1=>nx9812, B0
      =>que_out_14_2_1, B1=>nx9786, C0=>que_out_11_2_1, C1=>nx9760);
   ix8168 : aoi22 port map ( Y=>nx8167, A0=>que_out_13_2_1, A1=>nx9734, B0=>
      que_out_7_2_1, B1=>nx9708);
   ix8170 : aoi22 port map ( Y=>nx8169, A0=>que_out_12_2_1, A1=>nx9682, B0=>
      que_out_1_2_1, B1=>nx9656);
   ix3983 : or04 port map ( Y=>out_column_2_2, A0=>nx3978, A1=>nx3952, A2=>
      nx3924, A3=>nx3898);
   ix3979 : nand03 port map ( Y=>nx3978, A0=>nx8175, A1=>nx8177, A2=>nx8179
   );
   ix8176 : aoi222 port map ( Y=>nx8175, A0=>que_out_10_2_2, A1=>nx10306, B0
      =>que_out_6_2_2, B1=>nx10358, C0=>que_out_9_2_2, C1=>nx10332);
   ix8178 : aoi22 port map ( Y=>nx8177, A0=>que_out_5_2_2, A1=>nx10254, B0=>
      que_out_18_2_2, B1=>nx10280);
   ix8180 : aoi22 port map ( Y=>nx8179, A0=>que_out_17_2_2, A1=>nx10228, B0
      =>que_out_20_2_2, B1=>nx10202);
   ix3953 : nand03 port map ( Y=>nx3952, A0=>nx8183, A1=>nx8185, A2=>nx8187
   );
   ix8184 : aoi222 port map ( Y=>nx8183, A0=>que_out_19_2_2, A1=>nx10176, B0
      =>que_out_21_2_2, B1=>nx10150, C0=>que_out_8_2_2, C1=>nx10124);
   ix8186 : aoi22 port map ( Y=>nx8185, A0=>que_out_25_2_2, A1=>nx10072, B0
      =>que_out_16_2_2, B1=>nx10098);
   ix8188 : aoi22 port map ( Y=>nx8187, A0=>que_out_24_2_2, A1=>nx10046, B0
      =>que_out_22_2_2, B1=>nx10020);
   ix3925 : nand03 port map ( Y=>nx3924, A0=>nx8191, A1=>nx8193, A2=>nx8195
   );
   ix8192 : aoi222 port map ( Y=>nx8191, A0=>que_out_15_2_2, A1=>nx9968, B0
      =>que_out_3_2_2, B1=>nx9994, C0=>que_out_23_2_2, C1=>nx9942);
   ix8194 : aoi22 port map ( Y=>nx8193, A0=>que_out_27_2_2, A1=>nx9916, B0=>
      que_out_4_2_2, B1=>nx9890);
   ix8196 : aoi22 port map ( Y=>nx8195, A0=>que_out_0_2_2, A1=>nx9838, B0=>
      que_out_2_2_2, B1=>nx9864);
   ix3899 : nand03 port map ( Y=>nx3898, A0=>nx8199, A1=>nx8201, A2=>nx8203
   );
   ix8200 : aoi222 port map ( Y=>nx8199, A0=>que_out_26_2_2, A1=>nx9812, B0
      =>que_out_14_2_2, B1=>nx9786, C0=>que_out_11_2_2, C1=>nx9760);
   ix8202 : aoi22 port map ( Y=>nx8201, A0=>que_out_13_2_2, A1=>nx9734, B0=>
      que_out_7_2_2, B1=>nx9708);
   ix8204 : aoi22 port map ( Y=>nx8203, A0=>que_out_12_2_2, A1=>nx9682, B0=>
      que_out_1_2_2, B1=>nx9656);
   ix4093 : or04 port map ( Y=>out_column_2_3, A0=>nx4088, A1=>nx4062, A2=>
      nx4034, A3=>nx4008);
   ix4089 : nand03 port map ( Y=>nx4088, A0=>nx8209, A1=>nx8211, A2=>nx8213
   );
   ix8210 : aoi222 port map ( Y=>nx8209, A0=>que_out_10_2_3, A1=>nx10308, B0
      =>que_out_6_2_3, B1=>nx10360, C0=>que_out_9_2_3, C1=>nx10334);
   ix8212 : aoi22 port map ( Y=>nx8211, A0=>que_out_5_2_3, A1=>nx10256, B0=>
      que_out_18_2_3, B1=>nx10282);
   ix8214 : aoi22 port map ( Y=>nx8213, A0=>que_out_17_2_3, A1=>nx10230, B0
      =>que_out_20_2_3, B1=>nx10204);
   ix4063 : nand03 port map ( Y=>nx4062, A0=>nx8217, A1=>nx8219, A2=>nx8221
   );
   ix8218 : aoi222 port map ( Y=>nx8217, A0=>que_out_19_2_3, A1=>nx10178, B0
      =>que_out_21_2_3, B1=>nx10152, C0=>que_out_8_2_3, C1=>nx10126);
   ix8220 : aoi22 port map ( Y=>nx8219, A0=>que_out_25_2_3, A1=>nx10074, B0
      =>que_out_16_2_3, B1=>nx10100);
   ix8222 : aoi22 port map ( Y=>nx8221, A0=>que_out_24_2_3, A1=>nx10048, B0
      =>que_out_22_2_3, B1=>nx10022);
   ix4035 : nand03 port map ( Y=>nx4034, A0=>nx8225, A1=>nx8227, A2=>nx8229
   );
   ix8226 : aoi222 port map ( Y=>nx8225, A0=>que_out_15_2_3, A1=>nx9970, B0
      =>que_out_3_2_3, B1=>nx9996, C0=>que_out_23_2_3, C1=>nx9944);
   ix8228 : aoi22 port map ( Y=>nx8227, A0=>que_out_27_2_3, A1=>nx9918, B0=>
      que_out_4_2_3, B1=>nx9892);
   ix8230 : aoi22 port map ( Y=>nx8229, A0=>que_out_0_2_3, A1=>nx9840, B0=>
      que_out_2_2_3, B1=>nx9866);
   ix4009 : nand03 port map ( Y=>nx4008, A0=>nx8233, A1=>nx8235, A2=>nx8237
   );
   ix8234 : aoi222 port map ( Y=>nx8233, A0=>que_out_26_2_3, A1=>nx9814, B0
      =>que_out_14_2_3, B1=>nx9788, C0=>que_out_11_2_3, C1=>nx9762);
   ix8236 : aoi22 port map ( Y=>nx8235, A0=>que_out_13_2_3, A1=>nx9736, B0=>
      que_out_7_2_3, B1=>nx9710);
   ix8238 : aoi22 port map ( Y=>nx8237, A0=>que_out_12_2_3, A1=>nx9684, B0=>
      que_out_1_2_3, B1=>nx9658);
   ix4203 : or04 port map ( Y=>out_column_2_4, A0=>nx4198, A1=>nx4172, A2=>
      nx4144, A3=>nx4118);
   ix4199 : nand03 port map ( Y=>nx4198, A0=>nx8243, A1=>nx8245, A2=>nx8247
   );
   ix8244 : aoi222 port map ( Y=>nx8243, A0=>que_out_10_2_4, A1=>nx10308, B0
      =>que_out_6_2_4, B1=>nx10360, C0=>que_out_9_2_4, C1=>nx10334);
   ix8246 : aoi22 port map ( Y=>nx8245, A0=>que_out_5_2_4, A1=>nx10256, B0=>
      que_out_18_2_4, B1=>nx10282);
   ix8248 : aoi22 port map ( Y=>nx8247, A0=>que_out_17_2_4, A1=>nx10230, B0
      =>que_out_20_2_4, B1=>nx10204);
   ix4173 : nand03 port map ( Y=>nx4172, A0=>nx8251, A1=>nx8253, A2=>nx8255
   );
   ix8252 : aoi222 port map ( Y=>nx8251, A0=>que_out_19_2_4, A1=>nx10178, B0
      =>que_out_21_2_4, B1=>nx10152, C0=>que_out_8_2_4, C1=>nx10126);
   ix8254 : aoi22 port map ( Y=>nx8253, A0=>que_out_25_2_4, A1=>nx10074, B0
      =>que_out_16_2_4, B1=>nx10100);
   ix8256 : aoi22 port map ( Y=>nx8255, A0=>que_out_24_2_4, A1=>nx10048, B0
      =>que_out_22_2_4, B1=>nx10022);
   ix4145 : nand03 port map ( Y=>nx4144, A0=>nx8259, A1=>nx8261, A2=>nx8263
   );
   ix8260 : aoi222 port map ( Y=>nx8259, A0=>que_out_15_2_4, A1=>nx9970, B0
      =>que_out_3_2_4, B1=>nx9996, C0=>que_out_23_2_4, C1=>nx9944);
   ix8262 : aoi22 port map ( Y=>nx8261, A0=>que_out_27_2_4, A1=>nx9918, B0=>
      que_out_4_2_4, B1=>nx9892);
   ix8264 : aoi22 port map ( Y=>nx8263, A0=>que_out_0_2_4, A1=>nx9840, B0=>
      que_out_2_2_4, B1=>nx9866);
   ix4119 : nand03 port map ( Y=>nx4118, A0=>nx8267, A1=>nx8269, A2=>nx8271
   );
   ix8268 : aoi222 port map ( Y=>nx8267, A0=>que_out_26_2_4, A1=>nx9814, B0
      =>que_out_14_2_4, B1=>nx9788, C0=>que_out_11_2_4, C1=>nx9762);
   ix8270 : aoi22 port map ( Y=>nx8269, A0=>que_out_13_2_4, A1=>nx9736, B0=>
      que_out_7_2_4, B1=>nx9710);
   ix8272 : aoi22 port map ( Y=>nx8271, A0=>que_out_12_2_4, A1=>nx9684, B0=>
      que_out_1_2_4, B1=>nx9658);
   ix4313 : or04 port map ( Y=>out_column_2_5, A0=>nx4308, A1=>nx4282, A2=>
      nx4254, A3=>nx4228);
   ix4309 : nand03 port map ( Y=>nx4308, A0=>nx8277, A1=>nx8279, A2=>nx8281
   );
   ix8278 : aoi222 port map ( Y=>nx8277, A0=>que_out_10_2_5, A1=>nx10308, B0
      =>que_out_6_2_5, B1=>nx10360, C0=>que_out_9_2_5, C1=>nx10334);
   ix8280 : aoi22 port map ( Y=>nx8279, A0=>que_out_5_2_5, A1=>nx10256, B0=>
      que_out_18_2_5, B1=>nx10282);
   ix8282 : aoi22 port map ( Y=>nx8281, A0=>que_out_17_2_5, A1=>nx10230, B0
      =>que_out_20_2_5, B1=>nx10204);
   ix4283 : nand03 port map ( Y=>nx4282, A0=>nx8285, A1=>nx8287, A2=>nx8289
   );
   ix8286 : aoi222 port map ( Y=>nx8285, A0=>que_out_19_2_5, A1=>nx10178, B0
      =>que_out_21_2_5, B1=>nx10152, C0=>que_out_8_2_5, C1=>nx10126);
   ix8288 : aoi22 port map ( Y=>nx8287, A0=>que_out_25_2_5, A1=>nx10074, B0
      =>que_out_16_2_5, B1=>nx10100);
   ix8290 : aoi22 port map ( Y=>nx8289, A0=>que_out_24_2_5, A1=>nx10048, B0
      =>que_out_22_2_5, B1=>nx10022);
   ix4255 : nand03 port map ( Y=>nx4254, A0=>nx8293, A1=>nx8295, A2=>nx8297
   );
   ix8294 : aoi222 port map ( Y=>nx8293, A0=>que_out_15_2_5, A1=>nx9970, B0
      =>que_out_3_2_5, B1=>nx9996, C0=>que_out_23_2_5, C1=>nx9944);
   ix8296 : aoi22 port map ( Y=>nx8295, A0=>que_out_27_2_5, A1=>nx9918, B0=>
      que_out_4_2_5, B1=>nx9892);
   ix8298 : aoi22 port map ( Y=>nx8297, A0=>que_out_0_2_5, A1=>nx9840, B0=>
      que_out_2_2_5, B1=>nx9866);
   ix4229 : nand03 port map ( Y=>nx4228, A0=>nx8301, A1=>nx8303, A2=>nx8305
   );
   ix8302 : aoi222 port map ( Y=>nx8301, A0=>que_out_26_2_5, A1=>nx9814, B0
      =>que_out_14_2_5, B1=>nx9788, C0=>que_out_11_2_5, C1=>nx9762);
   ix8304 : aoi22 port map ( Y=>nx8303, A0=>que_out_13_2_5, A1=>nx9736, B0=>
      que_out_7_2_5, B1=>nx9710);
   ix8306 : aoi22 port map ( Y=>nx8305, A0=>que_out_12_2_5, A1=>nx9684, B0=>
      que_out_1_2_5, B1=>nx9658);
   ix4423 : or04 port map ( Y=>out_column_2_6, A0=>nx4418, A1=>nx4392, A2=>
      nx4364, A3=>nx4338);
   ix4419 : nand03 port map ( Y=>nx4418, A0=>nx8311, A1=>nx8313, A2=>nx8315
   );
   ix8312 : aoi222 port map ( Y=>nx8311, A0=>que_out_10_2_6, A1=>nx10308, B0
      =>que_out_6_2_6, B1=>nx10360, C0=>que_out_9_2_6, C1=>nx10334);
   ix8314 : aoi22 port map ( Y=>nx8313, A0=>que_out_5_2_6, A1=>nx10256, B0=>
      que_out_18_2_6, B1=>nx10282);
   ix8316 : aoi22 port map ( Y=>nx8315, A0=>que_out_17_2_6, A1=>nx10230, B0
      =>que_out_20_2_6, B1=>nx10204);
   ix4393 : nand03 port map ( Y=>nx4392, A0=>nx8319, A1=>nx8321, A2=>nx8323
   );
   ix8320 : aoi222 port map ( Y=>nx8319, A0=>que_out_19_2_6, A1=>nx10178, B0
      =>que_out_21_2_6, B1=>nx10152, C0=>que_out_8_2_6, C1=>nx10126);
   ix8322 : aoi22 port map ( Y=>nx8321, A0=>que_out_25_2_6, A1=>nx10074, B0
      =>que_out_16_2_6, B1=>nx10100);
   ix8324 : aoi22 port map ( Y=>nx8323, A0=>que_out_24_2_6, A1=>nx10048, B0
      =>que_out_22_2_6, B1=>nx10022);
   ix4365 : nand03 port map ( Y=>nx4364, A0=>nx8327, A1=>nx8329, A2=>nx8331
   );
   ix8328 : aoi222 port map ( Y=>nx8327, A0=>que_out_15_2_6, A1=>nx9970, B0
      =>que_out_3_2_6, B1=>nx9996, C0=>que_out_23_2_6, C1=>nx9944);
   ix8330 : aoi22 port map ( Y=>nx8329, A0=>que_out_27_2_6, A1=>nx9918, B0=>
      que_out_4_2_6, B1=>nx9892);
   ix8332 : aoi22 port map ( Y=>nx8331, A0=>que_out_0_2_6, A1=>nx9840, B0=>
      que_out_2_2_6, B1=>nx9866);
   ix4339 : nand03 port map ( Y=>nx4338, A0=>nx8335, A1=>nx8337, A2=>nx8339
   );
   ix8336 : aoi222 port map ( Y=>nx8335, A0=>que_out_26_2_6, A1=>nx9814, B0
      =>que_out_14_2_6, B1=>nx9788, C0=>que_out_11_2_6, C1=>nx9762);
   ix8338 : aoi22 port map ( Y=>nx8337, A0=>que_out_13_2_6, A1=>nx9736, B0=>
      que_out_7_2_6, B1=>nx9710);
   ix8340 : aoi22 port map ( Y=>nx8339, A0=>que_out_12_2_6, A1=>nx9684, B0=>
      que_out_1_2_6, B1=>nx9658);
   ix4533 : or04 port map ( Y=>out_column_2_7, A0=>nx4528, A1=>nx4502, A2=>
      nx4474, A3=>nx4448);
   ix4529 : nand03 port map ( Y=>nx4528, A0=>nx8345, A1=>nx8347, A2=>nx8349
   );
   ix8346 : aoi222 port map ( Y=>nx8345, A0=>que_out_10_2_7, A1=>nx10308, B0
      =>que_out_6_2_7, B1=>nx10360, C0=>que_out_9_2_7, C1=>nx10334);
   ix8348 : aoi22 port map ( Y=>nx8347, A0=>que_out_5_2_7, A1=>nx10256, B0=>
      que_out_18_2_7, B1=>nx10282);
   ix8350 : aoi22 port map ( Y=>nx8349, A0=>que_out_17_2_7, A1=>nx10230, B0
      =>que_out_20_2_7, B1=>nx10204);
   ix4503 : nand03 port map ( Y=>nx4502, A0=>nx8353, A1=>nx8355, A2=>nx8357
   );
   ix8354 : aoi222 port map ( Y=>nx8353, A0=>que_out_19_2_7, A1=>nx10178, B0
      =>que_out_21_2_7, B1=>nx10152, C0=>que_out_8_2_7, C1=>nx10126);
   ix8356 : aoi22 port map ( Y=>nx8355, A0=>que_out_25_2_7, A1=>nx10074, B0
      =>que_out_16_2_7, B1=>nx10100);
   ix8358 : aoi22 port map ( Y=>nx8357, A0=>que_out_24_2_7, A1=>nx10048, B0
      =>que_out_22_2_7, B1=>nx10022);
   ix4475 : nand03 port map ( Y=>nx4474, A0=>nx8361, A1=>nx8363, A2=>nx8365
   );
   ix8362 : aoi222 port map ( Y=>nx8361, A0=>que_out_15_2_7, A1=>nx9970, B0
      =>que_out_3_2_7, B1=>nx9996, C0=>que_out_23_2_7, C1=>nx9944);
   ix8364 : aoi22 port map ( Y=>nx8363, A0=>que_out_27_2_7, A1=>nx9918, B0=>
      que_out_4_2_7, B1=>nx9892);
   ix8366 : aoi22 port map ( Y=>nx8365, A0=>que_out_0_2_7, A1=>nx9840, B0=>
      que_out_2_2_7, B1=>nx9866);
   ix4449 : nand03 port map ( Y=>nx4448, A0=>nx8369, A1=>nx8371, A2=>nx8373
   );
   ix8370 : aoi222 port map ( Y=>nx8369, A0=>que_out_26_2_7, A1=>nx9814, B0
      =>que_out_14_2_7, B1=>nx9788, C0=>que_out_11_2_7, C1=>nx9762);
   ix8372 : aoi22 port map ( Y=>nx8371, A0=>que_out_13_2_7, A1=>nx9736, B0=>
      que_out_7_2_7, B1=>nx9710);
   ix8374 : aoi22 port map ( Y=>nx8373, A0=>que_out_12_2_7, A1=>nx9684, B0=>
      que_out_1_2_7, B1=>nx9658);
   ix4643 : or04 port map ( Y=>out_column_2_8, A0=>nx4638, A1=>nx4612, A2=>
      nx4584, A3=>nx4558);
   ix4639 : nand03 port map ( Y=>nx4638, A0=>nx8379, A1=>nx8381, A2=>nx8383
   );
   ix8380 : aoi222 port map ( Y=>nx8379, A0=>que_out_10_2_8, A1=>nx10308, B0
      =>que_out_6_2_8, B1=>nx10360, C0=>que_out_9_2_8, C1=>nx10334);
   ix8382 : aoi22 port map ( Y=>nx8381, A0=>que_out_5_2_8, A1=>nx10256, B0=>
      que_out_18_2_8, B1=>nx10282);
   ix8384 : aoi22 port map ( Y=>nx8383, A0=>que_out_17_2_8, A1=>nx10230, B0
      =>que_out_20_2_8, B1=>nx10204);
   ix4613 : nand03 port map ( Y=>nx4612, A0=>nx8387, A1=>nx8389, A2=>nx8391
   );
   ix8388 : aoi222 port map ( Y=>nx8387, A0=>que_out_19_2_8, A1=>nx10178, B0
      =>que_out_21_2_8, B1=>nx10152, C0=>que_out_8_2_8, C1=>nx10126);
   ix8390 : aoi22 port map ( Y=>nx8389, A0=>que_out_25_2_8, A1=>nx10074, B0
      =>que_out_16_2_8, B1=>nx10100);
   ix8392 : aoi22 port map ( Y=>nx8391, A0=>que_out_24_2_8, A1=>nx10048, B0
      =>que_out_22_2_8, B1=>nx10022);
   ix4585 : nand03 port map ( Y=>nx4584, A0=>nx8395, A1=>nx8397, A2=>nx8399
   );
   ix8396 : aoi222 port map ( Y=>nx8395, A0=>que_out_15_2_8, A1=>nx9970, B0
      =>que_out_3_2_8, B1=>nx9996, C0=>que_out_23_2_8, C1=>nx9944);
   ix8398 : aoi22 port map ( Y=>nx8397, A0=>que_out_27_2_8, A1=>nx9918, B0=>
      que_out_4_2_8, B1=>nx9892);
   ix8400 : aoi22 port map ( Y=>nx8399, A0=>que_out_0_2_8, A1=>nx9840, B0=>
      que_out_2_2_8, B1=>nx9866);
   ix4559 : nand03 port map ( Y=>nx4558, A0=>nx8403, A1=>nx8405, A2=>nx8407
   );
   ix8404 : aoi222 port map ( Y=>nx8403, A0=>que_out_26_2_8, A1=>nx9814, B0
      =>que_out_14_2_8, B1=>nx9788, C0=>que_out_11_2_8, C1=>nx9762);
   ix8406 : aoi22 port map ( Y=>nx8405, A0=>que_out_13_2_8, A1=>nx9736, B0=>
      que_out_7_2_8, B1=>nx9710);
   ix8408 : aoi22 port map ( Y=>nx8407, A0=>que_out_12_2_8, A1=>nx9684, B0=>
      que_out_1_2_8, B1=>nx9658);
   ix4753 : or04 port map ( Y=>out_column_2_9, A0=>nx4748, A1=>nx4722, A2=>
      nx4694, A3=>nx4668);
   ix4749 : nand03 port map ( Y=>nx4748, A0=>nx8413, A1=>nx8415, A2=>nx8417
   );
   ix8414 : aoi222 port map ( Y=>nx8413, A0=>que_out_10_2_9, A1=>nx10308, B0
      =>que_out_6_2_9, B1=>nx10360, C0=>que_out_9_2_9, C1=>nx10334);
   ix8416 : aoi22 port map ( Y=>nx8415, A0=>que_out_5_2_9, A1=>nx10256, B0=>
      que_out_18_2_9, B1=>nx10282);
   ix8418 : aoi22 port map ( Y=>nx8417, A0=>que_out_17_2_9, A1=>nx10230, B0
      =>que_out_20_2_9, B1=>nx10204);
   ix4723 : nand03 port map ( Y=>nx4722, A0=>nx8421, A1=>nx8423, A2=>nx8425
   );
   ix8422 : aoi222 port map ( Y=>nx8421, A0=>que_out_19_2_9, A1=>nx10178, B0
      =>que_out_21_2_9, B1=>nx10152, C0=>que_out_8_2_9, C1=>nx10126);
   ix8424 : aoi22 port map ( Y=>nx8423, A0=>que_out_25_2_9, A1=>nx10074, B0
      =>que_out_16_2_9, B1=>nx10100);
   ix8426 : aoi22 port map ( Y=>nx8425, A0=>que_out_24_2_9, A1=>nx10048, B0
      =>que_out_22_2_9, B1=>nx10022);
   ix4695 : nand03 port map ( Y=>nx4694, A0=>nx8429, A1=>nx8431, A2=>nx8433
   );
   ix8430 : aoi222 port map ( Y=>nx8429, A0=>que_out_15_2_9, A1=>nx9970, B0
      =>que_out_3_2_9, B1=>nx9996, C0=>que_out_23_2_9, C1=>nx9944);
   ix8432 : aoi22 port map ( Y=>nx8431, A0=>que_out_27_2_9, A1=>nx9918, B0=>
      que_out_4_2_9, B1=>nx9892);
   ix8434 : aoi22 port map ( Y=>nx8433, A0=>que_out_0_2_9, A1=>nx9840, B0=>
      que_out_2_2_9, B1=>nx9866);
   ix4669 : nand03 port map ( Y=>nx4668, A0=>nx8437, A1=>nx8439, A2=>nx8441
   );
   ix8438 : aoi222 port map ( Y=>nx8437, A0=>que_out_26_2_9, A1=>nx9814, B0
      =>que_out_14_2_9, B1=>nx9788, C0=>que_out_11_2_9, C1=>nx9762);
   ix8440 : aoi22 port map ( Y=>nx8439, A0=>que_out_13_2_9, A1=>nx9736, B0=>
      que_out_7_2_9, B1=>nx9710);
   ix8442 : aoi22 port map ( Y=>nx8441, A0=>que_out_12_2_9, A1=>nx9684, B0=>
      que_out_1_2_9, B1=>nx9658);
   ix4863 : or04 port map ( Y=>out_column_2_10, A0=>nx4858, A1=>nx4832, A2=>
      nx4804, A3=>nx4778);
   ix4859 : nand03 port map ( Y=>nx4858, A0=>nx8447, A1=>nx8449, A2=>nx8451
   );
   ix8448 : aoi222 port map ( Y=>nx8447, A0=>que_out_10_2_10, A1=>nx10310, 
      B0=>que_out_6_2_10, B1=>nx10362, C0=>que_out_9_2_10, C1=>nx10336);
   ix8450 : aoi22 port map ( Y=>nx8449, A0=>que_out_5_2_10, A1=>nx10258, B0
      =>que_out_18_2_10, B1=>nx10284);
   ix8452 : aoi22 port map ( Y=>nx8451, A0=>que_out_17_2_10, A1=>nx10232, B0
      =>que_out_20_2_10, B1=>nx10206);
   ix4833 : nand03 port map ( Y=>nx4832, A0=>nx8455, A1=>nx8457, A2=>nx8459
   );
   ix8456 : aoi222 port map ( Y=>nx8455, A0=>que_out_19_2_10, A1=>nx10180, 
      B0=>que_out_21_2_10, B1=>nx10154, C0=>que_out_8_2_10, C1=>nx10128);
   ix8458 : aoi22 port map ( Y=>nx8457, A0=>que_out_25_2_10, A1=>nx10076, B0
      =>que_out_16_2_10, B1=>nx10102);
   ix8460 : aoi22 port map ( Y=>nx8459, A0=>que_out_24_2_10, A1=>nx10050, B0
      =>que_out_22_2_10, B1=>nx10024);
   ix4805 : nand03 port map ( Y=>nx4804, A0=>nx8463, A1=>nx8465, A2=>nx8467
   );
   ix8464 : aoi222 port map ( Y=>nx8463, A0=>que_out_15_2_10, A1=>nx9972, B0
      =>que_out_3_2_10, B1=>nx9998, C0=>que_out_23_2_10, C1=>nx9946);
   ix8466 : aoi22 port map ( Y=>nx8465, A0=>que_out_27_2_10, A1=>nx9920, B0
      =>que_out_4_2_10, B1=>nx9894);
   ix8468 : aoi22 port map ( Y=>nx8467, A0=>que_out_0_2_10, A1=>nx9842, B0=>
      que_out_2_2_10, B1=>nx9868);
   ix4779 : nand03 port map ( Y=>nx4778, A0=>nx8471, A1=>nx8473, A2=>nx8475
   );
   ix8472 : aoi222 port map ( Y=>nx8471, A0=>que_out_26_2_10, A1=>nx9816, B0
      =>que_out_14_2_10, B1=>nx9790, C0=>que_out_11_2_10, C1=>nx9764);
   ix8474 : aoi22 port map ( Y=>nx8473, A0=>que_out_13_2_10, A1=>nx9738, B0
      =>que_out_7_2_10, B1=>nx9712);
   ix8476 : aoi22 port map ( Y=>nx8475, A0=>que_out_12_2_10, A1=>nx9686, B0
      =>que_out_1_2_10, B1=>nx9660);
   ix4973 : or04 port map ( Y=>out_column_2_11, A0=>nx4968, A1=>nx4942, A2=>
      nx4914, A3=>nx4888);
   ix4969 : nand03 port map ( Y=>nx4968, A0=>nx8481, A1=>nx8483, A2=>nx8485
   );
   ix8482 : aoi222 port map ( Y=>nx8481, A0=>que_out_10_2_11, A1=>nx10310, 
      B0=>que_out_6_2_11, B1=>nx10362, C0=>que_out_9_2_11, C1=>nx10336);
   ix8484 : aoi22 port map ( Y=>nx8483, A0=>que_out_5_2_11, A1=>nx10258, B0
      =>que_out_18_2_11, B1=>nx10284);
   ix8486 : aoi22 port map ( Y=>nx8485, A0=>que_out_17_2_11, A1=>nx10232, B0
      =>que_out_20_2_11, B1=>nx10206);
   ix4943 : nand03 port map ( Y=>nx4942, A0=>nx8489, A1=>nx8491, A2=>nx8493
   );
   ix8490 : aoi222 port map ( Y=>nx8489, A0=>que_out_19_2_11, A1=>nx10180, 
      B0=>que_out_21_2_11, B1=>nx10154, C0=>que_out_8_2_11, C1=>nx10128);
   ix8492 : aoi22 port map ( Y=>nx8491, A0=>que_out_25_2_11, A1=>nx10076, B0
      =>que_out_16_2_11, B1=>nx10102);
   ix8494 : aoi22 port map ( Y=>nx8493, A0=>que_out_24_2_11, A1=>nx10050, B0
      =>que_out_22_2_11, B1=>nx10024);
   ix4915 : nand03 port map ( Y=>nx4914, A0=>nx8497, A1=>nx8499, A2=>nx8501
   );
   ix8498 : aoi222 port map ( Y=>nx8497, A0=>que_out_15_2_11, A1=>nx9972, B0
      =>que_out_3_2_11, B1=>nx9998, C0=>que_out_23_2_11, C1=>nx9946);
   ix8500 : aoi22 port map ( Y=>nx8499, A0=>que_out_27_2_11, A1=>nx9920, B0
      =>que_out_4_2_11, B1=>nx9894);
   ix8502 : aoi22 port map ( Y=>nx8501, A0=>que_out_0_2_11, A1=>nx9842, B0=>
      que_out_2_2_11, B1=>nx9868);
   ix4889 : nand03 port map ( Y=>nx4888, A0=>nx8505, A1=>nx8507, A2=>nx8509
   );
   ix8506 : aoi222 port map ( Y=>nx8505, A0=>que_out_26_2_11, A1=>nx9816, B0
      =>que_out_14_2_11, B1=>nx9790, C0=>que_out_11_2_11, C1=>nx9764);
   ix8508 : aoi22 port map ( Y=>nx8507, A0=>que_out_13_2_11, A1=>nx9738, B0
      =>que_out_7_2_11, B1=>nx9712);
   ix8510 : aoi22 port map ( Y=>nx8509, A0=>que_out_12_2_11, A1=>nx9686, B0
      =>que_out_1_2_11, B1=>nx9660);
   ix5083 : or04 port map ( Y=>out_column_2_12, A0=>nx5078, A1=>nx5052, A2=>
      nx5024, A3=>nx4998);
   ix5079 : nand03 port map ( Y=>nx5078, A0=>nx8515, A1=>nx8517, A2=>nx8519
   );
   ix8516 : aoi222 port map ( Y=>nx8515, A0=>que_out_10_2_12, A1=>nx10310, 
      B0=>que_out_6_2_12, B1=>nx10362, C0=>que_out_9_2_12, C1=>nx10336);
   ix8518 : aoi22 port map ( Y=>nx8517, A0=>que_out_5_2_12, A1=>nx10258, B0
      =>que_out_18_2_12, B1=>nx10284);
   ix8520 : aoi22 port map ( Y=>nx8519, A0=>que_out_17_2_12, A1=>nx10232, B0
      =>que_out_20_2_12, B1=>nx10206);
   ix5053 : nand03 port map ( Y=>nx5052, A0=>nx8523, A1=>nx8525, A2=>nx8527
   );
   ix8524 : aoi222 port map ( Y=>nx8523, A0=>que_out_19_2_12, A1=>nx10180, 
      B0=>que_out_21_2_12, B1=>nx10154, C0=>que_out_8_2_12, C1=>nx10128);
   ix8526 : aoi22 port map ( Y=>nx8525, A0=>que_out_25_2_12, A1=>nx10076, B0
      =>que_out_16_2_12, B1=>nx10102);
   ix8528 : aoi22 port map ( Y=>nx8527, A0=>que_out_24_2_12, A1=>nx10050, B0
      =>que_out_22_2_12, B1=>nx10024);
   ix5025 : nand03 port map ( Y=>nx5024, A0=>nx8531, A1=>nx8533, A2=>nx8535
   );
   ix8532 : aoi222 port map ( Y=>nx8531, A0=>que_out_15_2_12, A1=>nx9972, B0
      =>que_out_3_2_12, B1=>nx9998, C0=>que_out_23_2_12, C1=>nx9946);
   ix8534 : aoi22 port map ( Y=>nx8533, A0=>que_out_27_2_12, A1=>nx9920, B0
      =>que_out_4_2_12, B1=>nx9894);
   ix8536 : aoi22 port map ( Y=>nx8535, A0=>que_out_0_2_12, A1=>nx9842, B0=>
      que_out_2_2_12, B1=>nx9868);
   ix4999 : nand03 port map ( Y=>nx4998, A0=>nx8539, A1=>nx8541, A2=>nx8543
   );
   ix8540 : aoi222 port map ( Y=>nx8539, A0=>que_out_26_2_12, A1=>nx9816, B0
      =>que_out_14_2_12, B1=>nx9790, C0=>que_out_11_2_12, C1=>nx9764);
   ix8542 : aoi22 port map ( Y=>nx8541, A0=>que_out_13_2_12, A1=>nx9738, B0
      =>que_out_7_2_12, B1=>nx9712);
   ix8544 : aoi22 port map ( Y=>nx8543, A0=>que_out_12_2_12, A1=>nx9686, B0
      =>que_out_1_2_12, B1=>nx9660);
   ix5193 : or04 port map ( Y=>out_column_2_13, A0=>nx5188, A1=>nx5162, A2=>
      nx5134, A3=>nx5108);
   ix5189 : nand03 port map ( Y=>nx5188, A0=>nx8549, A1=>nx8551, A2=>nx8553
   );
   ix8550 : aoi222 port map ( Y=>nx8549, A0=>que_out_10_2_13, A1=>nx10310, 
      B0=>que_out_6_2_13, B1=>nx10362, C0=>que_out_9_2_13, C1=>nx10336);
   ix8552 : aoi22 port map ( Y=>nx8551, A0=>que_out_5_2_13, A1=>nx10258, B0
      =>que_out_18_2_13, B1=>nx10284);
   ix8554 : aoi22 port map ( Y=>nx8553, A0=>que_out_17_2_13, A1=>nx10232, B0
      =>que_out_20_2_13, B1=>nx10206);
   ix5163 : nand03 port map ( Y=>nx5162, A0=>nx8557, A1=>nx8559, A2=>nx8561
   );
   ix8558 : aoi222 port map ( Y=>nx8557, A0=>que_out_19_2_13, A1=>nx10180, 
      B0=>que_out_21_2_13, B1=>nx10154, C0=>que_out_8_2_13, C1=>nx10128);
   ix8560 : aoi22 port map ( Y=>nx8559, A0=>que_out_25_2_13, A1=>nx10076, B0
      =>que_out_16_2_13, B1=>nx10102);
   ix8562 : aoi22 port map ( Y=>nx8561, A0=>que_out_24_2_13, A1=>nx10050, B0
      =>que_out_22_2_13, B1=>nx10024);
   ix5135 : nand03 port map ( Y=>nx5134, A0=>nx8565, A1=>nx8567, A2=>nx8569
   );
   ix8566 : aoi222 port map ( Y=>nx8565, A0=>que_out_15_2_13, A1=>nx9972, B0
      =>que_out_3_2_13, B1=>nx9998, C0=>que_out_23_2_13, C1=>nx9946);
   ix8568 : aoi22 port map ( Y=>nx8567, A0=>que_out_27_2_13, A1=>nx9920, B0
      =>que_out_4_2_13, B1=>nx9894);
   ix8570 : aoi22 port map ( Y=>nx8569, A0=>que_out_0_2_13, A1=>nx9842, B0=>
      que_out_2_2_13, B1=>nx9868);
   ix5109 : nand03 port map ( Y=>nx5108, A0=>nx8573, A1=>nx8575, A2=>nx8577
   );
   ix8574 : aoi222 port map ( Y=>nx8573, A0=>que_out_26_2_13, A1=>nx9816, B0
      =>que_out_14_2_13, B1=>nx9790, C0=>que_out_11_2_13, C1=>nx9764);
   ix8576 : aoi22 port map ( Y=>nx8575, A0=>que_out_13_2_13, A1=>nx9738, B0
      =>que_out_7_2_13, B1=>nx9712);
   ix8578 : aoi22 port map ( Y=>nx8577, A0=>que_out_12_2_13, A1=>nx9686, B0
      =>que_out_1_2_13, B1=>nx9660);
   ix5303 : or04 port map ( Y=>out_column_2_14, A0=>nx5298, A1=>nx5272, A2=>
      nx5244, A3=>nx5218);
   ix5299 : nand03 port map ( Y=>nx5298, A0=>nx8583, A1=>nx8585, A2=>nx8587
   );
   ix8584 : aoi222 port map ( Y=>nx8583, A0=>que_out_10_2_14, A1=>nx10310, 
      B0=>que_out_6_2_14, B1=>nx10362, C0=>que_out_9_2_14, C1=>nx10336);
   ix8586 : aoi22 port map ( Y=>nx8585, A0=>que_out_5_2_14, A1=>nx10258, B0
      =>que_out_18_2_14, B1=>nx10284);
   ix8588 : aoi22 port map ( Y=>nx8587, A0=>que_out_17_2_14, A1=>nx10232, B0
      =>que_out_20_2_14, B1=>nx10206);
   ix5273 : nand03 port map ( Y=>nx5272, A0=>nx8591, A1=>nx8593, A2=>nx8595
   );
   ix8592 : aoi222 port map ( Y=>nx8591, A0=>que_out_19_2_14, A1=>nx10180, 
      B0=>que_out_21_2_14, B1=>nx10154, C0=>que_out_8_2_14, C1=>nx10128);
   ix8594 : aoi22 port map ( Y=>nx8593, A0=>que_out_25_2_14, A1=>nx10076, B0
      =>que_out_16_2_14, B1=>nx10102);
   ix8596 : aoi22 port map ( Y=>nx8595, A0=>que_out_24_2_14, A1=>nx10050, B0
      =>que_out_22_2_14, B1=>nx10024);
   ix5245 : nand03 port map ( Y=>nx5244, A0=>nx8599, A1=>nx8601, A2=>nx8603
   );
   ix8600 : aoi222 port map ( Y=>nx8599, A0=>que_out_15_2_14, A1=>nx9972, B0
      =>que_out_3_2_14, B1=>nx9998, C0=>que_out_23_2_14, C1=>nx9946);
   ix8602 : aoi22 port map ( Y=>nx8601, A0=>que_out_27_2_14, A1=>nx9920, B0
      =>que_out_4_2_14, B1=>nx9894);
   ix8604 : aoi22 port map ( Y=>nx8603, A0=>que_out_0_2_14, A1=>nx9842, B0=>
      que_out_2_2_14, B1=>nx9868);
   ix5219 : nand03 port map ( Y=>nx5218, A0=>nx8607, A1=>nx8609, A2=>nx8611
   );
   ix8608 : aoi222 port map ( Y=>nx8607, A0=>que_out_26_2_14, A1=>nx9816, B0
      =>que_out_14_2_14, B1=>nx9790, C0=>que_out_11_2_14, C1=>nx9764);
   ix8610 : aoi22 port map ( Y=>nx8609, A0=>que_out_13_2_14, A1=>nx9738, B0
      =>que_out_7_2_14, B1=>nx9712);
   ix8612 : aoi22 port map ( Y=>nx8611, A0=>que_out_12_2_14, A1=>nx9686, B0
      =>que_out_1_2_14, B1=>nx9660);
   ix5413 : or04 port map ( Y=>out_column_2_15, A0=>nx5408, A1=>nx5382, A2=>
      nx5354, A3=>nx5328);
   ix5409 : nand03 port map ( Y=>nx5408, A0=>nx8617, A1=>nx8619, A2=>nx8621
   );
   ix8618 : aoi222 port map ( Y=>nx8617, A0=>que_out_10_2_15, A1=>nx10310, 
      B0=>que_out_6_2_15, B1=>nx10362, C0=>que_out_9_2_15, C1=>nx10336);
   ix8620 : aoi22 port map ( Y=>nx8619, A0=>que_out_5_2_15, A1=>nx10258, B0
      =>que_out_18_2_15, B1=>nx10284);
   ix8622 : aoi22 port map ( Y=>nx8621, A0=>que_out_17_2_15, A1=>nx10232, B0
      =>que_out_20_2_15, B1=>nx10206);
   ix5383 : nand03 port map ( Y=>nx5382, A0=>nx8625, A1=>nx8627, A2=>nx8629
   );
   ix8626 : aoi222 port map ( Y=>nx8625, A0=>que_out_19_2_15, A1=>nx10180, 
      B0=>que_out_21_2_15, B1=>nx10154, C0=>que_out_8_2_15, C1=>nx10128);
   ix8628 : aoi22 port map ( Y=>nx8627, A0=>que_out_25_2_15, A1=>nx10076, B0
      =>que_out_16_2_15, B1=>nx10102);
   ix8630 : aoi22 port map ( Y=>nx8629, A0=>que_out_24_2_15, A1=>nx10050, B0
      =>que_out_22_2_15, B1=>nx10024);
   ix5355 : nand03 port map ( Y=>nx5354, A0=>nx8633, A1=>nx8635, A2=>nx8637
   );
   ix8634 : aoi222 port map ( Y=>nx8633, A0=>que_out_15_2_15, A1=>nx9972, B0
      =>que_out_3_2_15, B1=>nx9998, C0=>que_out_23_2_15, C1=>nx9946);
   ix8636 : aoi22 port map ( Y=>nx8635, A0=>que_out_27_2_15, A1=>nx9920, B0
      =>que_out_4_2_15, B1=>nx9894);
   ix8638 : aoi22 port map ( Y=>nx8637, A0=>que_out_0_2_15, A1=>nx9842, B0=>
      que_out_2_2_15, B1=>nx9868);
   ix5329 : nand03 port map ( Y=>nx5328, A0=>nx8641, A1=>nx8643, A2=>nx8645
   );
   ix8642 : aoi222 port map ( Y=>nx8641, A0=>que_out_26_2_15, A1=>nx9816, B0
      =>que_out_14_2_15, B1=>nx9790, C0=>que_out_11_2_15, C1=>nx9764);
   ix8644 : aoi22 port map ( Y=>nx8643, A0=>que_out_13_2_15, A1=>nx9738, B0
      =>que_out_7_2_15, B1=>nx9712);
   ix8646 : aoi22 port map ( Y=>nx8645, A0=>que_out_12_2_15, A1=>nx9686, B0
      =>que_out_1_2_15, B1=>nx9660);
   ix5523 : or04 port map ( Y=>out_column_1_0, A0=>nx5518, A1=>nx5492, A2=>
      nx5464, A3=>nx5438);
   ix5519 : nand03 port map ( Y=>nx5518, A0=>nx8651, A1=>nx8653, A2=>nx8655
   );
   ix8652 : aoi222 port map ( Y=>nx8651, A0=>que_out_10_1_0, A1=>nx10310, B0
      =>que_out_6_1_0, B1=>nx10362, C0=>que_out_9_1_0, C1=>nx10336);
   ix8654 : aoi22 port map ( Y=>nx8653, A0=>que_out_5_1_0, A1=>nx10258, B0=>
      que_out_18_1_0, B1=>nx10284);
   ix8656 : aoi22 port map ( Y=>nx8655, A0=>que_out_17_1_0, A1=>nx10232, B0
      =>que_out_20_1_0, B1=>nx10206);
   ix5493 : nand03 port map ( Y=>nx5492, A0=>nx8659, A1=>nx8661, A2=>nx8663
   );
   ix8660 : aoi222 port map ( Y=>nx8659, A0=>que_out_19_1_0, A1=>nx10180, B0
      =>que_out_21_1_0, B1=>nx10154, C0=>que_out_8_1_0, C1=>nx10128);
   ix8662 : aoi22 port map ( Y=>nx8661, A0=>que_out_25_1_0, A1=>nx10076, B0
      =>que_out_16_1_0, B1=>nx10102);
   ix8664 : aoi22 port map ( Y=>nx8663, A0=>que_out_24_1_0, A1=>nx10050, B0
      =>que_out_22_1_0, B1=>nx10024);
   ix5465 : nand03 port map ( Y=>nx5464, A0=>nx8667, A1=>nx8669, A2=>nx8671
   );
   ix8668 : aoi222 port map ( Y=>nx8667, A0=>que_out_15_1_0, A1=>nx9972, B0
      =>que_out_3_1_0, B1=>nx9998, C0=>que_out_23_1_0, C1=>nx9946);
   ix8670 : aoi22 port map ( Y=>nx8669, A0=>que_out_27_1_0, A1=>nx9920, B0=>
      que_out_4_1_0, B1=>nx9894);
   ix8672 : aoi22 port map ( Y=>nx8671, A0=>que_out_0_1_0, A1=>nx9842, B0=>
      que_out_2_1_0, B1=>nx9868);
   ix5439 : nand03 port map ( Y=>nx5438, A0=>nx8675, A1=>nx8677, A2=>nx8679
   );
   ix8676 : aoi222 port map ( Y=>nx8675, A0=>que_out_26_1_0, A1=>nx9816, B0
      =>que_out_14_1_0, B1=>nx9790, C0=>que_out_11_1_0, C1=>nx9764);
   ix8678 : aoi22 port map ( Y=>nx8677, A0=>que_out_13_1_0, A1=>nx9738, B0=>
      que_out_7_1_0, B1=>nx9712);
   ix8680 : aoi22 port map ( Y=>nx8679, A0=>que_out_12_1_0, A1=>nx9686, B0=>
      que_out_1_1_0, B1=>nx9660);
   ix5633 : or04 port map ( Y=>out_column_1_1, A0=>nx5628, A1=>nx5602, A2=>
      nx5574, A3=>nx5548);
   ix5629 : nand03 port map ( Y=>nx5628, A0=>nx8685, A1=>nx8687, A2=>nx8689
   );
   ix8686 : aoi222 port map ( Y=>nx8685, A0=>que_out_10_1_1, A1=>nx10312, B0
      =>que_out_6_1_1, B1=>nx10364, C0=>que_out_9_1_1, C1=>nx10338);
   ix8688 : aoi22 port map ( Y=>nx8687, A0=>que_out_5_1_1, A1=>nx10260, B0=>
      que_out_18_1_1, B1=>nx10286);
   ix8690 : aoi22 port map ( Y=>nx8689, A0=>que_out_17_1_1, A1=>nx10234, B0
      =>que_out_20_1_1, B1=>nx10208);
   ix5603 : nand03 port map ( Y=>nx5602, A0=>nx8693, A1=>nx8695, A2=>nx8697
   );
   ix8694 : aoi222 port map ( Y=>nx8693, A0=>que_out_19_1_1, A1=>nx10182, B0
      =>que_out_21_1_1, B1=>nx10156, C0=>que_out_8_1_1, C1=>nx10130);
   ix8696 : aoi22 port map ( Y=>nx8695, A0=>que_out_25_1_1, A1=>nx10078, B0
      =>que_out_16_1_1, B1=>nx10104);
   ix8698 : aoi22 port map ( Y=>nx8697, A0=>que_out_24_1_1, A1=>nx10052, B0
      =>que_out_22_1_1, B1=>nx10026);
   ix5575 : nand03 port map ( Y=>nx5574, A0=>nx8701, A1=>nx8703, A2=>nx8705
   );
   ix8702 : aoi222 port map ( Y=>nx8701, A0=>que_out_15_1_1, A1=>nx9974, B0
      =>que_out_3_1_1, B1=>nx10000, C0=>que_out_23_1_1, C1=>nx9948);
   ix8704 : aoi22 port map ( Y=>nx8703, A0=>que_out_27_1_1, A1=>nx9922, B0=>
      que_out_4_1_1, B1=>nx9896);
   ix8706 : aoi22 port map ( Y=>nx8705, A0=>que_out_0_1_1, A1=>nx9844, B0=>
      que_out_2_1_1, B1=>nx9870);
   ix5549 : nand03 port map ( Y=>nx5548, A0=>nx8709, A1=>nx8711, A2=>nx8713
   );
   ix8710 : aoi222 port map ( Y=>nx8709, A0=>que_out_26_1_1, A1=>nx9818, B0
      =>que_out_14_1_1, B1=>nx9792, C0=>que_out_11_1_1, C1=>nx9766);
   ix8712 : aoi22 port map ( Y=>nx8711, A0=>que_out_13_1_1, A1=>nx9740, B0=>
      que_out_7_1_1, B1=>nx9714);
   ix8714 : aoi22 port map ( Y=>nx8713, A0=>que_out_12_1_1, A1=>nx9688, B0=>
      que_out_1_1_1, B1=>nx9662);
   ix5743 : or04 port map ( Y=>out_column_1_2, A0=>nx5738, A1=>nx5712, A2=>
      nx5684, A3=>nx5658);
   ix5739 : nand03 port map ( Y=>nx5738, A0=>nx8719, A1=>nx8721, A2=>nx8723
   );
   ix8720 : aoi222 port map ( Y=>nx8719, A0=>que_out_10_1_2, A1=>nx10312, B0
      =>que_out_6_1_2, B1=>nx10364, C0=>que_out_9_1_2, C1=>nx10338);
   ix8722 : aoi22 port map ( Y=>nx8721, A0=>que_out_5_1_2, A1=>nx10260, B0=>
      que_out_18_1_2, B1=>nx10286);
   ix8724 : aoi22 port map ( Y=>nx8723, A0=>que_out_17_1_2, A1=>nx10234, B0
      =>que_out_20_1_2, B1=>nx10208);
   ix5713 : nand03 port map ( Y=>nx5712, A0=>nx8727, A1=>nx8729, A2=>nx8731
   );
   ix8728 : aoi222 port map ( Y=>nx8727, A0=>que_out_19_1_2, A1=>nx10182, B0
      =>que_out_21_1_2, B1=>nx10156, C0=>que_out_8_1_2, C1=>nx10130);
   ix8730 : aoi22 port map ( Y=>nx8729, A0=>que_out_25_1_2, A1=>nx10078, B0
      =>que_out_16_1_2, B1=>nx10104);
   ix8732 : aoi22 port map ( Y=>nx8731, A0=>que_out_24_1_2, A1=>nx10052, B0
      =>que_out_22_1_2, B1=>nx10026);
   ix5685 : nand03 port map ( Y=>nx5684, A0=>nx8735, A1=>nx8737, A2=>nx8739
   );
   ix8736 : aoi222 port map ( Y=>nx8735, A0=>que_out_15_1_2, A1=>nx9974, B0
      =>que_out_3_1_2, B1=>nx10000, C0=>que_out_23_1_2, C1=>nx9948);
   ix8738 : aoi22 port map ( Y=>nx8737, A0=>que_out_27_1_2, A1=>nx9922, B0=>
      que_out_4_1_2, B1=>nx9896);
   ix8740 : aoi22 port map ( Y=>nx8739, A0=>que_out_0_1_2, A1=>nx9844, B0=>
      que_out_2_1_2, B1=>nx9870);
   ix5659 : nand03 port map ( Y=>nx5658, A0=>nx8743, A1=>nx8745, A2=>nx8747
   );
   ix8744 : aoi222 port map ( Y=>nx8743, A0=>que_out_26_1_2, A1=>nx9818, B0
      =>que_out_14_1_2, B1=>nx9792, C0=>que_out_11_1_2, C1=>nx9766);
   ix8746 : aoi22 port map ( Y=>nx8745, A0=>que_out_13_1_2, A1=>nx9740, B0=>
      que_out_7_1_2, B1=>nx9714);
   ix8748 : aoi22 port map ( Y=>nx8747, A0=>que_out_12_1_2, A1=>nx9688, B0=>
      que_out_1_1_2, B1=>nx9662);
   ix5853 : or04 port map ( Y=>out_column_1_3, A0=>nx5848, A1=>nx5822, A2=>
      nx5794, A3=>nx5768);
   ix5849 : nand03 port map ( Y=>nx5848, A0=>nx8753, A1=>nx8755, A2=>nx8757
   );
   ix8754 : aoi222 port map ( Y=>nx8753, A0=>que_out_10_1_3, A1=>nx10312, B0
      =>que_out_6_1_3, B1=>nx10364, C0=>que_out_9_1_3, C1=>nx10338);
   ix8756 : aoi22 port map ( Y=>nx8755, A0=>que_out_5_1_3, A1=>nx10260, B0=>
      que_out_18_1_3, B1=>nx10286);
   ix8758 : aoi22 port map ( Y=>nx8757, A0=>que_out_17_1_3, A1=>nx10234, B0
      =>que_out_20_1_3, B1=>nx10208);
   ix5823 : nand03 port map ( Y=>nx5822, A0=>nx8761, A1=>nx8763, A2=>nx8765
   );
   ix8762 : aoi222 port map ( Y=>nx8761, A0=>que_out_19_1_3, A1=>nx10182, B0
      =>que_out_21_1_3, B1=>nx10156, C0=>que_out_8_1_3, C1=>nx10130);
   ix8764 : aoi22 port map ( Y=>nx8763, A0=>que_out_25_1_3, A1=>nx10078, B0
      =>que_out_16_1_3, B1=>nx10104);
   ix8766 : aoi22 port map ( Y=>nx8765, A0=>que_out_24_1_3, A1=>nx10052, B0
      =>que_out_22_1_3, B1=>nx10026);
   ix5795 : nand03 port map ( Y=>nx5794, A0=>nx8769, A1=>nx8771, A2=>nx8773
   );
   ix8770 : aoi222 port map ( Y=>nx8769, A0=>que_out_15_1_3, A1=>nx9974, B0
      =>que_out_3_1_3, B1=>nx10000, C0=>que_out_23_1_3, C1=>nx9948);
   ix8772 : aoi22 port map ( Y=>nx8771, A0=>que_out_27_1_3, A1=>nx9922, B0=>
      que_out_4_1_3, B1=>nx9896);
   ix8774 : aoi22 port map ( Y=>nx8773, A0=>que_out_0_1_3, A1=>nx9844, B0=>
      que_out_2_1_3, B1=>nx9870);
   ix5769 : nand03 port map ( Y=>nx5768, A0=>nx8777, A1=>nx8779, A2=>nx8781
   );
   ix8778 : aoi222 port map ( Y=>nx8777, A0=>que_out_26_1_3, A1=>nx9818, B0
      =>que_out_14_1_3, B1=>nx9792, C0=>que_out_11_1_3, C1=>nx9766);
   ix8780 : aoi22 port map ( Y=>nx8779, A0=>que_out_13_1_3, A1=>nx9740, B0=>
      que_out_7_1_3, B1=>nx9714);
   ix8782 : aoi22 port map ( Y=>nx8781, A0=>que_out_12_1_3, A1=>nx9688, B0=>
      que_out_1_1_3, B1=>nx9662);
   ix5963 : or04 port map ( Y=>out_column_1_4, A0=>nx5958, A1=>nx5932, A2=>
      nx5904, A3=>nx5878);
   ix5959 : nand03 port map ( Y=>nx5958, A0=>nx8787, A1=>nx8789, A2=>nx8791
   );
   ix8788 : aoi222 port map ( Y=>nx8787, A0=>que_out_10_1_4, A1=>nx10312, B0
      =>que_out_6_1_4, B1=>nx10364, C0=>que_out_9_1_4, C1=>nx10338);
   ix8790 : aoi22 port map ( Y=>nx8789, A0=>que_out_5_1_4, A1=>nx10260, B0=>
      que_out_18_1_4, B1=>nx10286);
   ix8792 : aoi22 port map ( Y=>nx8791, A0=>que_out_17_1_4, A1=>nx10234, B0
      =>que_out_20_1_4, B1=>nx10208);
   ix5933 : nand03 port map ( Y=>nx5932, A0=>nx8795, A1=>nx8797, A2=>nx8799
   );
   ix8796 : aoi222 port map ( Y=>nx8795, A0=>que_out_19_1_4, A1=>nx10182, B0
      =>que_out_21_1_4, B1=>nx10156, C0=>que_out_8_1_4, C1=>nx10130);
   ix8798 : aoi22 port map ( Y=>nx8797, A0=>que_out_25_1_4, A1=>nx10078, B0
      =>que_out_16_1_4, B1=>nx10104);
   ix8800 : aoi22 port map ( Y=>nx8799, A0=>que_out_24_1_4, A1=>nx10052, B0
      =>que_out_22_1_4, B1=>nx10026);
   ix5905 : nand03 port map ( Y=>nx5904, A0=>nx8803, A1=>nx8805, A2=>nx8807
   );
   ix8804 : aoi222 port map ( Y=>nx8803, A0=>que_out_15_1_4, A1=>nx9974, B0
      =>que_out_3_1_4, B1=>nx10000, C0=>que_out_23_1_4, C1=>nx9948);
   ix8806 : aoi22 port map ( Y=>nx8805, A0=>que_out_27_1_4, A1=>nx9922, B0=>
      que_out_4_1_4, B1=>nx9896);
   ix8808 : aoi22 port map ( Y=>nx8807, A0=>que_out_0_1_4, A1=>nx9844, B0=>
      que_out_2_1_4, B1=>nx9870);
   ix5879 : nand03 port map ( Y=>nx5878, A0=>nx8811, A1=>nx8813, A2=>nx8815
   );
   ix8812 : aoi222 port map ( Y=>nx8811, A0=>que_out_26_1_4, A1=>nx9818, B0
      =>que_out_14_1_4, B1=>nx9792, C0=>que_out_11_1_4, C1=>nx9766);
   ix8814 : aoi22 port map ( Y=>nx8813, A0=>que_out_13_1_4, A1=>nx9740, B0=>
      que_out_7_1_4, B1=>nx9714);
   ix8816 : aoi22 port map ( Y=>nx8815, A0=>que_out_12_1_4, A1=>nx9688, B0=>
      que_out_1_1_4, B1=>nx9662);
   ix6073 : or04 port map ( Y=>out_column_1_5, A0=>nx6068, A1=>nx6042, A2=>
      nx6014, A3=>nx5988);
   ix6069 : nand03 port map ( Y=>nx6068, A0=>nx8821, A1=>nx8823, A2=>nx8825
   );
   ix8822 : aoi222 port map ( Y=>nx8821, A0=>que_out_10_1_5, A1=>nx10312, B0
      =>que_out_6_1_5, B1=>nx10364, C0=>que_out_9_1_5, C1=>nx10338);
   ix8824 : aoi22 port map ( Y=>nx8823, A0=>que_out_5_1_5, A1=>nx10260, B0=>
      que_out_18_1_5, B1=>nx10286);
   ix8826 : aoi22 port map ( Y=>nx8825, A0=>que_out_17_1_5, A1=>nx10234, B0
      =>que_out_20_1_5, B1=>nx10208);
   ix6043 : nand03 port map ( Y=>nx6042, A0=>nx8829, A1=>nx8831, A2=>nx8833
   );
   ix8830 : aoi222 port map ( Y=>nx8829, A0=>que_out_19_1_5, A1=>nx10182, B0
      =>que_out_21_1_5, B1=>nx10156, C0=>que_out_8_1_5, C1=>nx10130);
   ix8832 : aoi22 port map ( Y=>nx8831, A0=>que_out_25_1_5, A1=>nx10078, B0
      =>que_out_16_1_5, B1=>nx10104);
   ix8834 : aoi22 port map ( Y=>nx8833, A0=>que_out_24_1_5, A1=>nx10052, B0
      =>que_out_22_1_5, B1=>nx10026);
   ix6015 : nand03 port map ( Y=>nx6014, A0=>nx8837, A1=>nx8839, A2=>nx8841
   );
   ix8838 : aoi222 port map ( Y=>nx8837, A0=>que_out_15_1_5, A1=>nx9974, B0
      =>que_out_3_1_5, B1=>nx10000, C0=>que_out_23_1_5, C1=>nx9948);
   ix8840 : aoi22 port map ( Y=>nx8839, A0=>que_out_27_1_5, A1=>nx9922, B0=>
      que_out_4_1_5, B1=>nx9896);
   ix8842 : aoi22 port map ( Y=>nx8841, A0=>que_out_0_1_5, A1=>nx9844, B0=>
      que_out_2_1_5, B1=>nx9870);
   ix5989 : nand03 port map ( Y=>nx5988, A0=>nx8845, A1=>nx8847, A2=>nx8849
   );
   ix8846 : aoi222 port map ( Y=>nx8845, A0=>que_out_26_1_5, A1=>nx9818, B0
      =>que_out_14_1_5, B1=>nx9792, C0=>que_out_11_1_5, C1=>nx9766);
   ix8848 : aoi22 port map ( Y=>nx8847, A0=>que_out_13_1_5, A1=>nx9740, B0=>
      que_out_7_1_5, B1=>nx9714);
   ix8850 : aoi22 port map ( Y=>nx8849, A0=>que_out_12_1_5, A1=>nx9688, B0=>
      que_out_1_1_5, B1=>nx9662);
   ix6183 : or04 port map ( Y=>out_column_1_6, A0=>nx6178, A1=>nx6152, A2=>
      nx6124, A3=>nx6098);
   ix6179 : nand03 port map ( Y=>nx6178, A0=>nx8855, A1=>nx8857, A2=>nx8859
   );
   ix8856 : aoi222 port map ( Y=>nx8855, A0=>que_out_10_1_6, A1=>nx10312, B0
      =>que_out_6_1_6, B1=>nx10364, C0=>que_out_9_1_6, C1=>nx10338);
   ix8858 : aoi22 port map ( Y=>nx8857, A0=>que_out_5_1_6, A1=>nx10260, B0=>
      que_out_18_1_6, B1=>nx10286);
   ix8860 : aoi22 port map ( Y=>nx8859, A0=>que_out_17_1_6, A1=>nx10234, B0
      =>que_out_20_1_6, B1=>nx10208);
   ix6153 : nand03 port map ( Y=>nx6152, A0=>nx8863, A1=>nx8865, A2=>nx8867
   );
   ix8864 : aoi222 port map ( Y=>nx8863, A0=>que_out_19_1_6, A1=>nx10182, B0
      =>que_out_21_1_6, B1=>nx10156, C0=>que_out_8_1_6, C1=>nx10130);
   ix8866 : aoi22 port map ( Y=>nx8865, A0=>que_out_25_1_6, A1=>nx10078, B0
      =>que_out_16_1_6, B1=>nx10104);
   ix8868 : aoi22 port map ( Y=>nx8867, A0=>que_out_24_1_6, A1=>nx10052, B0
      =>que_out_22_1_6, B1=>nx10026);
   ix6125 : nand03 port map ( Y=>nx6124, A0=>nx8871, A1=>nx8873, A2=>nx8875
   );
   ix8872 : aoi222 port map ( Y=>nx8871, A0=>que_out_15_1_6, A1=>nx9974, B0
      =>que_out_3_1_6, B1=>nx10000, C0=>que_out_23_1_6, C1=>nx9948);
   ix8874 : aoi22 port map ( Y=>nx8873, A0=>que_out_27_1_6, A1=>nx9922, B0=>
      que_out_4_1_6, B1=>nx9896);
   ix8876 : aoi22 port map ( Y=>nx8875, A0=>que_out_0_1_6, A1=>nx9844, B0=>
      que_out_2_1_6, B1=>nx9870);
   ix6099 : nand03 port map ( Y=>nx6098, A0=>nx8879, A1=>nx8881, A2=>nx8883
   );
   ix8880 : aoi222 port map ( Y=>nx8879, A0=>que_out_26_1_6, A1=>nx9818, B0
      =>que_out_14_1_6, B1=>nx9792, C0=>que_out_11_1_6, C1=>nx9766);
   ix8882 : aoi22 port map ( Y=>nx8881, A0=>que_out_13_1_6, A1=>nx9740, B0=>
      que_out_7_1_6, B1=>nx9714);
   ix8884 : aoi22 port map ( Y=>nx8883, A0=>que_out_12_1_6, A1=>nx9688, B0=>
      que_out_1_1_6, B1=>nx9662);
   ix6293 : or04 port map ( Y=>out_column_1_7, A0=>nx6288, A1=>nx6262, A2=>
      nx6234, A3=>nx6208);
   ix6289 : nand03 port map ( Y=>nx6288, A0=>nx8889, A1=>nx8891, A2=>nx8893
   );
   ix8890 : aoi222 port map ( Y=>nx8889, A0=>que_out_10_1_7, A1=>nx10312, B0
      =>que_out_6_1_7, B1=>nx10364, C0=>que_out_9_1_7, C1=>nx10338);
   ix8892 : aoi22 port map ( Y=>nx8891, A0=>que_out_5_1_7, A1=>nx10260, B0=>
      que_out_18_1_7, B1=>nx10286);
   ix8894 : aoi22 port map ( Y=>nx8893, A0=>que_out_17_1_7, A1=>nx10234, B0
      =>que_out_20_1_7, B1=>nx10208);
   ix6263 : nand03 port map ( Y=>nx6262, A0=>nx8897, A1=>nx8899, A2=>nx8901
   );
   ix8898 : aoi222 port map ( Y=>nx8897, A0=>que_out_19_1_7, A1=>nx10182, B0
      =>que_out_21_1_7, B1=>nx10156, C0=>que_out_8_1_7, C1=>nx10130);
   ix8900 : aoi22 port map ( Y=>nx8899, A0=>que_out_25_1_7, A1=>nx10078, B0
      =>que_out_16_1_7, B1=>nx10104);
   ix8902 : aoi22 port map ( Y=>nx8901, A0=>que_out_24_1_7, A1=>nx10052, B0
      =>que_out_22_1_7, B1=>nx10026);
   ix6235 : nand03 port map ( Y=>nx6234, A0=>nx8905, A1=>nx8907, A2=>nx8909
   );
   ix8906 : aoi222 port map ( Y=>nx8905, A0=>que_out_15_1_7, A1=>nx9974, B0
      =>que_out_3_1_7, B1=>nx10000, C0=>que_out_23_1_7, C1=>nx9948);
   ix8908 : aoi22 port map ( Y=>nx8907, A0=>que_out_27_1_7, A1=>nx9922, B0=>
      que_out_4_1_7, B1=>nx9896);
   ix8910 : aoi22 port map ( Y=>nx8909, A0=>que_out_0_1_7, A1=>nx9844, B0=>
      que_out_2_1_7, B1=>nx9870);
   ix6209 : nand03 port map ( Y=>nx6208, A0=>nx8913, A1=>nx8915, A2=>nx8917
   );
   ix8914 : aoi222 port map ( Y=>nx8913, A0=>que_out_26_1_7, A1=>nx9818, B0
      =>que_out_14_1_7, B1=>nx9792, C0=>que_out_11_1_7, C1=>nx9766);
   ix8916 : aoi22 port map ( Y=>nx8915, A0=>que_out_13_1_7, A1=>nx9740, B0=>
      que_out_7_1_7, B1=>nx9714);
   ix8918 : aoi22 port map ( Y=>nx8917, A0=>que_out_12_1_7, A1=>nx9688, B0=>
      que_out_1_1_7, B1=>nx9662);
   ix6403 : or04 port map ( Y=>out_column_1_8, A0=>nx6398, A1=>nx6372, A2=>
      nx6344, A3=>nx6318);
   ix6399 : nand03 port map ( Y=>nx6398, A0=>nx8923, A1=>nx8925, A2=>nx8927
   );
   ix8924 : aoi222 port map ( Y=>nx8923, A0=>que_out_10_1_8, A1=>nx10314, B0
      =>que_out_6_1_8, B1=>nx10366, C0=>que_out_9_1_8, C1=>nx10340);
   ix8926 : aoi22 port map ( Y=>nx8925, A0=>que_out_5_1_8, A1=>nx10262, B0=>
      que_out_18_1_8, B1=>nx10288);
   ix8928 : aoi22 port map ( Y=>nx8927, A0=>que_out_17_1_8, A1=>nx10236, B0
      =>que_out_20_1_8, B1=>nx10210);
   ix6373 : nand03 port map ( Y=>nx6372, A0=>nx8931, A1=>nx8933, A2=>nx8935
   );
   ix8932 : aoi222 port map ( Y=>nx8931, A0=>que_out_19_1_8, A1=>nx10184, B0
      =>que_out_21_1_8, B1=>nx10158, C0=>que_out_8_1_8, C1=>nx10132);
   ix8934 : aoi22 port map ( Y=>nx8933, A0=>que_out_25_1_8, A1=>nx10080, B0
      =>que_out_16_1_8, B1=>nx10106);
   ix8936 : aoi22 port map ( Y=>nx8935, A0=>que_out_24_1_8, A1=>nx10054, B0
      =>que_out_22_1_8, B1=>nx10028);
   ix6345 : nand03 port map ( Y=>nx6344, A0=>nx8939, A1=>nx8941, A2=>nx8943
   );
   ix8940 : aoi222 port map ( Y=>nx8939, A0=>que_out_15_1_8, A1=>nx9976, B0
      =>que_out_3_1_8, B1=>nx10002, C0=>que_out_23_1_8, C1=>nx9950);
   ix8942 : aoi22 port map ( Y=>nx8941, A0=>que_out_27_1_8, A1=>nx9924, B0=>
      que_out_4_1_8, B1=>nx9898);
   ix8944 : aoi22 port map ( Y=>nx8943, A0=>que_out_0_1_8, A1=>nx9846, B0=>
      que_out_2_1_8, B1=>nx9872);
   ix6319 : nand03 port map ( Y=>nx6318, A0=>nx8947, A1=>nx8949, A2=>nx8951
   );
   ix8948 : aoi222 port map ( Y=>nx8947, A0=>que_out_26_1_8, A1=>nx9820, B0
      =>que_out_14_1_8, B1=>nx9794, C0=>que_out_11_1_8, C1=>nx9768);
   ix8950 : aoi22 port map ( Y=>nx8949, A0=>que_out_13_1_8, A1=>nx9742, B0=>
      que_out_7_1_8, B1=>nx9716);
   ix8952 : aoi22 port map ( Y=>nx8951, A0=>que_out_12_1_8, A1=>nx9690, B0=>
      que_out_1_1_8, B1=>nx9664);
   ix6513 : or04 port map ( Y=>out_column_1_9, A0=>nx6508, A1=>nx6482, A2=>
      nx6454, A3=>nx6428);
   ix6509 : nand03 port map ( Y=>nx6508, A0=>nx8955, A1=>nx8957, A2=>nx8959
   );
   ix8956 : aoi222 port map ( Y=>nx8955, A0=>que_out_10_1_9, A1=>nx10314, B0
      =>que_out_6_1_9, B1=>nx10366, C0=>que_out_9_1_9, C1=>nx10340);
   ix8958 : aoi22 port map ( Y=>nx8957, A0=>que_out_5_1_9, A1=>nx10262, B0=>
      que_out_18_1_9, B1=>nx10288);
   ix8960 : aoi22 port map ( Y=>nx8959, A0=>que_out_17_1_9, A1=>nx10236, B0
      =>que_out_20_1_9, B1=>nx10210);
   ix6483 : nand03 port map ( Y=>nx6482, A0=>nx8963, A1=>nx8965, A2=>nx8967
   );
   ix8964 : aoi222 port map ( Y=>nx8963, A0=>que_out_19_1_9, A1=>nx10184, B0
      =>que_out_21_1_9, B1=>nx10158, C0=>que_out_8_1_9, C1=>nx10132);
   ix8966 : aoi22 port map ( Y=>nx8965, A0=>que_out_25_1_9, A1=>nx10080, B0
      =>que_out_16_1_9, B1=>nx10106);
   ix8968 : aoi22 port map ( Y=>nx8967, A0=>que_out_24_1_9, A1=>nx10054, B0
      =>que_out_22_1_9, B1=>nx10028);
   ix6455 : nand03 port map ( Y=>nx6454, A0=>nx8970, A1=>nx8973, A2=>nx8975
   );
   ix8972 : aoi222 port map ( Y=>nx8970, A0=>que_out_15_1_9, A1=>nx9976, B0
      =>que_out_3_1_9, B1=>nx10002, C0=>que_out_23_1_9, C1=>nx9950);
   ix8974 : aoi22 port map ( Y=>nx8973, A0=>que_out_27_1_9, A1=>nx9924, B0=>
      que_out_4_1_9, B1=>nx9898);
   ix8976 : aoi22 port map ( Y=>nx8975, A0=>que_out_0_1_9, A1=>nx9846, B0=>
      que_out_2_1_9, B1=>nx9872);
   ix6429 : nand03 port map ( Y=>nx6428, A0=>nx8978, A1=>nx8981, A2=>nx8983
   );
   ix8980 : aoi222 port map ( Y=>nx8978, A0=>que_out_26_1_9, A1=>nx9820, B0
      =>que_out_14_1_9, B1=>nx9794, C0=>que_out_11_1_9, C1=>nx9768);
   ix8982 : aoi22 port map ( Y=>nx8981, A0=>que_out_13_1_9, A1=>nx9742, B0=>
      que_out_7_1_9, B1=>nx9716);
   ix8984 : aoi22 port map ( Y=>nx8983, A0=>que_out_12_1_9, A1=>nx9690, B0=>
      que_out_1_1_9, B1=>nx9664);
   ix6623 : or04 port map ( Y=>out_column_1_10, A0=>nx6618, A1=>nx6592, A2=>
      nx6564, A3=>nx6538);
   ix6619 : nand03 port map ( Y=>nx6618, A0=>nx8989, A1=>nx8991, A2=>nx8993
   );
   ix8990 : aoi222 port map ( Y=>nx8989, A0=>que_out_10_1_10, A1=>nx10314, 
      B0=>que_out_6_1_10, B1=>nx10366, C0=>que_out_9_1_10, C1=>nx10340);
   ix8992 : aoi22 port map ( Y=>nx8991, A0=>que_out_5_1_10, A1=>nx10262, B0
      =>que_out_18_1_10, B1=>nx10288);
   ix8994 : aoi22 port map ( Y=>nx8993, A0=>que_out_17_1_10, A1=>nx10236, B0
      =>que_out_20_1_10, B1=>nx10210);
   ix6593 : nand03 port map ( Y=>nx6592, A0=>nx8997, A1=>nx8999, A2=>nx9001
   );
   ix8998 : aoi222 port map ( Y=>nx8997, A0=>que_out_19_1_10, A1=>nx10184, 
      B0=>que_out_21_1_10, B1=>nx10158, C0=>que_out_8_1_10, C1=>nx10132);
   ix9000 : aoi22 port map ( Y=>nx8999, A0=>que_out_25_1_10, A1=>nx10080, B0
      =>que_out_16_1_10, B1=>nx10106);
   ix9002 : aoi22 port map ( Y=>nx9001, A0=>que_out_24_1_10, A1=>nx10054, B0
      =>que_out_22_1_10, B1=>nx10028);
   ix6565 : nand03 port map ( Y=>nx6564, A0=>nx9005, A1=>nx9007, A2=>nx9009
   );
   ix9006 : aoi222 port map ( Y=>nx9005, A0=>que_out_15_1_10, A1=>nx9976, B0
      =>que_out_3_1_10, B1=>nx10002, C0=>que_out_23_1_10, C1=>nx9950);
   ix9008 : aoi22 port map ( Y=>nx9007, A0=>que_out_27_1_10, A1=>nx9924, B0
      =>que_out_4_1_10, B1=>nx9898);
   ix9010 : aoi22 port map ( Y=>nx9009, A0=>que_out_0_1_10, A1=>nx9846, B0=>
      que_out_2_1_10, B1=>nx9872);
   ix6539 : nand03 port map ( Y=>nx6538, A0=>nx9013, A1=>nx9015, A2=>nx9017
   );
   ix9014 : aoi222 port map ( Y=>nx9013, A0=>que_out_26_1_10, A1=>nx9820, B0
      =>que_out_14_1_10, B1=>nx9794, C0=>que_out_11_1_10, C1=>nx9768);
   ix9016 : aoi22 port map ( Y=>nx9015, A0=>que_out_13_1_10, A1=>nx9742, B0
      =>que_out_7_1_10, B1=>nx9716);
   ix9018 : aoi22 port map ( Y=>nx9017, A0=>que_out_12_1_10, A1=>nx9690, B0
      =>que_out_1_1_10, B1=>nx9664);
   ix6733 : or04 port map ( Y=>out_column_1_11, A0=>nx6728, A1=>nx6702, A2=>
      nx6674, A3=>nx6648);
   ix6729 : nand03 port map ( Y=>nx6728, A0=>nx9023, A1=>nx9025, A2=>nx9027
   );
   ix9024 : aoi222 port map ( Y=>nx9023, A0=>que_out_10_1_11, A1=>nx10314, 
      B0=>que_out_6_1_11, B1=>nx10366, C0=>que_out_9_1_11, C1=>nx10340);
   ix9026 : aoi22 port map ( Y=>nx9025, A0=>que_out_5_1_11, A1=>nx10262, B0
      =>que_out_18_1_11, B1=>nx10288);
   ix9028 : aoi22 port map ( Y=>nx9027, A0=>que_out_17_1_11, A1=>nx10236, B0
      =>que_out_20_1_11, B1=>nx10210);
   ix6703 : nand03 port map ( Y=>nx6702, A0=>nx9031, A1=>nx9033, A2=>nx9035
   );
   ix9032 : aoi222 port map ( Y=>nx9031, A0=>que_out_19_1_11, A1=>nx10184, 
      B0=>que_out_21_1_11, B1=>nx10158, C0=>que_out_8_1_11, C1=>nx10132);
   ix9034 : aoi22 port map ( Y=>nx9033, A0=>que_out_25_1_11, A1=>nx10080, B0
      =>que_out_16_1_11, B1=>nx10106);
   ix9036 : aoi22 port map ( Y=>nx9035, A0=>que_out_24_1_11, A1=>nx10054, B0
      =>que_out_22_1_11, B1=>nx10028);
   ix6675 : nand03 port map ( Y=>nx6674, A0=>nx9039, A1=>nx9041, A2=>nx9043
   );
   ix9040 : aoi222 port map ( Y=>nx9039, A0=>que_out_15_1_11, A1=>nx9976, B0
      =>que_out_3_1_11, B1=>nx10002, C0=>que_out_23_1_11, C1=>nx9950);
   ix9042 : aoi22 port map ( Y=>nx9041, A0=>que_out_27_1_11, A1=>nx9924, B0
      =>que_out_4_1_11, B1=>nx9898);
   ix9044 : aoi22 port map ( Y=>nx9043, A0=>que_out_0_1_11, A1=>nx9846, B0=>
      que_out_2_1_11, B1=>nx9872);
   ix6649 : nand03 port map ( Y=>nx6648, A0=>nx9047, A1=>nx9049, A2=>nx9051
   );
   ix9048 : aoi222 port map ( Y=>nx9047, A0=>que_out_26_1_11, A1=>nx9820, B0
      =>que_out_14_1_11, B1=>nx9794, C0=>que_out_11_1_11, C1=>nx9768);
   ix9050 : aoi22 port map ( Y=>nx9049, A0=>que_out_13_1_11, A1=>nx9742, B0
      =>que_out_7_1_11, B1=>nx9716);
   ix9052 : aoi22 port map ( Y=>nx9051, A0=>que_out_12_1_11, A1=>nx9690, B0
      =>que_out_1_1_11, B1=>nx9664);
   ix6843 : or04 port map ( Y=>out_column_1_12, A0=>nx6838, A1=>nx6812, A2=>
      nx6784, A3=>nx6758);
   ix6839 : nand03 port map ( Y=>nx6838, A0=>nx9057, A1=>nx9059, A2=>nx9061
   );
   ix9058 : aoi222 port map ( Y=>nx9057, A0=>que_out_10_1_12, A1=>nx10314, 
      B0=>que_out_6_1_12, B1=>nx10366, C0=>que_out_9_1_12, C1=>nx10340);
   ix9060 : aoi22 port map ( Y=>nx9059, A0=>que_out_5_1_12, A1=>nx10262, B0
      =>que_out_18_1_12, B1=>nx10288);
   ix9062 : aoi22 port map ( Y=>nx9061, A0=>que_out_17_1_12, A1=>nx10236, B0
      =>que_out_20_1_12, B1=>nx10210);
   ix6813 : nand03 port map ( Y=>nx6812, A0=>nx9065, A1=>nx9067, A2=>nx9069
   );
   ix9066 : aoi222 port map ( Y=>nx9065, A0=>que_out_19_1_12, A1=>nx10184, 
      B0=>que_out_21_1_12, B1=>nx10158, C0=>que_out_8_1_12, C1=>nx10132);
   ix9068 : aoi22 port map ( Y=>nx9067, A0=>que_out_25_1_12, A1=>nx10080, B0
      =>que_out_16_1_12, B1=>nx10106);
   ix9070 : aoi22 port map ( Y=>nx9069, A0=>que_out_24_1_12, A1=>nx10054, B0
      =>que_out_22_1_12, B1=>nx10028);
   ix6785 : nand03 port map ( Y=>nx6784, A0=>nx9073, A1=>nx9075, A2=>nx9077
   );
   ix9074 : aoi222 port map ( Y=>nx9073, A0=>que_out_15_1_12, A1=>nx9976, B0
      =>que_out_3_1_12, B1=>nx10002, C0=>que_out_23_1_12, C1=>nx9950);
   ix9076 : aoi22 port map ( Y=>nx9075, A0=>que_out_27_1_12, A1=>nx9924, B0
      =>que_out_4_1_12, B1=>nx9898);
   ix9078 : aoi22 port map ( Y=>nx9077, A0=>que_out_0_1_12, A1=>nx9846, B0=>
      que_out_2_1_12, B1=>nx9872);
   ix6759 : nand03 port map ( Y=>nx6758, A0=>nx9081, A1=>nx9083, A2=>nx9085
   );
   ix9082 : aoi222 port map ( Y=>nx9081, A0=>que_out_26_1_12, A1=>nx9820, B0
      =>que_out_14_1_12, B1=>nx9794, C0=>que_out_11_1_12, C1=>nx9768);
   ix9084 : aoi22 port map ( Y=>nx9083, A0=>que_out_13_1_12, A1=>nx9742, B0
      =>que_out_7_1_12, B1=>nx9716);
   ix9086 : aoi22 port map ( Y=>nx9085, A0=>que_out_12_1_12, A1=>nx9690, B0
      =>que_out_1_1_12, B1=>nx9664);
   ix6953 : or04 port map ( Y=>out_column_1_13, A0=>nx6948, A1=>nx6922, A2=>
      nx6894, A3=>nx6868);
   ix6949 : nand03 port map ( Y=>nx6948, A0=>nx9090, A1=>nx9093, A2=>nx9095
   );
   ix9092 : aoi222 port map ( Y=>nx9090, A0=>que_out_10_1_13, A1=>nx10314, 
      B0=>que_out_6_1_13, B1=>nx10366, C0=>que_out_9_1_13, C1=>nx10340);
   ix9094 : aoi22 port map ( Y=>nx9093, A0=>que_out_5_1_13, A1=>nx10262, B0
      =>que_out_18_1_13, B1=>nx10288);
   ix9096 : aoi22 port map ( Y=>nx9095, A0=>que_out_17_1_13, A1=>nx10236, B0
      =>que_out_20_1_13, B1=>nx10210);
   ix6923 : nand03 port map ( Y=>nx6922, A0=>nx9098, A1=>nx9101, A2=>nx9103
   );
   ix9100 : aoi222 port map ( Y=>nx9098, A0=>que_out_19_1_13, A1=>nx10184, 
      B0=>que_out_21_1_13, B1=>nx10158, C0=>que_out_8_1_13, C1=>nx10132);
   ix9102 : aoi22 port map ( Y=>nx9101, A0=>que_out_25_1_13, A1=>nx10080, B0
      =>que_out_16_1_13, B1=>nx10106);
   ix9104 : aoi22 port map ( Y=>nx9103, A0=>que_out_24_1_13, A1=>nx10054, B0
      =>que_out_22_1_13, B1=>nx10028);
   ix6895 : nand03 port map ( Y=>nx6894, A0=>nx9106, A1=>nx9108, A2=>nx9110
   );
   ix9107 : aoi222 port map ( Y=>nx9106, A0=>que_out_15_1_13, A1=>nx9976, B0
      =>que_out_3_1_13, B1=>nx10002, C0=>que_out_23_1_13, C1=>nx9950);
   ix9109 : aoi22 port map ( Y=>nx9108, A0=>que_out_27_1_13, A1=>nx9924, B0
      =>que_out_4_1_13, B1=>nx9898);
   ix9111 : aoi22 port map ( Y=>nx9110, A0=>que_out_0_1_13, A1=>nx9846, B0=>
      que_out_2_1_13, B1=>nx9872);
   ix6869 : nand03 port map ( Y=>nx6868, A0=>nx9113, A1=>nx9115, A2=>nx9117
   );
   ix9114 : aoi222 port map ( Y=>nx9113, A0=>que_out_26_1_13, A1=>nx9820, B0
      =>que_out_14_1_13, B1=>nx9794, C0=>que_out_11_1_13, C1=>nx9768);
   ix9116 : aoi22 port map ( Y=>nx9115, A0=>que_out_13_1_13, A1=>nx9742, B0
      =>que_out_7_1_13, B1=>nx9716);
   ix9118 : aoi22 port map ( Y=>nx9117, A0=>que_out_12_1_13, A1=>nx9690, B0
      =>que_out_1_1_13, B1=>nx9664);
   ix7063 : or04 port map ( Y=>out_column_1_14, A0=>nx7058, A1=>nx7032, A2=>
      nx7004, A3=>nx6978);
   ix7059 : nand03 port map ( Y=>nx7058, A0=>nx9121, A1=>nx9123, A2=>nx9125
   );
   ix9122 : aoi222 port map ( Y=>nx9121, A0=>que_out_10_1_14, A1=>nx10314, 
      B0=>que_out_6_1_14, B1=>nx10366, C0=>que_out_9_1_14, C1=>nx10340);
   ix9124 : aoi22 port map ( Y=>nx9123, A0=>que_out_5_1_14, A1=>nx10262, B0
      =>que_out_18_1_14, B1=>nx10288);
   ix9126 : aoi22 port map ( Y=>nx9125, A0=>que_out_17_1_14, A1=>nx10236, B0
      =>que_out_20_1_14, B1=>nx10210);
   ix7033 : nand03 port map ( Y=>nx7032, A0=>nx9128, A1=>nx9130, A2=>nx9132
   );
   ix9129 : aoi222 port map ( Y=>nx9128, A0=>que_out_19_1_14, A1=>nx10184, 
      B0=>que_out_21_1_14, B1=>nx10158, C0=>que_out_8_1_14, C1=>nx10132);
   ix9131 : aoi22 port map ( Y=>nx9130, A0=>que_out_25_1_14, A1=>nx10080, B0
      =>que_out_16_1_14, B1=>nx10106);
   ix9133 : aoi22 port map ( Y=>nx9132, A0=>que_out_24_1_14, A1=>nx10054, B0
      =>que_out_22_1_14, B1=>nx10028);
   ix7005 : nand03 port map ( Y=>nx7004, A0=>nx9135, A1=>nx9137, A2=>nx9139
   );
   ix9136 : aoi222 port map ( Y=>nx9135, A0=>que_out_15_1_14, A1=>nx9976, B0
      =>que_out_3_1_14, B1=>nx10002, C0=>que_out_23_1_14, C1=>nx9950);
   ix9138 : aoi22 port map ( Y=>nx9137, A0=>que_out_27_1_14, A1=>nx9924, B0
      =>que_out_4_1_14, B1=>nx9898);
   ix9140 : aoi22 port map ( Y=>nx9139, A0=>que_out_0_1_14, A1=>nx9846, B0=>
      que_out_2_1_14, B1=>nx9872);
   ix6979 : nand03 port map ( Y=>nx6978, A0=>nx9142, A1=>nx9144, A2=>nx9146
   );
   ix9143 : aoi222 port map ( Y=>nx9142, A0=>que_out_26_1_14, A1=>nx9820, B0
      =>que_out_14_1_14, B1=>nx9794, C0=>que_out_11_1_14, C1=>nx9768);
   ix9145 : aoi22 port map ( Y=>nx9144, A0=>que_out_13_1_14, A1=>nx9742, B0
      =>que_out_7_1_14, B1=>nx9716);
   ix9147 : aoi22 port map ( Y=>nx9146, A0=>que_out_12_1_14, A1=>nx9690, B0
      =>que_out_1_1_14, B1=>nx9664);
   ix7173 : or04 port map ( Y=>out_column_1_15, A0=>nx7168, A1=>nx7142, A2=>
      nx7114, A3=>nx7088);
   ix7169 : nand03 port map ( Y=>nx7168, A0=>nx9150, A1=>nx9152, A2=>nx9154
   );
   ix9151 : aoi222 port map ( Y=>nx9150, A0=>que_out_10_1_15, A1=>nx10316, 
      B0=>que_out_6_1_15, B1=>nx10368, C0=>que_out_9_1_15, C1=>nx10342);
   ix9153 : aoi22 port map ( Y=>nx9152, A0=>que_out_5_1_15, A1=>nx10264, B0
      =>que_out_18_1_15, B1=>nx10290);
   ix9155 : aoi22 port map ( Y=>nx9154, A0=>que_out_17_1_15, A1=>nx10238, B0
      =>que_out_20_1_15, B1=>nx10212);
   ix7143 : nand03 port map ( Y=>nx7142, A0=>nx9157, A1=>nx9159, A2=>nx9161
   );
   ix9158 : aoi222 port map ( Y=>nx9157, A0=>que_out_19_1_15, A1=>nx10186, 
      B0=>que_out_21_1_15, B1=>nx10160, C0=>que_out_8_1_15, C1=>nx10134);
   ix9160 : aoi22 port map ( Y=>nx9159, A0=>que_out_25_1_15, A1=>nx10082, B0
      =>que_out_16_1_15, B1=>nx10108);
   ix9162 : aoi22 port map ( Y=>nx9161, A0=>que_out_24_1_15, A1=>nx10056, B0
      =>que_out_22_1_15, B1=>nx10030);
   ix7115 : nand03 port map ( Y=>nx7114, A0=>nx9164, A1=>nx9166, A2=>nx9168
   );
   ix9165 : aoi222 port map ( Y=>nx9164, A0=>que_out_15_1_15, A1=>nx9978, B0
      =>que_out_3_1_15, B1=>nx10004, C0=>que_out_23_1_15, C1=>nx9952);
   ix9167 : aoi22 port map ( Y=>nx9166, A0=>que_out_27_1_15, A1=>nx9926, B0
      =>que_out_4_1_15, B1=>nx9900);
   ix9169 : aoi22 port map ( Y=>nx9168, A0=>que_out_0_1_15, A1=>nx9848, B0=>
      que_out_2_1_15, B1=>nx9874);
   ix7089 : nand03 port map ( Y=>nx7088, A0=>nx9171, A1=>nx9173, A2=>nx9175
   );
   ix9172 : aoi222 port map ( Y=>nx9171, A0=>que_out_26_1_15, A1=>nx9822, B0
      =>que_out_14_1_15, B1=>nx9796, C0=>que_out_11_1_15, C1=>nx9770);
   ix9174 : aoi22 port map ( Y=>nx9173, A0=>que_out_13_1_15, A1=>nx9744, B0
      =>que_out_7_1_15, B1=>nx9718);
   ix9176 : aoi22 port map ( Y=>nx9175, A0=>que_out_12_1_15, A1=>nx9692, B0
      =>que_out_1_1_15, B1=>nx9666);
   ix7283 : or04 port map ( Y=>out_column_0_0, A0=>nx7278, A1=>nx7252, A2=>
      nx7224, A3=>nx7198);
   ix7279 : nand03 port map ( Y=>nx7278, A0=>nx9179, A1=>nx9181, A2=>nx9183
   );
   ix9180 : aoi222 port map ( Y=>nx9179, A0=>que_out_10_0_0, A1=>nx10316, B0
      =>que_out_6_0_0, B1=>nx10368, C0=>que_out_9_0_0, C1=>nx10342);
   ix9182 : aoi22 port map ( Y=>nx9181, A0=>que_out_5_0_0, A1=>nx10264, B0=>
      que_out_18_0_0, B1=>nx10290);
   ix9184 : aoi22 port map ( Y=>nx9183, A0=>que_out_17_0_0, A1=>nx10238, B0
      =>que_out_20_0_0, B1=>nx10212);
   ix7253 : nand03 port map ( Y=>nx7252, A0=>nx9186, A1=>nx9188, A2=>nx9190
   );
   ix9187 : aoi222 port map ( Y=>nx9186, A0=>que_out_19_0_0, A1=>nx10186, B0
      =>que_out_21_0_0, B1=>nx10160, C0=>que_out_8_0_0, C1=>nx10134);
   ix9189 : aoi22 port map ( Y=>nx9188, A0=>que_out_25_0_0, A1=>nx10082, B0
      =>que_out_16_0_0, B1=>nx10108);
   ix9191 : aoi22 port map ( Y=>nx9190, A0=>que_out_24_0_0, A1=>nx10056, B0
      =>que_out_22_0_0, B1=>nx10030);
   ix7225 : nand03 port map ( Y=>nx7224, A0=>nx9193, A1=>nx9195, A2=>nx9197
   );
   ix9194 : aoi222 port map ( Y=>nx9193, A0=>que_out_15_0_0, A1=>nx9978, B0
      =>que_out_3_0_0, B1=>nx10004, C0=>que_out_23_0_0, C1=>nx9952);
   ix9196 : aoi22 port map ( Y=>nx9195, A0=>que_out_27_0_0, A1=>nx9926, B0=>
      que_out_4_0_0, B1=>nx9900);
   ix9198 : aoi22 port map ( Y=>nx9197, A0=>que_out_0_0_0, A1=>nx9848, B0=>
      que_out_2_0_0, B1=>nx9874);
   ix7199 : nand03 port map ( Y=>nx7198, A0=>nx9200, A1=>nx9202, A2=>nx9204
   );
   ix9201 : aoi222 port map ( Y=>nx9200, A0=>que_out_26_0_0, A1=>nx9822, B0
      =>que_out_14_0_0, B1=>nx9796, C0=>que_out_11_0_0, C1=>nx9770);
   ix9203 : aoi22 port map ( Y=>nx9202, A0=>que_out_13_0_0, A1=>nx9744, B0=>
      que_out_7_0_0, B1=>nx9718);
   ix9205 : aoi22 port map ( Y=>nx9204, A0=>que_out_12_0_0, A1=>nx9692, B0=>
      que_out_1_0_0, B1=>nx9666);
   ix7393 : or04 port map ( Y=>out_column_0_1, A0=>nx7388, A1=>nx7362, A2=>
      nx7334, A3=>nx7308);
   ix7389 : nand03 port map ( Y=>nx7388, A0=>nx9208, A1=>nx9210, A2=>nx9212
   );
   ix9209 : aoi222 port map ( Y=>nx9208, A0=>que_out_10_0_1, A1=>nx10316, B0
      =>que_out_6_0_1, B1=>nx10368, C0=>que_out_9_0_1, C1=>nx10342);
   ix9211 : aoi22 port map ( Y=>nx9210, A0=>que_out_5_0_1, A1=>nx10264, B0=>
      que_out_18_0_1, B1=>nx10290);
   ix9213 : aoi22 port map ( Y=>nx9212, A0=>que_out_17_0_1, A1=>nx10238, B0
      =>que_out_20_0_1, B1=>nx10212);
   ix7363 : nand03 port map ( Y=>nx7362, A0=>nx9215, A1=>nx9217, A2=>nx9219
   );
   ix9216 : aoi222 port map ( Y=>nx9215, A0=>que_out_19_0_1, A1=>nx10186, B0
      =>que_out_21_0_1, B1=>nx10160, C0=>que_out_8_0_1, C1=>nx10134);
   ix9218 : aoi22 port map ( Y=>nx9217, A0=>que_out_25_0_1, A1=>nx10082, B0
      =>que_out_16_0_1, B1=>nx10108);
   ix9220 : aoi22 port map ( Y=>nx9219, A0=>que_out_24_0_1, A1=>nx10056, B0
      =>que_out_22_0_1, B1=>nx10030);
   ix7335 : nand03 port map ( Y=>nx7334, A0=>nx9222, A1=>nx9224, A2=>nx9226
   );
   ix9223 : aoi222 port map ( Y=>nx9222, A0=>que_out_15_0_1, A1=>nx9978, B0
      =>que_out_3_0_1, B1=>nx10004, C0=>que_out_23_0_1, C1=>nx9952);
   ix9225 : aoi22 port map ( Y=>nx9224, A0=>que_out_27_0_1, A1=>nx9926, B0=>
      que_out_4_0_1, B1=>nx9900);
   ix9227 : aoi22 port map ( Y=>nx9226, A0=>que_out_0_0_1, A1=>nx9848, B0=>
      que_out_2_0_1, B1=>nx9874);
   ix7309 : nand03 port map ( Y=>nx7308, A0=>nx9229, A1=>nx9231, A2=>nx9233
   );
   ix9230 : aoi222 port map ( Y=>nx9229, A0=>que_out_26_0_1, A1=>nx9822, B0
      =>que_out_14_0_1, B1=>nx9796, C0=>que_out_11_0_1, C1=>nx9770);
   ix9232 : aoi22 port map ( Y=>nx9231, A0=>que_out_13_0_1, A1=>nx9744, B0=>
      que_out_7_0_1, B1=>nx9718);
   ix9234 : aoi22 port map ( Y=>nx9233, A0=>que_out_12_0_1, A1=>nx9692, B0=>
      que_out_1_0_1, B1=>nx9666);
   ix7503 : or04 port map ( Y=>out_column_0_2, A0=>nx7498, A1=>nx7472, A2=>
      nx7444, A3=>nx7418);
   ix7499 : nand03 port map ( Y=>nx7498, A0=>nx9237, A1=>nx9239, A2=>nx9241
   );
   ix9238 : aoi222 port map ( Y=>nx9237, A0=>que_out_10_0_2, A1=>nx10316, B0
      =>que_out_6_0_2, B1=>nx10368, C0=>que_out_9_0_2, C1=>nx10342);
   ix9240 : aoi22 port map ( Y=>nx9239, A0=>que_out_5_0_2, A1=>nx10264, B0=>
      que_out_18_0_2, B1=>nx10290);
   ix9242 : aoi22 port map ( Y=>nx9241, A0=>que_out_17_0_2, A1=>nx10238, B0
      =>que_out_20_0_2, B1=>nx10212);
   ix7473 : nand03 port map ( Y=>nx7472, A0=>nx9244, A1=>nx9246, A2=>nx9248
   );
   ix9245 : aoi222 port map ( Y=>nx9244, A0=>que_out_19_0_2, A1=>nx10186, B0
      =>que_out_21_0_2, B1=>nx10160, C0=>que_out_8_0_2, C1=>nx10134);
   ix9247 : aoi22 port map ( Y=>nx9246, A0=>que_out_25_0_2, A1=>nx10082, B0
      =>que_out_16_0_2, B1=>nx10108);
   ix9249 : aoi22 port map ( Y=>nx9248, A0=>que_out_24_0_2, A1=>nx10056, B0
      =>que_out_22_0_2, B1=>nx10030);
   ix7445 : nand03 port map ( Y=>nx7444, A0=>nx9251, A1=>nx9253, A2=>nx9255
   );
   ix9252 : aoi222 port map ( Y=>nx9251, A0=>que_out_15_0_2, A1=>nx9978, B0
      =>que_out_3_0_2, B1=>nx10004, C0=>que_out_23_0_2, C1=>nx9952);
   ix9254 : aoi22 port map ( Y=>nx9253, A0=>que_out_27_0_2, A1=>nx9926, B0=>
      que_out_4_0_2, B1=>nx9900);
   ix9256 : aoi22 port map ( Y=>nx9255, A0=>que_out_0_0_2, A1=>nx9848, B0=>
      que_out_2_0_2, B1=>nx9874);
   ix7419 : nand03 port map ( Y=>nx7418, A0=>nx9258, A1=>nx9260, A2=>nx9262
   );
   ix9259 : aoi222 port map ( Y=>nx9258, A0=>que_out_26_0_2, A1=>nx9822, B0
      =>que_out_14_0_2, B1=>nx9796, C0=>que_out_11_0_2, C1=>nx9770);
   ix9261 : aoi22 port map ( Y=>nx9260, A0=>que_out_13_0_2, A1=>nx9744, B0=>
      que_out_7_0_2, B1=>nx9718);
   ix9263 : aoi22 port map ( Y=>nx9262, A0=>que_out_12_0_2, A1=>nx9692, B0=>
      que_out_1_0_2, B1=>nx9666);
   ix7613 : or04 port map ( Y=>out_column_0_3, A0=>nx7608, A1=>nx7582, A2=>
      nx7554, A3=>nx7528);
   ix7609 : nand03 port map ( Y=>nx7608, A0=>nx9266, A1=>nx9268, A2=>nx9270
   );
   ix9267 : aoi222 port map ( Y=>nx9266, A0=>que_out_10_0_3, A1=>nx10316, B0
      =>que_out_6_0_3, B1=>nx10368, C0=>que_out_9_0_3, C1=>nx10342);
   ix9269 : aoi22 port map ( Y=>nx9268, A0=>que_out_5_0_3, A1=>nx10264, B0=>
      que_out_18_0_3, B1=>nx10290);
   ix9271 : aoi22 port map ( Y=>nx9270, A0=>que_out_17_0_3, A1=>nx10238, B0
      =>que_out_20_0_3, B1=>nx10212);
   ix7583 : nand03 port map ( Y=>nx7582, A0=>nx9273, A1=>nx9275, A2=>nx9277
   );
   ix9274 : aoi222 port map ( Y=>nx9273, A0=>que_out_19_0_3, A1=>nx10186, B0
      =>que_out_21_0_3, B1=>nx10160, C0=>que_out_8_0_3, C1=>nx10134);
   ix9276 : aoi22 port map ( Y=>nx9275, A0=>que_out_25_0_3, A1=>nx10082, B0
      =>que_out_16_0_3, B1=>nx10108);
   ix9278 : aoi22 port map ( Y=>nx9277, A0=>que_out_24_0_3, A1=>nx10056, B0
      =>que_out_22_0_3, B1=>nx10030);
   ix7555 : nand03 port map ( Y=>nx7554, A0=>nx9280, A1=>nx9282, A2=>nx9284
   );
   ix9281 : aoi222 port map ( Y=>nx9280, A0=>que_out_15_0_3, A1=>nx9978, B0
      =>que_out_3_0_3, B1=>nx10004, C0=>que_out_23_0_3, C1=>nx9952);
   ix9283 : aoi22 port map ( Y=>nx9282, A0=>que_out_27_0_3, A1=>nx9926, B0=>
      que_out_4_0_3, B1=>nx9900);
   ix9285 : aoi22 port map ( Y=>nx9284, A0=>que_out_0_0_3, A1=>nx9848, B0=>
      que_out_2_0_3, B1=>nx9874);
   ix7529 : nand03 port map ( Y=>nx7528, A0=>nx9287, A1=>nx9289, A2=>nx9291
   );
   ix9288 : aoi222 port map ( Y=>nx9287, A0=>que_out_26_0_3, A1=>nx9822, B0
      =>que_out_14_0_3, B1=>nx9796, C0=>que_out_11_0_3, C1=>nx9770);
   ix9290 : aoi22 port map ( Y=>nx9289, A0=>que_out_13_0_3, A1=>nx9744, B0=>
      que_out_7_0_3, B1=>nx9718);
   ix9292 : aoi22 port map ( Y=>nx9291, A0=>que_out_12_0_3, A1=>nx9692, B0=>
      que_out_1_0_3, B1=>nx9666);
   ix7723 : or04 port map ( Y=>out_column_0_4, A0=>nx7718, A1=>nx7692, A2=>
      nx7664, A3=>nx7638);
   ix7719 : nand03 port map ( Y=>nx7718, A0=>nx9295, A1=>nx9297, A2=>nx9299
   );
   ix9296 : aoi222 port map ( Y=>nx9295, A0=>que_out_10_0_4, A1=>nx10316, B0
      =>que_out_6_0_4, B1=>nx10368, C0=>que_out_9_0_4, C1=>nx10342);
   ix9298 : aoi22 port map ( Y=>nx9297, A0=>que_out_5_0_4, A1=>nx10264, B0=>
      que_out_18_0_4, B1=>nx10290);
   ix9300 : aoi22 port map ( Y=>nx9299, A0=>que_out_17_0_4, A1=>nx10238, B0
      =>que_out_20_0_4, B1=>nx10212);
   ix7693 : nand03 port map ( Y=>nx7692, A0=>nx9302, A1=>nx9304, A2=>nx9306
   );
   ix9303 : aoi222 port map ( Y=>nx9302, A0=>que_out_19_0_4, A1=>nx10186, B0
      =>que_out_21_0_4, B1=>nx10160, C0=>que_out_8_0_4, C1=>nx10134);
   ix9305 : aoi22 port map ( Y=>nx9304, A0=>que_out_25_0_4, A1=>nx10082, B0
      =>que_out_16_0_4, B1=>nx10108);
   ix9307 : aoi22 port map ( Y=>nx9306, A0=>que_out_24_0_4, A1=>nx10056, B0
      =>que_out_22_0_4, B1=>nx10030);
   ix7665 : nand03 port map ( Y=>nx7664, A0=>nx9309, A1=>nx9311, A2=>nx9313
   );
   ix9310 : aoi222 port map ( Y=>nx9309, A0=>que_out_15_0_4, A1=>nx9978, B0
      =>que_out_3_0_4, B1=>nx10004, C0=>que_out_23_0_4, C1=>nx9952);
   ix9312 : aoi22 port map ( Y=>nx9311, A0=>que_out_27_0_4, A1=>nx9926, B0=>
      que_out_4_0_4, B1=>nx9900);
   ix9314 : aoi22 port map ( Y=>nx9313, A0=>que_out_0_0_4, A1=>nx9848, B0=>
      que_out_2_0_4, B1=>nx9874);
   ix7639 : nand03 port map ( Y=>nx7638, A0=>nx9316, A1=>nx9318, A2=>nx9320
   );
   ix9317 : aoi222 port map ( Y=>nx9316, A0=>que_out_26_0_4, A1=>nx9822, B0
      =>que_out_14_0_4, B1=>nx9796, C0=>que_out_11_0_4, C1=>nx9770);
   ix9319 : aoi22 port map ( Y=>nx9318, A0=>que_out_13_0_4, A1=>nx9744, B0=>
      que_out_7_0_4, B1=>nx9718);
   ix9321 : aoi22 port map ( Y=>nx9320, A0=>que_out_12_0_4, A1=>nx9692, B0=>
      que_out_1_0_4, B1=>nx9666);
   ix7833 : or04 port map ( Y=>out_column_0_5, A0=>nx7828, A1=>nx7802, A2=>
      nx7774, A3=>nx7748);
   ix7829 : nand03 port map ( Y=>nx7828, A0=>nx9324, A1=>nx9326, A2=>nx9328
   );
   ix9325 : aoi222 port map ( Y=>nx9324, A0=>que_out_10_0_5, A1=>nx10316, B0
      =>que_out_6_0_5, B1=>nx10368, C0=>que_out_9_0_5, C1=>nx10342);
   ix9327 : aoi22 port map ( Y=>nx9326, A0=>que_out_5_0_5, A1=>nx10264, B0=>
      que_out_18_0_5, B1=>nx10290);
   ix9329 : aoi22 port map ( Y=>nx9328, A0=>que_out_17_0_5, A1=>nx10238, B0
      =>que_out_20_0_5, B1=>nx10212);
   ix7803 : nand03 port map ( Y=>nx7802, A0=>nx9331, A1=>nx9333, A2=>nx9335
   );
   ix9332 : aoi222 port map ( Y=>nx9331, A0=>que_out_19_0_5, A1=>nx10186, B0
      =>que_out_21_0_5, B1=>nx10160, C0=>que_out_8_0_5, C1=>nx10134);
   ix9334 : aoi22 port map ( Y=>nx9333, A0=>que_out_25_0_5, A1=>nx10082, B0
      =>que_out_16_0_5, B1=>nx10108);
   ix9336 : aoi22 port map ( Y=>nx9335, A0=>que_out_24_0_5, A1=>nx10056, B0
      =>que_out_22_0_5, B1=>nx10030);
   ix7775 : nand03 port map ( Y=>nx7774, A0=>nx9338, A1=>nx9340, A2=>nx9342
   );
   ix9339 : aoi222 port map ( Y=>nx9338, A0=>que_out_15_0_5, A1=>nx9978, B0
      =>que_out_3_0_5, B1=>nx10004, C0=>que_out_23_0_5, C1=>nx9952);
   ix9341 : aoi22 port map ( Y=>nx9340, A0=>que_out_27_0_5, A1=>nx9926, B0=>
      que_out_4_0_5, B1=>nx9900);
   ix9343 : aoi22 port map ( Y=>nx9342, A0=>que_out_0_0_5, A1=>nx9848, B0=>
      que_out_2_0_5, B1=>nx9874);
   ix7749 : nand03 port map ( Y=>nx7748, A0=>nx9345, A1=>nx9347, A2=>nx9349
   );
   ix9346 : aoi222 port map ( Y=>nx9345, A0=>que_out_26_0_5, A1=>nx9822, B0
      =>que_out_14_0_5, B1=>nx9796, C0=>que_out_11_0_5, C1=>nx9770);
   ix9348 : aoi22 port map ( Y=>nx9347, A0=>que_out_13_0_5, A1=>nx9744, B0=>
      que_out_7_0_5, B1=>nx9718);
   ix9350 : aoi22 port map ( Y=>nx9349, A0=>que_out_12_0_5, A1=>nx9692, B0=>
      que_out_1_0_5, B1=>nx9666);
   ix7943 : or04 port map ( Y=>out_column_0_6, A0=>nx7938, A1=>nx7912, A2=>
      nx7884, A3=>nx7858);
   ix7939 : nand03 port map ( Y=>nx7938, A0=>nx9353, A1=>nx9355, A2=>nx9357
   );
   ix9354 : aoi222 port map ( Y=>nx9353, A0=>que_out_10_0_6, A1=>nx10318, B0
      =>que_out_6_0_6, B1=>nx10370, C0=>que_out_9_0_6, C1=>nx10344);
   ix9356 : aoi22 port map ( Y=>nx9355, A0=>que_out_5_0_6, A1=>nx10266, B0=>
      que_out_18_0_6, B1=>nx10292);
   ix9358 : aoi22 port map ( Y=>nx9357, A0=>que_out_17_0_6, A1=>nx10240, B0
      =>que_out_20_0_6, B1=>nx10214);
   ix7913 : nand03 port map ( Y=>nx7912, A0=>nx9360, A1=>nx9362, A2=>nx9364
   );
   ix9361 : aoi222 port map ( Y=>nx9360, A0=>que_out_19_0_6, A1=>nx10188, B0
      =>que_out_21_0_6, B1=>nx10162, C0=>que_out_8_0_6, C1=>nx10136);
   ix9363 : aoi22 port map ( Y=>nx9362, A0=>que_out_25_0_6, A1=>nx10084, B0
      =>que_out_16_0_6, B1=>nx10110);
   ix9365 : aoi22 port map ( Y=>nx9364, A0=>que_out_24_0_6, A1=>nx10058, B0
      =>que_out_22_0_6, B1=>nx10032);
   ix7885 : nand03 port map ( Y=>nx7884, A0=>nx9367, A1=>nx9369, A2=>nx9371
   );
   ix9368 : aoi222 port map ( Y=>nx9367, A0=>que_out_15_0_6, A1=>nx9980, B0
      =>que_out_3_0_6, B1=>nx10006, C0=>que_out_23_0_6, C1=>nx9954);
   ix9370 : aoi22 port map ( Y=>nx9369, A0=>que_out_27_0_6, A1=>nx9928, B0=>
      que_out_4_0_6, B1=>nx9902);
   ix9372 : aoi22 port map ( Y=>nx9371, A0=>que_out_0_0_6, A1=>nx9850, B0=>
      que_out_2_0_6, B1=>nx9876);
   ix7859 : nand03 port map ( Y=>nx7858, A0=>nx9374, A1=>nx9376, A2=>nx9378
   );
   ix9375 : aoi222 port map ( Y=>nx9374, A0=>que_out_26_0_6, A1=>nx9824, B0
      =>que_out_14_0_6, B1=>nx9798, C0=>que_out_11_0_6, C1=>nx9772);
   ix9377 : aoi22 port map ( Y=>nx9376, A0=>que_out_13_0_6, A1=>nx9746, B0=>
      que_out_7_0_6, B1=>nx9720);
   ix9379 : aoi22 port map ( Y=>nx9378, A0=>que_out_12_0_6, A1=>nx9694, B0=>
      que_out_1_0_6, B1=>nx9668);
   ix8053 : or04 port map ( Y=>out_column_0_7, A0=>nx8048, A1=>nx8022, A2=>
      nx7994, A3=>nx7968);
   ix8049 : nand03 port map ( Y=>nx8048, A0=>nx9382, A1=>nx9384, A2=>nx9386
   );
   ix9383 : aoi222 port map ( Y=>nx9382, A0=>que_out_10_0_7, A1=>nx10318, B0
      =>que_out_6_0_7, B1=>nx10370, C0=>que_out_9_0_7, C1=>nx10344);
   ix9385 : aoi22 port map ( Y=>nx9384, A0=>que_out_5_0_7, A1=>nx10266, B0=>
      que_out_18_0_7, B1=>nx10292);
   ix9387 : aoi22 port map ( Y=>nx9386, A0=>que_out_17_0_7, A1=>nx10240, B0
      =>que_out_20_0_7, B1=>nx10214);
   ix8023 : nand03 port map ( Y=>nx8022, A0=>nx9389, A1=>nx9391, A2=>nx9393
   );
   ix9390 : aoi222 port map ( Y=>nx9389, A0=>que_out_19_0_7, A1=>nx10188, B0
      =>que_out_21_0_7, B1=>nx10162, C0=>que_out_8_0_7, C1=>nx10136);
   ix9392 : aoi22 port map ( Y=>nx9391, A0=>que_out_25_0_7, A1=>nx10084, B0
      =>que_out_16_0_7, B1=>nx10110);
   ix9394 : aoi22 port map ( Y=>nx9393, A0=>que_out_24_0_7, A1=>nx10058, B0
      =>que_out_22_0_7, B1=>nx10032);
   ix7995 : nand03 port map ( Y=>nx7994, A0=>nx9396, A1=>nx9398, A2=>nx9400
   );
   ix9397 : aoi222 port map ( Y=>nx9396, A0=>que_out_15_0_7, A1=>nx9980, B0
      =>que_out_3_0_7, B1=>nx10006, C0=>que_out_23_0_7, C1=>nx9954);
   ix9399 : aoi22 port map ( Y=>nx9398, A0=>que_out_27_0_7, A1=>nx9928, B0=>
      que_out_4_0_7, B1=>nx9902);
   ix9401 : aoi22 port map ( Y=>nx9400, A0=>que_out_0_0_7, A1=>nx9850, B0=>
      que_out_2_0_7, B1=>nx9876);
   ix7969 : nand03 port map ( Y=>nx7968, A0=>nx9403, A1=>nx9405, A2=>nx9407
   );
   ix9404 : aoi222 port map ( Y=>nx9403, A0=>que_out_26_0_7, A1=>nx9824, B0
      =>que_out_14_0_7, B1=>nx9798, C0=>que_out_11_0_7, C1=>nx9772);
   ix9406 : aoi22 port map ( Y=>nx9405, A0=>que_out_13_0_7, A1=>nx9746, B0=>
      que_out_7_0_7, B1=>nx9720);
   ix9408 : aoi22 port map ( Y=>nx9407, A0=>que_out_12_0_7, A1=>nx9694, B0=>
      que_out_1_0_7, B1=>nx9668);
   ix8163 : or04 port map ( Y=>out_column_0_8, A0=>nx8158, A1=>nx8132, A2=>
      nx8104, A3=>nx8078);
   ix8159 : nand03 port map ( Y=>nx8158, A0=>nx9411, A1=>nx9413, A2=>nx9415
   );
   ix9412 : aoi222 port map ( Y=>nx9411, A0=>que_out_10_0_8, A1=>nx10318, B0
      =>que_out_6_0_8, B1=>nx10370, C0=>que_out_9_0_8, C1=>nx10344);
   ix9414 : aoi22 port map ( Y=>nx9413, A0=>que_out_5_0_8, A1=>nx10266, B0=>
      que_out_18_0_8, B1=>nx10292);
   ix9416 : aoi22 port map ( Y=>nx9415, A0=>que_out_17_0_8, A1=>nx10240, B0
      =>que_out_20_0_8, B1=>nx10214);
   ix8133 : nand03 port map ( Y=>nx8132, A0=>nx9418, A1=>nx9420, A2=>nx9422
   );
   ix9419 : aoi222 port map ( Y=>nx9418, A0=>que_out_19_0_8, A1=>nx10188, B0
      =>que_out_21_0_8, B1=>nx10162, C0=>que_out_8_0_8, C1=>nx10136);
   ix9421 : aoi22 port map ( Y=>nx9420, A0=>que_out_25_0_8, A1=>nx10084, B0
      =>que_out_16_0_8, B1=>nx10110);
   ix9423 : aoi22 port map ( Y=>nx9422, A0=>que_out_24_0_8, A1=>nx10058, B0
      =>que_out_22_0_8, B1=>nx10032);
   ix8105 : nand03 port map ( Y=>nx8104, A0=>nx9425, A1=>nx9427, A2=>nx9429
   );
   ix9426 : aoi222 port map ( Y=>nx9425, A0=>que_out_15_0_8, A1=>nx9980, B0
      =>que_out_3_0_8, B1=>nx10006, C0=>que_out_23_0_8, C1=>nx9954);
   ix9428 : aoi22 port map ( Y=>nx9427, A0=>que_out_27_0_8, A1=>nx9928, B0=>
      que_out_4_0_8, B1=>nx9902);
   ix9430 : aoi22 port map ( Y=>nx9429, A0=>que_out_0_0_8, A1=>nx9850, B0=>
      que_out_2_0_8, B1=>nx9876);
   ix8079 : nand03 port map ( Y=>nx8078, A0=>nx9432, A1=>nx9434, A2=>nx9436
   );
   ix9433 : aoi222 port map ( Y=>nx9432, A0=>que_out_26_0_8, A1=>nx9824, B0
      =>que_out_14_0_8, B1=>nx9798, C0=>que_out_11_0_8, C1=>nx9772);
   ix9435 : aoi22 port map ( Y=>nx9434, A0=>que_out_13_0_8, A1=>nx9746, B0=>
      que_out_7_0_8, B1=>nx9720);
   ix9437 : aoi22 port map ( Y=>nx9436, A0=>que_out_12_0_8, A1=>nx9694, B0=>
      que_out_1_0_8, B1=>nx9668);
   ix8273 : or04 port map ( Y=>out_column_0_9, A0=>nx8268, A1=>nx8242, A2=>
      nx8214, A3=>nx8188);
   ix8269 : nand03 port map ( Y=>nx8268, A0=>nx9440, A1=>nx9442, A2=>nx9444
   );
   ix9441 : aoi222 port map ( Y=>nx9440, A0=>que_out_10_0_9, A1=>nx10318, B0
      =>que_out_6_0_9, B1=>nx10370, C0=>que_out_9_0_9, C1=>nx10344);
   ix9443 : aoi22 port map ( Y=>nx9442, A0=>que_out_5_0_9, A1=>nx10266, B0=>
      que_out_18_0_9, B1=>nx10292);
   ix9445 : aoi22 port map ( Y=>nx9444, A0=>que_out_17_0_9, A1=>nx10240, B0
      =>que_out_20_0_9, B1=>nx10214);
   ix8243 : nand03 port map ( Y=>nx8242, A0=>nx9447, A1=>nx9449, A2=>nx9451
   );
   ix9448 : aoi222 port map ( Y=>nx9447, A0=>que_out_19_0_9, A1=>nx10188, B0
      =>que_out_21_0_9, B1=>nx10162, C0=>que_out_8_0_9, C1=>nx10136);
   ix9450 : aoi22 port map ( Y=>nx9449, A0=>que_out_25_0_9, A1=>nx10084, B0
      =>que_out_16_0_9, B1=>nx10110);
   ix9452 : aoi22 port map ( Y=>nx9451, A0=>que_out_24_0_9, A1=>nx10058, B0
      =>que_out_22_0_9, B1=>nx10032);
   ix8215 : nand03 port map ( Y=>nx8214, A0=>nx9454, A1=>nx9456, A2=>nx9458
   );
   ix9455 : aoi222 port map ( Y=>nx9454, A0=>que_out_15_0_9, A1=>nx9980, B0
      =>que_out_3_0_9, B1=>nx10006, C0=>que_out_23_0_9, C1=>nx9954);
   ix9457 : aoi22 port map ( Y=>nx9456, A0=>que_out_27_0_9, A1=>nx9928, B0=>
      que_out_4_0_9, B1=>nx9902);
   ix9459 : aoi22 port map ( Y=>nx9458, A0=>que_out_0_0_9, A1=>nx9850, B0=>
      que_out_2_0_9, B1=>nx9876);
   ix8189 : nand03 port map ( Y=>nx8188, A0=>nx9461, A1=>nx9463, A2=>nx9465
   );
   ix9462 : aoi222 port map ( Y=>nx9461, A0=>que_out_26_0_9, A1=>nx9824, B0
      =>que_out_14_0_9, B1=>nx9798, C0=>que_out_11_0_9, C1=>nx9772);
   ix9464 : aoi22 port map ( Y=>nx9463, A0=>que_out_13_0_9, A1=>nx9746, B0=>
      que_out_7_0_9, B1=>nx9720);
   ix9466 : aoi22 port map ( Y=>nx9465, A0=>que_out_12_0_9, A1=>nx9694, B0=>
      que_out_1_0_9, B1=>nx9668);
   ix8383 : or04 port map ( Y=>out_column_0_10, A0=>nx8378, A1=>nx8352, A2=>
      nx8324, A3=>nx8298);
   ix8379 : nand03 port map ( Y=>nx8378, A0=>nx9469, A1=>nx9471, A2=>nx9473
   );
   ix9470 : aoi222 port map ( Y=>nx9469, A0=>que_out_10_0_10, A1=>nx10318, 
      B0=>que_out_6_0_10, B1=>nx10370, C0=>que_out_9_0_10, C1=>nx10344);
   ix9472 : aoi22 port map ( Y=>nx9471, A0=>que_out_5_0_10, A1=>nx10266, B0
      =>que_out_18_0_10, B1=>nx10292);
   ix9474 : aoi22 port map ( Y=>nx9473, A0=>que_out_17_0_10, A1=>nx10240, B0
      =>que_out_20_0_10, B1=>nx10214);
   ix8353 : nand03 port map ( Y=>nx8352, A0=>nx9476, A1=>nx9478, A2=>nx9480
   );
   ix9477 : aoi222 port map ( Y=>nx9476, A0=>que_out_19_0_10, A1=>nx10188, 
      B0=>que_out_21_0_10, B1=>nx10162, C0=>que_out_8_0_10, C1=>nx10136);
   ix9479 : aoi22 port map ( Y=>nx9478, A0=>que_out_25_0_10, A1=>nx10084, B0
      =>que_out_16_0_10, B1=>nx10110);
   ix9481 : aoi22 port map ( Y=>nx9480, A0=>que_out_24_0_10, A1=>nx10058, B0
      =>que_out_22_0_10, B1=>nx10032);
   ix8325 : nand03 port map ( Y=>nx8324, A0=>nx9483, A1=>nx9485, A2=>nx9487
   );
   ix9484 : aoi222 port map ( Y=>nx9483, A0=>que_out_15_0_10, A1=>nx9980, B0
      =>que_out_3_0_10, B1=>nx10006, C0=>que_out_23_0_10, C1=>nx9954);
   ix9486 : aoi22 port map ( Y=>nx9485, A0=>que_out_27_0_10, A1=>nx9928, B0
      =>que_out_4_0_10, B1=>nx9902);
   ix9488 : aoi22 port map ( Y=>nx9487, A0=>que_out_0_0_10, A1=>nx9850, B0=>
      que_out_2_0_10, B1=>nx9876);
   ix8299 : nand03 port map ( Y=>nx8298, A0=>nx9490, A1=>nx9492, A2=>nx9494
   );
   ix9491 : aoi222 port map ( Y=>nx9490, A0=>que_out_26_0_10, A1=>nx9824, B0
      =>que_out_14_0_10, B1=>nx9798, C0=>que_out_11_0_10, C1=>nx9772);
   ix9493 : aoi22 port map ( Y=>nx9492, A0=>que_out_13_0_10, A1=>nx9746, B0
      =>que_out_7_0_10, B1=>nx9720);
   ix9495 : aoi22 port map ( Y=>nx9494, A0=>que_out_12_0_10, A1=>nx9694, B0
      =>que_out_1_0_10, B1=>nx9668);
   ix8493 : or04 port map ( Y=>out_column_0_11, A0=>nx8488, A1=>nx8462, A2=>
      nx8434, A3=>nx8408);
   ix8489 : nand03 port map ( Y=>nx8488, A0=>nx9498, A1=>nx9500, A2=>nx9502
   );
   ix9499 : aoi222 port map ( Y=>nx9498, A0=>que_out_10_0_11, A1=>nx10318, 
      B0=>que_out_6_0_11, B1=>nx10370, C0=>que_out_9_0_11, C1=>nx10344);
   ix9501 : aoi22 port map ( Y=>nx9500, A0=>que_out_5_0_11, A1=>nx10266, B0
      =>que_out_18_0_11, B1=>nx10292);
   ix9503 : aoi22 port map ( Y=>nx9502, A0=>que_out_17_0_11, A1=>nx10240, B0
      =>que_out_20_0_11, B1=>nx10214);
   ix8463 : nand03 port map ( Y=>nx8462, A0=>nx9505, A1=>nx9507, A2=>nx9509
   );
   ix9506 : aoi222 port map ( Y=>nx9505, A0=>que_out_19_0_11, A1=>nx10188, 
      B0=>que_out_21_0_11, B1=>nx10162, C0=>que_out_8_0_11, C1=>nx10136);
   ix9508 : aoi22 port map ( Y=>nx9507, A0=>que_out_25_0_11, A1=>nx10084, B0
      =>que_out_16_0_11, B1=>nx10110);
   ix9510 : aoi22 port map ( Y=>nx9509, A0=>que_out_24_0_11, A1=>nx10058, B0
      =>que_out_22_0_11, B1=>nx10032);
   ix8435 : nand03 port map ( Y=>nx8434, A0=>nx9512, A1=>nx9514, A2=>nx9516
   );
   ix9513 : aoi222 port map ( Y=>nx9512, A0=>que_out_15_0_11, A1=>nx9980, B0
      =>que_out_3_0_11, B1=>nx10006, C0=>que_out_23_0_11, C1=>nx9954);
   ix9515 : aoi22 port map ( Y=>nx9514, A0=>que_out_27_0_11, A1=>nx9928, B0
      =>que_out_4_0_11, B1=>nx9902);
   ix9517 : aoi22 port map ( Y=>nx9516, A0=>que_out_0_0_11, A1=>nx9850, B0=>
      que_out_2_0_11, B1=>nx9876);
   ix8409 : nand03 port map ( Y=>nx8408, A0=>nx9519, A1=>nx9521, A2=>nx9523
   );
   ix9520 : aoi222 port map ( Y=>nx9519, A0=>que_out_26_0_11, A1=>nx9824, B0
      =>que_out_14_0_11, B1=>nx9798, C0=>que_out_11_0_11, C1=>nx9772);
   ix9522 : aoi22 port map ( Y=>nx9521, A0=>que_out_13_0_11, A1=>nx9746, B0
      =>que_out_7_0_11, B1=>nx9720);
   ix9524 : aoi22 port map ( Y=>nx9523, A0=>que_out_12_0_11, A1=>nx9694, B0
      =>que_out_1_0_11, B1=>nx9668);
   ix8603 : or04 port map ( Y=>out_column_0_12, A0=>nx8598, A1=>nx8572, A2=>
      nx8544, A3=>nx8518);
   ix8599 : nand03 port map ( Y=>nx8598, A0=>nx9527, A1=>nx9529, A2=>nx9531
   );
   ix9528 : aoi222 port map ( Y=>nx9527, A0=>que_out_10_0_12, A1=>nx10318, 
      B0=>que_out_6_0_12, B1=>nx10370, C0=>que_out_9_0_12, C1=>nx10344);
   ix9530 : aoi22 port map ( Y=>nx9529, A0=>que_out_5_0_12, A1=>nx10266, B0
      =>que_out_18_0_12, B1=>nx10292);
   ix9532 : aoi22 port map ( Y=>nx9531, A0=>que_out_17_0_12, A1=>nx10240, B0
      =>que_out_20_0_12, B1=>nx10214);
   ix8573 : nand03 port map ( Y=>nx8572, A0=>nx9534, A1=>nx9536, A2=>nx9538
   );
   ix9535 : aoi222 port map ( Y=>nx9534, A0=>que_out_19_0_12, A1=>nx10188, 
      B0=>que_out_21_0_12, B1=>nx10162, C0=>que_out_8_0_12, C1=>nx10136);
   ix9537 : aoi22 port map ( Y=>nx9536, A0=>que_out_25_0_12, A1=>nx10084, B0
      =>que_out_16_0_12, B1=>nx10110);
   ix9539 : aoi22 port map ( Y=>nx9538, A0=>que_out_24_0_12, A1=>nx10058, B0
      =>que_out_22_0_12, B1=>nx10032);
   ix8545 : nand03 port map ( Y=>nx8544, A0=>nx9541, A1=>nx9543, A2=>nx9545
   );
   ix9542 : aoi222 port map ( Y=>nx9541, A0=>que_out_15_0_12, A1=>nx9980, B0
      =>que_out_3_0_12, B1=>nx10006, C0=>que_out_23_0_12, C1=>nx9954);
   ix9544 : aoi22 port map ( Y=>nx9543, A0=>que_out_27_0_12, A1=>nx9928, B0
      =>que_out_4_0_12, B1=>nx9902);
   ix9546 : aoi22 port map ( Y=>nx9545, A0=>que_out_0_0_12, A1=>nx9850, B0=>
      que_out_2_0_12, B1=>nx9876);
   ix8519 : nand03 port map ( Y=>nx8518, A0=>nx9548, A1=>nx9550, A2=>nx9552
   );
   ix9549 : aoi222 port map ( Y=>nx9548, A0=>que_out_26_0_12, A1=>nx9824, B0
      =>que_out_14_0_12, B1=>nx9798, C0=>que_out_11_0_12, C1=>nx9772);
   ix9551 : aoi22 port map ( Y=>nx9550, A0=>que_out_13_0_12, A1=>nx9746, B0
      =>que_out_7_0_12, B1=>nx9720);
   ix9553 : aoi22 port map ( Y=>nx9552, A0=>que_out_12_0_12, A1=>nx9694, B0
      =>que_out_1_0_12, B1=>nx9668);
   ix8713 : or04 port map ( Y=>out_column_0_13, A0=>nx8708, A1=>nx8682, A2=>
      nx8654, A3=>nx8628);
   ix8709 : nand03 port map ( Y=>nx8708, A0=>nx9556, A1=>nx9558, A2=>nx9560
   );
   ix9557 : aoi222 port map ( Y=>nx9556, A0=>que_out_10_0_13, A1=>nx10320, 
      B0=>que_out_6_0_13, B1=>nx10372, C0=>que_out_9_0_13, C1=>nx10346);
   ix9559 : aoi22 port map ( Y=>nx9558, A0=>que_out_5_0_13, A1=>nx10268, B0
      =>que_out_18_0_13, B1=>nx10294);
   ix9561 : aoi22 port map ( Y=>nx9560, A0=>que_out_17_0_13, A1=>nx10242, B0
      =>que_out_20_0_13, B1=>nx10216);
   ix8683 : nand03 port map ( Y=>nx8682, A0=>nx9563, A1=>nx9565, A2=>nx9567
   );
   ix9564 : aoi222 port map ( Y=>nx9563, A0=>que_out_19_0_13, A1=>nx10190, 
      B0=>que_out_21_0_13, B1=>nx10164, C0=>que_out_8_0_13, C1=>nx10138);
   ix9566 : aoi22 port map ( Y=>nx9565, A0=>que_out_25_0_13, A1=>nx10086, B0
      =>que_out_16_0_13, B1=>nx10112);
   ix9568 : aoi22 port map ( Y=>nx9567, A0=>que_out_24_0_13, A1=>nx10060, B0
      =>que_out_22_0_13, B1=>nx10034);
   ix8655 : nand03 port map ( Y=>nx8654, A0=>nx9570, A1=>nx9572, A2=>nx9574
   );
   ix9571 : aoi222 port map ( Y=>nx9570, A0=>que_out_15_0_13, A1=>nx9982, B0
      =>que_out_3_0_13, B1=>nx10008, C0=>que_out_23_0_13, C1=>nx9956);
   ix9573 : aoi22 port map ( Y=>nx9572, A0=>que_out_27_0_13, A1=>nx9930, B0
      =>que_out_4_0_13, B1=>nx9904);
   ix9575 : aoi22 port map ( Y=>nx9574, A0=>que_out_0_0_13, A1=>nx9852, B0=>
      que_out_2_0_13, B1=>nx9878);
   ix8629 : nand03 port map ( Y=>nx8628, A0=>nx9577, A1=>nx9579, A2=>nx9581
   );
   ix9578 : aoi222 port map ( Y=>nx9577, A0=>que_out_26_0_13, A1=>nx9826, B0
      =>que_out_14_0_13, B1=>nx9800, C0=>que_out_11_0_13, C1=>nx9774);
   ix9580 : aoi22 port map ( Y=>nx9579, A0=>que_out_13_0_13, A1=>nx9748, B0
      =>que_out_7_0_13, B1=>nx9722);
   ix9582 : aoi22 port map ( Y=>nx9581, A0=>que_out_12_0_13, A1=>nx9696, B0
      =>que_out_1_0_13, B1=>nx9670);
   ix8823 : or04 port map ( Y=>out_column_0_14, A0=>nx8818, A1=>nx8792, A2=>
      nx8764, A3=>nx8738);
   ix8819 : nand03 port map ( Y=>nx8818, A0=>nx9585, A1=>nx9587, A2=>nx9589
   );
   ix9586 : aoi222 port map ( Y=>nx9585, A0=>que_out_10_0_14, A1=>nx10320, 
      B0=>que_out_6_0_14, B1=>nx10372, C0=>que_out_9_0_14, C1=>nx10346);
   ix9588 : aoi22 port map ( Y=>nx9587, A0=>que_out_5_0_14, A1=>nx10268, B0
      =>que_out_18_0_14, B1=>nx10294);
   ix9590 : aoi22 port map ( Y=>nx9589, A0=>que_out_17_0_14, A1=>nx10242, B0
      =>que_out_20_0_14, B1=>nx10216);
   ix8793 : nand03 port map ( Y=>nx8792, A0=>nx9592, A1=>nx9594, A2=>nx9596
   );
   ix9593 : aoi222 port map ( Y=>nx9592, A0=>que_out_19_0_14, A1=>nx10190, 
      B0=>que_out_21_0_14, B1=>nx10164, C0=>que_out_8_0_14, C1=>nx10138);
   ix9595 : aoi22 port map ( Y=>nx9594, A0=>que_out_25_0_14, A1=>nx10086, B0
      =>que_out_16_0_14, B1=>nx10112);
   ix9597 : aoi22 port map ( Y=>nx9596, A0=>que_out_24_0_14, A1=>nx10060, B0
      =>que_out_22_0_14, B1=>nx10034);
   ix8765 : nand03 port map ( Y=>nx8764, A0=>nx9599, A1=>nx9601, A2=>nx9603
   );
   ix9600 : aoi222 port map ( Y=>nx9599, A0=>que_out_15_0_14, A1=>nx9982, B0
      =>que_out_3_0_14, B1=>nx10008, C0=>que_out_23_0_14, C1=>nx9956);
   ix9602 : aoi22 port map ( Y=>nx9601, A0=>que_out_27_0_14, A1=>nx9930, B0
      =>que_out_4_0_14, B1=>nx9904);
   ix9604 : aoi22 port map ( Y=>nx9603, A0=>que_out_0_0_14, A1=>nx9852, B0=>
      que_out_2_0_14, B1=>nx9878);
   ix8739 : nand03 port map ( Y=>nx8738, A0=>nx9606, A1=>nx9608, A2=>nx9610
   );
   ix9607 : aoi222 port map ( Y=>nx9606, A0=>que_out_26_0_14, A1=>nx9826, B0
      =>que_out_14_0_14, B1=>nx9800, C0=>que_out_11_0_14, C1=>nx9774);
   ix9609 : aoi22 port map ( Y=>nx9608, A0=>que_out_13_0_14, A1=>nx9748, B0
      =>que_out_7_0_14, B1=>nx9722);
   ix9611 : aoi22 port map ( Y=>nx9610, A0=>que_out_12_0_14, A1=>nx9696, B0
      =>que_out_1_0_14, B1=>nx9670);
   ix8933 : or04 port map ( Y=>out_column_0_15, A0=>nx8928, A1=>nx8902, A2=>
      nx8874, A3=>nx8848);
   ix8929 : nand03 port map ( Y=>nx8928, A0=>nx9614, A1=>nx9616, A2=>nx9618
   );
   ix9615 : aoi222 port map ( Y=>nx9614, A0=>que_out_10_0_15, A1=>nx10320, 
      B0=>que_out_6_0_15, B1=>nx10372, C0=>que_out_9_0_15, C1=>nx10346);
   ix9617 : aoi22 port map ( Y=>nx9616, A0=>que_out_5_0_15, A1=>nx10268, B0
      =>que_out_18_0_15, B1=>nx10294);
   ix9619 : aoi22 port map ( Y=>nx9618, A0=>que_out_17_0_15, A1=>nx10242, B0
      =>que_out_20_0_15, B1=>nx10216);
   ix8903 : nand03 port map ( Y=>nx8902, A0=>nx9621, A1=>nx9623, A2=>nx9625
   );
   ix9622 : aoi222 port map ( Y=>nx9621, A0=>que_out_19_0_15, A1=>nx10190, 
      B0=>que_out_21_0_15, B1=>nx10164, C0=>que_out_8_0_15, C1=>nx10138);
   ix9624 : aoi22 port map ( Y=>nx9623, A0=>que_out_25_0_15, A1=>nx10086, B0
      =>que_out_16_0_15, B1=>nx10112);
   ix9626 : aoi22 port map ( Y=>nx9625, A0=>que_out_24_0_15, A1=>nx10060, B0
      =>que_out_22_0_15, B1=>nx10034);
   ix8875 : nand03 port map ( Y=>nx8874, A0=>nx9628, A1=>nx9630, A2=>nx9632
   );
   ix9629 : aoi222 port map ( Y=>nx9628, A0=>que_out_15_0_15, A1=>nx9982, B0
      =>que_out_3_0_15, B1=>nx10008, C0=>que_out_23_0_15, C1=>nx9956);
   ix9631 : aoi22 port map ( Y=>nx9630, A0=>que_out_27_0_15, A1=>nx9930, B0
      =>que_out_4_0_15, B1=>nx9904);
   ix9633 : aoi22 port map ( Y=>nx9632, A0=>que_out_0_0_15, A1=>nx9852, B0=>
      que_out_2_0_15, B1=>nx9878);
   ix8849 : nand03 port map ( Y=>nx8848, A0=>nx9635, A1=>nx9637, A2=>nx9639
   );
   ix9636 : aoi222 port map ( Y=>nx9635, A0=>que_out_26_0_15, A1=>nx9826, B0
      =>que_out_14_0_15, B1=>nx9800, C0=>que_out_11_0_15, C1=>nx9774);
   ix9638 : aoi22 port map ( Y=>nx9637, A0=>que_out_13_0_15, A1=>nx9748, B0
      =>que_out_7_0_15, B1=>nx9722);
   ix9640 : aoi22 port map ( Y=>nx9639, A0=>que_out_12_0_15, A1=>nx9696, B0
      =>que_out_1_0_15, B1=>nx9670);
   ix6944 : inv02 port map ( Y=>nx6943, A=>nx88);
   ix9647 : inv02 port map ( Y=>nx9648, A=>nx10378);
   ix9649 : inv02 port map ( Y=>nx9650, A=>nx10378);
   ix9651 : inv02 port map ( Y=>nx9652, A=>nx10378);
   ix9653 : inv02 port map ( Y=>nx9654, A=>nx10378);
   ix9655 : inv02 port map ( Y=>nx9656, A=>nx10378);
   ix9657 : inv02 port map ( Y=>nx9658, A=>nx10378);
   ix9659 : inv02 port map ( Y=>nx9660, A=>nx10378);
   ix9661 : inv02 port map ( Y=>nx9662, A=>nx10380);
   ix9663 : inv02 port map ( Y=>nx9664, A=>nx10380);
   ix9665 : inv02 port map ( Y=>nx9666, A=>nx10380);
   ix9667 : inv02 port map ( Y=>nx9668, A=>nx10380);
   ix9669 : inv02 port map ( Y=>nx9670, A=>nx10380);
   ix9673 : inv02 port map ( Y=>nx9674, A=>nx10382);
   ix9675 : inv02 port map ( Y=>nx9676, A=>nx10382);
   ix9677 : inv02 port map ( Y=>nx9678, A=>nx10382);
   ix9679 : inv02 port map ( Y=>nx9680, A=>nx10382);
   ix9681 : inv02 port map ( Y=>nx9682, A=>nx10382);
   ix9683 : inv02 port map ( Y=>nx9684, A=>nx10382);
   ix9685 : inv02 port map ( Y=>nx9686, A=>nx10382);
   ix9687 : inv02 port map ( Y=>nx9688, A=>nx10384);
   ix9689 : inv02 port map ( Y=>nx9690, A=>nx10384);
   ix9691 : inv02 port map ( Y=>nx9692, A=>nx10384);
   ix9693 : inv02 port map ( Y=>nx9694, A=>nx10384);
   ix9695 : inv02 port map ( Y=>nx9696, A=>nx10384);
   ix9699 : inv02 port map ( Y=>nx9700, A=>nx10386);
   ix9701 : inv02 port map ( Y=>nx9702, A=>nx10386);
   ix9703 : inv02 port map ( Y=>nx9704, A=>nx10386);
   ix9705 : inv02 port map ( Y=>nx9706, A=>nx10386);
   ix9707 : inv02 port map ( Y=>nx9708, A=>nx10386);
   ix9709 : inv02 port map ( Y=>nx9710, A=>nx10386);
   ix9711 : inv02 port map ( Y=>nx9712, A=>nx10386);
   ix9713 : inv02 port map ( Y=>nx9714, A=>nx10388);
   ix9715 : inv02 port map ( Y=>nx9716, A=>nx10388);
   ix9717 : inv02 port map ( Y=>nx9718, A=>nx10388);
   ix9719 : inv02 port map ( Y=>nx9720, A=>nx10388);
   ix9721 : inv02 port map ( Y=>nx9722, A=>nx10388);
   ix9725 : inv02 port map ( Y=>nx9726, A=>nx10390);
   ix9727 : inv02 port map ( Y=>nx9728, A=>nx10390);
   ix9729 : inv02 port map ( Y=>nx9730, A=>nx10390);
   ix9731 : inv02 port map ( Y=>nx9732, A=>nx10390);
   ix9733 : inv02 port map ( Y=>nx9734, A=>nx10390);
   ix9735 : inv02 port map ( Y=>nx9736, A=>nx10390);
   ix9737 : inv02 port map ( Y=>nx9738, A=>nx10390);
   ix9739 : inv02 port map ( Y=>nx9740, A=>nx10392);
   ix9741 : inv02 port map ( Y=>nx9742, A=>nx10392);
   ix9743 : inv02 port map ( Y=>nx9744, A=>nx10392);
   ix9745 : inv02 port map ( Y=>nx9746, A=>nx10392);
   ix9747 : inv02 port map ( Y=>nx9748, A=>nx10392);
   ix9751 : inv02 port map ( Y=>nx9752, A=>nx10394);
   ix9753 : inv02 port map ( Y=>nx9754, A=>nx10394);
   ix9755 : inv02 port map ( Y=>nx9756, A=>nx10394);
   ix9757 : inv02 port map ( Y=>nx9758, A=>nx10394);
   ix9759 : inv02 port map ( Y=>nx9760, A=>nx10394);
   ix9761 : inv02 port map ( Y=>nx9762, A=>nx10394);
   ix9763 : inv02 port map ( Y=>nx9764, A=>nx10394);
   ix9765 : inv02 port map ( Y=>nx9766, A=>nx10396);
   ix9767 : inv02 port map ( Y=>nx9768, A=>nx10396);
   ix9769 : inv02 port map ( Y=>nx9770, A=>nx10396);
   ix9771 : inv02 port map ( Y=>nx9772, A=>nx10396);
   ix9773 : inv02 port map ( Y=>nx9774, A=>nx10396);
   ix9777 : inv02 port map ( Y=>nx9778, A=>nx10398);
   ix9779 : inv02 port map ( Y=>nx9780, A=>nx10398);
   ix9781 : inv02 port map ( Y=>nx9782, A=>nx10398);
   ix9783 : inv02 port map ( Y=>nx9784, A=>nx10398);
   ix9785 : inv02 port map ( Y=>nx9786, A=>nx10398);
   ix9787 : inv02 port map ( Y=>nx9788, A=>nx10398);
   ix9789 : inv02 port map ( Y=>nx9790, A=>nx10398);
   ix9791 : inv02 port map ( Y=>nx9792, A=>nx10400);
   ix9793 : inv02 port map ( Y=>nx9794, A=>nx10400);
   ix9795 : inv02 port map ( Y=>nx9796, A=>nx10400);
   ix9797 : inv02 port map ( Y=>nx9798, A=>nx10400);
   ix9799 : inv02 port map ( Y=>nx9800, A=>nx10400);
   ix9803 : inv02 port map ( Y=>nx9804, A=>nx10402);
   ix9805 : inv02 port map ( Y=>nx9806, A=>nx10402);
   ix9807 : inv02 port map ( Y=>nx9808, A=>nx10402);
   ix9809 : inv02 port map ( Y=>nx9810, A=>nx10402);
   ix9811 : inv02 port map ( Y=>nx9812, A=>nx10402);
   ix9813 : inv02 port map ( Y=>nx9814, A=>nx10402);
   ix9815 : inv02 port map ( Y=>nx9816, A=>nx10402);
   ix9817 : inv02 port map ( Y=>nx9818, A=>nx10404);
   ix9819 : inv02 port map ( Y=>nx9820, A=>nx10404);
   ix9821 : inv02 port map ( Y=>nx9822, A=>nx10404);
   ix9823 : inv02 port map ( Y=>nx9824, A=>nx10404);
   ix9825 : inv02 port map ( Y=>nx9826, A=>nx10404);
   ix9829 : inv02 port map ( Y=>nx9830, A=>nx10406);
   ix9831 : inv02 port map ( Y=>nx9832, A=>nx10406);
   ix9833 : inv02 port map ( Y=>nx9834, A=>nx10406);
   ix9835 : inv02 port map ( Y=>nx9836, A=>nx10406);
   ix9837 : inv02 port map ( Y=>nx9838, A=>nx10406);
   ix9839 : inv02 port map ( Y=>nx9840, A=>nx10406);
   ix9841 : inv02 port map ( Y=>nx9842, A=>nx10406);
   ix9843 : inv02 port map ( Y=>nx9844, A=>nx10408);
   ix9845 : inv02 port map ( Y=>nx9846, A=>nx10408);
   ix9847 : inv02 port map ( Y=>nx9848, A=>nx10408);
   ix9849 : inv02 port map ( Y=>nx9850, A=>nx10408);
   ix9851 : inv02 port map ( Y=>nx9852, A=>nx10408);
   ix9855 : inv02 port map ( Y=>nx9856, A=>nx10410);
   ix9857 : inv02 port map ( Y=>nx9858, A=>nx10410);
   ix9859 : inv02 port map ( Y=>nx9860, A=>nx10410);
   ix9861 : inv02 port map ( Y=>nx9862, A=>nx10410);
   ix9863 : inv02 port map ( Y=>nx9864, A=>nx10410);
   ix9865 : inv02 port map ( Y=>nx9866, A=>nx10410);
   ix9867 : inv02 port map ( Y=>nx9868, A=>nx10410);
   ix9869 : inv02 port map ( Y=>nx9870, A=>nx10412);
   ix9871 : inv02 port map ( Y=>nx9872, A=>nx10412);
   ix9873 : inv02 port map ( Y=>nx9874, A=>nx10412);
   ix9875 : inv02 port map ( Y=>nx9876, A=>nx10412);
   ix9877 : inv02 port map ( Y=>nx9878, A=>nx10412);
   ix9881 : inv02 port map ( Y=>nx9882, A=>nx10414);
   ix9883 : inv02 port map ( Y=>nx9884, A=>nx10414);
   ix9885 : inv02 port map ( Y=>nx9886, A=>nx10414);
   ix9887 : inv02 port map ( Y=>nx9888, A=>nx10414);
   ix9889 : inv02 port map ( Y=>nx9890, A=>nx10414);
   ix9891 : inv02 port map ( Y=>nx9892, A=>nx10414);
   ix9893 : inv02 port map ( Y=>nx9894, A=>nx10414);
   ix9895 : inv02 port map ( Y=>nx9896, A=>nx10416);
   ix9897 : inv02 port map ( Y=>nx9898, A=>nx10416);
   ix9899 : inv02 port map ( Y=>nx9900, A=>nx10416);
   ix9901 : inv02 port map ( Y=>nx9902, A=>nx10416);
   ix9903 : inv02 port map ( Y=>nx9904, A=>nx10416);
   ix9907 : inv02 port map ( Y=>nx9908, A=>nx10418);
   ix9909 : inv02 port map ( Y=>nx9910, A=>nx10418);
   ix9911 : inv02 port map ( Y=>nx9912, A=>nx10418);
   ix9913 : inv02 port map ( Y=>nx9914, A=>nx10418);
   ix9915 : inv02 port map ( Y=>nx9916, A=>nx10418);
   ix9917 : inv02 port map ( Y=>nx9918, A=>nx10418);
   ix9919 : inv02 port map ( Y=>nx9920, A=>nx10418);
   ix9921 : inv02 port map ( Y=>nx9922, A=>nx10420);
   ix9923 : inv02 port map ( Y=>nx9924, A=>nx10420);
   ix9925 : inv02 port map ( Y=>nx9926, A=>nx10420);
   ix9927 : inv02 port map ( Y=>nx9928, A=>nx10420);
   ix9929 : inv02 port map ( Y=>nx9930, A=>nx10420);
   ix9933 : inv02 port map ( Y=>nx9934, A=>nx10422);
   ix9935 : inv02 port map ( Y=>nx9936, A=>nx10422);
   ix9937 : inv02 port map ( Y=>nx9938, A=>nx10422);
   ix9939 : inv02 port map ( Y=>nx9940, A=>nx10422);
   ix9941 : inv02 port map ( Y=>nx9942, A=>nx10422);
   ix9943 : inv02 port map ( Y=>nx9944, A=>nx10422);
   ix9945 : inv02 port map ( Y=>nx9946, A=>nx10422);
   ix9947 : inv02 port map ( Y=>nx9948, A=>nx10424);
   ix9949 : inv02 port map ( Y=>nx9950, A=>nx10424);
   ix9951 : inv02 port map ( Y=>nx9952, A=>nx10424);
   ix9953 : inv02 port map ( Y=>nx9954, A=>nx10424);
   ix9955 : inv02 port map ( Y=>nx9956, A=>nx10424);
   ix9959 : inv02 port map ( Y=>nx9960, A=>nx10426);
   ix9961 : inv02 port map ( Y=>nx9962, A=>nx10426);
   ix9963 : inv02 port map ( Y=>nx9964, A=>nx10426);
   ix9965 : inv02 port map ( Y=>nx9966, A=>nx10426);
   ix9967 : inv02 port map ( Y=>nx9968, A=>nx10426);
   ix9969 : inv02 port map ( Y=>nx9970, A=>nx10426);
   ix9971 : inv02 port map ( Y=>nx9972, A=>nx10426);
   ix9973 : inv02 port map ( Y=>nx9974, A=>nx10428);
   ix9975 : inv02 port map ( Y=>nx9976, A=>nx10428);
   ix9977 : inv02 port map ( Y=>nx9978, A=>nx10428);
   ix9979 : inv02 port map ( Y=>nx9980, A=>nx10428);
   ix9981 : inv02 port map ( Y=>nx9982, A=>nx10428);
   ix9985 : inv02 port map ( Y=>nx9986, A=>nx10430);
   ix9987 : inv02 port map ( Y=>nx9988, A=>nx10430);
   ix9989 : inv02 port map ( Y=>nx9990, A=>nx10430);
   ix9991 : inv02 port map ( Y=>nx9992, A=>nx10430);
   ix9993 : inv02 port map ( Y=>nx9994, A=>nx10430);
   ix9995 : inv02 port map ( Y=>nx9996, A=>nx10430);
   ix9997 : inv02 port map ( Y=>nx9998, A=>nx10430);
   ix9999 : inv02 port map ( Y=>nx10000, A=>nx10432);
   ix10001 : inv02 port map ( Y=>nx10002, A=>nx10432);
   ix10003 : inv02 port map ( Y=>nx10004, A=>nx10432);
   ix10005 : inv02 port map ( Y=>nx10006, A=>nx10432);
   ix10007 : inv02 port map ( Y=>nx10008, A=>nx10432);
   ix10011 : inv02 port map ( Y=>nx10012, A=>nx10434);
   ix10013 : inv02 port map ( Y=>nx10014, A=>nx10434);
   ix10015 : inv02 port map ( Y=>nx10016, A=>nx10434);
   ix10017 : inv02 port map ( Y=>nx10018, A=>nx10434);
   ix10019 : inv02 port map ( Y=>nx10020, A=>nx10434);
   ix10021 : inv02 port map ( Y=>nx10022, A=>nx10434);
   ix10023 : inv02 port map ( Y=>nx10024, A=>nx10434);
   ix10025 : inv02 port map ( Y=>nx10026, A=>nx10436);
   ix10027 : inv02 port map ( Y=>nx10028, A=>nx10436);
   ix10029 : inv02 port map ( Y=>nx10030, A=>nx10436);
   ix10031 : inv02 port map ( Y=>nx10032, A=>nx10436);
   ix10033 : inv02 port map ( Y=>nx10034, A=>nx10436);
   ix10037 : inv02 port map ( Y=>nx10038, A=>nx10438);
   ix10039 : inv02 port map ( Y=>nx10040, A=>nx10438);
   ix10041 : inv02 port map ( Y=>nx10042, A=>nx10438);
   ix10043 : inv02 port map ( Y=>nx10044, A=>nx10438);
   ix10045 : inv02 port map ( Y=>nx10046, A=>nx10438);
   ix10047 : inv02 port map ( Y=>nx10048, A=>nx10438);
   ix10049 : inv02 port map ( Y=>nx10050, A=>nx10438);
   ix10051 : inv02 port map ( Y=>nx10052, A=>nx10440);
   ix10053 : inv02 port map ( Y=>nx10054, A=>nx10440);
   ix10055 : inv02 port map ( Y=>nx10056, A=>nx10440);
   ix10057 : inv02 port map ( Y=>nx10058, A=>nx10440);
   ix10059 : inv02 port map ( Y=>nx10060, A=>nx10440);
   ix10063 : inv02 port map ( Y=>nx10064, A=>nx10442);
   ix10065 : inv02 port map ( Y=>nx10066, A=>nx10442);
   ix10067 : inv02 port map ( Y=>nx10068, A=>nx10442);
   ix10069 : inv02 port map ( Y=>nx10070, A=>nx10442);
   ix10071 : inv02 port map ( Y=>nx10072, A=>nx10442);
   ix10073 : inv02 port map ( Y=>nx10074, A=>nx10442);
   ix10075 : inv02 port map ( Y=>nx10076, A=>nx10442);
   ix10077 : inv02 port map ( Y=>nx10078, A=>nx10444);
   ix10079 : inv02 port map ( Y=>nx10080, A=>nx10444);
   ix10081 : inv02 port map ( Y=>nx10082, A=>nx10444);
   ix10083 : inv02 port map ( Y=>nx10084, A=>nx10444);
   ix10085 : inv02 port map ( Y=>nx10086, A=>nx10444);
   ix10089 : inv02 port map ( Y=>nx10090, A=>nx10446);
   ix10091 : inv02 port map ( Y=>nx10092, A=>nx10446);
   ix10093 : inv02 port map ( Y=>nx10094, A=>nx10446);
   ix10095 : inv02 port map ( Y=>nx10096, A=>nx10446);
   ix10097 : inv02 port map ( Y=>nx10098, A=>nx10446);
   ix10099 : inv02 port map ( Y=>nx10100, A=>nx10446);
   ix10101 : inv02 port map ( Y=>nx10102, A=>nx10446);
   ix10103 : inv02 port map ( Y=>nx10104, A=>nx10448);
   ix10105 : inv02 port map ( Y=>nx10106, A=>nx10448);
   ix10107 : inv02 port map ( Y=>nx10108, A=>nx10448);
   ix10109 : inv02 port map ( Y=>nx10110, A=>nx10448);
   ix10111 : inv02 port map ( Y=>nx10112, A=>nx10448);
   ix10115 : inv02 port map ( Y=>nx10116, A=>nx10450);
   ix10117 : inv02 port map ( Y=>nx10118, A=>nx10450);
   ix10119 : inv02 port map ( Y=>nx10120, A=>nx10450);
   ix10121 : inv02 port map ( Y=>nx10122, A=>nx10450);
   ix10123 : inv02 port map ( Y=>nx10124, A=>nx10450);
   ix10125 : inv02 port map ( Y=>nx10126, A=>nx10450);
   ix10127 : inv02 port map ( Y=>nx10128, A=>nx10450);
   ix10129 : inv02 port map ( Y=>nx10130, A=>nx10452);
   ix10131 : inv02 port map ( Y=>nx10132, A=>nx10452);
   ix10133 : inv02 port map ( Y=>nx10134, A=>nx10452);
   ix10135 : inv02 port map ( Y=>nx10136, A=>nx10452);
   ix10137 : inv02 port map ( Y=>nx10138, A=>nx10452);
   ix10141 : inv02 port map ( Y=>nx10142, A=>nx10454);
   ix10143 : inv02 port map ( Y=>nx10144, A=>nx10454);
   ix10145 : inv02 port map ( Y=>nx10146, A=>nx10454);
   ix10147 : inv02 port map ( Y=>nx10148, A=>nx10454);
   ix10149 : inv02 port map ( Y=>nx10150, A=>nx10454);
   ix10151 : inv02 port map ( Y=>nx10152, A=>nx10454);
   ix10153 : inv02 port map ( Y=>nx10154, A=>nx10454);
   ix10155 : inv02 port map ( Y=>nx10156, A=>nx10456);
   ix10157 : inv02 port map ( Y=>nx10158, A=>nx10456);
   ix10159 : inv02 port map ( Y=>nx10160, A=>nx10456);
   ix10161 : inv02 port map ( Y=>nx10162, A=>nx10456);
   ix10163 : inv02 port map ( Y=>nx10164, A=>nx10456);
   ix10167 : inv02 port map ( Y=>nx10168, A=>nx10458);
   ix10169 : inv02 port map ( Y=>nx10170, A=>nx10458);
   ix10171 : inv02 port map ( Y=>nx10172, A=>nx10458);
   ix10173 : inv02 port map ( Y=>nx10174, A=>nx10458);
   ix10175 : inv02 port map ( Y=>nx10176, A=>nx10458);
   ix10177 : inv02 port map ( Y=>nx10178, A=>nx10458);
   ix10179 : inv02 port map ( Y=>nx10180, A=>nx10458);
   ix10181 : inv02 port map ( Y=>nx10182, A=>nx10460);
   ix10183 : inv02 port map ( Y=>nx10184, A=>nx10460);
   ix10185 : inv02 port map ( Y=>nx10186, A=>nx10460);
   ix10187 : inv02 port map ( Y=>nx10188, A=>nx10460);
   ix10189 : inv02 port map ( Y=>nx10190, A=>nx10460);
   ix10193 : inv02 port map ( Y=>nx10194, A=>nx10462);
   ix10195 : inv02 port map ( Y=>nx10196, A=>nx10462);
   ix10197 : inv02 port map ( Y=>nx10198, A=>nx10462);
   ix10199 : inv02 port map ( Y=>nx10200, A=>nx10462);
   ix10201 : inv02 port map ( Y=>nx10202, A=>nx10462);
   ix10203 : inv02 port map ( Y=>nx10204, A=>nx10462);
   ix10205 : inv02 port map ( Y=>nx10206, A=>nx10462);
   ix10207 : inv02 port map ( Y=>nx10208, A=>nx10464);
   ix10209 : inv02 port map ( Y=>nx10210, A=>nx10464);
   ix10211 : inv02 port map ( Y=>nx10212, A=>nx10464);
   ix10213 : inv02 port map ( Y=>nx10214, A=>nx10464);
   ix10215 : inv02 port map ( Y=>nx10216, A=>nx10464);
   ix10219 : inv02 port map ( Y=>nx10220, A=>nx10466);
   ix10221 : inv02 port map ( Y=>nx10222, A=>nx10466);
   ix10223 : inv02 port map ( Y=>nx10224, A=>nx10466);
   ix10225 : inv02 port map ( Y=>nx10226, A=>nx10466);
   ix10227 : inv02 port map ( Y=>nx10228, A=>nx10466);
   ix10229 : inv02 port map ( Y=>nx10230, A=>nx10466);
   ix10231 : inv02 port map ( Y=>nx10232, A=>nx10466);
   ix10233 : inv02 port map ( Y=>nx10234, A=>nx10468);
   ix10235 : inv02 port map ( Y=>nx10236, A=>nx10468);
   ix10237 : inv02 port map ( Y=>nx10238, A=>nx10468);
   ix10239 : inv02 port map ( Y=>nx10240, A=>nx10468);
   ix10241 : inv02 port map ( Y=>nx10242, A=>nx10468);
   ix10245 : inv02 port map ( Y=>nx10246, A=>nx10470);
   ix10247 : inv02 port map ( Y=>nx10248, A=>nx10470);
   ix10249 : inv02 port map ( Y=>nx10250, A=>nx10470);
   ix10251 : inv02 port map ( Y=>nx10252, A=>nx10470);
   ix10253 : inv02 port map ( Y=>nx10254, A=>nx10470);
   ix10255 : inv02 port map ( Y=>nx10256, A=>nx10470);
   ix10257 : inv02 port map ( Y=>nx10258, A=>nx10470);
   ix10259 : inv02 port map ( Y=>nx10260, A=>nx10472);
   ix10261 : inv02 port map ( Y=>nx10262, A=>nx10472);
   ix10263 : inv02 port map ( Y=>nx10264, A=>nx10472);
   ix10265 : inv02 port map ( Y=>nx10266, A=>nx10472);
   ix10267 : inv02 port map ( Y=>nx10268, A=>nx10472);
   ix10271 : inv02 port map ( Y=>nx10272, A=>nx10474);
   ix10273 : inv02 port map ( Y=>nx10274, A=>nx10474);
   ix10275 : inv02 port map ( Y=>nx10276, A=>nx10474);
   ix10277 : inv02 port map ( Y=>nx10278, A=>nx10474);
   ix10279 : inv02 port map ( Y=>nx10280, A=>nx10474);
   ix10281 : inv02 port map ( Y=>nx10282, A=>nx10474);
   ix10283 : inv02 port map ( Y=>nx10284, A=>nx10474);
   ix10285 : inv02 port map ( Y=>nx10286, A=>nx10476);
   ix10287 : inv02 port map ( Y=>nx10288, A=>nx10476);
   ix10289 : inv02 port map ( Y=>nx10290, A=>nx10476);
   ix10291 : inv02 port map ( Y=>nx10292, A=>nx10476);
   ix10293 : inv02 port map ( Y=>nx10294, A=>nx10476);
   ix10297 : inv02 port map ( Y=>nx10298, A=>nx10478);
   ix10299 : inv02 port map ( Y=>nx10300, A=>nx10478);
   ix10301 : inv02 port map ( Y=>nx10302, A=>nx10478);
   ix10303 : inv02 port map ( Y=>nx10304, A=>nx10478);
   ix10305 : inv02 port map ( Y=>nx10306, A=>nx10478);
   ix10307 : inv02 port map ( Y=>nx10308, A=>nx10478);
   ix10309 : inv02 port map ( Y=>nx10310, A=>nx10478);
   ix10311 : inv02 port map ( Y=>nx10312, A=>nx10480);
   ix10313 : inv02 port map ( Y=>nx10314, A=>nx10480);
   ix10315 : inv02 port map ( Y=>nx10316, A=>nx10480);
   ix10317 : inv02 port map ( Y=>nx10318, A=>nx10480);
   ix10319 : inv02 port map ( Y=>nx10320, A=>nx10480);
   ix10323 : inv02 port map ( Y=>nx10324, A=>nx10482);
   ix10325 : inv02 port map ( Y=>nx10326, A=>nx10482);
   ix10327 : inv02 port map ( Y=>nx10328, A=>nx10482);
   ix10329 : inv02 port map ( Y=>nx10330, A=>nx10482);
   ix10331 : inv02 port map ( Y=>nx10332, A=>nx10482);
   ix10333 : inv02 port map ( Y=>nx10334, A=>nx10482);
   ix10335 : inv02 port map ( Y=>nx10336, A=>nx10482);
   ix10337 : inv02 port map ( Y=>nx10338, A=>nx10484);
   ix10339 : inv02 port map ( Y=>nx10340, A=>nx10484);
   ix10341 : inv02 port map ( Y=>nx10342, A=>nx10484);
   ix10343 : inv02 port map ( Y=>nx10344, A=>nx10484);
   ix10345 : inv02 port map ( Y=>nx10346, A=>nx10484);
   ix10349 : inv02 port map ( Y=>nx10350, A=>nx10486);
   ix10351 : inv02 port map ( Y=>nx10352, A=>nx10486);
   ix10353 : inv02 port map ( Y=>nx10354, A=>nx10486);
   ix10355 : inv02 port map ( Y=>nx10356, A=>nx10486);
   ix10357 : inv02 port map ( Y=>nx10358, A=>nx10486);
   ix10359 : inv02 port map ( Y=>nx10360, A=>nx10486);
   ix10361 : inv02 port map ( Y=>nx10362, A=>nx10486);
   ix10363 : inv02 port map ( Y=>nx10364, A=>nx10488);
   ix10365 : inv02 port map ( Y=>nx10366, A=>nx10488);
   ix10367 : inv02 port map ( Y=>nx10368, A=>nx10488);
   ix10369 : inv02 port map ( Y=>nx10370, A=>nx10488);
   ix10371 : inv02 port map ( Y=>nx10372, A=>nx10488);
   ix10373 : buf02 port map ( Y=>nx10374, A=>nx6955);
   ix10375 : buf02 port map ( Y=>nx10376, A=>nx6955);
   ix10377 : inv02 port map ( Y=>nx10378, A=>nx14);
   ix10379 : inv02 port map ( Y=>nx10380, A=>nx14);
   ix10381 : inv02 port map ( Y=>nx10382, A=>nx30);
   ix10383 : inv02 port map ( Y=>nx10384, A=>nx30);
   ix10385 : inv02 port map ( Y=>nx10386, A=>nx42);
   ix10387 : inv02 port map ( Y=>nx10388, A=>nx42);
   ix10389 : inv02 port map ( Y=>nx10390, A=>nx48);
   ix10391 : inv02 port map ( Y=>nx10392, A=>nx48);
   ix10393 : inv02 port map ( Y=>nx10394, A=>nx64);
   ix10395 : inv02 port map ( Y=>nx10396, A=>nx64);
   ix10397 : inv02 port map ( Y=>nx10398, A=>nx68);
   ix10399 : inv02 port map ( Y=>nx10400, A=>nx68);
   ix10401 : inv02 port map ( Y=>nx10402, A=>nx74);
   ix10403 : inv02 port map ( Y=>nx10404, A=>nx74);
   ix10405 : inv02 port map ( Y=>nx10406, A=>nx90);
   ix10407 : inv02 port map ( Y=>nx10408, A=>nx90);
   ix10409 : inv02 port map ( Y=>nx10410, A=>nx94);
   ix10411 : inv02 port map ( Y=>nx10412, A=>nx94);
   ix10413 : inv02 port map ( Y=>nx10414, A=>nx100);
   ix10415 : inv02 port map ( Y=>nx10416, A=>nx100);
   ix10417 : inv02 port map ( Y=>nx10418, A=>nx104);
   ix10419 : inv02 port map ( Y=>nx10420, A=>nx104);
   ix10421 : inv02 port map ( Y=>nx10422, A=>nx114);
   ix10423 : inv02 port map ( Y=>nx10424, A=>nx114);
   ix10425 : inv02 port map ( Y=>nx10426, A=>nx118);
   ix10427 : inv02 port map ( Y=>nx10428, A=>nx118);
   ix10429 : inv02 port map ( Y=>nx10430, A=>nx122);
   ix10431 : inv02 port map ( Y=>nx10432, A=>nx122);
   ix10433 : inv02 port map ( Y=>nx10434, A=>nx136);
   ix10435 : inv02 port map ( Y=>nx10436, A=>nx136);
   ix10437 : inv02 port map ( Y=>nx10438, A=>nx144);
   ix10439 : inv02 port map ( Y=>nx10440, A=>nx144);
   ix10441 : inv02 port map ( Y=>nx10442, A=>nx150);
   ix10443 : inv02 port map ( Y=>nx10444, A=>nx150);
   ix10445 : inv02 port map ( Y=>nx10446, A=>nx158);
   ix10447 : inv02 port map ( Y=>nx10448, A=>nx158);
   ix10449 : inv02 port map ( Y=>nx10450, A=>nx166);
   ix10451 : inv02 port map ( Y=>nx10452, A=>nx166);
   ix10453 : inv02 port map ( Y=>nx10454, A=>nx172);
   ix10455 : inv02 port map ( Y=>nx10456, A=>nx172);
   ix10457 : inv02 port map ( Y=>nx10458, A=>nx180);
   ix10459 : inv02 port map ( Y=>nx10460, A=>nx180);
   ix10461 : inv02 port map ( Y=>nx10462, A=>nx192);
   ix10463 : inv02 port map ( Y=>nx10464, A=>nx192);
   ix10465 : inv02 port map ( Y=>nx10466, A=>nx200);
   ix10467 : inv02 port map ( Y=>nx10468, A=>nx200);
   ix10469 : inv02 port map ( Y=>nx10470, A=>nx206);
   ix10471 : inv02 port map ( Y=>nx10472, A=>nx206);
   ix10473 : inv02 port map ( Y=>nx10474, A=>nx214);
   ix10475 : inv02 port map ( Y=>nx10476, A=>nx214);
   ix10477 : inv02 port map ( Y=>nx10478, A=>nx222);
   ix10479 : inv02 port map ( Y=>nx10480, A=>nx222);
   ix10481 : inv02 port map ( Y=>nx10482, A=>nx226);
   ix10483 : inv02 port map ( Y=>nx10484, A=>nx226);
   ix10485 : inv02 port map ( Y=>nx10486, A=>nx230);
   ix10487 : inv02 port map ( Y=>nx10488, A=>nx230);
   ix8951 : nor02ii port map ( Y=>sel_que_0, A0=>nx6829, A1=>nx6885);
   ix8961 : nor02ii port map ( Y=>sel_que_1, A0=>nx6839, A1=>nx6885);
   ix8971 : nor02ii port map ( Y=>sel_que_2, A0=>nx6843, A1=>nx6885);
   ix8979 : nor02ii port map ( Y=>sel_que_3, A0=>nx6847, A1=>nx6885);
   ix8987 : nor02ii port map ( Y=>sel_que_4, A0=>nx6829, A1=>nx6905);
   ix8991 : nor02ii port map ( Y=>sel_que_5, A0=>nx6839, A1=>nx6905);
   ix8995 : nor02ii port map ( Y=>sel_que_6, A0=>nx6843, A1=>nx6905);
   ix8999 : nor02ii port map ( Y=>sel_que_7, A0=>nx6847, A1=>nx6905);
   ix9007 : nor02ii port map ( Y=>sel_que_8, A0=>nx6829, A1=>nx6915);
   ix9011 : nor02ii port map ( Y=>sel_que_9, A0=>nx6839, A1=>nx6915);
   ix9015 : nor02ii port map ( Y=>sel_que_10, A0=>nx6843, A1=>nx6915);
   ix9019 : nor02ii port map ( Y=>sel_que_11, A0=>nx6847, A1=>nx6915);
   ix9053 : nor02ii port map ( Y=>sel_que_17, A0=>nx6893, A1=>nx6885);
   ix9063 : nor02ii port map ( Y=>sel_que_18, A0=>nx6897, A1=>nx6885);
   ix9071 : nor02ii port map ( Y=>sel_que_19, A0=>nx6901, A1=>nx6885);
   ix6906 : nor02ii port map ( Y=>nx6905, A0=>cache_in_sel(3), A1=>
      cache_in_sel(2));
   ix9079 : nor02ii port map ( Y=>sel_que_21, A0=>nx6893, A1=>nx6905);
   ix9083 : nor02ii port map ( Y=>sel_que_22, A0=>nx6897, A1=>nx6905);
   ix9087 : nor02ii port map ( Y=>sel_que_23, A0=>nx6901, A1=>nx6905);
   ix6916 : nor02ii port map ( Y=>nx6915, A0=>cache_in_sel(2), A1=>
      cache_in_sel(3));
   ix9095 : nor02ii port map ( Y=>sel_que_25, A0=>nx6893, A1=>nx6915);
   ix9099 : nor02ii port map ( Y=>sel_que_26, A0=>nx6897, A1=>nx6915);
   ix9103 : nor02ii port map ( Y=>sel_que_27, A0=>nx6901, A1=>nx6915);
   ix223 : nor02ii port map ( Y=>nx222, A0=>nx6931, A1=>nx62);
   ix231 : nor02ii port map ( Y=>nx230, A0=>nx6945, A1=>nx88);
   ix207 : nor02ii port map ( Y=>nx206, A0=>nx10374, A1=>nx28);
   ix123 : nor02ii port map ( Y=>nx122, A0=>nx10374, A1=>nx62);
   ix65 : nor02ii port map ( Y=>nx64, A0=>nx6949, A1=>nx62);
   ix49 : nor02ii port map ( Y=>nx48, A0=>nx6949, A1=>nx28);
   ix31 : nor02ii port map ( Y=>nx30, A0=>nx6931, A1=>nx28);
   ix10493 : inv02 port map ( Y=>nx10494, A=>nx6937);
   ix10495 : inv02 port map ( Y=>nx10496, A=>nx6937);
   ix10497 : inv02 port map ( Y=>nx10498, A=>nx6939);
   ix10499 : inv02 port map ( Y=>nx10500, A=>nx6939);
   ix10501 : inv01 port map ( Y=>nx10502, A=>nx6961);
   ix10503 : inv01 port map ( Y=>nx10504, A=>nx6961);
   ix10505 : inv02 port map ( Y=>nx10506, A=>nx6833);
   ix10507 : inv02 port map ( Y=>nx10508, A=>nx6835);
   ix10509 : inv01 port map ( Y=>nx10510, A=>in_word(15));
   ix10511 : inv01 port map ( Y=>nx10512, A=>nx10510);
   ix10513 : inv01 port map ( Y=>nx10514, A=>nx10510);
   ix10515 : inv01 port map ( Y=>nx10516, A=>nx10510);
   ix10517 : inv01 port map ( Y=>nx10518, A=>nx10510);
   ix10519 : inv01 port map ( Y=>nx10520, A=>in_word(14));
   ix10521 : inv01 port map ( Y=>nx10522, A=>nx10520);
   ix10523 : inv01 port map ( Y=>nx10524, A=>nx10520);
   ix10525 : inv01 port map ( Y=>nx10526, A=>nx10520);
   ix10527 : inv01 port map ( Y=>nx10528, A=>nx10520);
   ix10529 : inv01 port map ( Y=>nx10530, A=>in_word(13));
   ix10531 : inv01 port map ( Y=>nx10532, A=>nx10530);
   ix10533 : inv01 port map ( Y=>nx10534, A=>nx10530);
   ix10535 : inv01 port map ( Y=>nx10536, A=>nx10530);
   ix10537 : inv01 port map ( Y=>nx10538, A=>nx10530);
   ix10539 : inv01 port map ( Y=>nx10540, A=>in_word(12));
   ix10541 : inv01 port map ( Y=>nx10542, A=>nx10540);
   ix10543 : inv01 port map ( Y=>nx10544, A=>nx10540);
   ix10545 : inv01 port map ( Y=>nx10546, A=>nx10540);
   ix10547 : inv01 port map ( Y=>nx10548, A=>nx10540);
   ix10549 : inv01 port map ( Y=>nx10550, A=>in_word(11));
   ix10551 : inv01 port map ( Y=>nx10552, A=>nx10550);
   ix10553 : inv01 port map ( Y=>nx10554, A=>nx10550);
   ix10555 : inv01 port map ( Y=>nx10556, A=>nx10550);
   ix10557 : inv01 port map ( Y=>nx10558, A=>nx10550);
   ix10559 : inv01 port map ( Y=>nx10560, A=>in_word(10));
   ix10561 : inv01 port map ( Y=>nx10562, A=>nx10560);
   ix10563 : inv01 port map ( Y=>nx10564, A=>nx10560);
   ix10565 : inv01 port map ( Y=>nx10566, A=>nx10560);
   ix10567 : inv01 port map ( Y=>nx10568, A=>nx10560);
   ix10569 : inv01 port map ( Y=>nx10570, A=>in_word(9));
   ix10571 : inv01 port map ( Y=>nx10572, A=>nx10570);
   ix10573 : inv01 port map ( Y=>nx10574, A=>nx10570);
   ix10575 : inv01 port map ( Y=>nx10576, A=>nx10570);
   ix10577 : inv01 port map ( Y=>nx10578, A=>nx10570);
   ix10579 : inv01 port map ( Y=>nx10580, A=>in_word(8));
   ix10581 : inv01 port map ( Y=>nx10582, A=>nx10580);
   ix10583 : inv01 port map ( Y=>nx10584, A=>nx10580);
   ix10585 : inv01 port map ( Y=>nx10586, A=>nx10580);
   ix10587 : inv01 port map ( Y=>nx10588, A=>nx10580);
   ix10589 : inv01 port map ( Y=>nx10590, A=>in_word(7));
   ix10591 : inv01 port map ( Y=>nx10592, A=>nx10590);
   ix10593 : inv01 port map ( Y=>nx10594, A=>nx10590);
   ix10595 : inv01 port map ( Y=>nx10596, A=>nx10590);
   ix10597 : inv01 port map ( Y=>nx10598, A=>nx10590);
   ix10599 : inv01 port map ( Y=>nx10600, A=>in_word(6));
   ix10601 : inv01 port map ( Y=>nx10602, A=>nx10600);
   ix10603 : inv01 port map ( Y=>nx10604, A=>nx10600);
   ix10605 : inv01 port map ( Y=>nx10606, A=>nx10600);
   ix10607 : inv01 port map ( Y=>nx10608, A=>nx10600);
   ix10609 : inv01 port map ( Y=>nx10610, A=>in_word(5));
   ix10611 : inv01 port map ( Y=>nx10612, A=>nx10610);
   ix10613 : inv01 port map ( Y=>nx10614, A=>nx10610);
   ix10615 : inv01 port map ( Y=>nx10616, A=>nx10610);
   ix10617 : inv01 port map ( Y=>nx10618, A=>nx10610);
   ix10619 : inv01 port map ( Y=>nx10620, A=>in_word(4));
   ix10621 : inv01 port map ( Y=>nx10622, A=>nx10620);
   ix10623 : inv01 port map ( Y=>nx10624, A=>nx10620);
   ix10625 : inv01 port map ( Y=>nx10626, A=>nx10620);
   ix10627 : inv01 port map ( Y=>nx10628, A=>nx10620);
   ix10629 : inv01 port map ( Y=>nx10630, A=>in_word(3));
   ix10631 : inv01 port map ( Y=>nx10632, A=>nx10630);
   ix10633 : inv01 port map ( Y=>nx10634, A=>nx10630);
   ix10635 : inv01 port map ( Y=>nx10636, A=>nx10630);
   ix10637 : inv01 port map ( Y=>nx10638, A=>nx10630);
   ix10639 : inv01 port map ( Y=>nx10640, A=>in_word(2));
   ix10641 : inv01 port map ( Y=>nx10642, A=>nx10640);
   ix10643 : inv01 port map ( Y=>nx10644, A=>nx10640);
   ix10645 : inv01 port map ( Y=>nx10646, A=>nx10640);
   ix10647 : inv01 port map ( Y=>nx10648, A=>nx10640);
   ix10649 : inv01 port map ( Y=>nx10650, A=>in_word(1));
   ix10651 : inv01 port map ( Y=>nx10652, A=>nx10650);
   ix10653 : inv01 port map ( Y=>nx10654, A=>nx10650);
   ix10655 : inv01 port map ( Y=>nx10656, A=>nx10650);
   ix10657 : inv01 port map ( Y=>nx10658, A=>nx10650);
   ix10659 : inv01 port map ( Y=>nx10660, A=>in_word(0));
   ix10661 : inv01 port map ( Y=>nx10662, A=>nx10660);
   ix10663 : inv01 port map ( Y=>nx10664, A=>nx10660);
   ix10665 : inv01 port map ( Y=>nx10666, A=>nx10660);
   ix10667 : inv01 port map ( Y=>nx10668, A=>nx10660);
   ix10689 : inv02 port map ( Y=>nx10690, A=>nx10742);
   ix10691 : inv02 port map ( Y=>nx10692, A=>nx10742);
   ix10693 : inv02 port map ( Y=>nx10694, A=>nx10742);
   ix10695 : inv02 port map ( Y=>nx10696, A=>nx10742);
   ix10697 : inv02 port map ( Y=>nx10698, A=>nx10742);
   ix10699 : inv02 port map ( Y=>nx10700, A=>nx10742);
   ix10701 : inv02 port map ( Y=>nx10702, A=>nx10742);
   ix10703 : inv02 port map ( Y=>nx10704, A=>nx10744);
   ix10705 : inv02 port map ( Y=>nx10706, A=>nx10744);
   ix10707 : inv02 port map ( Y=>nx10708, A=>nx10744);
   ix10709 : inv02 port map ( Y=>nx10710, A=>nx10744);
   ix10711 : inv02 port map ( Y=>nx10712, A=>nx10744);
   ix10713 : inv02 port map ( Y=>nx10714, A=>nx10746);
   ix10715 : inv02 port map ( Y=>nx10716, A=>nx10746);
   ix10717 : inv02 port map ( Y=>nx10718, A=>nx10746);
   ix10719 : inv02 port map ( Y=>nx10720, A=>nx10746);
   ix10721 : inv02 port map ( Y=>nx10722, A=>nx10746);
   ix10723 : inv02 port map ( Y=>nx10724, A=>nx10746);
   ix10725 : inv02 port map ( Y=>nx10726, A=>nx10746);
   ix10727 : inv02 port map ( Y=>nx10728, A=>nx10748);
   ix10729 : inv02 port map ( Y=>nx10730, A=>nx10748);
   ix10731 : inv02 port map ( Y=>nx10732, A=>nx10748);
   ix10733 : inv02 port map ( Y=>nx10734, A=>nx10748);
   ix10735 : inv02 port map ( Y=>nx10736, A=>nx10748);
   ix10741 : inv02 port map ( Y=>nx10742, A=>reset);
   ix10743 : inv02 port map ( Y=>nx10744, A=>reset);
   ix10745 : inv02 port map ( Y=>nx10746, A=>clk);
   ix10747 : inv02 port map ( Y=>nx10748, A=>clk);
end Dataflow ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity AdvancedCounter_16 is
   port (
      clk : IN std_logic ;
      reset : IN std_logic ;
      enable : IN std_logic ;
      mode_in : IN std_logic_vector (1 DOWNTO 0) ;
      max_val_in : IN std_logic_vector (15 DOWNTO 0) ;
      max_reached_out : OUT std_logic ;
      counter_out : OUT std_logic_vector (15 DOWNTO 0)) ;
end AdvancedCounter_16 ;

architecture behavioural_unfold_2902 of AdvancedCounter_16 is
   signal counter_out_0_EXMPLR, counter_out_15_EXMPLR, counter_out_14_EXMPLR, 
      nx149, counter_out_13_EXMPLR, counter_out_12_EXMPLR, nx152, 
      counter_out_11_EXMPLR, counter_out_10_EXMPLR, nx155, 
      counter_out_9_EXMPLR, counter_out_8_EXMPLR, nx157, 
      counter_out_7_EXMPLR, counter_out_6_EXMPLR, nx159, 
      counter_out_5_EXMPLR, counter_out_4_EXMPLR, nx161, 
      counter_out_3_EXMPLR, counter_out_2_EXMPLR, counter_out_1_EXMPLR, 
      counter_out_dup0_0, nx22, nx34, nx46, nx70, nx94, nx118, nx142, nx166, 
      nx174, nx192, nx206, nx224, nx246, nx173, nx183, nx193, nx203, nx213, 
      nx223, nx233, nx243, nx253, nx263, nx273, nx283, nx293, nx303, nx313, 
      nx323, nx339, nx344, nx348, nx350, nx353, nx358, nx362, nx364, nx367, 
      nx372, nx376, nx378, nx381, nx386, nx390, nx392, nx395, nx400, nx404, 
      nx406, nx409, nx414, nx419, nx424, nx428, nx430, nx436, nx439, nx445, 
      nx447, nx449, nx451, nx458, nx460, nx462, nx464, nx466, nx468, nx470, 
      nx472, nx474: std_logic ;

begin
   counter_out(15) <= counter_out_0_EXMPLR ;
   counter_out(14) <= counter_out_0_EXMPLR ;
   counter_out(13) <= counter_out_0_EXMPLR ;
   counter_out(12) <= counter_out_0_EXMPLR ;
   counter_out(11) <= counter_out_0_EXMPLR ;
   counter_out(10) <= counter_out_0_EXMPLR ;
   counter_out(9) <= counter_out_0_EXMPLR ;
   counter_out(8) <= counter_out_0_EXMPLR ;
   counter_out(7) <= counter_out_0_EXMPLR ;
   counter_out(6) <= counter_out_0_EXMPLR ;
   counter_out(5) <= counter_out_0_EXMPLR ;
   counter_out(4) <= counter_out_0_EXMPLR ;
   counter_out(3) <= counter_out_0_EXMPLR ;
   counter_out(2) <= counter_out_0_EXMPLR ;
   counter_out(1) <= counter_out_0_EXMPLR ;
   counter_out(0) <= counter_out_0_EXMPLR ;
   ix140 : fake_gnd port map ( Y=>counter_out_0_EXMPLR);
   ix251 : and04 port map ( Y=>max_reached_out, A0=>nx192, A1=>nx206, A2=>
      nx224, A3=>nx246);
   ix324 : mux21_ni port map ( Y=>nx323, A0=>counter_out_15_EXMPLR, A1=>
      nx174, S0=>nx474);
   ix314 : mux21_ni port map ( Y=>nx313, A0=>counter_out_14_EXMPLR, A1=>
      nx166, S0=>nx472);
   reg_counter_data_14 : dffr port map ( Q=>counter_out_14_EXMPLR, QB=>nx339, 
      D=>nx313, CLK=>clk, R=>nx462);
   ix345 : nand02 port map ( Y=>nx344, A0=>counter_out_13_EXMPLR, A1=>nx152
   );
   ix304 : mux21 port map ( Y=>nx303, A0=>nx348, A1=>nx350, S0=>nx472);
   reg_counter_data_13 : dffr port map ( Q=>counter_out_13_EXMPLR, QB=>nx348, 
      D=>nx303, CLK=>clk, R=>nx462);
   ix351 : oai21 port map ( Y=>nx350, A0=>nx152, A1=>counter_out_13_EXMPLR, 
      B0=>nx344);
   ix294 : mux21_ni port map ( Y=>nx293, A0=>counter_out_12_EXMPLR, A1=>
      nx142, S0=>nx472);
   reg_counter_data_12 : dffr port map ( Q=>counter_out_12_EXMPLR, QB=>nx353, 
      D=>nx293, CLK=>clk, R=>nx462);
   ix359 : nand02 port map ( Y=>nx358, A0=>counter_out_11_EXMPLR, A1=>nx155
   );
   ix284 : mux21 port map ( Y=>nx283, A0=>nx362, A1=>nx364, S0=>nx472);
   reg_counter_data_11 : dffr port map ( Q=>counter_out_11_EXMPLR, QB=>nx362, 
      D=>nx283, CLK=>clk, R=>nx462);
   ix365 : oai21 port map ( Y=>nx364, A0=>nx155, A1=>counter_out_11_EXMPLR, 
      B0=>nx358);
   ix274 : mux21_ni port map ( Y=>nx273, A0=>counter_out_10_EXMPLR, A1=>
      nx118, S0=>nx472);
   reg_counter_data_10 : dffr port map ( Q=>counter_out_10_EXMPLR, QB=>nx367, 
      D=>nx273, CLK=>clk, R=>nx462);
   ix373 : nand02 port map ( Y=>nx372, A0=>counter_out_9_EXMPLR, A1=>nx157);
   ix264 : mux21 port map ( Y=>nx263, A0=>nx376, A1=>nx378, S0=>nx472);
   reg_counter_data_9 : dffr port map ( Q=>counter_out_9_EXMPLR, QB=>nx376, 
      D=>nx263, CLK=>clk, R=>nx462);
   ix379 : oai21 port map ( Y=>nx378, A0=>nx157, A1=>counter_out_9_EXMPLR, 
      B0=>nx372);
   ix254 : mux21_ni port map ( Y=>nx253, A0=>counter_out_8_EXMPLR, A1=>nx94, 
      S0=>nx472);
   reg_counter_data_8 : dffr port map ( Q=>counter_out_8_EXMPLR, QB=>nx381, 
      D=>nx253, CLK=>clk, R=>nx462);
   ix387 : nand02 port map ( Y=>nx386, A0=>counter_out_7_EXMPLR, A1=>nx159);
   ix244 : mux21 port map ( Y=>nx243, A0=>nx390, A1=>nx392, S0=>nx470);
   reg_counter_data_7 : dffr port map ( Q=>counter_out_7_EXMPLR, QB=>nx390, 
      D=>nx243, CLK=>clk, R=>nx464);
   ix393 : oai21 port map ( Y=>nx392, A0=>nx159, A1=>counter_out_7_EXMPLR, 
      B0=>nx386);
   ix234 : mux21_ni port map ( Y=>nx233, A0=>counter_out_6_EXMPLR, A1=>nx70, 
      S0=>nx470);
   reg_counter_data_6 : dffr port map ( Q=>counter_out_6_EXMPLR, QB=>nx395, 
      D=>nx233, CLK=>clk, R=>nx464);
   ix401 : nand02 port map ( Y=>nx400, A0=>counter_out_5_EXMPLR, A1=>nx161);
   ix224 : mux21 port map ( Y=>nx223, A0=>nx404, A1=>nx406, S0=>nx470);
   reg_counter_data_5 : dffr port map ( Q=>counter_out_5_EXMPLR, QB=>nx404, 
      D=>nx223, CLK=>clk, R=>nx464);
   ix407 : oai21 port map ( Y=>nx406, A0=>nx161, A1=>counter_out_5_EXMPLR, 
      B0=>nx400);
   ix214 : mux21_ni port map ( Y=>nx213, A0=>counter_out_4_EXMPLR, A1=>nx46, 
      S0=>nx470);
   reg_counter_data_4 : dffr port map ( Q=>counter_out_4_EXMPLR, QB=>nx409, 
      D=>nx213, CLK=>clk, R=>nx464);
   ix47 : aoi21 port map ( Y=>nx46, A0=>nx414, A1=>nx409, B0=>nx161);
   ix415 : nand04 port map ( Y=>nx414, A0=>counter_out_3_EXMPLR, A1=>
      counter_out_2_EXMPLR, A2=>counter_out_1_EXMPLR, A3=>counter_out_dup0_0
   );
   reg_counter_data_3 : dffr port map ( Q=>counter_out_3_EXMPLR, QB=>OPEN, D
      =>nx203, CLK=>clk, R=>nx466);
   ix204 : mux21_ni port map ( Y=>nx203, A0=>counter_out_3_EXMPLR, A1=>nx34, 
      S0=>nx470);
   ix35 : xnor2 port map ( Y=>nx34, A0=>counter_out_3_EXMPLR, A1=>nx419);
   ix420 : nand03 port map ( Y=>nx419, A0=>counter_out_2_EXMPLR, A1=>
      counter_out_1_EXMPLR, A2=>counter_out_dup0_0);
   reg_counter_data_2 : dffr port map ( Q=>counter_out_2_EXMPLR, QB=>OPEN, D
      =>nx193, CLK=>clk, R=>nx464);
   ix194 : mux21_ni port map ( Y=>nx193, A0=>counter_out_2_EXMPLR, A1=>nx22, 
      S0=>nx470);
   ix23 : xnor2 port map ( Y=>nx22, A0=>counter_out_2_EXMPLR, A1=>nx424);
   ix184 : mux21 port map ( Y=>nx183, A0=>nx428, A1=>nx430, S0=>nx470);
   reg_counter_data_1 : dffr port map ( Q=>counter_out_1_EXMPLR, QB=>nx428, 
      D=>nx183, CLK=>clk, R=>nx464);
   ix431 : oai21 port map ( Y=>nx430, A0=>counter_out_dup0_0, A1=>
      counter_out_1_EXMPLR, B0=>nx424);
   reg_counter_data_0 : dffr port map ( Q=>counter_out_dup0_0, QB=>nx436, D
      =>nx173, CLK=>clk, R=>nx464);
   reg_counter_data_15 : dffr port map ( Q=>counter_out_15_EXMPLR, QB=>nx439, 
      D=>nx323, CLK=>clk, R=>nx466);
   ix247 : and04 port map ( Y=>nx246, A0=>nx445, A1=>nx447, A2=>nx449, A3=>
      nx451);
   ix448 : xnor2 port map ( Y=>nx447, A0=>counter_out_2_EXMPLR, A1=>
      max_val_in(2));
   ix450 : xnor2 port map ( Y=>nx449, A0=>counter_out_3_EXMPLR, A1=>
      max_val_in(3));
   ix193 : and04 port map ( Y=>nx192, A0=>nx439, A1=>nx339, A2=>nx348, A3=>
      nx353);
   ix175 : xor2 port map ( Y=>nx174, A0=>nx149, A1=>counter_out_15_EXMPLR);
   ix173 : nor02ii port map ( Y=>nx149, A0=>nx344, A1=>counter_out_14_EXMPLR
   );
   ix167 : xor2 port map ( Y=>nx166, A0=>nx339, A1=>nx344);
   ix149 : nor02ii port map ( Y=>nx152, A0=>nx358, A1=>counter_out_12_EXMPLR
   );
   ix143 : xor2 port map ( Y=>nx142, A0=>nx353, A1=>nx358);
   ix125 : nor02ii port map ( Y=>nx155, A0=>nx372, A1=>counter_out_10_EXMPLR
   );
   ix119 : xor2 port map ( Y=>nx118, A0=>nx367, A1=>nx372);
   ix101 : nor02ii port map ( Y=>nx157, A0=>nx386, A1=>counter_out_8_EXMPLR
   );
   ix95 : xor2 port map ( Y=>nx94, A0=>nx381, A1=>nx386);
   ix77 : nor02ii port map ( Y=>nx159, A0=>nx400, A1=>counter_out_6_EXMPLR);
   ix71 : xor2 port map ( Y=>nx70, A0=>nx395, A1=>nx400);
   ix53 : nor02ii port map ( Y=>nx161, A0=>nx414, A1=>counter_out_4_EXMPLR);
   ix425 : or02 port map ( Y=>nx424, A0=>nx428, A1=>nx436);
   ix174 : xnor2 port map ( Y=>nx173, A0=>nx436, A1=>nx474);
   ix207 : and04 port map ( Y=>nx206, A0=>nx362, A1=>nx367, A2=>nx376, A3=>
      nx381);
   ix225 : and04 port map ( Y=>nx224, A0=>nx390, A1=>nx395, A2=>nx404, A3=>
      nx458);
   ix217 : xnor2 port map ( Y=>nx458, A0=>max_val_in(0), A1=>
      counter_out_dup0_0);
   ix446 : xor2 port map ( Y=>nx445, A0=>nx428, A1=>max_val_in(1));
   ix452 : xor2 port map ( Y=>nx451, A0=>nx409, A1=>max_val_in(4));
   ix459 : inv01 port map ( Y=>nx460, A=>reset);
   ix461 : inv02 port map ( Y=>nx462, A=>nx460);
   ix463 : inv02 port map ( Y=>nx464, A=>nx460);
   ix465 : inv02 port map ( Y=>nx466, A=>nx460);
   ix467 : inv01 port map ( Y=>nx468, A=>enable);
   ix469 : inv02 port map ( Y=>nx470, A=>nx468);
   ix471 : inv02 port map ( Y=>nx472, A=>nx468);
   ix473 : inv02 port map ( Y=>nx474, A=>nx468);
end behavioural_unfold_2902 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Controller is
   port (
      clk : IN std_logic ;
      reset : IN std_logic ;
      io_ready_in : IN std_logic ;
      io_done_out : OUT std_logic ;
      mem_data_in : IN std_logic_vector (15 DOWNTO 0) ;
      mem_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
      mem_addr_out : OUT std_logic_vector (15 DOWNTO 0) ;
      mem_write_out : OUT std_logic ;
      mem_read_out : OUT std_logic ;
      wind_en : OUT std_logic ;
      wind_rst : OUT std_logic ;
      wind_col_in_4_15 : OUT std_logic ;
      wind_col_in_4_14 : OUT std_logic ;
      wind_col_in_4_13 : OUT std_logic ;
      wind_col_in_4_12 : OUT std_logic ;
      wind_col_in_4_11 : OUT std_logic ;
      wind_col_in_4_10 : OUT std_logic ;
      wind_col_in_4_9 : OUT std_logic ;
      wind_col_in_4_8 : OUT std_logic ;
      wind_col_in_4_7 : OUT std_logic ;
      wind_col_in_4_6 : OUT std_logic ;
      wind_col_in_4_5 : OUT std_logic ;
      wind_col_in_4_4 : OUT std_logic ;
      wind_col_in_4_3 : OUT std_logic ;
      wind_col_in_4_2 : OUT std_logic ;
      wind_col_in_4_1 : OUT std_logic ;
      wind_col_in_4_0 : OUT std_logic ;
      wind_col_in_3_15 : OUT std_logic ;
      wind_col_in_3_14 : OUT std_logic ;
      wind_col_in_3_13 : OUT std_logic ;
      wind_col_in_3_12 : OUT std_logic ;
      wind_col_in_3_11 : OUT std_logic ;
      wind_col_in_3_10 : OUT std_logic ;
      wind_col_in_3_9 : OUT std_logic ;
      wind_col_in_3_8 : OUT std_logic ;
      wind_col_in_3_7 : OUT std_logic ;
      wind_col_in_3_6 : OUT std_logic ;
      wind_col_in_3_5 : OUT std_logic ;
      wind_col_in_3_4 : OUT std_logic ;
      wind_col_in_3_3 : OUT std_logic ;
      wind_col_in_3_2 : OUT std_logic ;
      wind_col_in_3_1 : OUT std_logic ;
      wind_col_in_3_0 : OUT std_logic ;
      wind_col_in_2_15 : OUT std_logic ;
      wind_col_in_2_14 : OUT std_logic ;
      wind_col_in_2_13 : OUT std_logic ;
      wind_col_in_2_12 : OUT std_logic ;
      wind_col_in_2_11 : OUT std_logic ;
      wind_col_in_2_10 : OUT std_logic ;
      wind_col_in_2_9 : OUT std_logic ;
      wind_col_in_2_8 : OUT std_logic ;
      wind_col_in_2_7 : OUT std_logic ;
      wind_col_in_2_6 : OUT std_logic ;
      wind_col_in_2_5 : OUT std_logic ;
      wind_col_in_2_4 : OUT std_logic ;
      wind_col_in_2_3 : OUT std_logic ;
      wind_col_in_2_2 : OUT std_logic ;
      wind_col_in_2_1 : OUT std_logic ;
      wind_col_in_2_0 : OUT std_logic ;
      wind_col_in_1_15 : OUT std_logic ;
      wind_col_in_1_14 : OUT std_logic ;
      wind_col_in_1_13 : OUT std_logic ;
      wind_col_in_1_12 : OUT std_logic ;
      wind_col_in_1_11 : OUT std_logic ;
      wind_col_in_1_10 : OUT std_logic ;
      wind_col_in_1_9 : OUT std_logic ;
      wind_col_in_1_8 : OUT std_logic ;
      wind_col_in_1_7 : OUT std_logic ;
      wind_col_in_1_6 : OUT std_logic ;
      wind_col_in_1_5 : OUT std_logic ;
      wind_col_in_1_4 : OUT std_logic ;
      wind_col_in_1_3 : OUT std_logic ;
      wind_col_in_1_2 : OUT std_logic ;
      wind_col_in_1_1 : OUT std_logic ;
      wind_col_in_1_0 : OUT std_logic ;
      wind_col_in_0_15 : OUT std_logic ;
      wind_col_in_0_14 : OUT std_logic ;
      wind_col_in_0_13 : OUT std_logic ;
      wind_col_in_0_12 : OUT std_logic ;
      wind_col_in_0_11 : OUT std_logic ;
      wind_col_in_0_10 : OUT std_logic ;
      wind_col_in_0_9 : OUT std_logic ;
      wind_col_in_0_8 : OUT std_logic ;
      wind_col_in_0_7 : OUT std_logic ;
      wind_col_in_0_6 : OUT std_logic ;
      wind_col_in_0_5 : OUT std_logic ;
      wind_col_in_0_4 : OUT std_logic ;
      wind_col_in_0_3 : OUT std_logic ;
      wind_col_in_0_2 : OUT std_logic ;
      wind_col_in_0_1 : OUT std_logic ;
      wind_col_in_0_0 : OUT std_logic ;
      filter_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
      filter_ready_out : OUT std_logic ;
      filter_reset : OUT std_logic ;
      comp_unit_ready : OUT std_logic ;
      comp_unit_operation : OUT std_logic ;
      comp_unit_flt_size : OUT std_logic ;
      comp_unit_relu : OUT std_logic ;
      comp_unit_data1_out : OUT std_logic_vector (15 DOWNTO 0) ;
      comp_unit_data2_out : OUT std_logic_vector (15 DOWNTO 0) ;
      comp_unit_buffer_finished : IN std_logic ;
      comp_unit_finished : IN std_logic ;
      comp_unit_data1_in : IN std_logic_vector (15 DOWNTO 0) ;
      comp_unit_data2_in : IN std_logic_vector (15 DOWNTO 0) ;
      argmax_ready : OUT std_logic ;
      argmax_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
      argmax_data_in : IN std_logic_vector (15 DOWNTO 0)) ;
end Controller ;

architecture Mixed of Controller is
   component Cache_5_16_28_5
      port (
         in_word : IN std_logic_vector (15 DOWNTO 0) ;
         cache_in_sel : IN std_logic_vector (4 DOWNTO 0) ;
         cache_out_sel : IN std_logic_vector (4 DOWNTO 0) ;
         decoder_enable : IN std_logic ;
         out_column_0_15 : OUT std_logic ;
         out_column_0_14 : OUT std_logic ;
         out_column_0_13 : OUT std_logic ;
         out_column_0_12 : OUT std_logic ;
         out_column_0_11 : OUT std_logic ;
         out_column_0_10 : OUT std_logic ;
         out_column_0_9 : OUT std_logic ;
         out_column_0_8 : OUT std_logic ;
         out_column_0_7 : OUT std_logic ;
         out_column_0_6 : OUT std_logic ;
         out_column_0_5 : OUT std_logic ;
         out_column_0_4 : OUT std_logic ;
         out_column_0_3 : OUT std_logic ;
         out_column_0_2 : OUT std_logic ;
         out_column_0_1 : OUT std_logic ;
         out_column_0_0 : OUT std_logic ;
         out_column_1_15 : OUT std_logic ;
         out_column_1_14 : OUT std_logic ;
         out_column_1_13 : OUT std_logic ;
         out_column_1_12 : OUT std_logic ;
         out_column_1_11 : OUT std_logic ;
         out_column_1_10 : OUT std_logic ;
         out_column_1_9 : OUT std_logic ;
         out_column_1_8 : OUT std_logic ;
         out_column_1_7 : OUT std_logic ;
         out_column_1_6 : OUT std_logic ;
         out_column_1_5 : OUT std_logic ;
         out_column_1_4 : OUT std_logic ;
         out_column_1_3 : OUT std_logic ;
         out_column_1_2 : OUT std_logic ;
         out_column_1_1 : OUT std_logic ;
         out_column_1_0 : OUT std_logic ;
         out_column_2_15 : OUT std_logic ;
         out_column_2_14 : OUT std_logic ;
         out_column_2_13 : OUT std_logic ;
         out_column_2_12 : OUT std_logic ;
         out_column_2_11 : OUT std_logic ;
         out_column_2_10 : OUT std_logic ;
         out_column_2_9 : OUT std_logic ;
         out_column_2_8 : OUT std_logic ;
         out_column_2_7 : OUT std_logic ;
         out_column_2_6 : OUT std_logic ;
         out_column_2_5 : OUT std_logic ;
         out_column_2_4 : OUT std_logic ;
         out_column_2_3 : OUT std_logic ;
         out_column_2_2 : OUT std_logic ;
         out_column_2_1 : OUT std_logic ;
         out_column_2_0 : OUT std_logic ;
         out_column_3_15 : OUT std_logic ;
         out_column_3_14 : OUT std_logic ;
         out_column_3_13 : OUT std_logic ;
         out_column_3_12 : OUT std_logic ;
         out_column_3_11 : OUT std_logic ;
         out_column_3_10 : OUT std_logic ;
         out_column_3_9 : OUT std_logic ;
         out_column_3_8 : OUT std_logic ;
         out_column_3_7 : OUT std_logic ;
         out_column_3_6 : OUT std_logic ;
         out_column_3_5 : OUT std_logic ;
         out_column_3_4 : OUT std_logic ;
         out_column_3_3 : OUT std_logic ;
         out_column_3_2 : OUT std_logic ;
         out_column_3_1 : OUT std_logic ;
         out_column_3_0 : OUT std_logic ;
         out_column_4_15 : OUT std_logic ;
         out_column_4_14 : OUT std_logic ;
         out_column_4_13 : OUT std_logic ;
         out_column_4_12 : OUT std_logic ;
         out_column_4_11 : OUT std_logic ;
         out_column_4_10 : OUT std_logic ;
         out_column_4_9 : OUT std_logic ;
         out_column_4_8 : OUT std_logic ;
         out_column_4_7 : OUT std_logic ;
         out_column_4_6 : OUT std_logic ;
         out_column_4_5 : OUT std_logic ;
         out_column_4_4 : OUT std_logic ;
         out_column_4_3 : OUT std_logic ;
         out_column_4_2 : OUT std_logic ;
         out_column_4_1 : OUT std_logic ;
         out_column_4_0 : OUT std_logic ;
         clk : IN std_logic ;
         reset : IN std_logic) ;
   end component ;
   component AdvancedCounter_16
      port (
         clk : IN std_logic ;
         reset : IN std_logic ;
         enable : IN std_logic ;
         mode_in : IN std_logic_vector (1 DOWNTO 0) ;
         max_val_in : IN std_logic_vector (15 DOWNTO 0) ;
         max_reached_out : OUT std_logic ;
         counter_out : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   signal current_state_13, wind_width_count_4, wind_width_count_3, 
      wind_width_count_2, wind_width_count_1, wind_width_count_0, 
      cache_height_count_en, cache_height_ended, max_height_2, max_height_0, 
      cache_width_count_4, cache_width_count_3, cache_width_count_2, 
      cache_width_count_1, cache_width_count_0, cache_data_in_15, 
      cache_data_in_14, cache_data_in_13, cache_data_in_12, cache_data_in_11, 
      cache_data_in_10, cache_data_in_9, cache_data_in_8, cache_data_in_7, 
      cache_data_in_6, cache_data_in_5, cache_data_in_4, cache_data_in_3, 
      cache_data_in_2, cache_data_in_1, cache_data_in_0, cache_data_out_4_15, 
      cache_data_out_4_14, cache_data_out_4_13, cache_data_out_4_12, 
      cache_data_out_4_11, cache_data_out_4_10, cache_data_out_4_9, 
      cache_data_out_4_8, cache_data_out_4_7, cache_data_out_4_6, 
      cache_data_out_4_5, cache_data_out_4_4, cache_data_out_4_3, 
      cache_data_out_4_2, cache_data_out_4_1, cache_data_out_4_0, 
      cache_data_out_3_15, cache_data_out_3_14, cache_data_out_3_13, 
      cache_data_out_3_12, cache_data_out_3_11, cache_data_out_3_10, 
      cache_data_out_3_9, cache_data_out_3_8, cache_data_out_3_7, 
      cache_data_out_3_6, cache_data_out_3_5, cache_data_out_3_4, 
      cache_data_out_3_3, cache_data_out_3_2, cache_data_out_3_1, 
      cache_data_out_3_0, cache_data_out_2_15, cache_data_out_2_14, 
      cache_data_out_2_13, cache_data_out_2_12, cache_data_out_2_11, 
      cache_data_out_2_10, cache_data_out_2_9, cache_data_out_2_8, 
      cache_data_out_2_7, cache_data_out_2_6, cache_data_out_2_5, 
      cache_data_out_2_4, cache_data_out_2_3, cache_data_out_2_2, 
      cache_data_out_2_1, cache_data_out_2_0, cache_data_out_1_15, 
      cache_data_out_1_14, cache_data_out_1_13, cache_data_out_1_12, 
      cache_data_out_1_11, cache_data_out_1_10, cache_data_out_1_9, 
      cache_data_out_1_8, cache_data_out_1_7, cache_data_out_1_6, 
      cache_data_out_1_5, cache_data_out_1_4, cache_data_out_1_3, 
      cache_data_out_1_2, cache_data_out_1_1, cache_data_out_1_0, 
      cache_data_out_0_15, cache_data_out_0_14, cache_data_out_0_13, 
      cache_data_out_0_12, cache_data_out_0_11, cache_data_out_0_10, 
      cache_data_out_0_9, cache_data_out_0_8, cache_data_out_0_7, 
      cache_data_out_0_6, cache_data_out_0_5, cache_data_out_0_4, 
      cache_data_out_0_3, cache_data_out_0_2, cache_data_out_0_1, 
      cache_data_out_0_0, cache_load, cache_rst_actual, 
      comp_unit_flt_size_EXMPLR, max_height_4, max_height_3, max_height_1, 
      comp_unit_operation_EXMPLR, argmax_ready_EXMPLR, 
      filter_ready_out_EXMPLR, comp_unit_relu_EXMPLR, current_state_21, 
      layer_type_out_1, current_state_3, current_state_26, nflt_layer_out_3, 
      current_state_4, nflt_layer_out_1, nflt_layer_out_0, nx78, nx12873, 
      nx92, current_state_8, current_state_7, current_state_6, 
      current_state_5, nx118, current_state_2, nx134, nx140, nx148, nx12875, 
      current_state_24, ftc_cntrl_reg_out_12, current_state_16, 
      ftc_cntrl_reg_out_8, nx12877, nx158, ftc_cntrl_reg_out_14, 
      current_state_10, nx174, nx182, nx196, cntr1_inst_counter_out_1, 
      cntr1_inst_counter_out_0, nx206, cntr1_inst_counter_out_3, 
      cntr1_inst_counter_out_2, nx230, nx244, cntr1_inst_counter_out_4, 
      nx12882, nx262, nx276, nx278, flt_size_out_0, flt_size_out_2, 
      flt_size_out_1, nx308, nx310, nx316, nx330, nx12883, nx336, 
      ftc_cntrl_reg_out_13, nx362, ftc_cntrl_reg_out_11, nx12884, 
      window_width_cntr_counter_out_14, nx12885, 
      window_width_cntr_counter_out_13, window_width_cntr_counter_out_12, 
      nx12887, window_width_cntr_counter_out_11, 
      window_width_cntr_counter_out_10, nx12889, 
      window_width_cntr_counter_out_9, window_width_cntr_counter_out_8, 
      nx12891, window_width_cntr_counter_out_7, 
      window_width_cntr_counter_out_6, nx12893, 
      window_width_cntr_counter_out_5, nx378, nx384, nx392, nx400, nx408, 
      nx428, nx452, nx476, nx500, nx524, nx550, nx564, nx576, 
      img_width_out_0, nx582, new_width_out_0, nx602, nx604, nx612, 
      img_width_out_1, new_width_out_1, nx630, nx636, nx640, img_width_out_2, 
      new_width_out_2, nx674, img_width_out_3, new_width_out_3, nx704, 
      img_width_out_4, new_width_out_4, nx722, nx732, current_state_15, 
      write_offset_data_out_0, nx760, new_size_squared_out_0, 
      write_offset_data_out_1, nx780, new_size_squared_out_1, 
      write_offset_data_out_2, new_size_squared_out_2, 
      write_offset_data_out_3, nx832, new_size_squared_out_3, nx850, 
      write_offset_data_out_4, nx852, nx858, new_size_squared_out_4, 
      write_offset_data_out_5, new_size_squared_out_5, 
      write_offset_data_out_6, nx898, nx904, new_size_squared_out_6, 
      write_offset_data_out_7, new_size_squared_out_7, nx944, 
      write_offset_data_out_8, nx948, nx954, new_size_squared_out_8, 
      write_offset_data_out_9, new_size_squared_out_9, 
      write_offset_data_out_10, nx994, nx1000, new_size_squared_out_10, 
      write_offset_data_out_11, new_size_squared_out_11, nx1040, 
      write_offset_data_out_12, nx1042, nx1048, new_size_squared_out_12, 
      write_offset_data_out_13, new_size_squared_out_13, 
      write_offset_data_out_14, nx1088, nx1094, new_size_squared_out_14, 
      write_offset_data_out_15, new_size_squared_out_15, nx1128, nx1138, 
      ftc_cntrl_reg_out_9, nx1146, nx1154, nx1168, ftc_cntrl_reg_out_10, 
      nx1182, nx1206, nx1212, cache_width_cntr_counter_out_14, nx12896, 
      cache_width_cntr_counter_out_13, cache_width_cntr_counter_out_12, 
      nx12898, cache_width_cntr_counter_out_11, 
      cache_width_cntr_counter_out_10, nx12900, 
      cache_width_cntr_counter_out_9, cache_width_cntr_counter_out_8, 
      nx12902, cache_width_cntr_counter_out_7, 
      cache_width_cntr_counter_out_6, nx12904, nx1224, nx1230, nx1238, 
      nx1246, nx1254, cache_width_cntr_counter_out_5, nx1260, nx1280, nx1304, 
      nx1328, nx1352, nx1376, nx1402, nx1416, nx1434, nx1436, nx1438, nx1446, 
      nx1448, nx1456, nx1460, current_state_19, current_state_18, nx1478, 
      nx1484, nx1500, nx12906, nx1518, nx1524, nx1534, nx1546, 
      num_channels_counter_out_3, nflt_layer_temp_3, 
      num_channels_counter_out_2, nflt_layer_temp_2, nx12908, 
      num_channels_counter_out_1, nflt_layer_temp_1, 
      num_channels_counter_out_0, nflt_layer_temp_0, 
      max_num_channels_data_out_0, nx1608, nx1618, nx1642, nx1648, nx1660, 
      max_num_channels_data_out_2, nx1674, nx1686, 
      max_num_channels_data_out_3, nx1700, nx1712, 
      max_num_channels_data_out_4, nlayers_counter_out_0, nx12910, 
      nlayers_counter_out_2, nlayers_counter_out_1, nx1764, nx1780, nx1796, 
      nx12912, nx1838, nx1876, current_state_27, class_cntr_counter_out_3, 
      class_cntr_counter_out_2, class_cntr_counter_out_1, 
      class_cntr_counter_out_0, nx1904, nx1912, nx1926, nx1938, nx1946, 
      flt_bias_out_0, nx2128, nx2140, nx2142, flt_bias_out_1, nx2168, 
      flt_bias_out_2, nx2194, flt_bias_out_3, nx2220, flt_bias_out_4, nx2246, 
      flt_bias_out_5, nx2272, flt_bias_out_6, nx2298, flt_bias_out_7, nx2324, 
      flt_bias_out_8, nx2350, flt_bias_out_9, nx2376, flt_bias_out_10, 
      nx2402, flt_bias_out_11, nx2428, flt_bias_out_12, nx2454, 
      flt_bias_out_13, nx2480, flt_bias_out_14, nx2506, flt_bias_out_15, 
      nx2532, nx2546, ftc_cntrl_reg_out_15, nx2566, nx2580, nx2622, nx2642, 
      bias_offset_data_out_0, nx2664, nx2668, img_base_addr_0, 
      write_base_prev_data_out_0, nx2674, nx2678, img_addr_offset_0, nx2712, 
      nx2724, nx2738, nx2740, addr1_data_0, nx2754, nx2766, 
      write_base_data_out_1, addr1_data_1, nx2822, img_base_addr_1, 
      write_base_prev_data_out_1, img_addr_offset_1, bias_offset_data_out_1, 
      nx2874, nx2882, nx2892, write_base_data_out_2, nx2914, nx2924, nx2926, 
      nx2928, nx2932, addr1_data_2, nx2942, img_base_addr_2, 
      write_base_prev_data_out_2, nx2968, nx2974, img_addr_offset_2, nx2988, 
      nx2996, bias_offset_data_out_2, nx3016, write_base_data_out_3, nx3048, 
      nx3050, nx3060, nx3074, nx3076, nx3078, addr1_data_3, nx3092, 
      bias_offset_data_out_3, nx3122, img_base_addr_3, 
      write_base_prev_data_out_3, nx3146, img_addr_offset_3, nx3160, nx3168, 
      write_base_data_out_4, nx3206, addr1_data_4, nx3232, nx3238, nx3246, 
      img_base_addr_4, nx3264, nx3270, img_addr_offset_4, nx3278, nx3284, 
      nx3292, bias_offset_data_out_4, nx3312, write_base_data_out_5, nx3346, 
      nx3356, nx3360, nx3370, addr1_data_5, img_base_addr_5, 
      write_base_prev_data_out_5, nx3412, img_addr_offset_5, nx3434, 
      bias_offset_data_out_5, nx3454, nx3458, write_base_data_out_6, 
      addr1_data_6, nx3516, nx3522, nx3532, img_base_addr_6, nx3548, nx3554, 
      img_addr_offset_6, nx3562, nx3568, bias_offset_data_out_6, nx3608, 
      write_base_data_out_7, nx3630, nx3640, nx3654, addr1_data_7, 
      img_base_addr_7, write_base_prev_data_out_7, nx3696, img_addr_offset_7, 
      nx3718, bias_offset_data_out_7, nx3738, nx3742, write_base_data_out_8, 
      nx3780, addr1_data_8, nx3800, nx3806, nx3816, img_base_addr_8, nx3832, 
      nx3838, img_addr_offset_8, nx3846, nx3852, bias_offset_data_out_8, 
      nx3892, write_base_data_out_9, nx3914, nx3924, nx3938, addr1_data_9, 
      img_base_addr_9, write_base_prev_data_out_9, nx3980, img_addr_offset_9, 
      nx4002, bias_offset_data_out_9, nx4022, nx4026, nx4044, 
      write_base_data_out_10, addr1_data_10, nx4084, nx4090, nx4100, 
      img_base_addr_10, nx4116, nx4122, img_addr_offset_10, nx4130, nx4136, 
      bias_offset_data_out_10, nx4176, write_base_data_out_11, nx4198, 
      nx4208, nx4222, addr1_data_11, img_base_addr_11, 
      write_base_prev_data_out_11, nx4264, img_addr_offset_11, nx4286, 
      bias_offset_data_out_11, nx4306, write_base_data_out_12, addr1_data_12, 
      nx4368, nx4374, img_base_addr_12, nx4400, nx4406, img_addr_offset_12, 
      nx4414, nx4420, bias_offset_data_out_12, write_base_data_out_13, 
      nx4492, nx4506, addr1_data_13, nx4534, img_base_addr_13, 
      write_base_prev_data_out_13, nx4548, img_addr_offset_13, nx4568, 
      nx4570, bias_offset_data_out_13, nx4590, nx4594, 
      write_base_data_out_14, addr1_data_14, nx4652, nx4658, nx4668, 
      img_base_addr_14, nx4684, nx4690, img_addr_offset_14, nx4698, nx4704, 
      bias_offset_data_out_14, nx4744, nx4754, bias_offset_data_out_15, 
      write_base_data_out_15, nx4782, addr1_data_15, nx4802, nx4804, nx4812, 
      nx4816, nx4826, img_base_addr_15, write_base_prev_data_out_15, nx4834, 
      nx4850, nx12921, nx12931, nx12941, nx12951, nx12961, nx12971, nx12981, 
      nx12991, nx13001, nx13011, nx13021, nx13031, nx13041, nx13051, nx13061, 
      nx13071, nx13081, nx13091, nx13101, nx13111, nx13121, nx13131, nx13141, 
      nx13151, nx13161, nx13171, nx13181, nx13191, nx13201, nx13211, nx13221, 
      nx13231, nx13241, nx13251, nx13261, nx13271, nx13281, nx13291, nx13301, 
      nx13311, nx13321, nx13331, nx13341, nx13351, nx13361, nx13371, nx13381, 
      nx13391, nx13401, nx13411, nx13421, nx13431, nx13441, nx13451, nx13461, 
      nx13471, nx13481, nx13491, nx13501, nx13511, nx13521, nx13531, nx13541, 
      nx13551, nx13561, nx13571, nx13581, nx13591, nx13601, nx13611, nx13621, 
      nx13631, nx13641, nx13651, nx13661, nx13671, nx13681, nx13691, nx13701, 
      nx13711, nx13721, nx13731, nx13741, nx13751, nx13761, nx13771, nx13781, 
      nx13791, nx13801, nx13811, nx13821, nx13831, nx13841, nx13851, nx13861, 
      nx13871, nx13881, nx13891, nx13901, nx13911, nx13921, nx13931, nx13941, 
      nx13951, nx13961, nx13971, nx13981, nx13991, nx14001, nx14011, nx14021, 
      nx14031, nx14041, nx14051, nx14061, nx14071, nx14081, nx14091, nx14101, 
      nx14111, nx14121, nx14131, nx14141, nx14151, nx14161, nx14171, nx14181, 
      nx14191, nx14201, nx14211, nx14221, nx14231, nx14241, nx14251, nx14261, 
      nx14271, nx14281, nx14291, nx14301, nx14311, nx14321, nx14331, nx14341, 
      nx14351, nx14361, nx14371, nx14381, nx14391, nx14401, nx14411, nx14421, 
      nx14431, nx14441, nx14451, nx14461, nx14471, nx14481, nx14491, nx14501, 
      nx14511, nx14521, nx14531, nx14541, nx14551, nx14561, nx14571, nx14581, 
      nx14591, nx14601, nx14611, nx14621, nx14631, nx14641, nx14651, nx14661, 
      nx14671, nx14681, nx14691, nx14701, nx14711, nx14721, nx14731, nx14741, 
      nx14751, nx14761, nx14771, nx14781, nx14791, nx14801, nx14811, nx14821, 
      nx14831, nx14841, nx14851, nx14861, nx14871, nx14881, nx14891, nx14901, 
      nx14911, nx14921, nx14931, nx14941, nx14951, nx14961, nx14971, nx14981, 
      nx14991, nx15001, nx15011, nx15021, nx15031, nx15041, nx15051, nx15061, 
      nx15071, nx15081, nx15091, nx15101, nx15111, nx15121, nx15131, nx15141, 
      nx15161, nx15171, nx15181, nx15191, nx15201, nx15221, nx15231, nx15241, 
      nx15251, nx15261, nx15281, nx15291, nx15301, nx15311, nx15321, nx15331, 
      nx15351, nx15361, nx15371, nx15381, nx15392, nx15396, nx15402, nx15407, 
      nx15412, nx15416, nx15422, nx15426, nx15428, nx15432, nx15435, nx15445, 
      nx15450, nx15452, nx15460, nx15466, nx15470, nx15474, nx15479, nx15486, 
      nx15488, nx15491, nx15496, nx15500, nx15502, nx15504, nx15506, nx15508, 
      nx15512, nx15514, nx15516, nx15518, nx15523, nx15525, nx15527, nx15530, 
      nx15531, nx15533, nx15537, nx15541, nx15544, nx15546, nx15548, nx15554, 
      nx15559, nx15561, nx15563, nx15567, nx15571, nx15573, nx15575, nx15580, 
      nx15586, nx15588, nx15591, nx15596, nx15598, nx15602, nx15605, nx15609, 
      nx15614, nx15617, nx15619, nx15621, nx15626, nx15630, nx15635, nx15637, 
      nx15640, nx15644, nx15647, nx15653, nx15657, nx15660, nx15666, nx15670, 
      nx15673, nx15679, nx15683, nx15686, nx15692, nx15696, nx15711, nx15716, 
      nx15717, nx15720, nx15726, nx15730, nx15732, nx15735, nx15741, nx15745, 
      nx15750, nx15753, nx15756, nx15759, nx15763, nx15765, nx15768, nx15770, 
      nx15772, nx15774, nx15776, nx15781, nx15785, nx15786, nx15791, nx15795, 
      nx15797, nx15802, nx15806, nx15807, nx15812, nx15816, nx15818, nx15823, 
      nx15827, nx15828, nx15833, nx15837, nx15839, nx15844, nx15848, nx15849, 
      nx15854, nx15859, nx15861, nx15865, nx15868, nx15873, nx15876, nx15878, 
      nx15883, nx15885, nx15888, nx15890, nx15893, nx15898, nx15902, nx15904, 
      nx15907, nx15912, nx15916, nx15918, nx15921, nx15926, nx15930, nx15932, 
      nx15935, nx15940, nx15944, nx15946, nx15949, nx15954, nx15959, nx15970, 
      nx15974, nx15983, nx15989, nx15995, nx15997, nx16005, nx16013, nx16019, 
      nx16025, nx16028, nx16037, nx16039, nx16042, nx16046, nx16052, nx16055, 
      nx16063, nx16065, nx16067, nx16070, nx16075, nx16079, nx16081, nx16084, 
      nx16089, nx16093, nx16095, nx16098, nx16103, nx16107, nx16109, nx16112, 
      nx16117, nx16121, nx16123, nx16126, nx16131, nx16136, nx16148, nx16150, 
      nx16153, nx16155, nx16166, nx16172, nx16178, nx16180, nx16189, nx16191, 
      nx16196, nx16198, nx16202, nx16204, nx16213, nx16216, nx16222, nx16224, 
      nx16226, nx16228, nx16234, nx16239, nx16243, nx16247, nx16253, nx16258, 
      nx16262, nx16265, nx16269, nx16274, nx16278, nx16280, nx16282, nx16284, 
      nx16290, nx16299, nx16302, nx16305, nx16307, nx16313, nx16318, nx16324, 
      nx16327, nx16332, nx16334, nx16336, nx16338, nx16346, nx16348, nx16373, 
      nx16455, nx16459, nx16463, nx16507, nx16511, nx16514, nx16518, nx16521, 
      nx16524, nx16527, nx16530, nx16533, nx16536, nx16539, nx16542, nx16545, 
      nx16548, nx16551, nx16554, nx16557, nx16560, nx16563, nx16566, nx16569, 
      nx16572, nx16575, nx16578, nx16581, nx16584, nx16587, nx16590, nx16593, 
      nx16596, nx16599, nx16602, nx16605, nx16608, nx16610, nx16629, nx16715, 
      nx16721, nx16727, nx16729, nx16732, nx16736, nx16738, nx16742, nx16745, 
      nx16747, nx16756, nx16764, nx16768, nx16770, nx16774, nx16776, nx16780, 
      nx16786, nx16788, nx16791, nx16796, nx16798, nx16802, nx16804, nx16806, 
      nx16810, nx16812, nx16818, nx16820, nx16825, nx16829, nx16831, nx16833, 
      nx16835, nx16837, nx16839, nx16843, nx16846, nx16849, nx16852, nx16857, 
      nx16861, nx16863, nx16868, nx16870, nx16874, nx16878, nx16880, nx16895, 
      nx16906, nx16911, nx16915, nx16916, nx16924, nx16927, nx16931, nx16934, 
      nx16943, nx16945, nx16948, nx16956, nx16962, nx16967, nx16973, nx16976, 
      nx16978, nx16983, nx16993, nx17002, nx17004, nx17021, nx17031, nx17035, 
      nx17038, nx17042, nx17044, nx17047, nx17051, nx17054, nx17056, nx17060, 
      nx17065, nx17074, nx17076, nx17077, nx17081, nx17085, nx17089, nx17100, 
      nx17102, nx17104, nx17106, nx17110, nx17112, nx17114, nx17125, nx17135, 
      nx17138, nx17140, nx17147, nx17157, nx17161, nx17164, nx17168, nx17175, 
      nx17178, nx17183, nx17186, nx17188, nx17194, nx17199, nx17204, nx17210, 
      nx17214, nx17218, nx17229, nx17231, nx17233, nx17235, nx17239, nx17242, 
      nx17244, nx17255, nx17265, nx17268, nx17270, nx17277, nx17287, nx17291, 
      nx17294, nx17298, nx17307, nx17310, nx17312, nx17315, nx17321, nx17326, 
      nx17331, nx17337, nx17341, nx17345, nx17356, nx17358, nx17360, nx17362, 
      nx17366, nx17369, nx17371, nx17374, nx17377, nx17382, nx17392, nx17395, 
      nx17397, nx17404, nx17414, nx17418, nx17421, nx17425, nx17434, nx17437, 
      nx17439, nx17442, nx17448, nx17453, nx17458, nx17464, nx17468, nx17472, 
      nx17483, nx17485, nx17487, nx17489, nx17493, nx17496, nx17498, nx17509, 
      nx17519, nx17522, nx17541, nx17545, nx17548, nx17552, nx17561, nx17564, 
      nx17566, nx17575, nx17580, nx17591, nx17595, nx17599, nx17610, nx17612, 
      nx17614, nx17616, nx17620, nx17623, nx17625, nx17636, nx17641, nx17646, 
      nx17649, nx17658, nx17660, nx17663, nx17670, nx17671, nx17673, nx17677, 
      nx17679, nx17682, nx17685, nx17687, nx17692, nx17696, nx17700, nx17711, 
      nx17723, nx17726, nx17728, nx17737, nx17740, nx17744, nx17748, nx17751, 
      nx17754, nx17757, nx17760, nx17763, nx17766, nx17769, nx17772, nx17775, 
      nx17778, nx17781, nx17784, nx17787, nx17790, nx17793, nx17796, nx17803, 
      nx17805, nx17807, nx17809, nx17811, nx17813, nx17815, nx17817, nx17819, 
      nx17821, nx17823, nx17825, nx17827, nx17829, nx17831, nx17833, nx17835, 
      nx17837, nx17839, nx17841, nx17843, nx17845, nx17847, nx17855, nx17857, 
      nx17859, nx17863, nx17865, nx17869, nx17871, nx17873, nx17875, nx17877, 
      nx17879, nx17887, nx17893, nx17895, nx17897, nx17899, nx17907, nx17909, 
      nx17911, nx17913, nx17915, nx17917, nx17919, nx17921, nx17923, nx17927, 
      nx17929, nx17937, nx17939, nx17941, nx17943, nx17945, nx17947, nx17949, 
      nx17951, nx17959, nx17961, nx17963, nx17965, nx17971, nx17973, nx17975, 
      nx17979, nx17981, nx17983, nx17993, nx17995, nx17997, nx17999, nx18001, 
      nx18003, nx18005, nx18007, nx18011, nx18017, nx18021, nx18023, nx18027, 
      nx18029, nx18031, nx18033, nx18035, nx18037, nx18039, nx18041, nx18045, 
      nx18047, nx18049, nx18051, nx18053, nx18055, nx18059, nx18063, nx18065, 
      nx18067, nx18069, nx18077, nx18081, nx18085, nx18087, nx18089, nx18091, 
      nx18117, nx18119, nx18121, nx18137, nx18139, nx18141, nx18143, nx18151, 
      nx18153, nx18155, nx18157, nx18163, nx18165, nx18167, nx18169, nx18171, 
      nx18173, nx18175, nx18177, nx18179, nx18181, nx18183, nx18185, nx18187, 
      nx18189, nx18191, nx18193, nx18195, nx18197, nx18199, nx18201, nx18203, 
      nx18205, nx18207, nx18211, nx18217, nx18219, nx18225, nx18227, nx18229, 
      nx18231, nx18233, nx18235, nx18237, nx18239, nx18241, nx18243, nx18245, 
      nx18247, nx18249, nx18251, nx18253, nx18255, nx18257, nx18259, nx18261, 
      nx18263, nx18265, nx18269, nx18271, nx18273, nx18275, nx18277, nx18279, 
      nx18281, nx18283, nx18285, nx18287, nx18289, nx18291, nx18293, nx18295, 
      nx18297, nx18299, nx18301, nx18303, nx18305, nx18307, nx18309, nx18311, 
      nx18313, nx18315, nx18317, nx18319, nx18321, nx18323, nx18325, nx18327, 
      nx18329, nx18331, nx18333, nx18335, nx18339, nx18341, nx18343, nx18345, 
      nx18347, nx18349, nx18351, nx18353, nx18355, nx18357, nx18359, nx18361, 
      nx18363, nx18365, nx18367, nx18369, nx18371, nx18373, nx18375, nx18381, 
      nx18383, nx18385, nx17067, nx3366, nx16995, nx18543, nx18544, nx18545, 
      nx18546, nx18547, nx18548, nx18549, nx18550, nx18551, nx18552, nx18553, 
      nx15341, nx18554, nx18555, nx18556, nx18557, nx18558, nx18559, nx18560, 
      nx18561, nx18562, nx18009, nx18563, nx18564, nx18565, nx18566, nx18567, 
      nx18568, nx3046, nx16882, nx16885, nx16808, nx18569, nx18570, nx18571, 
      nx18572, nx18573, nx18574, nx18575, NOT_nx4768, nx18576, nx18577, 
      nx18578, nx18579, nx16888, nx18580, nx18581, nx18582, nx18583, nx18584, 
      nx18585, nx3444, nx18586, nx18587, nx17013, nx18588, nx17016, nx3112, 
      nx16891, nx18589, nx18590, nx16987, nx18591, nx18592, nx18593, nx18594, 
      nx18595, nx18596, nx18597, nx18598, nx18599, nx17118, nx18600, nx18601, 
      nx17121, nx3184, nx18602, nx18603, nx16990, nx18604, nx17656, nx18605, 
      nx18223, nx18606, nx18607, nx18608, nx18609, nx18610, nx18043, nx18611, 
      nx18612, nx18613, nx18614, nx18615, nx15271, nx18616, nx18617, nx18618, 
      nx18619, nx18620, nx18621, nx18622, nx18623, nx18624, nx18625, nx4612, 
      nx18626, nx17731, nx18627, nx18628, nx18629, nx17629, nx18630, nx18631, 
      nx17632, nx4328, nx18632, nx17502, nx17505, nx17529, nx18633, nx18634, 
      nx18635, nx18636, nx15151, nx18267, nx18337, nx18637, nx18638, nx18639, 
      nx18640, nx18641, nx18642, nx18643, nx18644, nx18645, nx18646, nx17023, 
      nx18647, nx3132, nx18648, nx16898, nx18649, nx16901, nx16814, nx18650, 
      nx18651, nx18652, nx18653, nx18654, nx18655, nx18656, nx18657, nx18658, 
      nx17127, nx18659, nx18660, nx18661, nx18662, nx18663, nx18664, nx18665, 
      nx18666, nx18667, nx18668, nx18669, nx18670, nx18671, nx18672, nx18673, 
      nx15211, nx17585, nx18674, nx18675, nx18676, nx18677, nx18678, nx17526, 
      nx18679, nx18680, nx17402, nx18681, nx18682, nx18683, nx18684, nx18685, 
      nx18686, nx18687, nx18688, nx4194, nx18689, nx18690, nx18691, nx18692, 
      nx17399, nx18693, nx18694, nx18695, nx18696, nx17272, nx18697, nx18698, 
      nx17275, nx3626, nx18699, nx18700, nx17145, nx18701, nx18702, nx18703, 
      nx18704, nx18705, nx18706, nx18707, nx18708, nx18709, nx18710, nx18711, 
      nx4502, nx18712, nx18713, nx18714, nx18715, nx18716, nx17556, nx4218, 
      nx17429, nx4168, nx18717, nx18718, nx18719, nx18720, nx18721, nx18722, 
      nx18723, nx18724, nx17638, nx18725, nx18726, nx18727, nx18728, nx18729, 
      nx18730, nx17511, nx18731, nx17514, nx4296, nx18732, nx18733, nx17384, 
      nx17387, nx18734, nx18735, nx18736, nx18737, nx18738, nx18739, nx18740, 
      nx18741, nx18742, NOT_nx3476, nx18743, nx18744, nx18745, nx18746, 
      nx18747, nx18748, nx18749, nx18750, nx3682, nx18751, nx18752, nx18753, 
      nx18754, nx18755, nx18756, nx3966, nx18757, nx18758, nx17279, nx18759, 
      nx17282, nx18760, nx18761, nx18762, nx17149, nx18763, nx17152, nx3398, 
      nx17026, nx18764, nx18765, nx18766, nx18767, nx18768, nx18769, nx3342, 
      nx18770, nx18771, nx17006, nx18772, nx18773, nx17009, nx18774, nx18775, 
      nx18776, nx18777, nx18778, nx18779, nx18780, nx4496, nx18781, nx17431, 
      nx18782, nx18783, nx18784, nx18785, nx18786, nx18787, nx18788, nx17323, 
      nx18789, nx18790, nx3934, nx18791, nx18792, nx3644, nx18793, nx18794, 
      nx18795, nx17196, nx3884, nx3928, nx17302, nx3650, nx17172, nx3600, 
      nx18796, nx18797, nx18798, nx18799, nx18800, nx18801, nx18802, nx18803, 
      nx18804, nx18805, nx18806, nx18807, NOT_nx3910, nx18808, nx18809, 
      nx18810, nx18811, nx18812, nx18813, nx18814, nx18815, nx18816, nx17531, 
      nx18817, nx17571, nx18818, nx18819, nx18820, nx18135, nx18821, nx18822, 
      nx18075, nx17536, nx18823, nx18824, nx18213, nx17977, nx4250, nx17450, 
      nx18825, nx17409, nx18826, nx18827, nx18828, nx18829, nx18830, nx18831, 
      nx18832, nx17247, nx17250, nx18833, nx18834, nx18835, nx18836, nx18837, 
      nx18838, nx17533, nx18839, nx17406, nx18840, nx18841, nx18842, nx18843, 
      nx3760, nx17577, nx4736, nx18844, nx18845, nx18846, nx18847, nx17257, 
      nx3728, nx17130, nx18848, nx18849, nx18850, nx18851, nx18852, nx18853, 
      nx18854, nx18855, nx4012, nx18856, nx18857, nx18858, nx17260, nx18859, 
      nx18860, nx18861, nx18862, nx18863, nx18864, nx18865, nx18866, nx16998, 
      nx18867, nx18868, nx3216, nx16937, nx18869, nx18870, nx18871, nx18872, 
      nx18873, nx18874, nx4580, nx18875, nx18876, nx18877, nx18878, nx18879, 
      nx18880, nx17142, nx18881, nx18882, nx18883, nx18884, nx18885, nx18886, 
      nx18887, nx18888, nx18889, nx18890, nx18891, nx18892, nx18893, nx18894, 
      nx18895, nx18896, nx18897, nx18898, nx18899, nx18900, nx18901, nx18902, 
      nx18903, nx18904, nx18905, nx18906, nx18907, nx18908, nx18909, nx18910, 
      nx18911, nx18912, nx18913, nx18914, nx18915, nx18916, nx19292, nx19294, 
      nx19296, nx19298, nx19300, nx19302, nx19308: std_logic ;
   
   signal DANGLING : std_logic_vector (15 downto 0 );

begin
   io_done_out <= comp_unit_relu_EXMPLR ;
   wind_rst <= comp_unit_relu_EXMPLR ;
   filter_ready_out <= filter_ready_out_EXMPLR ;
   filter_reset <= reset ;
   comp_unit_operation <= comp_unit_operation_EXMPLR ;
   comp_unit_flt_size <= comp_unit_flt_size_EXMPLR ;
   comp_unit_relu <= comp_unit_relu_EXMPLR ;
   argmax_ready <= argmax_ready_EXMPLR ;
   img_cache : Cache_5_16_28_5 port map ( in_word(15)=>cache_data_in_15, 
      in_word(14)=>cache_data_in_14, in_word(13)=>cache_data_in_13, 
      in_word(12)=>cache_data_in_12, in_word(11)=>cache_data_in_11, 
      in_word(10)=>cache_data_in_10, in_word(9)=>cache_data_in_9, in_word(8)
      =>cache_data_in_8, in_word(7)=>cache_data_in_7, in_word(6)=>
      cache_data_in_6, in_word(5)=>cache_data_in_5, in_word(4)=>
      cache_data_in_4, in_word(3)=>cache_data_in_3, in_word(2)=>
      cache_data_in_2, in_word(1)=>cache_data_in_1, in_word(0)=>
      cache_data_in_0, cache_in_sel(4)=>nx17815, cache_in_sel(3)=>
      cache_width_count_3, cache_in_sel(2)=>nx17819, cache_in_sel(1)=>
      cache_width_count_1, cache_in_sel(0)=>cache_width_count_0, 
      cache_out_sel(4)=>wind_width_count_4, cache_out_sel(3)=>
      wind_width_count_3, cache_out_sel(2)=>wind_width_count_2, 
      cache_out_sel(1)=>wind_width_count_1, cache_out_sel(0)=>nx17811, 
      decoder_enable=>cache_load, out_column_0_15=>cache_data_out_4_15, 
      out_column_0_14=>cache_data_out_4_14, out_column_0_13=>
      cache_data_out_4_13, out_column_0_12=>cache_data_out_4_12, 
      out_column_0_11=>cache_data_out_4_11, out_column_0_10=>
      cache_data_out_4_10, out_column_0_9=>cache_data_out_4_9, 
      out_column_0_8=>cache_data_out_4_8, out_column_0_7=>cache_data_out_4_7, 
      out_column_0_6=>cache_data_out_4_6, out_column_0_5=>cache_data_out_4_5, 
      out_column_0_4=>cache_data_out_4_4, out_column_0_3=>cache_data_out_4_3, 
      out_column_0_2=>cache_data_out_4_2, out_column_0_1=>cache_data_out_4_1, 
      out_column_0_0=>cache_data_out_4_0, out_column_1_15=>
      cache_data_out_3_15, out_column_1_14=>cache_data_out_3_14, 
      out_column_1_13=>cache_data_out_3_13, out_column_1_12=>
      cache_data_out_3_12, out_column_1_11=>cache_data_out_3_11, 
      out_column_1_10=>cache_data_out_3_10, out_column_1_9=>
      cache_data_out_3_9, out_column_1_8=>cache_data_out_3_8, out_column_1_7
      =>cache_data_out_3_7, out_column_1_6=>cache_data_out_3_6, 
      out_column_1_5=>cache_data_out_3_5, out_column_1_4=>cache_data_out_3_4, 
      out_column_1_3=>cache_data_out_3_3, out_column_1_2=>cache_data_out_3_2, 
      out_column_1_1=>cache_data_out_3_1, out_column_1_0=>cache_data_out_3_0, 
      out_column_2_15=>cache_data_out_2_15, out_column_2_14=>
      cache_data_out_2_14, out_column_2_13=>cache_data_out_2_13, 
      out_column_2_12=>cache_data_out_2_12, out_column_2_11=>
      cache_data_out_2_11, out_column_2_10=>cache_data_out_2_10, 
      out_column_2_9=>cache_data_out_2_9, out_column_2_8=>cache_data_out_2_8, 
      out_column_2_7=>cache_data_out_2_7, out_column_2_6=>cache_data_out_2_6, 
      out_column_2_5=>cache_data_out_2_5, out_column_2_4=>cache_data_out_2_4, 
      out_column_2_3=>cache_data_out_2_3, out_column_2_2=>cache_data_out_2_2, 
      out_column_2_1=>cache_data_out_2_1, out_column_2_0=>cache_data_out_2_0, 
      out_column_3_15=>cache_data_out_1_15, out_column_3_14=>
      cache_data_out_1_14, out_column_3_13=>cache_data_out_1_13, 
      out_column_3_12=>cache_data_out_1_12, out_column_3_11=>
      cache_data_out_1_11, out_column_3_10=>cache_data_out_1_10, 
      out_column_3_9=>cache_data_out_1_9, out_column_3_8=>cache_data_out_1_8, 
      out_column_3_7=>cache_data_out_1_7, out_column_3_6=>cache_data_out_1_6, 
      out_column_3_5=>cache_data_out_1_5, out_column_3_4=>cache_data_out_1_4, 
      out_column_3_3=>cache_data_out_1_3, out_column_3_2=>cache_data_out_1_2, 
      out_column_3_1=>cache_data_out_1_1, out_column_3_0=>cache_data_out_1_0, 
      out_column_4_15=>cache_data_out_0_15, out_column_4_14=>
      cache_data_out_0_14, out_column_4_13=>cache_data_out_0_13, 
      out_column_4_12=>cache_data_out_0_12, out_column_4_11=>
      cache_data_out_0_11, out_column_4_10=>cache_data_out_0_10, 
      out_column_4_9=>cache_data_out_0_9, out_column_4_8=>cache_data_out_0_8, 
      out_column_4_7=>cache_data_out_0_7, out_column_4_6=>cache_data_out_0_6, 
      out_column_4_5=>cache_data_out_0_5, out_column_4_4=>cache_data_out_0_4, 
      out_column_4_3=>cache_data_out_0_3, out_column_4_2=>cache_data_out_0_2, 
      out_column_4_1=>cache_data_out_0_1, out_column_4_0=>cache_data_out_0_0, 
      clk=>nx17823, reset=>cache_rst_actual);
   cache_height_cntr : AdvancedCounter_16 port map ( clk=>clk, reset=>
      nx17805, enable=>cache_height_count_en, mode_in(1)=>
      comp_unit_relu_EXMPLR, mode_in(0)=>comp_unit_relu_EXMPLR, 
      max_val_in(15)=>comp_unit_relu_EXMPLR, max_val_in(14)=>
      comp_unit_relu_EXMPLR, max_val_in(13)=>comp_unit_relu_EXMPLR, 
      max_val_in(12)=>comp_unit_relu_EXMPLR, max_val_in(11)=>
      comp_unit_relu_EXMPLR, max_val_in(10)=>comp_unit_relu_EXMPLR, 
      max_val_in(9)=>comp_unit_relu_EXMPLR, max_val_in(8)=>
      comp_unit_relu_EXMPLR, max_val_in(7)=>comp_unit_relu_EXMPLR, 
      max_val_in(6)=>comp_unit_relu_EXMPLR, max_val_in(5)=>
      comp_unit_relu_EXMPLR, max_val_in(4)=>max_height_4, max_val_in(3)=>
      max_height_3, max_val_in(2)=>max_height_2, max_val_in(1)=>max_height_1, 
      max_val_in(0)=>max_height_0, max_reached_out=>cache_height_ended, 
      counter_out(15)=>DANGLING(0), counter_out(14)=>DANGLING(1), 
      counter_out(13)=>DANGLING(2), counter_out(12)=>DANGLING(3), 
      counter_out(11)=>DANGLING(4), counter_out(10)=>DANGLING(5), 
      counter_out(9)=>DANGLING(6), counter_out(8)=>DANGLING(7), 
      counter_out(7)=>DANGLING(8), counter_out(6)=>DANGLING(9), 
      counter_out(5)=>DANGLING(10), counter_out(4)=>DANGLING(11), 
      counter_out(3)=>DANGLING(12), counter_out(2)=>DANGLING(13), 
      counter_out(1)=>DANGLING(14), counter_out(0)=>DANGLING(15));
   ix12710 : fake_gnd port map ( Y=>comp_unit_relu_EXMPLR);
   ix321 : oai21 port map ( Y=>filter_ready_out_EXMPLR, A0=>nx18255, A1=>
      nx15396, B0=>nx16313);
   reg_current_state_11 : dffr port map ( Q=>OPEN, QB=>nx15392, D=>nx17865, 
      CLK=>nx17823, R=>reset);
   ix15403 : nand04 port map ( Y=>nx15402, A0=>cntr1_inst_counter_out_3, A1
      =>cntr1_inst_counter_out_2, A2=>cntr1_inst_counter_out_1, A3=>
      cntr1_inst_counter_out_0);
   reg_cntr1_inst_counter_out_3 : dffr port map ( Q=>
      cntr1_inst_counter_out_3, QB=>OPEN, D=>nx13001, CLK=>clk, R=>nx17929);
   ix245 : xnor2 port map ( Y=>nx244, A0=>cntr1_inst_counter_out_3, A1=>
      nx15407);
   ix15408 : nand03 port map ( Y=>nx15407, A0=>cntr1_inst_counter_out_2, A1
      =>cntr1_inst_counter_out_1, A2=>cntr1_inst_counter_out_0);
   reg_cntr1_inst_counter_out_2 : dffr port map ( Q=>
      cntr1_inst_counter_out_2, QB=>OPEN, D=>nx12991, CLK=>clk, R=>nx17929);
   ix231 : xnor2 port map ( Y=>nx230, A0=>cntr1_inst_counter_out_2, A1=>
      nx15412);
   ix15413 : nand02 port map ( Y=>nx15412, A0=>cntr1_inst_counter_out_1, A1
      =>cntr1_inst_counter_out_0);
   reg_cntr1_inst_counter_out_1 : dffr port map ( Q=>
      cntr1_inst_counter_out_1, QB=>nx15416, D=>nx12981, CLK=>clk, R=>
      nx17929);
   ix183 : oai21 port map ( Y=>nx182, A0=>nx15422, A1=>nx15537, B0=>nx16302
   );
   ix13992 : mux21 port map ( Y=>nx13991, A0=>nx15426, A1=>nx15428, S0=>
      nx17973);
   num_channels_counter_out_4 : dffr port map ( Q=>OPEN, QB=>nx15426, D=>
      nx13991, CLK=>clk, R=>reset);
   ix15429 : aoi222 port map ( Y=>nx15428, A0=>max_num_channels_data_out_4, 
      A1=>nx1642, B0=>mem_data_in(4), B1=>nx17899, C0=>nx18271, C1=>nx1712);
   ix13982 : oai22 port map ( Y=>nx13981, A0=>nx15432, A1=>nx582, B0=>
      nx16299, B1=>nx15435);
   max_num_channels_inst_reg_q_4 : dffr port map ( Q=>
      max_num_channels_data_out_4, QB=>nx15432, D=>nx13981, CLK=>clk, R=>
      reset);
   ix119 : and02 port map ( Y=>nx118, A0=>current_state_8, A1=>nx15546);
   reg_current_state_8 : dffr port map ( Q=>current_state_8, QB=>OPEN, D=>
      nx17907, CLK=>nx17837, R=>reset);
   reg_current_state_7 : dffr port map ( Q=>current_state_7, QB=>OPEN, D=>
      current_state_6, CLK=>nx17835, R=>reset);
   reg_current_state_6 : dffr port map ( Q=>current_state_6, QB=>OPEN, D=>
      current_state_5, CLK=>nx17835, R=>reset);
   reg_current_state_5 : dffr port map ( Q=>current_state_5, QB=>OPEN, D=>
      nx17895, CLK=>nx17835, R=>reset);
   reg_current_state_4 : dffr port map ( Q=>current_state_4, QB=>OPEN, D=>
      current_state_3, CLK=>nx17835, R=>reset);
   reg_current_state_3 : dffr port map ( Q=>current_state_3, QB=>OPEN, D=>
      nx12910, CLK=>nx17835, R=>reset);
   reg_current_state_2 : dffr port map ( Q=>current_state_2, QB=>nx15445, D
      =>nx140, CLK=>nx17823, R=>reset);
   ix135 : oai21 port map ( Y=>nx134, A0=>io_ready_in, A1=>nx15450, B0=>
      nx15452);
   reg_current_state_1 : dffr port map ( Q=>OPEN, QB=>nx15450, D=>nx134, CLK
      =>nx17823, R=>reset);
   reg_current_state_0 : dffs_ni port map ( Q=>OPEN, QB=>nx15452, D=>
      comp_unit_relu_EXMPLR, CLK=>nx17823, S=>reset);
   ix1733 : nand02 port map ( Y=>nx12875, A0=>nx15460, A1=>nx15426);
   ix15461 : nor04 port map ( Y=>nx15460, A0=>num_channels_counter_out_0, A1
      =>num_channels_counter_out_1, A2=>num_channels_counter_out_2, A3=>
      num_channels_counter_out_3);
   ix13912 : mux21_ni port map ( Y=>nx13911, A0=>num_channels_counter_out_0, 
      A1=>nx1618, S0=>nx17973);
   ix1619 : mux21_ni port map ( Y=>nx1618, A0=>nx1608, A1=>nx15531, S0=>
      nx18269);
   ix1609 : nand03 port map ( Y=>nx1608, A0=>nx15466, A1=>nx15474, A2=>
      nx15445);
   ix15467 : oai21 port map ( Y=>nx15466, A0=>max_num_channels_data_out_0, 
      A1=>nx18151, B0=>nx17887);
   ix13902 : oai32 port map ( Y=>nx13901, A0=>nx15470, A1=>nx17897, A2=>
      nx17875, B0=>nx15474, B1=>nx18259);
   max_num_channels_inst_reg_q_0 : dffr port map ( Q=>
      max_num_channels_data_out_0, QB=>nx15470, D=>nx13901, CLK=>clk, R=>
      reset);
   reg_current_state_9 : dffr port map ( Q=>OPEN, QB=>nx15435, D=>nx118, CLK
      =>nx17823, R=>reset);
   reg_current_state_26 : dffr port map ( Q=>current_state_26, QB=>OPEN, D=>
      nx1796, CLK=>nx17823, R=>reset);
   ix15475 : aoi22 port map ( Y=>nx15474, A0=>mem_data_in(0), A1=>nx17897, 
      B0=>nx17875, B1=>nflt_layer_temp_0);
   nflt_layer_total_reg_q_0 : dffr port map ( Q=>nflt_layer_temp_0, QB=>OPEN, 
      D=>nx13891, CLK=>clk, R=>reset);
   ix13892 : mux21_ni port map ( Y=>nx13891, A0=>nflt_layer_temp_0, A1=>
      mem_data_in(0), S0=>nx17893);
   layer_type_reg_q_0 : dffr port map ( Q=>comp_unit_operation_EXMPLR, QB=>
      OPEN, D=>nx12961, CLK=>clk, R=>reset);
   ix12962 : mux21_ni port map ( Y=>nx12961, A0=>nx18151, A1=>mem_data_in(0), 
      S0=>current_state_3);
   reg_current_state_25 : dffr port map ( Q=>OPEN, QB=>nx15530, D=>nx92, CLK
      =>nx17825, R=>reset);
   ix12922 : oai32 port map ( Y=>nx12921, A0=>nx15488, A1=>nx17893, A2=>
      nx17887, B0=>nx15491, B1=>nx18263);
   reg_nflt_layer_out_0 : dffr port map ( Q=>nflt_layer_out_0, QB=>nx15488, 
      D=>nx12921, CLK=>clk, R=>reset);
   ix12932 : oai32 port map ( Y=>nx12931, A0=>nx15500, A1=>nx17893, A2=>
      nx17887, B0=>nx15502, B1=>nx18263);
   reg_nflt_layer_out_1 : dffr port map ( Q=>nflt_layer_out_1, QB=>nx15500, 
      D=>nx12931, CLK=>clk, R=>reset);
   ix15503 : mux21_ni port map ( Y=>nx15502, A0=>nx15504, A1=>nx15508, S0=>
      nx17893);
   ix15505 : aoi21 port map ( Y=>nx15504, A0=>nflt_layer_out_1, A1=>
      nflt_layer_out_0, B0=>nx15506);
   ix15509 : inv01 port map ( Y=>nx15508, A=>mem_data_in(1));
   ix12942 : oai32 port map ( Y=>nx12941, A0=>nx15512, A1=>nx17893, A2=>
      nx17887, B0=>nx15514, B1=>nx18263);
   nflt_layer_out_2 : dffr port map ( Q=>OPEN, QB=>nx15512, D=>nx12941, CLK
      =>clk, R=>reset);
   ix15515 : mux21_ni port map ( Y=>nx15514, A0=>nx15516, A1=>nx15518, S0=>
      nx17895);
   ix15519 : inv01 port map ( Y=>nx15518, A=>mem_data_in(2));
   reg_nflt_layer_out_3 : dffr port map ( Q=>nflt_layer_out_3, QB=>OPEN, D=>
      nx12951, CLK=>clk, R=>reset);
   ix12952 : mux21_ni port map ( Y=>nx12951, A0=>nx78, A1=>nflt_layer_out_3, 
      S0=>nx18263);
   ix79 : mux21 port map ( Y=>nx78, A0=>nx15523, A1=>nx15527, S0=>nx17895);
   ix15524 : xnor2 port map ( Y=>nx15523, A0=>nflt_layer_out_3, A1=>nx15525
   );
   ix15528 : inv01 port map ( Y=>nx15527, A=>mem_data_in(3));
   reg_num_channels_counter_out_0 : dffr port map ( Q=>
      num_channels_counter_out_0, QB=>nx15531, D=>nx13911, CLK=>clk, R=>
      reset);
   ix1547 : oai21 port map ( Y=>nx1546, A0=>nx15422, A1=>nx15537, B0=>
      nx18269);
   ix15538 : nand02 port map ( Y=>nx15537, A0=>current_state_24, A1=>nx15637
   );
   ix1535 : oai21 port map ( Y=>nx1534, A0=>nx15541, A1=>nx17847, B0=>
      nx15716);
   ix1519 : nand02 port map ( Y=>nx1518, A0=>nx15544, A1=>nx16065);
   ix15545 : aoi32 port map ( Y=>nx15544, A0=>nx15546, A1=>
      comp_unit_finished, A2=>current_state_19, B0=>nx15561, B1=>nx12906);
   ix14032 : mux21_ni port map ( Y=>nx14031, A0=>layer_type_out_1, A1=>
      mem_data_in(1), S0=>current_state_3);
   layer_type_reg_q_1 : dffr port map ( Q=>layer_type_out_1, QB=>nx15548, D
      =>nx14031, CLK=>clk, R=>reset);
   ix1501 : oai221 port map ( Y=>nx1500, A0=>nx18273, A1=>nx17847, B0=>
      comp_unit_finished, B1=>nx15573, C0=>nx18059);
   reg_current_state_17 : dffr port map ( Q=>OPEN, QB=>nx15554, D=>nx1478, 
      CLK=>nx17835, R=>reset);
   ix13342 : mux21 port map ( Y=>nx13341, A0=>nx15559, A1=>nx15575, S0=>
      nx18045);
   ix15560 : aoi32 port map ( Y=>nx15559, A0=>nx15561, A1=>
      ftc_cntrl_reg_out_11, A2=>current_state_21, B0=>ftc_cntrl_reg_out_8, 
      B1=>nx158);
   ix13072 : mux21_ni port map ( Y=>nx13071, A0=>nx362, A1=>
      ftc_cntrl_reg_out_14, S0=>nx18045);
   ix363 : oai22 port map ( Y=>nx362, A0=>nx15561, A1=>nx15567, B0=>nx15563, 
      B1=>nx16198);
   ix15568 : aoi21 port map ( Y=>nx15567, A0=>nx17873, A1=>nx15621, B0=>
      current_state_21);
   ix1839 : oai321 port map ( Y=>nx1838, A0=>nx15546, A1=>nx15571, A2=>
      nx15573, B0=>nx15575, B1=>nx15602, C0=>nx16196);
   ix15572 : inv01 port map ( Y=>nx15571, A=>comp_unit_finished);
   reg_current_state_19 : dffr port map ( Q=>current_state_19, QB=>nx15573, 
      D=>nx1500, CLK=>nx17825, R=>reset);
   ftc_cntrl_reg_reg_q_8 : dffr port map ( Q=>ftc_cntrl_reg_out_8, QB=>
      nx15575, D=>nx13341, CLK=>nx17825, R=>nx17805);
   reg_current_state_13 : dffr port map ( Q=>current_state_13, QB=>OPEN, D=>
      nx330, CLK=>nx17825, R=>reset);
   ix331 : oai22 port map ( Y=>nx330, A0=>nx18255, A1=>nx316, B0=>nx15598, 
      B1=>nx196);
   ix317 : nand04 port map ( Y=>nx316, A0=>nx15580, A1=>
      cntr1_inst_counter_out_0, A2=>cntr1_inst_counter_out_3, A3=>nx15596);
   ix15581 : nor03_2x port map ( Y=>nx15580, A0=>nx310, A1=>nx278, A2=>nx276
   );
   cntr1_inst_counter_out_5 : dffr port map ( Q=>OPEN, QB=>nx15586, D=>
      nx13021, CLK=>clk, R=>nx17929);
   reg_cntr1_inst_counter_out_4 : dffr port map ( Q=>
      cntr1_inst_counter_out_4, QB=>nx15591, D=>nx13011, CLK=>clk, R=>
      nx17929);
   reg_cntr1_inst_counter_out_0 : dffr port map ( Q=>
      cntr1_inst_counter_out_0, QB=>OPEN, D=>nx12971, CLK=>clk, R=>nx17929);
   ix12972 : xnor2 port map ( Y=>nx12971, A0=>cntr1_inst_counter_out_0, A1=>
      nx18255);
   reg_current_state_10 : dffr port map ( Q=>current_state_10, QB=>nx15598, 
      D=>nx182, CLK=>nx17825, R=>reset);
   ix197 : nand02 port map ( Y=>nx196, A0=>nx18151, A1=>nx15548);
   reg_current_state_20 : dffr port map ( Q=>OPEN, QB=>nx15605, D=>nx1838, 
      CLK=>nx17825, R=>reset);
   ix13852 : mux21 port map ( Y=>nx13851, A0=>nx15609, A1=>nx15621, S0=>
      nx18045);
   ix15610 : nand04 port map ( Y=>nx15609, A0=>nx1402, A1=>nx1416, A2=>
      nx1434, A3=>nx1456);
   cache_width_cntr_counter_out_15 : dffr port map ( Q=>OPEN, QB=>nx15614, D
      =>nx13841, CLK=>clk, R=>nx17961);
   ix1225 : nand02 port map ( Y=>nx1224, A0=>nx15617, A1=>nx16065);
   ix15618 : aoi21 port map ( Y=>nx15617, A0=>nx15619, A1=>nx17921, B0=>
      nx17807);
   ftc_cntrl_reg_reg_q_12 : dffr port map ( Q=>ftc_cntrl_reg_out_12, QB=>
      nx15621, D=>nx13851, CLK=>nx17825, R=>nx17805);
   ix337 : or02 port map ( Y=>nx336, A0=>nx12883, A1=>nx17805);
   reg_current_state_14 : dffr port map ( Q=>OPEN, QB=>nx15626, D=>nx336, 
      CLK=>nx17827, R=>reset);
   ix13062 : mux21_ni port map ( Y=>nx13061, A0=>cache_height_ended, A1=>
      ftc_cntrl_reg_out_13, S0=>nx18045);
   reg_current_state_15 : dffr port map ( Q=>current_state_15, QB=>nx15861, 
      D=>nx1138, CLK=>nx17833, R=>reset);
   ix1139 : oai22 port map ( Y=>nx1138, A0=>nx15635, A1=>nx15637, B0=>
      nx18279, B1=>nx15859);
   reg_current_state_24 : dffr port map ( Q=>current_state_24, QB=>nx15635, 
      D=>nx1534, CLK=>nx17827, R=>reset);
   ix15638 : nor04 port map ( Y=>nx15637, A0=>nx1128, A1=>nx1040, A2=>nx944, 
      A3=>nx850);
   ix1129 : nand04 port map ( Y=>nx1128, A0=>nx15640, A1=>nx15781, A2=>
      nx15786, A3=>nx15791);
   ix13652 : oai22 port map ( Y=>nx13651, A0=>nx15644, A1=>nx18053, B0=>
      nx15776, B1=>nx17951);
   reg_write_offset_reg_q_14 : dffr port map ( Q=>write_offset_data_out_14, 
      QB=>nx15647, D=>nx13631, CLK=>nx17827, R=>reset);
   ix15654 : nand02 port map ( Y=>nx15653, A0=>write_offset_data_out_13, A1
      =>nx1042);
   ix13612 : oai22 port map ( Y=>nx13611, A0=>nx15657, A1=>nx18053, B0=>
      nx15774, B1=>nx17949);
   ix15658 : oai21 port map ( Y=>nx15657, A0=>nx1042, A1=>
      write_offset_data_out_13, B0=>nx15653);
   reg_write_offset_reg_q_12 : dffr port map ( Q=>write_offset_data_out_12, 
      QB=>nx15660, D=>nx13591, CLK=>nx17827, R=>reset);
   ix15667 : nand02 port map ( Y=>nx15666, A0=>write_offset_data_out_11, A1
      =>nx994);
   ix13572 : oai22 port map ( Y=>nx13571, A0=>nx15670, A1=>nx18051, B0=>
      nx15772, B1=>nx17949);
   ix15671 : oai21 port map ( Y=>nx15670, A0=>nx994, A1=>
      write_offset_data_out_11, B0=>nx15666);
   reg_write_offset_reg_q_10 : dffr port map ( Q=>write_offset_data_out_10, 
      QB=>nx15673, D=>nx13551, CLK=>nx17827, R=>reset);
   ix15680 : nand02 port map ( Y=>nx15679, A0=>write_offset_data_out_9, A1=>
      nx948);
   ix13532 : oai22 port map ( Y=>nx13531, A0=>nx15683, A1=>nx18051, B0=>
      nx15770, B1=>nx17949);
   ix15684 : oai21 port map ( Y=>nx15683, A0=>nx948, A1=>
      write_offset_data_out_9, B0=>nx15679);
   reg_write_offset_reg_q_8 : dffr port map ( Q=>write_offset_data_out_8, QB
      =>nx15686, D=>nx13511, CLK=>nx17827, R=>reset);
   ix15693 : nand02 port map ( Y=>nx15692, A0=>write_offset_data_out_7, A1=>
      nx898);
   ix13492 : oai22 port map ( Y=>nx13491, A0=>nx15696, A1=>nx17947, B0=>
      nx15717, B1=>nx18051);
   reg_write_offset_reg_q_7 : dffr port map ( Q=>write_offset_data_out_7, QB
      =>nx15696, D=>nx13491, CLK=>nx17827, R=>reset);
   reg_current_state_22 : dffr port map ( Q=>OPEN, QB=>nx15541, D=>nx1518, 
      CLK=>nx17829, R=>reset);
   reg_current_state_23 : dffr port map ( Q=>OPEN, QB=>nx15716, D=>nx1524, 
      CLK=>nx17829, R=>reset);
   ix13032 : mux21_ni port map ( Y=>nx13031, A0=>flt_size_out_0, A1=>
      mem_data_in(0), S0=>current_state_5);
   flt_size_reg_q_0 : dffr port map ( Q=>flt_size_out_0, QB=>OPEN, D=>
      nx13031, CLK=>clk, R=>reset);
   flt_size_reg_q_2 : dffr port map ( Q=>flt_size_out_2, QB=>nx15711, D=>
      nx13041, CLK=>clk, R=>reset);
   ix13042 : mux21_ni port map ( Y=>nx13041, A0=>flt_size_out_2, A1=>
      mem_data_in(2), S0=>current_state_5);
   ix13052 : mux21_ni port map ( Y=>nx13051, A0=>flt_size_out_1, A1=>
      mem_data_in(1), S0=>current_state_5);
   flt_size_reg_q_1 : dffr port map ( Q=>flt_size_out_1, QB=>OPEN, D=>
      nx13051, CLK=>clk, R=>reset);
   ix15718 : oai21 port map ( Y=>nx15717, A0=>nx898, A1=>
      write_offset_data_out_7, B0=>nx15692);
   reg_write_offset_reg_q_6 : dffr port map ( Q=>write_offset_data_out_6, QB
      =>nx15720, D=>nx13471, CLK=>nx17829, R=>reset);
   ix15727 : nand02 port map ( Y=>nx15726, A0=>write_offset_data_out_5, A1=>
      nx852);
   ix13452 : oai22 port map ( Y=>nx13451, A0=>nx15730, A1=>nx17947, B0=>
      nx15732, B1=>nx18049);
   reg_write_offset_reg_q_5 : dffr port map ( Q=>write_offset_data_out_5, QB
      =>nx15730, D=>nx13451, CLK=>nx17829, R=>reset);
   ix15733 : oai21 port map ( Y=>nx15732, A0=>nx852, A1=>
      write_offset_data_out_5, B0=>nx15726);
   reg_write_offset_reg_q_4 : dffr port map ( Q=>write_offset_data_out_4, QB
      =>nx15735, D=>nx13431, CLK=>nx17829, R=>reset);
   reg_write_offset_reg_q_3 : dffr port map ( Q=>write_offset_data_out_3, QB
      =>nx15745, D=>nx13411, CLK=>nx17829, R=>reset);
   ix13392 : oai22 port map ( Y=>nx13391, A0=>nx15750, A1=>nx17947, B0=>
      nx15753, B1=>nx18049);
   ix15754 : oai21 port map ( Y=>nx15753, A0=>nx780, A1=>
      write_offset_data_out_2, B0=>nx15768);
   ix13372 : oai22 port map ( Y=>nx13371, A0=>nx15756, A1=>nx17947, B0=>
      nx15759, B1=>nx18049);
   ix15760 : oai21 port map ( Y=>nx15759, A0=>write_offset_data_out_0, A1=>
      write_offset_data_out_1, B0=>nx15765);
   reg_write_offset_reg_q_0 : dffr port map ( Q=>write_offset_data_out_0, QB
      =>nx15763, D=>nx13351, CLK=>nx17829, R=>reset);
   reg_write_offset_reg_q_1 : dffr port map ( Q=>write_offset_data_out_1, QB
      =>nx15756, D=>nx13371, CLK=>nx17831, R=>reset);
   reg_write_offset_reg_q_2 : dffr port map ( Q=>write_offset_data_out_2, QB
      =>nx15750, D=>nx13391, CLK=>nx17831, R=>reset);
   reg_write_offset_reg_q_9 : dffr port map ( Q=>write_offset_data_out_9, QB
      =>nx15770, D=>nx13531, CLK=>nx17831, R=>reset);
   reg_write_offset_reg_q_11 : dffr port map ( Q=>write_offset_data_out_11, 
      QB=>nx15772, D=>nx13571, CLK=>nx17831, R=>reset);
   reg_write_offset_reg_q_13 : dffr port map ( Q=>write_offset_data_out_13, 
      QB=>nx15774, D=>nx13611, CLK=>nx17831, R=>reset);
   reg_write_offset_reg_q_15 : dffr port map ( Q=>write_offset_data_out_15, 
      QB=>nx15776, D=>nx13651, CLK=>nx17831, R=>reset);
   new_size_squared_reg_q_15 : dffr port map ( Q=>new_size_squared_out_15, 
      QB=>OPEN, D=>nx13661, CLK=>clk, R=>reset);
   new_size_squared_reg_q_14 : dffr port map ( Q=>new_size_squared_out_14, 
      QB=>nx15785, D=>nx13641, CLK=>clk, R=>reset);
   new_size_squared_reg_q_13 : dffr port map ( Q=>new_size_squared_out_13, 
      QB=>OPEN, D=>nx13621, CLK=>clk, R=>reset);
   new_size_squared_reg_q_12 : dffr port map ( Q=>new_size_squared_out_12, 
      QB=>nx15795, D=>nx13601, CLK=>clk, R=>reset);
   ix1041 : nand04 port map ( Y=>nx1040, A0=>nx15797, A1=>nx15802, A2=>
      nx15807, A3=>nx15812);
   new_size_squared_reg_q_11 : dffr port map ( Q=>new_size_squared_out_11, 
      QB=>OPEN, D=>nx13581, CLK=>clk, R=>reset);
   new_size_squared_reg_q_10 : dffr port map ( Q=>new_size_squared_out_10, 
      QB=>nx15806, D=>nx13561, CLK=>clk, R=>reset);
   new_size_squared_reg_q_9 : dffr port map ( Q=>new_size_squared_out_9, QB
      =>OPEN, D=>nx13541, CLK=>clk, R=>reset);
   new_size_squared_reg_q_8 : dffr port map ( Q=>new_size_squared_out_8, QB
      =>nx15816, D=>nx13521, CLK=>clk, R=>reset);
   ix945 : nand04 port map ( Y=>nx944, A0=>nx15818, A1=>nx15823, A2=>nx15828, 
      A3=>nx15833);
   new_size_squared_reg_q_7 : dffr port map ( Q=>new_size_squared_out_7, QB
      =>OPEN, D=>nx13501, CLK=>clk, R=>reset);
   new_size_squared_reg_q_6 : dffr port map ( Q=>new_size_squared_out_6, QB
      =>nx15827, D=>nx13481, CLK=>clk, R=>reset);
   new_size_squared_reg_q_5 : dffr port map ( Q=>new_size_squared_out_5, QB
      =>OPEN, D=>nx13461, CLK=>clk, R=>reset);
   new_size_squared_reg_q_4 : dffr port map ( Q=>new_size_squared_out_4, QB
      =>nx15837, D=>nx13441, CLK=>clk, R=>reset);
   ix851 : nand04 port map ( Y=>nx850, A0=>nx15839, A1=>nx15844, A2=>nx15849, 
      A3=>nx15854);
   new_size_squared_reg_q_3 : dffr port map ( Q=>new_size_squared_out_3, QB
      =>OPEN, D=>nx13421, CLK=>clk, R=>reset);
   new_size_squared_reg_q_2 : dffr port map ( Q=>new_size_squared_out_2, QB
      =>nx15848, D=>nx13401, CLK=>clk, R=>reset);
   new_size_squared_reg_q_1 : dffr port map ( Q=>new_size_squared_out_1, QB
      =>OPEN, D=>nx13381, CLK=>clk, R=>reset);
   new_size_squared_reg_q_0 : dffr port map ( Q=>new_size_squared_out_0, QB
      =>OPEN, D=>nx13361, CLK=>clk, R=>reset);
   ftc_cntrl_reg_reg_q_13 : dffr port map ( Q=>ftc_cntrl_reg_out_13, QB=>
      nx15859, D=>nx13061, CLK=>nx17831, R=>nx17805);
   ix1169 : nand02 port map ( Y=>nx1168, A0=>nx18225, A1=>nx15878);
   ix13332 : mux21 port map ( Y=>nx13331, A0=>nx15868, A1=>nx15865, S0=>
      nx18045);
   ix15869 : nand04 port map ( Y=>nx15868, A0=>nx550, A1=>nx564, A2=>nx612, 
      A3=>nx732);
   window_width_cntr_counter_out_15 : dffr port map ( Q=>OPEN, QB=>nx15873, 
      D=>nx13221, CLK=>clk, R=>nx17939);
   ix379 : nand02 port map ( Y=>nx378, A0=>nx15876, A1=>nx15878);
   ix15877 : aoi22 port map ( Y=>nx15876, A0=>nx17921, A1=>
      ftc_cntrl_reg_out_13, B0=>nx17871, B1=>ftc_cntrl_reg_out_12);
   ix13672 : mux21_ni port map ( Y=>nx13671, A0=>nx1154, A1=>
      ftc_cntrl_reg_out_9, S0=>nx18045);
   ix1155 : oai21 port map ( Y=>nx1154, A0=>nx15883, A1=>nx15885, B0=>
      nx15876);
   ftc_cntrl_reg_reg_q_9 : dffr port map ( Q=>ftc_cntrl_reg_out_9, QB=>
      nx15883, D=>nx13671, CLK=>nx17833, R=>nx17805);
   ix15886 : aoi21 port map ( Y=>nx15885, A0=>nx18225, A1=>nx1146, B0=>
      nx17921);
   reg_current_state_16 : dffr port map ( Q=>current_state_16, QB=>nx15888, 
      D=>nx1168, CLK=>nx17833, R=>reset);
   reg_window_width_cntr_counter_out_14 : dffr port map ( Q=>
      window_width_cntr_counter_out_14, QB=>nx15893, D=>nx13211, CLK=>clk, R
      =>nx17939);
   ix15899 : nand02 port map ( Y=>nx15898, A0=>
      window_width_cntr_counter_out_13, A1=>nx12887);
   reg_window_width_cntr_counter_out_13 : dffr port map ( Q=>
      window_width_cntr_counter_out_13, QB=>nx15902, D=>nx13201, CLK=>clk, R
      =>nx17939);
   ix15905 : oai21 port map ( Y=>nx15904, A0=>nx12887, A1=>
      window_width_cntr_counter_out_13, B0=>nx15898);
   reg_window_width_cntr_counter_out_12 : dffr port map ( Q=>
      window_width_cntr_counter_out_12, QB=>nx15907, D=>nx13191, CLK=>clk, R
      =>nx17939);
   ix15913 : nand02 port map ( Y=>nx15912, A0=>
      window_width_cntr_counter_out_11, A1=>nx12889);
   reg_window_width_cntr_counter_out_11 : dffr port map ( Q=>
      window_width_cntr_counter_out_11, QB=>nx15916, D=>nx13181, CLK=>clk, R
      =>nx17939);
   ix15919 : oai21 port map ( Y=>nx15918, A0=>nx12889, A1=>
      window_width_cntr_counter_out_11, B0=>nx15912);
   reg_window_width_cntr_counter_out_10 : dffr port map ( Q=>
      window_width_cntr_counter_out_10, QB=>nx15921, D=>nx13171, CLK=>clk, R
      =>nx17939);
   ix15927 : nand02 port map ( Y=>nx15926, A0=>
      window_width_cntr_counter_out_9, A1=>nx12891);
   reg_window_width_cntr_counter_out_9 : dffr port map ( Q=>
      window_width_cntr_counter_out_9, QB=>nx15930, D=>nx13161, CLK=>clk, R
      =>nx17939);
   ix15933 : oai21 port map ( Y=>nx15932, A0=>nx12891, A1=>
      window_width_cntr_counter_out_9, B0=>nx15926);
   reg_window_width_cntr_counter_out_8 : dffr port map ( Q=>
      window_width_cntr_counter_out_8, QB=>nx15935, D=>nx13151, CLK=>clk, R
      =>nx17941);
   ix15941 : nand02 port map ( Y=>nx15940, A0=>
      window_width_cntr_counter_out_7, A1=>nx12893);
   reg_window_width_cntr_counter_out_7 : dffr port map ( Q=>
      window_width_cntr_counter_out_7, QB=>nx15944, D=>nx13141, CLK=>clk, R
      =>nx17941);
   ix15947 : oai21 port map ( Y=>nx15946, A0=>nx12893, A1=>
      window_width_cntr_counter_out_7, B0=>nx15940);
   reg_window_width_cntr_counter_out_6 : dffr port map ( Q=>
      window_width_cntr_counter_out_6, QB=>nx15949, D=>nx13131, CLK=>clk, R
      =>nx17941);
   reg_wind_width_count_4 : dffr port map ( Q=>wind_width_count_4, QB=>OPEN, 
      D=>nx14041, CLK=>clk, R=>nx17943);
   ix1877 : xnor2 port map ( Y=>nx1876, A0=>wind_width_count_4, A1=>nx15959
   );
   ix15960 : nand04 port map ( Y=>nx15959, A0=>wind_width_count_1, A1=>
      nx17811, A2=>wind_width_count_2, A3=>wind_width_count_3);
   reg_wind_width_count_1 : dffr port map ( Q=>wind_width_count_1, QB=>OPEN, 
      D=>nx13091, CLK=>clk, R=>nx17941);
   ix385 : xor2 port map ( Y=>nx384, A0=>wind_width_count_1, A1=>nx17811);
   reg_wind_width_count_0 : dffr port map ( Q=>wind_width_count_0, QB=>OPEN, 
      D=>nx13081, CLK=>clk, R=>nx17941);
   reg_current_state_21 : dffr port map ( Q=>current_state_21, QB=>nx15970, 
      D=>nx12877, CLK=>nx17833, R=>reset);
   ftc_cntrl_reg_reg_q_11 : dffr port map ( Q=>ftc_cntrl_reg_out_11, QB=>
      nx15865, D=>nx13331, CLK=>nx17833, R=>nx17805);
   ix1875 : oai22 port map ( Y=>nx12884, A0=>ftc_cntrl_reg_out_9, A1=>
      nx18225, B0=>nx15970, B1=>ftc_cntrl_reg_out_11);
   reg_wind_width_count_2 : dffr port map ( Q=>wind_width_count_2, QB=>OPEN, 
      D=>nx13101, CLK=>clk, R=>nx17941);
   ix393 : xnor2 port map ( Y=>nx392, A0=>wind_width_count_2, A1=>nx15983);
   ix15984 : nand02 port map ( Y=>nx15983, A0=>wind_width_count_1, A1=>
      nx17813);
   reg_wind_width_count_3 : dffr port map ( Q=>wind_width_count_3, QB=>OPEN, 
      D=>nx13111, CLK=>clk, R=>nx17941);
   ix401 : xnor2 port map ( Y=>nx400, A0=>wind_width_count_3, A1=>nx15989);
   ix15990 : nand03 port map ( Y=>nx15989, A0=>wind_width_count_1, A1=>
      nx17813, A2=>wind_width_count_2);
   reg_window_width_cntr_counter_out_5 : dffr port map ( Q=>
      window_width_cntr_counter_out_5, QB=>nx15995, D=>nx13121, CLK=>clk, R
      =>nx17943);
   ix15998 : oai21 port map ( Y=>nx15997, A0=>nx408, A1=>
      window_width_cntr_counter_out_5, B0=>nx15954);
   ix409 : nor02ii port map ( Y=>nx408, A0=>nx15959, A1=>wind_width_count_4
   );
   ix605 : xor2 port map ( Y=>nx604, A0=>nx602, A1=>nx17813);
   img_width_reg_q_0 : dffr port map ( Q=>img_width_out_0, QB=>nx16005, D=>
      nx13241, CLK=>clk, R=>reset);
   ix13232 : mux21_ni port map ( Y=>nx13231, A0=>new_width_out_0, A1=>
      mem_data_in(0), S0=>current_state_6);
   new_width_reg_q_0 : dffr port map ( Q=>new_width_out_0, QB=>OPEN, D=>
      nx13231, CLK=>clk, R=>reset);
   ix733 : and04 port map ( Y=>nx732, A0=>nx16013, A1=>nx16025, A2=>nx16039, 
      A3=>nx16052);
   ix16014 : xnor2 port map ( Y=>nx16013, A0=>wind_width_count_1, A1=>nx640
   );
   img_width_reg_q_1 : dffr port map ( Q=>img_width_out_1, QB=>nx16019, D=>
      nx13261, CLK=>clk, R=>reset);
   ix13252 : mux21_ni port map ( Y=>nx13251, A0=>new_width_out_1, A1=>
      mem_data_in(1), S0=>current_state_6);
   new_width_reg_q_1 : dffr port map ( Q=>new_width_out_1, QB=>OPEN, D=>
      nx13251, CLK=>clk, R=>reset);
   ix16026 : xnor2 port map ( Y=>nx16025, A0=>wind_width_count_2, A1=>nx674
   );
   ix675 : mux21 port map ( Y=>nx674, A0=>nx17845, A1=>nx18055, S0=>nx18225
   );
   ix16029 : aoi21 port map ( Y=>nx16028, A0=>img_width_out_2, A1=>nx630, B0
      =>nx16037);
   img_width_reg_q_2 : dffs_ni port map ( Q=>img_width_out_2, QB=>OPEN, D=>
      nx13281, CLK=>clk, S=>reset);
   ix13282 : ao221 port map ( Y=>nx13281, A0=>nx17875, A1=>new_width_out_2, 
      B0=>img_width_out_2, B1=>nx18259, C0=>nx17897);
   new_width_reg_q_2 : dffr port map ( Q=>new_width_out_2, QB=>OPEN, D=>
      nx13271, CLK=>clk, R=>reset);
   ix13272 : mux21_ni port map ( Y=>nx13271, A0=>new_width_out_2, A1=>
      mem_data_in(2), S0=>current_state_6);
   ix16038 : nor03_2x port map ( Y=>nx16037, A0=>img_width_out_0, A1=>
      img_width_out_1, A2=>img_width_out_2);
   ix16040 : xnor2 port map ( Y=>nx16039, A0=>wind_width_count_3, A1=>nx704
   );
   img_width_reg_q_3 : dffs_ni port map ( Q=>img_width_out_3, QB=>nx16046, D
      =>nx13301, CLK=>clk, S=>reset);
   ix13292 : mux21_ni port map ( Y=>nx13291, A0=>new_width_out_3, A1=>
      mem_data_in(3), S0=>current_state_6);
   new_width_reg_q_3 : dffr port map ( Q=>new_width_out_3, QB=>OPEN, D=>
      nx13291, CLK=>clk, R=>reset);
   ix16053 : xnor2 port map ( Y=>nx16052, A0=>wind_width_count_4, A1=>nx722
   );
   ix16056 : xnor2 port map ( Y=>nx16055, A0=>img_width_out_4, A1=>nx16063);
   img_width_reg_q_4 : dffs_ni port map ( Q=>img_width_out_4, QB=>OPEN, D=>
      nx13321, CLK=>clk, S=>reset);
   ix13322 : ao22 port map ( Y=>nx13321, A0=>nx17875, A1=>new_width_out_4, 
      B0=>img_width_out_4, B1=>nx18259);
   new_width_reg_q_4 : dffr port map ( Q=>new_width_out_4, QB=>OPEN, D=>
      nx13311, CLK=>clk, R=>reset);
   ix13312 : mux21_ni port map ( Y=>nx13311, A0=>new_width_out_4, A1=>
      mem_data_in(4), S0=>current_state_6);
   reg_cache_width_cntr_counter_out_14 : dffr port map ( Q=>
      cache_width_cntr_counter_out_14, QB=>nx16070, D=>nx13831, CLK=>clk, R
      =>nx17961);
   ix16076 : nand02 port map ( Y=>nx16075, A0=>
      cache_width_cntr_counter_out_13, A1=>nx12898);
   reg_cache_width_cntr_counter_out_13 : dffr port map ( Q=>
      cache_width_cntr_counter_out_13, QB=>nx16079, D=>nx13821, CLK=>clk, R
      =>nx17961);
   ix16082 : oai21 port map ( Y=>nx16081, A0=>nx12898, A1=>
      cache_width_cntr_counter_out_13, B0=>nx16075);
   reg_cache_width_cntr_counter_out_12 : dffr port map ( Q=>
      cache_width_cntr_counter_out_12, QB=>nx16084, D=>nx13811, CLK=>clk, R
      =>nx17961);
   ix16090 : nand02 port map ( Y=>nx16089, A0=>
      cache_width_cntr_counter_out_11, A1=>nx12900);
   reg_cache_width_cntr_counter_out_11 : dffr port map ( Q=>
      cache_width_cntr_counter_out_11, QB=>nx16093, D=>nx13801, CLK=>clk, R
      =>nx17961);
   ix16096 : oai21 port map ( Y=>nx16095, A0=>nx12900, A1=>
      cache_width_cntr_counter_out_11, B0=>nx16089);
   reg_cache_width_cntr_counter_out_10 : dffr port map ( Q=>
      cache_width_cntr_counter_out_10, QB=>nx16098, D=>nx13791, CLK=>clk, R
      =>nx17961);
   ix16104 : nand02 port map ( Y=>nx16103, A0=>
      cache_width_cntr_counter_out_9, A1=>nx12902);
   reg_cache_width_cntr_counter_out_9 : dffr port map ( Q=>
      cache_width_cntr_counter_out_9, QB=>nx16107, D=>nx13781, CLK=>clk, R=>
      nx17961);
   ix16110 : oai21 port map ( Y=>nx16109, A0=>nx12902, A1=>
      cache_width_cntr_counter_out_9, B0=>nx16103);
   reg_cache_width_cntr_counter_out_8 : dffr port map ( Q=>
      cache_width_cntr_counter_out_8, QB=>nx16112, D=>nx13771, CLK=>clk, R=>
      nx17963);
   ix16118 : nand02 port map ( Y=>nx16117, A0=>
      cache_width_cntr_counter_out_7, A1=>nx12904);
   reg_cache_width_cntr_counter_out_7 : dffr port map ( Q=>
      cache_width_cntr_counter_out_7, QB=>nx16121, D=>nx13761, CLK=>clk, R=>
      nx17963);
   ix16124 : oai21 port map ( Y=>nx16123, A0=>nx12904, A1=>
      cache_width_cntr_counter_out_7, B0=>nx16117);
   reg_cache_width_cntr_counter_out_6 : dffr port map ( Q=>
      cache_width_cntr_counter_out_6, QB=>nx16126, D=>nx13751, CLK=>clk, R=>
      nx17963);
   reg_cache_width_count_4 : dffr port map ( Q=>cache_width_count_4, QB=>
      OPEN, D=>nx13731, CLK=>clk, R=>nx17965);
   ix1255 : xnor2 port map ( Y=>nx1254, A0=>nx17815, A1=>nx16136);
   ix16137 : nand04 port map ( Y=>nx16136, A0=>cache_width_count_1, A1=>
      cache_width_count_0, A2=>nx17819, A3=>cache_width_count_3);
   reg_cache_width_count_1 : dffr port map ( Q=>cache_width_count_1, QB=>
      OPEN, D=>nx13701, CLK=>clk, R=>nx17963);
   ix1231 : xor2 port map ( Y=>nx1230, A0=>cache_width_count_1, A1=>
      cache_width_count_0);
   reg_cache_width_count_0 : dffr port map ( Q=>cache_width_count_0, QB=>
      OPEN, D=>nx13691, CLK=>clk, R=>nx17963);
   ix13682 : mux21_ni port map ( Y=>nx13681, A0=>nx1206, A1=>
      ftc_cntrl_reg_out_10, S0=>nx18045);
   ix1207 : oai21 port map ( Y=>nx1206, A0=>nx16148, A1=>nx16150, B0=>
      nx16155);
   ftc_cntrl_reg_reg_q_10 : dffr port map ( Q=>ftc_cntrl_reg_out_10, QB=>
      nx16148, D=>nx13681, CLK=>nx17833, R=>nx17807);
   ix1195 : nor03_2x port map ( Y=>cache_height_count_en, A0=>nx16153, A1=>
      ftc_cntrl_reg_out_13, A2=>nx15621);
   ix16156 : oai21 port map ( Y=>nx16155, A0=>nx17871, A1=>nx12883, B0=>
      nx15621);
   reg_cache_width_count_2 : dffr port map ( Q=>cache_width_count_2, QB=>
      OPEN, D=>nx13711, CLK=>clk, R=>nx17963);
   ix1239 : xnor2 port map ( Y=>nx1238, A0=>nx17819, A1=>nx16166);
   ix16167 : nand02 port map ( Y=>nx16166, A0=>cache_width_count_1, A1=>
      cache_width_count_0);
   reg_cache_width_count_3 : dffr port map ( Q=>cache_width_count_3, QB=>
      OPEN, D=>nx13721, CLK=>clk, R=>nx17963);
   ix1247 : xnor2 port map ( Y=>nx1246, A0=>cache_width_count_3, A1=>nx16172
   );
   ix16173 : nand03 port map ( Y=>nx16172, A0=>cache_width_count_1, A1=>
      cache_width_count_0, A2=>nx17821);
   reg_cache_width_cntr_counter_out_5 : dffr port map ( Q=>
      cache_width_cntr_counter_out_5, QB=>nx16178, D=>nx13741, CLK=>clk, R=>
      nx17965);
   ix16181 : oai21 port map ( Y=>nx16180, A0=>nx1260, A1=>
      cache_width_cntr_counter_out_5, B0=>nx16131);
   ix1261 : nor02ii port map ( Y=>nx1260, A0=>nx16136, A1=>nx17817);
   ix1457 : nor04 port map ( Y=>nx1456, A0=>nx1436, A1=>nx1438, A2=>nx1446, 
      A3=>nx1448);
   ix16190 : aoi21 port map ( Y=>nx16189, A0=>img_width_out_1, A1=>
      img_width_out_0, B0=>nx16191);
   ix1439 : xnor2 port map ( Y=>nx1438, A0=>nx17821, A1=>nx18055);
   ix1447 : xnor2 port map ( Y=>nx1446, A0=>cache_width_count_3, A1=>nx16042
   );
   ix1449 : xnor2 port map ( Y=>nx1448, A0=>nx17817, A1=>nx16055);
   ix16197 : aoi43 port map ( Y=>nx16196, A0=>nx15563, A1=>nx17845, A2=>
      nx17871, A3=>nx15621, B0=>nx15561, B1=>ftc_cntrl_reg_out_11, B2=>
      current_state_21);
   ix16199 : aoi22 port map ( Y=>nx16198, A0=>nx17921, A1=>nx15859, B0=>
      nx15970, B1=>nx16153);
   ftc_cntrl_reg_reg_q_14 : dffr port map ( Q=>ftc_cntrl_reg_out_14, QB=>
      nx15563, D=>nx13071, CLK=>nx17833, R=>nx17807);
   ix159 : nand02 port map ( Y=>nx158, A0=>nx16202, A1=>nx16204);
   ix16203 : oai21 port map ( Y=>nx16202, A0=>nx17873, A1=>nx15970, B0=>
      nx16065);
   ix16205 : aoi43 port map ( Y=>nx16204, A0=>nx17873, A1=>nx15621, A2=>
      nx15575, A3=>nx15561, B0=>current_state_21, B1=>nx15563, B2=>nx17845);
   reg_current_state_18 : dffr port map ( Q=>current_state_18, QB=>OPEN, D=>
      nx1484, CLK=>nx17835, R=>reset);
   reg_num_channels_counter_out_1 : dffr port map ( Q=>
      num_channels_counter_out_1, QB=>OPEN, D=>nx13931, CLK=>clk, R=>reset);
   ix13932 : mux21_ni port map ( Y=>nx13931, A0=>num_channels_counter_out_1, 
      A1=>nx1648, S0=>nx17973);
   ix1649 : oai321 port map ( Y=>nx1648, A0=>nx16213, A1=>nx18265, A2=>
      nx18151, B0=>nx148, B1=>nx16224, C0=>nx16228);
   max_num_channels_inst_reg_q_1 : dffr port map ( Q=>OPEN, QB=>nx16213, D=>
      nx13921, CLK=>clk, R=>reset);
   ix13922 : oai32 port map ( Y=>nx13921, A0=>nx16213, A1=>nx17897, A2=>
      nx17875, B0=>nx16216, B1=>nx18259);
   ix16217 : aoi22 port map ( Y=>nx16216, A0=>mem_data_in(1), A1=>nx17897, 
      B0=>nx17875, B1=>nflt_layer_temp_1);
   nflt_layer_total_reg_q_1 : dffr port map ( Q=>nflt_layer_temp_1, QB=>OPEN, 
      D=>nx13881, CLK=>clk, R=>reset);
   ix13882 : mux21_ni port map ( Y=>nx13881, A0=>nflt_layer_temp_1, A1=>
      mem_data_in(1), S0=>nx17895);
   ix16225 : aoi21 port map ( Y=>nx16224, A0=>num_channels_counter_out_1, A1
      =>num_channels_counter_out_0, B0=>nx16226);
   ix16229 : aoi22 port map ( Y=>nx16228, A0=>mem_data_in(1), A1=>nx17899, 
      B0=>nx17877, B1=>nflt_layer_temp_1);
   ix13952 : mux21_ni port map ( Y=>nx13951, A0=>num_channels_counter_out_2, 
      A1=>nx1674, S0=>nx17973);
   ix1675 : oai21 port map ( Y=>nx1674, A0=>nx16234, A1=>nx18269, B0=>
      nx16239);
   ix16235 : aoi22 port map ( Y=>nx16234, A0=>mem_data_in(2), A1=>nx17899, 
      B0=>nx17877, B1=>nflt_layer_temp_2);
   nflt_layer_total_reg_q_2 : dffr port map ( Q=>nflt_layer_temp_2, QB=>OPEN, 
      D=>nx13871, CLK=>clk, R=>reset);
   ix13872 : mux21_ni port map ( Y=>nx13871, A0=>nflt_layer_temp_2, A1=>
      mem_data_in(2), S0=>nx17895);
   ix16240 : aoi22 port map ( Y=>nx16239, A0=>max_num_channels_data_out_2, 
      A1=>nx1642, B0=>nx18269, B1=>nx1660);
   ix13942 : oai32 port map ( Y=>nx13941, A0=>nx16243, A1=>nx17899, A2=>
      nx17877, B0=>nx16234, B1=>nx18259);
   max_num_channels_inst_reg_q_2 : dffr port map ( Q=>
      max_num_channels_data_out_2, QB=>nx16243, D=>nx13941, CLK=>clk, R=>
      reset);
   ix1643 : nor02_2x port map ( Y=>nx1642, A0=>nx18265, A1=>nx18151);
   ix1661 : oai21 port map ( Y=>nx1660, A0=>nx16247, A1=>nx16226, B0=>
      nx12908);
   reg_num_channels_counter_out_2 : dffr port map ( Q=>
      num_channels_counter_out_2, QB=>nx16247, D=>nx13951, CLK=>clk, R=>
      reset);
   reg_num_channels_counter_out_3 : dffr port map ( Q=>
      num_channels_counter_out_3, QB=>OPEN, D=>nx13971, CLK=>clk, R=>reset);
   ix13972 : mux21_ni port map ( Y=>nx13971, A0=>num_channels_counter_out_3, 
      A1=>nx1700, S0=>nx17973);
   ix1701 : oai21 port map ( Y=>nx1700, A0=>nx16253, A1=>nx18269, B0=>
      nx16258);
   ix16254 : aoi22 port map ( Y=>nx16253, A0=>mem_data_in(3), A1=>nx17899, 
      B0=>nx17877, B1=>nflt_layer_temp_3);
   nflt_layer_total_reg_q_3 : dffr port map ( Q=>nflt_layer_temp_3, QB=>OPEN, 
      D=>nx13861, CLK=>clk, R=>reset);
   ix13862 : mux21_ni port map ( Y=>nx13861, A0=>nflt_layer_temp_3, A1=>
      mem_data_in(3), S0=>nx17895);
   ix16259 : aoi22 port map ( Y=>nx16258, A0=>max_num_channels_data_out_3, 
      A1=>nx1642, B0=>nx18269, B1=>nx1686);
   ix13962 : oai32 port map ( Y=>nx13961, A0=>nx16262, A1=>nx17899, A2=>
      nx17877, B0=>nx16253, B1=>nx18259);
   max_num_channels_inst_reg_q_3 : dffr port map ( Q=>
      max_num_channels_data_out_3, QB=>nx16262, D=>nx13961, CLK=>clk, R=>
      reset);
   ix1687 : xor2 port map ( Y=>nx1686, A0=>num_channels_counter_out_3, A1=>
      nx16265);
   ix16266 : nor03_2x port map ( Y=>nx16265, A0=>num_channels_counter_out_0, 
      A1=>num_channels_counter_out_1, A2=>num_channels_counter_out_2);
   ix16270 : nor03_2x port map ( Y=>nx16269, A0=>nlayers_counter_out_1, A1=>
      nlayers_counter_out_2, A2=>nx16278);
   reg_nlayers_counter_out_1 : dffr port map ( Q=>nlayers_counter_out_1, QB
      =>OPEN, D=>nx14011, CLK=>clk, R=>reset);
   ix14012 : mux21_ni port map ( Y=>nx14011, A0=>nx1764, A1=>
      nlayers_counter_out_1, S0=>nx16282);
   ix16275 : aoi21 port map ( Y=>nx16274, A0=>nlayers_counter_out_1, A1=>
      nlayers_counter_out_0, B0=>nx16284);
   ix14002 : oai32 port map ( Y=>nx14001, A0=>nx16278, A1=>current_state_2, 
      A2=>nx17877, B0=>nx16280, B1=>nx16282);
   reg_nlayers_counter_out_0 : dffr port map ( Q=>nlayers_counter_out_0, QB
      =>nx16278, D=>nx14001, CLK=>clk, R=>reset);
   reg_nlayers_counter_out_2 : dffr port map ( Q=>nlayers_counter_out_2, QB
      =>OPEN, D=>nx14021, CLK=>clk, R=>reset);
   ix14022 : mux21_ni port map ( Y=>nx14021, A0=>nx1780, A1=>
      nlayers_counter_out_2, S0=>nx16282);
   ix16291 : xnor2 port map ( Y=>nx16290, A0=>nlayers_counter_out_2, A1=>
      nx16284);
   ix16300 : inv01 port map ( Y=>nx16299, A=>mem_data_in(4));
   ix1713 : oai21 port map ( Y=>nx1712, A0=>nx15426, A1=>nx15460, B0=>
      nx12875);
   reg_current_state_12 : dffr port map ( Q=>OPEN, QB=>nx16302, D=>nx174, 
      CLK=>nx17837, R=>reset);
   ix175 : nand03 port map ( Y=>nx174, A0=>nx16305, A1=>nx15435, A2=>nx18265
   );
   ix16306 : oai21 port map ( Y=>nx16305, A0=>nx18151, A1=>nx15548, B0=>
      current_state_8);
   ix16308 : oai21 port map ( Y=>nx16307, A0=>cntr1_inst_counter_out_0, A1=>
      cntr1_inst_counter_out_1, B0=>nx15412);
   ix16314 : nand02 port map ( Y=>nx16313, A0=>current_state_10, A1=>nx196);
   ix1939 : nand02 port map ( Y=>nx1938, A0=>nx16318, A1=>nx18075);
   ix16319 : nand03 port map ( Y=>nx16318, A0=>nx12873, A1=>nx15486, A2=>
      nx16269);
   ix1737 : nor02_2x port map ( Y=>nx12873, A0=>nx12875, A1=>nx15537);
   reg_current_state_27 : dffr port map ( Q=>current_state_27, QB=>nx16327, 
      D=>nx1938, CLK=>nx17837, R=>reset);
   reg_class_cntr_counter_out_0 : dffr port map ( Q=>
      class_cntr_counter_out_0, QB=>nx16324, D=>nx14051, CLK=>nx17837, R=>
      reset);
   reg_class_cntr_counter_out_1 : dffr port map ( Q=>
      class_cntr_counter_out_1, QB=>nx16332, D=>nx14061, CLK=>nx17837, R=>
      reset);
   ix16335 : oai21 port map ( Y=>nx16334, A0=>class_cntr_counter_out_0, A1=>
      class_cntr_counter_out_1, B0=>nx16336);
   reg_class_cntr_counter_out_2 : dffr port map ( Q=>
      class_cntr_counter_out_2, QB=>nx16338, D=>nx14071, CLK=>nx17837, R=>
      reset);
   reg_class_cntr_counter_out_3 : dffr port map ( Q=>
      class_cntr_counter_out_3, QB=>nx16348, D=>nx14081, CLK=>nx17837, R=>
      reset);
   reg_flt_bias1_reg_q_0 : dff port map ( Q=>flt_bias_out_0, QB=>OPEN, D=>
      nx14101, CLK=>clk);
   ix14102 : mux21_ni port map ( Y=>nx14101, A0=>flt_bias_out_0, A1=>
      mem_data_in(0), S0=>nx17993);
   ix2129 : nor02_2x port map ( Y=>nx2128, A0=>nx16302, A1=>nx18153);
   ix14092 : oai21 port map ( Y=>nx14091, A0=>nx18297, A1=>nx182, B0=>
      nx16302);
   channel_zero_reg_q_0 : dffr port map ( Q=>OPEN, QB=>nx16373, D=>nx14091, 
      CLK=>clk, R=>reset);
   reg_flt_bias1_reg_q_1 : dff port map ( Q=>flt_bias_out_1, QB=>OPEN, D=>
      nx14121, CLK=>clk);
   ix14122 : mux21_ni port map ( Y=>nx14121, A0=>flt_bias_out_1, A1=>
      mem_data_in(1), S0=>nx17993);
   reg_flt_bias1_reg_q_2 : dff port map ( Q=>flt_bias_out_2, QB=>OPEN, D=>
      nx14141, CLK=>clk);
   ix14142 : mux21_ni port map ( Y=>nx14141, A0=>flt_bias_out_2, A1=>
      mem_data_in(2), S0=>nx17993);
   reg_flt_bias1_reg_q_3 : dff port map ( Q=>flt_bias_out_3, QB=>OPEN, D=>
      nx14161, CLK=>clk);
   ix14162 : mux21_ni port map ( Y=>nx14161, A0=>flt_bias_out_3, A1=>
      mem_data_in(3), S0=>nx17993);
   reg_flt_bias1_reg_q_4 : dff port map ( Q=>flt_bias_out_4, QB=>OPEN, D=>
      nx14181, CLK=>clk);
   ix14182 : mux21_ni port map ( Y=>nx14181, A0=>flt_bias_out_4, A1=>
      mem_data_in(4), S0=>nx17993);
   reg_flt_bias1_reg_q_5 : dff port map ( Q=>flt_bias_out_5, QB=>OPEN, D=>
      nx14201, CLK=>clk);
   ix14202 : mux21_ni port map ( Y=>nx14201, A0=>flt_bias_out_5, A1=>
      mem_data_in(5), S0=>nx17993);
   reg_flt_bias1_reg_q_6 : dff port map ( Q=>flt_bias_out_6, QB=>OPEN, D=>
      nx14221, CLK=>clk);
   ix14222 : mux21_ni port map ( Y=>nx14221, A0=>flt_bias_out_6, A1=>
      mem_data_in(6), S0=>nx17995);
   reg_flt_bias1_reg_q_7 : dff port map ( Q=>flt_bias_out_7, QB=>OPEN, D=>
      nx14241, CLK=>clk);
   ix14242 : mux21_ni port map ( Y=>nx14241, A0=>flt_bias_out_7, A1=>
      mem_data_in(7), S0=>nx17995);
   reg_flt_bias1_reg_q_8 : dff port map ( Q=>flt_bias_out_8, QB=>OPEN, D=>
      nx14261, CLK=>clk);
   ix14262 : mux21_ni port map ( Y=>nx14261, A0=>flt_bias_out_8, A1=>
      mem_data_in(8), S0=>nx17995);
   reg_flt_bias1_reg_q_9 : dff port map ( Q=>flt_bias_out_9, QB=>OPEN, D=>
      nx14281, CLK=>clk);
   ix14282 : mux21_ni port map ( Y=>nx14281, A0=>flt_bias_out_9, A1=>
      mem_data_in(9), S0=>nx17995);
   reg_flt_bias1_reg_q_10 : dff port map ( Q=>flt_bias_out_10, QB=>OPEN, D=>
      nx14301, CLK=>clk);
   ix14302 : mux21_ni port map ( Y=>nx14301, A0=>flt_bias_out_10, A1=>
      mem_data_in(10), S0=>nx17995);
   reg_flt_bias1_reg_q_11 : dff port map ( Q=>flt_bias_out_11, QB=>OPEN, D=>
      nx14321, CLK=>clk);
   ix14322 : mux21_ni port map ( Y=>nx14321, A0=>flt_bias_out_11, A1=>
      mem_data_in(11), S0=>nx17995);
   reg_flt_bias1_reg_q_12 : dff port map ( Q=>flt_bias_out_12, QB=>OPEN, D=>
      nx14341, CLK=>clk);
   ix14342 : mux21_ni port map ( Y=>nx14341, A0=>flt_bias_out_12, A1=>
      mem_data_in(12), S0=>nx2128);
   reg_flt_bias1_reg_q_13 : dff port map ( Q=>flt_bias_out_13, QB=>OPEN, D=>
      nx14361, CLK=>clk);
   ix14362 : mux21_ni port map ( Y=>nx14361, A0=>flt_bias_out_13, A1=>
      mem_data_in(13), S0=>nx2128);
   reg_flt_bias1_reg_q_14 : dff port map ( Q=>flt_bias_out_14, QB=>OPEN, D=>
      nx14381, CLK=>clk);
   ix14382 : mux21_ni port map ( Y=>nx14381, A0=>flt_bias_out_14, A1=>
      mem_data_in(14), S0=>nx2128);
   reg_flt_bias1_reg_q_15 : dff port map ( Q=>flt_bias_out_15, QB=>OPEN, D=>
      nx14401, CLK=>clk);
   ix14402 : mux21_ni port map ( Y=>nx14401, A0=>flt_bias_out_15, A1=>
      mem_data_in(15), S0=>nx2128);
   ix5153 : nor03_2x port map ( Y=>max_height_3, A0=>nx16042, A1=>nx17807, 
      A2=>nx17923);
   ix5157 : nor03_2x port map ( Y=>max_height_4, A0=>nx16055, A1=>nx17807, 
      A2=>nx17923);
   ix4861 : or02 port map ( Y=>cache_rst_actual, A0=>nx17809, A1=>reset);
   ix2619 : nand02 port map ( Y=>cache_load, A0=>nx16455, A1=>nx18081);
   ix14422 : mux21 port map ( Y=>nx14421, A0=>nx16459, A1=>nx16463, S0=>
      nx18047);
   ix16460 : aoi32 port map ( Y=>nx16459, A0=>nx1460, A1=>cache_height_ended, 
      A2=>nx17873, B0=>ftc_cntrl_reg_out_15, B1=>nx2566);
   ix2567 : nand03 port map ( Y=>nx2566, A0=>ftc_cntrl_reg_out_13, A1=>
      nx15605, A2=>nx17923);
   ftc_cntrl_reg_reg_q_15 : dffr port map ( Q=>ftc_cntrl_reg_out_15, QB=>
      nx16463, D=>nx14421, CLK=>nx17839, R=>nx17809);
   ix1183 : nor03_2x port map ( Y=>nx1182, A0=>ftc_cntrl_reg_out_12, A1=>
      nx18279, A2=>ftc_cntrl_reg_out_13);
   ix5143 : nand02 port map ( Y=>max_height_0, A0=>nx16507, A1=>
      img_width_out_0);
   ix5149 : nand02 port map ( Y=>max_height_2, A0=>nx16507, A1=>nx18055);
   ix2153 : oai21 port map ( Y=>comp_unit_data1_out(0), A0=>nx18063, A1=>
      nx16511, B0=>nx16514);
   bias1_reg_reg_q_0 : dffr port map ( Q=>OPEN, QB=>nx16511, D=>nx14111, CLK
      =>clk, R=>reset);
   ix16515 : nand02 port map ( Y=>nx16514, A0=>nx2140, A1=>nx17997);
   ix2179 : oai21 port map ( Y=>comp_unit_data1_out(1), A0=>nx18063, A1=>
      nx16518, B0=>nx16521);
   bias1_reg_reg_q_1 : dffr port map ( Q=>OPEN, QB=>nx16518, D=>nx14131, CLK
      =>clk, R=>reset);
   ix16522 : nand02 port map ( Y=>nx16521, A0=>nx2168, A1=>nx17997);
   ix2205 : oai21 port map ( Y=>comp_unit_data1_out(2), A0=>nx18063, A1=>
      nx16524, B0=>nx16527);
   bias1_reg_reg_q_2 : dffr port map ( Q=>OPEN, QB=>nx16524, D=>nx14151, CLK
      =>clk, R=>reset);
   ix16528 : nand02 port map ( Y=>nx16527, A0=>nx2194, A1=>nx17997);
   ix2231 : oai21 port map ( Y=>comp_unit_data1_out(3), A0=>nx18063, A1=>
      nx16530, B0=>nx16533);
   bias1_reg_reg_q_3 : dffr port map ( Q=>OPEN, QB=>nx16530, D=>nx14171, CLK
      =>clk, R=>reset);
   ix16534 : nand02 port map ( Y=>nx16533, A0=>nx2220, A1=>nx17997);
   ix2257 : oai21 port map ( Y=>comp_unit_data1_out(4), A0=>nx18065, A1=>
      nx16536, B0=>nx16539);
   bias1_reg_reg_q_4 : dffr port map ( Q=>OPEN, QB=>nx16536, D=>nx14191, CLK
      =>clk, R=>reset);
   ix16540 : nand02 port map ( Y=>nx16539, A0=>nx2246, A1=>nx17997);
   ix2283 : oai21 port map ( Y=>comp_unit_data1_out(5), A0=>nx18065, A1=>
      nx16542, B0=>nx16545);
   bias1_reg_reg_q_5 : dffr port map ( Q=>OPEN, QB=>nx16542, D=>nx14211, CLK
      =>clk, R=>reset);
   ix16546 : nand02 port map ( Y=>nx16545, A0=>nx2272, A1=>nx17997);
   ix2309 : oai21 port map ( Y=>comp_unit_data1_out(6), A0=>nx18065, A1=>
      nx16548, B0=>nx16551);
   bias1_reg_reg_q_6 : dffr port map ( Q=>OPEN, QB=>nx16548, D=>nx14231, CLK
      =>clk, R=>reset);
   ix16552 : nand02 port map ( Y=>nx16551, A0=>nx2298, A1=>nx17997);
   ix2335 : oai21 port map ( Y=>comp_unit_data1_out(7), A0=>nx18065, A1=>
      nx16554, B0=>nx16557);
   bias1_reg_reg_q_7 : dffr port map ( Q=>OPEN, QB=>nx16554, D=>nx14251, CLK
      =>clk, R=>reset);
   ix16558 : nand02 port map ( Y=>nx16557, A0=>nx2324, A1=>nx17999);
   ix2361 : oai21 port map ( Y=>comp_unit_data1_out(8), A0=>nx18065, A1=>
      nx16560, B0=>nx16563);
   bias1_reg_reg_q_8 : dffr port map ( Q=>OPEN, QB=>nx16560, D=>nx14271, CLK
      =>clk, R=>reset);
   ix16564 : nand02 port map ( Y=>nx16563, A0=>nx2350, A1=>nx17999);
   ix2387 : oai21 port map ( Y=>comp_unit_data1_out(9), A0=>nx18065, A1=>
      nx16566, B0=>nx16569);
   bias1_reg_reg_q_9 : dffr port map ( Q=>OPEN, QB=>nx16566, D=>nx14291, CLK
      =>clk, R=>reset);
   ix16570 : nand02 port map ( Y=>nx16569, A0=>nx2376, A1=>nx17999);
   ix2413 : oai21 port map ( Y=>comp_unit_data1_out(10), A0=>nx18067, A1=>
      nx16572, B0=>nx16575);
   bias1_reg_reg_q_10 : dffr port map ( Q=>OPEN, QB=>nx16572, D=>nx14311, 
      CLK=>clk, R=>reset);
   ix16576 : nand02 port map ( Y=>nx16575, A0=>nx2402, A1=>nx17999);
   ix2439 : oai21 port map ( Y=>comp_unit_data1_out(11), A0=>nx18067, A1=>
      nx16578, B0=>nx16581);
   bias1_reg_reg_q_11 : dffr port map ( Q=>OPEN, QB=>nx16578, D=>nx14331, 
      CLK=>clk, R=>reset);
   ix16582 : nand02 port map ( Y=>nx16581, A0=>nx2428, A1=>nx17999);
   ix2465 : oai21 port map ( Y=>comp_unit_data1_out(12), A0=>nx18067, A1=>
      nx16584, B0=>nx16587);
   bias1_reg_reg_q_12 : dffr port map ( Q=>OPEN, QB=>nx16584, D=>nx14351, 
      CLK=>clk, R=>reset);
   ix16588 : nand02 port map ( Y=>nx16587, A0=>nx2454, A1=>nx17999);
   ix2491 : oai21 port map ( Y=>comp_unit_data1_out(13), A0=>nx18067, A1=>
      nx16590, B0=>nx16593);
   bias1_reg_reg_q_13 : dffr port map ( Q=>OPEN, QB=>nx16590, D=>nx14371, 
      CLK=>clk, R=>reset);
   ix16594 : nand02 port map ( Y=>nx16593, A0=>nx2480, A1=>nx17999);
   ix2517 : oai21 port map ( Y=>comp_unit_data1_out(14), A0=>nx18067, A1=>
      nx16596, B0=>nx16599);
   bias1_reg_reg_q_14 : dffr port map ( Q=>OPEN, QB=>nx16596, D=>nx14391, 
      CLK=>clk, R=>reset);
   ix16600 : nand02 port map ( Y=>nx16599, A0=>nx2506, A1=>nx18001);
   ix2543 : oai21 port map ( Y=>comp_unit_data1_out(15), A0=>nx18067, A1=>
      nx16602, B0=>nx16605);
   bias1_reg_reg_q_15 : dffr port map ( Q=>OPEN, QB=>nx16602, D=>nx14411, 
      CLK=>clk, R=>reset);
   ix16606 : nand02 port map ( Y=>nx16605, A0=>nx2532, A1=>nx18001);
   ix2117 : oai21 port map ( Y=>comp_unit_ready, A0=>nx18273, A1=>nx196, B0
      =>nx16608);
   ix16609 : aoi21 port map ( Y=>nx16608, A0=>nx17971, A1=>nx18305, B0=>
      nx18233);
   ix16611 : nand03 port map ( Y=>nx16610, A0=>flt_size_out_0, A1=>nx15711, 
      A2=>flt_size_out_1);
   ix4883 : aoi21 port map ( Y=>mem_read_out, A0=>nx16715, A1=>nx16721, B0=>
      reset);
   ix16722 : nor04 port map ( Y=>nx16721, A0=>nx18003, A1=>nx17869, A2=>
      nx2754, A3=>nx2128);
   ix2755 : nand02 port map ( Y=>nx2754, A0=>nx16727, A1=>nx16729);
   ix16728 : nor04 port map ( Y=>nx16727, A0=>current_state_2, A1=>
      current_state_3, A2=>nx17895, A3=>current_state_5);
   ix16730 : nor04 port map ( Y=>nx16729, A0=>current_state_6, A1=>nx17907, 
      A2=>current_state_8, A3=>nx17899);
   ix4867 : aoi21 port map ( Y=>mem_write_out, A0=>nx18053, A1=>nx18883, B0
      =>reset);
   reg_current_state_28 : dffr port map ( Q=>OPEN, QB=>nx16732, D=>nx1946, 
      CLK=>nx17839, R=>reset);
   ix2779 : nand04 port map ( Y=>mem_addr_out(0), A0=>nx16736, A1=>nx16756, 
      A2=>nx16780, A3=>nx16788);
   ix16737 : aoi221 port map ( Y=>nx16736, A0=>nx16738, A1=>nx17855, B0=>
      addr1_data_0, B1=>nx18037, C0=>nx2740);
   ix16739 : oai21 port map ( Y=>nx16738, A0=>class_cntr_counter_out_0, A1=>
      nx18007, B0=>nx16747);
   ix14432 : oai33 port map ( Y=>nx14431, A0=>nx16742, A1=>nx2622, A2=>
      nx18069, B0=>nx16745, B1=>nx17887, B2=>nx17879);
   reg_write_base_reg_q_0 : dffr port map ( Q=>OPEN, QB=>nx16745, D=>nx14431, 
      CLK=>nx17839, R=>reset);
   reg_addr1_data_0 : dffr port map ( Q=>addr1_data_0, QB=>OPEN, D=>nx14481, 
      CLK=>clk, R=>reset);
   ix2767 : nand02 port map ( Y=>nx2766, A0=>nx16313, A1=>nx18121);
   ix2741 : nor02_2x port map ( Y=>nx2740, A0=>nx18883, A1=>nx16738);
   ix16757 : oai21 port map ( Y=>nx16756, A0=>img_addr_offset_0, A1=>
      img_base_addr_0, B0=>nx2724);
   reg_img_addr_offset_0 : dffr port map ( Q=>img_addr_offset_0, QB=>OPEN, D
      =>nx14471, CLK=>clk, R=>nx18031);
   ix2713 : or02 port map ( Y=>nx2712, A0=>nx12873, A1=>reset);
   img_base_addr_inst_reg_q_0 : dffs_ni port map ( Q=>img_base_addr_0, QB=>
      OPEN, D=>nx14461, CLK=>clk, S=>reset);
   reg_write_base_prev_reg_q_0 : dffr port map ( Q=>
      write_base_prev_data_out_0, QB=>nx16764, D=>nx14451, CLK=>clk, R=>
      reset);
   ix16769 : nand04 port map ( Y=>nx16768, A0=>nx16770, A1=>nx2678, A2=>
      nx16774, A3=>nx16776);
   ix2679 : nor02_2x port map ( Y=>nx2678, A0=>nx16302, A1=>nx2674);
   ix16777 : xnor2 port map ( Y=>nx16776, A0=>nflt_layer_temp_3, A1=>
      nflt_layer_out_3);
   ix2725 : aoi21 port map ( Y=>nx2724, A0=>img_base_addr_0, A1=>
      img_addr_offset_0, B0=>nx18085);
   ix16781 : oai21 port map ( Y=>nx16780, A0=>nx18007, A1=>
      bias_offset_data_out_0, B0=>nx2668);
   reg_bias_offset_reg_q_0 : dffr port map ( Q=>bias_offset_data_out_0, QB=>
      OPEN, D=>nx14441, CLK=>clk, R=>reset);
   ix2669 : aoi21 port map ( Y=>nx2668, A0=>bias_offset_data_out_0, A1=>
      nx18007, B0=>nx18135);
   ix16787 : nand02 port map ( Y=>nx16786, A0=>nx18233, A1=>nx18297);
   ix16789 : oai221 port map ( Y=>nx16788, A0=>nx18011, A1=>nx18229, B0=>
      write_offset_data_out_0, B1=>nx18007, C0=>nx16791);
   ix2885 : or02 port map ( Y=>mem_addr_out(1), A0=>nx2882, A1=>nx2822);
   ix2883 : oai222 port map ( Y=>nx2882, A0=>nx2874, A1=>nx18075, B0=>
      nx16810, B1=>nx18085, C0=>nx16835, C1=>nx18135);
   ix2875 : nand02 port map ( Y=>nx2874, A0=>nx16796, A1=>nx16738);
   ix16797 : xnor2 port map ( Y=>nx16796, A0=>nx16747, A1=>nx16798);
   reg_write_base_reg_q_1 : dffr port map ( Q=>write_base_data_out_1, QB=>
      nx16802, D=>nx14491, CLK=>nx17839, R=>reset);
   ix16805 : xnor2 port map ( Y=>nx16804, A0=>nx16806, A1=>nx16808);
   ix16807 : nand02 port map ( Y=>nx16806, A0=>new_size_squared_out_0, A1=>
      nx18009);
   ix16811 : xnor2 port map ( Y=>nx16810, A0=>nx16812, A1=>nx16814);
   ix16813 : nand02 port map ( Y=>nx16812, A0=>img_base_addr_0, A1=>
      img_addr_offset_0);
   img_base_addr_inst_reg_q_1 : dffs_ni port map ( Q=>img_base_addr_1, QB=>
      nx16818, D=>nx14521, CLK=>clk, S=>reset);
   ix16821 : aoi21 port map ( Y=>nx16820, A0=>write_base_prev_data_out_1, A1
      =>write_base_prev_data_out_0, B0=>nx16825);
   reg_write_base_prev_reg_q_1 : dffr port map ( Q=>
      write_base_prev_data_out_1, QB=>OPEN, D=>nx14511, CLK=>clk, R=>reset);
   ix16830 : oai21 port map ( Y=>nx16829, A0=>img_addr_offset_0, A1=>
      img_addr_offset_1, B0=>nx16831);
   ix16832 : nand02 port map ( Y=>nx16831, A0=>img_addr_offset_1, A1=>
      img_addr_offset_0);
   reg_img_addr_offset_1 : dffr port map ( Q=>img_addr_offset_1, QB=>nx16833, 
      D=>nx14531, CLK=>clk, R=>nx18031);
   ix16836 : xnor2 port map ( Y=>nx16835, A0=>nx16837, A1=>nx16839);
   ix16838 : nand02 port map ( Y=>nx16837, A0=>bias_offset_data_out_0, A1=>
      nx18009);
   reg_bias_offset_reg_q_1 : dffr port map ( Q=>bias_offset_data_out_1, QB=>
      nx16843, D=>nx14541, CLK=>clk, R=>reset);
   ix2823 : oai222 port map ( Y=>nx2822, A0=>nx16846, A1=>nx18139, B0=>
      nx16796, B1=>nx16857, C0=>nx16861, C1=>nx18143);
   ix16850 : oai21 port map ( Y=>nx16849, A0=>addr1_data_0, A1=>addr1_data_1, 
      B0=>nx16852);
   reg_addr1_data_1 : dffr port map ( Q=>addr1_data_1, QB=>nx16846, D=>
      nx14501, CLK=>clk, R=>reset);
   ix16853 : nand02 port map ( Y=>nx16852, A0=>addr1_data_1, A1=>
      addr1_data_0);
   ix16858 : aoi21 port map ( Y=>nx16857, A0=>nx2738, A1=>nx17855, B0=>
      nx17975);
   ix16862 : xnor2 port map ( Y=>nx16861, A0=>nx16791, A1=>nx16863);
   ix3031 : nand02 port map ( Y=>mem_addr_out(2), A0=>nx16868, A1=>nx16916);
   ix16869 : aoi222 port map ( Y=>nx16868, A0=>nx16870, A1=>nx17855, B0=>
      nx3016, B1=>nx18021, C0=>nx2996, C1=>nx18003);
   ix16871 : nor02_2x port map ( Y=>nx16870, A0=>nx2928, A1=>nx2874);
   ix2929 : xnor2 port map ( Y=>nx2928, A0=>nx2924, A1=>nx16874);
   ix2925 : oai22 port map ( Y=>nx2924, A0=>nx16747, A1=>nx16798, B0=>
      nx16332, B1=>nx16802);
   reg_write_base_reg_q_2 : dffr port map ( Q=>write_base_data_out_2, QB=>
      nx16878, D=>nx14551, CLK=>nx17839, R=>reset);
   ix16881 : xnor2 port map ( Y=>nx16880, A0=>nx16882, A1=>nx16885);
   ix3017 : xor2 port map ( Y=>nx3016, A0=>nx16888, A1=>nx16891);
   reg_bias_offset_reg_q_2 : dffr port map ( Q=>bias_offset_data_out_2, QB=>
      nx16895, D=>nx14601, CLK=>clk, R=>reset);
   ix2997 : xor2 port map ( Y=>nx2996, A0=>nx16898, A1=>nx16901);
   img_base_addr_inst_reg_q_2 : dffs_ni port map ( Q=>img_base_addr_2, QB=>
      nx16911, D=>nx14581, CLK=>clk, S=>reset);
   ix2975 : oai21 port map ( Y=>nx2974, A0=>nx16906, A1=>nx16825, B0=>nx2968
   );
   reg_write_base_prev_reg_q_2 : dffr port map ( Q=>
      write_base_prev_data_out_2, QB=>nx16906, D=>nx14571, CLK=>clk, R=>
      reset);
   reg_img_addr_offset_2 : dffr port map ( Q=>img_addr_offset_2, QB=>nx16915, 
      D=>nx14591, CLK=>clk, R=>nx18031);
   ix16917 : aoi222 port map ( Y=>nx16916, A0=>addr1_data_2, A1=>nx18037, B0
      =>nx2914, B1=>nx18017, C0=>nx2928, C1=>nx2932);
   reg_addr1_data_2 : dffr port map ( Q=>addr1_data_2, QB=>OPEN, D=>nx14561, 
      CLK=>clk, R=>reset);
   ix2943 : xnor2 port map ( Y=>nx2942, A0=>addr1_data_2, A1=>nx16852);
   ix2915 : xnor2 port map ( Y=>nx2914, A0=>nx2892, A1=>nx16924);
   ix2893 : oai22 port map ( Y=>nx2892, A0=>nx16791, A1=>nx16863, B0=>
      nx15756, B1=>nx16802);
   ix2643 : nand02 port map ( Y=>nx2642, A0=>nx18313, A1=>nx18053);
   ix3177 : nand02 port map ( Y=>mem_addr_out(3), A0=>nx16931, A1=>nx16973);
   ix16932 : aoi222 port map ( Y=>nx16931, A0=>nx17975, A1=>nx3074, B0=>
      nx3168, B1=>nx18003, C0=>nx3122, C1=>nx18021);
   ix16935 : aoi22 port map ( Y=>nx16934, A0=>class_cntr_counter_out_2, A1=>
      write_base_data_out_2, B0=>nx2924, B1=>nx2926);
   reg_write_base_reg_q_3 : dffs_ni port map ( Q=>write_base_data_out_3, QB
      =>nx16945, D=>nx14611, CLK=>nx17839, S=>reset);
   ix3051 : xnor2 port map ( Y=>nx3050, A0=>nx3046, A1=>nx16943);
   ix3169 : xnor2 port map ( Y=>nx3168, A0=>nx3132, A1=>nx16948);
   ix16949 : xnor2 port map ( Y=>nx16948, A0=>img_base_addr_3, A1=>
      img_addr_offset_3);
   img_base_addr_inst_reg_q_3 : dffr port map ( Q=>img_base_addr_3, QB=>OPEN, 
      D=>nx14651, CLK=>clk, R=>reset);
   ix3147 : xor2 port map ( Y=>nx3146, A0=>write_base_prev_data_out_3, A1=>
      nx16956);
   reg_write_base_prev_reg_q_3 : dffr port map ( Q=>
      write_base_prev_data_out_3, QB=>OPEN, D=>nx14641, CLK=>clk, R=>reset);
   ix16957 : nor03_2x port map ( Y=>nx16956, A0=>write_base_prev_data_out_0, 
      A1=>write_base_prev_data_out_1, A2=>write_base_prev_data_out_2);
   reg_img_addr_offset_3 : dffr port map ( Q=>img_addr_offset_3, QB=>OPEN, D
      =>nx14661, CLK=>clk, R=>nx18031);
   ix3161 : xnor2 port map ( Y=>nx3160, A0=>img_addr_offset_3, A1=>nx16962);
   ix16963 : nand03 port map ( Y=>nx16962, A0=>img_addr_offset_2, A1=>
      img_addr_offset_1, A2=>nx18027);
   ix3123 : xnor2 port map ( Y=>nx3122, A0=>nx3112, A1=>nx16967);
   reg_bias_offset_reg_q_3 : dffr port map ( Q=>bias_offset_data_out_3, QB=>
      OPEN, D=>nx14631, CLK=>clk, R=>reset);
   ix16974 : aoi322 port map ( Y=>nx16973, A0=>nx3076, A1=>nx16978, A2=>
      nx17855, B0=>addr1_data_3, B1=>nx18037, C0=>nx3060, C1=>nx18017);
   ix3077 : nand02 port map ( Y=>nx3076, A0=>nx16976, A1=>nx16870);
   ix16977 : xnor2 port map ( Y=>nx16976, A0=>nx16934, A1=>nx16937);
   reg_addr1_data_3 : dffr port map ( Q=>addr1_data_3, QB=>OPEN, D=>nx14621, 
      CLK=>clk, R=>reset);
   ix3093 : xnor2 port map ( Y=>nx3092, A0=>addr1_data_3, A1=>nx16983);
   ix16984 : nand03 port map ( Y=>nx16983, A0=>addr1_data_2, A1=>
      addr1_data_1, A2=>addr1_data_0);
   ix3061 : xor2 port map ( Y=>nx3060, A0=>nx16987, A1=>nx16990);
   ix3327 : nand02 port map ( Y=>mem_addr_out(4), A0=>nx16993, A1=>nx17047);
   ix16994 : aoi222 port map ( Y=>nx16993, A0=>nx16995, A1=>nx17855, B0=>
      nx3312, B1=>nx18021, C0=>nx3292, C1=>nx18003);
   ix3079 : nor02_2x port map ( Y=>nx3078, A0=>nx16870, A1=>nx16976);
   reg_write_base_reg_q_4 : dffr port map ( Q=>write_base_data_out_4, QB=>
      nx17002, D=>nx14671, CLK=>nx17839, R=>reset);
   ix17005 : xnor2 port map ( Y=>nx17004, A0=>nx17006, A1=>nx17009);
   ix3313 : xor2 port map ( Y=>nx3312, A0=>nx17013, A1=>nx17016);
   reg_bias_offset_reg_q_4 : dffr port map ( Q=>bias_offset_data_out_4, QB=>
      nx17021, D=>nx14721, CLK=>clk, R=>reset);
   ix859 : aoi21 port map ( Y=>nx858, A0=>nx15741, A1=>nx15735, B0=>nx852);
   ix3293 : xor2 port map ( Y=>nx3292, A0=>nx17023, A1=>nx17026);
   img_base_addr_inst_reg_q_4 : dffs_ni port map ( Q=>img_base_addr_4, QB=>
      nx17038, D=>nx14701, CLK=>clk, S=>reset);
   ix3271 : oai21 port map ( Y=>nx3270, A0=>nx17031, A1=>nx17035, B0=>nx3264
   );
   reg_write_base_prev_reg_q_4 : dffr port map ( Q=>OPEN, QB=>nx17031, D=>
      nx14691, CLK=>clk, R=>reset);
   ix17036 : nor04 port map ( Y=>nx17035, A0=>write_base_prev_data_out_0, A1
      =>write_base_prev_data_out_1, A2=>write_base_prev_data_out_2, A3=>
      write_base_prev_data_out_3);
   ix3265 : nand02 port map ( Y=>nx3264, A0=>nx17035, A1=>nx17031);
   ix3285 : aoi21 port map ( Y=>nx3284, A0=>nx17042, A1=>nx17044, B0=>nx3278
   );
   ix17043 : nand04 port map ( Y=>nx17042, A0=>img_addr_offset_3, A1=>
      img_addr_offset_2, A2=>img_addr_offset_1, A3=>nx18027);
   reg_img_addr_offset_4 : dffr port map ( Q=>img_addr_offset_4, QB=>nx17044, 
      D=>nx14711, CLK=>clk, R=>nx18031);
   ix17048 : aoi21 port map ( Y=>nx17047, A0=>nx3206, A1=>nx18017, B0=>
      nx3246);
   ix3207 : xnor2 port map ( Y=>nx3206, A0=>nx3184, A1=>nx17051);
   ix3247 : oai22 port map ( Y=>nx3246, A0=>nx16998, A1=>nx17054, B0=>
      nx17056, B1=>nx18139);
   ix17055 : aoi21 port map ( Y=>nx17054, A0=>nx3078, A1=>nx17855, B0=>
      nx17975);
   ix3239 : aoi21 port map ( Y=>nx3238, A0=>nx17060, A1=>nx17056, B0=>nx3232
   );
   ix17061 : nand04 port map ( Y=>nx17060, A0=>addr1_data_3, A1=>
      addr1_data_2, A2=>addr1_data_1, A3=>addr1_data_0);
   reg_addr1_data_4 : dffr port map ( Q=>addr1_data_4, QB=>nx17056, D=>
      nx14681, CLK=>clk, R=>reset);
   ix3469 : nand02 port map ( Y=>mem_addr_out(5), A0=>nx17065, A1=>nx17106);
   ix17066 : aoi222 port map ( Y=>nx17065, A0=>nx18543, A1=>nx17857, B0=>
      nx3454, B1=>nx18021, C0=>nx3434, C1=>nx18003);
   reg_write_base_reg_q_5 : dffs_ni port map ( Q=>write_base_data_out_5, QB
      =>nx17076, D=>nx14731, CLK=>nx17841, S=>reset);
   ix3347 : xnor2 port map ( Y=>nx3346, A0=>nx3342, A1=>nx17074);
   ix17078 : nand02 port map ( Y=>nx17077, A0=>write_base_data_out_4, A1=>
      nx3216);
   ix3455 : xnor2 port map ( Y=>nx3454, A0=>nx3444, A1=>nx17081);
   reg_bias_offset_reg_q_5 : dffr port map ( Q=>bias_offset_data_out_5, QB=>
      nx17085, D=>nx14781, CLK=>clk, R=>reset);
   ix3435 : xnor2 port map ( Y=>nx3434, A0=>nx3398, A1=>nx17089);
   img_base_addr_inst_reg_q_5 : dffr port map ( Q=>img_base_addr_5, QB=>OPEN, 
      D=>nx14761, CLK=>clk, R=>reset);
   ix3413 : xnor2 port map ( Y=>nx3412, A0=>write_base_prev_data_out_5, A1=>
      nx3264);
   reg_write_base_prev_reg_q_5 : dffr port map ( Q=>
      write_base_prev_data_out_5, QB=>OPEN, D=>nx14751, CLK=>clk, R=>reset);
   ix17101 : oai21 port map ( Y=>nx17100, A0=>nx3278, A1=>img_addr_offset_5, 
      B0=>nx17102);
   ix17103 : nand02 port map ( Y=>nx17102, A0=>img_addr_offset_5, A1=>nx3278
   );
   reg_img_addr_offset_5 : dffr port map ( Q=>img_addr_offset_5, QB=>nx17104, 
      D=>nx14771, CLK=>clk, R=>nx18031);
   ix17107 : aoi222 port map ( Y=>nx17106, A0=>addr1_data_5, A1=>nx18037, B0
      =>nx3366, B1=>nx3370, C0=>nx3356, C1=>nx18017);
   ix17111 : oai21 port map ( Y=>nx17110, A0=>nx3232, A1=>addr1_data_5, B0=>
      nx17112);
   ix17113 : nand02 port map ( Y=>nx17112, A0=>addr1_data_5, A1=>nx3232);
   reg_addr1_data_5 : dffr port map ( Q=>addr1_data_5, QB=>nx17114, D=>
      nx14741, CLK=>clk, R=>reset);
   ix3371 : oai21 port map ( Y=>nx3370, A0=>nx16995, A1=>nx18075, B0=>
      nx18883);
   ix3357 : xor2 port map ( Y=>nx3356, A0=>nx17118, A1=>nx17121);
   ix3611 : or02 port map ( Y=>mem_addr_out(6), A0=>nx3608, A1=>nx3532);
   ix3609 : oai222 port map ( Y=>nx3608, A0=>nx17125, A1=>nx18135, B0=>
      nx17147, B1=>nx18087, C0=>nx3600, C1=>nx18075);
   ix17126 : xnor2 port map ( Y=>nx17125, A0=>nx17127, A1=>nx17130);
   reg_bias_offset_reg_q_6 : dffr port map ( Q=>bias_offset_data_out_6, QB=>
      nx17135, D=>nx14841, CLK=>clk, R=>reset);
   ix905 : aoi21 port map ( Y=>nx904, A0=>nx15726, A1=>nx15720, B0=>nx898);
   reg_write_base_reg_q_6 : dffs_ni port map ( Q=>write_base_data_out_6, QB
      =>nx17138, D=>nx14791, CLK=>nx17841, S=>reset);
   ix17141 : xnor2 port map ( Y=>nx17140, A0=>nx17142, A1=>nx17145);
   ix17148 : xnor2 port map ( Y=>nx17147, A0=>nx17149, A1=>nx17152);
   img_base_addr_inst_reg_q_6 : dffs_ni port map ( Q=>img_base_addr_6, QB=>
      nx17164, D=>nx14821, CLK=>clk, S=>reset);
   ix3555 : oai21 port map ( Y=>nx3554, A0=>nx17157, A1=>nx17161, B0=>nx3548
   );
   reg_write_base_prev_reg_q_6 : dffr port map ( Q=>OPEN, QB=>nx17157, D=>
      nx14811, CLK=>clk, R=>reset);
   ix17162 : nor02_2x port map ( Y=>nx17161, A0=>nx3264, A1=>
      write_base_prev_data_out_5);
   ix3549 : nand02 port map ( Y=>nx3548, A0=>nx17161, A1=>nx17157);
   ix3569 : aoi21 port map ( Y=>nx3568, A0=>nx17102, A1=>nx17168, B0=>nx3562
   );
   reg_img_addr_offset_6 : dffr port map ( Q=>img_addr_offset_6, QB=>nx17168, 
      D=>nx14831, CLK=>clk, R=>nx18031);
   ix17176 : nand02 port map ( Y=>nx17175, A0=>write_base_data_out_6, A1=>
      nx3360);
   ix3533 : oai222 port map ( Y=>nx3532, A0=>nx17172, A1=>nx17178, B0=>
      nx17183, B1=>nx18143, C0=>nx17188, C1=>nx18139);
   ix17179 : aoi21 port map ( Y=>nx17178, A0=>nx3458, A1=>nx17857, B0=>
      nx17975);
   ix17184 : xor2 port map ( Y=>nx17183, A0=>nx18597, A1=>nx17186);
   reg_addr1_data_6 : dffr port map ( Q=>addr1_data_6, QB=>nx17188, D=>
      nx14801, CLK=>clk, R=>reset);
   ix3753 : nand02 port map ( Y=>mem_addr_out(7), A0=>nx17194, A1=>nx17235);
   ix17195 : aoi222 port map ( Y=>nx17194, A0=>nx17196, A1=>nx17857, B0=>
      nx3738, B1=>nx18021, C0=>nx3718, C1=>nx18003);
   ix3631 : xnor2 port map ( Y=>nx3630, A0=>nx3626, A1=>nx17204);
   reg_write_base_reg_q_7 : dffr port map ( Q=>write_base_data_out_7, QB=>
      nx17199, D=>nx14851, CLK=>nx17841, R=>reset);
   ix3739 : xnor2 port map ( Y=>nx3738, A0=>nx3728, A1=>nx17210);
   reg_bias_offset_reg_q_7 : dffr port map ( Q=>bias_offset_data_out_7, QB=>
      nx17214, D=>nx14901, CLK=>clk, R=>reset);
   ix3719 : xnor2 port map ( Y=>nx3718, A0=>nx18760, A1=>nx17218);
   img_base_addr_inst_reg_q_7 : dffr port map ( Q=>img_base_addr_7, QB=>OPEN, 
      D=>nx14881, CLK=>clk, R=>reset);
   ix3697 : xnor2 port map ( Y=>nx3696, A0=>write_base_prev_data_out_7, A1=>
      nx3548);
   reg_write_base_prev_reg_q_7 : dffr port map ( Q=>
      write_base_prev_data_out_7, QB=>OPEN, D=>nx14871, CLK=>clk, R=>reset);
   ix17230 : oai21 port map ( Y=>nx17229, A0=>nx3562, A1=>img_addr_offset_7, 
      B0=>nx17231);
   ix17232 : nand02 port map ( Y=>nx17231, A0=>img_addr_offset_7, A1=>nx3562
   );
   reg_img_addr_offset_7 : dffr port map ( Q=>img_addr_offset_7, QB=>nx17233, 
      D=>nx14891, CLK=>clk, R=>nx18033);
   ix17236 : aoi222 port map ( Y=>nx17235, A0=>addr1_data_7, A1=>nx18037, B0
      =>nx3640, B1=>nx18017, C0=>nx3650, C1=>nx3654);
   ix17240 : oai21 port map ( Y=>nx17239, A0=>nx3516, A1=>addr1_data_7, B0=>
      nx17242);
   ix17243 : nand02 port map ( Y=>nx17242, A0=>addr1_data_7, A1=>nx3516);
   reg_addr1_data_7 : dffr port map ( Q=>addr1_data_7, QB=>nx17244, D=>
      nx14861, CLK=>clk, R=>reset);
   ix3641 : xor2 port map ( Y=>nx3640, A0=>nx17247, A1=>nx17250);
   ix3895 : or02 port map ( Y=>mem_addr_out(8), A0=>nx3892, A1=>nx3816);
   ix3893 : oai222 port map ( Y=>nx3892, A0=>nx17255, A1=>nx18135, B0=>
      nx17277, B1=>nx18089, C0=>nx3884, C1=>nx18075);
   ix17256 : xnor2 port map ( Y=>nx17255, A0=>nx17257, A1=>nx17260);
   reg_bias_offset_reg_q_8 : dffr port map ( Q=>bias_offset_data_out_8, QB=>
      nx17265, D=>nx14961, CLK=>clk, R=>reset);
   ix955 : aoi21 port map ( Y=>nx954, A0=>nx15692, A1=>nx15686, B0=>nx948);
   reg_write_base_reg_q_8 : dffs_ni port map ( Q=>write_base_data_out_8, QB
      =>nx17268, D=>nx14911, CLK=>nx17841, S=>reset);
   ix17271 : xnor2 port map ( Y=>nx17270, A0=>nx17272, A1=>nx17275);
   ix17278 : xnor2 port map ( Y=>nx17277, A0=>nx17279, A1=>nx17282);
   img_base_addr_inst_reg_q_8 : dffr port map ( Q=>img_base_addr_8, QB=>
      nx17294, D=>nx14941, CLK=>clk, R=>reset);
   ix3839 : oai21 port map ( Y=>nx3838, A0=>nx17287, A1=>nx17291, B0=>nx3832
   );
   reg_write_base_prev_reg_q_8 : dffr port map ( Q=>OPEN, QB=>nx17287, D=>
      nx14931, CLK=>clk, R=>reset);
   ix17292 : nor02_2x port map ( Y=>nx17291, A0=>nx3548, A1=>
      write_base_prev_data_out_7);
   ix3833 : nand02 port map ( Y=>nx3832, A0=>nx17291, A1=>nx17287);
   ix3853 : aoi21 port map ( Y=>nx3852, A0=>nx17231, A1=>nx17298, B0=>nx3846
   );
   reg_img_addr_offset_8 : dffr port map ( Q=>img_addr_offset_8, QB=>nx17298, 
      D=>nx14951, CLK=>clk, R=>nx18033);
   ix3817 : oai222 port map ( Y=>nx3816, A0=>nx17307, A1=>nx18143, B0=>
      nx17302, B1=>nx17312, C0=>nx17315, C1=>nx18139);
   ix17308 : xor2 port map ( Y=>nx17307, A0=>nx3760, A1=>nx17310);
   ix17313 : aoi21 port map ( Y=>nx17312, A0=>nx3742, A1=>nx17857, B0=>
      nx17975);
   reg_addr1_data_8 : dffr port map ( Q=>addr1_data_8, QB=>nx17315, D=>
      nx14921, CLK=>clk, R=>reset);
   ix4037 : nand02 port map ( Y=>mem_addr_out(9), A0=>nx17321, A1=>nx17362);
   ix17322 : aoi222 port map ( Y=>nx17321, A0=>nx17323, A1=>nx17857, B0=>
      nx4022, B1=>nx18021, C0=>nx4002, C1=>nx18003);
   ix3915 : xnor2 port map ( Y=>nx3914, A0=>nx18694, A1=>nx17331);
   reg_write_base_reg_q_9 : dffs_ni port map ( Q=>write_base_data_out_9, QB
      =>nx17326, D=>nx14971, CLK=>nx17841, S=>reset);
   ix4023 : xnor2 port map ( Y=>nx4022, A0=>nx4012, A1=>nx17337);
   reg_bias_offset_reg_q_9 : dffr port map ( Q=>bias_offset_data_out_9, QB=>
      nx17341, D=>nx15021, CLK=>clk, R=>reset);
   ix4003 : xnor2 port map ( Y=>nx4002, A0=>nx3966, A1=>nx17345);
   img_base_addr_inst_reg_q_9 : dffr port map ( Q=>img_base_addr_9, QB=>OPEN, 
      D=>nx15001, CLK=>clk, R=>reset);
   ix3981 : xnor2 port map ( Y=>nx3980, A0=>write_base_prev_data_out_9, A1=>
      nx3832);
   reg_write_base_prev_reg_q_9 : dffr port map ( Q=>
      write_base_prev_data_out_9, QB=>OPEN, D=>nx14991, CLK=>clk, R=>reset);
   ix17357 : oai21 port map ( Y=>nx17356, A0=>nx3846, A1=>img_addr_offset_9, 
      B0=>nx17358);
   ix17359 : nand02 port map ( Y=>nx17358, A0=>img_addr_offset_9, A1=>nx3846
   );
   reg_img_addr_offset_9 : dffr port map ( Q=>img_addr_offset_9, QB=>nx17360, 
      D=>nx15011, CLK=>clk, R=>nx18033);
   ix17363 : aoi222 port map ( Y=>nx17362, A0=>addr1_data_9, A1=>nx18037, B0
      =>nx3924, B1=>nx18017, C0=>nx3934, C1=>nx3938);
   ix17367 : oai21 port map ( Y=>nx17366, A0=>nx3800, A1=>addr1_data_9, B0=>
      nx17369);
   ix17370 : nand02 port map ( Y=>nx17369, A0=>addr1_data_9, A1=>nx3800);
   reg_addr1_data_9 : dffr port map ( Q=>addr1_data_9, QB=>nx17371, D=>
      nx14981, CLK=>clk, R=>reset);
   ix3925 : xor2 port map ( Y=>nx3924, A0=>nx17374, A1=>nx17377);
   ix17375 : aoi22 port map ( Y=>nx17374, A0=>write_offset_data_out_8, A1=>
      nx18897, B0=>nx3760, B1=>nx3780);
   ix4179 : or02 port map ( Y=>mem_addr_out(10), A0=>nx4176, A1=>nx4100);
   ix4177 : oai222 port map ( Y=>nx4176, A0=>nx17382, A1=>nx18135, B0=>
      nx17404, B1=>nx18089, C0=>nx4168, C1=>nx18075);
   ix17383 : xnor2 port map ( Y=>nx17382, A0=>nx17384, A1=>nx17387);
   reg_bias_offset_reg_q_10 : dffr port map ( Q=>bias_offset_data_out_10, QB
      =>nx17392, D=>nx15081, CLK=>clk, R=>reset);
   ix1001 : aoi21 port map ( Y=>nx1000, A0=>nx15679, A1=>nx15673, B0=>nx994
   );
   reg_write_base_reg_q_10 : dffr port map ( Q=>write_base_data_out_10, QB=>
      nx17395, D=>nx15031, CLK=>nx17841, R=>reset);
   ix17398 : xnor2 port map ( Y=>nx17397, A0=>nx17399, A1=>nx17402);
   ix17405 : xnor2 port map ( Y=>nx17404, A0=>nx17406, A1=>nx17409);
   img_base_addr_inst_reg_q_10 : dffr port map ( Q=>img_base_addr_10, QB=>
      nx17421, D=>nx15061, CLK=>clk, R=>reset);
   ix4123 : oai21 port map ( Y=>nx4122, A0=>nx17414, A1=>nx17418, B0=>nx4116
   );
   reg_write_base_prev_reg_q_10 : dffr port map ( Q=>OPEN, QB=>nx17414, D=>
      nx15051, CLK=>clk, R=>reset);
   ix17419 : nor02_2x port map ( Y=>nx17418, A0=>nx3832, A1=>
      write_base_prev_data_out_9);
   ix4117 : nand02 port map ( Y=>nx4116, A0=>nx17418, A1=>nx17414);
   ix4137 : aoi21 port map ( Y=>nx4136, A0=>nx17358, A1=>nx17425, B0=>nx4130
   );
   reg_img_addr_offset_10 : dffr port map ( Q=>img_addr_offset_10, QB=>
      nx17425, D=>nx15071, CLK=>clk, R=>nx18033);
   ix4101 : oai222 port map ( Y=>nx4100, A0=>nx17434, A1=>nx18143, B0=>
      nx17429, B1=>nx17439, C0=>nx17442, C1=>nx18139);
   ix17435 : xor2 port map ( Y=>nx17434, A0=>nx4044, A1=>nx17437);
   ix4045 : oai22 port map ( Y=>nx4044, A0=>nx17374, A1=>nx17377, B0=>
      nx15770, B1=>nx17326);
   ix17440 : aoi21 port map ( Y=>nx17439, A0=>nx4026, A1=>nx17859, B0=>
      nx17977);
   reg_addr1_data_10 : dffr port map ( Q=>addr1_data_10, QB=>nx17442, D=>
      nx15041, CLK=>clk, R=>reset);
   ix4321 : nand02 port map ( Y=>mem_addr_out(11), A0=>nx17448, A1=>nx17489
   );
   ix17449 : aoi222 port map ( Y=>nx17448, A0=>nx17450, A1=>nx17859, B0=>
      nx4306, B1=>nx18023, C0=>nx4286, C1=>nx18005);
   ix4199 : xnor2 port map ( Y=>nx4198, A0=>nx4194, A1=>nx17458);
   reg_write_base_reg_q_11 : dffs_ni port map ( Q=>write_base_data_out_11, 
      QB=>nx17453, D=>nx15091, CLK=>nx17841, S=>reset);
   ix4307 : xnor2 port map ( Y=>nx4306, A0=>nx4296, A1=>nx17464);
   reg_bias_offset_reg_q_11 : dffr port map ( Q=>bias_offset_data_out_11, QB
      =>nx17468, D=>nx15141, CLK=>clk, R=>reset);
   ix4287 : xnor2 port map ( Y=>nx4286, A0=>nx4250, A1=>nx17472);
   img_base_addr_inst_reg_q_11 : dffs_ni port map ( Q=>img_base_addr_11, QB
      =>OPEN, D=>nx15121, CLK=>clk, S=>reset);
   ix4265 : xnor2 port map ( Y=>nx4264, A0=>write_base_prev_data_out_11, A1
      =>nx4116);
   reg_write_base_prev_reg_q_11 : dffr port map ( Q=>
      write_base_prev_data_out_11, QB=>OPEN, D=>nx15111, CLK=>clk, R=>reset
   );
   ix17484 : oai21 port map ( Y=>nx17483, A0=>nx4130, A1=>img_addr_offset_11, 
      B0=>nx17485);
   ix17486 : nand02 port map ( Y=>nx17485, A0=>img_addr_offset_11, A1=>
      nx4130);
   reg_img_addr_offset_11 : dffr port map ( Q=>img_addr_offset_11, QB=>
      nx17487, D=>nx15131, CLK=>clk, R=>nx18033);
   ix17490 : aoi222 port map ( Y=>nx17489, A0=>addr1_data_11, A1=>nx18037, 
      B0=>nx4218, B1=>nx4222, C0=>nx4208, C1=>nx18017);
   ix17494 : oai21 port map ( Y=>nx17493, A0=>nx4084, A1=>addr1_data_11, B0
      =>nx17496);
   ix17497 : nand02 port map ( Y=>nx17496, A0=>addr1_data_11, A1=>nx4084);
   reg_addr1_data_11 : dffr port map ( Q=>addr1_data_11, QB=>nx17498, D=>
      nx15101, CLK=>clk, R=>reset);
   ix4209 : xor2 port map ( Y=>nx4208, A0=>nx17502, A1=>nx17505);
   ix17510 : xnor2 port map ( Y=>nx17509, A0=>nx17511, A1=>nx17514);
   reg_bias_offset_reg_q_12 : dffr port map ( Q=>bias_offset_data_out_12, QB
      =>nx17519, D=>nx15201, CLK=>clk, R=>reset);
   ix1049 : aoi21 port map ( Y=>nx1048, A0=>nx15666, A1=>nx15660, B0=>nx1042
   );
   reg_write_base_reg_q_12 : dffs_ni port map ( Q=>write_base_data_out_12, 
      QB=>nx17522, D=>nx15151, CLK=>nx17843, S=>reset);
   img_base_addr_inst_reg_q_12 : dffs_ni port map ( Q=>img_base_addr_12, QB
      =>nx17548, D=>nx15181, CLK=>clk, S=>reset);
   ix4407 : oai21 port map ( Y=>nx4406, A0=>nx17541, A1=>nx17545, B0=>nx4400
   );
   reg_write_base_prev_reg_q_12 : dffr port map ( Q=>OPEN, QB=>nx17541, D=>
      nx15171, CLK=>clk, R=>reset);
   ix17546 : nor02_2x port map ( Y=>nx17545, A0=>nx4116, A1=>
      write_base_prev_data_out_11);
   ix4401 : nand02 port map ( Y=>nx4400, A0=>nx17545, A1=>nx17541);
   ix4421 : aoi21 port map ( Y=>nx4420, A0=>nx17485, A1=>nx17552, B0=>nx4414
   );
   reg_img_addr_offset_12 : dffr port map ( Q=>img_addr_offset_12, QB=>
      nx17552, D=>nx15191, CLK=>clk, R=>nx18033);
   ix17562 : xor2 port map ( Y=>nx17561, A0=>nx4328, A1=>nx17564);
   reg_addr1_data_12 : dffr port map ( Q=>addr1_data_12, QB=>nx17566, D=>
      nx15161, CLK=>clk, R=>reset);
   ix4605 : nand02 port map ( Y=>mem_addr_out(13), A0=>nx17575, A1=>nx17616
   );
   ix17576 : aoi222 port map ( Y=>nx17575, A0=>nx17577, A1=>nx17859, B0=>
      nx4590, B1=>nx18023, C0=>nx4570, C1=>nx18005);
   reg_write_base_reg_q_13 : dffr port map ( Q=>write_base_data_out_13, QB=>
      nx17580, D=>nx15211, CLK=>nx17843, R=>reset);
   ix4591 : xnor2 port map ( Y=>nx4590, A0=>nx18726, A1=>nx17591);
   reg_bias_offset_reg_q_13 : dffr port map ( Q=>bias_offset_data_out_13, QB
      =>nx17595, D=>nx15261, CLK=>clk, R=>reset);
   ix4571 : xnor2 port map ( Y=>nx4570, A0=>nx4534, A1=>nx17599);
   ix4535 : oai22 port map ( Y=>nx4534, A0=>nx18838, A1=>nx17536, B0=>
      nx17552, B1=>nx17548);
   img_base_addr_inst_reg_q_13 : dffr port map ( Q=>img_base_addr_13, QB=>
      OPEN, D=>nx15241, CLK=>clk, R=>reset);
   ix4549 : xnor2 port map ( Y=>nx4548, A0=>write_base_prev_data_out_13, A1
      =>nx4400);
   reg_write_base_prev_reg_q_13 : dffr port map ( Q=>
      write_base_prev_data_out_13, QB=>OPEN, D=>nx15231, CLK=>clk, R=>reset
   );
   ix17611 : oai21 port map ( Y=>nx17610, A0=>nx4414, A1=>img_addr_offset_13, 
      B0=>nx17612);
   ix17613 : nand02 port map ( Y=>nx17612, A0=>img_addr_offset_13, A1=>
      nx4414);
   reg_img_addr_offset_13 : dffr port map ( Q=>img_addr_offset_13, QB=>
      nx17614, D=>nx15251, CLK=>clk, R=>nx18033);
   ix17617 : aoi222 port map ( Y=>nx17616, A0=>addr1_data_13, A1=>nx18039, 
      B0=>nx4502, B1=>nx4506, C0=>nx4492, C1=>nx2642);
   ix17621 : oai21 port map ( Y=>nx17620, A0=>nx4368, A1=>addr1_data_13, B0
      =>nx17623);
   ix17624 : nand02 port map ( Y=>nx17623, A0=>addr1_data_13, A1=>nx4368);
   reg_addr1_data_13 : dffr port map ( Q=>addr1_data_13, QB=>nx17625, D=>
      nx15221, CLK=>clk, R=>reset);
   ix4493 : xor2 port map ( Y=>nx4492, A0=>nx17629, A1=>nx17632);
   ix4747 : or02 port map ( Y=>mem_addr_out(14), A0=>nx4744, A1=>nx4668);
   ix4745 : oai222 port map ( Y=>nx4744, A0=>nx17636, A1=>nx18135, B0=>
      nx17658, B1=>nx18091, C0=>nx4736, C1=>nx18339);
   ix17637 : xnor2 port map ( Y=>nx17636, A0=>nx17638, A1=>nx17641);
   reg_bias_offset_reg_q_14 : dffr port map ( Q=>bias_offset_data_out_14, QB
      =>nx17646, D=>nx15321, CLK=>clk, R=>reset);
   reg_write_base_reg_q_14 : dffr port map ( Q=>write_base_data_out_14, QB=>
      nx17649, D=>nx15271, CLK=>nx17843, R=>reset);
   ix17659 : xnor2 port map ( Y=>nx17658, A0=>nx17660, A1=>nx17663);
   ix17661 : aoi22 port map ( Y=>nx17660, A0=>img_addr_offset_13, A1=>
      img_base_addr_13, B0=>nx4534, B1=>nx4568);
   img_base_addr_inst_reg_q_14 : dffr port map ( Q=>img_base_addr_14, QB=>
      nx17673, D=>nx15301, CLK=>clk, R=>reset);
   reg_write_base_prev_reg_q_14 : dffr port map ( Q=>OPEN, QB=>nx17670, D=>
      nx15291, CLK=>clk, R=>reset);
   ix17672 : nor02_2x port map ( Y=>nx17671, A0=>nx4400, A1=>
      write_base_prev_data_out_13);
   reg_img_addr_offset_14 : dffr port map ( Q=>img_addr_offset_14, QB=>
      nx17677, D=>nx15311, CLK=>clk, R=>nx18035);
   ix4669 : oai222 port map ( Y=>nx4668, A0=>nx17682, A1=>nx18143, B0=>
      nx17687, B1=>nx18139, C0=>nx17679, C1=>nx17692);
   ix17683 : xor2 port map ( Y=>nx17682, A0=>nx18627, A1=>nx17685);
   reg_addr1_data_14 : dffr port map ( Q=>addr1_data_14, QB=>nx17687, D=>
      nx15281, CLK=>clk, R=>reset);
   ix17693 : aoi21 port map ( Y=>nx17692, A0=>nx4594, A1=>nx17859, B0=>
      nx17977);
   ix4859 : nand02 port map ( Y=>mem_addr_out(15), A0=>nx17696, A1=>nx17728
   );
   ix17697 : aoi222 port map ( Y=>nx17696, A0=>nx4816, A1=>nx18381, B0=>
      nx17977, B1=>nx4812, C0=>nx4850, C1=>nx18005);
   ix4817 : xnor2 port map ( Y=>nx4816, A0=>nx4736, A1=>nx4812);
   ix4813 : xnor2 port map ( Y=>nx4812, A0=>nx17700, A1=>
      write_base_data_out_15);
   ix17701 : nand02 port map ( Y=>nx17700, A0=>write_base_data_out_14, A1=>
      nx4496);
   reg_write_base_reg_q_15 : dffs_ni port map ( Q=>write_base_data_out_15, 
      QB=>OPEN, D=>nx15341, CLK=>nx17843, S=>reset);
   ix4851 : xnor2 port map ( Y=>nx4850, A0=>nx4826, A1=>nx17711);
   ix4827 : oai22 port map ( Y=>nx4826, A0=>nx17660, A1=>nx17663, B0=>
      nx17677, B1=>nx17673);
   img_base_addr_inst_reg_q_15 : dffs_ni port map ( Q=>img_base_addr_15, QB
      =>OPEN, D=>nx15371, CLK=>clk, S=>reset);
   ix4835 : xnor2 port map ( Y=>nx4834, A0=>write_base_prev_data_out_15, A1
      =>nx4684);
   reg_write_base_prev_reg_q_15 : dffr port map ( Q=>
      write_base_prev_data_out_15, QB=>OPEN, D=>nx15361, CLK=>clk, R=>reset
   );
   ix4685 : nand02 port map ( Y=>nx4684, A0=>nx17671, A1=>nx17670);
   img_addr_offset_15 : dffr port map ( Q=>OPEN, QB=>nx17726, D=>nx15381, 
      CLK=>clk, R=>nx18035);
   ix17729 : aoi222 port map ( Y=>nx17728, A0=>nx4804, A1=>nx2642, B0=>
      addr1_data_15, B1=>nx18039, C0=>nx4782, C1=>nx18023);
   ix4805 : xnor2 port map ( Y=>nx4804, A0=>nx17731, A1=>nx4802);
   reg_addr1_data_15 : dffr port map ( Q=>addr1_data_15, QB=>nx17740, D=>
      nx15351, CLK=>clk, R=>reset);
   ix4783 : xnor2 port map ( Y=>nx4782, A0=>nx4754, A1=>nx17744);
   ix4755 : oai22 port map ( Y=>nx4754, A0=>nx18725, A1=>nx17641, B0=>
      nx18915, B1=>nx17646);
   reg_bias_offset_reg_q_15 : dffr port map ( Q=>bias_offset_data_out_15, QB
      =>nx17748, D=>nx15331, CLK=>clk, R=>reset);
   ix1961 : inv01 port map ( Y=>mem_data_out(0), A=>nx17751);
   ix17752 : aoi222 port map ( Y=>nx17751, A0=>comp_unit_data2_in(0), A1=>
      nx17909, B0=>comp_unit_data1_in(0), B1=>nx17915, C0=>argmax_data_in(0), 
      C1=>nx17979);
   ix1971 : inv01 port map ( Y=>mem_data_out(1), A=>nx17754);
   ix17755 : aoi222 port map ( Y=>nx17754, A0=>comp_unit_data2_in(1), A1=>
      nx17909, B0=>comp_unit_data1_in(1), B1=>nx17915, C0=>argmax_data_in(1), 
      C1=>nx17979);
   ix1981 : inv01 port map ( Y=>mem_data_out(2), A=>nx17757);
   ix17758 : aoi222 port map ( Y=>nx17757, A0=>comp_unit_data2_in(2), A1=>
      nx17909, B0=>comp_unit_data1_in(2), B1=>nx17915, C0=>argmax_data_in(2), 
      C1=>nx17979);
   ix1991 : inv01 port map ( Y=>mem_data_out(3), A=>nx17760);
   ix17761 : aoi222 port map ( Y=>nx17760, A0=>comp_unit_data2_in(3), A1=>
      nx17909, B0=>comp_unit_data1_in(3), B1=>nx17915, C0=>argmax_data_in(3), 
      C1=>nx17979);
   ix2001 : inv01 port map ( Y=>mem_data_out(4), A=>nx17763);
   ix17764 : aoi222 port map ( Y=>nx17763, A0=>comp_unit_data2_in(4), A1=>
      nx17909, B0=>comp_unit_data1_in(4), B1=>nx17915, C0=>argmax_data_in(4), 
      C1=>nx17979);
   ix2011 : inv01 port map ( Y=>mem_data_out(5), A=>nx17766);
   ix17767 : aoi222 port map ( Y=>nx17766, A0=>comp_unit_data2_in(5), A1=>
      nx17909, B0=>comp_unit_data1_in(5), B1=>nx17917, C0=>argmax_data_in(5), 
      C1=>nx17979);
   ix2021 : inv01 port map ( Y=>mem_data_out(6), A=>nx17769);
   ix17770 : aoi222 port map ( Y=>nx17769, A0=>comp_unit_data2_in(6), A1=>
      nx17911, B0=>comp_unit_data1_in(6), B1=>nx17917, C0=>argmax_data_in(6), 
      C1=>nx17979);
   ix2031 : inv01 port map ( Y=>mem_data_out(7), A=>nx17772);
   ix17773 : aoi222 port map ( Y=>nx17772, A0=>comp_unit_data2_in(7), A1=>
      nx17911, B0=>comp_unit_data1_in(7), B1=>nx17917, C0=>argmax_data_in(7), 
      C1=>nx17981);
   ix2041 : inv01 port map ( Y=>mem_data_out(8), A=>nx17775);
   ix17776 : aoi222 port map ( Y=>nx17775, A0=>comp_unit_data2_in(8), A1=>
      nx17911, B0=>comp_unit_data1_in(8), B1=>nx17917, C0=>argmax_data_in(8), 
      C1=>nx17981);
   ix2051 : inv01 port map ( Y=>mem_data_out(9), A=>nx17778);
   ix17779 : aoi222 port map ( Y=>nx17778, A0=>comp_unit_data2_in(9), A1=>
      nx17911, B0=>comp_unit_data1_in(9), B1=>nx17917, C0=>argmax_data_in(9), 
      C1=>nx17981);
   ix2061 : inv01 port map ( Y=>mem_data_out(10), A=>nx17781);
   ix17782 : aoi222 port map ( Y=>nx17781, A0=>comp_unit_data2_in(10), A1=>
      nx17911, B0=>comp_unit_data1_in(10), B1=>nx17917, C0=>
      argmax_data_in(10), C1=>nx17981);
   ix2071 : inv01 port map ( Y=>mem_data_out(11), A=>nx17784);
   ix17785 : aoi222 port map ( Y=>nx17784, A0=>comp_unit_data2_in(11), A1=>
      nx17911, B0=>comp_unit_data1_in(11), B1=>nx17917, C0=>
      argmax_data_in(11), C1=>nx17981);
   ix2081 : inv01 port map ( Y=>mem_data_out(12), A=>nx17787);
   ix17788 : aoi222 port map ( Y=>nx17787, A0=>comp_unit_data2_in(12), A1=>
      nx17911, B0=>comp_unit_data1_in(12), B1=>nx17919, C0=>
      argmax_data_in(12), C1=>nx17981);
   ix2091 : inv01 port map ( Y=>mem_data_out(13), A=>nx17790);
   ix17791 : aoi222 port map ( Y=>nx17790, A0=>comp_unit_data2_in(13), A1=>
      nx17913, B0=>comp_unit_data1_in(13), B1=>nx17919, C0=>
      argmax_data_in(13), C1=>nx17981);
   ix2101 : inv01 port map ( Y=>mem_data_out(14), A=>nx17793);
   ix17794 : aoi222 port map ( Y=>nx17793, A0=>comp_unit_data2_in(14), A1=>
      nx17913, B0=>comp_unit_data1_in(14), B1=>nx17919, C0=>
      argmax_data_in(14), C1=>nx17983);
   ix2111 : inv01 port map ( Y=>mem_data_out(15), A=>nx17796);
   ix17797 : aoi222 port map ( Y=>nx17796, A0=>comp_unit_data2_in(15), A1=>
      nx17913, B0=>comp_unit_data1_in(15), B1=>nx17919, C0=>
      argmax_data_in(15), C1=>nx17983);
   ix4595 : inv01 port map ( Y=>nx4594, A=>nx17577);
   ix4569 : inv01 port map ( Y=>nx4568, A=>nx17599);
   ix4027 : inv01 port map ( Y=>nx4026, A=>nx17323);
   ix3781 : inv01 port map ( Y=>nx3780, A=>nx17310);
   ix3743 : inv01 port map ( Y=>nx3742, A=>nx17196);
   ix3459 : inv01 port map ( Y=>nx3458, A=>nx18543);
   ix16979 : inv01 port map ( Y=>nx16978, A=>nx3078);
   ix3075 : inv01 port map ( Y=>nx3074, A=>nx16976);
   ix3049 : inv01 port map ( Y=>nx3048, A=>nx16943);
   ix2969 : inv01 port map ( Y=>nx2968, A=>nx16956);
   ix2927 : inv01 port map ( Y=>nx2926, A=>nx16874);
   ix2739 : inv01 port map ( Y=>nx2738, A=>nx16738);
   ix2665 : inv01 port map ( Y=>nx2664, A=>nx16786);
   ix2623 : inv01 port map ( Y=>nx2622, A=>nx16806);
   ix16630 : inv01 port map ( Y=>nx16629, A=>nx2546);
   ix1803 : inv01 port map ( Y=>nx12910, A=>nx16282);
   ix1681 : inv01 port map ( Y=>nx12908, A=>nx16265);
   ix1461 : inv01 port map ( Y=>nx1460, A=>nx15609);
   ix15620 : inv01 port map ( Y=>nx15619, A=>nx1182);
   ix781 : inv01 port map ( Y=>nx780, A=>nx15765);
   ix637 : inv01 port map ( Y=>nx636, A=>nx16189);
   ix631 : inv01 port map ( Y=>nx630, A=>nx16191);
   ix583 : inv01 port map ( Y=>nx582, A=>nx15479);
   ix15975 : inv01 port map ( Y=>nx15974, A=>nx576);
   ix15397 : inv01 port map ( Y=>nx15396, A=>nx316);
   ix1859 : inv01 port map ( Y=>nx12877, A=>nx16204);
   ix15423 : inv01 port map ( Y=>nx15422, A=>nx12875);
   ix149 : inv01 port map ( Y=>nx148, A=>nx15533);
   ix303 : inv01 port map ( Y=>comp_unit_flt_size_EXMPLR, A=>nx16610);
   ix17802 : inv01 port map ( Y=>nx17803, A=>current_state_13);
   ix17804 : inv02 port map ( Y=>nx17805, A=>nx17803);
   ix17806 : inv02 port map ( Y=>nx17807, A=>nx17803);
   ix17808 : inv02 port map ( Y=>nx17809, A=>nx17803);
   ix17810 : buf02 port map ( Y=>nx17811, A=>wind_width_count_0);
   ix17812 : buf02 port map ( Y=>nx17813, A=>wind_width_count_0);
   ix17814 : buf02 port map ( Y=>nx17815, A=>cache_width_count_4);
   ix17816 : buf02 port map ( Y=>nx17817, A=>cache_width_count_4);
   ix17818 : buf02 port map ( Y=>nx17819, A=>cache_width_count_2);
   ix17820 : buf02 port map ( Y=>nx17821, A=>cache_width_count_2);
   ix17822 : inv02 port map ( Y=>nx17823, A=>clk);
   ix17824 : inv02 port map ( Y=>nx17825, A=>clk);
   ix17826 : inv02 port map ( Y=>nx17827, A=>clk);
   ix17828 : inv02 port map ( Y=>nx17829, A=>clk);
   ix17830 : inv02 port map ( Y=>nx17831, A=>clk);
   ix17832 : inv02 port map ( Y=>nx17833, A=>clk);
   ix17834 : inv02 port map ( Y=>nx17835, A=>clk);
   ix17836 : inv02 port map ( Y=>nx17837, A=>clk);
   ix17838 : inv02 port map ( Y=>nx17839, A=>clk);
   ix17840 : inv02 port map ( Y=>nx17841, A=>clk);
   ix17842 : inv02 port map ( Y=>nx17843, A=>clk);
   ix17844 : inv02 port map ( Y=>nx17845, A=>nx18305);
   ix17846 : inv02 port map ( Y=>nx17847, A=>nx18305);
   ix17854 : inv02 port map ( Y=>nx17855, A=>nx18339);
   ix17856 : inv02 port map ( Y=>nx17857, A=>nx18339);
   ix17858 : inv02 port map ( Y=>nx17859, A=>nx18339);
   ix17862 : inv01 port map ( Y=>nx17863, A=>filter_ready_out_EXMPLR);
   ix17864 : inv02 port map ( Y=>nx17865, A=>nx18319);
   ix17868 : inv02 port map ( Y=>nx17869, A=>nx18319);
   ix17870 : inv02 port map ( Y=>nx17871, A=>nx15605);
   ix17872 : inv02 port map ( Y=>nx17873, A=>nx15605);
   ix17874 : inv02 port map ( Y=>nx17875, A=>nx18333);
   ix17876 : inv02 port map ( Y=>nx17877, A=>nx18333);
   ix17878 : inv02 port map ( Y=>nx17879, A=>nx18333);
   ix17886 : inv02 port map ( Y=>nx17887, A=>nx15530);
   ix17892 : buf02 port map ( Y=>nx17893, A=>current_state_4);
   ix17894 : buf02 port map ( Y=>nx17895, A=>current_state_4);
   ix17896 : inv02 port map ( Y=>nx17897, A=>nx15435);
   ix17898 : inv02 port map ( Y=>nx17899, A=>nx15435);
   ix17906 : inv02 port map ( Y=>nx17907, A=>nx18323);
   ix17908 : inv02 port map ( Y=>nx17909, A=>nx15716);
   ix17910 : inv02 port map ( Y=>nx17911, A=>nx15716);
   ix17912 : inv02 port map ( Y=>nx17913, A=>nx15716);
   ix17914 : inv02 port map ( Y=>nx17915, A=>nx15541);
   ix17916 : inv02 port map ( Y=>nx17917, A=>nx15541);
   ix17918 : inv02 port map ( Y=>nx17919, A=>nx15541);
   ix17920 : inv02 port map ( Y=>nx17921, A=>nx15626);
   ix17922 : inv02 port map ( Y=>nx17923, A=>nx18279);
   ix17926 : inv02 port map ( Y=>nx17927, A=>nx15392);
   ix17928 : buf02 port map ( Y=>nx17929, A=>nx206);
   ix17936 : inv01 port map ( Y=>nx17937, A=>nx378);
   ix17938 : inv02 port map ( Y=>nx17939, A=>nx17937);
   ix17940 : inv02 port map ( Y=>nx17941, A=>nx17937);
   ix17942 : inv02 port map ( Y=>nx17943, A=>nx17937);
   ix17946 : inv02 port map ( Y=>nx17947, A=>nx17945);
   ix17948 : inv02 port map ( Y=>nx17949, A=>nx18329);
   ix17950 : inv02 port map ( Y=>nx17951, A=>nx18329);
   ix17958 : inv01 port map ( Y=>nx17959, A=>nx1224);
   ix17960 : inv02 port map ( Y=>nx17961, A=>nx17959);
   ix17962 : inv02 port map ( Y=>nx17963, A=>nx17959);
   ix17964 : inv02 port map ( Y=>nx17965, A=>nx17959);
   ix17970 : inv02 port map ( Y=>nx17971, A=>nx15554);
   ix17972 : buf02 port map ( Y=>nx17973, A=>nx1546);
   ix17974 : inv02 port map ( Y=>nx17975, A=>nx16732);
   ix17978 : inv02 port map ( Y=>nx17979, A=>nx18883);
   ix17980 : inv02 port map ( Y=>nx17981, A=>nx18884);
   ix17982 : inv02 port map ( Y=>nx17983, A=>nx18884);
   ix17992 : nor02_2x port map ( Y=>nx17993, A0=>nx16302, A1=>nx18153);
   ix17994 : nor02_2x port map ( Y=>nx17995, A0=>nx16302, A1=>nx18153);
   ix17996 : inv02 port map ( Y=>nx17997, A=>nx18117);
   ix17998 : inv02 port map ( Y=>nx17999, A=>nx18117);
   ix18000 : inv02 port map ( Y=>nx18001, A=>nx18117);
   ix18002 : inv02 port map ( Y=>nx18003, A=>nx18091);
   ix18004 : inv02 port map ( Y=>nx18005, A=>nx18091);
   ix18006 : inv02 port map ( Y=>nx18007, A=>nx16745);
   ix18010 : inv02 port map ( Y=>nx18011, A=>nx16927);
   ix18016 : inv02 port map ( Y=>nx18017, A=>nx18143);
   ix18020 : inv02 port map ( Y=>nx18021, A=>nx18137);
   ix18022 : inv02 port map ( Y=>nx18023, A=>nx18137);
   ix18026 : buf02 port map ( Y=>nx18027, A=>img_addr_offset_0);
   ix18028 : inv01 port map ( Y=>nx18029, A=>nx2712);
   ix18030 : inv02 port map ( Y=>nx18031, A=>nx18029);
   ix18032 : inv02 port map ( Y=>nx18033, A=>nx18029);
   ix18034 : inv02 port map ( Y=>nx18035, A=>nx18029);
   ix18036 : inv02 port map ( Y=>nx18037, A=>nx18141);
   ix18038 : inv02 port map ( Y=>nx18039, A=>nx18141);
   ix18040 : inv02 port map ( Y=>nx18041, A=>nx18911);
   ix18044 : buf02 port map ( Y=>nx18045, A=>nx15630);
   ix18046 : buf02 port map ( Y=>nx18047, A=>nx15630);
   ix18048 : inv02 port map ( Y=>nx18049, A=>nx760);
   ix18050 : inv02 port map ( Y=>nx18051, A=>nx18229);
   ix18052 : inv02 port map ( Y=>nx18053, A=>nx18229);
   ix18054 : buf02 port map ( Y=>nx18055, A=>nx16028);
   ix18058 : inv01 port map ( Y=>nx18059, A=>current_state_18);
   ix18062 : inv01 port map ( Y=>nx18063, A=>nx18233);
   ix18064 : inv01 port map ( Y=>nx18065, A=>nx18233);
   ix18066 : inv01 port map ( Y=>nx18067, A=>nx18233);
   ix18068 : inv02 port map ( Y=>nx18069, A=>nx19308);
   ix18076 : inv02 port map ( Y=>nx18077, A=>nx18381);
   ix18080 : inv02 port map ( Y=>nx18081, A=>nx2580);
   ix18084 : inv02 port map ( Y=>nx18085, A=>nx18243);
   ix18086 : inv02 port map ( Y=>nx18087, A=>nx18243);
   ix18088 : inv02 port map ( Y=>nx18089, A=>nx18243);
   ix18090 : inv02 port map ( Y=>nx18091, A=>nx18243);
   ix18116 : inv02 port map ( Y=>nx18117, A=>nx2142);
   ix18120 : inv02 port map ( Y=>nx18121, A=>nx18119);
   ix18136 : inv02 port map ( Y=>nx18137, A=>nx2664);
   ix18138 : inv02 port map ( Y=>nx18139, A=>nx2766);
   ix18140 : inv02 port map ( Y=>nx18141, A=>nx2766);
   ix18142 : inv02 port map ( Y=>nx18143, A=>nx2642);
   ix18150 : buf02 port map ( Y=>nx18151, A=>comp_unit_operation_EXMPLR);
   ix18152 : buf02 port map ( Y=>nx18153, A=>comp_unit_operation_EXMPLR);
   ix18154 : inv01 port map ( Y=>nx18155, A=>nx18385);
   ix18156 : inv01 port map ( Y=>nx18157, A=>nx18385);
   ix311 : xnor2 port map ( Y=>nx310, A0=>nx15591, A1=>nx308);
   ix13012 : mux21_ni port map ( Y=>nx13011, A0=>nx262, A1=>
      cntr1_inst_counter_out_4, S0=>nx18255);
   ix263 : xor2 port map ( Y=>nx262, A0=>nx15591, A1=>nx15402);
   ix13002 : mux21_ni port map ( Y=>nx13001, A0=>nx244, A1=>
      cntr1_inst_counter_out_3, S0=>nx18255);
   ix12992 : mux21_ni port map ( Y=>nx12991, A0=>nx230, A1=>
      cntr1_inst_counter_out_2, S0=>nx18255);
   ix12982 : mux21 port map ( Y=>nx12981, A0=>nx16307, A1=>nx15416, S0=>
      nx18255);
   ix207 : nand02 port map ( Y=>nx206, A0=>nx16313, A1=>nx17803);
   ix141 : nor02ii port map ( Y=>nx140, A0=>nx15450, A1=>io_ready_in);
   ix1797 : and03 port map ( Y=>nx1796, A0=>nx12873, A1=>nx15486, A2=>
      nx18163);
   ix18162 : inv01 port map ( Y=>nx18163, A=>nx16269);
   ix15480 : and02 port map ( Y=>nx15479, A0=>nx15435, A1=>nx18333);
   ix93 : nor02ii port map ( Y=>nx92, A0=>nx15486, A1=>nx12873);
   ix15487 : and04 port map ( Y=>nx15486, A0=>nflt_layer_out_0, A1=>nx15500, 
      A2=>nx15512, A3=>nx18165);
   ix18164 : inv01 port map ( Y=>nx18165, A=>nflt_layer_out_3);
   ix15492 : mux21 port map ( Y=>nx15491, A0=>nx15488, A1=>mem_data_in(0), 
      S0=>nx17893);
   ix15497 : nor02ii port map ( Y=>nx15496, A0=>nx17893, A1=>nx18265);
   ix15507 : and02 port map ( Y=>nx15506, A0=>nx15488, A1=>nx15500);
   ix15517 : xor2 port map ( Y=>nx15516, A0=>nx15512, A1=>nx15506);
   ix15526 : and03 port map ( Y=>nx15525, A0=>nx15488, A1=>nx15500, A2=>
      nx15512);
   ix15534 : and03 port map ( Y=>nx15533, A0=>nx15445, A1=>nx15435, A2=>
      nx19302);
   ix15547 : nor02ii port map ( Y=>nx15546, A0=>nx18151, A1=>
      layer_type_out_1);
   ix1479 : ao32 port map ( Y=>nx1478, A0=>nx15575, A1=>current_state_15, A2
      =>nx15883, B0=>current_state_16, B1=>ftc_cntrl_reg_out_11);
   ix15562 : or02 port map ( Y=>nx15561, A0=>ftc_cntrl_reg_out_14, A1=>
      nx18305);
   ix279 : xor2 port map ( Y=>nx278, A0=>nx18257, A1=>
      cntr1_inst_counter_out_2);
   ix277 : xnor2 port map ( Y=>nx276, A0=>nx18257, A1=>nx15586);
   ix13022 : mux21 port map ( Y=>nx13021, A0=>nx15588, A1=>nx15586, S0=>
      nx18257);
   ix15589 : xor2 port map ( Y=>nx15588, A0=>nx15586, A1=>nx12882);
   ix269 : nor02ii port map ( Y=>nx12882, A0=>nx15402, A1=>
      cntr1_inst_counter_out_4);
   ix15597 : xnor2 port map ( Y=>nx15596, A0=>nx18257, A1=>
      cntr1_inst_counter_out_1);
   ix15603 : nor02ii port map ( Y=>nx15602, A0=>nx12912, A1=>nx15861);
   ix1847 : nor02ii port map ( Y=>nx12912, A0=>nx15605, A1=>nx15621);
   ix1403 : and04 port map ( Y=>nx1402, A0=>nx15614, A1=>nx16070, A2=>
      nx16079, A3=>nx16084);
   ix13842 : mux21 port map ( Y=>nx13841, A0=>nx16067, A1=>nx15614, S0=>
      nx18289);
   ix349 : nor02ii port map ( Y=>nx12883, A0=>nx18279, A1=>nx15859);
   ix15631 : and04 port map ( Y=>nx15630, A0=>nx16153, A1=>nx15861, A2=>
      nx15888, A3=>nx15970);
   ix15641 : xor2 port map ( Y=>nx15640, A0=>nx15776, A1=>
      new_size_squared_out_15);
   ix15645 : xor2 port map ( Y=>nx15644, A0=>nx15776, A1=>nx1088);
   ix1089 : nor02ii port map ( Y=>nx1088, A0=>nx15653, A1=>
      write_offset_data_out_14);
   ix13632 : ao22 port map ( Y=>nx13631, A0=>nx1094, A1=>nx18229, B0=>
      write_offset_data_out_14, B1=>nx18329);
   ix1043 : nor02ii port map ( Y=>nx1042, A0=>nx15666, A1=>
      write_offset_data_out_12);
   ix13592 : ao22 port map ( Y=>nx13591, A0=>nx1048, A1=>nx18229, B0=>
      write_offset_data_out_12, B1=>nx18329);
   ix995 : nor02ii port map ( Y=>nx994, A0=>nx15679, A1=>
      write_offset_data_out_10);
   ix13552 : ao22 port map ( Y=>nx13551, A0=>nx1000, A1=>nx18229, B0=>
      write_offset_data_out_10, B1=>nx18329);
   ix949 : nor02ii port map ( Y=>nx948, A0=>nx15692, A1=>
      write_offset_data_out_8);
   ix13512 : ao22 port map ( Y=>nx13511, A0=>nx954, A1=>nx18231, B0=>
      write_offset_data_out_8, B1=>nx18329);
   ix763 : nor02ii port map ( Y=>nx17945, A0=>nx18231, A1=>nx15537);
   ix15700 : nand02 port map ( Y=>nx760, A0=>nx15541, A1=>nx15716);
   ix1525 : nor02_2x port map ( Y=>nx1524, A0=>nx15541, A1=>nx18305);
   ix899 : nor02ii port map ( Y=>nx898, A0=>nx15726, A1=>
      write_offset_data_out_6);
   ix13472 : ao22 port map ( Y=>nx13471, A0=>nx904, A1=>nx18231, B0=>
      write_offset_data_out_6, B1=>nx18329);
   ix853 : nor02ii port map ( Y=>nx852, A0=>nx15741, A1=>
      write_offset_data_out_4);
   ix13432 : ao22 port map ( Y=>nx13431, A0=>write_offset_data_out_4, A1=>
      nx18331, B0=>nx858, B1=>nx18231);
   ix15742 : or04 port map ( Y=>nx15741, A0=>nx15745, A1=>nx15750, A2=>
      nx15756, A3=>nx15763);
   ix13412 : ao22 port map ( Y=>nx13411, A0=>write_offset_data_out_3, A1=>
      nx18331, B0=>nx832, B1=>nx18231);
   ix13352 : mux21_ni port map ( Y=>nx13351, A0=>nx18331, A1=>nx18231, S0=>
      nx15763);
   ix15766 : or02 port map ( Y=>nx15765, A0=>nx15756, A1=>nx15763);
   ix15769 : or03 port map ( Y=>nx15768, A0=>nx15750, A1=>nx15756, A2=>
      nx15763);
   ix13662 : mux21_ni port map ( Y=>nx13661, A0=>mem_data_in(15), A1=>
      new_size_squared_out_15, S0=>nx18323);
   ix15782 : xnor2 port map ( Y=>nx15781, A0=>nx15647, A1=>nx15785);
   ix13642 : mux21_ni port map ( Y=>nx13641, A0=>mem_data_in(14), A1=>
      new_size_squared_out_14, S0=>nx18323);
   ix15787 : xor2 port map ( Y=>nx15786, A0=>nx15774, A1=>
      new_size_squared_out_13);
   ix13622 : mux21_ni port map ( Y=>nx13621, A0=>mem_data_in(13), A1=>
      new_size_squared_out_13, S0=>nx18323);
   ix15792 : xnor2 port map ( Y=>nx15791, A0=>nx15660, A1=>nx15795);
   ix13602 : mux21_ni port map ( Y=>nx13601, A0=>mem_data_in(12), A1=>
      new_size_squared_out_12, S0=>nx18323);
   ix15798 : xor2 port map ( Y=>nx15797, A0=>nx15772, A1=>
      new_size_squared_out_11);
   ix13582 : mux21_ni port map ( Y=>nx13581, A0=>mem_data_in(11), A1=>
      new_size_squared_out_11, S0=>nx18323);
   ix15803 : xnor2 port map ( Y=>nx15802, A0=>nx15673, A1=>nx15806);
   ix13562 : mux21_ni port map ( Y=>nx13561, A0=>mem_data_in(10), A1=>
      new_size_squared_out_10, S0=>nx18323);
   ix15808 : xor2 port map ( Y=>nx15807, A0=>nx15770, A1=>
      new_size_squared_out_9);
   ix13542 : mux21_ni port map ( Y=>nx13541, A0=>mem_data_in(9), A1=>
      new_size_squared_out_9, S0=>nx18325);
   ix15813 : xnor2 port map ( Y=>nx15812, A0=>nx15686, A1=>nx15816);
   ix13522 : mux21_ni port map ( Y=>nx13521, A0=>mem_data_in(8), A1=>
      new_size_squared_out_8, S0=>nx18325);
   ix15819 : xor2 port map ( Y=>nx15818, A0=>nx15696, A1=>
      new_size_squared_out_7);
   ix13502 : mux21_ni port map ( Y=>nx13501, A0=>mem_data_in(7), A1=>
      new_size_squared_out_7, S0=>nx18325);
   ix15824 : xnor2 port map ( Y=>nx15823, A0=>nx15720, A1=>nx15827);
   ix13482 : mux21_ni port map ( Y=>nx13481, A0=>mem_data_in(6), A1=>
      new_size_squared_out_6, S0=>nx18325);
   ix15829 : xor2 port map ( Y=>nx15828, A0=>nx15730, A1=>
      new_size_squared_out_5);
   ix13462 : mux21_ni port map ( Y=>nx13461, A0=>mem_data_in(5), A1=>
      new_size_squared_out_5, S0=>nx18325);
   ix15834 : xnor2 port map ( Y=>nx15833, A0=>nx15735, A1=>nx15837);
   ix13442 : mux21_ni port map ( Y=>nx13441, A0=>mem_data_in(4), A1=>
      new_size_squared_out_4, S0=>nx18325);
   ix15840 : xor2 port map ( Y=>nx15839, A0=>nx15745, A1=>
      new_size_squared_out_3);
   ix13422 : mux21_ni port map ( Y=>nx13421, A0=>mem_data_in(3), A1=>
      new_size_squared_out_3, S0=>nx18325);
   ix15845 : xnor2 port map ( Y=>nx15844, A0=>nx15750, A1=>nx15848);
   ix13402 : mux21_ni port map ( Y=>nx13401, A0=>mem_data_in(2), A1=>
      new_size_squared_out_2, S0=>nx18327);
   ix15850 : xor2 port map ( Y=>nx15849, A0=>nx15756, A1=>
      new_size_squared_out_1);
   ix13382 : mux21_ni port map ( Y=>nx13381, A0=>mem_data_in(1), A1=>
      new_size_squared_out_1, S0=>nx18327);
   ix15855 : xor2 port map ( Y=>nx15854, A0=>nx15763, A1=>
      new_size_squared_out_0);
   ix13362 : mux21_ni port map ( Y=>nx13361, A0=>mem_data_in(0), A1=>
      new_size_squared_out_0, S0=>nx18327);
   ix577 : or02 port map ( Y=>nx576, A0=>ftc_cntrl_reg_out_11, A1=>nx15888);
   ix551 : and04 port map ( Y=>nx550, A0=>nx15873, A1=>nx15893, A2=>nx15902, 
      A3=>nx15907);
   ix13222 : mux21 port map ( Y=>nx13221, A0=>nx15890, A1=>nx15873, S0=>
      nx18283);
   ix15879 : or03 port map ( Y=>nx15878, A0=>ftc_cntrl_reg_out_8, A1=>
      nx15861, A2=>nx15883);
   ix1147 : ao21 port map ( Y=>nx1146, A0=>nx18279, A1=>nx15605, B0=>
      current_state_16);
   ix15891 : xor2 port map ( Y=>nx15890, A0=>nx15873, A1=>nx12885);
   ix531 : nor02ii port map ( Y=>nx12885, A0=>nx15898, A1=>
      window_width_cntr_counter_out_14);
   ix13212 : mux21_ni port map ( Y=>nx13211, A0=>nx524, A1=>
      window_width_cntr_counter_out_14, S0=>nx18283);
   ix525 : xor2 port map ( Y=>nx524, A0=>nx15893, A1=>nx15898);
   ix13202 : mux21 port map ( Y=>nx13201, A0=>nx15904, A1=>nx15902, S0=>
      nx18283);
   ix507 : nor02ii port map ( Y=>nx12887, A0=>nx15912, A1=>
      window_width_cntr_counter_out_12);
   ix13192 : mux21_ni port map ( Y=>nx13191, A0=>nx500, A1=>
      window_width_cntr_counter_out_12, S0=>nx18283);
   ix501 : xor2 port map ( Y=>nx500, A0=>nx15907, A1=>nx15912);
   ix13182 : mux21 port map ( Y=>nx13181, A0=>nx15918, A1=>nx15916, S0=>
      nx18283);
   ix483 : nor02ii port map ( Y=>nx12889, A0=>nx15926, A1=>
      window_width_cntr_counter_out_10);
   ix13172 : mux21_ni port map ( Y=>nx13171, A0=>nx476, A1=>
      window_width_cntr_counter_out_10, S0=>nx18283);
   ix477 : xor2 port map ( Y=>nx476, A0=>nx15921, A1=>nx15926);
   ix13162 : mux21 port map ( Y=>nx13161, A0=>nx15932, A1=>nx15930, S0=>
      nx18283);
   ix459 : nor02ii port map ( Y=>nx12891, A0=>nx15940, A1=>
      window_width_cntr_counter_out_8);
   ix13152 : mux21_ni port map ( Y=>nx13151, A0=>nx452, A1=>
      window_width_cntr_counter_out_8, S0=>nx18285);
   ix453 : xor2 port map ( Y=>nx452, A0=>nx15935, A1=>nx15940);
   ix13142 : mux21 port map ( Y=>nx13141, A0=>nx15946, A1=>nx15944, S0=>
      nx18285);
   ix435 : nor02ii port map ( Y=>nx12893, A0=>nx15954, A1=>
      window_width_cntr_counter_out_6);
   ix13132 : mux21_ni port map ( Y=>nx13131, A0=>nx428, A1=>
      window_width_cntr_counter_out_6, S0=>nx18285);
   ix429 : xor2 port map ( Y=>nx428, A0=>nx15949, A1=>nx15954);
   ix15955 : or03 port map ( Y=>nx15954, A0=>nx18167, A1=>nx15995, A2=>
      nx15959);
   ix18166 : inv01 port map ( Y=>nx18167, A=>wind_width_count_4);
   ix14042 : mux21_ni port map ( Y=>nx14041, A0=>nx1876, A1=>
      wind_width_count_4, S0=>nx18285);
   ix13092 : mux21_ni port map ( Y=>nx13091, A0=>nx384, A1=>
      wind_width_count_1, S0=>nx18285);
   ix13082 : xor2 port map ( Y=>nx13081, A0=>nx17811, A1=>nx12884);
   ix13102 : mux21_ni port map ( Y=>nx13101, A0=>nx392, A1=>
      wind_width_count_2, S0=>nx18285);
   ix13112 : mux21_ni port map ( Y=>nx13111, A0=>nx400, A1=>
      wind_width_count_3, S0=>nx18285);
   ix13122 : mux21 port map ( Y=>nx13121, A0=>nx15997, A1=>nx15995, S0=>
      nx18287);
   ix565 : and04 port map ( Y=>nx564, A0=>nx15916, A1=>nx15921, A2=>nx15930, 
      A3=>nx15935);
   ix613 : and04 port map ( Y=>nx612, A0=>nx15944, A1=>nx15949, A2=>nx15995, 
      A3=>nx18169);
   ix18168 : inv01 port map ( Y=>nx18169, A=>nx604);
   ix603 : mux21 port map ( Y=>nx602, A0=>nx18305, A1=>img_width_out_0, S0=>
      nx18225);
   ix13242 : ao221 port map ( Y=>nx13241, A0=>img_width_out_0, A1=>nx18259, 
      B0=>nx18911, B1=>new_width_out_0, C0=>nx17897);
   ix641 : mux21 port map ( Y=>nx640, A0=>nx18305, A1=>nx16189, S0=>nx18225
   );
   ix13262 : ao22 port map ( Y=>nx13261, A0=>img_width_out_1, A1=>nx18261, 
      B0=>nx18911, B1=>new_width_out_1);
   ix705 : nor02ii port map ( Y=>nx704, A0=>nx16042, A1=>nx18225);
   ix16043 : xor2 port map ( Y=>nx16042, A0=>nx16046, A1=>nx16037);
   ix13302 : ao22 port map ( Y=>nx13301, A0=>img_width_out_3, A1=>nx18261, 
      B0=>nx18911, B1=>new_width_out_3);
   ix723 : nor02ii port map ( Y=>nx722, A0=>nx16055, A1=>nx18227);
   ix16064 : and04 port map ( Y=>nx16063, A0=>nx16005, A1=>nx16019, A2=>
      nx18171, A3=>nx16046);
   ix18170 : inv01 port map ( Y=>nx18171, A=>img_width_out_2);
   ix16066 : or02 port map ( Y=>nx16065, A0=>nx15605, A1=>nx15621);
   ix16068 : xor2 port map ( Y=>nx16067, A0=>nx15614, A1=>nx12896);
   ix1383 : nor02ii port map ( Y=>nx12896, A0=>nx16075, A1=>
      cache_width_cntr_counter_out_14);
   ix13832 : mux21_ni port map ( Y=>nx13831, A0=>nx1376, A1=>
      cache_width_cntr_counter_out_14, S0=>nx18289);
   ix1377 : xor2 port map ( Y=>nx1376, A0=>nx16070, A1=>nx16075);
   ix13822 : mux21 port map ( Y=>nx13821, A0=>nx16081, A1=>nx16079, S0=>
      nx18289);
   ix1359 : nor02ii port map ( Y=>nx12898, A0=>nx16089, A1=>
      cache_width_cntr_counter_out_12);
   ix13812 : mux21_ni port map ( Y=>nx13811, A0=>nx1352, A1=>
      cache_width_cntr_counter_out_12, S0=>nx18289);
   ix1353 : xor2 port map ( Y=>nx1352, A0=>nx16084, A1=>nx16089);
   ix13802 : mux21 port map ( Y=>nx13801, A0=>nx16095, A1=>nx16093, S0=>
      nx18289);
   ix1335 : nor02ii port map ( Y=>nx12900, A0=>nx16103, A1=>
      cache_width_cntr_counter_out_10);
   ix13792 : mux21_ni port map ( Y=>nx13791, A0=>nx1328, A1=>
      cache_width_cntr_counter_out_10, S0=>nx18289);
   ix1329 : xor2 port map ( Y=>nx1328, A0=>nx16098, A1=>nx16103);
   ix13782 : mux21 port map ( Y=>nx13781, A0=>nx16109, A1=>nx16107, S0=>
      nx18289);
   ix1311 : nor02ii port map ( Y=>nx12902, A0=>nx16117, A1=>
      cache_width_cntr_counter_out_8);
   ix13772 : mux21_ni port map ( Y=>nx13771, A0=>nx1304, A1=>
      cache_width_cntr_counter_out_8, S0=>nx18291);
   ix1305 : xor2 port map ( Y=>nx1304, A0=>nx16112, A1=>nx16117);
   ix13762 : mux21 port map ( Y=>nx13761, A0=>nx16123, A1=>nx16121, S0=>
      nx18291);
   ix1287 : nor02ii port map ( Y=>nx12904, A0=>nx16131, A1=>
      cache_width_cntr_counter_out_6);
   ix13752 : mux21_ni port map ( Y=>nx13751, A0=>nx1280, A1=>
      cache_width_cntr_counter_out_6, S0=>nx18291);
   ix1281 : xor2 port map ( Y=>nx1280, A0=>nx16126, A1=>nx16131);
   ix16132 : or03 port map ( Y=>nx16131, A0=>nx18173, A1=>nx16178, A2=>
      nx16136);
   ix18172 : inv01 port map ( Y=>nx18173, A=>nx17817);
   ix13732 : mux21_ni port map ( Y=>nx13731, A0=>nx1254, A1=>nx17815, S0=>
      nx18291);
   ix13702 : mux21_ni port map ( Y=>nx13701, A0=>nx1230, A1=>
      cache_width_count_1, S0=>nx18291);
   ix13692 : xor2 port map ( Y=>nx13691, A0=>cache_width_count_0, A1=>
      nx18383);
   ix16151 : mux21_ni port map ( Y=>nx16150, A0=>cache_height_count_en, A1=>
      nx17871, S0=>nx18279);
   ix16154 : and02 port map ( Y=>nx16153, A0=>nx18279, A1=>nx15605);
   ix1213 : nor02ii port map ( Y=>nx1212, A0=>nx16155, A1=>
      ftc_cntrl_reg_out_10);
   ix13712 : mux21_ni port map ( Y=>nx13711, A0=>nx1238, A1=>nx17819, S0=>
      nx18291);
   ix13722 : mux21_ni port map ( Y=>nx13721, A0=>nx1246, A1=>
      cache_width_count_3, S0=>nx18291);
   ix13742 : mux21 port map ( Y=>nx13741, A0=>nx16180, A1=>nx16178, S0=>
      nx18293);
   ix1417 : and04 port map ( Y=>nx1416, A0=>nx16093, A1=>nx16098, A2=>
      nx16107, A3=>nx16112);
   ix1435 : and04 port map ( Y=>nx1434, A0=>nx16121, A1=>nx16126, A2=>
      nx16178, A3=>nx18175);
   ix1427 : xnor2 port map ( Y=>nx18175, A0=>nx16005, A1=>
      cache_width_count_0);
   ix1437 : xor2 port map ( Y=>nx1436, A0=>cache_width_count_1, A1=>nx636);
   ix16192 : and02 port map ( Y=>nx16191, A0=>nx16005, A1=>nx16019);
   ix1485 : nor02_2x port map ( Y=>nx1484, A0=>nx18273, A1=>nx18307);
   ix1867 : and02 port map ( Y=>nx12906, A0=>current_state_21, A1=>nx15865);
   ix16223 : and02 port map ( Y=>nx16222, A0=>nx18265, A1=>nx18333);
   ix16227 : nor02ii port map ( Y=>nx16226, A0=>num_channels_counter_out_1, 
      A1=>nx15531);
   ix1765 : mux21 port map ( Y=>nx1764, A0=>nx15508, A1=>nx16274, S0=>
      nx15445);
   ix16281 : mux21 port map ( Y=>nx16280, A0=>mem_data_in(0), A1=>nx16278, 
      S0=>nx15445);
   ix16283 : and02 port map ( Y=>nx16282, A0=>nx15445, A1=>nx18333);
   ix16285 : nor02ii port map ( Y=>nx16284, A0=>nlayers_counter_out_1, A1=>
      nx16278);
   ix1781 : mux21 port map ( Y=>nx1780, A0=>nx15518, A1=>nx16290, S0=>
      nx15445);
   ix309 : or02 port map ( Y=>nx308, A0=>nx18307, A1=>nx18257);
   ix16322 : nor02ii port map ( Y=>argmax_ready_EXMPLR, A0=>nx16327, A1=>
      nx1926);
   ix1927 : or04 port map ( Y=>nx1926, A0=>class_cntr_counter_out_0, A1=>
      nx16332, A2=>class_cntr_counter_out_2, A3=>nx18887);
   ix14052 : mux21 port map ( Y=>nx14051, A0=>current_state_27, A1=>nx18339, 
      S0=>nx16324);
   ix14062 : mux21 port map ( Y=>nx14061, A0=>nx16334, A1=>nx16332, S0=>
      nx18339);
   ix16337 : or02 port map ( Y=>nx16336, A0=>nx16332, A1=>nx16324);
   ix14072 : mux21_ni port map ( Y=>nx14071, A0=>nx1904, A1=>
      class_cntr_counter_out_2, S0=>nx18339);
   ix1905 : xor2 port map ( Y=>nx1904, A0=>nx16338, A1=>nx16336);
   ix14082 : mux21_ni port map ( Y=>nx14081, A0=>nx1912, A1=>
      class_cntr_counter_out_3, S0=>nx18341);
   ix1913 : xor2 port map ( Y=>nx1912, A0=>nx18887, A1=>nx16346);
   ix16347 : or03 port map ( Y=>nx16346, A0=>nx16338, A1=>nx16332, A2=>
      nx16324);
   ix4917 : nor02ii port map ( Y=>argmax_data_out(0), A0=>nx18341, A1=>
      mem_data_in(0));
   ix4919 : nor02ii port map ( Y=>argmax_data_out(1), A0=>nx18341, A1=>
      mem_data_in(1));
   ix4921 : nor02ii port map ( Y=>argmax_data_out(2), A0=>nx18341, A1=>
      mem_data_in(2));
   ix4923 : nor02ii port map ( Y=>argmax_data_out(3), A0=>nx18341, A1=>
      mem_data_in(3));
   ix4925 : nor02ii port map ( Y=>argmax_data_out(4), A0=>nx18341, A1=>
      mem_data_in(4));
   ix4927 : nor02ii port map ( Y=>argmax_data_out(5), A0=>nx18341, A1=>
      mem_data_in(5));
   ix4929 : nor02ii port map ( Y=>argmax_data_out(6), A0=>nx18343, A1=>
      mem_data_in(6));
   ix4931 : nor02ii port map ( Y=>argmax_data_out(7), A0=>nx18343, A1=>
      mem_data_in(7));
   ix4933 : nor02ii port map ( Y=>argmax_data_out(8), A0=>nx18343, A1=>
      mem_data_in(8));
   ix4935 : nor02ii port map ( Y=>argmax_data_out(9), A0=>nx18343, A1=>
      mem_data_in(9));
   ix4937 : nor02ii port map ( Y=>argmax_data_out(10), A0=>nx18343, A1=>
      mem_data_in(10));
   ix4939 : nor02ii port map ( Y=>argmax_data_out(11), A0=>nx18343, A1=>
      mem_data_in(11));
   ix4941 : nor02ii port map ( Y=>argmax_data_out(12), A0=>nx18343, A1=>
      mem_data_in(12));
   ix4943 : nor02ii port map ( Y=>argmax_data_out(13), A0=>nx18345, A1=>
      mem_data_in(13));
   ix4945 : nor02ii port map ( Y=>argmax_data_out(14), A0=>nx18345, A1=>
      mem_data_in(14));
   ix4947 : nor02ii port map ( Y=>argmax_data_out(15), A0=>nx18345, A1=>
      mem_data_in(15));
   ix4949 : and02 port map ( Y=>comp_unit_data2_out(0), A0=>nx18233, A1=>
      nx2140);
   ix2141 : mux21_ni port map ( Y=>nx2140, A0=>flt_bias_out_0, A1=>
      mem_data_in(0), S0=>nx18297);
   ix4951 : and02 port map ( Y=>comp_unit_data2_out(1), A0=>nx18233, A1=>
      nx2168);
   ix2169 : mux21_ni port map ( Y=>nx2168, A0=>flt_bias_out_1, A1=>
      mem_data_in(1), S0=>nx18297);
   ix4953 : and02 port map ( Y=>comp_unit_data2_out(2), A0=>nx18235, A1=>
      nx2194);
   ix2195 : mux21_ni port map ( Y=>nx2194, A0=>flt_bias_out_2, A1=>
      mem_data_in(2), S0=>nx18297);
   ix4955 : and02 port map ( Y=>comp_unit_data2_out(3), A0=>nx18235, A1=>
      nx2220);
   ix2221 : mux21_ni port map ( Y=>nx2220, A0=>flt_bias_out_3, A1=>
      mem_data_in(3), S0=>nx18297);
   ix4957 : and02 port map ( Y=>comp_unit_data2_out(4), A0=>nx18235, A1=>
      nx2246);
   ix2247 : mux21_ni port map ( Y=>nx2246, A0=>flt_bias_out_4, A1=>
      mem_data_in(4), S0=>nx18297);
   ix4959 : and02 port map ( Y=>comp_unit_data2_out(5), A0=>nx18235, A1=>
      nx2272);
   ix2273 : mux21_ni port map ( Y=>nx2272, A0=>flt_bias_out_5, A1=>
      mem_data_in(5), S0=>nx18299);
   ix4961 : and02 port map ( Y=>comp_unit_data2_out(6), A0=>nx18235, A1=>
      nx2298);
   ix2299 : mux21_ni port map ( Y=>nx2298, A0=>flt_bias_out_6, A1=>
      mem_data_in(6), S0=>nx18299);
   ix4963 : and02 port map ( Y=>comp_unit_data2_out(7), A0=>nx18235, A1=>
      nx2324);
   ix2325 : mux21_ni port map ( Y=>nx2324, A0=>flt_bias_out_7, A1=>
      mem_data_in(7), S0=>nx18299);
   ix4965 : and02 port map ( Y=>comp_unit_data2_out(8), A0=>nx18235, A1=>
      nx2350);
   ix2351 : mux21_ni port map ( Y=>nx2350, A0=>flt_bias_out_8, A1=>
      mem_data_in(8), S0=>nx18299);
   ix4967 : and02 port map ( Y=>comp_unit_data2_out(9), A0=>nx18237, A1=>
      nx2376);
   ix2377 : mux21_ni port map ( Y=>nx2376, A0=>flt_bias_out_9, A1=>
      mem_data_in(9), S0=>nx18299);
   ix4969 : and02 port map ( Y=>comp_unit_data2_out(10), A0=>nx18237, A1=>
      nx2402);
   ix2403 : mux21_ni port map ( Y=>nx2402, A0=>flt_bias_out_10, A1=>
      mem_data_in(10), S0=>nx18299);
   ix4971 : and02 port map ( Y=>comp_unit_data2_out(11), A0=>nx18237, A1=>
      nx2428);
   ix2429 : mux21_ni port map ( Y=>nx2428, A0=>flt_bias_out_11, A1=>
      mem_data_in(11), S0=>nx18299);
   ix4973 : and02 port map ( Y=>comp_unit_data2_out(12), A0=>nx18237, A1=>
      nx2454);
   ix2455 : mux21_ni port map ( Y=>nx2454, A0=>flt_bias_out_12, A1=>
      mem_data_in(12), S0=>nx18301);
   ix4975 : and02 port map ( Y=>comp_unit_data2_out(13), A0=>nx18237, A1=>
      nx2480);
   ix2481 : mux21_ni port map ( Y=>nx2480, A0=>flt_bias_out_13, A1=>
      mem_data_in(13), S0=>nx18301);
   ix4977 : and02 port map ( Y=>comp_unit_data2_out(14), A0=>nx18237, A1=>
      nx2506);
   ix2507 : mux21_ni port map ( Y=>nx2506, A0=>flt_bias_out_14, A1=>
      mem_data_in(14), S0=>nx18301);
   ix4979 : and02 port map ( Y=>comp_unit_data2_out(15), A0=>nx18237, A1=>
      nx2532);
   ix2533 : mux21_ni port map ( Y=>nx2532, A0=>flt_bias_out_15, A1=>
      mem_data_in(15), S0=>nx18301);
   ix5147 : and03 port map ( Y=>max_height_1, A0=>nx636, A1=>nx17803, A2=>
      nx18281);
   ix16456 : or03 port map ( Y=>nx16455, A0=>nx18307, A1=>nx15605, A2=>
      nx16463);
   ix16466 : ao21 port map ( Y=>nx2580, A0=>nx16463, A1=>nx12912, B0=>nx1182
   );
   ix2583 : and02 port map ( Y=>cache_data_in_0, A0=>mem_data_in(0), A1=>
      nx18243);
   ix2585 : and02 port map ( Y=>cache_data_in_1, A0=>mem_data_in(1), A1=>
      nx18243);
   ix2587 : and02 port map ( Y=>cache_data_in_2, A0=>mem_data_in(2), A1=>
      nx18243);
   ix2589 : and02 port map ( Y=>cache_data_in_3, A0=>mem_data_in(3), A1=>
      nx18245);
   ix2591 : and02 port map ( Y=>cache_data_in_4, A0=>mem_data_in(4), A1=>
      nx18245);
   ix2593 : and02 port map ( Y=>cache_data_in_5, A0=>mem_data_in(5), A1=>
      nx18245);
   ix2595 : and02 port map ( Y=>cache_data_in_6, A0=>mem_data_in(6), A1=>
      nx18245);
   ix2597 : and02 port map ( Y=>cache_data_in_7, A0=>mem_data_in(7), A1=>
      nx18245);
   ix2599 : and02 port map ( Y=>cache_data_in_8, A0=>mem_data_in(8), A1=>
      nx18245);
   ix2601 : and02 port map ( Y=>cache_data_in_9, A0=>mem_data_in(9), A1=>
      nx18245);
   ix2603 : and02 port map ( Y=>cache_data_in_10, A0=>mem_data_in(10), A1=>
      nx18247);
   ix2605 : and02 port map ( Y=>cache_data_in_11, A0=>mem_data_in(11), A1=>
      nx18247);
   ix2607 : and02 port map ( Y=>cache_data_in_12, A0=>mem_data_in(12), A1=>
      nx18247);
   ix2609 : and02 port map ( Y=>cache_data_in_13, A0=>mem_data_in(13), A1=>
      nx18247);
   ix2611 : and02 port map ( Y=>cache_data_in_14, A0=>mem_data_in(14), A1=>
      nx18247);
   ix2613 : and02 port map ( Y=>cache_data_in_15, A0=>mem_data_in(15), A1=>
      nx18247);
   ix16508 : and02 port map ( Y=>nx16507, A0=>nx17803, A1=>nx18281);
   ix14112 : mux21 port map ( Y=>nx14111, A0=>nx16514, A1=>nx16511, S0=>
      nx18273);
   ix14132 : mux21 port map ( Y=>nx14131, A0=>nx16521, A1=>nx16518, S0=>
      nx18273);
   ix14152 : mux21 port map ( Y=>nx14151, A0=>nx16527, A1=>nx16524, S0=>
      nx18273);
   ix14172 : mux21 port map ( Y=>nx14171, A0=>nx16533, A1=>nx16530, S0=>
      nx18273);
   ix14192 : mux21 port map ( Y=>nx14191, A0=>nx16539, A1=>nx16536, S0=>
      nx18275);
   ix14212 : mux21 port map ( Y=>nx14211, A0=>nx16545, A1=>nx16542, S0=>
      nx18275);
   ix14232 : mux21 port map ( Y=>nx14231, A0=>nx16551, A1=>nx16548, S0=>
      nx18275);
   ix14252 : mux21 port map ( Y=>nx14251, A0=>nx16557, A1=>nx16554, S0=>
      nx18275);
   ix14272 : mux21 port map ( Y=>nx14271, A0=>nx16563, A1=>nx16560, S0=>
      nx18275);
   ix14292 : mux21 port map ( Y=>nx14291, A0=>nx16569, A1=>nx16566, S0=>
      nx18275);
   ix14312 : mux21 port map ( Y=>nx14311, A0=>nx16575, A1=>nx16572, S0=>
      nx18275);
   ix14332 : mux21 port map ( Y=>nx14331, A0=>nx16581, A1=>nx16578, S0=>
      nx18277);
   ix14352 : mux21 port map ( Y=>nx14351, A0=>nx16587, A1=>nx16584, S0=>
      nx18277);
   ix14372 : mux21 port map ( Y=>nx14371, A0=>nx16593, A1=>nx16590, S0=>
      nx18277);
   ix14392 : mux21 port map ( Y=>nx14391, A0=>nx16599, A1=>nx16596, S0=>
      nx18277);
   ix14412 : mux21 port map ( Y=>nx14411, A0=>nx16605, A1=>nx16602, S0=>
      nx18277);
   ix4885 : nor02ii port map ( Y=>filter_data_out(0), A0=>nx18319, A1=>
      mem_data_in(0));
   ix4887 : nor02ii port map ( Y=>filter_data_out(1), A0=>nx18319, A1=>
      mem_data_in(1));
   ix4889 : nor02ii port map ( Y=>filter_data_out(2), A0=>nx18319, A1=>
      mem_data_in(2));
   ix4891 : nor02ii port map ( Y=>filter_data_out(3), A0=>nx18319, A1=>
      mem_data_in(3));
   ix4893 : nor02ii port map ( Y=>filter_data_out(4), A0=>nx18319, A1=>
      mem_data_in(4));
   ix4895 : nor02ii port map ( Y=>filter_data_out(5), A0=>nx18321, A1=>
      mem_data_in(5));
   ix4897 : nor02ii port map ( Y=>filter_data_out(6), A0=>nx18321, A1=>
      mem_data_in(6));
   ix4899 : nor02ii port map ( Y=>filter_data_out(7), A0=>nx18321, A1=>
      mem_data_in(7));
   ix4901 : nor02ii port map ( Y=>filter_data_out(8), A0=>nx18321, A1=>
      mem_data_in(8));
   ix4903 : nor02ii port map ( Y=>filter_data_out(9), A0=>nx18321, A1=>
      mem_data_in(9));
   ix4905 : nor02ii port map ( Y=>filter_data_out(10), A0=>nx18321, A1=>
      mem_data_in(10));
   ix4907 : nor02ii port map ( Y=>filter_data_out(11), A0=>nx18321, A1=>
      mem_data_in(11));
   ix4909 : nor02ii port map ( Y=>filter_data_out(12), A0=>nx17863, A1=>
      mem_data_in(12));
   ix4911 : nor02ii port map ( Y=>filter_data_out(13), A0=>nx17863, A1=>
      mem_data_in(13));
   ix4913 : nor02ii port map ( Y=>filter_data_out(14), A0=>nx17863, A1=>
      mem_data_in(14));
   ix4915 : nor02ii port map ( Y=>filter_data_out(15), A0=>nx17863, A1=>
      mem_data_in(15));
   ix4981 : and02 port map ( Y=>wind_col_in_0_0, A0=>nx18359, A1=>
      cache_data_out_0_0);
   ix4983 : and02 port map ( Y=>wind_col_in_0_1, A0=>nx18359, A1=>
      cache_data_out_0_1);
   ix4985 : and02 port map ( Y=>wind_col_in_0_2, A0=>nx18359, A1=>
      cache_data_out_0_2);
   ix4987 : and02 port map ( Y=>wind_col_in_0_3, A0=>nx18359, A1=>
      cache_data_out_0_3);
   ix4989 : and02 port map ( Y=>wind_col_in_0_4, A0=>nx18359, A1=>
      cache_data_out_0_4);
   ix4991 : and02 port map ( Y=>wind_col_in_0_5, A0=>nx18359, A1=>
      cache_data_out_0_5);
   ix4993 : and02 port map ( Y=>wind_col_in_0_6, A0=>nx18359, A1=>
      cache_data_out_0_6);
   ix4995 : and02 port map ( Y=>wind_col_in_0_7, A0=>nx18361, A1=>
      cache_data_out_0_7);
   ix4997 : and02 port map ( Y=>wind_col_in_0_8, A0=>nx18361, A1=>
      cache_data_out_0_8);
   ix4999 : and02 port map ( Y=>wind_col_in_0_9, A0=>nx18361, A1=>
      cache_data_out_0_9);
   ix5001 : and02 port map ( Y=>wind_col_in_0_10, A0=>nx18361, A1=>
      cache_data_out_0_10);
   ix5003 : and02 port map ( Y=>wind_col_in_0_11, A0=>nx18361, A1=>
      cache_data_out_0_11);
   ix5005 : and02 port map ( Y=>wind_col_in_0_12, A0=>nx18361, A1=>
      cache_data_out_0_12);
   ix5007 : and02 port map ( Y=>wind_col_in_0_13, A0=>nx18361, A1=>
      cache_data_out_0_13);
   ix5009 : and02 port map ( Y=>wind_col_in_0_14, A0=>nx18363, A1=>
      cache_data_out_0_14);
   ix5011 : and02 port map ( Y=>wind_col_in_0_15, A0=>nx18363, A1=>
      cache_data_out_0_15);
   ix5013 : and02 port map ( Y=>wind_col_in_1_0, A0=>nx18363, A1=>
      cache_data_out_1_0);
   ix5015 : and02 port map ( Y=>wind_col_in_1_1, A0=>nx18363, A1=>
      cache_data_out_1_1);
   ix5017 : and02 port map ( Y=>wind_col_in_1_2, A0=>nx18363, A1=>
      cache_data_out_1_2);
   ix5019 : and02 port map ( Y=>wind_col_in_1_3, A0=>nx18363, A1=>
      cache_data_out_1_3);
   ix5021 : and02 port map ( Y=>wind_col_in_1_4, A0=>nx18363, A1=>
      cache_data_out_1_4);
   ix5023 : and02 port map ( Y=>wind_col_in_1_5, A0=>nx18365, A1=>
      cache_data_out_1_5);
   ix5025 : and02 port map ( Y=>wind_col_in_1_6, A0=>nx18365, A1=>
      cache_data_out_1_6);
   ix5027 : and02 port map ( Y=>wind_col_in_1_7, A0=>nx18365, A1=>
      cache_data_out_1_7);
   ix5029 : and02 port map ( Y=>wind_col_in_1_8, A0=>nx18365, A1=>
      cache_data_out_1_8);
   ix5031 : and02 port map ( Y=>wind_col_in_1_9, A0=>nx18365, A1=>
      cache_data_out_1_9);
   ix5033 : and02 port map ( Y=>wind_col_in_1_10, A0=>nx18365, A1=>
      cache_data_out_1_10);
   ix5035 : and02 port map ( Y=>wind_col_in_1_11, A0=>nx18365, A1=>
      cache_data_out_1_11);
   ix5037 : and02 port map ( Y=>wind_col_in_1_12, A0=>nx18367, A1=>
      cache_data_out_1_12);
   ix5039 : and02 port map ( Y=>wind_col_in_1_13, A0=>nx18367, A1=>
      cache_data_out_1_13);
   ix5041 : and02 port map ( Y=>wind_col_in_1_14, A0=>nx18367, A1=>
      cache_data_out_1_14);
   ix5043 : and02 port map ( Y=>wind_col_in_1_15, A0=>nx18367, A1=>
      cache_data_out_1_15);
   ix5045 : and02 port map ( Y=>wind_col_in_2_0, A0=>nx18367, A1=>
      cache_data_out_2_0);
   ix5047 : and02 port map ( Y=>wind_col_in_2_1, A0=>nx18367, A1=>
      cache_data_out_2_1);
   ix5049 : and02 port map ( Y=>wind_col_in_2_2, A0=>nx18367, A1=>
      cache_data_out_2_2);
   ix5051 : and02 port map ( Y=>wind_col_in_2_3, A0=>nx18155, A1=>
      cache_data_out_2_3);
   ix5053 : and02 port map ( Y=>wind_col_in_2_4, A0=>nx18155, A1=>
      cache_data_out_2_4);
   ix5055 : and02 port map ( Y=>wind_col_in_2_5, A0=>nx18155, A1=>
      cache_data_out_2_5);
   ix5057 : and02 port map ( Y=>wind_col_in_2_6, A0=>nx18155, A1=>
      cache_data_out_2_6);
   ix5059 : and02 port map ( Y=>wind_col_in_2_7, A0=>nx18155, A1=>
      cache_data_out_2_7);
   ix5061 : and02 port map ( Y=>wind_col_in_2_8, A0=>nx18155, A1=>
      cache_data_out_2_8);
   ix5063 : and02 port map ( Y=>wind_col_in_2_9, A0=>nx18155, A1=>
      cache_data_out_2_9);
   ix5065 : and02 port map ( Y=>wind_col_in_2_10, A0=>nx18369, A1=>
      cache_data_out_2_10);
   ix5067 : and02 port map ( Y=>wind_col_in_2_11, A0=>nx18369, A1=>
      cache_data_out_2_11);
   ix5069 : and02 port map ( Y=>wind_col_in_2_12, A0=>nx18369, A1=>
      cache_data_out_2_12);
   ix5071 : and02 port map ( Y=>wind_col_in_2_13, A0=>nx18369, A1=>
      cache_data_out_2_13);
   ix5073 : and02 port map ( Y=>wind_col_in_2_14, A0=>nx18369, A1=>
      cache_data_out_2_14);
   ix5075 : and02 port map ( Y=>wind_col_in_2_15, A0=>nx18369, A1=>
      cache_data_out_2_15);
   ix5077 : and02 port map ( Y=>wind_col_in_3_0, A0=>nx18369, A1=>
      cache_data_out_3_0);
   ix5079 : and02 port map ( Y=>wind_col_in_3_1, A0=>nx18371, A1=>
      cache_data_out_3_1);
   ix5081 : and02 port map ( Y=>wind_col_in_3_2, A0=>nx18371, A1=>
      cache_data_out_3_2);
   ix5083 : and02 port map ( Y=>wind_col_in_3_3, A0=>nx18371, A1=>
      cache_data_out_3_3);
   ix5085 : and02 port map ( Y=>wind_col_in_3_4, A0=>nx18371, A1=>
      cache_data_out_3_4);
   ix5087 : and02 port map ( Y=>wind_col_in_3_5, A0=>nx18371, A1=>
      cache_data_out_3_5);
   ix5089 : and02 port map ( Y=>wind_col_in_3_6, A0=>nx18371, A1=>
      cache_data_out_3_6);
   ix5091 : and02 port map ( Y=>wind_col_in_3_7, A0=>nx18371, A1=>
      cache_data_out_3_7);
   ix5093 : and02 port map ( Y=>wind_col_in_3_8, A0=>nx18373, A1=>
      cache_data_out_3_8);
   ix5095 : and02 port map ( Y=>wind_col_in_3_9, A0=>nx18373, A1=>
      cache_data_out_3_9);
   ix5097 : and02 port map ( Y=>wind_col_in_3_10, A0=>nx18373, A1=>
      cache_data_out_3_10);
   ix5099 : and02 port map ( Y=>wind_col_in_3_11, A0=>nx18373, A1=>
      cache_data_out_3_11);
   ix5101 : and02 port map ( Y=>wind_col_in_3_12, A0=>nx18373, A1=>
      cache_data_out_3_12);
   ix5103 : and02 port map ( Y=>wind_col_in_3_13, A0=>nx18373, A1=>
      cache_data_out_3_13);
   ix5105 : and02 port map ( Y=>wind_col_in_3_14, A0=>nx18373, A1=>
      cache_data_out_3_14);
   ix5107 : and02 port map ( Y=>wind_col_in_3_15, A0=>nx18375, A1=>
      cache_data_out_3_15);
   ix5109 : and02 port map ( Y=>wind_col_in_4_0, A0=>nx18375, A1=>
      cache_data_out_4_0);
   ix5111 : and02 port map ( Y=>wind_col_in_4_1, A0=>nx18375, A1=>
      cache_data_out_4_1);
   ix5113 : and02 port map ( Y=>wind_col_in_4_2, A0=>nx18375, A1=>
      cache_data_out_4_2);
   ix5115 : and02 port map ( Y=>wind_col_in_4_3, A0=>nx18375, A1=>
      cache_data_out_4_3);
   ix5117 : and02 port map ( Y=>wind_col_in_4_4, A0=>nx18375, A1=>
      cache_data_out_4_4);
   ix5119 : and02 port map ( Y=>wind_col_in_4_5, A0=>nx18375, A1=>
      cache_data_out_4_5);
   ix5121 : and02 port map ( Y=>wind_col_in_4_6, A0=>nx18157, A1=>
      cache_data_out_4_6);
   ix5123 : and02 port map ( Y=>wind_col_in_4_7, A0=>nx18157, A1=>
      cache_data_out_4_7);
   ix5125 : and02 port map ( Y=>wind_col_in_4_8, A0=>nx18157, A1=>
      cache_data_out_4_8);
   ix5127 : and02 port map ( Y=>wind_col_in_4_9, A0=>nx18157, A1=>
      cache_data_out_4_9);
   ix5129 : and02 port map ( Y=>wind_col_in_4_10, A0=>nx18157, A1=>
      cache_data_out_4_10);
   ix5131 : and02 port map ( Y=>wind_col_in_4_11, A0=>nx18157, A1=>
      cache_data_out_4_11);
   ix5133 : and02 port map ( Y=>wind_col_in_4_12, A0=>nx18157, A1=>
      cache_data_out_4_12);
   ix5135 : and02 port map ( Y=>wind_col_in_4_13, A0=>nx2546, A1=>
      cache_data_out_4_13);
   ix5137 : and02 port map ( Y=>wind_col_in_4_14, A0=>nx2546, A1=>
      cache_data_out_4_14);
   ix5139 : and02 port map ( Y=>wind_col_in_4_15, A0=>nx2546, A1=>
      cache_data_out_4_15);
   ix2555 : or03 port map ( Y=>wind_en, A0=>nx15974, A1=>nx18385, A2=>
      nx12906);
   ix2547 : or03 port map ( Y=>nx2546, A0=>nx15865, A1=>nx15970, A2=>nx18307
   );
   ix16716 : and03 port map ( Y=>nx16715, A0=>nx18137, A1=>nx18345, A2=>
      nx18313);
   ix2641 : nand02 port map ( Y=>nx16927, A0=>nx18301, A1=>nx18239);
   ix16720 : nor02ii port map ( Y=>nx2142, A0=>nx18277, A1=>nx196);
   ix1947 : nor02_2x port map ( Y=>nx1946, A0=>nx1926, A1=>nx16327);
   ix16743 : nor02ii port map ( Y=>nx16742, A0=>new_size_squared_out_0, A1=>
      nx16745);
   ix16748 : or02 port map ( Y=>nx16747, A0=>nx16745, A1=>nx16324);
   ix14482 : xor2 port map ( Y=>nx14481, A0=>addr1_data_0, A1=>nx18347);
   ix16752 : or03 port map ( Y=>nx18119, A0=>nx2128, A1=>nx17927, A2=>nx2754
   );
   ix14472 : xor2 port map ( Y=>nx14471, A0=>img_addr_offset_0, A1=>nx18247
   );
   ix14462 : mux21_ni port map ( Y=>nx14461, A0=>nx16764, A1=>
      img_base_addr_0, S0=>nx18333);
   ix14452 : mux21 port map ( Y=>nx14451, A0=>nx16764, A1=>nx16745, S0=>
      nx18353);
   ix16771 : xor2 port map ( Y=>nx16770, A0=>nflt_layer_temp_1, A1=>nx15500
   );
   ix2675 : xor2 port map ( Y=>nx2674, A0=>nflt_layer_temp_0, A1=>
      nflt_layer_out_0);
   ix16775 : xor2 port map ( Y=>nx16774, A0=>nflt_layer_temp_2, A1=>nx15512
   );
   ix14442 : mux21_ni port map ( Y=>nx14441, A0=>nx15763, A1=>
      bias_offset_data_out_0, S0=>nx18313);
   ix16792 : or02 port map ( Y=>nx16791, A0=>nx16745, A1=>nx15763);
   ix16799 : xnor2 port map ( Y=>nx16798, A0=>nx16802, A1=>nx16332);
   ix14492 : ao32 port map ( Y=>nx14491, A0=>write_base_data_out_1, A1=>
      nx18265, A2=>nx18335, B0=>nx19308, B1=>nx18177);
   ix18176 : inv01 port map ( Y=>nx18177, A=>nx16804);
   ix14522 : mux21 port map ( Y=>nx14521, A0=>nx16820, A1=>nx16818, S0=>
      nx18335);
   ix14512 : mux21_ni port map ( Y=>nx14511, A0=>write_base_prev_data_out_1, 
      A1=>write_base_data_out_1, S0=>nx18353);
   ix16826 : nor02ii port map ( Y=>nx16825, A0=>write_base_prev_data_out_1, 
      A1=>nx16764);
   ix14532 : mux21 port map ( Y=>nx14531, A0=>nx16833, A1=>nx16829, S0=>
      nx18249);
   ix16840 : xnor2 port map ( Y=>nx16839, A0=>nx16843, A1=>nx16802);
   ix14542 : ao32 port map ( Y=>nx14541, A0=>nx18179, A1=>nx18301, A2=>
      nx18239, B0=>bias_offset_data_out_1, B1=>nx18313);
   ix18178 : inv01 port map ( Y=>nx18179, A=>nx15759);
   ix14502 : mux21 port map ( Y=>nx14501, A0=>nx16846, A1=>nx16849, S0=>
      nx18347);
   ix16864 : xnor2 port map ( Y=>nx16863, A0=>nx16802, A1=>nx15756);
   ix16875 : xnor2 port map ( Y=>nx16874, A0=>nx18885, A1=>nx16338);
   ix14552 : ao32 port map ( Y=>nx14551, A0=>write_base_data_out_2, A1=>
      nx18265, A2=>nx18335, B0=>nx19308, B1=>nx18181);
   ix18180 : inv01 port map ( Y=>nx18181, A=>nx16880);
   ix14602 : ao32 port map ( Y=>nx14601, A0=>nx18183, A1=>nx18301, A2=>
      nx18239, B0=>bias_offset_data_out_2, B1=>nx18313);
   ix18182 : inv01 port map ( Y=>nx18183, A=>nx15753);
   ix14582 : mux21_ni port map ( Y=>nx14581, A0=>nx2974, A1=>img_base_addr_2, 
      S0=>nx18335);
   ix14572 : mux21 port map ( Y=>nx14571, A0=>nx16906, A1=>nx18885, S0=>
      nx18353);
   ix14592 : mux21_ni port map ( Y=>nx14591, A0=>img_addr_offset_2, A1=>
      nx2988, S0=>nx18249);
   ix2989 : xor2 port map ( Y=>nx2988, A0=>nx16915, A1=>nx16831);
   ix14562 : mux21_ni port map ( Y=>nx14561, A0=>addr1_data_2, A1=>nx2942, 
      S0=>nx18347);
   ix16925 : xnor2 port map ( Y=>nx16924, A0=>nx18885, A1=>nx15750);
   ix2933 : oai21 port map ( Y=>nx2932, A0=>nx18185, A1=>nx18345, B0=>
      nx18311);
   ix18184 : inv01 port map ( Y=>nx18185, A=>nx2874);
   ix14612 : mux21_ni port map ( Y=>nx14611, A0=>write_base_data_out_3, A1=>
      nx3050, S0=>nx19308);
   ix16944 : xor2 port map ( Y=>nx16943, A0=>new_size_squared_out_3, A1=>
      nx18889);
   ix14652 : mux21_ni port map ( Y=>nx14651, A0=>nx3146, A1=>img_base_addr_3, 
      S0=>nx18335);
   ix14642 : mux21_ni port map ( Y=>nx14641, A0=>write_base_prev_data_out_3, 
      A1=>write_base_data_out_3, S0=>nx18353);
   ix14662 : mux21_ni port map ( Y=>nx14661, A0=>img_addr_offset_3, A1=>
      nx3160, S0=>nx18249);
   ix16968 : xor2 port map ( Y=>nx16967, A0=>bias_offset_data_out_3, A1=>
      nx18889);
   ix14632 : mux21_ni port map ( Y=>nx14631, A0=>nx832, A1=>
      bias_offset_data_out_3, S0=>nx18313);
   ix833 : xor2 port map ( Y=>nx832, A0=>nx15745, A1=>nx15768);
   ix14622 : mux21_ni port map ( Y=>nx14621, A0=>addr1_data_3, A1=>nx3092, 
      S0=>nx18347);
   ix14672 : ao32 port map ( Y=>nx14671, A0=>write_base_data_out_4, A1=>
      nx18267, A2=>nx18335, B0=>nx19308, B1=>nx18187);
   ix18186 : inv01 port map ( Y=>nx18187, A=>nx17004);
   ix14722 : mux21_ni port map ( Y=>nx14721, A0=>nx858, A1=>
      bias_offset_data_out_4, S0=>nx18313);
   ix14702 : mux21_ni port map ( Y=>nx14701, A0=>nx3270, A1=>img_base_addr_4, 
      S0=>nx18335);
   ix14692 : mux21 port map ( Y=>nx14691, A0=>nx17031, A1=>nx18891, S0=>
      nx18353);
   ix14712 : mux21_ni port map ( Y=>nx14711, A0=>img_addr_offset_4, A1=>
      nx3284, S0=>nx18249);
   ix3279 : nor02ii port map ( Y=>nx3278, A0=>nx17042, A1=>img_addr_offset_4
   );
   ix17052 : xnor2 port map ( Y=>nx17051, A0=>nx18891, A1=>nx15735);
   ix14682 : mux21_ni port map ( Y=>nx14681, A0=>addr1_data_4, A1=>nx3238, 
      S0=>nx18347);
   ix3233 : nor02ii port map ( Y=>nx3232, A0=>nx17060, A1=>addr1_data_4);
   ix14732 : mux21_ni port map ( Y=>nx14731, A0=>write_base_data_out_5, A1=>
      nx3346, S0=>nx19308);
   ix17075 : xor2 port map ( Y=>nx17074, A0=>new_size_squared_out_5, A1=>
      nx17076);
   ix17082 : xnor2 port map ( Y=>nx17081, A0=>nx17085, A1=>nx17076);
   ix14782 : ao32 port map ( Y=>nx14781, A0=>nx18189, A1=>nx18303, A2=>
      nx18239, B0=>bias_offset_data_out_5, B1=>nx18315);
   ix18188 : inv01 port map ( Y=>nx18189, A=>nx15732);
   ix17090 : xor2 port map ( Y=>nx17089, A0=>img_base_addr_5, A1=>nx17104);
   ix14762 : mux21_ni port map ( Y=>nx14761, A0=>nx3412, A1=>img_base_addr_5, 
      S0=>nx18041);
   ix14752 : mux21_ni port map ( Y=>nx14751, A0=>write_base_prev_data_out_5, 
      A1=>write_base_data_out_5, S0=>nx18353);
   ix14772 : mux21 port map ( Y=>nx14771, A0=>nx17104, A1=>nx17100, S0=>
      nx18249);
   ix14742 : mux21 port map ( Y=>nx14741, A0=>nx17114, A1=>nx17110, S0=>
      nx18347);
   ix14842 : mux21_ni port map ( Y=>nx14841, A0=>nx904, A1=>
      bias_offset_data_out_6, S0=>nx18315);
   ix14792 : ao32 port map ( Y=>nx14791, A0=>write_base_data_out_6, A1=>
      nx18267, A2=>nx18041, B0=>nx19308, B1=>nx18191);
   ix18190 : inv01 port map ( Y=>nx18191, A=>nx17140);
   ix14822 : mux21_ni port map ( Y=>nx14821, A0=>nx3554, A1=>img_base_addr_6, 
      S0=>nx18041);
   ix14812 : mux21 port map ( Y=>nx14811, A0=>nx17157, A1=>nx18893, S0=>
      nx18353);
   ix14832 : mux21_ni port map ( Y=>nx14831, A0=>img_addr_offset_6, A1=>
      nx3568, S0=>nx18249);
   ix3563 : nor02ii port map ( Y=>nx3562, A0=>nx17102, A1=>img_addr_offset_6
   );
   ix3361 : nor02ii port map ( Y=>nx3360, A0=>nx17077, A1=>
      write_base_data_out_5);
   ix17187 : xnor2 port map ( Y=>nx17186, A0=>nx18893, A1=>nx15720);
   ix14802 : mux21_ni port map ( Y=>nx14801, A0=>addr1_data_6, A1=>nx3522, 
      S0=>nx18347);
   ix3523 : xor2 port map ( Y=>nx3522, A0=>nx17188, A1=>nx17112);
   ix14852 : mux21_ni port map ( Y=>nx14851, A0=>nx18895, A1=>nx3630, S0=>
      nx19294);
   ix17205 : xor2_2x port map ( Y=>nx17204, A0=>new_size_squared_out_7, A1=>
      nx17199);
   ix17211 : xnor2 port map ( Y=>nx17210, A0=>nx17214, A1=>nx17199);
   ix14902 : ao32 port map ( Y=>nx14901, A0=>nx18193, A1=>nx18303, A2=>
      nx18239, B0=>bias_offset_data_out_7, B1=>nx18315);
   ix18192 : inv01 port map ( Y=>nx18193, A=>nx15717);
   ix17219 : xor2 port map ( Y=>nx17218, A0=>img_base_addr_7, A1=>nx17233);
   ix14882 : mux21_ni port map ( Y=>nx14881, A0=>nx3696, A1=>img_base_addr_7, 
      S0=>nx18041);
   ix14872 : mux21_ni port map ( Y=>nx14871, A0=>write_base_prev_data_out_7, 
      A1=>nx18895, S0=>nx18355);
   ix14892 : mux21 port map ( Y=>nx14891, A0=>nx17233, A1=>nx17229, S0=>
      nx18249);
   ix14862 : mux21 port map ( Y=>nx14861, A0=>nx17244, A1=>nx17239, S0=>
      nx18349);
   ix3517 : nor02ii port map ( Y=>nx3516, A0=>nx17112, A1=>addr1_data_6);
   ix3655 : oai21 port map ( Y=>nx3654, A0=>nx18195, A1=>nx18345, B0=>
      nx18311);
   ix18194 : inv01 port map ( Y=>nx18195, A=>nx3600);
   ix14962 : mux21_ni port map ( Y=>nx14961, A0=>nx954, A1=>
      bias_offset_data_out_8, S0=>nx18315);
   ix14912 : ao32 port map ( Y=>nx14911, A0=>nx18897, A1=>nx18267, A2=>
      nx18337, B0=>nx19294, B1=>nx18197);
   ix18196 : inv01 port map ( Y=>nx18197, A=>nx17270);
   ix14942 : mux21_ni port map ( Y=>nx14941, A0=>nx3838, A1=>img_base_addr_8, 
      S0=>nx18337);
   ix14932 : mux21 port map ( Y=>nx14931, A0=>nx17287, A1=>nx18899, S0=>
      nx18355);
   ix14952 : mux21_ni port map ( Y=>nx14951, A0=>img_addr_offset_8, A1=>
      nx3852, S0=>nx18251);
   ix3847 : nor02ii port map ( Y=>nx3846, A0=>nx17231, A1=>img_addr_offset_8
   );
   ix17311 : xnor2 port map ( Y=>nx17310, A0=>nx18899, A1=>nx15686);
   ix14922 : mux21_ni port map ( Y=>nx14921, A0=>addr1_data_8, A1=>nx3806, 
      S0=>nx18349);
   ix3807 : xor2 port map ( Y=>nx3806, A0=>nx17315, A1=>nx17242);
   ix14972 : mux21_ni port map ( Y=>nx14971, A0=>nx18901, A1=>nx3914, S0=>
      nx19294);
   ix17332 : xor2 port map ( Y=>nx17331, A0=>new_size_squared_out_9, A1=>
      nx17326);
   ix17338 : xnor2 port map ( Y=>nx17337, A0=>nx17341, A1=>nx17326);
   ix15022 : ao32 port map ( Y=>nx15021, A0=>nx18199, A1=>nx18303, A2=>
      nx18239, B0=>bias_offset_data_out_9, B1=>nx18315);
   ix18198 : inv01 port map ( Y=>nx18199, A=>nx15683);
   ix17346 : xor2 port map ( Y=>nx17345, A0=>img_base_addr_9, A1=>nx17360);
   ix15002 : mux21_ni port map ( Y=>nx15001, A0=>nx3980, A1=>img_base_addr_9, 
      S0=>nx18337);
   ix14992 : mux21_ni port map ( Y=>nx14991, A0=>write_base_prev_data_out_9, 
      A1=>nx18901, S0=>nx18355);
   ix15012 : mux21 port map ( Y=>nx15011, A0=>nx17360, A1=>nx17356, S0=>
      nx18251);
   ix14982 : mux21 port map ( Y=>nx14981, A0=>nx17371, A1=>nx17366, S0=>
      nx18349);
   ix3801 : nor02ii port map ( Y=>nx3800, A0=>nx17242, A1=>addr1_data_8);
   ix17378 : xnor2 port map ( Y=>nx17377, A0=>nx17326, A1=>nx15770);
   ix3939 : oai21 port map ( Y=>nx3938, A0=>nx18201, A1=>nx18345, B0=>
      nx18311);
   ix18200 : inv01 port map ( Y=>nx18201, A=>nx3884);
   ix15082 : mux21_ni port map ( Y=>nx15081, A0=>nx1000, A1=>
      bias_offset_data_out_10, S0=>nx18315);
   ix15032 : ao32 port map ( Y=>nx15031, A0=>write_base_data_out_10, A1=>
      nx18267, A2=>nx18337, B0=>nx19294, B1=>nx18203);
   ix18202 : inv01 port map ( Y=>nx18203, A=>nx17397);
   ix15062 : mux21_ni port map ( Y=>nx15061, A0=>nx4122, A1=>
      img_base_addr_10, S0=>nx18337);
   ix15052 : mux21 port map ( Y=>nx15051, A0=>nx17414, A1=>nx18903, S0=>
      nx18355);
   ix15072 : mux21_ni port map ( Y=>nx15071, A0=>img_addr_offset_10, A1=>
      nx4136, S0=>nx18251);
   ix4131 : nor02ii port map ( Y=>nx4130, A0=>nx17358, A1=>
      img_addr_offset_10);
   ix17438 : xnor2 port map ( Y=>nx17437, A0=>nx18903, A1=>nx15673);
   ix15042 : mux21_ni port map ( Y=>nx15041, A0=>addr1_data_10, A1=>nx4090, 
      S0=>nx18349);
   ix4091 : xor2 port map ( Y=>nx4090, A0=>nx17442, A1=>nx17369);
   ix15092 : mux21_ni port map ( Y=>nx15091, A0=>nx18905, A1=>nx4198, S0=>
      nx19294);
   ix17459 : xor2 port map ( Y=>nx17458, A0=>new_size_squared_out_11, A1=>
      nx18907);
   ix17465 : xnor2 port map ( Y=>nx17464, A0=>nx17468, A1=>nx18907);
   ix15142 : ao32 port map ( Y=>nx15141, A0=>nx18205, A1=>nx18303, A2=>
      nx18239, B0=>bias_offset_data_out_11, B1=>nx18315);
   ix18204 : inv01 port map ( Y=>nx18205, A=>nx15670);
   ix17473 : xor2 port map ( Y=>nx17472, A0=>img_base_addr_11, A1=>nx17487);
   ix15122 : mux21_ni port map ( Y=>nx15121, A0=>nx4264, A1=>
      img_base_addr_11, S0=>nx18337);
   ix15112 : mux21_ni port map ( Y=>nx15111, A0=>write_base_prev_data_out_11, 
      A1=>nx18905, S0=>nx18355);
   ix15132 : mux21 port map ( Y=>nx15131, A0=>nx17487, A1=>nx17483, S0=>
      nx18251);
   ix15102 : mux21 port map ( Y=>nx15101, A0=>nx17498, A1=>nx17493, S0=>
      nx18349);
   ix4085 : nor02ii port map ( Y=>nx4084, A0=>nx17369, A1=>addr1_data_10);
   ix4223 : oai21 port map ( Y=>nx4222, A0=>nx18207, A1=>nx18077, B0=>
      nx18311);
   ix18206 : inv01 port map ( Y=>nx18207, A=>nx4168);
   ix15202 : mux21_ni port map ( Y=>nx15201, A0=>nx1048, A1=>
      bias_offset_data_out_12, S0=>nx18317);
   ix15182 : mux21_ni port map ( Y=>nx15181, A0=>nx4406, A1=>
      img_base_addr_12, S0=>nx18043);
   ix15172 : mux21 port map ( Y=>nx15171, A0=>nx17541, A1=>nx18909, S0=>
      nx18355);
   ix15192 : mux21_ni port map ( Y=>nx15191, A0=>img_addr_offset_12, A1=>
      nx4420, S0=>nx18251);
   ix4415 : nor02ii port map ( Y=>nx4414, A0=>nx17485, A1=>
      img_addr_offset_12);
   ix17565 : xnor2 port map ( Y=>nx17564, A0=>nx18909, A1=>nx15660);
   ix15162 : mux21_ni port map ( Y=>nx15161, A0=>addr1_data_12, A1=>nx4374, 
      S0=>nx18349);
   ix4375 : xor2 port map ( Y=>nx4374, A0=>nx17566, A1=>nx17496);
   ix17592 : xnor2 port map ( Y=>nx17591, A0=>nx17595, A1=>nx18913);
   ix15262 : ao32 port map ( Y=>nx15261, A0=>nx18211, A1=>nx18303, A2=>
      nx18241, B0=>bias_offset_data_out_13, B1=>nx18317);
   ix18210 : inv01 port map ( Y=>nx18211, A=>nx15657);
   ix17600 : xor2 port map ( Y=>nx17599, A0=>img_base_addr_13, A1=>nx17614);
   ix15242 : mux21_ni port map ( Y=>nx15241, A0=>nx4548, A1=>
      img_base_addr_13, S0=>nx18043);
   ix15232 : mux21_ni port map ( Y=>nx15231, A0=>write_base_prev_data_out_13, 
      A1=>write_base_data_out_13, S0=>nx18355);
   ix15252 : mux21 port map ( Y=>nx15251, A0=>nx17614, A1=>nx17610, S0=>
      nx18251);
   ix15222 : mux21 port map ( Y=>nx15221, A0=>nx17625, A1=>nx17620, S0=>
      nx18349);
   ix4369 : nor02ii port map ( Y=>nx4368, A0=>nx17496, A1=>addr1_data_12);
   ix4507 : oai21 port map ( Y=>nx4506, A0=>nx18213, A1=>nx18077, B0=>
      nx18311);
   ix17642 : xnor2 port map ( Y=>nx17641, A0=>nx17646, A1=>nx18915);
   ix15322 : mux21_ni port map ( Y=>nx15321, A0=>nx1094, A1=>
      bias_offset_data_out_14, S0=>nx18317);
   ix1095 : xor2 port map ( Y=>nx1094, A0=>nx15647, A1=>nx15653);
   ix17664 : xnor2 port map ( Y=>nx17663, A0=>nx17673, A1=>nx17677);
   ix15302 : mux21_ni port map ( Y=>nx15301, A0=>nx4690, A1=>
      img_base_addr_14, S0=>nx18043);
   ix4691 : xnor2 port map ( Y=>nx4690, A0=>nx17670, A1=>nx17671);
   ix15292 : mux21 port map ( Y=>nx15291, A0=>nx17670, A1=>nx18915, S0=>
      nx18357);
   ix15312 : mux21_ni port map ( Y=>nx15311, A0=>img_addr_offset_14, A1=>
      nx4704, S0=>nx18251);
   ix4705 : xor2 port map ( Y=>nx4704, A0=>nx17677, A1=>nx17612);
   ix17680 : xor2 port map ( Y=>nx17679, A0=>nx18915, A1=>nx4496);
   ix17686 : xnor2 port map ( Y=>nx17685, A0=>nx18916, A1=>nx15647);
   ix15282 : mux21_ni port map ( Y=>nx15281, A0=>addr1_data_14, A1=>nx4658, 
      S0=>nx18351);
   ix4659 : xor2 port map ( Y=>nx4658, A0=>nx17687, A1=>nx17623);
   ix17712 : xor2 port map ( Y=>nx17711, A0=>img_base_addr_15, A1=>nx17726);
   ix15372 : mux21_ni port map ( Y=>nx15371, A0=>nx4834, A1=>
      img_base_addr_15, S0=>nx18043);
   ix15362 : mux21_ni port map ( Y=>nx15361, A0=>write_base_prev_data_out_15, 
      A1=>write_base_data_out_15, S0=>nx18357);
   ix15382 : mux21 port map ( Y=>nx15381, A0=>nx17726, A1=>nx17723, S0=>
      nx18253);
   ix17724 : xor2 port map ( Y=>nx17723, A0=>nx17726, A1=>nx4698);
   ix4699 : nor02ii port map ( Y=>nx4698, A0=>nx17612, A1=>
      img_addr_offset_14);
   ix4803 : xor2 port map ( Y=>nx4802, A0=>write_base_data_out_15, A1=>
      write_offset_data_out_15);
   ix15352 : mux21 port map ( Y=>nx15351, A0=>nx17740, A1=>nx17737, S0=>
      nx18351);
   ix17738 : xor2 port map ( Y=>nx17737, A0=>nx17740, A1=>nx4652);
   ix4653 : nor02ii port map ( Y=>nx4652, A0=>nx17623, A1=>addr1_data_14);
   ix17745 : xor2 port map ( Y=>nx17744, A0=>nx17748, A1=>
      write_base_data_out_15);
   ix15332 : ao32 port map ( Y=>nx15331, A0=>nx18217, A1=>nx18303, A2=>
      nx18241, B0=>bias_offset_data_out_15, B1=>nx18317);
   ix18216 : inv01 port map ( Y=>nx18217, A=>nx15644);
   ix18218 : inv02 port map ( Y=>nx18219, A=>nx16222);
   ix18224 : inv02 port map ( Y=>nx18225, A=>nx15974);
   ix18226 : inv02 port map ( Y=>nx18227, A=>nx15974);
   ix18228 : inv01 port map ( Y=>nx18229, A=>nx18049);
   ix18230 : inv01 port map ( Y=>nx18231, A=>nx18049);
   ix18232 : inv01 port map ( Y=>nx18233, A=>nx18059);
   ix18234 : inv01 port map ( Y=>nx18235, A=>nx18059);
   ix18236 : inv01 port map ( Y=>nx18237, A=>nx18059);
   ix18238 : inv02 port map ( Y=>nx18239, A=>nx18117);
   ix18240 : inv02 port map ( Y=>nx18241, A=>nx18117);
   ix18242 : inv02 port map ( Y=>nx18243, A=>nx18081);
   ix18244 : inv02 port map ( Y=>nx18245, A=>nx18081);
   ix18246 : inv02 port map ( Y=>nx18247, A=>nx18081);
   ix18248 : inv02 port map ( Y=>nx18249, A=>nx18081);
   ix18250 : inv02 port map ( Y=>nx18251, A=>nx18081);
   ix18252 : inv02 port map ( Y=>nx18253, A=>nx18081);
   ix18254 : inv02 port map ( Y=>nx18255, A=>nx17927);
   ix18256 : inv02 port map ( Y=>nx18257, A=>nx17927);
   ix18258 : inv02 port map ( Y=>nx18259, A=>nx582);
   ix18260 : inv02 port map ( Y=>nx18261, A=>nx582);
   ix18262 : buf02 port map ( Y=>nx18263, A=>nx15496);
   ix18264 : inv02 port map ( Y=>nx18265, A=>nx17887);
   ix18268 : inv01 port map ( Y=>nx18269, A=>nx148);
   ix18270 : inv01 port map ( Y=>nx18271, A=>nx148);
   ix18272 : inv02 port map ( Y=>nx18273, A=>nx17971);
   ix18274 : inv02 port map ( Y=>nx18275, A=>nx17971);
   ix18276 : inv02 port map ( Y=>nx18277, A=>nx17971);
   ix18278 : inv02 port map ( Y=>nx18279, A=>nx17921);
   ix18280 : inv02 port map ( Y=>nx18281, A=>nx17921);
   ix18282 : inv02 port map ( Y=>nx18283, A=>nx12884);
   ix18284 : inv02 port map ( Y=>nx18285, A=>nx12884);
   ix18286 : inv02 port map ( Y=>nx18287, A=>nx12884);
   ix18288 : inv02 port map ( Y=>nx18289, A=>nx1212);
   ix18290 : inv02 port map ( Y=>nx18291, A=>nx18383);
   ix18292 : inv02 port map ( Y=>nx18293, A=>nx18383);
   ix18294 : inv01 port map ( Y=>nx18295, A=>nx16373);
   ix18296 : inv02 port map ( Y=>nx18297, A=>nx18295);
   ix18298 : inv02 port map ( Y=>nx18299, A=>nx18295);
   ix18300 : inv02 port map ( Y=>nx18301, A=>nx18295);
   ix18302 : inv02 port map ( Y=>nx18303, A=>nx18295);
   ix18304 : inv02 port map ( Y=>nx18305, A=>comp_unit_flt_size_EXMPLR);
   ix18306 : inv02 port map ( Y=>nx18307, A=>comp_unit_flt_size_EXMPLR);
   ix18308 : inv02 port map ( Y=>nx18309, A=>nx17975);
   ix18310 : inv02 port map ( Y=>nx18311, A=>nx17975);
   ix18312 : inv02 port map ( Y=>nx18313, A=>nx18011);
   ix18314 : inv02 port map ( Y=>nx18315, A=>nx18011);
   ix18316 : inv02 port map ( Y=>nx18317, A=>nx18011);
   ix18318 : inv01 port map ( Y=>nx18319, A=>filter_ready_out_EXMPLR);
   ix18320 : inv01 port map ( Y=>nx18321, A=>filter_ready_out_EXMPLR);
   ix18322 : inv02 port map ( Y=>nx18323, A=>current_state_7);
   ix18324 : inv02 port map ( Y=>nx18325, A=>current_state_7);
   ix18326 : inv02 port map ( Y=>nx18327, A=>current_state_7);
   ix18328 : inv02 port map ( Y=>nx18329, A=>nx17947);
   ix18330 : inv02 port map ( Y=>nx18331, A=>nx17947);
   ix18332 : inv02 port map ( Y=>nx18333, A=>nx18912);
   ix18334 : inv02 port map ( Y=>nx18335, A=>nx18912);
   ix18338 : inv02 port map ( Y=>nx18339, A=>nx18381);
   ix18340 : inv02 port map ( Y=>nx18341, A=>nx18381);
   ix18342 : inv02 port map ( Y=>nx18343, A=>nx18381);
   ix18344 : inv02 port map ( Y=>nx18345, A=>nx18381);
   ix18346 : inv02 port map ( Y=>nx18347, A=>nx18121);
   ix18348 : inv02 port map ( Y=>nx18349, A=>nx18121);
   ix18350 : inv02 port map ( Y=>nx18351, A=>nx18121);
   ix18352 : inv02 port map ( Y=>nx18353, A=>nx16768);
   ix18354 : inv02 port map ( Y=>nx18355, A=>nx16768);
   ix18356 : inv02 port map ( Y=>nx18357, A=>nx16768);
   ix18358 : inv01 port map ( Y=>nx18359, A=>nx18385);
   ix18360 : inv01 port map ( Y=>nx18361, A=>nx18385);
   ix18362 : inv01 port map ( Y=>nx18363, A=>nx18385);
   ix18364 : inv01 port map ( Y=>nx18365, A=>nx18385);
   ix18366 : inv01 port map ( Y=>nx18367, A=>nx16629);
   ix18368 : inv01 port map ( Y=>nx18369, A=>nx16629);
   ix18370 : inv01 port map ( Y=>nx18371, A=>nx16629);
   ix18372 : inv01 port map ( Y=>nx18373, A=>nx16629);
   ix18374 : inv01 port map ( Y=>nx18375, A=>nx16629);
   ix18380 : inv02 port map ( Y=>nx18381, A=>nx18075);
   ix18382 : inv01 port map ( Y=>nx18383, A=>nx18289);
   ix18384 : inv01 port map ( Y=>nx18385, A=>nx2546);
   ix17068 : nor02ii port map ( Y=>nx17067, A0=>nx3366, A1=>nx16995);
   ix3367 : xor2 port map ( Y=>nx3366, A0=>nx17076, A1=>nx17077);
   ix16996 : nor02ii port map ( Y=>nx16995, A0=>nx3078, A1=>nx18867);
   ix18917 : buf04 port map ( Y=>nx18543, A=>nx17067);
   ix18918 : inv02 port map ( Y=>nx18544, A=>new_size_squared_out_15);
   ix18919 : inv02 port map ( Y=>nx18545, A=>write_base_data_out_15);
   ix18920 : oai32 port map ( Y=>nx18546, A0=>nx19302, A1=>nx18544, A2=>
      write_base_data_out_15, B0=>nx18545, B1=>new_size_squared_out_15);
   ix18921 : and02 port map ( Y=>nx18547, A0=>nx18909, A1=>nx15795);
   ix18922 : nor02_2x port map ( Y=>nx18548, A0=>nx18909, A1=>nx15795);
   ix18923 : and02 port map ( Y=>nx18549, A0=>nx18916, A1=>nx15785);
   ix18924 : inv02 port map ( Y=>nx18550, A=>write_base_data_out_13);
   ix18925 : inv02 port map ( Y=>nx18551, A=>new_size_squared_out_13);
   ix18926 : aoi32 port map ( Y=>nx18552, A0=>nx18223, A1=>nx18545, A2=>
      nx18544, B0=>write_base_data_out_15, B1=>new_size_squared_out_15);
   ix18927 : nor02_2x port map ( Y=>nx18553, A0=>NOT_nx4768, A1=>nx18552);
   reg_nx15341 : ao221 port map ( Y=>nx15341, A0=>nx18546, A1=>NOT_nx4768, 
      B0=>write_base_data_out_15, B1=>nx19302, C0=>nx18553);
   ix18928 : and02 port map ( Y=>nx18554, A0=>write_base_data_out_13, A1=>
      new_size_squared_out_13);
   ix18929 : inv02 port map ( Y=>nx18555, A=>nx17585);
   ix18930 : inv01 port map ( Y=>nx18556, A=>nx18916);
   ix18931 : inv02 port map ( Y=>nx18557, A=>nx15785);
   ix18932 : inv02 port map ( Y=>nx18558, A=>nx18909);
   ix18933 : inv02 port map ( Y=>nx18559, A=>nx15795);
   ix18934 : inv01 port map ( Y=>nx18560, A=>nx18885);
   ix18935 : inv02 port map ( Y=>nx18561, A=>nx15848);
   ix18936 : nand02_2x port map ( Y=>nx18562, A0=>nx18886, A1=>nx15848);
   reg_nx18009 : inv02 port map ( Y=>nx18009, A=>nx16745);
   ix18937 : inv02 port map ( Y=>nx18563, A=>nx16802);
   ix18938 : nand03_2x port map ( Y=>nx18564, A0=>new_size_squared_out_0, A1
      =>nx18009, A2=>nx18563);
   ix18939 : inv02 port map ( Y=>nx18565, A=>new_size_squared_out_1);
   ix18940 : nand02_2x port map ( Y=>nx18566, A0=>new_size_squared_out_1, A1
      =>nx18563);
   ix18941 : nand03_2x port map ( Y=>nx18567, A0=>nx18566, A1=>
      new_size_squared_out_0, A2=>nx18009);
   ix18942 : inv02 port map ( Y=>nx18568, A=>write_base_data_out_1);
   reg_nx3046 : inv01 port map ( Y=>nx3046, A=>nx18877);
   reg_nx16882 : inv01 port map ( Y=>nx16882, A=>nx18774);
   reg_nx16885 : oai22 port map ( Y=>nx16885, A0=>nx18560, A1=>nx18561, B0=>
      nx18886, B1=>nx15848);
   reg_nx16808 : oai22 port map ( Y=>nx16808, A0=>nx18563, A1=>
      new_size_squared_out_1, B0=>nx18565, B1=>nx16802);
   ix18943 : nor02_2x port map ( Y=>nx18569, A0=>nx18549, A1=>nx17585);
   ix18944 : nor02_2x port map ( Y=>nx18570, A0=>nx18547, A1=>nx17458);
   ix18945 : inv02 port map ( Y=>nx18571, A=>nx18905);
   ix18946 : inv02 port map ( Y=>nx18572, A=>new_size_squared_out_11);
   ix18947 : nor03_2x port map ( Y=>nx18573, A0=>nx18547, A1=>nx18571, A2=>
      nx18572);
   ix18948 : or02 port map ( Y=>nx18574, A0=>nx18573, A1=>nx18548);
   ix18949 : oai32 port map ( Y=>nx18575, A0=>nx18549, A1=>nx18550, A2=>
      nx18551, B0=>nx18916, B1=>nx15785);
   reg_NOT_nx4768 : aoi321 port map ( Y=>NOT_nx4768, A0=>nx18689, A1=>
      nx18569, A2=>nx18570, B0=>nx18574, B1=>nx18569, C0=>nx18575);
   ix18950 : inv01 port map ( Y=>nx18576, A=>nx18547);
   ix18951 : and02 port map ( Y=>nx18577, A0=>nx18905, A1=>
      new_size_squared_out_11);
   ix18952 : inv02 port map ( Y=>nx18578, A=>nx17458);
   ix18953 : inv02 port map ( Y=>nx18579, A=>nx16839);
   reg_nx16888 : aoi32 port map ( Y=>nx16888, A0=>nx18579, A1=>
      bias_offset_data_out_0, A2=>nx18009, B0=>write_base_data_out_1, B1=>
      bias_offset_data_out_1);
   ix18954 : and02 port map ( Y=>nx18580, A0=>nx18886, A1=>nx16895);
   ix18955 : nor02_2x port map ( Y=>nx18581, A0=>nx16888, A1=>nx18580);
   ix18956 : nor02_2x port map ( Y=>nx18582, A0=>nx18886, A1=>nx16895);
   ix18957 : and02 port map ( Y=>nx18583, A0=>nx18891, A1=>nx17021);
   ix18958 : inv02 port map ( Y=>nx18584, A=>write_base_data_out_3);
   ix18959 : inv02 port map ( Y=>nx18585, A=>bias_offset_data_out_3);
   reg_nx3444 : inv01 port map ( Y=>nx3444, A=>nx18657);
   ix18960 : and02 port map ( Y=>nx18586, A0=>write_base_data_out_3, A1=>
      bias_offset_data_out_3);
   ix18961 : inv02 port map ( Y=>nx18587, A=>nx16967);
   reg_nx17013 : oai32 port map ( Y=>nx17013, A0=>nx18586, A1=>nx18581, A2=>
      nx18582, B0=>nx18587, B1=>nx18586);
   ix18962 : nor02_2x port map ( Y=>nx18588, A0=>nx18891, A1=>nx17021);
   reg_nx17016 : ao21 port map ( Y=>nx17016, A0=>nx18891, A1=>nx17021, B0=>
      nx18588);
   reg_nx3112 : inv02 port map ( Y=>nx3112, A=>nx18660);
   reg_nx16891 : ao21 port map ( Y=>nx16891, A0=>nx18886, A1=>nx16895, B0=>
      nx18582);
   ix18963 : nand02_2x port map ( Y=>nx18589, A0=>write_offset_data_out_6, 
      A1=>write_base_data_out_6);
   ix18964 : inv02 port map ( Y=>nx18590, A=>nx16924);
   reg_nx16987 : aoi22 port map ( Y=>nx16987, A0=>write_offset_data_out_2, 
      A1=>write_base_data_out_2, B0=>nx2892, B1=>nx18590);
   ix18965 : and02 port map ( Y=>nx18591, A0=>nx15745, A1=>nx18889);
   ix18966 : nor02_2x port map ( Y=>nx18592, A0=>nx16987, A1=>nx18591);
   ix18967 : nor02_2x port map ( Y=>nx18593, A0=>nx15745, A1=>nx18889);
   ix18968 : and02 port map ( Y=>nx18594, A0=>nx15730, A1=>nx17076);
   ix18969 : inv02 port map ( Y=>nx18595, A=>write_offset_data_out_4);
   ix18970 : inv02 port map ( Y=>nx18596, A=>write_base_data_out_4);
   ix18971 : inv01 port map ( Y=>nx18597, A=>NOT_nx3476);
   ix18972 : and02 port map ( Y=>nx18598, A0=>write_offset_data_out_4, A1=>
      write_base_data_out_4);
   ix18973 : inv02 port map ( Y=>nx18599, A=>nx17051);
   reg_nx17118 : oai32 port map ( Y=>nx17118, A0=>nx18598, A1=>nx18592, A2=>
      nx18593, B0=>nx18599, B1=>nx18598);
   ix18974 : inv02 port map ( Y=>nx18600, A=>nx15730);
   ix18975 : inv02 port map ( Y=>nx18601, A=>nx17076);
   reg_nx17121 : oai22 port map ( Y=>nx17121, A0=>nx18600, A1=>nx18601, B0=>
      nx15730, B1=>nx17076);
   reg_nx3184 : inv01 port map ( Y=>nx3184, A=>nx18743);
   ix18976 : inv02 port map ( Y=>nx18602, A=>nx15745);
   ix18977 : inv02 port map ( Y=>nx18603, A=>nx18889);
   reg_nx16990 : oai22 port map ( Y=>nx16990, A0=>nx18602, A1=>nx18603, B0=>
      nx15745, B1=>nx18890);
   ix18978 : aoi22 port map ( Y=>nx18604, A0=>nx18576, A1=>nx18577, B0=>
      nx18690, B1=>nx18570);
   reg_nx17656 : oai22 port map ( Y=>nx17656, A0=>nx18556, A1=>nx18557, B0=>
      nx18916, B1=>nx15785);
   ix18979 : inv02 port map ( Y=>nx18605, A=>nx17656);
   reg_nx18223 : inv01 port map ( Y=>nx18223, A=>nx19302);
   ix18980 : nand02_2x port map ( Y=>nx18606, A0=>nx18223, A1=>nx18555);
   ix18981 : inv01 port map ( Y=>nx18607, A=>nx18604);
   ix18982 : inv02 port map ( Y=>nx18608, A=>nx18554);
   ix18983 : inv02 port map ( Y=>nx18609, A=>nx18548);
   ix18984 : nand04_2x port map ( Y=>nx18610, A0=>nx18605, A1=>nx18223, A2=>
      nx18608, A3=>nx18609);
   reg_nx18043 : inv02 port map ( Y=>nx18043, A=>nx18912);
   ix18985 : aoi21 port map ( Y=>nx18611, A0=>nx18548, A1=>nx18555, B0=>
      nx18554);
   ix18986 : inv02 port map ( Y=>nx18612, A=>nx18555);
   ix18987 : nand03_2x port map ( Y=>nx18613, A0=>nx18605, A1=>nx18608, A2=>
      nx18612);
   ix18988 : oai21 port map ( Y=>nx18614, A0=>nx18605, A1=>nx18611, B0=>
      nx18613);
   ix18989 : aoi32 port map ( Y=>nx18615, A0=>write_base_data_out_14, A1=>
      nx18267, A2=>nx18043, B0=>nx18223, B1=>nx18614);
   reg_nx15271 : oai321 port map ( Y=>nx15271, A0=>nx18604, A1=>nx18605, A2
      =>nx18606, B0=>nx18607, B1=>nx18610, C0=>nx18615);
   ix18990 : nand02_2x port map ( Y=>nx18616, A0=>write_offset_data_out_14, 
      A1=>write_base_data_out_14);
   ix18991 : inv02 port map ( Y=>nx18617, A=>nx15772);
   ix18992 : inv02 port map ( Y=>nx18618, A=>nx18907);
   ix18993 : nand02_2x port map ( Y=>nx18619, A0=>nx15772, A1=>nx18907);
   ix18994 : and02 port map ( Y=>nx18620, A0=>write_offset_data_out_10, A1=>
      write_base_data_out_10);
   ix18995 : aoi21 port map ( Y=>nx18621, A0=>nx15772, A1=>nx18908, B0=>
      nx17437);
   ix18996 : aoi222 port map ( Y=>nx18622, A0=>nx18617, A1=>nx18618, B0=>
      nx18619, B1=>nx18620, C0=>nx4044, C1=>nx18621);
   ix18997 : and02 port map ( Y=>nx18623, A0=>nx15774, A1=>nx18913);
   ix18998 : inv02 port map ( Y=>nx18624, A=>write_offset_data_out_12);
   ix18999 : inv02 port map ( Y=>nx18625, A=>write_base_data_out_12);
   reg_nx4612 : oai332 port map ( Y=>nx4612, A0=>nx18622, A1=>nx18623, A2=>
      nx17564, B0=>nx18623, B1=>nx18624, B2=>nx18625, C0=>nx15774, C1=>
      nx18913);
   ix19000 : inv02 port map ( Y=>nx18626, A=>nx4612);
   reg_nx17731 : ao22 port map ( Y=>nx17731, A0=>nx18616, A1=>nx18626, B0=>
      nx17685, B1=>nx18616);
   ix19001 : inv01 port map ( Y=>nx18627, A=>nx18626);
   ix19002 : oai21 port map ( Y=>nx18628, A0=>nx18624, A1=>nx18625, B0=>
      nx17564);
   ix19003 : oai21 port map ( Y=>nx18629, A0=>nx18624, A1=>nx18625, B0=>
      nx18622);
   reg_nx17629 : nand02_2x port map ( Y=>nx17629, A0=>nx18628, A1=>nx18629);
   ix19004 : inv02 port map ( Y=>nx18630, A=>nx15774);
   ix19005 : inv01 port map ( Y=>nx18631, A=>nx18913);
   reg_nx17632 : oai22 port map ( Y=>nx17632, A0=>nx18630, A1=>nx18631, B0=>
      nx15774, B1=>nx18913);
   reg_nx4328 : inv01 port map ( Y=>nx4328, A=>nx18622);
   ix19006 : inv02 port map ( Y=>nx18632, A=>nx17437);
   reg_nx17502 : oai22 port map ( Y=>nx17502, A0=>nx18620, A1=>nx4044, B0=>
      nx18632, B1=>nx18620);
   reg_nx17505 : oai22 port map ( Y=>nx17505, A0=>nx18617, A1=>nx18618, B0=>
      nx15772, B1=>nx18908);
   reg_nx17529 : oai22 port map ( Y=>nx17529, A0=>nx18558, A1=>nx18559, B0=>
      nx18910, B1=>nx15795);
   ix19007 : inv02 port map ( Y=>nx18633, A=>nx17529);
   ix19008 : inv02 port map ( Y=>nx18634, A=>write_base_data_out_12);
   ix19009 : or02 port map ( Y=>nx18635, A0=>nx17887, A1=>nx18912);
   ix19010 : nand03_2x port map ( Y=>nx18636, A0=>nx17526, A1=>nx19294, A2=>
      nx18633);
   reg_nx15151 : oai321 port map ( Y=>nx15151, A0=>nx18679, A1=>nx19302, A2
      =>nx18633, B0=>nx18634, B1=>nx18635, C0=>nx18636);
   reg_nx18267 : inv02 port map ( Y=>nx18267, A=>nx17887);
   reg_nx18337 : inv02 port map ( Y=>nx18337, A=>nx18912);
   ix19011 : nand02_2x port map ( Y=>nx18637, A0=>img_addr_offset_3, A1=>
      img_base_addr_3);
   ix19012 : nand02_2x port map ( Y=>nx18638, A0=>nx16915, A1=>nx16911);
   ix19013 : inv02 port map ( Y=>nx18639, A=>nx16818);
   ix19014 : inv02 port map ( Y=>nx18640, A=>nx16833);
   ix19015 : aoi22 port map ( Y=>nx18641, A0=>nx16818, A1=>nx16833, B0=>
      nx18639, B1=>nx18640);
   ix19016 : and02 port map ( Y=>nx18642, A0=>img_base_addr_0, A1=>
      img_addr_offset_0);
   ix19017 : inv02 port map ( Y=>nx18643, A=>nx16915);
   ix19018 : inv02 port map ( Y=>nx18644, A=>nx16911);
   ix19019 : aoi332 port map ( Y=>nx18645, A0=>nx18638, A1=>
      img_addr_offset_1, A2=>img_base_addr_1, B0=>nx18641, B1=>nx18638, B2=>
      nx18642, C0=>nx18643, C1=>nx18644);
   ix19020 : aoi22 port map ( Y=>nx18646, A0=>nx18637, A1=>nx18645, B0=>
      nx16948, B1=>nx18637);
   reg_nx17023 : inv01 port map ( Y=>nx17023, A=>nx18646);
   ix19021 : inv01 port map ( Y=>nx18647, A=>nx18646);
   reg_nx3132 : inv02 port map ( Y=>nx3132, A=>nx18645);
   ix19022 : and02 port map ( Y=>nx18648, A0=>img_addr_offset_1, A1=>
      img_base_addr_1);
   reg_nx16898 : oai22 port map ( Y=>nx16898, A0=>nx18641, A1=>nx18648, B0=>
      nx18648, B1=>nx18642);
   ix19023 : nor02_2x port map ( Y=>nx18649, A0=>nx16915, A1=>nx16911);
   reg_nx16901 : ao21 port map ( Y=>nx16901, A0=>nx16915, A1=>nx16911, B0=>
      nx18649);
   reg_nx16814 : oai22 port map ( Y=>nx16814, A0=>nx18639, A1=>nx18640, B0=>
      nx16818, B1=>nx16833);
   ix19024 : nand02_2x port map ( Y=>nx18650, A0=>write_base_data_out_5, A1
      =>bias_offset_data_out_5);
   ix19025 : inv01 port map ( Y=>nx18651, A=>nx18583);
   ix19026 : inv02 port map ( Y=>nx18652, A=>nx16967);
   ix19027 : inv01 port map ( Y=>nx18653, A=>nx18891);
   ix19028 : inv02 port map ( Y=>nx18654, A=>nx17021);
   ix19029 : inv02 port map ( Y=>nx18655, A=>nx18582);
   ix19030 : oai22 port map ( Y=>nx18656, A0=>nx18655, A1=>nx16967, B0=>
      nx18584, B1=>nx18585);
   ix19031 : aoi322 port map ( Y=>nx18657, A0=>nx18651, A1=>nx18581, A2=>
      nx18652, B0=>nx18653, B1=>nx18654, C0=>nx18656, C1=>nx18651);
   ix19032 : aoi22 port map ( Y=>nx18658, A0=>nx17081, A1=>nx18650, B0=>
      nx18650, B1=>nx18657);
   reg_nx17127 : inv02 port map ( Y=>nx17127, A=>nx18658);
   ix19033 : inv02 port map ( Y=>nx18659, A=>nx18658);
   ix19034 : nor02_2x port map ( Y=>nx18660, A0=>nx18581, A1=>nx18582);
   ix19035 : nand02_2x port map ( Y=>nx18661, A0=>nx18903, A1=>nx15806);
   ix19036 : inv01 port map ( Y=>nx18662, A=>nx18547);
   ix19037 : and02 port map ( Y=>nx18663, A0=>nx18578, A1=>nx18662);
   ix19038 : nor02_2x port map ( Y=>nx18664, A0=>nx18903, A1=>nx15806);
   ix19039 : inv02 port map ( Y=>nx18665, A=>nx18577);
   ix19040 : oai22 port map ( Y=>nx18666, A0=>nx18910, A1=>nx15795, B0=>
      nx18665, B1=>nx18547);
   ix19041 : aoi321 port map ( Y=>nx18667, A0=>nx18692, A1=>nx18661, A2=>
      nx18663, B0=>nx18663, B1=>nx18664, C0=>nx18666);
   ix19042 : inv02 port map ( Y=>nx18668, A=>new_size_squared_out_13);
   ix19043 : inv01 port map ( Y=>nx18669, A=>nx18913);
   ix19044 : aoi22 port map ( Y=>nx18670, A0=>nx18914, A1=>nx18668, B0=>
      new_size_squared_out_13, B1=>nx18669);
   ix19045 : inv02 port map ( Y=>nx18671, A=>write_base_data_out_13);
   ix19046 : oai22 port map ( Y=>nx18672, A0=>nx18668, A1=>nx18669, B0=>
      new_size_squared_out_13, B1=>nx18914);
   ix19047 : nand03_2x port map ( Y=>nx18673, A0=>nx18667, A1=>nx19294, A2=>
      nx18672);
   reg_nx15211 : oai321 port map ( Y=>nx15211, A0=>nx18667, A1=>nx19302, A2
      =>nx18670, B0=>nx18671, B1=>nx19296, C0=>nx18673);
   reg_nx17585 : oai22 port map ( Y=>nx17585, A0=>nx18669, A1=>
      new_size_squared_out_13, B0=>nx18668, B1=>nx18914);
   ix19048 : inv01 port map ( Y=>nx18674, A=>nx18903);
   ix19049 : inv02 port map ( Y=>nx18675, A=>nx15806);
   ix19050 : oai21 port map ( Y=>nx18676, A0=>nx18674, A1=>nx18675, B0=>
      nx18578);
   ix19051 : nor02_2x port map ( Y=>nx18677, A0=>nx18664, A1=>nx18577);
   ix19052 : aoi22 port map ( Y=>nx18678, A0=>nx18676, A1=>nx18665, B0=>
      nx18693, B1=>nx18677);
   reg_nx17526 : inv02 port map ( Y=>nx17526, A=>nx18678);
   ix19053 : inv02 port map ( Y=>nx18679, A=>nx18678);
   ix19054 : and02 port map ( Y=>nx18680, A0=>nx18903, A1=>nx15806);
   reg_nx17402 : ao21 port map ( Y=>nx17402, A0=>nx18904, A1=>nx15806, B0=>
      nx18664);
   ix19055 : and02 port map ( Y=>nx18681, A0=>nx18893, A1=>nx15827);
   ix19056 : nor02_2x port map ( Y=>nx18682, A0=>nx18681, A1=>nx18881);
   ix19057 : nor02_2x port map ( Y=>nx18683, A0=>nx18893, A1=>nx15827);
   ix19058 : and02 port map ( Y=>nx18684, A0=>nx18899, A1=>nx15816);
   ix19059 : inv02 port map ( Y=>nx18685, A=>nx18895);
   ix19060 : inv02 port map ( Y=>nx18686, A=>new_size_squared_out_7);
   ix19061 : inv02 port map ( Y=>nx18687, A=>nx18901);
   ix19062 : inv02 port map ( Y=>nx18688, A=>new_size_squared_out_9);
   reg_nx4194 : inv01 port map ( Y=>nx4194, A=>nx18805);
   ix19063 : inv01 port map ( Y=>nx18689, A=>nx18805);
   ix19064 : inv01 port map ( Y=>nx18690, A=>nx18805);
   ix19065 : nand02_2x port map ( Y=>nx18691, A0=>nx18901, A1=>
      new_size_squared_out_9);
   ix19066 : aoi22 port map ( Y=>nx18692, A0=>nx18691, A1=>NOT_nx3910, B0=>
      nx17331, B1=>nx18691);
   reg_nx17399 : inv02 port map ( Y=>nx17399, A=>nx18692);
   ix19067 : inv02 port map ( Y=>nx18693, A=>nx18692);
   ix19068 : inv01 port map ( Y=>nx18694, A=>NOT_nx3910);
   ix19069 : and02 port map ( Y=>nx18695, A0=>nx18895, A1=>
      new_size_squared_out_7);
   ix19070 : inv02 port map ( Y=>nx18696, A=>nx17204);
   reg_nx17272 : oai32 port map ( Y=>nx17272, A0=>nx18695, A1=>nx18682, A2=>
      nx18683, B0=>nx18696, B1=>nx18695);
   ix19071 : inv02 port map ( Y=>nx18697, A=>nx18899);
   ix19072 : inv02 port map ( Y=>nx18698, A=>nx15816);
   reg_nx17275 : oai22 port map ( Y=>nx17275, A0=>nx18697, A1=>nx18698, B0=>
      nx18899, B1=>nx15816);
   reg_nx3626 : oai22 port map ( Y=>nx3626, A0=>nx18893, A1=>nx15827, B0=>
      nx18681, B1=>nx18882);
   ix19073 : inv02 port map ( Y=>nx18699, A=>nx18894);
   ix19074 : inv02 port map ( Y=>nx18700, A=>nx15827);
   reg_nx17145 : oai22 port map ( Y=>nx17145, A0=>nx18699, A1=>nx18700, B0=>
      nx18894, B1=>nx15827);
   ix19075 : inv02 port map ( Y=>nx18701, A=>nx18905);
   ix19076 : inv02 port map ( Y=>nx18702, A=>write_base_data_out_12);
   ix19077 : inv02 port map ( Y=>nx18703, A=>write_base_data_out_13);
   ix19078 : inv02 port map ( Y=>nx18704, A=>nx3928);
   ix19079 : inv01 port map ( Y=>nx18705, A=>nx18914);
   ix19080 : inv02 port map ( Y=>nx18706, A=>nx18908);
   ix19081 : nor04_2x port map ( Y=>nx18707, A0=>write_base_data_out_12, A1
      =>write_base_data_out_10, A2=>nx18705, A3=>nx18706);
   ix19082 : and03 port map ( Y=>nx18708, A0=>nx17431, A1=>nx18704, A2=>
      nx18707);
   ix19083 : oai21 port map ( Y=>nx18709, A0=>nx4496, A1=>nx18708, B0=>
      nx17323);
   ix19084 : and02 port map ( Y=>nx18710, A0=>write_base_data_out_12, A1=>
      nx18906);
   ix19085 : inv01 port map ( Y=>nx18711, A=>nx17431);
   reg_nx4502 : oai422 port map ( Y=>nx4502, A0=>nx17431, A1=>nx18701, A2=>
      nx18702, A3=>write_base_data_out_13, B0=>nx18710, B1=>nx18914, C0=>
      nx18711, C1=>nx18914);
   ix19086 : nor02_2x port map ( Y=>nx18712, A0=>nx18701, A1=>nx17431);
   ix19087 : oai32 port map ( Y=>nx18713, A0=>nx18717, A1=>nx18701, A2=>
      write_base_data_out_12, B0=>nx18702, B1=>nx18712);
   ix19088 : inv02 port map ( Y=>nx18714, A=>write_base_data_out_10);
   ix19089 : nand04_2x port map ( Y=>nx18715, A0=>nx18717, A1=>nx18704, A2=>
      nx18908, A3=>nx18714);
   ix19090 : oai21 port map ( Y=>nx18716, A0=>nx18701, A1=>nx18717, B0=>
      nx18715);
   reg_nx17556 : oai322 port map ( Y=>nx17556, A0=>nx18717, A1=>nx18702, A2
      =>nx18701, B0=>nx18906, B1=>write_base_data_out_12, C0=>nx18711, C1=>
      write_base_data_out_12);
   reg_nx4218 : oai22 port map ( Y=>nx4218, A0=>nx18717, A1=>nx18906, B0=>
      nx18711, B1=>nx18908);
   reg_nx17429 : oai21 port map ( Y=>nx17429, A0=>nx3928, A1=>
      write_base_data_out_10, B0=>nx18717);
   reg_nx4168 : nand02_2x port map ( Y=>nx4168, A0=>nx17429, A1=>nx17323);
   ix19091 : buf02 port map ( Y=>nx18717, A=>nx17431);
   ix19092 : nand02_2x port map ( Y=>nx18718, A0=>write_base_data_out_13, A1
      =>bias_offset_data_out_13);
   ix19093 : nand02_2x port map ( Y=>nx18719, A0=>nx18904, A1=>nx17392);
   ix19094 : aoi21 port map ( Y=>nx18720, A0=>nx18904, A1=>nx17392, B0=>
      nx17337);
   ix19095 : nor02_2x port map ( Y=>nx18721, A0=>nx18904, A1=>nx17392);
   ix19096 : and02 port map ( Y=>nx18722, A0=>nx18910, A1=>nx17519);
   ix19097 : inv02 port map ( Y=>nx18723, A=>nx18906);
   ix19098 : inv02 port map ( Y=>nx18724, A=>bias_offset_data_out_11);
   reg_nx17638 : inv02 port map ( Y=>nx17638, A=>nx18851);
   ix19099 : inv02 port map ( Y=>nx18725, A=>nx18851);
   ix19100 : inv02 port map ( Y=>nx18726, A=>nx18850);
   ix19101 : nand02_2x port map ( Y=>nx18727, A0=>nx18906, A1=>
      bias_offset_data_out_11);
   ix19102 : inv02 port map ( Y=>nx18728, A=>nx17464);
   ix19103 : and02 port map ( Y=>nx18729, A0=>nx18906, A1=>
      bias_offset_data_out_11);
   ix19104 : nor02_2x port map ( Y=>nx18730, A0=>nx18728, A1=>nx18729);
   reg_nx17511 : ao21 port map ( Y=>nx17511, A0=>nx18727, A1=>nx18875, B0=>
      nx18730);
   ix19105 : nor02_2x port map ( Y=>nx18731, A0=>nx18910, A1=>nx17519);
   reg_nx17514 : ao21 port map ( Y=>nx17514, A0=>nx18910, A1=>nx17519, B0=>
      nx18731);
   reg_nx4296 : inv02 port map ( Y=>nx4296, A=>nx18875);
   ix19106 : and02 port map ( Y=>nx18732, A0=>nx18901, A1=>
      bias_offset_data_out_9);
   ix19107 : inv02 port map ( Y=>nx18733, A=>nx17337);
   reg_nx17384 : oai22 port map ( Y=>nx17384, A0=>nx18732, A1=>nx18857, B0=>
      nx18733, B1=>nx18732);
   reg_nx17387 : ao21 port map ( Y=>nx17387, A0=>nx18904, A1=>nx17392, B0=>
      nx18721);
   ix19108 : nor02_2x port map ( Y=>nx18734, A0=>nx17186, A1=>nx18594);
   ix19109 : inv02 port map ( Y=>nx18735, A=>nx17051);
   ix19110 : inv02 port map ( Y=>nx18736, A=>nx18593);
   ix19111 : oai22 port map ( Y=>nx18737, A0=>nx18736, A1=>nx17051, B0=>
      nx18595, B1=>nx18596);
   ix19112 : or02 port map ( Y=>nx18738, A0=>nx15730, A1=>nx17076);
   ix19113 : oai21 port map ( Y=>nx18739, A0=>nx17186, A1=>nx18738, B0=>
      nx18589);
   ix19114 : inv01 port map ( Y=>nx18740, A=>nx18594);
   ix19115 : inv02 port map ( Y=>nx18741, A=>nx15730);
   ix19116 : inv02 port map ( Y=>nx18742, A=>nx17076);
   reg_NOT_nx3476 : aoi322 port map ( Y=>NOT_nx3476, A0=>nx18740, A1=>
      nx18592, A2=>nx18735, B0=>nx18741, B1=>nx18742, C0=>nx18737, C1=>
      nx18740);
   ix19117 : nor02_2x port map ( Y=>nx18743, A0=>nx18593, A1=>nx18592);
   ix19118 : and02 port map ( Y=>nx18744, A0=>nx17044, A1=>nx17038);
   ix19119 : nor02_2x port map ( Y=>nx18745, A0=>nx18744, A1=>nx18647);
   ix19120 : nor02_2x port map ( Y=>nx18746, A0=>nx17044, A1=>nx17038);
   ix19121 : nor02_2x port map ( Y=>nx18747, A0=>nx18745, A1=>nx18746);
   ix19122 : and02 port map ( Y=>nx18748, A0=>nx17168, A1=>nx17164);
   ix19123 : inv02 port map ( Y=>nx18749, A=>img_addr_offset_5);
   ix19124 : inv02 port map ( Y=>nx18750, A=>img_base_addr_5);
   reg_nx3682 : oai332 port map ( Y=>nx3682, A0=>nx18747, A1=>nx18748, A2=>
      nx17089, B0=>nx18748, B1=>nx18749, B2=>nx18750, C0=>nx17168, C1=>
      nx17164);
   ix19125 : inv01 port map ( Y=>nx18751, A=>nx3682);
   ix19126 : and02 port map ( Y=>nx18752, A0=>nx17298, A1=>nx17294);
   ix19127 : inv02 port map ( Y=>nx18753, A=>img_addr_offset_7);
   ix19128 : inv02 port map ( Y=>nx18754, A=>img_base_addr_7);
   ix19129 : oai332 port map ( Y=>nx18755, A0=>nx18751, A1=>nx18752, A2=>
      nx17218, B0=>nx18752, B1=>nx18753, B2=>nx18754, C0=>nx17298, C1=>
      nx17294);
   ix19130 : inv02 port map ( Y=>nx18756, A=>nx18755);
   reg_nx3966 : inv02 port map ( Y=>nx3966, A=>nx18756);
   ix19131 : oai21 port map ( Y=>nx18757, A0=>nx18753, A1=>nx18754, B0=>
      nx17218);
   ix19132 : oai21 port map ( Y=>nx18758, A0=>nx18753, A1=>nx18754, B0=>
      nx18751);
   reg_nx17279 : nand02_2x port map ( Y=>nx17279, A0=>nx18757, A1=>nx18758);
   ix19133 : nor02_2x port map ( Y=>nx18759, A0=>nx17298, A1=>nx17294);
   reg_nx17282 : ao21 port map ( Y=>nx17282, A0=>nx17298, A1=>nx17294, B0=>
      nx18759);
   ix19134 : inv02 port map ( Y=>nx18760, A=>nx18751);
   ix19135 : and02 port map ( Y=>nx18761, A0=>img_addr_offset_5, A1=>
      img_base_addr_5);
   ix19136 : inv02 port map ( Y=>nx18762, A=>nx17089);
   reg_nx17149 : oai32 port map ( Y=>nx17149, A0=>nx18761, A1=>nx18745, A2=>
      nx18746, B0=>nx18762, B1=>nx18761);
   ix19137 : nor02_2x port map ( Y=>nx18763, A0=>nx17168, A1=>nx17164);
   reg_nx17152 : ao21 port map ( Y=>nx17152, A0=>nx17168, A1=>nx17164, B0=>
      nx18763);
   reg_nx3398 : oai22 port map ( Y=>nx3398, A0=>nx17044, A1=>nx17038, B0=>
      nx18744, B1=>nx18647);
   reg_nx17026 : ao21 port map ( Y=>nx17026, A0=>nx17044, A1=>nx17038, B0=>
      nx18746);
   ix19138 : nand02_2x port map ( Y=>nx18764, A0=>nx18567, A1=>nx18568);
   ix19139 : nand02_2x port map ( Y=>nx18765, A0=>nx18564, A1=>nx18565);
   ix19140 : inv02 port map ( Y=>nx18766, A=>nx3048);
   ix19141 : and02 port map ( Y=>nx18767, A0=>nx18891, A1=>nx15837);
   ix19142 : inv02 port map ( Y=>nx18768, A=>write_base_data_out_3);
   ix19143 : inv02 port map ( Y=>nx18769, A=>new_size_squared_out_3);
   reg_nx3342 : inv01 port map ( Y=>nx3342, A=>nx18879);
   ix19144 : ao21 port map ( Y=>nx18770, A0=>write_base_data_out_3, A1=>
      new_size_squared_out_3, B0=>nx3048);
   ix19145 : oai21 port map ( Y=>nx18771, A0=>nx18768, A1=>nx18769, B0=>
      nx18877);
   reg_nx17006 : nand02_2x port map ( Y=>nx17006, A0=>nx18770, A1=>nx18771);
   ix19146 : inv01 port map ( Y=>nx18772, A=>nx18891);
   ix19147 : inv02 port map ( Y=>nx18773, A=>nx15837);
   reg_nx17009 : oai22 port map ( Y=>nx17009, A0=>nx18772, A1=>nx18773, B0=>
      nx18892, B1=>nx15837);
   ix19148 : aoi22 port map ( Y=>nx18774, A0=>nx18564, A1=>nx18565, B0=>
      nx18567, B1=>nx18568);
   ix19149 : inv02 port map ( Y=>nx18775, A=>nx18902);
   ix19150 : inv02 port map ( Y=>nx18776, A=>write_base_data_out_10);
   ix19151 : inv02 port map ( Y=>nx18777, A=>nx18897);
   ix19152 : nor04_2x port map ( Y=>nx18778, A0=>nx18775, A1=>nx18703, A2=>
      nx18776, A3=>nx18777);
   ix19153 : inv01 port map ( Y=>nx18779, A=>nx18701);
   ix19154 : inv02 port map ( Y=>nx18780, A=>nx18702);
   reg_nx4496 : and04 port map ( Y=>nx4496, A0=>nx3644, A1=>nx18778, A2=>
      nx18779, A3=>nx18780);
   ix19155 : and02 port map ( Y=>nx18781, A0=>write_base_data_out_10, A1=>
      nx18897);
   reg_nx17431 : nand03_2x port map ( Y=>nx17431, A0=>nx3644, A1=>nx18902, 
      A2=>nx18781);
   ix19156 : inv02 port map ( Y=>nx18782, A=>nx17067);
   ix19157 : inv02 port map ( Y=>nx18783, A=>nx3360);
   ix19158 : nor02_2x port map ( Y=>nx18784, A0=>nx18897, A1=>
      write_base_data_out_6);
   ix19159 : and02 port map ( Y=>nx18785, A0=>nx17326, A1=>nx17199);
   ix19160 : inv01 port map ( Y=>nx18786, A=>nx18796);
   ix19161 : and02 port map ( Y=>nx18787, A0=>nx18898, A1=>nx18896);
   ix19162 : aoi43 port map ( Y=>nx18788, A0=>nx18796, A1=>nx18783, A2=>
      nx18784, A3=>nx18785, B0=>nx18786, B1=>nx18902, B2=>nx18787);
   reg_nx17323 : nor02_2x port map ( Y=>nx17323, A0=>nx18782, A1=>nx18788);
   ix19163 : inv02 port map ( Y=>nx18789, A=>nx18902);
   ix19164 : nand02_2x port map ( Y=>nx18790, A0=>nx18789, A1=>nx18787);
   reg_nx3934 : oai222 port map ( Y=>nx3934, A0=>nx18786, A1=>nx17326, B0=>
      nx18787, B1=>nx17326, C0=>nx18796, C1=>nx18790);
   ix19165 : inv02 port map ( Y=>nx18791, A=>nx18896);
   ix19166 : inv02 port map ( Y=>nx18792, A=>nx18898);
   reg_nx3644 : nor02_2x port map ( Y=>nx3644, A0=>nx18791, A1=>nx18796);
   ix19167 : inv02 port map ( Y=>nx18793, A=>write_base_data_out_6);
   ix19168 : and04 port map ( Y=>nx18794, A0=>nx18796, A1=>nx18783, A2=>
      nx17199, A3=>nx18793);
   ix19169 : nor02_2x port map ( Y=>nx18795, A0=>nx18794, A1=>nx3644);
   reg_nx17196 : nor02_2x port map ( Y=>nx17196, A0=>nx18782, A1=>nx18795);
   reg_nx3884 : oai321 port map ( Y=>nx3884, A0=>nx18797, A1=>nx18791, A2=>
      nx18898, B0=>nx18792, B1=>nx3644, C0=>nx17196);
   reg_nx3928 : nor04_2x port map ( Y=>nx3928, A0=>nx18797, A1=>nx18789, A2
      =>nx18792, A3=>nx18791);
   reg_nx17302 : oai322 port map ( Y=>nx17302, A0=>nx18797, A1=>nx18792, A2
      =>nx18791, B0=>nx18898, B1=>nx18896, C0=>nx18786, C1=>nx18898);
   reg_nx3650 : oai22 port map ( Y=>nx3650, A0=>nx18797, A1=>nx18896, B0=>
      nx18786, B1=>nx17199);
   reg_nx17172 : oai21 port map ( Y=>nx17172, A0=>nx3360, A1=>
      write_base_data_out_6, B0=>nx18797);
   reg_nx3600 : nand02_2x port map ( Y=>nx3600, A0=>nx17067, A1=>nx17172);
   ix19170 : buf04 port map ( Y=>nx18796, A=>nx17175);
   ix19171 : buf04 port map ( Y=>nx18797, A=>nx17175);
   ix19172 : inv02 port map ( Y=>nx18798, A=>nx18683);
   ix19173 : oai332 port map ( Y=>nx18799, A0=>nx18684, A1=>nx18798, A2=>
      nx17204, B0=>nx18684, B1=>nx18685, B2=>nx18686, C0=>nx18900, C1=>
      nx15816);
   ix19174 : nor02_2x port map ( Y=>nx18800, A0=>nx18680, A1=>nx17331);
   ix19175 : inv01 port map ( Y=>nx18801, A=>nx18684);
   ix19176 : inv02 port map ( Y=>nx18802, A=>nx17204);
   ix19177 : nand03_2x port map ( Y=>nx18803, A0=>nx18682, A1=>nx18801, A2=>
      nx18802);
   ix19178 : oai332 port map ( Y=>nx18804, A0=>nx18803, A1=>nx18680, A2=>
      nx17331, B0=>nx18687, B1=>nx18680, B2=>nx18688, C0=>nx18904, C1=>
      nx15806);
   ix19179 : aoi21 port map ( Y=>nx18805, A0=>nx19298, A1=>nx18800, B0=>
      nx19300);
   ix19180 : oai22 port map ( Y=>nx18806, A0=>nx18798, A1=>nx17204, B0=>
      nx18685, B1=>nx18686);
   ix19181 : nor02_2x port map ( Y=>nx18807, A0=>nx18900, A1=>nx15816);
   reg_NOT_nx3910 : aoi321 port map ( Y=>NOT_nx3910, A0=>nx18801, A1=>
      nx18682, A2=>nx18802, B0=>nx18806, B1=>nx18801, C0=>nx18807);
   ix19182 : inv02 port map ( Y=>nx18808, A=>img_addr_offset_11);
   ix19183 : inv02 port map ( Y=>nx18809, A=>img_base_addr_11);
   ix19184 : oai21 port map ( Y=>nx18810, A0=>nx18808, A1=>nx18809, B0=>
      nx17472);
   ix19185 : and02 port map ( Y=>nx18811, A0=>nx17425, A1=>nx17421);
   ix19186 : inv02 port map ( Y=>nx18812, A=>nx17548);
   ix19187 : inv02 port map ( Y=>nx18813, A=>nx17552);
   ix19188 : aoi22 port map ( Y=>nx18814, A0=>nx17548, A1=>nx17552, B0=>
      nx18812, B1=>nx18813);
   ix19189 : oai22 port map ( Y=>nx18815, A0=>nx18813, A1=>nx17548, B0=>
      nx18812, B1=>nx17552);
   ix19190 : nand02_2x port map ( Y=>nx18816, A0=>nx18815, A1=>nx17533);
   reg_nx17531 : oai21 port map ( Y=>nx17531, A0=>nx18839, A1=>nx18814, B0=>
      nx18816);
   ix19191 : inv02 port map ( Y=>nx18817, A=>nx17859);
   reg_nx17571 : ao32 port map ( Y=>nx17571, A0=>nx18716, A1=>nx18884, A2=>
      nx17323, B0=>nx18884, B1=>nx18817);
   ix19192 : nor02ii port map ( Y=>nx18818, A0=>nx18713, A1=>nx18716);
   ix19193 : inv01 port map ( Y=>nx18819, A=>nx17561);
   ix19194 : inv02 port map ( Y=>nx18820, A=>nx18143);
   reg_nx18135 : inv02 port map ( Y=>nx18135, A=>nx2664);
   ix19195 : oai22 port map ( Y=>nx18821, A0=>nx18135, A1=>nx17509, B0=>
      nx17566, B1=>nx18139);
   ix19196 : aoi321 port map ( Y=>nx18822, A0=>nx18818, A1=>
      argmax_ready_EXMPLR, A2=>nx17323, B0=>nx18819, B1=>nx18820, C0=>
      nx18821);
   reg_mem_addr_out_12 : oai221 port map ( Y=>mem_addr_out(12), A0=>nx18091, 
      A1=>nx17531, B0=>nx17556, B1=>nx17571, C0=>nx18822);
   reg_nx18075 : inv02 port map ( Y=>nx18075, A=>argmax_ready_EXMPLR);
   reg_nx17536 : oai22 port map ( Y=>nx17536, A0=>nx18812, A1=>nx18813, B0=>
      nx17548, B1=>nx17552);
   ix19197 : inv01 port map ( Y=>nx18823, A=>nx18716);
   ix19198 : inv02 port map ( Y=>nx18824, A=>nx17323);
   reg_nx18213 : nor03_2x port map ( Y=>nx18213, A0=>nx18713, A1=>nx18823, 
      A2=>nx18824);
   reg_nx17977 : inv02 port map ( Y=>nx17977, A=>nx18884);
   reg_nx4250 : oai22 port map ( Y=>nx4250, A0=>nx17425, A1=>nx17421, B0=>
      nx18811, B1=>nx17406);
   reg_nx17450 : and02 port map ( Y=>nx17450, A0=>nx18716, A1=>nx17323);
   ix19199 : nor02_2x port map ( Y=>nx18825, A0=>nx17425, A1=>nx17421);
   reg_nx17409 : ao21 port map ( Y=>nx17409, A0=>nx17425, A1=>nx17421, B0=>
      nx18825);
   ix19200 : inv02 port map ( Y=>nx18826, A=>nx15696);
   ix19201 : inv02 port map ( Y=>nx18827, A=>nx17199);
   ix19202 : nand02_2x port map ( Y=>nx18828, A0=>nx15696, A1=>nx17199);
   ix19203 : or02 port map ( Y=>nx18829, A0=>nx18737, A1=>nx18739);
   ix19204 : aoi21 port map ( Y=>nx18830, A0=>nx18592, A1=>nx18735, B0=>
      nx18829);
   ix19205 : nor02_2x port map ( Y=>nx18831, A0=>nx18739, A1=>nx18734);
   ix19206 : and02 port map ( Y=>nx18832, A0=>nx18592, A1=>nx18735);
   reg_nx17247 : oai32 port map ( Y=>nx17247, A0=>nx18832, A1=>nx18737, A2=>
      nx18739, B0=>nx18739, B1=>nx18734);
   reg_nx17250 : oai22 port map ( Y=>nx17250, A0=>nx18826, A1=>nx18827, B0=>
      nx15696, B1=>nx17199);
   ix19207 : inv02 port map ( Y=>nx18833, A=>nx18756);
   ix19208 : inv02 port map ( Y=>nx18834, A=>nx17345);
   ix19209 : nor02ii port map ( Y=>nx18835, A0=>nx18811, A1=>nx18810);
   ix19210 : oai22 port map ( Y=>nx18836, A0=>nx17425, A1=>nx17421, B0=>
      nx18808, B1=>nx18809);
   ix19211 : and02 port map ( Y=>nx18837, A0=>img_addr_offset_9, A1=>
      img_base_addr_9);
   ix19212 : aoi322 port map ( Y=>nx18838, A0=>nx18833, A1=>nx18834, A2=>
      nx18835, B0=>nx18810, B1=>nx18836, C0=>nx18835, C1=>nx18837);
   reg_nx17533 : inv02 port map ( Y=>nx17533, A=>nx18838);
   ix19213 : inv02 port map ( Y=>nx18839, A=>nx18838);
   reg_nx17406 : oai22 port map ( Y=>nx17406, A0=>nx18833, A1=>nx18837, B0=>
      nx18834, B1=>nx18837);
   ix19214 : nand02_2x port map ( Y=>nx18840, A0=>nx18826, A1=>nx18827);
   ix19215 : nor02ii port map ( Y=>nx18841, A0=>nx18831, A1=>nx18828);
   ix19216 : and02 port map ( Y=>nx18842, A0=>nx18826, A1=>nx18827);
   ix19217 : nor02_2x port map ( Y=>nx18843, A0=>nx18841, A1=>nx18842);
   reg_nx3760 : aoi21 port map ( Y=>nx3760, A0=>nx18830, A1=>nx18840, B0=>
      nx18843);
   reg_nx17577 : inv01 port map ( Y=>nx17577, A=>nx18709);
   reg_nx4736 : nand02_2x port map ( Y=>nx4736, A0=>nx17679, A1=>nx17577);
   ix19218 : nand02_2x port map ( Y=>nx18844, A0=>nx18896, A1=>
      bias_offset_data_out_7);
   ix19219 : and02 port map ( Y=>nx18845, A0=>nx18894, A1=>nx17135);
   ix19220 : nor02_2x port map ( Y=>nx18846, A0=>nx18894, A1=>nx17135);
   ix19221 : aoi22 port map ( Y=>nx18847, A0=>nx18844, A1=>nx18849, B0=>
      nx17210, B1=>nx18844);
   reg_nx17257 : inv01 port map ( Y=>nx17257, A=>nx18847);
   reg_nx3728 : oai22 port map ( Y=>nx3728, A0=>nx18894, A1=>nx17135, B0=>
      nx18845, B1=>nx18659);
   reg_nx17130 : ao21 port map ( Y=>nx17130, A0=>nx18894, A1=>nx17135, B0=>
      nx18846);
   ix19222 : inv02 port map ( Y=>nx18848, A=>nx18846);
   ix19223 : ao22 port map ( Y=>nx18849, A0=>nx18845, A1=>nx18848, B0=>
      nx18659, B1=>nx18848);
   ix19224 : inv02 port map ( Y=>nx18850, A=>nx4580);
   ix19225 : oai21 port map ( Y=>nx18851, A0=>nx18850, A1=>nx17591, B0=>
      nx18718);
   ix19226 : inv02 port map ( Y=>nx18852, A=>nx18900);
   ix19227 : inv02 port map ( Y=>nx18853, A=>nx17265);
   ix19228 : nand02_2x port map ( Y=>nx18854, A0=>nx18900, A1=>nx17265);
   ix19229 : aoi22 port map ( Y=>nx18855, A0=>nx18852, A1=>nx18853, B0=>
      nx18847, B1=>nx18854);
   reg_nx4012 : inv02 port map ( Y=>nx4012, A=>nx18855);
   ix19230 : inv02 port map ( Y=>nx18856, A=>nx18855);
   ix19231 : inv02 port map ( Y=>nx18857, A=>nx18855);
   ix19232 : nor02_2x port map ( Y=>nx18858, A0=>nx18900, A1=>nx17265);
   reg_nx17260 : ao21 port map ( Y=>nx17260, A0=>nx18900, A1=>nx17265, B0=>
      nx18858);
   ix19233 : oai22 port map ( Y=>nx18859, A0=>nx18892, A1=>nx18890, B0=>
      nx18892, B1=>nx18887);
   ix19234 : inv01 port map ( Y=>nx18860, A=>nx16934);
   ix19235 : ao22 port map ( Y=>nx18861, A0=>nx18892, A1=>nx18890, B0=>
      nx18892, B1=>nx18887);
   ix19236 : inv01 port map ( Y=>nx18862, A=>nx18888);
   ix19237 : inv01 port map ( Y=>nx18863, A=>nx18892);
   ix19238 : inv02 port map ( Y=>nx18864, A=>nx18890);
   ix19239 : oai33 port map ( Y=>nx18865, A0=>nx18862, A1=>nx18863, A2=>
      nx18864, B0=>nx18888, B1=>nx18892, B2=>nx18890);
   ix19240 : aoi221 port map ( Y=>nx18866, A0=>nx18859, A1=>nx18860, B0=>
      nx16934, B1=>nx18861, C0=>nx18865);
   reg_nx16998 : inv01 port map ( Y=>nx16998, A=>nx18866);
   ix19241 : inv01 port map ( Y=>nx18867, A=>nx18866);
   ix19242 : and02 port map ( Y=>nx18868, A0=>nx18888, A1=>nx18890);
   reg_nx3216 : oai22 port map ( Y=>nx3216, A0=>nx18888, A1=>nx18890, B0=>
      nx18868, B1=>nx16934);
   reg_nx16937 : oai22 port map ( Y=>nx16937, A0=>nx18862, A1=>nx18864, B0=>
      nx18888, B1=>nx18890);
   ix19243 : nor02_2x port map ( Y=>nx18869, A0=>nx18722, A1=>nx17464);
   ix19244 : nand03_2x port map ( Y=>nx18870, A0=>nx18869, A1=>nx18856, A2=>
      nx18720);
   ix19245 : and03 port map ( Y=>nx18871, A0=>nx18719, A1=>nx18902, A2=>
      bias_offset_data_out_9);
   ix19246 : nor02_2x port map ( Y=>nx18872, A0=>nx18871, A1=>nx18721);
   ix19247 : oai332 port map ( Y=>nx18873, A0=>nx18872, A1=>nx18722, A2=>
      nx17464, B0=>nx18723, B1=>nx18722, B2=>nx18724, C0=>nx18910, C1=>
      nx17519);
   ix19248 : inv02 port map ( Y=>nx18874, A=>nx18873);
   reg_nx4580 : nand02_2x port map ( Y=>nx4580, A0=>nx18870, A1=>nx18874);
   ix19249 : aoi321 port map ( Y=>nx18875, A0=>nx18719, A1=>nx18902, A2=>
      bias_offset_data_out_9, B0=>nx18856, B1=>nx18720, C0=>nx18721);
   ix19250 : nand02_2x port map ( Y=>nx18876, A0=>write_base_data_out_5, A1
      =>new_size_squared_out_5);
   ix19251 : aoi32 port map ( Y=>nx18877, A0=>nx18764, A1=>nx18562, A2=>
      nx18765, B0=>nx18560, B1=>nx18561);
   ix19252 : oai332 port map ( Y=>nx18878, A0=>nx18877, A1=>nx18767, A2=>
      nx18766, B0=>nx18767, B1=>nx18768, B2=>nx18769, C0=>nx18892, C1=>
      nx15837);
   ix19253 : inv02 port map ( Y=>nx18879, A=>nx18878);
   ix19254 : aoi22 port map ( Y=>nx18880, A0=>nx17074, A1=>nx18876, B0=>
      nx18876, B1=>nx18879);
   reg_nx17142 : inv02 port map ( Y=>nx17142, A=>nx18880);
   ix19255 : inv02 port map ( Y=>nx18881, A=>nx18880);
   ix19256 : inv02 port map ( Y=>nx18882, A=>nx18880);
   ix19257 : buf16 port map ( Y=>nx18883, A=>nx18309);
   ix19258 : buf16 port map ( Y=>nx18884, A=>nx18309);
   ix19259 : buf16 port map ( Y=>nx18885, A=>nx16878);
   ix19260 : buf16 port map ( Y=>nx18886, A=>nx16878);
   ix19261 : buf16 port map ( Y=>nx18887, A=>nx16348);
   ix19262 : buf16 port map ( Y=>nx18888, A=>nx16348);
   ix19263 : buf16 port map ( Y=>nx18889, A=>nx16945);
   ix19264 : buf16 port map ( Y=>nx18890, A=>nx16945);
   ix19265 : buf16 port map ( Y=>nx18891, A=>nx17002);
   ix19266 : buf16 port map ( Y=>nx18892, A=>nx17002);
   ix19267 : buf16 port map ( Y=>nx18893, A=>nx17138);
   ix19268 : buf16 port map ( Y=>nx18894, A=>nx17138);
   ix19269 : buf16 port map ( Y=>nx18895, A=>write_base_data_out_7);
   ix19270 : buf16 port map ( Y=>nx18896, A=>write_base_data_out_7);
   ix19271 : buf16 port map ( Y=>nx18897, A=>write_base_data_out_8);
   ix19272 : buf16 port map ( Y=>nx18898, A=>write_base_data_out_8);
   ix19273 : buf16 port map ( Y=>nx18899, A=>nx17268);
   ix19274 : buf16 port map ( Y=>nx18900, A=>nx17268);
   ix19275 : buf16 port map ( Y=>nx18901, A=>write_base_data_out_9);
   ix19276 : buf16 port map ( Y=>nx18902, A=>write_base_data_out_9);
   ix19277 : buf16 port map ( Y=>nx18903, A=>nx17395);
   ix19278 : buf16 port map ( Y=>nx18904, A=>nx17395);
   ix19279 : buf16 port map ( Y=>nx18905, A=>write_base_data_out_11);
   ix19280 : buf16 port map ( Y=>nx18906, A=>write_base_data_out_11);
   ix19281 : buf16 port map ( Y=>nx18907, A=>nx17453);
   ix19282 : buf16 port map ( Y=>nx18908, A=>nx17453);
   ix19283 : buf16 port map ( Y=>nx18909, A=>nx17522);
   ix19284 : buf16 port map ( Y=>nx18910, A=>nx17522);
   ix19285 : buf16 port map ( Y=>nx18911, A=>current_state_26);
   ix19286 : buf16 port map ( Y=>nx18912, A=>current_state_26);
   ix19287 : buf16 port map ( Y=>nx18913, A=>nx17580);
   ix19288 : buf16 port map ( Y=>nx18914, A=>nx17580);
   ix19289 : buf16 port map ( Y=>nx18915, A=>nx17649);
   ix19290 : buf16 port map ( Y=>nx18916, A=>nx17649);
   ix19291 : inv02 port map ( Y=>nx19292, A=>nx18219);
   ix19293 : inv02 port map ( Y=>nx19294, A=>nx19292);
   ix19295 : inv02 port map ( Y=>nx19296, A=>nx19292);
   ix19297 : buf02 port map ( Y=>nx19298, A=>nx18799);
   ix19299 : buf02 port map ( Y=>nx19300, A=>nx18804);
   ix19301 : inv02 port map ( Y=>nx19302, A=>nx18219);
   ix19307 : inv02 port map ( Y=>nx19308, A=>nx16222);
end Mixed ;

