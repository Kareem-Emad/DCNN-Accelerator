library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library dcnn;

entity Ram is
	port (
		clk 					: in std_logic; -- the clock
		read_in					: in std_logic;
		write_in 				: in std_logic;
		address_in              : in std_logic_vector(15 downto 0); -- 256 addresses.
		data_in                 : in std_logic_vector(15 downto 0);
		data_out                : out std_logic_vector(15 downto 0));
end entity Ram;

architecture Behavioral of Ram is
	type ram_type is array (0 to 65536-1) of std_logic_vector(15 downto 0);
	signal ram : ram_type := (
		--R0=0,...,R5=5
		0 => X"0001", -- number of layers
		-- Start of Layer 1
		1 => X"0000", -- layer type (0: Conv, 1: Pool, 2: FC)
		2 => X"0002", -- Number of filters in layer
		3 => X"0003", -- Filter size
		4 => X"001A", -- New Layer Width
		5 => X"02A4", -- (New Layer Width)^2
		6 => X"0548", -- (New Layer Width)^2 * Number of filters in layer
		7 => X"1235", -- bias of filter 1
		8 => X"0001", -- start of filter 1
		9 => X"0002",
		10 => X"0003",
		11 => X"0004",
		12 => X"0005",
		13 => X"0006",
		14 => X"0007",
		15 => X"0008", 
		16 => X"0009", -- end of filter 1
		17 => X"AAAA", -- filter 2 bias
		18 => X"000B", -- start of filter 2
		19 => X"000C",
		20 => X"000D",
		21 => X"000E",
		22 => X"000F",
		23 => X"0010",
		24 => X"0011", -- end of filter 2
		-- start of image
		39000 => X"0001",
		39001 => X"0002",
		39002 => X"0003",
		39003 => X"0004",
		39004 => X"0005",
		39005 => X"0006",
		39006 => X"0007",
		39007 => X"0008",
		39008 => X"0009",
		39009 => X"0010",
		39010 => X"0011",
		39011 => X"0012",
		39012 => X"0013",
		39013 => X"0014",
		39014 => X"0015",
		39015 => X"0016",
		39016 => X"0017",
		39017 => X"0018",
		39018 => X"0019",
		39019 => X"0020",
		39020 => X"0021",
		39021 => X"0022",
		39022 => X"0023",
		39023 => X"0024",
		39024 => X"0025",
		39025 => X"0026",
		39026 => X"0027",
		39027 => X"0028",
		39028 => X"0001",
		39029 => X"0002",
		39030 => X"0003",
		39031 => X"0004",
		39032 => X"0005",
		39033 => X"0006",
		39034 => X"0007",
		39035 => X"0008",
		39036 => X"0009",
		39037 => X"0010",
		39038 => X"0011",
		39039 => X"0012",
		39040 => X"0013",
		39041 => X"0014",
		39042 => X"0015",
		39043 => X"0016",
		39044 => X"0017",
		39045 => X"0018",
		39046 => X"0019",
		39047 => X"0020",
		39048 => X"0021",
		39049 => X"0022",
		39050 => X"0023",
		39051 => X"0024",
		39052 => X"0025",
		39053 => X"0026",
		39054 => X"0027",
		39055 => X"0028",
		39056 => X"0001",
		39057 => X"0002",
		39058 => X"0003",
		39059 => X"0004",
		39060 => X"0005",
		39061 => X"0006",
		39062 => X"0007",
		39063 => X"0008",
		39064 => X"0009",
		39065 => X"0010",
		39066 => X"0011",
		39067 => X"0012",
		39068 => X"0013",
		39069 => X"0014",
		39070 => X"0015",
		39071 => X"0016",
		39072 => X"0017",
		39073 => X"0018",
		39074 => X"0019",
		39075 => X"0020",
		39076 => X"0021",
		39077 => X"0022",
		39078 => X"0023",
		39079 => X"0024",
		39080 => X"0025",
		39081 => X"0026",
		39082 => X"0027",
		39083 => X"0028",
		39084 => X"0001",
		39085 => X"0002",
		39086 => X"0003",
		39087 => X"0004",
		39088 => X"0005",
		39089 => X"0006",
		39090 => X"0007",
		39091 => X"0008",
		39092 => X"0009",
		39093 => X"0010",
		39094 => X"0011",
		39095 => X"0012",
		39096 => X"0013",
		39097 => X"0014",
		39098 => X"0015",
		39099 => X"0016",
		39100 => X"0017",
		39101 => X"0018",
		39102 => X"0019",
		39103 => X"0020",
		39104 => X"0021",
		39105 => X"0022",
		39106 => X"0023",
		39107 => X"0024",
		39108 => X"0025",
		39109 => X"0026",
		39110 => X"0027",
		39111 => X"0028",
		39112 => X"0001",
		39113 => X"0002",
		39114 => X"0003",
		39115 => X"0004",
		39116 => X"0005",
		39117 => X"0006",
		39118 => X"0007",
		39119 => X"0008",
		39120 => X"0009",
		39121 => X"0010",
		39122 => X"0011",
		39123 => X"0012",
		39124 => X"0013",
		39125 => X"0014",
		39126 => X"0015",
		39127 => X"0016",
		39128 => X"0017",
		39129 => X"0018",
		39130 => X"0019",
		39131 => X"0020",
		39132 => X"0021",
		39133 => X"0022",
		39134 => X"0023",
		39135 => X"0024",
		39136 => X"0025",
		39137 => X"0026",
		39138 => X"0027",
		39139 => X"0028",
		39140 => X"0002",
		39141 => X"0004",
		39142 => X"0006",
		39143 => X"0008",
		39144 => X"0010",
		39145 => X"0012",
		39146 => X"0014",
		39147 => X"0016",
		39148 => X"0018",
		39149 => X"0020",
		39150 => X"0022",
		39151 => X"0024",
		39152 => X"0026",
		39153 => X"0028",
		39154 => X"0030",
		39155 => X"0032",
		39156 => X"0034",
		39157 => X"0036",
		39158 => X"0038",
		39159 => X"0040",
		39160 => X"0042",
		39161 => X"0044",
		39162 => X"0046",
		39163 => X"0048",
		39164 => X"0050",
		39165 => X"0052",
		39166 => X"0054",
		39167 => X"0056",
		39168 => X"0002",
		39169 => X"0004",
		39170 => X"0006",
		39171 => X"0008",
		39172 => X"0010",
		39173 => X"0012",
		39174 => X"0014",
		39175 => X"0016",
		39176 => X"0018",
		39177 => X"0020",
		39178 => X"0022",
		39179 => X"0024",
		39180 => X"0026",
		39181 => X"0028",
		39182 => X"0030",
		39183 => X"0032",
		39184 => X"0034",
		39185 => X"0036",
		39186 => X"0038",
		39187 => X"0040",
		39188 => X"0042",
		39189 => X"0044",
		39190 => X"0046",
		39191 => X"0048",
		39192 => X"0050",
		39193 => X"0052",
		39194 => X"0054",
		39195 => X"0056",
		39196 => X"0002",
		39197 => X"0004",
		39198 => X"0006",
		39199 => X"0008",
		39200 => X"0010",
		39201 => X"0012",
		39202 => X"0014",
		39203 => X"0016",
		39204 => X"0018",
		39205 => X"0020",
		39206 => X"0022",
		39207 => X"0024",
		39208 => X"0026",
		39209 => X"0028",
		39210 => X"0030",
		39211 => X"0032",
		39212 => X"0034",
		39213 => X"0036",
		39214 => X"0038",
		39215 => X"0040",
		39216 => X"0042",
		39217 => X"0044",
		39218 => X"0046",
		39219 => X"0048",
		39220 => X"0050",
		39221 => X"0052",
		39222 => X"0054",
		39223 => X"0056",
		39224 => X"0002",
		39225 => X"0004",
		39226 => X"0006",
		39227 => X"0008",
		39228 => X"0010",
		39229 => X"0012",
		39230 => X"0014",
		39231 => X"0016",
		39232 => X"0018",
		39233 => X"0020",
		39234 => X"0022",
		39235 => X"0024",
		39236 => X"0026",
		39237 => X"0028",
		39238 => X"0030",
		39239 => X"0032",
		39240 => X"0034",
		39241 => X"0036",
		39242 => X"0038",
		39243 => X"0040",
		39244 => X"0042",
		39245 => X"0044",
		39246 => X"0046",
		39247 => X"0048",
		39248 => X"0050",
		39249 => X"0052",
		39250 => X"0054",
		39251 => X"0056",
		39252 => X"0002",
		39253 => X"0004",
		39254 => X"0006",
		39255 => X"0008",
		39256 => X"0010",
		39257 => X"0012",
		39258 => X"0014",
		39259 => X"0016",
		39260 => X"0018",
		39261 => X"0020",
		39262 => X"0022",
		39263 => X"0024",
		39264 => X"0026",
		39265 => X"0028",
		39266 => X"0030",
		39267 => X"0032",
		39268 => X"0034",
		39269 => X"0036",
		39270 => X"0038",
		39271 => X"0040",
		39272 => X"0042",
		39273 => X"0044",
		39274 => X"0046",
		39275 => X"0048",
		39276 => X"0050",
		39277 => X"0052",
		39278 => X"0054",
		39279 => X"0056",
		39280 => X"0003",
		39281 => X"0006",
		39282 => X"0009",
		39283 => X"0012",
		39284 => X"0015",
		39285 => X"0018",
		39286 => X"0021",
		39287 => X"0024",
		39288 => X"0027",
		39289 => X"0030",
		39290 => X"0033",
		39291 => X"0036",
		39292 => X"0039",
		39293 => X"0042",
		39294 => X"0045",
		39295 => X"0048",
		39296 => X"0051",
		39297 => X"0054",
		39298 => X"0057",
		39299 => X"0060",
		39300 => X"0063",
		39301 => X"0066",
		39302 => X"0069",
		39303 => X"0072",
		39304 => X"0075",
		39305 => X"0078",
		39306 => X"0081",
		39307 => X"0084",
		39308 => X"0003",
		39309 => X"0006",
		39310 => X"0009",
		39311 => X"0012",
		39312 => X"0015",
		39313 => X"0018",
		39314 => X"0021",
		39315 => X"0024",
		39316 => X"0027",
		39317 => X"0030",
		39318 => X"0033",
		39319 => X"0036",
		39320 => X"0039",
		39321 => X"0042",
		39322 => X"0045",
		39323 => X"0048",
		39324 => X"0051",
		39325 => X"0054",
		39326 => X"0057",
		39327 => X"0060",
		39328 => X"0063",
		39329 => X"0066",
		39330 => X"0069",
		39331 => X"0072",
		39332 => X"0075",
		39333 => X"0078",
		39334 => X"0081",
		39335 => X"0084",
		39336 => X"0003",
		39337 => X"0006",
		39338 => X"0009",
		39339 => X"0012",
		39340 => X"0015",
		39341 => X"0018",
		39342 => X"0021",
		39343 => X"0024",
		39344 => X"0027",
		39345 => X"0030",
		39346 => X"0033",
		39347 => X"0036",
		39348 => X"0039",
		39349 => X"0042",
		39350 => X"0045",
		39351 => X"0048",
		39352 => X"0051",
		39353 => X"0054",
		39354 => X"0057",
		39355 => X"0060",
		39356 => X"0063",
		39357 => X"0066",
		39358 => X"0069",
		39359 => X"0072",
		39360 => X"0075",
		39361 => X"0078",
		39362 => X"0081",
		39363 => X"0084",
		39364 => X"0003",
		39365 => X"0006",
		39366 => X"0009",
		39367 => X"0012",
		39368 => X"0015",
		39369 => X"0018",
		39370 => X"0021",
		39371 => X"0024",
		39372 => X"0027",
		39373 => X"0030",
		39374 => X"0033",
		39375 => X"0036",
		39376 => X"0039",
		39377 => X"0042",
		39378 => X"0045",
		39379 => X"0048",
		39380 => X"0051",
		39381 => X"0054",
		39382 => X"0057",
		39383 => X"0060",
		39384 => X"0063",
		39385 => X"0066",
		39386 => X"0069",
		39387 => X"0072",
		39388 => X"0075",
		39389 => X"0078",
		39390 => X"0081",
		39391 => X"0084",
		39392 => X"0003",
		39393 => X"0006",
		39394 => X"0009",
		39395 => X"0012",
		39396 => X"0015",
		39397 => X"0018",
		39398 => X"0021",
		39399 => X"0024",
		39400 => X"0027",
		39401 => X"0030",
		39402 => X"0033",
		39403 => X"0036",
		39404 => X"0039",
		39405 => X"0042",
		39406 => X"0045",
		39407 => X"0048",
		39408 => X"0051",
		39409 => X"0054",
		39410 => X"0057",
		39411 => X"0060",
		39412 => X"0063",
		39413 => X"0066",
		39414 => X"0069",
		39415 => X"0072",
		39416 => X"0075",
		39417 => X"0078",
		39418 => X"0081",
		39419 => X"0084",
		39420 => X"0004",
		39421 => X"0008",
		39422 => X"0012",
		39423 => X"0016",
		39424 => X"0020",
		39425 => X"0024",
		39426 => X"0028",
		39427 => X"0032",
		39428 => X"0036",
		39429 => X"0040",
		39430 => X"0044",
		39431 => X"0048",
		39432 => X"0052",
		39433 => X"0056",
		39434 => X"0060",
		39435 => X"0064",
		39436 => X"0068",
		39437 => X"0072",
		39438 => X"0076",
		39439 => X"0080",
		39440 => X"0084",
		39441 => X"0088",
		39442 => X"0092",
		39443 => X"0096",
		39444 => X"0100",
		39445 => X"0104",
		39446 => X"0108",
		39447 => X"0112",
		39448 => X"0004",
		39449 => X"0008",
		39450 => X"0012",
		39451 => X"0016",
		39452 => X"0020",
		39453 => X"0024",
		39454 => X"0028",
		39455 => X"0032",
		39456 => X"0036",
		39457 => X"0040",
		39458 => X"0044",
		39459 => X"0048",
		39460 => X"0052",
		39461 => X"0056",
		39462 => X"0060",
		39463 => X"0064",
		39464 => X"0068",
		39465 => X"0072",
		39466 => X"0076",
		39467 => X"0080",
		39468 => X"0084",
		39469 => X"0088",
		39470 => X"0092",
		39471 => X"0096",
		39472 => X"0100",
		39473 => X"0104",
		39474 => X"0108",
		39475 => X"0112",
		39476 => X"0004",
		39477 => X"0008",
		39478 => X"0012",
		39479 => X"0016",
		39480 => X"0020",
		39481 => X"0024",
		39482 => X"0028",
		39483 => X"0032",
		39484 => X"0036",
		39485 => X"0040",
		39486 => X"0044",
		39487 => X"0048",
		39488 => X"0052",
		39489 => X"0056",
		39490 => X"0060",
		39491 => X"0064",
		39492 => X"0068",
		39493 => X"0072",
		39494 => X"0076",
		39495 => X"0080",
		39496 => X"0084",
		39497 => X"0088",
		39498 => X"0092",
		39499 => X"0096",
		39500 => X"0100",
		39501 => X"0104",
		39502 => X"0108",
		39503 => X"0112",
		39504 => X"0004",
		39505 => X"0008",
		39506 => X"0012",
		39507 => X"0016",
		39508 => X"0020",
		39509 => X"0024",
		39510 => X"0028",
		39511 => X"0032",
		39512 => X"0036",
		39513 => X"0040",
		39514 => X"0044",
		39515 => X"0048",
		39516 => X"0052",
		39517 => X"0056",
		39518 => X"0060",
		39519 => X"0064",
		39520 => X"0068",
		39521 => X"0072",
		39522 => X"0076",
		39523 => X"0080",
		39524 => X"0084",
		39525 => X"0088",
		39526 => X"0092",
		39527 => X"0096",
		39528 => X"0100",
		39529 => X"0104",
		39530 => X"0108",
		39531 => X"0112",
		39532 => X"0004",
		39533 => X"0008",
		39534 => X"0012",
		39535 => X"0016",
		39536 => X"0020",
		39537 => X"0024",
		39538 => X"0028",
		39539 => X"0032",
		39540 => X"0036",
		39541 => X"0040",
		39542 => X"0044",
		39543 => X"0048",
		39544 => X"0052",
		39545 => X"0056",
		39546 => X"0060",
		39547 => X"0064",
		39548 => X"0068",
		39549 => X"0072",
		39550 => X"0076",
		39551 => X"0080",
		39552 => X"0084",
		39553 => X"0088",
		39554 => X"0092",
		39555 => X"0096",
		39556 => X"0100",
		39557 => X"0104",
		39558 => X"0108",
		39559 => X"0112",
		39560 => X"0005",
		39561 => X"0010",
		39562 => X"0015",
		39563 => X"0020",
		39564 => X"0025",
		39565 => X"0030",
		39566 => X"0035",
		39567 => X"0040",
		39568 => X"0045",
		39569 => X"0050",
		39570 => X"0055",
		39571 => X"0060",
		39572 => X"0065",
		39573 => X"0070",
		39574 => X"0075",
		39575 => X"0080",
		39576 => X"0085",
		39577 => X"0090",
		39578 => X"0095",
		39579 => X"0100",
		39580 => X"0105",
		39581 => X"0110",
		39582 => X"0115",
		39583 => X"0120",
		39584 => X"0125",
		39585 => X"0130",
		39586 => X"0135",
		39587 => X"0140",
		39588 => X"0005",
		39589 => X"0010",
		39590 => X"0015",
		39591 => X"0020",
		39592 => X"0025",
		39593 => X"0030",
		39594 => X"0035",
		39595 => X"0040",
		39596 => X"0045",
		39597 => X"0050",
		39598 => X"0055",
		39599 => X"0060",
		39600 => X"0065",
		39601 => X"0070",
		39602 => X"0075",
		39603 => X"0080",
		39604 => X"0085",
		39605 => X"0090",
		39606 => X"0095",
		39607 => X"0100",
		39608 => X"0105",
		39609 => X"0110",
		39610 => X"0115",
		39611 => X"0120",
		39612 => X"0125",
		39613 => X"0130",
		39614 => X"0135",
		39615 => X"0140",
		39616 => X"0005",
		39617 => X"0010",
		39618 => X"0015",
		39619 => X"0020",
		39620 => X"0025",
		39621 => X"0030",
		39622 => X"0035",
		39623 => X"0040",
		39624 => X"0045",
		39625 => X"0050",
		39626 => X"0055",
		39627 => X"0060",
		39628 => X"0065",
		39629 => X"0070",
		39630 => X"0075",
		39631 => X"0080",
		39632 => X"0085",
		39633 => X"0090",
		39634 => X"0095",
		39635 => X"0100",
		39636 => X"0105",
		39637 => X"0110",
		39638 => X"0115",
		39639 => X"0120",
		39640 => X"0125",
		39641 => X"0130",
		39642 => X"0135",
		39643 => X"0140",
		39644 => X"0005",
		39645 => X"0010",
		39646 => X"0015",
		39647 => X"0020",
		39648 => X"0025",
		39649 => X"0030",
		39650 => X"0035",
		39651 => X"0040",
		39652 => X"0045",
		39653 => X"0050",
		39654 => X"0055",
		39655 => X"0060",
		39656 => X"0065",
		39657 => X"0070",
		39658 => X"0075",
		39659 => X"0080",
		39660 => X"0085",
		39661 => X"0090",
		39662 => X"0095",
		39663 => X"0100",
		39664 => X"0105",
		39665 => X"0110",
		39666 => X"0115",
		39667 => X"0120",
		39668 => X"0125",
		39669 => X"0130",
		39670 => X"0135",
		39671 => X"0140",
		39672 => X"0005",
		39673 => X"0010",
		39674 => X"0015",
		39675 => X"0020",
		39676 => X"0025",
		39677 => X"0030",
		39678 => X"0035",
		39679 => X"0040",
		39680 => X"0045",
		39681 => X"0050",
		39682 => X"0055",
		39683 => X"0060",
		39684 => X"0065",
		39685 => X"0070",
		39686 => X"0075",
		39687 => X"0080",
		39688 => X"0085",
		39689 => X"0090",
		39690 => X"0095",
		39691 => X"0100",
		39692 => X"0105",
		39693 => X"0110",
		39694 => X"0115",
		39695 => X"0120",
		39696 => X"0125",
		39697 => X"0130",
		39698 => X"0135",
		39699 => X"0140",
		39700 => X"0006",
		39701 => X"0012",
		39702 => X"0018",
		39703 => X"0024",
		39704 => X"0030",
		39705 => X"0036",
		39706 => X"0042",
		39707 => X"0048",
		39708 => X"0054",
		39709 => X"0060",
		39710 => X"0066",
		39711 => X"0072",
		39712 => X"0078",
		39713 => X"0084",
		39714 => X"0090",
		39715 => X"0096",
		39716 => X"0102",
		39717 => X"0108",
		39718 => X"0114",
		39719 => X"0120",
		39720 => X"0126",
		39721 => X"0132",
		39722 => X"0138",
		39723 => X"0144",
		39724 => X"0150",
		39725 => X"0156",
		39726 => X"0162",
		39727 => X"0168",
		39728 => X"0006",
		39729 => X"0012",
		39730 => X"0018",
		39731 => X"0024",
		39732 => X"0030",
		39733 => X"0036",
		39734 => X"0042",
		39735 => X"0048",
		39736 => X"0054",
		39737 => X"0060",
		39738 => X"0066",
		39739 => X"0072",
		39740 => X"0078",
		39741 => X"0084",
		39742 => X"0090",
		39743 => X"0096",
		39744 => X"0102",
		39745 => X"0108",
		39746 => X"0114",
		39747 => X"0120",
		39748 => X"0126",
		39749 => X"0132",
		39750 => X"0138",
		39751 => X"0144",
		39752 => X"0150",
		39753 => X"0156",
		39754 => X"0162",
		39755 => X"0168",
		39756 => X"0006",
		39757 => X"0012",
		39758 => X"0018",
		39759 => X"0024",
		39760 => X"0030",
		39761 => X"0036",
		39762 => X"0042",
		39763 => X"0048",
		39764 => X"0054",
		39765 => X"0060",
		39766 => X"0066",
		39767 => X"0072",
		39768 => X"0078",
		39769 => X"0084",
		39770 => X"0090",
		39771 => X"0096",
		39772 => X"0102",
		39773 => X"0108",
		39774 => X"0114",
		39775 => X"0120",
		39776 => X"0126",
		39777 => X"0132",
		39778 => X"0138",
		39779 => X"0144",
		39780 => X"0150",
		39781 => X"0156",
		39782 => X"0162",
		39783 => X"0168",

		-- start of output data
		39784 => X"1202",
		39785 => X"2101",
		others => X"BBBB"
	);
	begin
		-- Inputs data into the RAM on the falling edge of the clock.
		process(clk) is
			begin
				if falling_edge(clk) then  
					if write_in = '1' then
						ram(to_integer(unsigned(address_in))) <= data_in;
					end if;
				end if;
		end process;

		-- Outputs data asynchronously when the output is applied.
		data_out <= ram(to_integer(unsigned(address_in))) when (read_in = '1') else (15 downto 0 => '0');
end Behavioral;