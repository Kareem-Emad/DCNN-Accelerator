//
// Verilog description for cell DCNNChip, 
// Sun May 12 02:11:46 2019
//
// LeonardoSpectrum Level 3, 2018a.2 
//


module DCNNChip ( clk, reset, io_ready_in, io_done_out, mem_read_out, 
                  mem_write_out, mem_addr_out, mem_data_in, mem_data_out ) ;

    input clk ;
    input reset ;
    input io_ready_in ;
    output io_done_out ;
    output mem_read_out ;
    output mem_write_out ;
    output [15:0]mem_addr_out ;
    input [15:0]mem_data_in ;
    output [15:0]mem_data_out ;

    wire image_wind_en, image_wind_col_4__15, image_wind_col_4__14, 
         image_wind_col_4__13, image_wind_col_4__12, image_wind_col_4__11, 
         image_wind_col_4__10, image_wind_col_4__9, image_wind_col_4__8, 
         image_wind_col_4__7, image_wind_col_4__6, image_wind_col_4__5, 
         image_wind_col_4__4, image_wind_col_4__3, image_wind_col_4__2, 
         image_wind_col_4__1, image_wind_col_4__0, image_wind_col_3__15, 
         image_wind_col_3__14, image_wind_col_3__13, image_wind_col_3__12, 
         image_wind_col_3__11, image_wind_col_3__10, image_wind_col_3__9, 
         image_wind_col_3__8, image_wind_col_3__7, image_wind_col_3__6, 
         image_wind_col_3__5, image_wind_col_3__4, image_wind_col_3__3, 
         image_wind_col_3__2, image_wind_col_3__1, image_wind_col_3__0, 
         image_wind_col_2__15, image_wind_col_2__14, image_wind_col_2__13, 
         image_wind_col_2__12, image_wind_col_2__11, image_wind_col_2__10, 
         image_wind_col_2__9, image_wind_col_2__8, image_wind_col_2__7, 
         image_wind_col_2__6, image_wind_col_2__5, image_wind_col_2__4, 
         image_wind_col_2__3, image_wind_col_2__2, image_wind_col_2__1, 
         image_wind_col_2__0, image_wind_col_1__15, image_wind_col_1__14, 
         image_wind_col_1__13, image_wind_col_1__12, image_wind_col_1__11, 
         image_wind_col_1__10, image_wind_col_1__9, image_wind_col_1__8, 
         image_wind_col_1__7, image_wind_col_1__6, image_wind_col_1__5, 
         image_wind_col_1__4, image_wind_col_1__3, image_wind_col_1__2, 
         image_wind_col_1__1, image_wind_col_1__0, image_wind_col_0__15, 
         image_wind_col_0__14, image_wind_col_0__13, image_wind_col_0__12, 
         image_wind_col_0__11, image_wind_col_0__10, image_wind_col_0__9, 
         image_wind_col_0__8, image_wind_col_0__7, image_wind_col_0__6, 
         image_wind_col_0__5, image_wind_col_0__4, image_wind_col_0__3, 
         image_wind_col_0__2, image_wind_col_0__1, image_wind_col_0__0, 
         filter_window_ready, filter_window_data_15, filter_window_data_14, 
         filter_window_data_13, filter_window_data_12, filter_window_data_11, 
         filter_window_data_10, filter_window_data_9, filter_window_data_8, 
         filter_window_data_7, filter_window_data_6, filter_window_data_5, 
         filter_window_data_4, filter_window_data_3, filter_window_data_2, 
         filter_window_data_1, filter_window_data_0, comp_unit_ready, 
         comp_unit_operation, comp_unit_relu, comp_unit_flt_size, 
         comp_unit_finished, comp_unit_bias_1_15, comp_unit_bias_1_14, 
         comp_unit_bias_1_13, comp_unit_bias_1_12, comp_unit_bias_1_11, 
         comp_unit_bias_1_10, comp_unit_bias_1_9, comp_unit_bias_1_8, 
         comp_unit_bias_1_7, comp_unit_bias_1_6, comp_unit_bias_1_5, 
         comp_unit_bias_1_4, comp_unit_bias_1_3, comp_unit_bias_1_2, 
         comp_unit_bias_1_1, comp_unit_bias_1_0, comp_unit_bias_2_15, 
         comp_unit_bias_2_14, comp_unit_bias_2_13, comp_unit_bias_2_12, 
         comp_unit_bias_2_11, comp_unit_bias_2_10, comp_unit_bias_2_9, 
         comp_unit_bias_2_8, comp_unit_bias_2_7, comp_unit_bias_2_6, 
         comp_unit_bias_2_5, comp_unit_bias_2_4, comp_unit_bias_2_3, 
         comp_unit_bias_2_2, comp_unit_bias_2_1, comp_unit_bias_2_0, 
         comp_unit_result_1_15, comp_unit_result_1_14, comp_unit_result_1_13, 
         comp_unit_result_1_12, comp_unit_result_1_11, comp_unit_result_1_10, 
         comp_unit_result_1_9, comp_unit_result_1_8, comp_unit_result_1_7, 
         comp_unit_result_1_6, comp_unit_result_1_5, comp_unit_result_1_4, 
         comp_unit_result_1_3, comp_unit_result_1_2, comp_unit_result_1_1, 
         comp_unit_result_1_0, comp_unit_result_2_15, comp_unit_result_2_14, 
         comp_unit_result_2_13, comp_unit_result_2_12, comp_unit_result_2_11, 
         comp_unit_result_2_10, comp_unit_result_2_9, comp_unit_result_2_8, 
         comp_unit_result_2_7, comp_unit_result_2_6, comp_unit_result_2_5, 
         comp_unit_result_2_4, comp_unit_result_2_3, comp_unit_result_2_2, 
         comp_unit_result_2_1, comp_unit_result_2_0, controller_bias_1_15, 
         controller_bias_1_14, controller_bias_1_13, controller_bias_1_12, 
         controller_bias_1_11, controller_bias_1_10, controller_bias_1_9, 
         controller_bias_1_8, controller_bias_1_7, controller_bias_1_6, 
         controller_bias_1_5, controller_bias_1_4, controller_bias_1_3, 
         controller_bias_1_2, controller_bias_1_1, controller_bias_1_0, 
         controller_bias_2_15, controller_bias_2_14, controller_bias_2_13, 
         controller_bias_2_12, controller_bias_2_11, controller_bias_2_10, 
         controller_bias_2_9, controller_bias_2_8, controller_bias_2_7, 
         controller_bias_2_6, controller_bias_2_5, controller_bias_2_4, 
         controller_bias_2_3, controller_bias_2_2, controller_bias_2_1, 
         controller_bias_2_0, controller_result_1_15, controller_result_1_14, 
         controller_result_1_13, controller_result_1_12, controller_result_1_11, 
         controller_result_1_10, controller_result_1_9, controller_result_1_8, 
         controller_result_1_7, controller_result_1_6, controller_result_1_5, 
         controller_result_1_4, controller_result_1_3, controller_result_1_2, 
         controller_result_1_1, controller_result_1_0, controller_result_2_15, 
         controller_result_2_14, controller_result_2_13, controller_result_2_12, 
         controller_result_2_11, controller_result_2_10, controller_result_2_9, 
         controller_result_2_8, controller_result_2_7, controller_result_2_6, 
         controller_result_2_5, controller_result_2_4, controller_result_2_3, 
         controller_result_2_2, controller_result_2_1, controller_result_2_0, 
         argmax_ready, argmax_data_outof_controller_15, 
         argmax_data_outof_controller_14, argmax_data_outof_controller_13, 
         argmax_data_outof_controller_12, argmax_data_outof_controller_11, 
         argmax_data_outof_controller_10, argmax_data_outof_controller_9, 
         argmax_data_outof_controller_8, argmax_data_outof_controller_7, 
         argmax_data_outof_controller_6, argmax_data_outof_controller_5, 
         argmax_data_outof_controller_4, argmax_data_outof_controller_3, 
         argmax_data_outof_controller_2, argmax_data_outof_controller_1, 
         argmax_data_outof_controller_0, argmax_data_out_3, argmax_data_out_2, 
         argmax_data_out_1, argmax_data_out_0, PWR, flt_size_out_0, nx495, nx584, 
         nx594, nx610, nx612, nx614, nx616, nx618, nx620, nx622, nx624, nx626, 
         nx628, nx630, nx632;
    wire [4:0] \$dummy ;




    Controller_16_16_5_16 controller_inst (.clk (clk), .reset (reset), .io_ready_in (
                          io_ready_in), .io_done_out (\$dummy [0]), .mem_data_in (
                          {mem_data_in[15],mem_data_in[14],mem_data_in[13],
                          mem_data_in[12],mem_data_in[11],mem_data_in[10],
                          mem_data_in[9],mem_data_in[8],mem_data_in[7],
                          mem_data_in[6],mem_data_in[5],mem_data_in[4],
                          mem_data_in[3],mem_data_in[2],mem_data_in[1],
                          mem_data_in[0]}), .mem_data_out ({mem_data_out[15],
                          mem_data_out[14],mem_data_out[13],mem_data_out[12],
                          mem_data_out[11],mem_data_out[10],mem_data_out[9],
                          mem_data_out[8],mem_data_out[7],mem_data_out[6],
                          mem_data_out[5],mem_data_out[4],mem_data_out[3],
                          mem_data_out[2],mem_data_out[1],mem_data_out[0]}), .mem_addr_out (
                          {mem_addr_out[15],mem_addr_out[14],mem_addr_out[13],
                          mem_addr_out[12],mem_addr_out[11],mem_addr_out[10],
                          mem_addr_out[9],mem_addr_out[8],mem_addr_out[7],
                          mem_addr_out[6],mem_addr_out[5],mem_addr_out[4],
                          mem_addr_out[3],mem_addr_out[2],mem_addr_out[1],
                          mem_addr_out[0]}), .mem_write_out (mem_write_out), .mem_read_out (
                          mem_read_out), .wind_en (image_wind_en), .wind_rst (
                          \$dummy [1]), .wind_col_in_4__15 (image_wind_col_4__15
                          ), .wind_col_in_4__14 (image_wind_col_4__14), .wind_col_in_4__13 (
                          image_wind_col_4__13), .wind_col_in_4__12 (
                          image_wind_col_4__12), .wind_col_in_4__11 (
                          image_wind_col_4__11), .wind_col_in_4__10 (
                          image_wind_col_4__10), .wind_col_in_4__9 (
                          image_wind_col_4__9), .wind_col_in_4__8 (
                          image_wind_col_4__8), .wind_col_in_4__7 (
                          image_wind_col_4__7), .wind_col_in_4__6 (
                          image_wind_col_4__6), .wind_col_in_4__5 (
                          image_wind_col_4__5), .wind_col_in_4__4 (
                          image_wind_col_4__4), .wind_col_in_4__3 (
                          image_wind_col_4__3), .wind_col_in_4__2 (
                          image_wind_col_4__2), .wind_col_in_4__1 (
                          image_wind_col_4__1), .wind_col_in_4__0 (
                          image_wind_col_4__0), .wind_col_in_3__15 (
                          image_wind_col_3__15), .wind_col_in_3__14 (
                          image_wind_col_3__14), .wind_col_in_3__13 (
                          image_wind_col_3__13), .wind_col_in_3__12 (
                          image_wind_col_3__12), .wind_col_in_3__11 (
                          image_wind_col_3__11), .wind_col_in_3__10 (
                          image_wind_col_3__10), .wind_col_in_3__9 (
                          image_wind_col_3__9), .wind_col_in_3__8 (
                          image_wind_col_3__8), .wind_col_in_3__7 (
                          image_wind_col_3__7), .wind_col_in_3__6 (
                          image_wind_col_3__6), .wind_col_in_3__5 (
                          image_wind_col_3__5), .wind_col_in_3__4 (
                          image_wind_col_3__4), .wind_col_in_3__3 (
                          image_wind_col_3__3), .wind_col_in_3__2 (
                          image_wind_col_3__2), .wind_col_in_3__1 (
                          image_wind_col_3__1), .wind_col_in_3__0 (
                          image_wind_col_3__0), .wind_col_in_2__15 (
                          image_wind_col_2__15), .wind_col_in_2__14 (
                          image_wind_col_2__14), .wind_col_in_2__13 (
                          image_wind_col_2__13), .wind_col_in_2__12 (
                          image_wind_col_2__12), .wind_col_in_2__11 (
                          image_wind_col_2__11), .wind_col_in_2__10 (
                          image_wind_col_2__10), .wind_col_in_2__9 (
                          image_wind_col_2__9), .wind_col_in_2__8 (
                          image_wind_col_2__8), .wind_col_in_2__7 (
                          image_wind_col_2__7), .wind_col_in_2__6 (
                          image_wind_col_2__6), .wind_col_in_2__5 (
                          image_wind_col_2__5), .wind_col_in_2__4 (
                          image_wind_col_2__4), .wind_col_in_2__3 (
                          image_wind_col_2__3), .wind_col_in_2__2 (
                          image_wind_col_2__2), .wind_col_in_2__1 (
                          image_wind_col_2__1), .wind_col_in_2__0 (
                          image_wind_col_2__0), .wind_col_in_1__15 (
                          image_wind_col_1__15), .wind_col_in_1__14 (
                          image_wind_col_1__14), .wind_col_in_1__13 (
                          image_wind_col_1__13), .wind_col_in_1__12 (
                          image_wind_col_1__12), .wind_col_in_1__11 (
                          image_wind_col_1__11), .wind_col_in_1__10 (
                          image_wind_col_1__10), .wind_col_in_1__9 (
                          image_wind_col_1__9), .wind_col_in_1__8 (
                          image_wind_col_1__8), .wind_col_in_1__7 (
                          image_wind_col_1__7), .wind_col_in_1__6 (
                          image_wind_col_1__6), .wind_col_in_1__5 (
                          image_wind_col_1__5), .wind_col_in_1__4 (
                          image_wind_col_1__4), .wind_col_in_1__3 (
                          image_wind_col_1__3), .wind_col_in_1__2 (
                          image_wind_col_1__2), .wind_col_in_1__1 (
                          image_wind_col_1__1), .wind_col_in_1__0 (
                          image_wind_col_1__0), .wind_col_in_0__15 (
                          image_wind_col_0__15), .wind_col_in_0__14 (
                          image_wind_col_0__14), .wind_col_in_0__13 (
                          image_wind_col_0__13), .wind_col_in_0__12 (
                          image_wind_col_0__12), .wind_col_in_0__11 (
                          image_wind_col_0__11), .wind_col_in_0__10 (
                          image_wind_col_0__10), .wind_col_in_0__9 (
                          image_wind_col_0__9), .wind_col_in_0__8 (
                          image_wind_col_0__8), .wind_col_in_0__7 (
                          image_wind_col_0__7), .wind_col_in_0__6 (
                          image_wind_col_0__6), .wind_col_in_0__5 (
                          image_wind_col_0__5), .wind_col_in_0__4 (
                          image_wind_col_0__4), .wind_col_in_0__3 (
                          image_wind_col_0__3), .wind_col_in_0__2 (
                          image_wind_col_0__2), .wind_col_in_0__1 (
                          image_wind_col_0__1), .wind_col_in_0__0 (
                          image_wind_col_0__0), .filter_data_out ({
                          filter_window_data_15,filter_window_data_14,
                          filter_window_data_13,filter_window_data_12,
                          filter_window_data_11,filter_window_data_10,
                          filter_window_data_9,filter_window_data_8,
                          filter_window_data_7,filter_window_data_6,
                          filter_window_data_5,filter_window_data_4,
                          filter_window_data_3,filter_window_data_2,
                          filter_window_data_1,filter_window_data_0}), .filter_ready_out (
                          filter_window_ready), .filter_reset (\$dummy [2]), .comp_unit_ready (
                          comp_unit_ready), .comp_unit_operation (
                          comp_unit_operation), .comp_unit_flt_size (
                          comp_unit_flt_size), .comp_unit_relu (comp_unit_relu)
                          , .comp_unit_data1_out ({controller_bias_1_15,
                          controller_bias_1_14,controller_bias_1_13,
                          controller_bias_1_12,controller_bias_1_11,
                          controller_bias_1_10,controller_bias_1_9,
                          controller_bias_1_8,controller_bias_1_7,
                          controller_bias_1_6,controller_bias_1_5,
                          controller_bias_1_4,controller_bias_1_3,
                          controller_bias_1_2,controller_bias_1_1,
                          controller_bias_1_0}), .comp_unit_data2_out ({
                          controller_bias_2_15,controller_bias_2_14,
                          controller_bias_2_13,controller_bias_2_12,
                          controller_bias_2_11,controller_bias_2_10,
                          controller_bias_2_9,controller_bias_2_8,
                          controller_bias_2_7,controller_bias_2_6,
                          controller_bias_2_5,controller_bias_2_4,
                          controller_bias_2_3,controller_bias_2_2,
                          controller_bias_2_1,controller_bias_2_0}), .comp_unit_buffer_finished (
                          io_done_out), .comp_unit_finished (comp_unit_finished)
                          , .comp_unit_data1_in ({controller_result_1_15,
                          controller_result_1_14,controller_result_1_13,
                          controller_result_1_12,controller_result_1_11,
                          controller_result_1_10,controller_result_1_9,
                          controller_result_1_8,controller_result_1_7,
                          controller_result_1_6,controller_result_1_5,
                          controller_result_1_4,controller_result_1_3,
                          controller_result_1_2,controller_result_1_1,
                          controller_result_1_0}), .comp_unit_data2_in ({
                          controller_result_2_15,controller_result_2_14,
                          controller_result_2_13,controller_result_2_12,
                          controller_result_2_11,controller_result_2_10,
                          controller_result_2_9,controller_result_2_8,
                          controller_result_2_7,controller_result_2_6,
                          controller_result_2_5,controller_result_2_4,
                          controller_result_2_3,controller_result_2_2,
                          controller_result_2_1,controller_result_2_0}), .argmax_ready (
                          argmax_ready), .argmax_data_out ({
                          argmax_data_outof_controller_15,
                          argmax_data_outof_controller_14,
                          argmax_data_outof_controller_13,
                          argmax_data_outof_controller_12,
                          argmax_data_outof_controller_11,
                          argmax_data_outof_controller_10,
                          argmax_data_outof_controller_9,
                          argmax_data_outof_controller_8,
                          argmax_data_outof_controller_7,
                          argmax_data_outof_controller_6,
                          argmax_data_outof_controller_5,
                          argmax_data_outof_controller_4,
                          argmax_data_outof_controller_3,
                          argmax_data_outof_controller_2,
                          argmax_data_outof_controller_1,
                          argmax_data_outof_controller_0}), .argmax_data_in ({
                          io_done_out,io_done_out,io_done_out,io_done_out,
                          io_done_out,io_done_out,io_done_out,io_done_out,
                          io_done_out,io_done_out,io_done_out,io_done_out,
                          argmax_data_out_3,argmax_data_out_2,argmax_data_out_1,
                          argmax_data_out_0})) ;
    ComputationBlock computation_block_inst (.img_data_col_0 ({
                     image_wind_col_0__15,image_wind_col_0__14,
                     image_wind_col_0__13,image_wind_col_0__12,
                     image_wind_col_0__11,image_wind_col_0__10,
                     image_wind_col_0__9,image_wind_col_0__8,image_wind_col_0__7
                     ,image_wind_col_0__6,image_wind_col_0__5,
                     image_wind_col_0__4,image_wind_col_0__3,image_wind_col_0__2
                     ,image_wind_col_0__1,image_wind_col_0__0}), .img_data_col_1 (
                     {image_wind_col_1__15,image_wind_col_1__14,
                     image_wind_col_1__13,image_wind_col_1__12,
                     image_wind_col_1__11,image_wind_col_1__10,
                     image_wind_col_1__9,image_wind_col_1__8,image_wind_col_1__7
                     ,image_wind_col_1__6,image_wind_col_1__5,
                     image_wind_col_1__4,image_wind_col_1__3,image_wind_col_1__2
                     ,image_wind_col_1__1,image_wind_col_1__0}), .img_data_col_2 (
                     {image_wind_col_2__15,image_wind_col_2__14,
                     image_wind_col_2__13,image_wind_col_2__12,
                     image_wind_col_2__11,image_wind_col_2__10,
                     image_wind_col_2__9,image_wind_col_2__8,image_wind_col_2__7
                     ,image_wind_col_2__6,image_wind_col_2__5,
                     image_wind_col_2__4,image_wind_col_2__3,image_wind_col_2__2
                     ,image_wind_col_2__1,image_wind_col_2__0}), .img_data_col_3 (
                     {image_wind_col_3__15,image_wind_col_3__14,
                     image_wind_col_3__13,image_wind_col_3__12,
                     image_wind_col_3__11,image_wind_col_3__10,
                     image_wind_col_3__9,image_wind_col_3__8,image_wind_col_3__7
                     ,image_wind_col_3__6,image_wind_col_3__5,
                     image_wind_col_3__4,image_wind_col_3__3,image_wind_col_3__2
                     ,image_wind_col_3__1,image_wind_col_3__0}), .img_data_col_4 (
                     {image_wind_col_4__15,image_wind_col_4__14,
                     image_wind_col_4__13,image_wind_col_4__12,
                     image_wind_col_4__11,image_wind_col_4__10,
                     image_wind_col_4__9,image_wind_col_4__8,image_wind_col_4__7
                     ,image_wind_col_4__6,image_wind_col_4__5,
                     image_wind_col_4__4,image_wind_col_4__3,image_wind_col_4__2
                     ,image_wind_col_4__1,image_wind_col_4__0}), .img_load (
                     image_wind_en), .img_reset (io_done_out), .filter_data_word (
                     {filter_window_data_15,filter_window_data_14,
                     filter_window_data_13,filter_window_data_12,
                     filter_window_data_11,filter_window_data_10,
                     filter_window_data_9,filter_window_data_8,
                     filter_window_data_7,filter_window_data_6,
                     filter_window_data_5,filter_window_data_4,
                     filter_window_data_3,filter_window_data_2,
                     filter_window_data_1,filter_window_data_0}), .filter_load (
                     filter_window_ready), .filter_reset (reset), .start (
                     comp_unit_ready), .operation (comp_unit_operation), .compute_relu (
                     comp_unit_relu), .filter_size (comp_unit_flt_size), .output1_init (
                     {comp_unit_bias_1_15,comp_unit_bias_1_14,
                     comp_unit_bias_1_13,comp_unit_bias_1_12,comp_unit_bias_1_11
                     ,comp_unit_bias_1_10,comp_unit_bias_1_9,comp_unit_bias_1_8,
                     comp_unit_bias_1_7,comp_unit_bias_1_6,comp_unit_bias_1_5,
                     comp_unit_bias_1_4,comp_unit_bias_1_3,comp_unit_bias_1_2,
                     comp_unit_bias_1_1,comp_unit_bias_1_0}), .output2_init ({
                     comp_unit_bias_2_15,comp_unit_bias_2_14,comp_unit_bias_2_13
                     ,comp_unit_bias_2_12,comp_unit_bias_2_11,
                     comp_unit_bias_2_10,comp_unit_bias_2_9,comp_unit_bias_2_8,
                     comp_unit_bias_2_7,comp_unit_bias_2_6,comp_unit_bias_2_5,
                     comp_unit_bias_2_4,comp_unit_bias_2_3,comp_unit_bias_2_2,
                     comp_unit_bias_2_1,comp_unit_bias_2_0}), .output1 ({
                     comp_unit_result_1_15,comp_unit_result_1_14,
                     comp_unit_result_1_13,comp_unit_result_1_12,
                     comp_unit_result_1_11,comp_unit_result_1_10,
                     comp_unit_result_1_9,comp_unit_result_1_8,
                     comp_unit_result_1_7,comp_unit_result_1_6,
                     comp_unit_result_1_5,comp_unit_result_1_4,
                     comp_unit_result_1_3,comp_unit_result_1_2,
                     comp_unit_result_1_1,comp_unit_result_1_0}), .output2 ({
                     comp_unit_result_2_15,comp_unit_result_2_14,
                     comp_unit_result_2_13,comp_unit_result_2_12,
                     comp_unit_result_2_11,comp_unit_result_2_10,
                     comp_unit_result_2_9,comp_unit_result_2_8,
                     comp_unit_result_2_7,comp_unit_result_2_6,
                     comp_unit_result_2_5,comp_unit_result_2_4,
                     comp_unit_result_2_3,comp_unit_result_2_2,
                     comp_unit_result_2_1,comp_unit_result_2_0}), .buffer_ready (
                     \$dummy [3]), .ready (comp_unit_finished), .clk (clk), .en (
                     PWR), .reset (io_done_out)) ;
    ArgMax argmax_inst (.inp ({argmax_data_outof_controller_15,
           argmax_data_outof_controller_14,argmax_data_outof_controller_13,
           argmax_data_outof_controller_12,argmax_data_outof_controller_11,
           argmax_data_outof_controller_10,argmax_data_outof_controller_9,
           argmax_data_outof_controller_8,argmax_data_outof_controller_7,
           argmax_data_outof_controller_6,argmax_data_outof_controller_5,
           argmax_data_outof_controller_4,argmax_data_outof_controller_3,
           argmax_data_outof_controller_2,argmax_data_outof_controller_1,
           argmax_data_outof_controller_0}), .en (argmax_ready), .clk (clk), .rst (
           reset), .ans ({argmax_data_out_3,argmax_data_out_2,argmax_data_out_1,
           argmax_data_out_0})) ;
    fake_vcc ix415 (.Y (PWR)) ;
    fake_gnd ix413 (.Y (io_done_out)) ;
    dffr flt_size_reg_reg_q_0 (.Q (flt_size_out_0), .QB (\$dummy [4]), .D (nx495
         ), .CLK (clk), .R (reset)) ;
    mux21_ni ix496 (.Y (nx495), .A0 (nx584), .A1 (comp_unit_flt_size), .S0 (
             comp_unit_ready)) ;
    inv02 ix583 (.Y (nx584), .A (nx612)) ;
    mux21_ni ix11 (.Y (controller_result_2_0), .A0 (comp_unit_result_1_0), .A1 (
             comp_unit_result_2_0), .S0 (nx612)) ;
    mux21_ni ix19 (.Y (controller_result_2_1), .A0 (comp_unit_result_1_1), .A1 (
             comp_unit_result_2_1), .S0 (nx612)) ;
    mux21_ni ix27 (.Y (controller_result_2_2), .A0 (comp_unit_result_1_2), .A1 (
             comp_unit_result_2_2), .S0 (nx612)) ;
    mux21_ni ix35 (.Y (controller_result_2_3), .A0 (comp_unit_result_1_3), .A1 (
             comp_unit_result_2_3), .S0 (nx612)) ;
    mux21_ni ix43 (.Y (controller_result_2_4), .A0 (comp_unit_result_1_4), .A1 (
             comp_unit_result_2_4), .S0 (nx612)) ;
    mux21_ni ix51 (.Y (controller_result_2_5), .A0 (comp_unit_result_1_5), .A1 (
             comp_unit_result_2_5), .S0 (nx612)) ;
    mux21_ni ix59 (.Y (controller_result_2_6), .A0 (comp_unit_result_1_6), .A1 (
             comp_unit_result_2_6), .S0 (nx614)) ;
    mux21_ni ix67 (.Y (controller_result_2_7), .A0 (comp_unit_result_1_7), .A1 (
             comp_unit_result_2_7), .S0 (nx614)) ;
    mux21_ni ix75 (.Y (controller_result_2_8), .A0 (comp_unit_result_1_8), .A1 (
             comp_unit_result_2_8), .S0 (nx614)) ;
    mux21_ni ix83 (.Y (controller_result_2_9), .A0 (comp_unit_result_1_9), .A1 (
             comp_unit_result_2_9), .S0 (nx614)) ;
    mux21_ni ix91 (.Y (controller_result_2_10), .A0 (comp_unit_result_1_10), .A1 (
             comp_unit_result_2_10), .S0 (nx614)) ;
    mux21_ni ix99 (.Y (controller_result_2_11), .A0 (comp_unit_result_1_11), .A1 (
             comp_unit_result_2_11), .S0 (nx614)) ;
    mux21_ni ix107 (.Y (controller_result_2_12), .A0 (comp_unit_result_1_12), .A1 (
             comp_unit_result_2_12), .S0 (nx614)) ;
    mux21_ni ix115 (.Y (controller_result_2_13), .A0 (comp_unit_result_1_13), .A1 (
             comp_unit_result_2_13), .S0 (nx616)) ;
    mux21_ni ix123 (.Y (controller_result_2_14), .A0 (comp_unit_result_1_14), .A1 (
             comp_unit_result_2_14), .S0 (nx616)) ;
    mux21_ni ix131 (.Y (controller_result_2_15), .A0 (comp_unit_result_1_15), .A1 (
             comp_unit_result_2_15), .S0 (nx616)) ;
    mux21_ni ix139 (.Y (controller_result_1_0), .A0 (comp_unit_result_2_0), .A1 (
             comp_unit_result_1_0), .S0 (nx616)) ;
    mux21_ni ix147 (.Y (controller_result_1_1), .A0 (comp_unit_result_2_1), .A1 (
             comp_unit_result_1_1), .S0 (nx616)) ;
    mux21_ni ix155 (.Y (controller_result_1_2), .A0 (comp_unit_result_2_2), .A1 (
             comp_unit_result_1_2), .S0 (nx616)) ;
    mux21_ni ix163 (.Y (controller_result_1_3), .A0 (comp_unit_result_2_3), .A1 (
             comp_unit_result_1_3), .S0 (nx616)) ;
    mux21_ni ix171 (.Y (controller_result_1_4), .A0 (comp_unit_result_2_4), .A1 (
             comp_unit_result_1_4), .S0 (nx618)) ;
    mux21_ni ix179 (.Y (controller_result_1_5), .A0 (comp_unit_result_2_5), .A1 (
             comp_unit_result_1_5), .S0 (nx618)) ;
    mux21_ni ix187 (.Y (controller_result_1_6), .A0 (comp_unit_result_2_6), .A1 (
             comp_unit_result_1_6), .S0 (nx618)) ;
    mux21_ni ix195 (.Y (controller_result_1_7), .A0 (comp_unit_result_2_7), .A1 (
             comp_unit_result_1_7), .S0 (nx618)) ;
    mux21_ni ix203 (.Y (controller_result_1_8), .A0 (comp_unit_result_2_8), .A1 (
             comp_unit_result_1_8), .S0 (nx618)) ;
    mux21_ni ix211 (.Y (controller_result_1_9), .A0 (comp_unit_result_2_9), .A1 (
             comp_unit_result_1_9), .S0 (nx618)) ;
    mux21_ni ix219 (.Y (controller_result_1_10), .A0 (comp_unit_result_2_10), .A1 (
             comp_unit_result_1_10), .S0 (nx618)) ;
    mux21_ni ix227 (.Y (controller_result_1_11), .A0 (comp_unit_result_2_11), .A1 (
             comp_unit_result_1_11), .S0 (nx620)) ;
    mux21_ni ix235 (.Y (controller_result_1_12), .A0 (comp_unit_result_2_12), .A1 (
             comp_unit_result_1_12), .S0 (nx620)) ;
    mux21_ni ix243 (.Y (controller_result_1_13), .A0 (comp_unit_result_2_13), .A1 (
             comp_unit_result_1_13), .S0 (nx620)) ;
    mux21_ni ix251 (.Y (controller_result_1_14), .A0 (comp_unit_result_2_14), .A1 (
             comp_unit_result_1_14), .S0 (nx620)) ;
    mux21_ni ix259 (.Y (controller_result_1_15), .A0 (comp_unit_result_2_15), .A1 (
             comp_unit_result_1_15), .S0 (nx620)) ;
    mux21_ni ix269 (.Y (comp_unit_bias_2_0), .A0 (controller_bias_2_0), .A1 (
             controller_bias_1_0), .S0 (nx624)) ;
    nand02 ix545 (.Y (nx594), .A0 (nx620), .A1 (nx610)) ;
    inv01 ix609 (.Y (nx610), .A (comp_unit_flt_size)) ;
    mux21_ni ix277 (.Y (comp_unit_bias_2_1), .A0 (controller_bias_2_1), .A1 (
             controller_bias_1_1), .S0 (nx624)) ;
    mux21_ni ix285 (.Y (comp_unit_bias_2_2), .A0 (controller_bias_2_2), .A1 (
             controller_bias_1_2), .S0 (nx624)) ;
    mux21_ni ix293 (.Y (comp_unit_bias_2_3), .A0 (controller_bias_2_3), .A1 (
             controller_bias_1_3), .S0 (nx624)) ;
    mux21_ni ix301 (.Y (comp_unit_bias_2_4), .A0 (controller_bias_2_4), .A1 (
             controller_bias_1_4), .S0 (nx624)) ;
    mux21_ni ix309 (.Y (comp_unit_bias_2_5), .A0 (controller_bias_2_5), .A1 (
             controller_bias_1_5), .S0 (nx624)) ;
    mux21_ni ix317 (.Y (comp_unit_bias_2_6), .A0 (controller_bias_2_6), .A1 (
             controller_bias_1_6), .S0 (nx624)) ;
    mux21_ni ix325 (.Y (comp_unit_bias_2_7), .A0 (controller_bias_2_7), .A1 (
             controller_bias_1_7), .S0 (nx626)) ;
    mux21_ni ix333 (.Y (comp_unit_bias_2_8), .A0 (controller_bias_2_8), .A1 (
             controller_bias_1_8), .S0 (nx626)) ;
    mux21_ni ix341 (.Y (comp_unit_bias_2_9), .A0 (controller_bias_2_9), .A1 (
             controller_bias_1_9), .S0 (nx626)) ;
    mux21_ni ix349 (.Y (comp_unit_bias_2_10), .A0 (controller_bias_2_10), .A1 (
             controller_bias_1_10), .S0 (nx626)) ;
    mux21_ni ix357 (.Y (comp_unit_bias_2_11), .A0 (controller_bias_2_11), .A1 (
             controller_bias_1_11), .S0 (nx626)) ;
    mux21_ni ix365 (.Y (comp_unit_bias_2_12), .A0 (controller_bias_2_12), .A1 (
             controller_bias_1_12), .S0 (nx626)) ;
    mux21_ni ix373 (.Y (comp_unit_bias_2_13), .A0 (controller_bias_2_13), .A1 (
             controller_bias_1_13), .S0 (nx626)) ;
    mux21_ni ix381 (.Y (comp_unit_bias_2_14), .A0 (controller_bias_2_14), .A1 (
             controller_bias_1_14), .S0 (nx628)) ;
    mux21_ni ix389 (.Y (comp_unit_bias_2_15), .A0 (controller_bias_2_15), .A1 (
             controller_bias_1_15), .S0 (nx628)) ;
    mux21_ni ix397 (.Y (comp_unit_bias_1_0), .A0 (controller_bias_1_0), .A1 (
             controller_bias_2_0), .S0 (nx628)) ;
    mux21_ni ix405 (.Y (comp_unit_bias_1_1), .A0 (controller_bias_1_1), .A1 (
             controller_bias_2_1), .S0 (nx628)) ;
    mux21_ni ix417 (.Y (comp_unit_bias_1_2), .A0 (controller_bias_1_2), .A1 (
             controller_bias_2_2), .S0 (nx628)) ;
    mux21_ni ix421 (.Y (comp_unit_bias_1_3), .A0 (controller_bias_1_3), .A1 (
             controller_bias_2_3), .S0 (nx628)) ;
    mux21_ni ix429 (.Y (comp_unit_bias_1_4), .A0 (controller_bias_1_4), .A1 (
             controller_bias_2_4), .S0 (nx628)) ;
    mux21_ni ix437 (.Y (comp_unit_bias_1_5), .A0 (controller_bias_1_5), .A1 (
             controller_bias_2_5), .S0 (nx630)) ;
    mux21_ni ix445 (.Y (comp_unit_bias_1_6), .A0 (controller_bias_1_6), .A1 (
             controller_bias_2_6), .S0 (nx630)) ;
    mux21_ni ix453 (.Y (comp_unit_bias_1_7), .A0 (controller_bias_1_7), .A1 (
             controller_bias_2_7), .S0 (nx630)) ;
    mux21_ni ix461 (.Y (comp_unit_bias_1_8), .A0 (controller_bias_1_8), .A1 (
             controller_bias_2_8), .S0 (nx630)) ;
    mux21_ni ix469 (.Y (comp_unit_bias_1_9), .A0 (controller_bias_1_9), .A1 (
             controller_bias_2_9), .S0 (nx630)) ;
    mux21_ni ix477 (.Y (comp_unit_bias_1_10), .A0 (controller_bias_1_10), .A1 (
             controller_bias_2_10), .S0 (nx630)) ;
    mux21_ni ix485 (.Y (comp_unit_bias_1_11), .A0 (controller_bias_1_11), .A1 (
             controller_bias_2_11), .S0 (nx630)) ;
    mux21_ni ix493 (.Y (comp_unit_bias_1_12), .A0 (controller_bias_1_12), .A1 (
             controller_bias_2_12), .S0 (nx632)) ;
    mux21_ni ix501 (.Y (comp_unit_bias_1_13), .A0 (controller_bias_1_13), .A1 (
             controller_bias_2_13), .S0 (nx632)) ;
    mux21_ni ix509 (.Y (comp_unit_bias_1_14), .A0 (controller_bias_1_14), .A1 (
             controller_bias_2_14), .S0 (nx632)) ;
    mux21_ni ix517 (.Y (comp_unit_bias_1_15), .A0 (controller_bias_1_15), .A1 (
             controller_bias_2_15), .S0 (nx632)) ;
    inv02 ix611 (.Y (nx612), .A (flt_size_out_0)) ;
    inv02 ix613 (.Y (nx614), .A (flt_size_out_0)) ;
    inv02 ix615 (.Y (nx616), .A (flt_size_out_0)) ;
    inv02 ix617 (.Y (nx618), .A (flt_size_out_0)) ;
    inv02 ix619 (.Y (nx620), .A (flt_size_out_0)) ;
    inv01 ix621 (.Y (nx622), .A (nx594)) ;
    inv02 ix623 (.Y (nx624), .A (nx622)) ;
    inv02 ix625 (.Y (nx626), .A (nx622)) ;
    inv02 ix627 (.Y (nx628), .A (nx622)) ;
    inv02 ix629 (.Y (nx630), .A (nx622)) ;
    inv02 ix631 (.Y (nx632), .A (nx622)) ;
endmodule


module ArgMax ( inp, en, clk, rst, ans ) ;

    input [15:0]inp ;
    input en ;
    input clk ;
    input rst ;
    output [3:0]ans ;

    wire reg_val_out_15, reg_val_out_14, reg_val_out_13, reg_val_out_12, 
         reg_val_out_11, reg_val_out_10, reg_val_out_9, reg_val_out_8, 
         reg_val_out_7, reg_val_out_6, reg_val_out_5, reg_val_out_4, 
         reg_val_out_3, reg_val_out_2, reg_val_out_1, reg_val_out_0, 
         compare_in1_inverted_15, compare_in1_inverted_14, 
         compare_in1_inverted_13, compare_in1_inverted_12, 
         compare_in1_inverted_11, compare_in1_inverted_10, 
         compare_in1_inverted_9, compare_in1_inverted_8, compare_in1_inverted_7, 
         compare_in1_inverted_6, compare_in1_inverted_5, compare_in1_inverted_4, 
         compare_in1_inverted_3, compare_in1_inverted_2, compare_in1_inverted_1, 
         compare_in1_inverted_0, compare_sub_res_15, tmp_15, curr_idx_0, nx54, 
         reg_idx_out_0, curr_idx_1, reg_idx_out_1, curr_idx_2, nx98, 
         reg_idx_out_2, curr_idx_3, nx157, reg_idx_out_3, nx140, nx152, nx164, 
         nx176, nx188, nx200, nx212, nx224, nx236, nx248, nx260, nx272, nx284, 
         nx296, nx308, nx165, nx175, nx185, nx195, nx205, nx215, nx225, nx235, 
         nx245, nx255, nx265, nx275, nx285, nx295, nx305, nx315, nx325, nx335, 
         nx345, nx355, nx365, nx375, nx385, nx395, nx405, nx411, nx482, nx484, 
         nx486, nx503, nx556, nx558, nx560, nx562, nx564, nx566, nx568, nx570;
    wire [37:0] \$dummy ;




    NAdder_16 compare_DoSubtraction (.a ({reg_val_out_15,reg_val_out_14,
              reg_val_out_13,reg_val_out_12,reg_val_out_11,reg_val_out_10,
              reg_val_out_9,reg_val_out_8,reg_val_out_7,reg_val_out_6,
              reg_val_out_5,reg_val_out_4,reg_val_out_3,reg_val_out_2,
              reg_val_out_1,reg_val_out_0}), .b ({compare_in1_inverted_15,
              compare_in1_inverted_14,compare_in1_inverted_13,
              compare_in1_inverted_12,compare_in1_inverted_11,
              compare_in1_inverted_10,compare_in1_inverted_9,
              compare_in1_inverted_8,compare_in1_inverted_7,
              compare_in1_inverted_6,compare_in1_inverted_5,
              compare_in1_inverted_4,compare_in1_inverted_3,
              compare_in1_inverted_2,compare_in1_inverted_1,
              compare_in1_inverted_0}), .cin (tmp_15), .s ({compare_sub_res_15,
              \$dummy [0],\$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],
              \$dummy [5],\$dummy [6],\$dummy [7],\$dummy [8],\$dummy [9],
              \$dummy [10],\$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14]})
              , .cout (\$dummy [15])) ;
    fake_vcc ix115 (.Y (tmp_15)) ;
    dffr valReg_reg_q_0 (.Q (reg_val_out_0), .QB (\$dummy [16]), .D (nx255), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix256 (.Y (nx255), .A0 (reg_val_out_0), .A1 (nx140), .S0 (nx558)) ;
    oai22 ix55 (.Y (nx54), .A0 (compare_sub_res_15), .A1 (nx405), .B0 (
          compare_in1_inverted_15), .B1 (reg_val_out_15)) ;
    aoi21 ix176 (.Y (nx175), .A0 (nx558), .A1 (compare_in1_inverted_15), .B0 (
          nx411)) ;
    inv01 ix410 (.Y (compare_in1_inverted_15), .A (inp[15])) ;
    dffs_ni valReg_reg_q_15 (.Q (reg_val_out_15), .QB (nx411), .D (nx175), .CLK (
            clk), .S (rst)) ;
    dffr valReg_reg_q_1 (.Q (reg_val_out_1), .QB (\$dummy [17]), .D (nx265), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix266 (.Y (nx265), .A0 (reg_val_out_1), .A1 (nx152), .S0 (nx558)) ;
    dffr valReg_reg_q_2 (.Q (reg_val_out_2), .QB (\$dummy [18]), .D (nx275), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix276 (.Y (nx275), .A0 (reg_val_out_2), .A1 (nx164), .S0 (nx558)) ;
    dffr valReg_reg_q_3 (.Q (reg_val_out_3), .QB (\$dummy [19]), .D (nx285), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix286 (.Y (nx285), .A0 (reg_val_out_3), .A1 (nx176), .S0 (nx558)) ;
    dffr valReg_reg_q_4 (.Q (reg_val_out_4), .QB (\$dummy [20]), .D (nx295), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix296 (.Y (nx295), .A0 (reg_val_out_4), .A1 (nx188), .S0 (nx558)) ;
    dffr valReg_reg_q_5 (.Q (reg_val_out_5), .QB (\$dummy [21]), .D (nx305), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix306 (.Y (nx305), .A0 (reg_val_out_5), .A1 (nx200), .S0 (nx558)) ;
    dffr valReg_reg_q_6 (.Q (reg_val_out_6), .QB (\$dummy [22]), .D (nx315), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix316 (.Y (nx315), .A0 (reg_val_out_6), .A1 (nx212), .S0 (nx560)) ;
    dffr valReg_reg_q_7 (.Q (reg_val_out_7), .QB (\$dummy [23]), .D (nx325), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix326 (.Y (nx325), .A0 (reg_val_out_7), .A1 (nx224), .S0 (nx560)) ;
    dffr valReg_reg_q_8 (.Q (reg_val_out_8), .QB (\$dummy [24]), .D (nx335), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix336 (.Y (nx335), .A0 (reg_val_out_8), .A1 (nx236), .S0 (nx560)) ;
    dffr valReg_reg_q_9 (.Q (reg_val_out_9), .QB (\$dummy [25]), .D (nx345), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix346 (.Y (nx345), .A0 (reg_val_out_9), .A1 (nx248), .S0 (nx560)) ;
    dffr valReg_reg_q_10 (.Q (reg_val_out_10), .QB (\$dummy [26]), .D (nx355), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix356 (.Y (nx355), .A0 (reg_val_out_10), .A1 (nx260), .S0 (nx560)
             ) ;
    dffr valReg_reg_q_11 (.Q (reg_val_out_11), .QB (\$dummy [27]), .D (nx365), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix366 (.Y (nx365), .A0 (reg_val_out_11), .A1 (nx272), .S0 (nx560)
             ) ;
    dffr valReg_reg_q_12 (.Q (reg_val_out_12), .QB (\$dummy [28]), .D (nx375), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix376 (.Y (nx375), .A0 (reg_val_out_12), .A1 (nx284), .S0 (nx560)
             ) ;
    dffr valReg_reg_q_13 (.Q (reg_val_out_13), .QB (\$dummy [29]), .D (nx385), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix386 (.Y (nx385), .A0 (reg_val_out_13), .A1 (nx296), .S0 (nx562)
             ) ;
    dffr valReg_reg_q_14 (.Q (reg_val_out_14), .QB (\$dummy [30]), .D (nx395), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix396 (.Y (nx395), .A0 (reg_val_out_14), .A1 (nx308), .S0 (nx562)
             ) ;
    dffr reg_curr_idx_0 (.Q (curr_idx_0), .QB (\$dummy [31]), .D (nx165), .CLK (
         clk), .R (rst)) ;
    dffr idxReg_reg_q_0 (.Q (reg_idx_out_0), .QB (\$dummy [32]), .D (nx185), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix186 (.Y (nx185), .A0 (reg_idx_out_0), .A1 (ans[0]), .S0 (nx562)
             ) ;
    mux21 ix196 (.Y (nx195), .A0 (nx482), .A1 (nx484), .S0 (nx562)) ;
    dffr reg_curr_idx_1 (.Q (curr_idx_1), .QB (nx482), .D (nx195), .CLK (clk), .R (
         rst)) ;
    oai21 ix485 (.Y (nx484), .A0 (curr_idx_0), .A1 (curr_idx_1), .B0 (nx486)) ;
    nand02 ix487 (.Y (nx486), .A0 (curr_idx_1), .A1 (curr_idx_0)) ;
    dffr idxReg_reg_q_1 (.Q (reg_idx_out_1), .QB (\$dummy [33]), .D (nx205), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix206 (.Y (nx205), .A0 (reg_idx_out_1), .A1 (ans[1]), .S0 (nx562)
             ) ;
    dffr reg_curr_idx_2 (.Q (curr_idx_2), .QB (\$dummy [34]), .D (nx215), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix216 (.Y (nx215), .A0 (curr_idx_2), .A1 (nx98), .S0 (nx562)) ;
    xnor2 ix99 (.Y (nx98), .A0 (curr_idx_2), .A1 (nx486)) ;
    dffr idxReg_reg_q_2 (.Q (reg_idx_out_2), .QB (\$dummy [35]), .D (nx225), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix226 (.Y (nx225), .A0 (reg_idx_out_2), .A1 (ans[2]), .S0 (nx562)
             ) ;
    dffr reg_curr_idx_3 (.Q (curr_idx_3), .QB (\$dummy [36]), .D (nx235), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix236 (.Y (nx235), .A0 (curr_idx_3), .A1 (nx157), .S0 (nx564)) ;
    xnor2 ix120 (.Y (nx157), .A0 (curr_idx_3), .A1 (nx503)) ;
    nand03 ix504 (.Y (nx503), .A0 (curr_idx_2), .A1 (curr_idx_1), .A2 (
           curr_idx_0)) ;
    dffr idxReg_reg_q_3 (.Q (reg_idx_out_3), .QB (\$dummy [37]), .D (nx245), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix246 (.Y (nx245), .A0 (reg_idx_out_3), .A1 (ans[3]), .S0 (nx564)
             ) ;
    inv01 ix510 (.Y (compare_in1_inverted_0), .A (inp[0])) ;
    inv01 ix512 (.Y (compare_in1_inverted_1), .A (inp[1])) ;
    inv01 ix514 (.Y (compare_in1_inverted_2), .A (inp[2])) ;
    inv01 ix516 (.Y (compare_in1_inverted_3), .A (inp[3])) ;
    inv01 ix518 (.Y (compare_in1_inverted_4), .A (inp[4])) ;
    inv01 ix520 (.Y (compare_in1_inverted_5), .A (inp[5])) ;
    inv01 ix522 (.Y (compare_in1_inverted_6), .A (inp[6])) ;
    inv01 ix524 (.Y (compare_in1_inverted_7), .A (inp[7])) ;
    inv01 ix526 (.Y (compare_in1_inverted_8), .A (inp[8])) ;
    inv01 ix528 (.Y (compare_in1_inverted_9), .A (inp[9])) ;
    inv01 ix530 (.Y (compare_in1_inverted_10), .A (inp[10])) ;
    inv01 ix532 (.Y (compare_in1_inverted_11), .A (inp[11])) ;
    inv01 ix534 (.Y (compare_in1_inverted_12), .A (inp[12])) ;
    inv01 ix536 (.Y (compare_in1_inverted_13), .A (inp[13])) ;
    inv01 ix538 (.Y (compare_in1_inverted_14), .A (inp[14])) ;
    mux21_ni ix141 (.Y (nx140), .A0 (reg_val_out_0), .A1 (inp[0]), .S0 (nx566)
             ) ;
    xnor2 ix406 (.Y (nx405), .A0 (inp[15]), .A1 (nx411)) ;
    mux21_ni ix153 (.Y (nx152), .A0 (reg_val_out_1), .A1 (inp[1]), .S0 (nx566)
             ) ;
    mux21_ni ix165 (.Y (nx164), .A0 (reg_val_out_2), .A1 (inp[2]), .S0 (nx566)
             ) ;
    mux21_ni ix177 (.Y (nx176), .A0 (reg_val_out_3), .A1 (inp[3]), .S0 (nx566)
             ) ;
    mux21_ni ix189 (.Y (nx188), .A0 (reg_val_out_4), .A1 (inp[4]), .S0 (nx566)
             ) ;
    mux21_ni ix201 (.Y (nx200), .A0 (reg_val_out_5), .A1 (inp[5]), .S0 (nx566)
             ) ;
    mux21_ni ix213 (.Y (nx212), .A0 (reg_val_out_6), .A1 (inp[6]), .S0 (nx566)
             ) ;
    mux21_ni ix225 (.Y (nx224), .A0 (reg_val_out_7), .A1 (inp[7]), .S0 (nx568)
             ) ;
    mux21_ni ix237 (.Y (nx236), .A0 (reg_val_out_8), .A1 (inp[8]), .S0 (nx568)
             ) ;
    mux21_ni ix249 (.Y (nx248), .A0 (reg_val_out_9), .A1 (inp[9]), .S0 (nx568)
             ) ;
    mux21_ni ix261 (.Y (nx260), .A0 (reg_val_out_10), .A1 (inp[10]), .S0 (nx568)
             ) ;
    mux21_ni ix273 (.Y (nx272), .A0 (reg_val_out_11), .A1 (inp[11]), .S0 (nx568)
             ) ;
    mux21_ni ix285 (.Y (nx284), .A0 (reg_val_out_12), .A1 (inp[12]), .S0 (nx568)
             ) ;
    mux21_ni ix297 (.Y (nx296), .A0 (reg_val_out_13), .A1 (inp[13]), .S0 (nx568)
             ) ;
    mux21_ni ix309 (.Y (nx308), .A0 (reg_val_out_14), .A1 (inp[14]), .S0 (nx570)
             ) ;
    mux21_ni ix67 (.Y (ans[0]), .A0 (reg_idx_out_0), .A1 (curr_idx_0), .S0 (
             nx570)) ;
    xor2 ix166 (.Y (nx165), .A0 (curr_idx_0), .A1 (nx564)) ;
    mux21_ni ix91 (.Y (ans[1]), .A0 (reg_idx_out_1), .A1 (curr_idx_1), .S0 (
             nx570)) ;
    mux21_ni ix119 (.Y (ans[2]), .A0 (reg_idx_out_2), .A1 (curr_idx_2), .S0 (
             nx570)) ;
    mux21_ni ix133 (.Y (ans[3]), .A0 (reg_idx_out_3), .A1 (curr_idx_3), .S0 (
             nx570)) ;
    inv01 ix555 (.Y (nx556), .A (en)) ;
    inv02 ix557 (.Y (nx558), .A (nx556)) ;
    inv02 ix559 (.Y (nx560), .A (nx556)) ;
    inv02 ix561 (.Y (nx562), .A (nx556)) ;
    inv02 ix563 (.Y (nx564), .A (nx556)) ;
    inv02 ix565 (.Y (nx566), .A (nx54)) ;
    inv02 ix567 (.Y (nx568), .A (nx54)) ;
    inv02 ix569 (.Y (nx570), .A (nx54)) ;
endmodule


module NAdder_16 ( a, b, cin, s, cout ) ;

    input [15:0]a ;
    input [15:0]b ;
    input cin ;
    output [15:0]s ;
    output cout ;

    wire nx12, nx16, nx61, nx103, nx105, nx125, nx127, nx129, nx135, nx152, 
         nx153, nx154, nx155, nx156, nx157, nx158, nx159, nx160, nx161, nx162, 
         nx163, nx164, nx165, nx166, nx167, nx168, nx169, nx170, nx38, nx171, 
         nx172, nx173, nx174, nx175, nx176, nx177, nx62, nx178, nx179, nx180, 
         nx97, nx181, nx182, nx183, nx184, nx185, nx186, nx98, nx223, nx225;



    assign s[13] = s[14] ;
    assign s[12] = s[14] ;
    assign s[11] = s[14] ;
    assign s[10] = s[14] ;
    assign s[9] = s[14] ;
    assign s[8] = s[14] ;
    assign s[7] = s[14] ;
    assign s[6] = s[14] ;
    assign s[5] = s[14] ;
    assign s[4] = s[14] ;
    assign s[3] = s[14] ;
    assign s[2] = s[14] ;
    assign s[1] = s[14] ;
    assign s[0] = s[14] ;
    assign cout = s[14] ;
    fake_gnd ix25 (.Y (s[14])) ;
    xor2 ix13 (.Y (nx12), .A0 (a[8]), .A1 (b[8])) ;
    xnor2 ix104 (.Y (nx103), .A0 (a[7]), .A1 (b[7])) ;
    aoi22 ix106 (.Y (nx105), .A0 (b[6]), .A1 (a[6]), .B0 (nx16), .B1 (nx225)) ;
    xor2 ix17 (.Y (nx16), .A0 (a[6]), .A1 (b[6])) ;
    xor2 ix27 (.Y (nx61), .A0 (a[2]), .A1 (b[2])) ;
    xnor2 ix126 (.Y (nx125), .A0 (a[1]), .A1 (b[1])) ;
    nor02_2x ix128 (.Y (nx127), .A0 (b[0]), .A1 (a[0])) ;
    nand02 ix130 (.Y (nx129), .A0 (b[1]), .A1 (a[1])) ;
    nand02 ix136 (.Y (nx135), .A0 (b[7]), .A1 (a[7])) ;
    or02 ix187 (.Y (nx152), .A0 (a[13]), .A1 (b[13])) ;
    nor02_2x ix188 (.Y (nx153), .A0 (a[11]), .A1 (b[11])) ;
    nand02_2x ix189 (.Y (nx154), .A0 (a[11]), .A1 (b[11])) ;
    inv02 ix190 (.Y (nx155), .A (a[12])) ;
    inv02 ix191 (.Y (nx156), .A (b[12])) ;
    aoi22 ix192 (.Y (nx157), .A0 (b[12]), .A1 (nx155), .B0 (a[12]), .B1 (nx156)
          ) ;
    nor02_2x ix193 (.Y (nx158), .A0 (a[13]), .A1 (b[13])) ;
    nor02_2x ix194 (.Y (nx159), .A0 (nx157), .A1 (nx158)) ;
    aoi322 ix195 (.Y (nx160), .A0 (nx152), .A1 (b[12]), .A2 (a[12]), .B0 (a[13])
           , .B1 (b[13]), .C0 (nx98), .C1 (nx159)) ;
    inv02 ix196 (.Y (nx161), .A (a[15])) ;
    inv02 ix197 (.Y (nx162), .A (b[15])) ;
    aoi22 ix198 (.Y (nx163), .A0 (b[15]), .A1 (nx161), .B0 (a[15]), .B1 (nx162)
          ) ;
    and02 ix199 (.Y (nx164), .A0 (b[14]), .A1 (a[14])) ;
    nor02_2x ix200 (.Y (nx165), .A0 (nx223), .A1 (nx164)) ;
    oai21 ix201 (.Y (nx166), .A0 (b[14]), .A1 (a[14]), .B0 (nx223)) ;
    nor03_2x ix202 (.Y (nx167), .A0 (nx223), .A1 (b[14]), .A2 (a[14])) ;
    aoi21 ix203 (.Y (nx168), .A0 (nx223), .A1 (nx164), .B0 (nx167)) ;
    oai21 ix204 (.Y (nx169), .A0 (nx160), .A1 (nx166), .B0 (nx168)) ;
    ao21 reg_s_15 (.Y (s[15]), .A0 (nx160), .A1 (nx165), .B0 (nx169)) ;
    or02 ix205 (.Y (nx170), .A0 (a[3]), .A1 (b[3])) ;
    oai21 reg_nx38 (.Y (nx38), .A0 (nx125), .A1 (nx127), .B0 (nx129)) ;
    aoi332 ix206 (.Y (nx171), .A0 (nx170), .A1 (b[2]), .A2 (a[2]), .B0 (nx38), .B1 (
           nx61), .B2 (nx170), .C0 (a[3]), .C1 (b[3])) ;
    inv02 ix207 (.Y (nx172), .A (a[4])) ;
    inv02 ix208 (.Y (nx173), .A (b[4])) ;
    aoi22 ix209 (.Y (nx174), .A0 (b[4]), .A1 (nx172), .B0 (a[4]), .B1 (nx173)) ;
    nor02_2x ix210 (.Y (nx175), .A0 (a[5]), .A1 (b[5])) ;
    inv02 ix211 (.Y (nx176), .A (a[5])) ;
    inv02 ix212 (.Y (nx177), .A (b[5])) ;
    oai332 reg_nx62 (.Y (nx62), .A0 (nx171), .A1 (nx174), .A2 (nx175), .B0 (
           nx175), .B1 (nx173), .B2 (nx172), .C0 (nx176), .C1 (nx177)) ;
    nor02_2x ix213 (.Y (nx178), .A0 (nx103), .A1 (nx105)) ;
    inv02 ix214 (.Y (nx179), .A (nx135)) ;
    and02 ix215 (.Y (nx180), .A0 (b[8]), .A1 (a[8])) ;
    oai32 reg_nx97 (.Y (nx97), .A0 (nx178), .A1 (nx179), .A2 (nx180), .B0 (nx180
          ), .B1 (nx12)) ;
    nor02_2x ix216 (.Y (nx181), .A0 (a[9]), .A1 (b[9])) ;
    and02 ix217 (.Y (nx182), .A0 (a[9]), .A1 (b[9])) ;
    nor02_2x ix218 (.Y (nx183), .A0 (b[10]), .A1 (a[10])) ;
    or04 ix219 (.Y (nx184), .A0 (nx181), .A1 (nx182), .A2 (nx183), .A3 (nx153)
         ) ;
    or02 ix220 (.Y (nx185), .A0 (b[10]), .A1 (a[10])) ;
    aoi22 ix221 (.Y (nx186), .A0 (nx185), .A1 (nx182), .B0 (b[10]), .B1 (a[10])
          ) ;
    oai221 reg_nx98 (.Y (nx98), .A0 (nx97), .A1 (nx184), .B0 (nx186), .B1 (nx153
           ), .C0 (nx154)) ;
    buf02 ix222 (.Y (nx223), .A (nx163)) ;
    buf02 ix224 (.Y (nx225), .A (nx62)) ;
endmodule


module ComputationBlock ( img_data_col_0, img_data_col_1, img_data_col_2, 
                          img_data_col_3, img_data_col_4, img_load, img_reset, 
                          filter_data_word, filter_load, filter_reset, start, 
                          operation, compute_relu, filter_size, output1_init, 
                          output2_init, output1, output2, buffer_ready, ready, 
                          clk, en, reset ) ;

    input [15:0]img_data_col_0 ;
    input [15:0]img_data_col_1 ;
    input [15:0]img_data_col_2 ;
    input [15:0]img_data_col_3 ;
    input [15:0]img_data_col_4 ;
    input img_load ;
    input img_reset ;
    input [15:0]filter_data_word ;
    input filter_load ;
    input filter_reset ;
    input start ;
    input operation ;
    input compute_relu ;
    input filter_size ;
    input [15:0]output1_init ;
    input [15:0]output2_init ;
    output [15:0]output1 ;
    output [15:0]output2 ;
    output buffer_ready ;
    output ready ;
    input clk ;
    input en ;
    input reset ;

    wire img_data_0__15, img_data_0__14, img_data_0__13, img_data_0__12, 
         img_data_0__11, img_data_0__10, img_data_0__9, img_data_0__8, 
         img_data_0__7, img_data_0__6, img_data_0__5, img_data_0__4, 
         img_data_0__3, img_data_0__2, img_data_0__1, img_data_0__0, 
         img_data_1__15, img_data_1__14, img_data_1__13, img_data_1__12, 
         img_data_1__11, img_data_1__10, img_data_1__9, img_data_1__8, 
         img_data_1__7, img_data_1__6, img_data_1__5, img_data_1__4, 
         img_data_1__3, img_data_1__2, img_data_1__1, img_data_1__0, 
         img_data_2__15, img_data_2__14, img_data_2__13, img_data_2__12, 
         img_data_2__11, img_data_2__10, img_data_2__9, img_data_2__8, 
         img_data_2__7, img_data_2__6, img_data_2__5, img_data_2__4, 
         img_data_2__3, img_data_2__2, img_data_2__1, img_data_2__0, 
         img_data_3__15, img_data_3__14, img_data_3__13, img_data_3__12, 
         img_data_3__11, img_data_3__10, img_data_3__9, img_data_3__8, 
         img_data_3__7, img_data_3__6, img_data_3__5, img_data_3__4, 
         img_data_3__3, img_data_3__2, img_data_3__1, img_data_3__0, 
         img_data_4__15, img_data_4__14, img_data_4__13, img_data_4__12, 
         img_data_4__11, img_data_4__10, img_data_4__9, img_data_4__8, 
         img_data_4__7, img_data_4__6, img_data_4__5, img_data_4__4, 
         img_data_4__3, img_data_4__2, img_data_4__1, img_data_4__0, 
         img_data_5__15, img_data_5__14, img_data_5__13, img_data_5__12, 
         img_data_5__11, img_data_5__10, img_data_5__9, img_data_5__8, 
         img_data_5__7, img_data_5__6, img_data_5__5, img_data_5__4, 
         img_data_5__3, img_data_5__2, img_data_5__1, img_data_5__0, 
         img_data_6__15, img_data_6__14, img_data_6__13, img_data_6__12, 
         img_data_6__11, img_data_6__10, img_data_6__9, img_data_6__8, 
         img_data_6__7, img_data_6__6, img_data_6__5, img_data_6__4, 
         img_data_6__3, img_data_6__2, img_data_6__1, img_data_6__0, 
         img_data_7__15, img_data_7__14, img_data_7__13, img_data_7__12, 
         img_data_7__11, img_data_7__10, img_data_7__9, img_data_7__8, 
         img_data_7__7, img_data_7__6, img_data_7__5, img_data_7__4, 
         img_data_7__3, img_data_7__2, img_data_7__1, img_data_7__0, 
         img_data_8__15, img_data_8__14, img_data_8__13, img_data_8__12, 
         img_data_8__11, img_data_8__10, img_data_8__9, img_data_8__8, 
         img_data_8__7, img_data_8__6, img_data_8__5, img_data_8__4, 
         img_data_8__3, img_data_8__2, img_data_8__1, img_data_8__0, 
         img_data_9__15, img_data_9__14, img_data_9__13, img_data_9__12, 
         img_data_9__11, img_data_9__10, img_data_9__9, img_data_9__8, 
         img_data_9__7, img_data_9__6, img_data_9__5, img_data_9__4, 
         img_data_9__3, img_data_9__2, img_data_9__1, img_data_9__0, 
         img_data_10__15, img_data_10__14, img_data_10__13, img_data_10__12, 
         img_data_10__11, img_data_10__10, img_data_10__9, img_data_10__8, 
         img_data_10__7, img_data_10__6, img_data_10__5, img_data_10__4, 
         img_data_10__3, img_data_10__2, img_data_10__1, img_data_10__0, 
         img_data_11__15, img_data_11__14, img_data_11__13, img_data_11__12, 
         img_data_11__11, img_data_11__10, img_data_11__9, img_data_11__8, 
         img_data_11__7, img_data_11__6, img_data_11__5, img_data_11__4, 
         img_data_11__3, img_data_11__2, img_data_11__1, img_data_11__0, 
         img_data_12__15, img_data_12__14, img_data_12__13, img_data_12__12, 
         img_data_12__11, img_data_12__10, img_data_12__9, img_data_12__8, 
         img_data_12__7, img_data_12__6, img_data_12__5, img_data_12__4, 
         img_data_12__3, img_data_12__2, img_data_12__1, img_data_12__0, 
         img_data_13__15, img_data_13__14, img_data_13__13, img_data_13__12, 
         img_data_13__11, img_data_13__10, img_data_13__9, img_data_13__8, 
         img_data_13__7, img_data_13__6, img_data_13__5, img_data_13__4, 
         img_data_13__3, img_data_13__2, img_data_13__1, img_data_13__0, 
         img_data_14__15, img_data_14__14, img_data_14__13, img_data_14__12, 
         img_data_14__11, img_data_14__10, img_data_14__9, img_data_14__8, 
         img_data_14__7, img_data_14__6, img_data_14__5, img_data_14__4, 
         img_data_14__3, img_data_14__2, img_data_14__1, img_data_14__0, 
         img_data_15__15, img_data_15__14, img_data_15__13, img_data_15__12, 
         img_data_15__11, img_data_15__10, img_data_15__9, img_data_15__8, 
         img_data_15__7, img_data_15__6, img_data_15__5, img_data_15__4, 
         img_data_15__3, img_data_15__2, img_data_15__1, img_data_15__0, 
         img_data_16__15, img_data_16__14, img_data_16__13, img_data_16__12, 
         img_data_16__11, img_data_16__10, img_data_16__9, img_data_16__8, 
         img_data_16__7, img_data_16__6, img_data_16__5, img_data_16__4, 
         img_data_16__3, img_data_16__2, img_data_16__1, img_data_16__0, 
         img_data_17__15, img_data_17__14, img_data_17__13, img_data_17__12, 
         img_data_17__11, img_data_17__10, img_data_17__9, img_data_17__8, 
         img_data_17__7, img_data_17__6, img_data_17__5, img_data_17__4, 
         img_data_17__3, img_data_17__2, img_data_17__1, img_data_17__0, 
         img_data_18__15, img_data_18__14, img_data_18__13, img_data_18__12, 
         img_data_18__11, img_data_18__10, img_data_18__9, img_data_18__8, 
         img_data_18__7, img_data_18__6, img_data_18__5, img_data_18__4, 
         img_data_18__3, img_data_18__2, img_data_18__1, img_data_18__0, 
         img_data_19__15, img_data_19__14, img_data_19__13, img_data_19__12, 
         img_data_19__11, img_data_19__10, img_data_19__9, img_data_19__8, 
         img_data_19__7, img_data_19__6, img_data_19__5, img_data_19__4, 
         img_data_19__3, img_data_19__2, img_data_19__1, img_data_19__0, 
         img_data_20__15, img_data_20__14, img_data_20__13, img_data_20__12, 
         img_data_20__11, img_data_20__10, img_data_20__9, img_data_20__8, 
         img_data_20__7, img_data_20__6, img_data_20__5, img_data_20__4, 
         img_data_20__3, img_data_20__2, img_data_20__1, img_data_20__0, 
         img_data_21__15, img_data_21__14, img_data_21__13, img_data_21__12, 
         img_data_21__11, img_data_21__10, img_data_21__9, img_data_21__8, 
         img_data_21__7, img_data_21__6, img_data_21__5, img_data_21__4, 
         img_data_21__3, img_data_21__2, img_data_21__1, img_data_21__0, 
         img_data_22__15, img_data_22__14, img_data_22__13, img_data_22__12, 
         img_data_22__11, img_data_22__10, img_data_22__9, img_data_22__8, 
         img_data_22__7, img_data_22__6, img_data_22__5, img_data_22__4, 
         img_data_22__3, img_data_22__2, img_data_22__1, img_data_22__0, 
         img_data_23__15, img_data_23__14, img_data_23__13, img_data_23__12, 
         img_data_23__11, img_data_23__10, img_data_23__9, img_data_23__8, 
         img_data_23__7, img_data_23__6, img_data_23__5, img_data_23__4, 
         img_data_23__3, img_data_23__2, img_data_23__1, img_data_23__0, 
         img_data_24__15, img_data_24__14, img_data_24__13, img_data_24__12, 
         img_data_24__11, img_data_24__10, img_data_24__9, img_data_24__8, 
         img_data_24__7, img_data_24__6, img_data_24__5, img_data_24__4, 
         img_data_24__3, img_data_24__2, img_data_24__1, img_data_24__0, 
         filter_data_0__15, filter_data_0__14, filter_data_0__13, 
         filter_data_0__12, filter_data_0__11, filter_data_0__10, 
         filter_data_0__9, filter_data_0__8, filter_data_0__7, filter_data_0__6, 
         filter_data_0__5, filter_data_0__4, filter_data_0__3, filter_data_0__2, 
         filter_data_0__1, filter_data_0__0, filter_data_1__15, 
         filter_data_1__14, filter_data_1__13, filter_data_1__12, 
         filter_data_1__11, filter_data_1__10, filter_data_1__9, 
         filter_data_1__8, filter_data_1__7, filter_data_1__6, filter_data_1__5, 
         filter_data_1__4, filter_data_1__3, filter_data_1__2, filter_data_1__1, 
         filter_data_1__0, filter_data_2__15, filter_data_2__14, 
         filter_data_2__13, filter_data_2__12, filter_data_2__11, 
         filter_data_2__10, filter_data_2__9, filter_data_2__8, filter_data_2__7, 
         filter_data_2__6, filter_data_2__5, filter_data_2__4, filter_data_2__3, 
         filter_data_2__2, filter_data_2__1, filter_data_2__0, filter_data_3__15, 
         filter_data_3__14, filter_data_3__13, filter_data_3__12, 
         filter_data_3__11, filter_data_3__10, filter_data_3__9, 
         filter_data_3__8, filter_data_3__7, filter_data_3__6, filter_data_3__5, 
         filter_data_3__4, filter_data_3__3, filter_data_3__2, filter_data_3__1, 
         filter_data_3__0, filter_data_4__15, filter_data_4__14, 
         filter_data_4__13, filter_data_4__12, filter_data_4__11, 
         filter_data_4__10, filter_data_4__9, filter_data_4__8, filter_data_4__7, 
         filter_data_4__6, filter_data_4__5, filter_data_4__4, filter_data_4__3, 
         filter_data_4__2, filter_data_4__1, filter_data_4__0, filter_data_5__15, 
         filter_data_5__14, filter_data_5__13, filter_data_5__12, 
         filter_data_5__11, filter_data_5__10, filter_data_5__9, 
         filter_data_5__8, filter_data_5__7, filter_data_5__6, filter_data_5__5, 
         filter_data_5__4, filter_data_5__3, filter_data_5__2, filter_data_5__1, 
         filter_data_5__0, filter_data_6__15, filter_data_6__14, 
         filter_data_6__13, filter_data_6__12, filter_data_6__11, 
         filter_data_6__10, filter_data_6__9, filter_data_6__8, filter_data_6__7, 
         filter_data_6__6, filter_data_6__5, filter_data_6__4, filter_data_6__3, 
         filter_data_6__2, filter_data_6__1, filter_data_6__0, filter_data_7__15, 
         filter_data_7__14, filter_data_7__13, filter_data_7__12, 
         filter_data_7__11, filter_data_7__10, filter_data_7__9, 
         filter_data_7__8, filter_data_7__7, filter_data_7__6, filter_data_7__5, 
         filter_data_7__4, filter_data_7__3, filter_data_7__2, filter_data_7__1, 
         filter_data_7__0, filter_data_8__15, filter_data_8__14, 
         filter_data_8__13, filter_data_8__12, filter_data_8__11, 
         filter_data_8__10, filter_data_8__9, filter_data_8__8, filter_data_8__7, 
         filter_data_8__6, filter_data_8__5, filter_data_8__4, filter_data_8__3, 
         filter_data_8__2, filter_data_8__1, filter_data_8__0, filter_data_9__15, 
         filter_data_9__14, filter_data_9__13, filter_data_9__12, 
         filter_data_9__11, filter_data_9__10, filter_data_9__9, 
         filter_data_9__8, filter_data_9__7, filter_data_9__6, filter_data_9__5, 
         filter_data_9__4, filter_data_9__3, filter_data_9__2, filter_data_9__1, 
         filter_data_9__0, filter_data_10__15, filter_data_10__14, 
         filter_data_10__13, filter_data_10__12, filter_data_10__11, 
         filter_data_10__10, filter_data_10__9, filter_data_10__8, 
         filter_data_10__7, filter_data_10__6, filter_data_10__5, 
         filter_data_10__4, filter_data_10__3, filter_data_10__2, 
         filter_data_10__1, filter_data_10__0, filter_data_11__15, 
         filter_data_11__14, filter_data_11__13, filter_data_11__12, 
         filter_data_11__11, filter_data_11__10, filter_data_11__9, 
         filter_data_11__8, filter_data_11__7, filter_data_11__6, 
         filter_data_11__5, filter_data_11__4, filter_data_11__3, 
         filter_data_11__2, filter_data_11__1, filter_data_11__0, 
         filter_data_12__15, filter_data_12__14, filter_data_12__13, 
         filter_data_12__12, filter_data_12__11, filter_data_12__10, 
         filter_data_12__9, filter_data_12__8, filter_data_12__7, 
         filter_data_12__6, filter_data_12__5, filter_data_12__4, 
         filter_data_12__3, filter_data_12__2, filter_data_12__1, 
         filter_data_12__0, filter_data_13__15, filter_data_13__14, 
         filter_data_13__13, filter_data_13__12, filter_data_13__11, 
         filter_data_13__10, filter_data_13__9, filter_data_13__8, 
         filter_data_13__7, filter_data_13__6, filter_data_13__5, 
         filter_data_13__4, filter_data_13__3, filter_data_13__2, 
         filter_data_13__1, filter_data_13__0, filter_data_14__15, 
         filter_data_14__14, filter_data_14__13, filter_data_14__12, 
         filter_data_14__11, filter_data_14__10, filter_data_14__9, 
         filter_data_14__8, filter_data_14__7, filter_data_14__6, 
         filter_data_14__5, filter_data_14__4, filter_data_14__3, 
         filter_data_14__2, filter_data_14__1, filter_data_14__0, 
         filter_data_15__15, filter_data_15__14, filter_data_15__13, 
         filter_data_15__12, filter_data_15__11, filter_data_15__10, 
         filter_data_15__9, filter_data_15__8, filter_data_15__7, 
         filter_data_15__6, filter_data_15__5, filter_data_15__4, 
         filter_data_15__3, filter_data_15__2, filter_data_15__1, 
         filter_data_15__0, filter_data_16__15, filter_data_16__14, 
         filter_data_16__13, filter_data_16__12, filter_data_16__11, 
         filter_data_16__10, filter_data_16__9, filter_data_16__8, 
         filter_data_16__7, filter_data_16__6, filter_data_16__5, 
         filter_data_16__4, filter_data_16__3, filter_data_16__2, 
         filter_data_16__1, filter_data_16__0, filter_data_17__15, 
         filter_data_17__14, filter_data_17__13, filter_data_17__12, 
         filter_data_17__11, filter_data_17__10, filter_data_17__9, 
         filter_data_17__8, filter_data_17__7, filter_data_17__6, 
         filter_data_17__5, filter_data_17__4, filter_data_17__3, 
         filter_data_17__2, filter_data_17__1, filter_data_17__0, 
         filter_data_18__15, filter_data_18__14, filter_data_18__13, 
         filter_data_18__12, filter_data_18__11, filter_data_18__10, 
         filter_data_18__9, filter_data_18__8, filter_data_18__7, 
         filter_data_18__6, filter_data_18__5, filter_data_18__4, 
         filter_data_18__3, filter_data_18__2, filter_data_18__1, 
         filter_data_18__0, filter_data_19__15, filter_data_19__14, 
         filter_data_19__13, filter_data_19__12, filter_data_19__11, 
         filter_data_19__10, filter_data_19__9, filter_data_19__8, 
         filter_data_19__7, filter_data_19__6, filter_data_19__5, 
         filter_data_19__4, filter_data_19__3, filter_data_19__2, 
         filter_data_19__1, filter_data_19__0, filter_data_20__15, 
         filter_data_20__14, filter_data_20__13, filter_data_20__12, 
         filter_data_20__11, filter_data_20__10, filter_data_20__9, 
         filter_data_20__8, filter_data_20__7, filter_data_20__6, 
         filter_data_20__5, filter_data_20__4, filter_data_20__3, 
         filter_data_20__2, filter_data_20__1, filter_data_20__0, 
         filter_data_21__15, filter_data_21__14, filter_data_21__13, 
         filter_data_21__12, filter_data_21__11, filter_data_21__10, 
         filter_data_21__9, filter_data_21__8, filter_data_21__7, 
         filter_data_21__6, filter_data_21__5, filter_data_21__4, 
         filter_data_21__3, filter_data_21__2, filter_data_21__1, 
         filter_data_21__0, filter_data_22__15, filter_data_22__14, 
         filter_data_22__13, filter_data_22__12, filter_data_22__11, 
         filter_data_22__10, filter_data_22__9, filter_data_22__8, 
         filter_data_22__7, filter_data_22__6, filter_data_22__5, 
         filter_data_22__4, filter_data_22__3, filter_data_22__2, 
         filter_data_22__1, filter_data_22__0, filter_data_23__15, 
         filter_data_23__14, filter_data_23__13, filter_data_23__12, 
         filter_data_23__11, filter_data_23__10, filter_data_23__9, 
         filter_data_23__8, filter_data_23__7, filter_data_23__6, 
         filter_data_23__5, filter_data_23__4, filter_data_23__3, 
         filter_data_23__2, filter_data_23__1, filter_data_23__0, 
         filter_data_24__15, filter_data_24__14, filter_data_24__13, 
         filter_data_24__12, filter_data_24__11, filter_data_24__10, 
         filter_data_24__9, filter_data_24__8, filter_data_24__7, 
         filter_data_24__6, filter_data_24__5, filter_data_24__4, 
         filter_data_24__3, filter_data_24__2, filter_data_24__1, 
         filter_data_24__0, d_cache_arr_0__31, d_cache_arr_0__30, 
         d_cache_arr_0__29, d_cache_arr_0__28, d_cache_arr_0__27, 
         d_cache_arr_0__26, d_cache_arr_0__25, d_cache_arr_0__24, 
         d_cache_arr_0__23, d_cache_arr_0__22, d_cache_arr_0__21, 
         d_cache_arr_0__20, d_cache_arr_0__19, d_cache_arr_0__18, 
         d_cache_arr_0__17, d_cache_arr_0__16, d_cache_arr_0__15, 
         d_cache_arr_0__14, d_cache_arr_0__13, d_cache_arr_0__12, 
         d_cache_arr_0__11, d_cache_arr_0__10, d_cache_arr_0__9, 
         d_cache_arr_0__8, d_cache_arr_0__7, d_cache_arr_0__6, d_cache_arr_0__5, 
         d_cache_arr_0__4, d_cache_arr_0__3, d_cache_arr_0__2, d_cache_arr_0__1, 
         d_cache_arr_0__0, d_cache_arr_1__31, d_cache_arr_1__30, 
         d_cache_arr_1__29, d_cache_arr_1__28, d_cache_arr_1__27, 
         d_cache_arr_1__26, d_cache_arr_1__25, d_cache_arr_1__24, 
         d_cache_arr_1__23, d_cache_arr_1__22, d_cache_arr_1__21, 
         d_cache_arr_1__20, d_cache_arr_1__19, d_cache_arr_1__18, 
         d_cache_arr_1__17, d_cache_arr_1__16, d_cache_arr_1__15, 
         d_cache_arr_1__14, d_cache_arr_1__13, d_cache_arr_1__12, 
         d_cache_arr_1__11, d_cache_arr_1__10, d_cache_arr_1__9, 
         d_cache_arr_1__8, d_cache_arr_1__7, d_cache_arr_1__6, d_cache_arr_1__5, 
         d_cache_arr_1__4, d_cache_arr_1__3, d_cache_arr_1__2, d_cache_arr_1__1, 
         d_cache_arr_1__0, d_cache_arr_2__31, d_cache_arr_2__30, 
         d_cache_arr_2__29, d_cache_arr_2__28, d_cache_arr_2__27, 
         d_cache_arr_2__26, d_cache_arr_2__25, d_cache_arr_2__24, 
         d_cache_arr_2__23, d_cache_arr_2__22, d_cache_arr_2__21, 
         d_cache_arr_2__20, d_cache_arr_2__19, d_cache_arr_2__18, 
         d_cache_arr_2__17, d_cache_arr_2__16, d_cache_arr_2__15, 
         d_cache_arr_2__14, d_cache_arr_2__13, d_cache_arr_2__12, 
         d_cache_arr_2__11, d_cache_arr_2__10, d_cache_arr_2__9, 
         d_cache_arr_2__8, d_cache_arr_2__7, d_cache_arr_2__6, d_cache_arr_2__5, 
         d_cache_arr_2__4, d_cache_arr_2__3, d_cache_arr_2__2, d_cache_arr_2__1, 
         d_cache_arr_2__0, d_cache_arr_3__31, d_cache_arr_3__30, 
         d_cache_arr_3__29, d_cache_arr_3__28, d_cache_arr_3__27, 
         d_cache_arr_3__26, d_cache_arr_3__25, d_cache_arr_3__24, 
         d_cache_arr_3__23, d_cache_arr_3__22, d_cache_arr_3__21, 
         d_cache_arr_3__20, d_cache_arr_3__19, d_cache_arr_3__18, 
         d_cache_arr_3__17, d_cache_arr_3__16, d_cache_arr_3__15, 
         d_cache_arr_3__14, d_cache_arr_3__13, d_cache_arr_3__12, 
         d_cache_arr_3__11, d_cache_arr_3__10, d_cache_arr_3__9, 
         d_cache_arr_3__8, d_cache_arr_3__7, d_cache_arr_3__6, d_cache_arr_3__5, 
         d_cache_arr_3__4, d_cache_arr_3__3, d_cache_arr_3__2, d_cache_arr_3__1, 
         d_cache_arr_3__0, d_cache_arr_4__31, d_cache_arr_4__30, 
         d_cache_arr_4__29, d_cache_arr_4__28, d_cache_arr_4__27, 
         d_cache_arr_4__26, d_cache_arr_4__25, d_cache_arr_4__24, 
         d_cache_arr_4__23, d_cache_arr_4__22, d_cache_arr_4__21, 
         d_cache_arr_4__20, d_cache_arr_4__19, d_cache_arr_4__18, 
         d_cache_arr_4__17, d_cache_arr_4__16, d_cache_arr_4__15, 
         d_cache_arr_4__14, d_cache_arr_4__13, d_cache_arr_4__12, 
         d_cache_arr_4__11, d_cache_arr_4__10, d_cache_arr_4__9, 
         d_cache_arr_4__8, d_cache_arr_4__7, d_cache_arr_4__6, d_cache_arr_4__5, 
         d_cache_arr_4__4, d_cache_arr_4__3, d_cache_arr_4__2, d_cache_arr_4__1, 
         d_cache_arr_4__0, d_cache_arr_5__31, d_cache_arr_5__30, 
         d_cache_arr_5__29, d_cache_arr_5__28, d_cache_arr_5__27, 
         d_cache_arr_5__26, d_cache_arr_5__25, d_cache_arr_5__24, 
         d_cache_arr_5__23, d_cache_arr_5__22, d_cache_arr_5__21, 
         d_cache_arr_5__20, d_cache_arr_5__19, d_cache_arr_5__18, 
         d_cache_arr_5__17, d_cache_arr_5__16, d_cache_arr_5__15, 
         d_cache_arr_5__14, d_cache_arr_5__13, d_cache_arr_5__12, 
         d_cache_arr_5__11, d_cache_arr_5__10, d_cache_arr_5__9, 
         d_cache_arr_5__8, d_cache_arr_5__7, d_cache_arr_5__6, d_cache_arr_5__5, 
         d_cache_arr_5__4, d_cache_arr_5__3, d_cache_arr_5__2, d_cache_arr_5__1, 
         d_cache_arr_5__0, d_cache_arr_6__31, d_cache_arr_6__30, 
         d_cache_arr_6__29, d_cache_arr_6__28, d_cache_arr_6__27, 
         d_cache_arr_6__26, d_cache_arr_6__25, d_cache_arr_6__24, 
         d_cache_arr_6__23, d_cache_arr_6__22, d_cache_arr_6__21, 
         d_cache_arr_6__20, d_cache_arr_6__19, d_cache_arr_6__18, 
         d_cache_arr_6__17, d_cache_arr_6__16, d_cache_arr_6__15, 
         d_cache_arr_6__14, d_cache_arr_6__13, d_cache_arr_6__12, 
         d_cache_arr_6__11, d_cache_arr_6__10, d_cache_arr_6__9, 
         d_cache_arr_6__8, d_cache_arr_6__7, d_cache_arr_6__6, d_cache_arr_6__5, 
         d_cache_arr_6__4, d_cache_arr_6__3, d_cache_arr_6__2, d_cache_arr_6__1, 
         d_cache_arr_6__0, d_cache_arr_7__31, d_cache_arr_7__30, 
         d_cache_arr_7__29, d_cache_arr_7__28, d_cache_arr_7__27, 
         d_cache_arr_7__26, d_cache_arr_7__25, d_cache_arr_7__24, 
         d_cache_arr_7__23, d_cache_arr_7__22, d_cache_arr_7__21, 
         d_cache_arr_7__20, d_cache_arr_7__19, d_cache_arr_7__18, 
         d_cache_arr_7__17, d_cache_arr_7__16, d_cache_arr_7__15, 
         d_cache_arr_7__14, d_cache_arr_7__13, d_cache_arr_7__12, 
         d_cache_arr_7__11, d_cache_arr_7__10, d_cache_arr_7__9, 
         d_cache_arr_7__8, d_cache_arr_7__7, d_cache_arr_7__6, d_cache_arr_7__5, 
         d_cache_arr_7__4, d_cache_arr_7__3, d_cache_arr_7__2, d_cache_arr_7__1, 
         d_cache_arr_7__0, d_cache_arr_8__31, d_cache_arr_8__30, 
         d_cache_arr_8__29, d_cache_arr_8__28, d_cache_arr_8__27, 
         d_cache_arr_8__26, d_cache_arr_8__25, d_cache_arr_8__24, 
         d_cache_arr_8__23, d_cache_arr_8__22, d_cache_arr_8__21, 
         d_cache_arr_8__20, d_cache_arr_8__19, d_cache_arr_8__18, 
         d_cache_arr_8__17, d_cache_arr_8__16, d_cache_arr_8__15, 
         d_cache_arr_8__14, d_cache_arr_8__13, d_cache_arr_8__12, 
         d_cache_arr_8__11, d_cache_arr_8__10, d_cache_arr_8__9, 
         d_cache_arr_8__8, d_cache_arr_8__7, d_cache_arr_8__6, d_cache_arr_8__5, 
         d_cache_arr_8__4, d_cache_arr_8__3, d_cache_arr_8__2, d_cache_arr_8__1, 
         d_cache_arr_8__0, d_cache_arr_9__31, d_cache_arr_9__30, 
         d_cache_arr_9__29, d_cache_arr_9__28, d_cache_arr_9__27, 
         d_cache_arr_9__26, d_cache_arr_9__25, d_cache_arr_9__24, 
         d_cache_arr_9__23, d_cache_arr_9__22, d_cache_arr_9__21, 
         d_cache_arr_9__20, d_cache_arr_9__19, d_cache_arr_9__18, 
         d_cache_arr_9__17, d_cache_arr_9__16, d_cache_arr_9__15, 
         d_cache_arr_9__14, d_cache_arr_9__13, d_cache_arr_9__12, 
         d_cache_arr_9__11, d_cache_arr_9__10, d_cache_arr_9__9, 
         d_cache_arr_9__8, d_cache_arr_9__7, d_cache_arr_9__6, d_cache_arr_9__5, 
         d_cache_arr_9__4, d_cache_arr_9__3, d_cache_arr_9__2, d_cache_arr_9__1, 
         d_cache_arr_9__0, d_cache_arr_10__31, d_cache_arr_10__30, 
         d_cache_arr_10__29, d_cache_arr_10__28, d_cache_arr_10__27, 
         d_cache_arr_10__26, d_cache_arr_10__25, d_cache_arr_10__24, 
         d_cache_arr_10__23, d_cache_arr_10__22, d_cache_arr_10__21, 
         d_cache_arr_10__20, d_cache_arr_10__19, d_cache_arr_10__18, 
         d_cache_arr_10__17, d_cache_arr_10__16, d_cache_arr_10__15, 
         d_cache_arr_10__14, d_cache_arr_10__13, d_cache_arr_10__12, 
         d_cache_arr_10__11, d_cache_arr_10__10, d_cache_arr_10__9, 
         d_cache_arr_10__8, d_cache_arr_10__7, d_cache_arr_10__6, 
         d_cache_arr_10__5, d_cache_arr_10__4, d_cache_arr_10__3, 
         d_cache_arr_10__2, d_cache_arr_10__1, d_cache_arr_10__0, 
         d_cache_arr_11__31, d_cache_arr_11__30, d_cache_arr_11__29, 
         d_cache_arr_11__28, d_cache_arr_11__27, d_cache_arr_11__26, 
         d_cache_arr_11__25, d_cache_arr_11__24, d_cache_arr_11__23, 
         d_cache_arr_11__22, d_cache_arr_11__21, d_cache_arr_11__20, 
         d_cache_arr_11__19, d_cache_arr_11__18, d_cache_arr_11__17, 
         d_cache_arr_11__16, d_cache_arr_11__15, d_cache_arr_11__14, 
         d_cache_arr_11__13, d_cache_arr_11__12, d_cache_arr_11__11, 
         d_cache_arr_11__10, d_cache_arr_11__9, d_cache_arr_11__8, 
         d_cache_arr_11__7, d_cache_arr_11__6, d_cache_arr_11__5, 
         d_cache_arr_11__4, d_cache_arr_11__3, d_cache_arr_11__2, 
         d_cache_arr_11__1, d_cache_arr_11__0, d_cache_arr_12__31, 
         d_cache_arr_12__30, d_cache_arr_12__29, d_cache_arr_12__28, 
         d_cache_arr_12__27, d_cache_arr_12__26, d_cache_arr_12__25, 
         d_cache_arr_12__24, d_cache_arr_12__23, d_cache_arr_12__22, 
         d_cache_arr_12__21, d_cache_arr_12__20, d_cache_arr_12__19, 
         d_cache_arr_12__18, d_cache_arr_12__17, d_cache_arr_12__16, 
         d_cache_arr_12__15, d_cache_arr_12__14, d_cache_arr_12__13, 
         d_cache_arr_12__12, d_cache_arr_12__11, d_cache_arr_12__10, 
         d_cache_arr_12__9, d_cache_arr_12__8, d_cache_arr_12__7, 
         d_cache_arr_12__6, d_cache_arr_12__5, d_cache_arr_12__4, 
         d_cache_arr_12__3, d_cache_arr_12__2, d_cache_arr_12__1, 
         d_cache_arr_12__0, d_cache_arr_13__31, d_cache_arr_13__30, 
         d_cache_arr_13__29, d_cache_arr_13__28, d_cache_arr_13__27, 
         d_cache_arr_13__26, d_cache_arr_13__25, d_cache_arr_13__24, 
         d_cache_arr_13__23, d_cache_arr_13__22, d_cache_arr_13__21, 
         d_cache_arr_13__20, d_cache_arr_13__19, d_cache_arr_13__18, 
         d_cache_arr_13__17, d_cache_arr_13__16, d_cache_arr_13__15, 
         d_cache_arr_13__14, d_cache_arr_13__13, d_cache_arr_13__12, 
         d_cache_arr_13__11, d_cache_arr_13__10, d_cache_arr_13__9, 
         d_cache_arr_13__8, d_cache_arr_13__7, d_cache_arr_13__6, 
         d_cache_arr_13__5, d_cache_arr_13__4, d_cache_arr_13__3, 
         d_cache_arr_13__2, d_cache_arr_13__1, d_cache_arr_13__0, 
         d_cache_arr_14__31, d_cache_arr_14__30, d_cache_arr_14__29, 
         d_cache_arr_14__28, d_cache_arr_14__27, d_cache_arr_14__26, 
         d_cache_arr_14__25, d_cache_arr_14__24, d_cache_arr_14__23, 
         d_cache_arr_14__22, d_cache_arr_14__21, d_cache_arr_14__20, 
         d_cache_arr_14__19, d_cache_arr_14__18, d_cache_arr_14__17, 
         d_cache_arr_14__16, d_cache_arr_14__15, d_cache_arr_14__14, 
         d_cache_arr_14__13, d_cache_arr_14__12, d_cache_arr_14__11, 
         d_cache_arr_14__10, d_cache_arr_14__9, d_cache_arr_14__8, 
         d_cache_arr_14__7, d_cache_arr_14__6, d_cache_arr_14__5, 
         d_cache_arr_14__4, d_cache_arr_14__3, d_cache_arr_14__2, 
         d_cache_arr_14__1, d_cache_arr_14__0, d_cache_arr_15__31, 
         d_cache_arr_15__30, d_cache_arr_15__29, d_cache_arr_15__28, 
         d_cache_arr_15__27, d_cache_arr_15__26, d_cache_arr_15__25, 
         d_cache_arr_15__24, d_cache_arr_15__23, d_cache_arr_15__22, 
         d_cache_arr_15__21, d_cache_arr_15__20, d_cache_arr_15__19, 
         d_cache_arr_15__18, d_cache_arr_15__17, d_cache_arr_15__16, 
         d_cache_arr_15__15, d_cache_arr_15__14, d_cache_arr_15__13, 
         d_cache_arr_15__12, d_cache_arr_15__11, d_cache_arr_15__10, 
         d_cache_arr_15__9, d_cache_arr_15__8, d_cache_arr_15__7, 
         d_cache_arr_15__6, d_cache_arr_15__5, d_cache_arr_15__4, 
         d_cache_arr_15__3, d_cache_arr_15__2, d_cache_arr_15__1, 
         d_cache_arr_15__0, d_cache_arr_16__31, d_cache_arr_16__30, 
         d_cache_arr_16__29, d_cache_arr_16__28, d_cache_arr_16__27, 
         d_cache_arr_16__26, d_cache_arr_16__25, d_cache_arr_16__24, 
         d_cache_arr_16__23, d_cache_arr_16__22, d_cache_arr_16__21, 
         d_cache_arr_16__20, d_cache_arr_16__19, d_cache_arr_16__18, 
         d_cache_arr_16__17, d_cache_arr_16__16, d_cache_arr_16__15, 
         d_cache_arr_16__14, d_cache_arr_16__13, d_cache_arr_16__12, 
         d_cache_arr_16__11, d_cache_arr_16__10, d_cache_arr_16__9, 
         d_cache_arr_16__8, d_cache_arr_16__7, d_cache_arr_16__6, 
         d_cache_arr_16__5, d_cache_arr_16__4, d_cache_arr_16__3, 
         d_cache_arr_16__2, d_cache_arr_16__1, d_cache_arr_16__0, 
         d_cache_arr_17__31, d_cache_arr_17__30, d_cache_arr_17__29, 
         d_cache_arr_17__28, d_cache_arr_17__27, d_cache_arr_17__26, 
         d_cache_arr_17__25, d_cache_arr_17__24, d_cache_arr_17__23, 
         d_cache_arr_17__22, d_cache_arr_17__21, d_cache_arr_17__20, 
         d_cache_arr_17__19, d_cache_arr_17__18, d_cache_arr_17__17, 
         d_cache_arr_17__16, d_cache_arr_17__15, d_cache_arr_17__14, 
         d_cache_arr_17__13, d_cache_arr_17__12, d_cache_arr_17__11, 
         d_cache_arr_17__10, d_cache_arr_17__9, d_cache_arr_17__8, 
         d_cache_arr_17__7, d_cache_arr_17__6, d_cache_arr_17__5, 
         d_cache_arr_17__4, d_cache_arr_17__3, d_cache_arr_17__2, 
         d_cache_arr_17__1, d_cache_arr_17__0, d_cache_arr_18__31, 
         d_cache_arr_18__30, d_cache_arr_18__29, d_cache_arr_18__28, 
         d_cache_arr_18__27, d_cache_arr_18__26, d_cache_arr_18__25, 
         d_cache_arr_18__24, d_cache_arr_18__23, d_cache_arr_18__22, 
         d_cache_arr_18__21, d_cache_arr_18__20, d_cache_arr_18__19, 
         d_cache_arr_18__18, d_cache_arr_18__17, d_cache_arr_18__16, 
         d_cache_arr_18__15, d_cache_arr_18__14, d_cache_arr_18__13, 
         d_cache_arr_18__12, d_cache_arr_18__11, d_cache_arr_18__10, 
         d_cache_arr_18__9, d_cache_arr_18__8, d_cache_arr_18__7, 
         d_cache_arr_18__6, d_cache_arr_18__5, d_cache_arr_18__4, 
         d_cache_arr_18__3, d_cache_arr_18__2, d_cache_arr_18__1, 
         d_cache_arr_18__0, d_cache_arr_19__31, d_cache_arr_19__30, 
         d_cache_arr_19__29, d_cache_arr_19__28, d_cache_arr_19__27, 
         d_cache_arr_19__26, d_cache_arr_19__25, d_cache_arr_19__24, 
         d_cache_arr_19__23, d_cache_arr_19__22, d_cache_arr_19__21, 
         d_cache_arr_19__20, d_cache_arr_19__19, d_cache_arr_19__18, 
         d_cache_arr_19__17, d_cache_arr_19__16, d_cache_arr_19__15, 
         d_cache_arr_19__14, d_cache_arr_19__13, d_cache_arr_19__12, 
         d_cache_arr_19__11, d_cache_arr_19__10, d_cache_arr_19__9, 
         d_cache_arr_19__8, d_cache_arr_19__7, d_cache_arr_19__6, 
         d_cache_arr_19__5, d_cache_arr_19__4, d_cache_arr_19__3, 
         d_cache_arr_19__2, d_cache_arr_19__1, d_cache_arr_19__0, 
         d_cache_arr_20__31, d_cache_arr_20__30, d_cache_arr_20__29, 
         d_cache_arr_20__28, d_cache_arr_20__27, d_cache_arr_20__26, 
         d_cache_arr_20__25, d_cache_arr_20__24, d_cache_arr_20__23, 
         d_cache_arr_20__22, d_cache_arr_20__21, d_cache_arr_20__20, 
         d_cache_arr_20__19, d_cache_arr_20__18, d_cache_arr_20__17, 
         d_cache_arr_20__16, d_cache_arr_20__15, d_cache_arr_20__14, 
         d_cache_arr_20__13, d_cache_arr_20__12, d_cache_arr_20__11, 
         d_cache_arr_20__10, d_cache_arr_20__9, d_cache_arr_20__8, 
         d_cache_arr_20__7, d_cache_arr_20__6, d_cache_arr_20__5, 
         d_cache_arr_20__4, d_cache_arr_20__3, d_cache_arr_20__2, 
         d_cache_arr_20__1, d_cache_arr_20__0, d_cache_arr_21__31, 
         d_cache_arr_21__30, d_cache_arr_21__29, d_cache_arr_21__28, 
         d_cache_arr_21__27, d_cache_arr_21__26, d_cache_arr_21__25, 
         d_cache_arr_21__24, d_cache_arr_21__23, d_cache_arr_21__22, 
         d_cache_arr_21__21, d_cache_arr_21__20, d_cache_arr_21__19, 
         d_cache_arr_21__18, d_cache_arr_21__17, d_cache_arr_21__16, 
         d_cache_arr_21__15, d_cache_arr_21__14, d_cache_arr_21__13, 
         d_cache_arr_21__12, d_cache_arr_21__11, d_cache_arr_21__10, 
         d_cache_arr_21__9, d_cache_arr_21__8, d_cache_arr_21__7, 
         d_cache_arr_21__6, d_cache_arr_21__5, d_cache_arr_21__4, 
         d_cache_arr_21__3, d_cache_arr_21__2, d_cache_arr_21__1, 
         d_cache_arr_21__0, d_cache_arr_22__31, d_cache_arr_22__30, 
         d_cache_arr_22__29, d_cache_arr_22__28, d_cache_arr_22__27, 
         d_cache_arr_22__26, d_cache_arr_22__25, d_cache_arr_22__24, 
         d_cache_arr_22__23, d_cache_arr_22__22, d_cache_arr_22__21, 
         d_cache_arr_22__20, d_cache_arr_22__19, d_cache_arr_22__18, 
         d_cache_arr_22__17, d_cache_arr_22__16, d_cache_arr_22__15, 
         d_cache_arr_22__14, d_cache_arr_22__13, d_cache_arr_22__12, 
         d_cache_arr_22__11, d_cache_arr_22__10, d_cache_arr_22__9, 
         d_cache_arr_22__8, d_cache_arr_22__7, d_cache_arr_22__6, 
         d_cache_arr_22__5, d_cache_arr_22__4, d_cache_arr_22__3, 
         d_cache_arr_22__2, d_cache_arr_22__1, d_cache_arr_22__0, 
         d_cache_arr_23__31, d_cache_arr_23__30, d_cache_arr_23__29, 
         d_cache_arr_23__28, d_cache_arr_23__27, d_cache_arr_23__26, 
         d_cache_arr_23__25, d_cache_arr_23__24, d_cache_arr_23__23, 
         d_cache_arr_23__22, d_cache_arr_23__21, d_cache_arr_23__20, 
         d_cache_arr_23__19, d_cache_arr_23__18, d_cache_arr_23__17, 
         d_cache_arr_23__16, d_cache_arr_23__15, d_cache_arr_23__14, 
         d_cache_arr_23__13, d_cache_arr_23__12, d_cache_arr_23__11, 
         d_cache_arr_23__10, d_cache_arr_23__9, d_cache_arr_23__8, 
         d_cache_arr_23__7, d_cache_arr_23__6, d_cache_arr_23__5, 
         d_cache_arr_23__4, d_cache_arr_23__3, d_cache_arr_23__2, 
         d_cache_arr_23__1, d_cache_arr_23__0, d_cache_arr_24__31, 
         d_cache_arr_24__30, d_cache_arr_24__29, d_cache_arr_24__28, 
         d_cache_arr_24__27, d_cache_arr_24__26, d_cache_arr_24__25, 
         d_cache_arr_24__24, d_cache_arr_24__23, d_cache_arr_24__22, 
         d_cache_arr_24__21, d_cache_arr_24__20, d_cache_arr_24__19, 
         d_cache_arr_24__18, d_cache_arr_24__17, d_cache_arr_24__16, 
         d_cache_arr_24__15, d_cache_arr_24__14, d_cache_arr_24__13, 
         d_cache_arr_24__12, d_cache_arr_24__11, d_cache_arr_24__10, 
         d_cache_arr_24__9, d_cache_arr_24__8, d_cache_arr_24__7, 
         d_cache_arr_24__6, d_cache_arr_24__5, d_cache_arr_24__4, 
         d_cache_arr_24__3, d_cache_arr_24__2, d_cache_arr_24__1, 
         d_cache_arr_24__0, q_cache_arr_0__31, q_cache_arr_0__30, 
         q_cache_arr_0__29, q_cache_arr_0__28, q_cache_arr_0__27, 
         q_cache_arr_0__26, q_cache_arr_0__25, q_cache_arr_0__24, 
         q_cache_arr_0__23, q_cache_arr_0__22, q_cache_arr_0__21, 
         q_cache_arr_0__20, q_cache_arr_0__19, q_cache_arr_0__18, 
         q_cache_arr_0__17, q_cache_arr_0__16, q_cache_arr_0__15, 
         q_cache_arr_0__14, q_cache_arr_0__13, q_cache_arr_0__12, 
         q_cache_arr_0__11, q_cache_arr_0__10, q_cache_arr_0__9, 
         q_cache_arr_0__8, q_cache_arr_0__7, q_cache_arr_0__6, q_cache_arr_0__5, 
         q_cache_arr_0__4, q_cache_arr_0__3, q_cache_arr_0__2, q_cache_arr_0__1, 
         q_cache_arr_0__0, q_cache_arr_1__31, q_cache_arr_1__30, 
         q_cache_arr_1__29, q_cache_arr_1__28, q_cache_arr_1__27, 
         q_cache_arr_1__26, q_cache_arr_1__25, q_cache_arr_1__24, 
         q_cache_arr_1__23, q_cache_arr_1__22, q_cache_arr_1__21, 
         q_cache_arr_1__20, q_cache_arr_1__19, q_cache_arr_1__18, 
         q_cache_arr_1__17, q_cache_arr_1__16, q_cache_arr_1__15, 
         q_cache_arr_1__14, q_cache_arr_1__13, q_cache_arr_1__12, 
         q_cache_arr_1__11, q_cache_arr_1__10, q_cache_arr_1__9, 
         q_cache_arr_1__8, q_cache_arr_1__7, q_cache_arr_1__6, q_cache_arr_1__5, 
         q_cache_arr_1__4, q_cache_arr_1__3, q_cache_arr_1__2, q_cache_arr_1__1, 
         q_cache_arr_1__0, q_cache_arr_2__31, q_cache_arr_2__30, 
         q_cache_arr_2__29, q_cache_arr_2__28, q_cache_arr_2__27, 
         q_cache_arr_2__26, q_cache_arr_2__25, q_cache_arr_2__24, 
         q_cache_arr_2__23, q_cache_arr_2__22, q_cache_arr_2__21, 
         q_cache_arr_2__20, q_cache_arr_2__19, q_cache_arr_2__18, 
         q_cache_arr_2__17, q_cache_arr_2__16, q_cache_arr_2__15, 
         q_cache_arr_2__14, q_cache_arr_2__13, q_cache_arr_2__12, 
         q_cache_arr_2__11, q_cache_arr_2__10, q_cache_arr_2__9, 
         q_cache_arr_2__8, q_cache_arr_2__7, q_cache_arr_2__6, q_cache_arr_2__5, 
         q_cache_arr_2__4, q_cache_arr_2__3, q_cache_arr_2__2, q_cache_arr_2__1, 
         q_cache_arr_2__0, q_cache_arr_3__31, q_cache_arr_3__30, 
         q_cache_arr_3__29, q_cache_arr_3__28, q_cache_arr_3__27, 
         q_cache_arr_3__26, q_cache_arr_3__25, q_cache_arr_3__24, 
         q_cache_arr_3__23, q_cache_arr_3__22, q_cache_arr_3__21, 
         q_cache_arr_3__20, q_cache_arr_3__19, q_cache_arr_3__18, 
         q_cache_arr_3__17, q_cache_arr_3__16, q_cache_arr_3__15, 
         q_cache_arr_3__14, q_cache_arr_3__13, q_cache_arr_3__12, 
         q_cache_arr_3__11, q_cache_arr_3__10, q_cache_arr_3__9, 
         q_cache_arr_3__8, q_cache_arr_3__7, q_cache_arr_3__6, q_cache_arr_3__5, 
         q_cache_arr_3__4, q_cache_arr_3__3, q_cache_arr_3__2, q_cache_arr_3__1, 
         q_cache_arr_3__0, q_cache_arr_4__31, q_cache_arr_4__30, 
         q_cache_arr_4__29, q_cache_arr_4__28, q_cache_arr_4__27, 
         q_cache_arr_4__26, q_cache_arr_4__25, q_cache_arr_4__24, 
         q_cache_arr_4__23, q_cache_arr_4__22, q_cache_arr_4__21, 
         q_cache_arr_4__20, q_cache_arr_4__19, q_cache_arr_4__18, 
         q_cache_arr_4__17, q_cache_arr_4__16, q_cache_arr_4__15, 
         q_cache_arr_4__14, q_cache_arr_4__13, q_cache_arr_4__12, 
         q_cache_arr_4__11, q_cache_arr_4__10, q_cache_arr_4__9, 
         q_cache_arr_4__8, q_cache_arr_4__7, q_cache_arr_4__6, q_cache_arr_4__5, 
         q_cache_arr_4__4, q_cache_arr_4__3, q_cache_arr_4__2, q_cache_arr_4__1, 
         q_cache_arr_4__0, q_cache_arr_5__31, q_cache_arr_5__30, 
         q_cache_arr_5__29, q_cache_arr_5__28, q_cache_arr_5__27, 
         q_cache_arr_5__26, q_cache_arr_5__25, q_cache_arr_5__24, 
         q_cache_arr_5__23, q_cache_arr_5__22, q_cache_arr_5__21, 
         q_cache_arr_5__20, q_cache_arr_5__19, q_cache_arr_5__18, 
         q_cache_arr_5__17, q_cache_arr_5__16, q_cache_arr_5__15, 
         q_cache_arr_5__14, q_cache_arr_5__13, q_cache_arr_5__12, 
         q_cache_arr_5__11, q_cache_arr_5__10, q_cache_arr_5__9, 
         q_cache_arr_5__8, q_cache_arr_5__7, q_cache_arr_5__6, q_cache_arr_5__5, 
         q_cache_arr_5__4, q_cache_arr_5__3, q_cache_arr_5__2, q_cache_arr_5__1, 
         q_cache_arr_5__0, q_cache_arr_6__31, q_cache_arr_6__30, 
         q_cache_arr_6__29, q_cache_arr_6__28, q_cache_arr_6__27, 
         q_cache_arr_6__26, q_cache_arr_6__25, q_cache_arr_6__24, 
         q_cache_arr_6__23, q_cache_arr_6__22, q_cache_arr_6__21, 
         q_cache_arr_6__20, q_cache_arr_6__19, q_cache_arr_6__18, 
         q_cache_arr_6__17, q_cache_arr_6__16, q_cache_arr_6__15, 
         q_cache_arr_6__14, q_cache_arr_6__13, q_cache_arr_6__12, 
         q_cache_arr_6__11, q_cache_arr_6__10, q_cache_arr_6__9, 
         q_cache_arr_6__8, q_cache_arr_6__7, q_cache_arr_6__6, q_cache_arr_6__5, 
         q_cache_arr_6__4, q_cache_arr_6__3, q_cache_arr_6__2, q_cache_arr_6__1, 
         q_cache_arr_6__0, q_cache_arr_7__31, q_cache_arr_7__30, 
         q_cache_arr_7__29, q_cache_arr_7__28, q_cache_arr_7__27, 
         q_cache_arr_7__26, q_cache_arr_7__25, q_cache_arr_7__24, 
         q_cache_arr_7__23, q_cache_arr_7__22, q_cache_arr_7__21, 
         q_cache_arr_7__20, q_cache_arr_7__19, q_cache_arr_7__18, 
         q_cache_arr_7__17, q_cache_arr_7__16, q_cache_arr_7__15, 
         q_cache_arr_7__14, q_cache_arr_7__13, q_cache_arr_7__12, 
         q_cache_arr_7__11, q_cache_arr_7__10, q_cache_arr_7__9, 
         q_cache_arr_7__8, q_cache_arr_7__7, q_cache_arr_7__6, q_cache_arr_7__5, 
         q_cache_arr_7__4, q_cache_arr_7__3, q_cache_arr_7__2, q_cache_arr_7__1, 
         q_cache_arr_7__0, q_cache_arr_8__31, q_cache_arr_8__30, 
         q_cache_arr_8__29, q_cache_arr_8__28, q_cache_arr_8__27, 
         q_cache_arr_8__26, q_cache_arr_8__25, q_cache_arr_8__24, 
         q_cache_arr_8__23, q_cache_arr_8__22, q_cache_arr_8__21, 
         q_cache_arr_8__20, q_cache_arr_8__19, q_cache_arr_8__18, 
         q_cache_arr_8__17, q_cache_arr_8__16, q_cache_arr_8__15, 
         q_cache_arr_8__14, q_cache_arr_8__13, q_cache_arr_8__12, 
         q_cache_arr_8__11, q_cache_arr_8__10, q_cache_arr_8__9, 
         q_cache_arr_8__8, q_cache_arr_8__7, q_cache_arr_8__6, q_cache_arr_8__5, 
         q_cache_arr_8__4, q_cache_arr_8__3, q_cache_arr_8__2, q_cache_arr_8__1, 
         q_cache_arr_8__0, q_cache_arr_9__31, q_cache_arr_9__30, 
         q_cache_arr_9__29, q_cache_arr_9__28, q_cache_arr_9__27, 
         q_cache_arr_9__26, q_cache_arr_9__25, q_cache_arr_9__24, 
         q_cache_arr_9__23, q_cache_arr_9__22, q_cache_arr_9__21, 
         q_cache_arr_9__20, q_cache_arr_9__19, q_cache_arr_9__18, 
         q_cache_arr_9__17, q_cache_arr_9__16, q_cache_arr_9__15, 
         q_cache_arr_9__14, q_cache_arr_9__13, q_cache_arr_9__12, 
         q_cache_arr_9__11, q_cache_arr_9__10, q_cache_arr_9__9, 
         q_cache_arr_9__8, q_cache_arr_9__7, q_cache_arr_9__6, q_cache_arr_9__5, 
         q_cache_arr_9__4, q_cache_arr_9__3, q_cache_arr_9__2, q_cache_arr_9__1, 
         q_cache_arr_9__0, q_cache_arr_10__31, q_cache_arr_10__30, 
         q_cache_arr_10__29, q_cache_arr_10__28, q_cache_arr_10__27, 
         q_cache_arr_10__26, q_cache_arr_10__25, q_cache_arr_10__24, 
         q_cache_arr_10__23, q_cache_arr_10__22, q_cache_arr_10__21, 
         q_cache_arr_10__20, q_cache_arr_10__19, q_cache_arr_10__18, 
         q_cache_arr_10__17, q_cache_arr_10__16, q_cache_arr_10__15, 
         q_cache_arr_10__14, q_cache_arr_10__13, q_cache_arr_10__12, 
         q_cache_arr_10__11, q_cache_arr_10__10, q_cache_arr_10__9, 
         q_cache_arr_10__8, q_cache_arr_10__7, q_cache_arr_10__6, 
         q_cache_arr_10__5, q_cache_arr_10__4, q_cache_arr_10__3, 
         q_cache_arr_10__2, q_cache_arr_10__1, q_cache_arr_10__0, 
         q_cache_arr_11__31, q_cache_arr_11__30, q_cache_arr_11__29, 
         q_cache_arr_11__28, q_cache_arr_11__27, q_cache_arr_11__26, 
         q_cache_arr_11__25, q_cache_arr_11__24, q_cache_arr_11__23, 
         q_cache_arr_11__22, q_cache_arr_11__21, q_cache_arr_11__20, 
         q_cache_arr_11__19, q_cache_arr_11__18, q_cache_arr_11__17, 
         q_cache_arr_11__16, q_cache_arr_11__15, q_cache_arr_11__14, 
         q_cache_arr_11__13, q_cache_arr_11__12, q_cache_arr_11__11, 
         q_cache_arr_11__10, q_cache_arr_11__9, q_cache_arr_11__8, 
         q_cache_arr_11__7, q_cache_arr_11__6, q_cache_arr_11__5, 
         q_cache_arr_11__4, q_cache_arr_11__3, q_cache_arr_11__2, 
         q_cache_arr_11__1, q_cache_arr_11__0, q_cache_arr_12__31, 
         q_cache_arr_12__30, q_cache_arr_12__29, q_cache_arr_12__28, 
         q_cache_arr_12__27, q_cache_arr_12__26, q_cache_arr_12__25, 
         q_cache_arr_12__24, q_cache_arr_12__23, q_cache_arr_12__22, 
         q_cache_arr_12__21, q_cache_arr_12__20, q_cache_arr_12__19, 
         q_cache_arr_12__18, q_cache_arr_12__17, q_cache_arr_12__16, 
         q_cache_arr_12__15, q_cache_arr_12__14, q_cache_arr_12__13, 
         q_cache_arr_12__12, q_cache_arr_12__11, q_cache_arr_12__10, 
         q_cache_arr_12__9, q_cache_arr_12__8, q_cache_arr_12__7, 
         q_cache_arr_12__6, q_cache_arr_12__5, q_cache_arr_12__4, 
         q_cache_arr_12__3, q_cache_arr_12__2, q_cache_arr_12__1, 
         q_cache_arr_12__0, q_cache_arr_13__31, q_cache_arr_13__30, 
         q_cache_arr_13__29, q_cache_arr_13__28, q_cache_arr_13__27, 
         q_cache_arr_13__26, q_cache_arr_13__25, q_cache_arr_13__24, 
         q_cache_arr_13__23, q_cache_arr_13__22, q_cache_arr_13__21, 
         q_cache_arr_13__20, q_cache_arr_13__19, q_cache_arr_13__18, 
         q_cache_arr_13__17, q_cache_arr_13__16, q_cache_arr_13__15, 
         q_cache_arr_13__14, q_cache_arr_13__13, q_cache_arr_13__12, 
         q_cache_arr_13__11, q_cache_arr_13__10, q_cache_arr_13__9, 
         q_cache_arr_13__8, q_cache_arr_13__7, q_cache_arr_13__6, 
         q_cache_arr_13__5, q_cache_arr_13__4, q_cache_arr_13__3, 
         q_cache_arr_13__2, q_cache_arr_13__1, q_cache_arr_13__0, 
         q_cache_arr_14__31, q_cache_arr_14__30, q_cache_arr_14__29, 
         q_cache_arr_14__28, q_cache_arr_14__27, q_cache_arr_14__26, 
         q_cache_arr_14__25, q_cache_arr_14__24, q_cache_arr_14__23, 
         q_cache_arr_14__22, q_cache_arr_14__21, q_cache_arr_14__20, 
         q_cache_arr_14__19, q_cache_arr_14__18, q_cache_arr_14__17, 
         q_cache_arr_14__16, q_cache_arr_14__15, q_cache_arr_14__14, 
         q_cache_arr_14__13, q_cache_arr_14__12, q_cache_arr_14__11, 
         q_cache_arr_14__10, q_cache_arr_14__9, q_cache_arr_14__8, 
         q_cache_arr_14__7, q_cache_arr_14__6, q_cache_arr_14__5, 
         q_cache_arr_14__4, q_cache_arr_14__3, q_cache_arr_14__2, 
         q_cache_arr_14__1, q_cache_arr_14__0, q_cache_arr_15__31, 
         q_cache_arr_15__30, q_cache_arr_15__29, q_cache_arr_15__28, 
         q_cache_arr_15__27, q_cache_arr_15__26, q_cache_arr_15__25, 
         q_cache_arr_15__24, q_cache_arr_15__23, q_cache_arr_15__22, 
         q_cache_arr_15__21, q_cache_arr_15__20, q_cache_arr_15__19, 
         q_cache_arr_15__18, q_cache_arr_15__17, q_cache_arr_15__16, 
         q_cache_arr_15__15, q_cache_arr_15__14, q_cache_arr_15__13, 
         q_cache_arr_15__12, q_cache_arr_15__11, q_cache_arr_15__10, 
         q_cache_arr_15__9, q_cache_arr_15__8, q_cache_arr_15__7, 
         q_cache_arr_15__6, q_cache_arr_15__5, q_cache_arr_15__4, 
         q_cache_arr_15__3, q_cache_arr_15__2, q_cache_arr_15__1, 
         q_cache_arr_15__0, q_cache_arr_16__31, q_cache_arr_16__30, 
         q_cache_arr_16__29, q_cache_arr_16__28, q_cache_arr_16__27, 
         q_cache_arr_16__26, q_cache_arr_16__25, q_cache_arr_16__24, 
         q_cache_arr_16__23, q_cache_arr_16__22, q_cache_arr_16__21, 
         q_cache_arr_16__20, q_cache_arr_16__19, q_cache_arr_16__18, 
         q_cache_arr_16__17, q_cache_arr_16__16, q_cache_arr_16__15, 
         q_cache_arr_16__14, q_cache_arr_16__13, q_cache_arr_16__12, 
         q_cache_arr_16__11, q_cache_arr_16__10, q_cache_arr_16__9, 
         q_cache_arr_16__8, q_cache_arr_16__7, q_cache_arr_16__6, 
         q_cache_arr_16__5, q_cache_arr_16__4, q_cache_arr_16__3, 
         q_cache_arr_16__2, q_cache_arr_16__1, q_cache_arr_16__0, 
         q_cache_arr_17__31, q_cache_arr_17__30, q_cache_arr_17__29, 
         q_cache_arr_17__28, q_cache_arr_17__27, q_cache_arr_17__26, 
         q_cache_arr_17__25, q_cache_arr_17__24, q_cache_arr_17__23, 
         q_cache_arr_17__22, q_cache_arr_17__21, q_cache_arr_17__20, 
         q_cache_arr_17__19, q_cache_arr_17__18, q_cache_arr_17__17, 
         q_cache_arr_17__16, q_cache_arr_17__15, q_cache_arr_17__14, 
         q_cache_arr_17__13, q_cache_arr_17__12, q_cache_arr_17__11, 
         q_cache_arr_17__10, q_cache_arr_17__9, q_cache_arr_17__8, 
         q_cache_arr_17__7, q_cache_arr_17__6, q_cache_arr_17__5, 
         q_cache_arr_17__4, q_cache_arr_17__3, q_cache_arr_17__2, 
         q_cache_arr_17__1, q_cache_arr_17__0, q_cache_arr_18__31, 
         q_cache_arr_18__30, q_cache_arr_18__29, q_cache_arr_18__28, 
         q_cache_arr_18__27, q_cache_arr_18__26, q_cache_arr_18__25, 
         q_cache_arr_18__24, q_cache_arr_18__23, q_cache_arr_18__22, 
         q_cache_arr_18__21, q_cache_arr_18__20, q_cache_arr_18__19, 
         q_cache_arr_18__18, q_cache_arr_18__17, q_cache_arr_18__16, 
         q_cache_arr_18__15, q_cache_arr_18__14, q_cache_arr_18__13, 
         q_cache_arr_18__12, q_cache_arr_18__11, q_cache_arr_18__10, 
         q_cache_arr_18__9, q_cache_arr_18__8, q_cache_arr_18__7, 
         q_cache_arr_18__6, q_cache_arr_18__5, q_cache_arr_18__4, 
         q_cache_arr_18__3, q_cache_arr_18__2, q_cache_arr_18__1, 
         q_cache_arr_18__0, q_cache_arr_19__31, q_cache_arr_19__30, 
         q_cache_arr_19__29, q_cache_arr_19__28, q_cache_arr_19__27, 
         q_cache_arr_19__26, q_cache_arr_19__25, q_cache_arr_19__24, 
         q_cache_arr_19__23, q_cache_arr_19__22, q_cache_arr_19__21, 
         q_cache_arr_19__20, q_cache_arr_19__19, q_cache_arr_19__18, 
         q_cache_arr_19__17, q_cache_arr_19__16, q_cache_arr_19__15, 
         q_cache_arr_19__14, q_cache_arr_19__13, q_cache_arr_19__12, 
         q_cache_arr_19__11, q_cache_arr_19__10, q_cache_arr_19__9, 
         q_cache_arr_19__8, q_cache_arr_19__7, q_cache_arr_19__6, 
         q_cache_arr_19__5, q_cache_arr_19__4, q_cache_arr_19__3, 
         q_cache_arr_19__2, q_cache_arr_19__1, q_cache_arr_19__0, 
         q_cache_arr_20__31, q_cache_arr_20__30, q_cache_arr_20__29, 
         q_cache_arr_20__28, q_cache_arr_20__27, q_cache_arr_20__26, 
         q_cache_arr_20__25, q_cache_arr_20__24, q_cache_arr_20__23, 
         q_cache_arr_20__22, q_cache_arr_20__21, q_cache_arr_20__20, 
         q_cache_arr_20__19, q_cache_arr_20__18, q_cache_arr_20__17, 
         q_cache_arr_20__16, q_cache_arr_20__15, q_cache_arr_20__14, 
         q_cache_arr_20__13, q_cache_arr_20__12, q_cache_arr_20__11, 
         q_cache_arr_20__10, q_cache_arr_20__9, q_cache_arr_20__8, 
         q_cache_arr_20__7, q_cache_arr_20__6, q_cache_arr_20__5, 
         q_cache_arr_20__4, q_cache_arr_20__3, q_cache_arr_20__2, 
         q_cache_arr_20__1, q_cache_arr_20__0, q_cache_arr_21__31, 
         q_cache_arr_21__30, q_cache_arr_21__29, q_cache_arr_21__28, 
         q_cache_arr_21__27, q_cache_arr_21__26, q_cache_arr_21__25, 
         q_cache_arr_21__24, q_cache_arr_21__23, q_cache_arr_21__22, 
         q_cache_arr_21__21, q_cache_arr_21__20, q_cache_arr_21__19, 
         q_cache_arr_21__18, q_cache_arr_21__17, q_cache_arr_21__16, 
         q_cache_arr_21__15, q_cache_arr_21__14, q_cache_arr_21__13, 
         q_cache_arr_21__12, q_cache_arr_21__11, q_cache_arr_21__10, 
         q_cache_arr_21__9, q_cache_arr_21__8, q_cache_arr_21__7, 
         q_cache_arr_21__6, q_cache_arr_21__5, q_cache_arr_21__4, 
         q_cache_arr_21__3, q_cache_arr_21__2, q_cache_arr_21__1, 
         q_cache_arr_21__0, q_cache_arr_22__31, q_cache_arr_22__30, 
         q_cache_arr_22__29, q_cache_arr_22__28, q_cache_arr_22__27, 
         q_cache_arr_22__26, q_cache_arr_22__25, q_cache_arr_22__24, 
         q_cache_arr_22__23, q_cache_arr_22__22, q_cache_arr_22__21, 
         q_cache_arr_22__20, q_cache_arr_22__19, q_cache_arr_22__18, 
         q_cache_arr_22__17, q_cache_arr_22__16, q_cache_arr_22__15, 
         q_cache_arr_22__14, q_cache_arr_22__13, q_cache_arr_22__12, 
         q_cache_arr_22__11, q_cache_arr_22__10, q_cache_arr_22__9, 
         q_cache_arr_22__8, q_cache_arr_22__7, q_cache_arr_22__6, 
         q_cache_arr_22__5, q_cache_arr_22__4, q_cache_arr_22__3, 
         q_cache_arr_22__2, q_cache_arr_22__1, q_cache_arr_22__0, 
         q_cache_arr_23__31, q_cache_arr_23__30, q_cache_arr_23__29, 
         q_cache_arr_23__28, q_cache_arr_23__27, q_cache_arr_23__26, 
         q_cache_arr_23__25, q_cache_arr_23__24, q_cache_arr_23__23, 
         q_cache_arr_23__22, q_cache_arr_23__21, q_cache_arr_23__20, 
         q_cache_arr_23__19, q_cache_arr_23__18, q_cache_arr_23__17, 
         q_cache_arr_23__16, q_cache_arr_23__15, q_cache_arr_23__14, 
         q_cache_arr_23__13, q_cache_arr_23__12, q_cache_arr_23__11, 
         q_cache_arr_23__10, q_cache_arr_23__9, q_cache_arr_23__8, 
         q_cache_arr_23__7, q_cache_arr_23__6, q_cache_arr_23__5, 
         q_cache_arr_23__4, q_cache_arr_23__3, q_cache_arr_23__2, 
         q_cache_arr_23__1, q_cache_arr_23__0, q_cache_arr_24__31, 
         q_cache_arr_24__30, q_cache_arr_24__29, q_cache_arr_24__28, 
         q_cache_arr_24__27, q_cache_arr_24__26, q_cache_arr_24__25, 
         q_cache_arr_24__24, q_cache_arr_24__23, q_cache_arr_24__22, 
         q_cache_arr_24__21, q_cache_arr_24__20, q_cache_arr_24__19, 
         q_cache_arr_24__18, q_cache_arr_24__17, q_cache_arr_24__16, 
         q_cache_arr_24__15, q_cache_arr_24__14, q_cache_arr_24__13, 
         q_cache_arr_24__12, q_cache_arr_24__11, q_cache_arr_24__10, 
         q_cache_arr_24__9, q_cache_arr_24__8, q_cache_arr_24__7, 
         q_cache_arr_24__6, q_cache_arr_24__5, q_cache_arr_24__4, 
         q_cache_arr_24__3, q_cache_arr_24__2, q_cache_arr_24__1, 
         q_cache_arr_24__0, img_load_tmp, filter_load_tmp, ready_tmp, 
         buffer_ready_tmp, comp_pipe_rst, comp_pipe_en, output1_init_q_15, 
         output1_init_q_14, output1_init_q_13, output1_init_q_12, 
         output1_init_q_11, output1_init_q_10, output1_init_q_9, 
         output1_init_q_8, output1_init_q_7, output1_init_q_6, output1_init_q_5, 
         output1_init_q_4, output1_init_q_3, output1_init_q_2, output1_init_q_1, 
         output1_init_q_0, output2_init_q_15, output2_init_q_14, 
         output2_init_q_13, output2_init_q_12, output2_init_q_11, 
         output2_init_q_10, output2_init_q_9, output2_init_q_8, output2_init_q_7, 
         output2_init_q_6, output2_init_q_5, output2_init_q_4, output2_init_q_3, 
         output2_init_q_2, output2_init_q_1, output2_init_q_0, filter_size_q, 
         operation_q, compute_relu_q, semi_ready, nx4, nx10, NOT_nx4, 
         buffer_ready_dup0, nx302, nx201, nx211, nx221, nx231, nx241, nx251, 
         nx261, nx271, nx281, nx291, nx301, nx311, nx321, nx331, nx341, nx351, 
         nx361, nx371, nx381, nx391, nx401, nx411, nx421, nx431, nx441, nx451, 
         nx461, nx471, nx481, nx491, nx501, nx511, nx521, nx531, nx541, nx551, 
         nx561, nx571, nx581, nx591, nx601, nx611, nx621, nx631, nx641, nx651, 
         nx661, nx671, nx681, nx691, nx701, nx711, nx721, nx731, nx741, nx751, 
         nx761, nx771, nx781, nx791, nx801, nx811, nx821, nx831, nx841, nx851, 
         nx861, nx875, nx879, nx996, nx1103, nx1105, nx1107, nx1109, nx1111, 
         nx1113, nx1115, nx1117, nx1119, nx1121, nx1131, nx1133, nx1137, nx1139, 
         nx1141, nx1143, nx1145, nx1147, nx1151, nx1161, nx1167, nx1169, nx1171, 
         nx1173, nx1175, nx1177, nx1179, nx1181, nx1183, nx1185, nx1187, nx1189, 
         nx1191, nx1193, nx1195;
    wire [70:0] \$dummy ;




    ComputationPipeline gen_comp_pipeline (.img_data_0__15 (img_data_0__15), .img_data_0__14 (
                        img_data_0__14), .img_data_0__13 (img_data_0__13), .img_data_0__12 (
                        img_data_0__12), .img_data_0__11 (img_data_0__11), .img_data_0__10 (
                        img_data_0__10), .img_data_0__9 (img_data_0__9), .img_data_0__8 (
                        img_data_0__8), .img_data_0__7 (img_data_0__7), .img_data_0__6 (
                        img_data_0__6), .img_data_0__5 (img_data_0__5), .img_data_0__4 (
                        img_data_0__4), .img_data_0__3 (img_data_0__3), .img_data_0__2 (
                        img_data_0__2), .img_data_0__1 (img_data_0__1), .img_data_0__0 (
                        img_data_0__0), .img_data_1__15 (nx1103), .img_data_1__14 (
                        img_data_1__14), .img_data_1__13 (img_data_1__13), .img_data_1__12 (
                        img_data_1__12), .img_data_1__11 (img_data_1__11), .img_data_1__10 (
                        img_data_1__10), .img_data_1__9 (img_data_1__9), .img_data_1__8 (
                        img_data_1__8), .img_data_1__7 (img_data_1__7), .img_data_1__6 (
                        img_data_1__6), .img_data_1__5 (img_data_1__5), .img_data_1__4 (
                        img_data_1__4), .img_data_1__3 (img_data_1__3), .img_data_1__2 (
                        img_data_1__2), .img_data_1__1 (img_data_1__1), .img_data_1__0 (
                        img_data_1__0), .img_data_2__15 (nx1105), .img_data_2__14 (
                        img_data_2__14), .img_data_2__13 (img_data_2__13), .img_data_2__12 (
                        img_data_2__12), .img_data_2__11 (img_data_2__11), .img_data_2__10 (
                        img_data_2__10), .img_data_2__9 (img_data_2__9), .img_data_2__8 (
                        img_data_2__8), .img_data_2__7 (img_data_2__7), .img_data_2__6 (
                        img_data_2__6), .img_data_2__5 (img_data_2__5), .img_data_2__4 (
                        img_data_2__4), .img_data_2__3 (img_data_2__3), .img_data_2__2 (
                        img_data_2__2), .img_data_2__1 (img_data_2__1), .img_data_2__0 (
                        img_data_2__0), .img_data_3__15 (img_data_3__15), .img_data_3__14 (
                        img_data_3__14), .img_data_3__13 (img_data_3__13), .img_data_3__12 (
                        img_data_3__12), .img_data_3__11 (img_data_3__11), .img_data_3__10 (
                        img_data_3__10), .img_data_3__9 (img_data_3__9), .img_data_3__8 (
                        img_data_3__8), .img_data_3__7 (img_data_3__7), .img_data_3__6 (
                        img_data_3__6), .img_data_3__5 (img_data_3__5), .img_data_3__4 (
                        img_data_3__4), .img_data_3__3 (img_data_3__3), .img_data_3__2 (
                        img_data_3__2), .img_data_3__1 (img_data_3__1), .img_data_3__0 (
                        img_data_3__0), .img_data_4__15 (img_data_4__15), .img_data_4__14 (
                        img_data_4__14), .img_data_4__13 (img_data_4__13), .img_data_4__12 (
                        img_data_4__12), .img_data_4__11 (img_data_4__11), .img_data_4__10 (
                        img_data_4__10), .img_data_4__9 (img_data_4__9), .img_data_4__8 (
                        img_data_4__8), .img_data_4__7 (img_data_4__7), .img_data_4__6 (
                        img_data_4__6), .img_data_4__5 (img_data_4__5), .img_data_4__4 (
                        img_data_4__4), .img_data_4__3 (img_data_4__3), .img_data_4__2 (
                        img_data_4__2), .img_data_4__1 (img_data_4__1), .img_data_4__0 (
                        img_data_4__0), .img_data_5__15 (img_data_5__15), .img_data_5__14 (
                        img_data_5__14), .img_data_5__13 (img_data_5__13), .img_data_5__12 (
                        img_data_5__12), .img_data_5__11 (img_data_5__11), .img_data_5__10 (
                        img_data_5__10), .img_data_5__9 (img_data_5__9), .img_data_5__8 (
                        img_data_5__8), .img_data_5__7 (img_data_5__7), .img_data_5__6 (
                        img_data_5__6), .img_data_5__5 (img_data_5__5), .img_data_5__4 (
                        img_data_5__4), .img_data_5__3 (img_data_5__3), .img_data_5__2 (
                        img_data_5__2), .img_data_5__1 (img_data_5__1), .img_data_5__0 (
                        img_data_5__0), .img_data_6__15 (nx1107), .img_data_6__14 (
                        img_data_6__14), .img_data_6__13 (img_data_6__13), .img_data_6__12 (
                        img_data_6__12), .img_data_6__11 (img_data_6__11), .img_data_6__10 (
                        img_data_6__10), .img_data_6__9 (img_data_6__9), .img_data_6__8 (
                        img_data_6__8), .img_data_6__7 (img_data_6__7), .img_data_6__6 (
                        img_data_6__6), .img_data_6__5 (img_data_6__5), .img_data_6__4 (
                        img_data_6__4), .img_data_6__3 (img_data_6__3), .img_data_6__2 (
                        img_data_6__2), .img_data_6__1 (img_data_6__1), .img_data_6__0 (
                        img_data_6__0), .img_data_7__15 (img_data_7__15), .img_data_7__14 (
                        img_data_7__14), .img_data_7__13 (img_data_7__13), .img_data_7__12 (
                        img_data_7__12), .img_data_7__11 (img_data_7__11), .img_data_7__10 (
                        img_data_7__10), .img_data_7__9 (img_data_7__9), .img_data_7__8 (
                        img_data_7__8), .img_data_7__7 (img_data_7__7), .img_data_7__6 (
                        img_data_7__6), .img_data_7__5 (img_data_7__5), .img_data_7__4 (
                        img_data_7__4), .img_data_7__3 (img_data_7__3), .img_data_7__2 (
                        img_data_7__2), .img_data_7__1 (img_data_7__1), .img_data_7__0 (
                        img_data_7__0), .img_data_8__15 (img_data_8__15), .img_data_8__14 (
                        img_data_8__14), .img_data_8__13 (img_data_8__13), .img_data_8__12 (
                        img_data_8__12), .img_data_8__11 (img_data_8__11), .img_data_8__10 (
                        img_data_8__10), .img_data_8__9 (img_data_8__9), .img_data_8__8 (
                        img_data_8__8), .img_data_8__7 (img_data_8__7), .img_data_8__6 (
                        img_data_8__6), .img_data_8__5 (img_data_8__5), .img_data_8__4 (
                        img_data_8__4), .img_data_8__3 (img_data_8__3), .img_data_8__2 (
                        img_data_8__2), .img_data_8__1 (img_data_8__1), .img_data_8__0 (
                        img_data_8__0), .img_data_9__15 (img_data_9__15), .img_data_9__14 (
                        img_data_9__14), .img_data_9__13 (img_data_9__13), .img_data_9__12 (
                        img_data_9__12), .img_data_9__11 (img_data_9__11), .img_data_9__10 (
                        img_data_9__10), .img_data_9__9 (img_data_9__9), .img_data_9__8 (
                        img_data_9__8), .img_data_9__7 (img_data_9__7), .img_data_9__6 (
                        img_data_9__6), .img_data_9__5 (img_data_9__5), .img_data_9__4 (
                        img_data_9__4), .img_data_9__3 (img_data_9__3), .img_data_9__2 (
                        img_data_9__2), .img_data_9__1 (img_data_9__1), .img_data_9__0 (
                        img_data_9__0), .img_data_10__15 (img_data_10__15), .img_data_10__14 (
                        img_data_10__14), .img_data_10__13 (img_data_10__13), .img_data_10__12 (
                        img_data_10__12), .img_data_10__11 (img_data_10__11), .img_data_10__10 (
                        img_data_10__10), .img_data_10__9 (img_data_10__9), .img_data_10__8 (
                        img_data_10__8), .img_data_10__7 (img_data_10__7), .img_data_10__6 (
                        img_data_10__6), .img_data_10__5 (img_data_10__5), .img_data_10__4 (
                        img_data_10__4), .img_data_10__3 (img_data_10__3), .img_data_10__2 (
                        img_data_10__2), .img_data_10__1 (img_data_10__1), .img_data_10__0 (
                        img_data_10__0), .img_data_11__15 (img_data_11__15), .img_data_11__14 (
                        img_data_11__14), .img_data_11__13 (img_data_11__13), .img_data_11__12 (
                        img_data_11__12), .img_data_11__11 (img_data_11__11), .img_data_11__10 (
                        img_data_11__10), .img_data_11__9 (img_data_11__9), .img_data_11__8 (
                        img_data_11__8), .img_data_11__7 (img_data_11__7), .img_data_11__6 (
                        img_data_11__6), .img_data_11__5 (img_data_11__5), .img_data_11__4 (
                        img_data_11__4), .img_data_11__3 (img_data_11__3), .img_data_11__2 (
                        img_data_11__2), .img_data_11__1 (img_data_11__1), .img_data_11__0 (
                        img_data_11__0), .img_data_12__15 (img_data_12__15), .img_data_12__14 (
                        img_data_12__14), .img_data_12__13 (img_data_12__13), .img_data_12__12 (
                        img_data_12__12), .img_data_12__11 (img_data_12__11), .img_data_12__10 (
                        img_data_12__10), .img_data_12__9 (img_data_12__9), .img_data_12__8 (
                        img_data_12__8), .img_data_12__7 (img_data_12__7), .img_data_12__6 (
                        img_data_12__6), .img_data_12__5 (img_data_12__5), .img_data_12__4 (
                        img_data_12__4), .img_data_12__3 (img_data_12__3), .img_data_12__2 (
                        img_data_12__2), .img_data_12__1 (img_data_12__1), .img_data_12__0 (
                        img_data_12__0), .img_data_13__15 (img_data_13__15), .img_data_13__14 (
                        img_data_13__14), .img_data_13__13 (img_data_13__13), .img_data_13__12 (
                        img_data_13__12), .img_data_13__11 (img_data_13__11), .img_data_13__10 (
                        img_data_13__10), .img_data_13__9 (img_data_13__9), .img_data_13__8 (
                        img_data_13__8), .img_data_13__7 (img_data_13__7), .img_data_13__6 (
                        img_data_13__6), .img_data_13__5 (img_data_13__5), .img_data_13__4 (
                        img_data_13__4), .img_data_13__3 (img_data_13__3), .img_data_13__2 (
                        img_data_13__2), .img_data_13__1 (img_data_13__1), .img_data_13__0 (
                        img_data_13__0), .img_data_14__15 (img_data_14__15), .img_data_14__14 (
                        img_data_14__14), .img_data_14__13 (img_data_14__13), .img_data_14__12 (
                        img_data_14__12), .img_data_14__11 (img_data_14__11), .img_data_14__10 (
                        img_data_14__10), .img_data_14__9 (img_data_14__9), .img_data_14__8 (
                        img_data_14__8), .img_data_14__7 (img_data_14__7), .img_data_14__6 (
                        img_data_14__6), .img_data_14__5 (img_data_14__5), .img_data_14__4 (
                        img_data_14__4), .img_data_14__3 (img_data_14__3), .img_data_14__2 (
                        img_data_14__2), .img_data_14__1 (img_data_14__1), .img_data_14__0 (
                        img_data_14__0), .img_data_15__15 (img_data_15__15), .img_data_15__14 (
                        img_data_15__14), .img_data_15__13 (img_data_15__13), .img_data_15__12 (
                        img_data_15__12), .img_data_15__11 (img_data_15__11), .img_data_15__10 (
                        img_data_15__10), .img_data_15__9 (img_data_15__9), .img_data_15__8 (
                        img_data_15__8), .img_data_15__7 (img_data_15__7), .img_data_15__6 (
                        img_data_15__6), .img_data_15__5 (img_data_15__5), .img_data_15__4 (
                        img_data_15__4), .img_data_15__3 (img_data_15__3), .img_data_15__2 (
                        img_data_15__2), .img_data_15__1 (img_data_15__1), .img_data_15__0 (
                        img_data_15__0), .img_data_16__15 (img_data_16__15), .img_data_16__14 (
                        img_data_16__14), .img_data_16__13 (img_data_16__13), .img_data_16__12 (
                        img_data_16__12), .img_data_16__11 (img_data_16__11), .img_data_16__10 (
                        img_data_16__10), .img_data_16__9 (img_data_16__9), .img_data_16__8 (
                        img_data_16__8), .img_data_16__7 (img_data_16__7), .img_data_16__6 (
                        img_data_16__6), .img_data_16__5 (img_data_16__5), .img_data_16__4 (
                        img_data_16__4), .img_data_16__3 (img_data_16__3), .img_data_16__2 (
                        img_data_16__2), .img_data_16__1 (img_data_16__1), .img_data_16__0 (
                        img_data_16__0), .img_data_17__15 (img_data_17__15), .img_data_17__14 (
                        img_data_17__14), .img_data_17__13 (img_data_17__13), .img_data_17__12 (
                        img_data_17__12), .img_data_17__11 (img_data_17__11), .img_data_17__10 (
                        img_data_17__10), .img_data_17__9 (img_data_17__9), .img_data_17__8 (
                        img_data_17__8), .img_data_17__7 (img_data_17__7), .img_data_17__6 (
                        img_data_17__6), .img_data_17__5 (img_data_17__5), .img_data_17__4 (
                        img_data_17__4), .img_data_17__3 (img_data_17__3), .img_data_17__2 (
                        img_data_17__2), .img_data_17__1 (img_data_17__1), .img_data_17__0 (
                        img_data_17__0), .img_data_18__15 (img_data_18__15), .img_data_18__14 (
                        img_data_18__14), .img_data_18__13 (img_data_18__13), .img_data_18__12 (
                        img_data_18__12), .img_data_18__11 (img_data_18__11), .img_data_18__10 (
                        img_data_18__10), .img_data_18__9 (img_data_18__9), .img_data_18__8 (
                        img_data_18__8), .img_data_18__7 (img_data_18__7), .img_data_18__6 (
                        img_data_18__6), .img_data_18__5 (img_data_18__5), .img_data_18__4 (
                        img_data_18__4), .img_data_18__3 (img_data_18__3), .img_data_18__2 (
                        img_data_18__2), .img_data_18__1 (img_data_18__1), .img_data_18__0 (
                        img_data_18__0), .img_data_19__15 (img_data_19__15), .img_data_19__14 (
                        img_data_19__14), .img_data_19__13 (img_data_19__13), .img_data_19__12 (
                        img_data_19__12), .img_data_19__11 (img_data_19__11), .img_data_19__10 (
                        img_data_19__10), .img_data_19__9 (img_data_19__9), .img_data_19__8 (
                        img_data_19__8), .img_data_19__7 (img_data_19__7), .img_data_19__6 (
                        img_data_19__6), .img_data_19__5 (img_data_19__5), .img_data_19__4 (
                        img_data_19__4), .img_data_19__3 (img_data_19__3), .img_data_19__2 (
                        img_data_19__2), .img_data_19__1 (img_data_19__1), .img_data_19__0 (
                        img_data_19__0), .img_data_20__15 (img_data_20__15), .img_data_20__14 (
                        img_data_20__14), .img_data_20__13 (img_data_20__13), .img_data_20__12 (
                        img_data_20__12), .img_data_20__11 (img_data_20__11), .img_data_20__10 (
                        img_data_20__10), .img_data_20__9 (img_data_20__9), .img_data_20__8 (
                        img_data_20__8), .img_data_20__7 (img_data_20__7), .img_data_20__6 (
                        img_data_20__6), .img_data_20__5 (img_data_20__5), .img_data_20__4 (
                        img_data_20__4), .img_data_20__3 (img_data_20__3), .img_data_20__2 (
                        img_data_20__2), .img_data_20__1 (img_data_20__1), .img_data_20__0 (
                        img_data_20__0), .img_data_21__15 (img_data_21__15), .img_data_21__14 (
                        img_data_21__14), .img_data_21__13 (img_data_21__13), .img_data_21__12 (
                        img_data_21__12), .img_data_21__11 (img_data_21__11), .img_data_21__10 (
                        img_data_21__10), .img_data_21__9 (img_data_21__9), .img_data_21__8 (
                        img_data_21__8), .img_data_21__7 (img_data_21__7), .img_data_21__6 (
                        img_data_21__6), .img_data_21__5 (img_data_21__5), .img_data_21__4 (
                        img_data_21__4), .img_data_21__3 (img_data_21__3), .img_data_21__2 (
                        img_data_21__2), .img_data_21__1 (img_data_21__1), .img_data_21__0 (
                        img_data_21__0), .img_data_22__15 (img_data_22__15), .img_data_22__14 (
                        img_data_22__14), .img_data_22__13 (img_data_22__13), .img_data_22__12 (
                        img_data_22__12), .img_data_22__11 (img_data_22__11), .img_data_22__10 (
                        img_data_22__10), .img_data_22__9 (img_data_22__9), .img_data_22__8 (
                        img_data_22__8), .img_data_22__7 (img_data_22__7), .img_data_22__6 (
                        img_data_22__6), .img_data_22__5 (img_data_22__5), .img_data_22__4 (
                        img_data_22__4), .img_data_22__3 (img_data_22__3), .img_data_22__2 (
                        img_data_22__2), .img_data_22__1 (img_data_22__1), .img_data_22__0 (
                        img_data_22__0), .img_data_23__15 (img_data_23__15), .img_data_23__14 (
                        img_data_23__14), .img_data_23__13 (img_data_23__13), .img_data_23__12 (
                        img_data_23__12), .img_data_23__11 (img_data_23__11), .img_data_23__10 (
                        img_data_23__10), .img_data_23__9 (img_data_23__9), .img_data_23__8 (
                        img_data_23__8), .img_data_23__7 (img_data_23__7), .img_data_23__6 (
                        img_data_23__6), .img_data_23__5 (img_data_23__5), .img_data_23__4 (
                        img_data_23__4), .img_data_23__3 (img_data_23__3), .img_data_23__2 (
                        img_data_23__2), .img_data_23__1 (img_data_23__1), .img_data_23__0 (
                        img_data_23__0), .img_data_24__15 (img_data_24__15), .img_data_24__14 (
                        img_data_24__14), .img_data_24__13 (img_data_24__13), .img_data_24__12 (
                        img_data_24__12), .img_data_24__11 (img_data_24__11), .img_data_24__10 (
                        img_data_24__10), .img_data_24__9 (img_data_24__9), .img_data_24__8 (
                        img_data_24__8), .img_data_24__7 (img_data_24__7), .img_data_24__6 (
                        img_data_24__6), .img_data_24__5 (img_data_24__5), .img_data_24__4 (
                        img_data_24__4), .img_data_24__3 (img_data_24__3), .img_data_24__2 (
                        img_data_24__2), .img_data_24__1 (img_data_24__1), .img_data_24__0 (
                        img_data_24__0), .filter_data_0__15 (filter_data_0__15)
                        , .filter_data_0__14 (filter_data_0__14), .filter_data_0__13 (
                        filter_data_0__13), .filter_data_0__12 (
                        filter_data_0__12), .filter_data_0__11 (
                        filter_data_0__11), .filter_data_0__10 (
                        filter_data_0__10), .filter_data_0__9 (filter_data_0__9)
                        , .filter_data_0__8 (filter_data_0__8), .filter_data_0__7 (
                        filter_data_0__7), .filter_data_0__6 (filter_data_0__6)
                        , .filter_data_0__5 (filter_data_0__5), .filter_data_0__4 (
                        filter_data_0__4), .filter_data_0__3 (filter_data_0__3)
                        , .filter_data_0__2 (filter_data_0__2), .filter_data_0__1 (
                        filter_data_0__1), .filter_data_0__0 (filter_data_0__0)
                        , .filter_data_1__15 (filter_data_1__15), .filter_data_1__14 (
                        filter_data_1__14), .filter_data_1__13 (
                        filter_data_1__13), .filter_data_1__12 (
                        filter_data_1__12), .filter_data_1__11 (
                        filter_data_1__11), .filter_data_1__10 (
                        filter_data_1__10), .filter_data_1__9 (filter_data_1__9)
                        , .filter_data_1__8 (filter_data_1__8), .filter_data_1__7 (
                        filter_data_1__7), .filter_data_1__6 (filter_data_1__6)
                        , .filter_data_1__5 (filter_data_1__5), .filter_data_1__4 (
                        filter_data_1__4), .filter_data_1__3 (filter_data_1__3)
                        , .filter_data_1__2 (filter_data_1__2), .filter_data_1__1 (
                        filter_data_1__1), .filter_data_1__0 (filter_data_1__0)
                        , .filter_data_2__15 (filter_data_2__15), .filter_data_2__14 (
                        filter_data_2__14), .filter_data_2__13 (
                        filter_data_2__13), .filter_data_2__12 (
                        filter_data_2__12), .filter_data_2__11 (
                        filter_data_2__11), .filter_data_2__10 (
                        filter_data_2__10), .filter_data_2__9 (filter_data_2__9)
                        , .filter_data_2__8 (filter_data_2__8), .filter_data_2__7 (
                        filter_data_2__7), .filter_data_2__6 (filter_data_2__6)
                        , .filter_data_2__5 (filter_data_2__5), .filter_data_2__4 (
                        filter_data_2__4), .filter_data_2__3 (filter_data_2__3)
                        , .filter_data_2__2 (filter_data_2__2), .filter_data_2__1 (
                        filter_data_2__1), .filter_data_2__0 (filter_data_2__0)
                        , .filter_data_3__15 (filter_data_3__15), .filter_data_3__14 (
                        filter_data_3__14), .filter_data_3__13 (
                        filter_data_3__13), .filter_data_3__12 (
                        filter_data_3__12), .filter_data_3__11 (
                        filter_data_3__11), .filter_data_3__10 (
                        filter_data_3__10), .filter_data_3__9 (filter_data_3__9)
                        , .filter_data_3__8 (filter_data_3__8), .filter_data_3__7 (
                        filter_data_3__7), .filter_data_3__6 (filter_data_3__6)
                        , .filter_data_3__5 (filter_data_3__5), .filter_data_3__4 (
                        filter_data_3__4), .filter_data_3__3 (filter_data_3__3)
                        , .filter_data_3__2 (filter_data_3__2), .filter_data_3__1 (
                        filter_data_3__1), .filter_data_3__0 (filter_data_3__0)
                        , .filter_data_4__15 (filter_data_4__15), .filter_data_4__14 (
                        filter_data_4__14), .filter_data_4__13 (
                        filter_data_4__13), .filter_data_4__12 (
                        filter_data_4__12), .filter_data_4__11 (
                        filter_data_4__11), .filter_data_4__10 (
                        filter_data_4__10), .filter_data_4__9 (filter_data_4__9)
                        , .filter_data_4__8 (filter_data_4__8), .filter_data_4__7 (
                        filter_data_4__7), .filter_data_4__6 (filter_data_4__6)
                        , .filter_data_4__5 (filter_data_4__5), .filter_data_4__4 (
                        filter_data_4__4), .filter_data_4__3 (filter_data_4__3)
                        , .filter_data_4__2 (filter_data_4__2), .filter_data_4__1 (
                        filter_data_4__1), .filter_data_4__0 (filter_data_4__0)
                        , .filter_data_5__15 (filter_data_5__15), .filter_data_5__14 (
                        filter_data_5__14), .filter_data_5__13 (
                        filter_data_5__13), .filter_data_5__12 (
                        filter_data_5__12), .filter_data_5__11 (
                        filter_data_5__11), .filter_data_5__10 (
                        filter_data_5__10), .filter_data_5__9 (filter_data_5__9)
                        , .filter_data_5__8 (filter_data_5__8), .filter_data_5__7 (
                        filter_data_5__7), .filter_data_5__6 (filter_data_5__6)
                        , .filter_data_5__5 (filter_data_5__5), .filter_data_5__4 (
                        filter_data_5__4), .filter_data_5__3 (filter_data_5__3)
                        , .filter_data_5__2 (filter_data_5__2), .filter_data_5__1 (
                        filter_data_5__1), .filter_data_5__0 (filter_data_5__0)
                        , .filter_data_6__15 (filter_data_6__15), .filter_data_6__14 (
                        filter_data_6__14), .filter_data_6__13 (
                        filter_data_6__13), .filter_data_6__12 (
                        filter_data_6__12), .filter_data_6__11 (
                        filter_data_6__11), .filter_data_6__10 (
                        filter_data_6__10), .filter_data_6__9 (filter_data_6__9)
                        , .filter_data_6__8 (filter_data_6__8), .filter_data_6__7 (
                        filter_data_6__7), .filter_data_6__6 (filter_data_6__6)
                        , .filter_data_6__5 (filter_data_6__5), .filter_data_6__4 (
                        filter_data_6__4), .filter_data_6__3 (filter_data_6__3)
                        , .filter_data_6__2 (filter_data_6__2), .filter_data_6__1 (
                        filter_data_6__1), .filter_data_6__0 (filter_data_6__0)
                        , .filter_data_7__15 (filter_data_7__15), .filter_data_7__14 (
                        filter_data_7__14), .filter_data_7__13 (
                        filter_data_7__13), .filter_data_7__12 (
                        filter_data_7__12), .filter_data_7__11 (
                        filter_data_7__11), .filter_data_7__10 (
                        filter_data_7__10), .filter_data_7__9 (filter_data_7__9)
                        , .filter_data_7__8 (filter_data_7__8), .filter_data_7__7 (
                        filter_data_7__7), .filter_data_7__6 (filter_data_7__6)
                        , .filter_data_7__5 (filter_data_7__5), .filter_data_7__4 (
                        filter_data_7__4), .filter_data_7__3 (filter_data_7__3)
                        , .filter_data_7__2 (filter_data_7__2), .filter_data_7__1 (
                        filter_data_7__1), .filter_data_7__0 (filter_data_7__0)
                        , .filter_data_8__15 (filter_data_8__15), .filter_data_8__14 (
                        filter_data_8__14), .filter_data_8__13 (
                        filter_data_8__13), .filter_data_8__12 (
                        filter_data_8__12), .filter_data_8__11 (
                        filter_data_8__11), .filter_data_8__10 (
                        filter_data_8__10), .filter_data_8__9 (filter_data_8__9)
                        , .filter_data_8__8 (filter_data_8__8), .filter_data_8__7 (
                        filter_data_8__7), .filter_data_8__6 (filter_data_8__6)
                        , .filter_data_8__5 (filter_data_8__5), .filter_data_8__4 (
                        filter_data_8__4), .filter_data_8__3 (filter_data_8__3)
                        , .filter_data_8__2 (filter_data_8__2), .filter_data_8__1 (
                        filter_data_8__1), .filter_data_8__0 (filter_data_8__0)
                        , .filter_data_9__15 (filter_data_9__15), .filter_data_9__14 (
                        filter_data_9__14), .filter_data_9__13 (
                        filter_data_9__13), .filter_data_9__12 (
                        filter_data_9__12), .filter_data_9__11 (
                        filter_data_9__11), .filter_data_9__10 (
                        filter_data_9__10), .filter_data_9__9 (filter_data_9__9)
                        , .filter_data_9__8 (filter_data_9__8), .filter_data_9__7 (
                        filter_data_9__7), .filter_data_9__6 (filter_data_9__6)
                        , .filter_data_9__5 (filter_data_9__5), .filter_data_9__4 (
                        filter_data_9__4), .filter_data_9__3 (filter_data_9__3)
                        , .filter_data_9__2 (filter_data_9__2), .filter_data_9__1 (
                        filter_data_9__1), .filter_data_9__0 (filter_data_9__0)
                        , .filter_data_10__15 (filter_data_10__15), .filter_data_10__14 (
                        filter_data_10__14), .filter_data_10__13 (
                        filter_data_10__13), .filter_data_10__12 (
                        filter_data_10__12), .filter_data_10__11 (
                        filter_data_10__11), .filter_data_10__10 (
                        filter_data_10__10), .filter_data_10__9 (
                        filter_data_10__9), .filter_data_10__8 (
                        filter_data_10__8), .filter_data_10__7 (
                        filter_data_10__7), .filter_data_10__6 (
                        filter_data_10__6), .filter_data_10__5 (
                        filter_data_10__5), .filter_data_10__4 (
                        filter_data_10__4), .filter_data_10__3 (
                        filter_data_10__3), .filter_data_10__2 (
                        filter_data_10__2), .filter_data_10__1 (
                        filter_data_10__1), .filter_data_10__0 (
                        filter_data_10__0), .filter_data_11__15 (
                        filter_data_11__15), .filter_data_11__14 (
                        filter_data_11__14), .filter_data_11__13 (
                        filter_data_11__13), .filter_data_11__12 (
                        filter_data_11__12), .filter_data_11__11 (
                        filter_data_11__11), .filter_data_11__10 (
                        filter_data_11__10), .filter_data_11__9 (
                        filter_data_11__9), .filter_data_11__8 (
                        filter_data_11__8), .filter_data_11__7 (
                        filter_data_11__7), .filter_data_11__6 (
                        filter_data_11__6), .filter_data_11__5 (
                        filter_data_11__5), .filter_data_11__4 (
                        filter_data_11__4), .filter_data_11__3 (
                        filter_data_11__3), .filter_data_11__2 (
                        filter_data_11__2), .filter_data_11__1 (
                        filter_data_11__1), .filter_data_11__0 (
                        filter_data_11__0), .filter_data_12__15 (
                        filter_data_12__15), .filter_data_12__14 (
                        filter_data_12__14), .filter_data_12__13 (
                        filter_data_12__13), .filter_data_12__12 (
                        filter_data_12__12), .filter_data_12__11 (
                        filter_data_12__11), .filter_data_12__10 (
                        filter_data_12__10), .filter_data_12__9 (
                        filter_data_12__9), .filter_data_12__8 (
                        filter_data_12__8), .filter_data_12__7 (
                        filter_data_12__7), .filter_data_12__6 (
                        filter_data_12__6), .filter_data_12__5 (
                        filter_data_12__5), .filter_data_12__4 (
                        filter_data_12__4), .filter_data_12__3 (
                        filter_data_12__3), .filter_data_12__2 (
                        filter_data_12__2), .filter_data_12__1 (
                        filter_data_12__1), .filter_data_12__0 (
                        filter_data_12__0), .filter_data_13__15 (
                        filter_data_13__15), .filter_data_13__14 (
                        filter_data_13__14), .filter_data_13__13 (
                        filter_data_13__13), .filter_data_13__12 (
                        filter_data_13__12), .filter_data_13__11 (
                        filter_data_13__11), .filter_data_13__10 (
                        filter_data_13__10), .filter_data_13__9 (
                        filter_data_13__9), .filter_data_13__8 (
                        filter_data_13__8), .filter_data_13__7 (
                        filter_data_13__7), .filter_data_13__6 (
                        filter_data_13__6), .filter_data_13__5 (
                        filter_data_13__5), .filter_data_13__4 (
                        filter_data_13__4), .filter_data_13__3 (
                        filter_data_13__3), .filter_data_13__2 (
                        filter_data_13__2), .filter_data_13__1 (
                        filter_data_13__1), .filter_data_13__0 (
                        filter_data_13__0), .filter_data_14__15 (
                        filter_data_14__15), .filter_data_14__14 (
                        filter_data_14__14), .filter_data_14__13 (
                        filter_data_14__13), .filter_data_14__12 (
                        filter_data_14__12), .filter_data_14__11 (
                        filter_data_14__11), .filter_data_14__10 (
                        filter_data_14__10), .filter_data_14__9 (
                        filter_data_14__9), .filter_data_14__8 (
                        filter_data_14__8), .filter_data_14__7 (
                        filter_data_14__7), .filter_data_14__6 (
                        filter_data_14__6), .filter_data_14__5 (
                        filter_data_14__5), .filter_data_14__4 (
                        filter_data_14__4), .filter_data_14__3 (
                        filter_data_14__3), .filter_data_14__2 (
                        filter_data_14__2), .filter_data_14__1 (
                        filter_data_14__1), .filter_data_14__0 (
                        filter_data_14__0), .filter_data_15__15 (
                        filter_data_15__15), .filter_data_15__14 (
                        filter_data_15__14), .filter_data_15__13 (
                        filter_data_15__13), .filter_data_15__12 (
                        filter_data_15__12), .filter_data_15__11 (
                        filter_data_15__11), .filter_data_15__10 (
                        filter_data_15__10), .filter_data_15__9 (
                        filter_data_15__9), .filter_data_15__8 (
                        filter_data_15__8), .filter_data_15__7 (
                        filter_data_15__7), .filter_data_15__6 (
                        filter_data_15__6), .filter_data_15__5 (
                        filter_data_15__5), .filter_data_15__4 (
                        filter_data_15__4), .filter_data_15__3 (
                        filter_data_15__3), .filter_data_15__2 (
                        filter_data_15__2), .filter_data_15__1 (
                        filter_data_15__1), .filter_data_15__0 (
                        filter_data_15__0), .filter_data_16__15 (
                        filter_data_16__15), .filter_data_16__14 (
                        filter_data_16__14), .filter_data_16__13 (
                        filter_data_16__13), .filter_data_16__12 (
                        filter_data_16__12), .filter_data_16__11 (
                        filter_data_16__11), .filter_data_16__10 (
                        filter_data_16__10), .filter_data_16__9 (
                        filter_data_16__9), .filter_data_16__8 (
                        filter_data_16__8), .filter_data_16__7 (
                        filter_data_16__7), .filter_data_16__6 (
                        filter_data_16__6), .filter_data_16__5 (
                        filter_data_16__5), .filter_data_16__4 (
                        filter_data_16__4), .filter_data_16__3 (
                        filter_data_16__3), .filter_data_16__2 (
                        filter_data_16__2), .filter_data_16__1 (
                        filter_data_16__1), .filter_data_16__0 (
                        filter_data_16__0), .filter_data_17__15 (
                        filter_data_17__15), .filter_data_17__14 (
                        filter_data_17__14), .filter_data_17__13 (
                        filter_data_17__13), .filter_data_17__12 (
                        filter_data_17__12), .filter_data_17__11 (
                        filter_data_17__11), .filter_data_17__10 (
                        filter_data_17__10), .filter_data_17__9 (
                        filter_data_17__9), .filter_data_17__8 (
                        filter_data_17__8), .filter_data_17__7 (
                        filter_data_17__7), .filter_data_17__6 (
                        filter_data_17__6), .filter_data_17__5 (
                        filter_data_17__5), .filter_data_17__4 (
                        filter_data_17__4), .filter_data_17__3 (
                        filter_data_17__3), .filter_data_17__2 (
                        filter_data_17__2), .filter_data_17__1 (
                        filter_data_17__1), .filter_data_17__0 (
                        filter_data_17__0), .filter_data_18__15 (
                        filter_data_18__15), .filter_data_18__14 (
                        filter_data_18__14), .filter_data_18__13 (
                        filter_data_18__13), .filter_data_18__12 (
                        filter_data_18__12), .filter_data_18__11 (
                        filter_data_18__11), .filter_data_18__10 (
                        filter_data_18__10), .filter_data_18__9 (
                        filter_data_18__9), .filter_data_18__8 (
                        filter_data_18__8), .filter_data_18__7 (
                        filter_data_18__7), .filter_data_18__6 (
                        filter_data_18__6), .filter_data_18__5 (
                        filter_data_18__5), .filter_data_18__4 (
                        filter_data_18__4), .filter_data_18__3 (
                        filter_data_18__3), .filter_data_18__2 (
                        filter_data_18__2), .filter_data_18__1 (
                        filter_data_18__1), .filter_data_18__0 (
                        filter_data_18__0), .filter_data_19__15 (
                        filter_data_19__15), .filter_data_19__14 (
                        filter_data_19__14), .filter_data_19__13 (
                        filter_data_19__13), .filter_data_19__12 (
                        filter_data_19__12), .filter_data_19__11 (
                        filter_data_19__11), .filter_data_19__10 (
                        filter_data_19__10), .filter_data_19__9 (
                        filter_data_19__9), .filter_data_19__8 (
                        filter_data_19__8), .filter_data_19__7 (
                        filter_data_19__7), .filter_data_19__6 (
                        filter_data_19__6), .filter_data_19__5 (
                        filter_data_19__5), .filter_data_19__4 (
                        filter_data_19__4), .filter_data_19__3 (
                        filter_data_19__3), .filter_data_19__2 (
                        filter_data_19__2), .filter_data_19__1 (
                        filter_data_19__1), .filter_data_19__0 (
                        filter_data_19__0), .filter_data_20__15 (
                        filter_data_20__15), .filter_data_20__14 (
                        filter_data_20__14), .filter_data_20__13 (
                        filter_data_20__13), .filter_data_20__12 (
                        filter_data_20__12), .filter_data_20__11 (
                        filter_data_20__11), .filter_data_20__10 (
                        filter_data_20__10), .filter_data_20__9 (
                        filter_data_20__9), .filter_data_20__8 (
                        filter_data_20__8), .filter_data_20__7 (
                        filter_data_20__7), .filter_data_20__6 (
                        filter_data_20__6), .filter_data_20__5 (
                        filter_data_20__5), .filter_data_20__4 (
                        filter_data_20__4), .filter_data_20__3 (
                        filter_data_20__3), .filter_data_20__2 (
                        filter_data_20__2), .filter_data_20__1 (
                        filter_data_20__1), .filter_data_20__0 (
                        filter_data_20__0), .filter_data_21__15 (
                        filter_data_21__15), .filter_data_21__14 (
                        filter_data_21__14), .filter_data_21__13 (
                        filter_data_21__13), .filter_data_21__12 (
                        filter_data_21__12), .filter_data_21__11 (
                        filter_data_21__11), .filter_data_21__10 (
                        filter_data_21__10), .filter_data_21__9 (
                        filter_data_21__9), .filter_data_21__8 (
                        filter_data_21__8), .filter_data_21__7 (
                        filter_data_21__7), .filter_data_21__6 (
                        filter_data_21__6), .filter_data_21__5 (
                        filter_data_21__5), .filter_data_21__4 (
                        filter_data_21__4), .filter_data_21__3 (
                        filter_data_21__3), .filter_data_21__2 (
                        filter_data_21__2), .filter_data_21__1 (
                        filter_data_21__1), .filter_data_21__0 (
                        filter_data_21__0), .filter_data_22__15 (
                        filter_data_22__15), .filter_data_22__14 (
                        filter_data_22__14), .filter_data_22__13 (
                        filter_data_22__13), .filter_data_22__12 (
                        filter_data_22__12), .filter_data_22__11 (
                        filter_data_22__11), .filter_data_22__10 (
                        filter_data_22__10), .filter_data_22__9 (
                        filter_data_22__9), .filter_data_22__8 (
                        filter_data_22__8), .filter_data_22__7 (
                        filter_data_22__7), .filter_data_22__6 (
                        filter_data_22__6), .filter_data_22__5 (
                        filter_data_22__5), .filter_data_22__4 (
                        filter_data_22__4), .filter_data_22__3 (
                        filter_data_22__3), .filter_data_22__2 (
                        filter_data_22__2), .filter_data_22__1 (
                        filter_data_22__1), .filter_data_22__0 (
                        filter_data_22__0), .filter_data_23__15 (
                        filter_data_23__15), .filter_data_23__14 (
                        filter_data_23__14), .filter_data_23__13 (
                        filter_data_23__13), .filter_data_23__12 (
                        filter_data_23__12), .filter_data_23__11 (
                        filter_data_23__11), .filter_data_23__10 (
                        filter_data_23__10), .filter_data_23__9 (
                        filter_data_23__9), .filter_data_23__8 (
                        filter_data_23__8), .filter_data_23__7 (
                        filter_data_23__7), .filter_data_23__6 (
                        filter_data_23__6), .filter_data_23__5 (
                        filter_data_23__5), .filter_data_23__4 (
                        filter_data_23__4), .filter_data_23__3 (
                        filter_data_23__3), .filter_data_23__2 (
                        filter_data_23__2), .filter_data_23__1 (
                        filter_data_23__1), .filter_data_23__0 (
                        filter_data_23__0), .filter_data_24__15 (
                        filter_data_24__15), .filter_data_24__14 (
                        filter_data_24__14), .filter_data_24__13 (
                        filter_data_24__13), .filter_data_24__12 (
                        filter_data_24__12), .filter_data_24__11 (
                        filter_data_24__11), .filter_data_24__10 (
                        filter_data_24__10), .filter_data_24__9 (
                        filter_data_24__9), .filter_data_24__8 (
                        filter_data_24__8), .filter_data_24__7 (
                        filter_data_24__7), .filter_data_24__6 (
                        filter_data_24__6), .filter_data_24__5 (
                        filter_data_24__5), .filter_data_24__4 (
                        filter_data_24__4), .filter_data_24__3 (
                        filter_data_24__3), .filter_data_24__2 (
                        filter_data_24__2), .filter_data_24__1 (
                        filter_data_24__1), .filter_data_24__0 (
                        filter_data_24__0), .d_arr_0__31 (d_cache_arr_0__31), .d_arr_0__30 (
                        d_cache_arr_0__30), .d_arr_0__29 (d_cache_arr_0__29), .d_arr_0__28 (
                        d_cache_arr_0__28), .d_arr_0__27 (d_cache_arr_0__27), .d_arr_0__26 (
                        d_cache_arr_0__26), .d_arr_0__25 (d_cache_arr_0__25), .d_arr_0__24 (
                        d_cache_arr_0__24), .d_arr_0__23 (d_cache_arr_0__23), .d_arr_0__22 (
                        d_cache_arr_0__22), .d_arr_0__21 (d_cache_arr_0__21), .d_arr_0__20 (
                        d_cache_arr_0__20), .d_arr_0__19 (d_cache_arr_0__19), .d_arr_0__18 (
                        d_cache_arr_0__18), .d_arr_0__17 (d_cache_arr_0__17), .d_arr_0__16 (
                        d_cache_arr_0__16), .d_arr_0__15 (d_cache_arr_0__15), .d_arr_0__14 (
                        d_cache_arr_0__14), .d_arr_0__13 (d_cache_arr_0__13), .d_arr_0__12 (
                        d_cache_arr_0__12), .d_arr_0__11 (d_cache_arr_0__11), .d_arr_0__10 (
                        d_cache_arr_0__10), .d_arr_0__9 (d_cache_arr_0__9), .d_arr_0__8 (
                        d_cache_arr_0__8), .d_arr_0__7 (d_cache_arr_0__7), .d_arr_0__6 (
                        d_cache_arr_0__6), .d_arr_0__5 (d_cache_arr_0__5), .d_arr_0__4 (
                        d_cache_arr_0__4), .d_arr_0__3 (d_cache_arr_0__3), .d_arr_0__2 (
                        d_cache_arr_0__2), .d_arr_0__1 (d_cache_arr_0__1), .d_arr_0__0 (
                        d_cache_arr_0__0), .d_arr_1__31 (d_cache_arr_1__31), .d_arr_1__30 (
                        d_cache_arr_1__30), .d_arr_1__29 (d_cache_arr_1__29), .d_arr_1__28 (
                        d_cache_arr_1__28), .d_arr_1__27 (d_cache_arr_1__27), .d_arr_1__26 (
                        d_cache_arr_1__26), .d_arr_1__25 (d_cache_arr_1__25), .d_arr_1__24 (
                        d_cache_arr_1__24), .d_arr_1__23 (d_cache_arr_1__23), .d_arr_1__22 (
                        d_cache_arr_1__22), .d_arr_1__21 (d_cache_arr_1__21), .d_arr_1__20 (
                        d_cache_arr_1__20), .d_arr_1__19 (d_cache_arr_1__19), .d_arr_1__18 (
                        d_cache_arr_1__18), .d_arr_1__17 (d_cache_arr_1__17), .d_arr_1__16 (
                        d_cache_arr_1__16), .d_arr_1__15 (d_cache_arr_1__15), .d_arr_1__14 (
                        d_cache_arr_1__14), .d_arr_1__13 (d_cache_arr_1__13), .d_arr_1__12 (
                        d_cache_arr_1__12), .d_arr_1__11 (d_cache_arr_1__11), .d_arr_1__10 (
                        d_cache_arr_1__10), .d_arr_1__9 (d_cache_arr_1__9), .d_arr_1__8 (
                        d_cache_arr_1__8), .d_arr_1__7 (d_cache_arr_1__7), .d_arr_1__6 (
                        d_cache_arr_1__6), .d_arr_1__5 (d_cache_arr_1__5), .d_arr_1__4 (
                        d_cache_arr_1__4), .d_arr_1__3 (d_cache_arr_1__3), .d_arr_1__2 (
                        d_cache_arr_1__2), .d_arr_1__1 (d_cache_arr_1__1), .d_arr_1__0 (
                        d_cache_arr_1__0), .d_arr_2__31 (d_cache_arr_2__31), .d_arr_2__30 (
                        d_cache_arr_2__30), .d_arr_2__29 (d_cache_arr_2__29), .d_arr_2__28 (
                        d_cache_arr_2__28), .d_arr_2__27 (d_cache_arr_2__27), .d_arr_2__26 (
                        d_cache_arr_2__26), .d_arr_2__25 (d_cache_arr_2__25), .d_arr_2__24 (
                        d_cache_arr_2__24), .d_arr_2__23 (d_cache_arr_2__23), .d_arr_2__22 (
                        d_cache_arr_2__22), .d_arr_2__21 (d_cache_arr_2__21), .d_arr_2__20 (
                        d_cache_arr_2__20), .d_arr_2__19 (d_cache_arr_2__19), .d_arr_2__18 (
                        d_cache_arr_2__18), .d_arr_2__17 (d_cache_arr_2__17), .d_arr_2__16 (
                        d_cache_arr_2__16), .d_arr_2__15 (d_cache_arr_2__15), .d_arr_2__14 (
                        d_cache_arr_2__14), .d_arr_2__13 (d_cache_arr_2__13), .d_arr_2__12 (
                        d_cache_arr_2__12), .d_arr_2__11 (d_cache_arr_2__11), .d_arr_2__10 (
                        d_cache_arr_2__10), .d_arr_2__9 (d_cache_arr_2__9), .d_arr_2__8 (
                        d_cache_arr_2__8), .d_arr_2__7 (d_cache_arr_2__7), .d_arr_2__6 (
                        d_cache_arr_2__6), .d_arr_2__5 (d_cache_arr_2__5), .d_arr_2__4 (
                        d_cache_arr_2__4), .d_arr_2__3 (d_cache_arr_2__3), .d_arr_2__2 (
                        d_cache_arr_2__2), .d_arr_2__1 (d_cache_arr_2__1), .d_arr_2__0 (
                        d_cache_arr_2__0), .d_arr_3__31 (d_cache_arr_3__31), .d_arr_3__30 (
                        d_cache_arr_3__30), .d_arr_3__29 (d_cache_arr_3__29), .d_arr_3__28 (
                        d_cache_arr_3__28), .d_arr_3__27 (d_cache_arr_3__27), .d_arr_3__26 (
                        d_cache_arr_3__26), .d_arr_3__25 (d_cache_arr_3__25), .d_arr_3__24 (
                        d_cache_arr_3__24), .d_arr_3__23 (d_cache_arr_3__23), .d_arr_3__22 (
                        d_cache_arr_3__22), .d_arr_3__21 (d_cache_arr_3__21), .d_arr_3__20 (
                        d_cache_arr_3__20), .d_arr_3__19 (d_cache_arr_3__19), .d_arr_3__18 (
                        d_cache_arr_3__18), .d_arr_3__17 (d_cache_arr_3__17), .d_arr_3__16 (
                        d_cache_arr_3__16), .d_arr_3__15 (d_cache_arr_3__15), .d_arr_3__14 (
                        d_cache_arr_3__14), .d_arr_3__13 (d_cache_arr_3__13), .d_arr_3__12 (
                        d_cache_arr_3__12), .d_arr_3__11 (d_cache_arr_3__11), .d_arr_3__10 (
                        d_cache_arr_3__10), .d_arr_3__9 (d_cache_arr_3__9), .d_arr_3__8 (
                        d_cache_arr_3__8), .d_arr_3__7 (d_cache_arr_3__7), .d_arr_3__6 (
                        d_cache_arr_3__6), .d_arr_3__5 (d_cache_arr_3__5), .d_arr_3__4 (
                        d_cache_arr_3__4), .d_arr_3__3 (d_cache_arr_3__3), .d_arr_3__2 (
                        d_cache_arr_3__2), .d_arr_3__1 (d_cache_arr_3__1), .d_arr_3__0 (
                        d_cache_arr_3__0), .d_arr_4__31 (d_cache_arr_4__31), .d_arr_4__30 (
                        d_cache_arr_4__30), .d_arr_4__29 (d_cache_arr_4__29), .d_arr_4__28 (
                        d_cache_arr_4__28), .d_arr_4__27 (d_cache_arr_4__27), .d_arr_4__26 (
                        d_cache_arr_4__26), .d_arr_4__25 (d_cache_arr_4__25), .d_arr_4__24 (
                        d_cache_arr_4__24), .d_arr_4__23 (d_cache_arr_4__23), .d_arr_4__22 (
                        d_cache_arr_4__22), .d_arr_4__21 (d_cache_arr_4__21), .d_arr_4__20 (
                        d_cache_arr_4__20), .d_arr_4__19 (d_cache_arr_4__19), .d_arr_4__18 (
                        d_cache_arr_4__18), .d_arr_4__17 (d_cache_arr_4__17), .d_arr_4__16 (
                        d_cache_arr_4__16), .d_arr_4__15 (d_cache_arr_4__15), .d_arr_4__14 (
                        d_cache_arr_4__14), .d_arr_4__13 (d_cache_arr_4__13), .d_arr_4__12 (
                        d_cache_arr_4__12), .d_arr_4__11 (d_cache_arr_4__11), .d_arr_4__10 (
                        d_cache_arr_4__10), .d_arr_4__9 (d_cache_arr_4__9), .d_arr_4__8 (
                        d_cache_arr_4__8), .d_arr_4__7 (d_cache_arr_4__7), .d_arr_4__6 (
                        d_cache_arr_4__6), .d_arr_4__5 (d_cache_arr_4__5), .d_arr_4__4 (
                        d_cache_arr_4__4), .d_arr_4__3 (d_cache_arr_4__3), .d_arr_4__2 (
                        d_cache_arr_4__2), .d_arr_4__1 (d_cache_arr_4__1), .d_arr_4__0 (
                        d_cache_arr_4__0), .d_arr_5__31 (d_cache_arr_5__31), .d_arr_5__30 (
                        d_cache_arr_5__30), .d_arr_5__29 (d_cache_arr_5__29), .d_arr_5__28 (
                        d_cache_arr_5__28), .d_arr_5__27 (d_cache_arr_5__27), .d_arr_5__26 (
                        d_cache_arr_5__26), .d_arr_5__25 (d_cache_arr_5__25), .d_arr_5__24 (
                        d_cache_arr_5__24), .d_arr_5__23 (d_cache_arr_5__23), .d_arr_5__22 (
                        d_cache_arr_5__22), .d_arr_5__21 (d_cache_arr_5__21), .d_arr_5__20 (
                        d_cache_arr_5__20), .d_arr_5__19 (d_cache_arr_5__19), .d_arr_5__18 (
                        d_cache_arr_5__18), .d_arr_5__17 (d_cache_arr_5__17), .d_arr_5__16 (
                        d_cache_arr_5__16), .d_arr_5__15 (d_cache_arr_5__15), .d_arr_5__14 (
                        d_cache_arr_5__14), .d_arr_5__13 (d_cache_arr_5__13), .d_arr_5__12 (
                        d_cache_arr_5__12), .d_arr_5__11 (d_cache_arr_5__11), .d_arr_5__10 (
                        d_cache_arr_5__10), .d_arr_5__9 (d_cache_arr_5__9), .d_arr_5__8 (
                        d_cache_arr_5__8), .d_arr_5__7 (d_cache_arr_5__7), .d_arr_5__6 (
                        d_cache_arr_5__6), .d_arr_5__5 (d_cache_arr_5__5), .d_arr_5__4 (
                        d_cache_arr_5__4), .d_arr_5__3 (d_cache_arr_5__3), .d_arr_5__2 (
                        d_cache_arr_5__2), .d_arr_5__1 (d_cache_arr_5__1), .d_arr_5__0 (
                        d_cache_arr_5__0), .d_arr_6__31 (d_cache_arr_6__31), .d_arr_6__30 (
                        d_cache_arr_6__30), .d_arr_6__29 (d_cache_arr_6__29), .d_arr_6__28 (
                        d_cache_arr_6__28), .d_arr_6__27 (d_cache_arr_6__27), .d_arr_6__26 (
                        d_cache_arr_6__26), .d_arr_6__25 (d_cache_arr_6__25), .d_arr_6__24 (
                        d_cache_arr_6__24), .d_arr_6__23 (d_cache_arr_6__23), .d_arr_6__22 (
                        d_cache_arr_6__22), .d_arr_6__21 (d_cache_arr_6__21), .d_arr_6__20 (
                        d_cache_arr_6__20), .d_arr_6__19 (d_cache_arr_6__19), .d_arr_6__18 (
                        d_cache_arr_6__18), .d_arr_6__17 (d_cache_arr_6__17), .d_arr_6__16 (
                        d_cache_arr_6__16), .d_arr_6__15 (d_cache_arr_6__15), .d_arr_6__14 (
                        d_cache_arr_6__14), .d_arr_6__13 (d_cache_arr_6__13), .d_arr_6__12 (
                        d_cache_arr_6__12), .d_arr_6__11 (d_cache_arr_6__11), .d_arr_6__10 (
                        d_cache_arr_6__10), .d_arr_6__9 (d_cache_arr_6__9), .d_arr_6__8 (
                        d_cache_arr_6__8), .d_arr_6__7 (d_cache_arr_6__7), .d_arr_6__6 (
                        d_cache_arr_6__6), .d_arr_6__5 (d_cache_arr_6__5), .d_arr_6__4 (
                        d_cache_arr_6__4), .d_arr_6__3 (d_cache_arr_6__3), .d_arr_6__2 (
                        d_cache_arr_6__2), .d_arr_6__1 (d_cache_arr_6__1), .d_arr_6__0 (
                        d_cache_arr_6__0), .d_arr_7__31 (d_cache_arr_7__31), .d_arr_7__30 (
                        d_cache_arr_7__30), .d_arr_7__29 (d_cache_arr_7__29), .d_arr_7__28 (
                        d_cache_arr_7__28), .d_arr_7__27 (d_cache_arr_7__27), .d_arr_7__26 (
                        d_cache_arr_7__26), .d_arr_7__25 (d_cache_arr_7__25), .d_arr_7__24 (
                        d_cache_arr_7__24), .d_arr_7__23 (d_cache_arr_7__23), .d_arr_7__22 (
                        d_cache_arr_7__22), .d_arr_7__21 (d_cache_arr_7__21), .d_arr_7__20 (
                        d_cache_arr_7__20), .d_arr_7__19 (d_cache_arr_7__19), .d_arr_7__18 (
                        d_cache_arr_7__18), .d_arr_7__17 (d_cache_arr_7__17), .d_arr_7__16 (
                        d_cache_arr_7__16), .d_arr_7__15 (d_cache_arr_7__15), .d_arr_7__14 (
                        d_cache_arr_7__14), .d_arr_7__13 (d_cache_arr_7__13), .d_arr_7__12 (
                        d_cache_arr_7__12), .d_arr_7__11 (d_cache_arr_7__11), .d_arr_7__10 (
                        d_cache_arr_7__10), .d_arr_7__9 (d_cache_arr_7__9), .d_arr_7__8 (
                        d_cache_arr_7__8), .d_arr_7__7 (d_cache_arr_7__7), .d_arr_7__6 (
                        d_cache_arr_7__6), .d_arr_7__5 (d_cache_arr_7__5), .d_arr_7__4 (
                        d_cache_arr_7__4), .d_arr_7__3 (d_cache_arr_7__3), .d_arr_7__2 (
                        d_cache_arr_7__2), .d_arr_7__1 (d_cache_arr_7__1), .d_arr_7__0 (
                        d_cache_arr_7__0), .d_arr_8__31 (d_cache_arr_8__31), .d_arr_8__30 (
                        d_cache_arr_8__30), .d_arr_8__29 (d_cache_arr_8__29), .d_arr_8__28 (
                        d_cache_arr_8__28), .d_arr_8__27 (d_cache_arr_8__27), .d_arr_8__26 (
                        d_cache_arr_8__26), .d_arr_8__25 (d_cache_arr_8__25), .d_arr_8__24 (
                        d_cache_arr_8__24), .d_arr_8__23 (d_cache_arr_8__23), .d_arr_8__22 (
                        d_cache_arr_8__22), .d_arr_8__21 (d_cache_arr_8__21), .d_arr_8__20 (
                        d_cache_arr_8__20), .d_arr_8__19 (d_cache_arr_8__19), .d_arr_8__18 (
                        d_cache_arr_8__18), .d_arr_8__17 (d_cache_arr_8__17), .d_arr_8__16 (
                        d_cache_arr_8__16), .d_arr_8__15 (d_cache_arr_8__15), .d_arr_8__14 (
                        d_cache_arr_8__14), .d_arr_8__13 (d_cache_arr_8__13), .d_arr_8__12 (
                        d_cache_arr_8__12), .d_arr_8__11 (d_cache_arr_8__11), .d_arr_8__10 (
                        d_cache_arr_8__10), .d_arr_8__9 (d_cache_arr_8__9), .d_arr_8__8 (
                        d_cache_arr_8__8), .d_arr_8__7 (d_cache_arr_8__7), .d_arr_8__6 (
                        d_cache_arr_8__6), .d_arr_8__5 (d_cache_arr_8__5), .d_arr_8__4 (
                        d_cache_arr_8__4), .d_arr_8__3 (d_cache_arr_8__3), .d_arr_8__2 (
                        d_cache_arr_8__2), .d_arr_8__1 (d_cache_arr_8__1), .d_arr_8__0 (
                        d_cache_arr_8__0), .d_arr_9__31 (d_cache_arr_9__31), .d_arr_9__30 (
                        d_cache_arr_9__30), .d_arr_9__29 (d_cache_arr_9__29), .d_arr_9__28 (
                        d_cache_arr_9__28), .d_arr_9__27 (d_cache_arr_9__27), .d_arr_9__26 (
                        d_cache_arr_9__26), .d_arr_9__25 (d_cache_arr_9__25), .d_arr_9__24 (
                        d_cache_arr_9__24), .d_arr_9__23 (d_cache_arr_9__23), .d_arr_9__22 (
                        d_cache_arr_9__22), .d_arr_9__21 (d_cache_arr_9__21), .d_arr_9__20 (
                        d_cache_arr_9__20), .d_arr_9__19 (d_cache_arr_9__19), .d_arr_9__18 (
                        d_cache_arr_9__18), .d_arr_9__17 (d_cache_arr_9__17), .d_arr_9__16 (
                        d_cache_arr_9__16), .d_arr_9__15 (d_cache_arr_9__15), .d_arr_9__14 (
                        d_cache_arr_9__14), .d_arr_9__13 (d_cache_arr_9__13), .d_arr_9__12 (
                        d_cache_arr_9__12), .d_arr_9__11 (d_cache_arr_9__11), .d_arr_9__10 (
                        d_cache_arr_9__10), .d_arr_9__9 (d_cache_arr_9__9), .d_arr_9__8 (
                        d_cache_arr_9__8), .d_arr_9__7 (d_cache_arr_9__7), .d_arr_9__6 (
                        d_cache_arr_9__6), .d_arr_9__5 (d_cache_arr_9__5), .d_arr_9__4 (
                        d_cache_arr_9__4), .d_arr_9__3 (d_cache_arr_9__3), .d_arr_9__2 (
                        d_cache_arr_9__2), .d_arr_9__1 (d_cache_arr_9__1), .d_arr_9__0 (
                        d_cache_arr_9__0), .d_arr_10__31 (d_cache_arr_10__31), .d_arr_10__30 (
                        d_cache_arr_10__30), .d_arr_10__29 (d_cache_arr_10__29)
                        , .d_arr_10__28 (d_cache_arr_10__28), .d_arr_10__27 (
                        d_cache_arr_10__27), .d_arr_10__26 (d_cache_arr_10__26)
                        , .d_arr_10__25 (d_cache_arr_10__25), .d_arr_10__24 (
                        d_cache_arr_10__24), .d_arr_10__23 (d_cache_arr_10__23)
                        , .d_arr_10__22 (d_cache_arr_10__22), .d_arr_10__21 (
                        d_cache_arr_10__21), .d_arr_10__20 (d_cache_arr_10__20)
                        , .d_arr_10__19 (d_cache_arr_10__19), .d_arr_10__18 (
                        d_cache_arr_10__18), .d_arr_10__17 (d_cache_arr_10__17)
                        , .d_arr_10__16 (d_cache_arr_10__16), .d_arr_10__15 (
                        d_cache_arr_10__15), .d_arr_10__14 (d_cache_arr_10__14)
                        , .d_arr_10__13 (d_cache_arr_10__13), .d_arr_10__12 (
                        d_cache_arr_10__12), .d_arr_10__11 (d_cache_arr_10__11)
                        , .d_arr_10__10 (d_cache_arr_10__10), .d_arr_10__9 (
                        d_cache_arr_10__9), .d_arr_10__8 (d_cache_arr_10__8), .d_arr_10__7 (
                        d_cache_arr_10__7), .d_arr_10__6 (d_cache_arr_10__6), .d_arr_10__5 (
                        d_cache_arr_10__5), .d_arr_10__4 (d_cache_arr_10__4), .d_arr_10__3 (
                        d_cache_arr_10__3), .d_arr_10__2 (d_cache_arr_10__2), .d_arr_10__1 (
                        d_cache_arr_10__1), .d_arr_10__0 (d_cache_arr_10__0), .d_arr_11__31 (
                        d_cache_arr_11__31), .d_arr_11__30 (d_cache_arr_11__30)
                        , .d_arr_11__29 (d_cache_arr_11__29), .d_arr_11__28 (
                        d_cache_arr_11__28), .d_arr_11__27 (d_cache_arr_11__27)
                        , .d_arr_11__26 (d_cache_arr_11__26), .d_arr_11__25 (
                        d_cache_arr_11__25), .d_arr_11__24 (d_cache_arr_11__24)
                        , .d_arr_11__23 (d_cache_arr_11__23), .d_arr_11__22 (
                        d_cache_arr_11__22), .d_arr_11__21 (d_cache_arr_11__21)
                        , .d_arr_11__20 (d_cache_arr_11__20), .d_arr_11__19 (
                        d_cache_arr_11__19), .d_arr_11__18 (d_cache_arr_11__18)
                        , .d_arr_11__17 (d_cache_arr_11__17), .d_arr_11__16 (
                        d_cache_arr_11__16), .d_arr_11__15 (d_cache_arr_11__15)
                        , .d_arr_11__14 (d_cache_arr_11__14), .d_arr_11__13 (
                        d_cache_arr_11__13), .d_arr_11__12 (d_cache_arr_11__12)
                        , .d_arr_11__11 (d_cache_arr_11__11), .d_arr_11__10 (
                        d_cache_arr_11__10), .d_arr_11__9 (d_cache_arr_11__9), .d_arr_11__8 (
                        d_cache_arr_11__8), .d_arr_11__7 (d_cache_arr_11__7), .d_arr_11__6 (
                        d_cache_arr_11__6), .d_arr_11__5 (d_cache_arr_11__5), .d_arr_11__4 (
                        d_cache_arr_11__4), .d_arr_11__3 (d_cache_arr_11__3), .d_arr_11__2 (
                        d_cache_arr_11__2), .d_arr_11__1 (d_cache_arr_11__1), .d_arr_11__0 (
                        d_cache_arr_11__0), .d_arr_12__31 (d_cache_arr_12__31), 
                        .d_arr_12__30 (d_cache_arr_12__30), .d_arr_12__29 (
                        d_cache_arr_12__29), .d_arr_12__28 (d_cache_arr_12__28)
                        , .d_arr_12__27 (d_cache_arr_12__27), .d_arr_12__26 (
                        d_cache_arr_12__26), .d_arr_12__25 (d_cache_arr_12__25)
                        , .d_arr_12__24 (d_cache_arr_12__24), .d_arr_12__23 (
                        d_cache_arr_12__23), .d_arr_12__22 (d_cache_arr_12__22)
                        , .d_arr_12__21 (d_cache_arr_12__21), .d_arr_12__20 (
                        d_cache_arr_12__20), .d_arr_12__19 (d_cache_arr_12__19)
                        , .d_arr_12__18 (d_cache_arr_12__18), .d_arr_12__17 (
                        d_cache_arr_12__17), .d_arr_12__16 (d_cache_arr_12__16)
                        , .d_arr_12__15 (d_cache_arr_12__15), .d_arr_12__14 (
                        d_cache_arr_12__14), .d_arr_12__13 (d_cache_arr_12__13)
                        , .d_arr_12__12 (d_cache_arr_12__12), .d_arr_12__11 (
                        d_cache_arr_12__11), .d_arr_12__10 (d_cache_arr_12__10)
                        , .d_arr_12__9 (d_cache_arr_12__9), .d_arr_12__8 (
                        d_cache_arr_12__8), .d_arr_12__7 (d_cache_arr_12__7), .d_arr_12__6 (
                        d_cache_arr_12__6), .d_arr_12__5 (d_cache_arr_12__5), .d_arr_12__4 (
                        d_cache_arr_12__4), .d_arr_12__3 (d_cache_arr_12__3), .d_arr_12__2 (
                        d_cache_arr_12__2), .d_arr_12__1 (d_cache_arr_12__1), .d_arr_12__0 (
                        d_cache_arr_12__0), .d_arr_13__31 (d_cache_arr_13__31), 
                        .d_arr_13__30 (d_cache_arr_13__30), .d_arr_13__29 (
                        d_cache_arr_13__29), .d_arr_13__28 (d_cache_arr_13__28)
                        , .d_arr_13__27 (d_cache_arr_13__27), .d_arr_13__26 (
                        d_cache_arr_13__26), .d_arr_13__25 (d_cache_arr_13__25)
                        , .d_arr_13__24 (d_cache_arr_13__24), .d_arr_13__23 (
                        d_cache_arr_13__23), .d_arr_13__22 (d_cache_arr_13__22)
                        , .d_arr_13__21 (d_cache_arr_13__21), .d_arr_13__20 (
                        d_cache_arr_13__20), .d_arr_13__19 (d_cache_arr_13__19)
                        , .d_arr_13__18 (d_cache_arr_13__18), .d_arr_13__17 (
                        d_cache_arr_13__17), .d_arr_13__16 (d_cache_arr_13__16)
                        , .d_arr_13__15 (d_cache_arr_13__15), .d_arr_13__14 (
                        d_cache_arr_13__14), .d_arr_13__13 (d_cache_arr_13__13)
                        , .d_arr_13__12 (d_cache_arr_13__12), .d_arr_13__11 (
                        d_cache_arr_13__11), .d_arr_13__10 (d_cache_arr_13__10)
                        , .d_arr_13__9 (d_cache_arr_13__9), .d_arr_13__8 (
                        d_cache_arr_13__8), .d_arr_13__7 (d_cache_arr_13__7), .d_arr_13__6 (
                        d_cache_arr_13__6), .d_arr_13__5 (d_cache_arr_13__5), .d_arr_13__4 (
                        d_cache_arr_13__4), .d_arr_13__3 (d_cache_arr_13__3), .d_arr_13__2 (
                        d_cache_arr_13__2), .d_arr_13__1 (d_cache_arr_13__1), .d_arr_13__0 (
                        d_cache_arr_13__0), .d_arr_14__31 (d_cache_arr_14__31), 
                        .d_arr_14__30 (d_cache_arr_14__30), .d_arr_14__29 (
                        d_cache_arr_14__29), .d_arr_14__28 (d_cache_arr_14__28)
                        , .d_arr_14__27 (d_cache_arr_14__27), .d_arr_14__26 (
                        d_cache_arr_14__26), .d_arr_14__25 (d_cache_arr_14__25)
                        , .d_arr_14__24 (d_cache_arr_14__24), .d_arr_14__23 (
                        d_cache_arr_14__23), .d_arr_14__22 (d_cache_arr_14__22)
                        , .d_arr_14__21 (d_cache_arr_14__21), .d_arr_14__20 (
                        d_cache_arr_14__20), .d_arr_14__19 (d_cache_arr_14__19)
                        , .d_arr_14__18 (d_cache_arr_14__18), .d_arr_14__17 (
                        d_cache_arr_14__17), .d_arr_14__16 (d_cache_arr_14__16)
                        , .d_arr_14__15 (d_cache_arr_14__15), .d_arr_14__14 (
                        d_cache_arr_14__14), .d_arr_14__13 (d_cache_arr_14__13)
                        , .d_arr_14__12 (d_cache_arr_14__12), .d_arr_14__11 (
                        d_cache_arr_14__11), .d_arr_14__10 (d_cache_arr_14__10)
                        , .d_arr_14__9 (d_cache_arr_14__9), .d_arr_14__8 (
                        d_cache_arr_14__8), .d_arr_14__7 (d_cache_arr_14__7), .d_arr_14__6 (
                        d_cache_arr_14__6), .d_arr_14__5 (d_cache_arr_14__5), .d_arr_14__4 (
                        d_cache_arr_14__4), .d_arr_14__3 (d_cache_arr_14__3), .d_arr_14__2 (
                        d_cache_arr_14__2), .d_arr_14__1 (d_cache_arr_14__1), .d_arr_14__0 (
                        d_cache_arr_14__0), .d_arr_15__31 (d_cache_arr_15__31), 
                        .d_arr_15__30 (d_cache_arr_15__30), .d_arr_15__29 (
                        d_cache_arr_15__29), .d_arr_15__28 (d_cache_arr_15__28)
                        , .d_arr_15__27 (d_cache_arr_15__27), .d_arr_15__26 (
                        d_cache_arr_15__26), .d_arr_15__25 (d_cache_arr_15__25)
                        , .d_arr_15__24 (d_cache_arr_15__24), .d_arr_15__23 (
                        d_cache_arr_15__23), .d_arr_15__22 (d_cache_arr_15__22)
                        , .d_arr_15__21 (d_cache_arr_15__21), .d_arr_15__20 (
                        d_cache_arr_15__20), .d_arr_15__19 (d_cache_arr_15__19)
                        , .d_arr_15__18 (d_cache_arr_15__18), .d_arr_15__17 (
                        d_cache_arr_15__17), .d_arr_15__16 (d_cache_arr_15__16)
                        , .d_arr_15__15 (d_cache_arr_15__15), .d_arr_15__14 (
                        d_cache_arr_15__14), .d_arr_15__13 (d_cache_arr_15__13)
                        , .d_arr_15__12 (d_cache_arr_15__12), .d_arr_15__11 (
                        d_cache_arr_15__11), .d_arr_15__10 (d_cache_arr_15__10)
                        , .d_arr_15__9 (d_cache_arr_15__9), .d_arr_15__8 (
                        d_cache_arr_15__8), .d_arr_15__7 (d_cache_arr_15__7), .d_arr_15__6 (
                        d_cache_arr_15__6), .d_arr_15__5 (d_cache_arr_15__5), .d_arr_15__4 (
                        d_cache_arr_15__4), .d_arr_15__3 (d_cache_arr_15__3), .d_arr_15__2 (
                        d_cache_arr_15__2), .d_arr_15__1 (d_cache_arr_15__1), .d_arr_15__0 (
                        d_cache_arr_15__0), .d_arr_16__31 (d_cache_arr_16__31), 
                        .d_arr_16__30 (d_cache_arr_16__30), .d_arr_16__29 (
                        d_cache_arr_16__29), .d_arr_16__28 (d_cache_arr_16__28)
                        , .d_arr_16__27 (d_cache_arr_16__27), .d_arr_16__26 (
                        d_cache_arr_16__26), .d_arr_16__25 (d_cache_arr_16__25)
                        , .d_arr_16__24 (d_cache_arr_16__24), .d_arr_16__23 (
                        d_cache_arr_16__23), .d_arr_16__22 (d_cache_arr_16__22)
                        , .d_arr_16__21 (d_cache_arr_16__21), .d_arr_16__20 (
                        d_cache_arr_16__20), .d_arr_16__19 (d_cache_arr_16__19)
                        , .d_arr_16__18 (d_cache_arr_16__18), .d_arr_16__17 (
                        d_cache_arr_16__17), .d_arr_16__16 (d_cache_arr_16__16)
                        , .d_arr_16__15 (d_cache_arr_16__15), .d_arr_16__14 (
                        d_cache_arr_16__14), .d_arr_16__13 (d_cache_arr_16__13)
                        , .d_arr_16__12 (d_cache_arr_16__12), .d_arr_16__11 (
                        d_cache_arr_16__11), .d_arr_16__10 (d_cache_arr_16__10)
                        , .d_arr_16__9 (d_cache_arr_16__9), .d_arr_16__8 (
                        d_cache_arr_16__8), .d_arr_16__7 (d_cache_arr_16__7), .d_arr_16__6 (
                        d_cache_arr_16__6), .d_arr_16__5 (d_cache_arr_16__5), .d_arr_16__4 (
                        d_cache_arr_16__4), .d_arr_16__3 (d_cache_arr_16__3), .d_arr_16__2 (
                        d_cache_arr_16__2), .d_arr_16__1 (d_cache_arr_16__1), .d_arr_16__0 (
                        d_cache_arr_16__0), .d_arr_17__31 (d_cache_arr_17__31), 
                        .d_arr_17__30 (d_cache_arr_17__30), .d_arr_17__29 (
                        d_cache_arr_17__29), .d_arr_17__28 (d_cache_arr_17__28)
                        , .d_arr_17__27 (d_cache_arr_17__27), .d_arr_17__26 (
                        d_cache_arr_17__26), .d_arr_17__25 (d_cache_arr_17__25)
                        , .d_arr_17__24 (d_cache_arr_17__24), .d_arr_17__23 (
                        d_cache_arr_17__23), .d_arr_17__22 (d_cache_arr_17__22)
                        , .d_arr_17__21 (d_cache_arr_17__21), .d_arr_17__20 (
                        d_cache_arr_17__20), .d_arr_17__19 (d_cache_arr_17__19)
                        , .d_arr_17__18 (d_cache_arr_17__18), .d_arr_17__17 (
                        d_cache_arr_17__17), .d_arr_17__16 (d_cache_arr_17__16)
                        , .d_arr_17__15 (d_cache_arr_17__15), .d_arr_17__14 (
                        d_cache_arr_17__14), .d_arr_17__13 (d_cache_arr_17__13)
                        , .d_arr_17__12 (d_cache_arr_17__12), .d_arr_17__11 (
                        d_cache_arr_17__11), .d_arr_17__10 (d_cache_arr_17__10)
                        , .d_arr_17__9 (d_cache_arr_17__9), .d_arr_17__8 (
                        d_cache_arr_17__8), .d_arr_17__7 (d_cache_arr_17__7), .d_arr_17__6 (
                        d_cache_arr_17__6), .d_arr_17__5 (d_cache_arr_17__5), .d_arr_17__4 (
                        d_cache_arr_17__4), .d_arr_17__3 (d_cache_arr_17__3), .d_arr_17__2 (
                        d_cache_arr_17__2), .d_arr_17__1 (d_cache_arr_17__1), .d_arr_17__0 (
                        d_cache_arr_17__0), .d_arr_18__31 (d_cache_arr_18__31), 
                        .d_arr_18__30 (d_cache_arr_18__30), .d_arr_18__29 (
                        d_cache_arr_18__29), .d_arr_18__28 (d_cache_arr_18__28)
                        , .d_arr_18__27 (d_cache_arr_18__27), .d_arr_18__26 (
                        d_cache_arr_18__26), .d_arr_18__25 (d_cache_arr_18__25)
                        , .d_arr_18__24 (d_cache_arr_18__24), .d_arr_18__23 (
                        d_cache_arr_18__23), .d_arr_18__22 (d_cache_arr_18__22)
                        , .d_arr_18__21 (d_cache_arr_18__21), .d_arr_18__20 (
                        d_cache_arr_18__20), .d_arr_18__19 (d_cache_arr_18__19)
                        , .d_arr_18__18 (d_cache_arr_18__18), .d_arr_18__17 (
                        d_cache_arr_18__17), .d_arr_18__16 (d_cache_arr_18__16)
                        , .d_arr_18__15 (d_cache_arr_18__15), .d_arr_18__14 (
                        d_cache_arr_18__14), .d_arr_18__13 (d_cache_arr_18__13)
                        , .d_arr_18__12 (d_cache_arr_18__12), .d_arr_18__11 (
                        d_cache_arr_18__11), .d_arr_18__10 (d_cache_arr_18__10)
                        , .d_arr_18__9 (d_cache_arr_18__9), .d_arr_18__8 (
                        d_cache_arr_18__8), .d_arr_18__7 (d_cache_arr_18__7), .d_arr_18__6 (
                        d_cache_arr_18__6), .d_arr_18__5 (d_cache_arr_18__5), .d_arr_18__4 (
                        d_cache_arr_18__4), .d_arr_18__3 (d_cache_arr_18__3), .d_arr_18__2 (
                        d_cache_arr_18__2), .d_arr_18__1 (d_cache_arr_18__1), .d_arr_18__0 (
                        d_cache_arr_18__0), .d_arr_19__31 (d_cache_arr_19__31), 
                        .d_arr_19__30 (d_cache_arr_19__30), .d_arr_19__29 (
                        d_cache_arr_19__29), .d_arr_19__28 (d_cache_arr_19__28)
                        , .d_arr_19__27 (d_cache_arr_19__27), .d_arr_19__26 (
                        d_cache_arr_19__26), .d_arr_19__25 (d_cache_arr_19__25)
                        , .d_arr_19__24 (d_cache_arr_19__24), .d_arr_19__23 (
                        d_cache_arr_19__23), .d_arr_19__22 (d_cache_arr_19__22)
                        , .d_arr_19__21 (d_cache_arr_19__21), .d_arr_19__20 (
                        d_cache_arr_19__20), .d_arr_19__19 (d_cache_arr_19__19)
                        , .d_arr_19__18 (d_cache_arr_19__18), .d_arr_19__17 (
                        d_cache_arr_19__17), .d_arr_19__16 (d_cache_arr_19__16)
                        , .d_arr_19__15 (d_cache_arr_19__15), .d_arr_19__14 (
                        d_cache_arr_19__14), .d_arr_19__13 (d_cache_arr_19__13)
                        , .d_arr_19__12 (d_cache_arr_19__12), .d_arr_19__11 (
                        d_cache_arr_19__11), .d_arr_19__10 (d_cache_arr_19__10)
                        , .d_arr_19__9 (d_cache_arr_19__9), .d_arr_19__8 (
                        d_cache_arr_19__8), .d_arr_19__7 (d_cache_arr_19__7), .d_arr_19__6 (
                        d_cache_arr_19__6), .d_arr_19__5 (d_cache_arr_19__5), .d_arr_19__4 (
                        d_cache_arr_19__4), .d_arr_19__3 (d_cache_arr_19__3), .d_arr_19__2 (
                        d_cache_arr_19__2), .d_arr_19__1 (d_cache_arr_19__1), .d_arr_19__0 (
                        d_cache_arr_19__0), .d_arr_20__31 (d_cache_arr_20__31), 
                        .d_arr_20__30 (d_cache_arr_20__30), .d_arr_20__29 (
                        d_cache_arr_20__29), .d_arr_20__28 (d_cache_arr_20__28)
                        , .d_arr_20__27 (d_cache_arr_20__27), .d_arr_20__26 (
                        d_cache_arr_20__26), .d_arr_20__25 (d_cache_arr_20__25)
                        , .d_arr_20__24 (d_cache_arr_20__24), .d_arr_20__23 (
                        d_cache_arr_20__23), .d_arr_20__22 (d_cache_arr_20__22)
                        , .d_arr_20__21 (d_cache_arr_20__21), .d_arr_20__20 (
                        d_cache_arr_20__20), .d_arr_20__19 (d_cache_arr_20__19)
                        , .d_arr_20__18 (d_cache_arr_20__18), .d_arr_20__17 (
                        d_cache_arr_20__17), .d_arr_20__16 (d_cache_arr_20__16)
                        , .d_arr_20__15 (d_cache_arr_20__15), .d_arr_20__14 (
                        d_cache_arr_20__14), .d_arr_20__13 (d_cache_arr_20__13)
                        , .d_arr_20__12 (d_cache_arr_20__12), .d_arr_20__11 (
                        d_cache_arr_20__11), .d_arr_20__10 (d_cache_arr_20__10)
                        , .d_arr_20__9 (d_cache_arr_20__9), .d_arr_20__8 (
                        d_cache_arr_20__8), .d_arr_20__7 (d_cache_arr_20__7), .d_arr_20__6 (
                        d_cache_arr_20__6), .d_arr_20__5 (d_cache_arr_20__5), .d_arr_20__4 (
                        d_cache_arr_20__4), .d_arr_20__3 (d_cache_arr_20__3), .d_arr_20__2 (
                        d_cache_arr_20__2), .d_arr_20__1 (d_cache_arr_20__1), .d_arr_20__0 (
                        d_cache_arr_20__0), .d_arr_21__31 (d_cache_arr_21__31), 
                        .d_arr_21__30 (d_cache_arr_21__30), .d_arr_21__29 (
                        d_cache_arr_21__29), .d_arr_21__28 (d_cache_arr_21__28)
                        , .d_arr_21__27 (d_cache_arr_21__27), .d_arr_21__26 (
                        d_cache_arr_21__26), .d_arr_21__25 (d_cache_arr_21__25)
                        , .d_arr_21__24 (d_cache_arr_21__24), .d_arr_21__23 (
                        d_cache_arr_21__23), .d_arr_21__22 (d_cache_arr_21__22)
                        , .d_arr_21__21 (d_cache_arr_21__21), .d_arr_21__20 (
                        d_cache_arr_21__20), .d_arr_21__19 (d_cache_arr_21__19)
                        , .d_arr_21__18 (d_cache_arr_21__18), .d_arr_21__17 (
                        d_cache_arr_21__17), .d_arr_21__16 (d_cache_arr_21__16)
                        , .d_arr_21__15 (d_cache_arr_21__15), .d_arr_21__14 (
                        d_cache_arr_21__14), .d_arr_21__13 (d_cache_arr_21__13)
                        , .d_arr_21__12 (d_cache_arr_21__12), .d_arr_21__11 (
                        d_cache_arr_21__11), .d_arr_21__10 (d_cache_arr_21__10)
                        , .d_arr_21__9 (d_cache_arr_21__9), .d_arr_21__8 (
                        d_cache_arr_21__8), .d_arr_21__7 (d_cache_arr_21__7), .d_arr_21__6 (
                        d_cache_arr_21__6), .d_arr_21__5 (d_cache_arr_21__5), .d_arr_21__4 (
                        d_cache_arr_21__4), .d_arr_21__3 (d_cache_arr_21__3), .d_arr_21__2 (
                        d_cache_arr_21__2), .d_arr_21__1 (d_cache_arr_21__1), .d_arr_21__0 (
                        d_cache_arr_21__0), .d_arr_22__31 (d_cache_arr_22__31), 
                        .d_arr_22__30 (d_cache_arr_22__30), .d_arr_22__29 (
                        d_cache_arr_22__29), .d_arr_22__28 (d_cache_arr_22__28)
                        , .d_arr_22__27 (d_cache_arr_22__27), .d_arr_22__26 (
                        d_cache_arr_22__26), .d_arr_22__25 (d_cache_arr_22__25)
                        , .d_arr_22__24 (d_cache_arr_22__24), .d_arr_22__23 (
                        d_cache_arr_22__23), .d_arr_22__22 (d_cache_arr_22__22)
                        , .d_arr_22__21 (d_cache_arr_22__21), .d_arr_22__20 (
                        d_cache_arr_22__20), .d_arr_22__19 (d_cache_arr_22__19)
                        , .d_arr_22__18 (d_cache_arr_22__18), .d_arr_22__17 (
                        d_cache_arr_22__17), .d_arr_22__16 (d_cache_arr_22__16)
                        , .d_arr_22__15 (d_cache_arr_22__15), .d_arr_22__14 (
                        d_cache_arr_22__14), .d_arr_22__13 (d_cache_arr_22__13)
                        , .d_arr_22__12 (d_cache_arr_22__12), .d_arr_22__11 (
                        d_cache_arr_22__11), .d_arr_22__10 (d_cache_arr_22__10)
                        , .d_arr_22__9 (d_cache_arr_22__9), .d_arr_22__8 (
                        d_cache_arr_22__8), .d_arr_22__7 (d_cache_arr_22__7), .d_arr_22__6 (
                        d_cache_arr_22__6), .d_arr_22__5 (d_cache_arr_22__5), .d_arr_22__4 (
                        d_cache_arr_22__4), .d_arr_22__3 (d_cache_arr_22__3), .d_arr_22__2 (
                        d_cache_arr_22__2), .d_arr_22__1 (d_cache_arr_22__1), .d_arr_22__0 (
                        d_cache_arr_22__0), .d_arr_23__31 (d_cache_arr_23__31), 
                        .d_arr_23__30 (d_cache_arr_23__30), .d_arr_23__29 (
                        d_cache_arr_23__29), .d_arr_23__28 (d_cache_arr_23__28)
                        , .d_arr_23__27 (d_cache_arr_23__27), .d_arr_23__26 (
                        d_cache_arr_23__26), .d_arr_23__25 (d_cache_arr_23__25)
                        , .d_arr_23__24 (d_cache_arr_23__24), .d_arr_23__23 (
                        d_cache_arr_23__23), .d_arr_23__22 (d_cache_arr_23__22)
                        , .d_arr_23__21 (d_cache_arr_23__21), .d_arr_23__20 (
                        d_cache_arr_23__20), .d_arr_23__19 (d_cache_arr_23__19)
                        , .d_arr_23__18 (d_cache_arr_23__18), .d_arr_23__17 (
                        d_cache_arr_23__17), .d_arr_23__16 (d_cache_arr_23__16)
                        , .d_arr_23__15 (d_cache_arr_23__15), .d_arr_23__14 (
                        d_cache_arr_23__14), .d_arr_23__13 (d_cache_arr_23__13)
                        , .d_arr_23__12 (d_cache_arr_23__12), .d_arr_23__11 (
                        d_cache_arr_23__11), .d_arr_23__10 (d_cache_arr_23__10)
                        , .d_arr_23__9 (d_cache_arr_23__9), .d_arr_23__8 (
                        d_cache_arr_23__8), .d_arr_23__7 (d_cache_arr_23__7), .d_arr_23__6 (
                        d_cache_arr_23__6), .d_arr_23__5 (d_cache_arr_23__5), .d_arr_23__4 (
                        d_cache_arr_23__4), .d_arr_23__3 (d_cache_arr_23__3), .d_arr_23__2 (
                        d_cache_arr_23__2), .d_arr_23__1 (d_cache_arr_23__1), .d_arr_23__0 (
                        d_cache_arr_23__0), .d_arr_24__31 (d_cache_arr_24__31), 
                        .d_arr_24__30 (d_cache_arr_24__30), .d_arr_24__29 (
                        d_cache_arr_24__29), .d_arr_24__28 (d_cache_arr_24__28)
                        , .d_arr_24__27 (d_cache_arr_24__27), .d_arr_24__26 (
                        d_cache_arr_24__26), .d_arr_24__25 (d_cache_arr_24__25)
                        , .d_arr_24__24 (d_cache_arr_24__24), .d_arr_24__23 (
                        d_cache_arr_24__23), .d_arr_24__22 (d_cache_arr_24__22)
                        , .d_arr_24__21 (d_cache_arr_24__21), .d_arr_24__20 (
                        d_cache_arr_24__20), .d_arr_24__19 (d_cache_arr_24__19)
                        , .d_arr_24__18 (d_cache_arr_24__18), .d_arr_24__17 (
                        d_cache_arr_24__17), .d_arr_24__16 (d_cache_arr_24__16)
                        , .d_arr_24__15 (d_cache_arr_24__15), .d_arr_24__14 (
                        d_cache_arr_24__14), .d_arr_24__13 (d_cache_arr_24__13)
                        , .d_arr_24__12 (d_cache_arr_24__12), .d_arr_24__11 (
                        d_cache_arr_24__11), .d_arr_24__10 (d_cache_arr_24__10)
                        , .d_arr_24__9 (d_cache_arr_24__9), .d_arr_24__8 (
                        d_cache_arr_24__8), .d_arr_24__7 (d_cache_arr_24__7), .d_arr_24__6 (
                        d_cache_arr_24__6), .d_arr_24__5 (d_cache_arr_24__5), .d_arr_24__4 (
                        d_cache_arr_24__4), .d_arr_24__3 (d_cache_arr_24__3), .d_arr_24__2 (
                        d_cache_arr_24__2), .d_arr_24__1 (d_cache_arr_24__1), .d_arr_24__0 (
                        d_cache_arr_24__0), .q_arr_0__31 (q_cache_arr_0__31), .q_arr_0__30 (
                        q_cache_arr_0__30), .q_arr_0__29 (q_cache_arr_0__29), .q_arr_0__28 (
                        q_cache_arr_0__28), .q_arr_0__27 (q_cache_arr_0__27), .q_arr_0__26 (
                        q_cache_arr_0__26), .q_arr_0__25 (q_cache_arr_0__25), .q_arr_0__24 (
                        q_cache_arr_0__24), .q_arr_0__23 (q_cache_arr_0__23), .q_arr_0__22 (
                        q_cache_arr_0__22), .q_arr_0__21 (q_cache_arr_0__21), .q_arr_0__20 (
                        q_cache_arr_0__20), .q_arr_0__19 (q_cache_arr_0__19), .q_arr_0__18 (
                        q_cache_arr_0__18), .q_arr_0__17 (q_cache_arr_0__17), .q_arr_0__16 (
                        q_cache_arr_0__16), .q_arr_0__15 (q_cache_arr_0__15), .q_arr_0__14 (
                        q_cache_arr_0__14), .q_arr_0__13 (q_cache_arr_0__13), .q_arr_0__12 (
                        q_cache_arr_0__12), .q_arr_0__11 (q_cache_arr_0__11), .q_arr_0__10 (
                        q_cache_arr_0__10), .q_arr_0__9 (q_cache_arr_0__9), .q_arr_0__8 (
                        q_cache_arr_0__8), .q_arr_0__7 (q_cache_arr_0__7), .q_arr_0__6 (
                        q_cache_arr_0__6), .q_arr_0__5 (q_cache_arr_0__5), .q_arr_0__4 (
                        q_cache_arr_0__4), .q_arr_0__3 (q_cache_arr_0__3), .q_arr_0__2 (
                        q_cache_arr_0__2), .q_arr_0__1 (q_cache_arr_0__1), .q_arr_0__0 (
                        q_cache_arr_0__0), .q_arr_1__31 (q_cache_arr_1__31), .q_arr_1__30 (
                        q_cache_arr_1__30), .q_arr_1__29 (q_cache_arr_1__29), .q_arr_1__28 (
                        q_cache_arr_1__28), .q_arr_1__27 (q_cache_arr_1__27), .q_arr_1__26 (
                        q_cache_arr_1__26), .q_arr_1__25 (q_cache_arr_1__25), .q_arr_1__24 (
                        q_cache_arr_1__24), .q_arr_1__23 (q_cache_arr_1__23), .q_arr_1__22 (
                        q_cache_arr_1__22), .q_arr_1__21 (q_cache_arr_1__21), .q_arr_1__20 (
                        q_cache_arr_1__20), .q_arr_1__19 (q_cache_arr_1__19), .q_arr_1__18 (
                        q_cache_arr_1__18), .q_arr_1__17 (q_cache_arr_1__17), .q_arr_1__16 (
                        q_cache_arr_1__16), .q_arr_1__15 (q_cache_arr_1__15), .q_arr_1__14 (
                        q_cache_arr_1__14), .q_arr_1__13 (q_cache_arr_1__13), .q_arr_1__12 (
                        q_cache_arr_1__12), .q_arr_1__11 (q_cache_arr_1__11), .q_arr_1__10 (
                        q_cache_arr_1__10), .q_arr_1__9 (q_cache_arr_1__9), .q_arr_1__8 (
                        q_cache_arr_1__8), .q_arr_1__7 (q_cache_arr_1__7), .q_arr_1__6 (
                        q_cache_arr_1__6), .q_arr_1__5 (q_cache_arr_1__5), .q_arr_1__4 (
                        q_cache_arr_1__4), .q_arr_1__3 (q_cache_arr_1__3), .q_arr_1__2 (
                        q_cache_arr_1__2), .q_arr_1__1 (q_cache_arr_1__1), .q_arr_1__0 (
                        q_cache_arr_1__0), .q_arr_2__31 (q_cache_arr_2__31), .q_arr_2__30 (
                        q_cache_arr_2__30), .q_arr_2__29 (q_cache_arr_2__29), .q_arr_2__28 (
                        q_cache_arr_2__28), .q_arr_2__27 (q_cache_arr_2__27), .q_arr_2__26 (
                        q_cache_arr_2__26), .q_arr_2__25 (q_cache_arr_2__25), .q_arr_2__24 (
                        q_cache_arr_2__24), .q_arr_2__23 (q_cache_arr_2__23), .q_arr_2__22 (
                        q_cache_arr_2__22), .q_arr_2__21 (q_cache_arr_2__21), .q_arr_2__20 (
                        q_cache_arr_2__20), .q_arr_2__19 (q_cache_arr_2__19), .q_arr_2__18 (
                        q_cache_arr_2__18), .q_arr_2__17 (q_cache_arr_2__17), .q_arr_2__16 (
                        q_cache_arr_2__16), .q_arr_2__15 (q_cache_arr_2__15), .q_arr_2__14 (
                        q_cache_arr_2__14), .q_arr_2__13 (q_cache_arr_2__13), .q_arr_2__12 (
                        q_cache_arr_2__12), .q_arr_2__11 (q_cache_arr_2__11), .q_arr_2__10 (
                        q_cache_arr_2__10), .q_arr_2__9 (q_cache_arr_2__9), .q_arr_2__8 (
                        q_cache_arr_2__8), .q_arr_2__7 (q_cache_arr_2__7), .q_arr_2__6 (
                        q_cache_arr_2__6), .q_arr_2__5 (q_cache_arr_2__5), .q_arr_2__4 (
                        q_cache_arr_2__4), .q_arr_2__3 (q_cache_arr_2__3), .q_arr_2__2 (
                        q_cache_arr_2__2), .q_arr_2__1 (q_cache_arr_2__1), .q_arr_2__0 (
                        q_cache_arr_2__0), .q_arr_3__31 (q_cache_arr_3__31), .q_arr_3__30 (
                        q_cache_arr_3__30), .q_arr_3__29 (q_cache_arr_3__29), .q_arr_3__28 (
                        q_cache_arr_3__28), .q_arr_3__27 (q_cache_arr_3__27), .q_arr_3__26 (
                        q_cache_arr_3__26), .q_arr_3__25 (q_cache_arr_3__25), .q_arr_3__24 (
                        q_cache_arr_3__24), .q_arr_3__23 (q_cache_arr_3__23), .q_arr_3__22 (
                        q_cache_arr_3__22), .q_arr_3__21 (q_cache_arr_3__21), .q_arr_3__20 (
                        q_cache_arr_3__20), .q_arr_3__19 (q_cache_arr_3__19), .q_arr_3__18 (
                        q_cache_arr_3__18), .q_arr_3__17 (q_cache_arr_3__17), .q_arr_3__16 (
                        q_cache_arr_3__16), .q_arr_3__15 (q_cache_arr_3__15), .q_arr_3__14 (
                        q_cache_arr_3__14), .q_arr_3__13 (q_cache_arr_3__13), .q_arr_3__12 (
                        q_cache_arr_3__12), .q_arr_3__11 (q_cache_arr_3__11), .q_arr_3__10 (
                        q_cache_arr_3__10), .q_arr_3__9 (q_cache_arr_3__9), .q_arr_3__8 (
                        q_cache_arr_3__8), .q_arr_3__7 (q_cache_arr_3__7), .q_arr_3__6 (
                        q_cache_arr_3__6), .q_arr_3__5 (q_cache_arr_3__5), .q_arr_3__4 (
                        q_cache_arr_3__4), .q_arr_3__3 (q_cache_arr_3__3), .q_arr_3__2 (
                        q_cache_arr_3__2), .q_arr_3__1 (q_cache_arr_3__1), .q_arr_3__0 (
                        q_cache_arr_3__0), .q_arr_4__31 (q_cache_arr_4__31), .q_arr_4__30 (
                        q_cache_arr_4__30), .q_arr_4__29 (q_cache_arr_4__29), .q_arr_4__28 (
                        q_cache_arr_4__28), .q_arr_4__27 (q_cache_arr_4__27), .q_arr_4__26 (
                        q_cache_arr_4__26), .q_arr_4__25 (q_cache_arr_4__25), .q_arr_4__24 (
                        q_cache_arr_4__24), .q_arr_4__23 (q_cache_arr_4__23), .q_arr_4__22 (
                        q_cache_arr_4__22), .q_arr_4__21 (q_cache_arr_4__21), .q_arr_4__20 (
                        q_cache_arr_4__20), .q_arr_4__19 (q_cache_arr_4__19), .q_arr_4__18 (
                        q_cache_arr_4__18), .q_arr_4__17 (q_cache_arr_4__17), .q_arr_4__16 (
                        q_cache_arr_4__16), .q_arr_4__15 (q_cache_arr_4__15), .q_arr_4__14 (
                        q_cache_arr_4__14), .q_arr_4__13 (q_cache_arr_4__13), .q_arr_4__12 (
                        q_cache_arr_4__12), .q_arr_4__11 (q_cache_arr_4__11), .q_arr_4__10 (
                        q_cache_arr_4__10), .q_arr_4__9 (q_cache_arr_4__9), .q_arr_4__8 (
                        q_cache_arr_4__8), .q_arr_4__7 (q_cache_arr_4__7), .q_arr_4__6 (
                        q_cache_arr_4__6), .q_arr_4__5 (q_cache_arr_4__5), .q_arr_4__4 (
                        q_cache_arr_4__4), .q_arr_4__3 (q_cache_arr_4__3), .q_arr_4__2 (
                        q_cache_arr_4__2), .q_arr_4__1 (q_cache_arr_4__1), .q_arr_4__0 (
                        q_cache_arr_4__0), .q_arr_5__31 (q_cache_arr_5__31), .q_arr_5__30 (
                        q_cache_arr_5__30), .q_arr_5__29 (q_cache_arr_5__29), .q_arr_5__28 (
                        q_cache_arr_5__28), .q_arr_5__27 (q_cache_arr_5__27), .q_arr_5__26 (
                        q_cache_arr_5__26), .q_arr_5__25 (q_cache_arr_5__25), .q_arr_5__24 (
                        q_cache_arr_5__24), .q_arr_5__23 (q_cache_arr_5__23), .q_arr_5__22 (
                        q_cache_arr_5__22), .q_arr_5__21 (q_cache_arr_5__21), .q_arr_5__20 (
                        q_cache_arr_5__20), .q_arr_5__19 (q_cache_arr_5__19), .q_arr_5__18 (
                        q_cache_arr_5__18), .q_arr_5__17 (q_cache_arr_5__17), .q_arr_5__16 (
                        q_cache_arr_5__16), .q_arr_5__15 (q_cache_arr_5__15), .q_arr_5__14 (
                        q_cache_arr_5__14), .q_arr_5__13 (q_cache_arr_5__13), .q_arr_5__12 (
                        q_cache_arr_5__12), .q_arr_5__11 (q_cache_arr_5__11), .q_arr_5__10 (
                        q_cache_arr_5__10), .q_arr_5__9 (q_cache_arr_5__9), .q_arr_5__8 (
                        q_cache_arr_5__8), .q_arr_5__7 (q_cache_arr_5__7), .q_arr_5__6 (
                        q_cache_arr_5__6), .q_arr_5__5 (q_cache_arr_5__5), .q_arr_5__4 (
                        q_cache_arr_5__4), .q_arr_5__3 (q_cache_arr_5__3), .q_arr_5__2 (
                        q_cache_arr_5__2), .q_arr_5__1 (q_cache_arr_5__1), .q_arr_5__0 (
                        q_cache_arr_5__0), .q_arr_6__31 (q_cache_arr_6__31), .q_arr_6__30 (
                        q_cache_arr_6__30), .q_arr_6__29 (q_cache_arr_6__29), .q_arr_6__28 (
                        q_cache_arr_6__28), .q_arr_6__27 (q_cache_arr_6__27), .q_arr_6__26 (
                        q_cache_arr_6__26), .q_arr_6__25 (q_cache_arr_6__25), .q_arr_6__24 (
                        q_cache_arr_6__24), .q_arr_6__23 (q_cache_arr_6__23), .q_arr_6__22 (
                        q_cache_arr_6__22), .q_arr_6__21 (q_cache_arr_6__21), .q_arr_6__20 (
                        q_cache_arr_6__20), .q_arr_6__19 (q_cache_arr_6__19), .q_arr_6__18 (
                        q_cache_arr_6__18), .q_arr_6__17 (q_cache_arr_6__17), .q_arr_6__16 (
                        q_cache_arr_6__16), .q_arr_6__15 (q_cache_arr_6__15), .q_arr_6__14 (
                        q_cache_arr_6__14), .q_arr_6__13 (q_cache_arr_6__13), .q_arr_6__12 (
                        q_cache_arr_6__12), .q_arr_6__11 (q_cache_arr_6__11), .q_arr_6__10 (
                        q_cache_arr_6__10), .q_arr_6__9 (q_cache_arr_6__9), .q_arr_6__8 (
                        q_cache_arr_6__8), .q_arr_6__7 (q_cache_arr_6__7), .q_arr_6__6 (
                        q_cache_arr_6__6), .q_arr_6__5 (q_cache_arr_6__5), .q_arr_6__4 (
                        q_cache_arr_6__4), .q_arr_6__3 (q_cache_arr_6__3), .q_arr_6__2 (
                        q_cache_arr_6__2), .q_arr_6__1 (q_cache_arr_6__1), .q_arr_6__0 (
                        q_cache_arr_6__0), .q_arr_7__31 (q_cache_arr_7__31), .q_arr_7__30 (
                        q_cache_arr_7__30), .q_arr_7__29 (q_cache_arr_7__29), .q_arr_7__28 (
                        q_cache_arr_7__28), .q_arr_7__27 (q_cache_arr_7__27), .q_arr_7__26 (
                        q_cache_arr_7__26), .q_arr_7__25 (q_cache_arr_7__25), .q_arr_7__24 (
                        q_cache_arr_7__24), .q_arr_7__23 (q_cache_arr_7__23), .q_arr_7__22 (
                        q_cache_arr_7__22), .q_arr_7__21 (q_cache_arr_7__21), .q_arr_7__20 (
                        q_cache_arr_7__20), .q_arr_7__19 (q_cache_arr_7__19), .q_arr_7__18 (
                        q_cache_arr_7__18), .q_arr_7__17 (q_cache_arr_7__17), .q_arr_7__16 (
                        q_cache_arr_7__16), .q_arr_7__15 (q_cache_arr_7__15), .q_arr_7__14 (
                        q_cache_arr_7__14), .q_arr_7__13 (q_cache_arr_7__13), .q_arr_7__12 (
                        q_cache_arr_7__12), .q_arr_7__11 (q_cache_arr_7__11), .q_arr_7__10 (
                        q_cache_arr_7__10), .q_arr_7__9 (q_cache_arr_7__9), .q_arr_7__8 (
                        q_cache_arr_7__8), .q_arr_7__7 (q_cache_arr_7__7), .q_arr_7__6 (
                        q_cache_arr_7__6), .q_arr_7__5 (q_cache_arr_7__5), .q_arr_7__4 (
                        q_cache_arr_7__4), .q_arr_7__3 (q_cache_arr_7__3), .q_arr_7__2 (
                        q_cache_arr_7__2), .q_arr_7__1 (q_cache_arr_7__1), .q_arr_7__0 (
                        q_cache_arr_7__0), .q_arr_8__31 (q_cache_arr_8__31), .q_arr_8__30 (
                        q_cache_arr_8__30), .q_arr_8__29 (q_cache_arr_8__29), .q_arr_8__28 (
                        q_cache_arr_8__28), .q_arr_8__27 (q_cache_arr_8__27), .q_arr_8__26 (
                        q_cache_arr_8__26), .q_arr_8__25 (q_cache_arr_8__25), .q_arr_8__24 (
                        q_cache_arr_8__24), .q_arr_8__23 (q_cache_arr_8__23), .q_arr_8__22 (
                        q_cache_arr_8__22), .q_arr_8__21 (q_cache_arr_8__21), .q_arr_8__20 (
                        q_cache_arr_8__20), .q_arr_8__19 (q_cache_arr_8__19), .q_arr_8__18 (
                        q_cache_arr_8__18), .q_arr_8__17 (q_cache_arr_8__17), .q_arr_8__16 (
                        q_cache_arr_8__16), .q_arr_8__15 (q_cache_arr_8__15), .q_arr_8__14 (
                        q_cache_arr_8__14), .q_arr_8__13 (q_cache_arr_8__13), .q_arr_8__12 (
                        q_cache_arr_8__12), .q_arr_8__11 (q_cache_arr_8__11), .q_arr_8__10 (
                        q_cache_arr_8__10), .q_arr_8__9 (q_cache_arr_8__9), .q_arr_8__8 (
                        q_cache_arr_8__8), .q_arr_8__7 (q_cache_arr_8__7), .q_arr_8__6 (
                        q_cache_arr_8__6), .q_arr_8__5 (q_cache_arr_8__5), .q_arr_8__4 (
                        q_cache_arr_8__4), .q_arr_8__3 (q_cache_arr_8__3), .q_arr_8__2 (
                        q_cache_arr_8__2), .q_arr_8__1 (q_cache_arr_8__1), .q_arr_8__0 (
                        q_cache_arr_8__0), .q_arr_9__31 (q_cache_arr_9__31), .q_arr_9__30 (
                        q_cache_arr_9__30), .q_arr_9__29 (q_cache_arr_9__29), .q_arr_9__28 (
                        q_cache_arr_9__28), .q_arr_9__27 (q_cache_arr_9__27), .q_arr_9__26 (
                        q_cache_arr_9__26), .q_arr_9__25 (q_cache_arr_9__25), .q_arr_9__24 (
                        q_cache_arr_9__24), .q_arr_9__23 (q_cache_arr_9__23), .q_arr_9__22 (
                        q_cache_arr_9__22), .q_arr_9__21 (q_cache_arr_9__21), .q_arr_9__20 (
                        q_cache_arr_9__20), .q_arr_9__19 (q_cache_arr_9__19), .q_arr_9__18 (
                        q_cache_arr_9__18), .q_arr_9__17 (q_cache_arr_9__17), .q_arr_9__16 (
                        q_cache_arr_9__16), .q_arr_9__15 (q_cache_arr_9__15), .q_arr_9__14 (
                        q_cache_arr_9__14), .q_arr_9__13 (q_cache_arr_9__13), .q_arr_9__12 (
                        q_cache_arr_9__12), .q_arr_9__11 (q_cache_arr_9__11), .q_arr_9__10 (
                        q_cache_arr_9__10), .q_arr_9__9 (q_cache_arr_9__9), .q_arr_9__8 (
                        q_cache_arr_9__8), .q_arr_9__7 (q_cache_arr_9__7), .q_arr_9__6 (
                        q_cache_arr_9__6), .q_arr_9__5 (q_cache_arr_9__5), .q_arr_9__4 (
                        q_cache_arr_9__4), .q_arr_9__3 (q_cache_arr_9__3), .q_arr_9__2 (
                        q_cache_arr_9__2), .q_arr_9__1 (q_cache_arr_9__1), .q_arr_9__0 (
                        q_cache_arr_9__0), .q_arr_10__31 (q_cache_arr_10__31), .q_arr_10__30 (
                        q_cache_arr_10__30), .q_arr_10__29 (q_cache_arr_10__29)
                        , .q_arr_10__28 (q_cache_arr_10__28), .q_arr_10__27 (
                        q_cache_arr_10__27), .q_arr_10__26 (q_cache_arr_10__26)
                        , .q_arr_10__25 (q_cache_arr_10__25), .q_arr_10__24 (
                        q_cache_arr_10__24), .q_arr_10__23 (q_cache_arr_10__23)
                        , .q_arr_10__22 (q_cache_arr_10__22), .q_arr_10__21 (
                        q_cache_arr_10__21), .q_arr_10__20 (q_cache_arr_10__20)
                        , .q_arr_10__19 (q_cache_arr_10__19), .q_arr_10__18 (
                        q_cache_arr_10__18), .q_arr_10__17 (q_cache_arr_10__17)
                        , .q_arr_10__16 (q_cache_arr_10__16), .q_arr_10__15 (
                        q_cache_arr_10__15), .q_arr_10__14 (q_cache_arr_10__14)
                        , .q_arr_10__13 (q_cache_arr_10__13), .q_arr_10__12 (
                        q_cache_arr_10__12), .q_arr_10__11 (q_cache_arr_10__11)
                        , .q_arr_10__10 (q_cache_arr_10__10), .q_arr_10__9 (
                        q_cache_arr_10__9), .q_arr_10__8 (q_cache_arr_10__8), .q_arr_10__7 (
                        q_cache_arr_10__7), .q_arr_10__6 (q_cache_arr_10__6), .q_arr_10__5 (
                        q_cache_arr_10__5), .q_arr_10__4 (q_cache_arr_10__4), .q_arr_10__3 (
                        q_cache_arr_10__3), .q_arr_10__2 (q_cache_arr_10__2), .q_arr_10__1 (
                        q_cache_arr_10__1), .q_arr_10__0 (q_cache_arr_10__0), .q_arr_11__31 (
                        q_cache_arr_11__31), .q_arr_11__30 (q_cache_arr_11__30)
                        , .q_arr_11__29 (q_cache_arr_11__29), .q_arr_11__28 (
                        q_cache_arr_11__28), .q_arr_11__27 (q_cache_arr_11__27)
                        , .q_arr_11__26 (q_cache_arr_11__26), .q_arr_11__25 (
                        q_cache_arr_11__25), .q_arr_11__24 (q_cache_arr_11__24)
                        , .q_arr_11__23 (q_cache_arr_11__23), .q_arr_11__22 (
                        q_cache_arr_11__22), .q_arr_11__21 (q_cache_arr_11__21)
                        , .q_arr_11__20 (q_cache_arr_11__20), .q_arr_11__19 (
                        q_cache_arr_11__19), .q_arr_11__18 (q_cache_arr_11__18)
                        , .q_arr_11__17 (q_cache_arr_11__17), .q_arr_11__16 (
                        q_cache_arr_11__16), .q_arr_11__15 (q_cache_arr_11__15)
                        , .q_arr_11__14 (q_cache_arr_11__14), .q_arr_11__13 (
                        q_cache_arr_11__13), .q_arr_11__12 (q_cache_arr_11__12)
                        , .q_arr_11__11 (q_cache_arr_11__11), .q_arr_11__10 (
                        q_cache_arr_11__10), .q_arr_11__9 (q_cache_arr_11__9), .q_arr_11__8 (
                        q_cache_arr_11__8), .q_arr_11__7 (q_cache_arr_11__7), .q_arr_11__6 (
                        q_cache_arr_11__6), .q_arr_11__5 (q_cache_arr_11__5), .q_arr_11__4 (
                        q_cache_arr_11__4), .q_arr_11__3 (q_cache_arr_11__3), .q_arr_11__2 (
                        q_cache_arr_11__2), .q_arr_11__1 (q_cache_arr_11__1), .q_arr_11__0 (
                        q_cache_arr_11__0), .q_arr_12__31 (q_cache_arr_12__31), 
                        .q_arr_12__30 (q_cache_arr_12__30), .q_arr_12__29 (
                        q_cache_arr_12__29), .q_arr_12__28 (q_cache_arr_12__28)
                        , .q_arr_12__27 (q_cache_arr_12__27), .q_arr_12__26 (
                        q_cache_arr_12__26), .q_arr_12__25 (q_cache_arr_12__25)
                        , .q_arr_12__24 (q_cache_arr_12__24), .q_arr_12__23 (
                        q_cache_arr_12__23), .q_arr_12__22 (q_cache_arr_12__22)
                        , .q_arr_12__21 (q_cache_arr_12__21), .q_arr_12__20 (
                        q_cache_arr_12__20), .q_arr_12__19 (q_cache_arr_12__19)
                        , .q_arr_12__18 (q_cache_arr_12__18), .q_arr_12__17 (
                        q_cache_arr_12__17), .q_arr_12__16 (q_cache_arr_12__16)
                        , .q_arr_12__15 (q_cache_arr_12__15), .q_arr_12__14 (
                        q_cache_arr_12__14), .q_arr_12__13 (q_cache_arr_12__13)
                        , .q_arr_12__12 (q_cache_arr_12__12), .q_arr_12__11 (
                        q_cache_arr_12__11), .q_arr_12__10 (q_cache_arr_12__10)
                        , .q_arr_12__9 (q_cache_arr_12__9), .q_arr_12__8 (
                        q_cache_arr_12__8), .q_arr_12__7 (q_cache_arr_12__7), .q_arr_12__6 (
                        q_cache_arr_12__6), .q_arr_12__5 (q_cache_arr_12__5), .q_arr_12__4 (
                        q_cache_arr_12__4), .q_arr_12__3 (q_cache_arr_12__3), .q_arr_12__2 (
                        q_cache_arr_12__2), .q_arr_12__1 (q_cache_arr_12__1), .q_arr_12__0 (
                        q_cache_arr_12__0), .q_arr_13__31 (q_cache_arr_13__31), 
                        .q_arr_13__30 (q_cache_arr_13__30), .q_arr_13__29 (
                        q_cache_arr_13__29), .q_arr_13__28 (q_cache_arr_13__28)
                        , .q_arr_13__27 (q_cache_arr_13__27), .q_arr_13__26 (
                        q_cache_arr_13__26), .q_arr_13__25 (q_cache_arr_13__25)
                        , .q_arr_13__24 (q_cache_arr_13__24), .q_arr_13__23 (
                        q_cache_arr_13__23), .q_arr_13__22 (q_cache_arr_13__22)
                        , .q_arr_13__21 (q_cache_arr_13__21), .q_arr_13__20 (
                        q_cache_arr_13__20), .q_arr_13__19 (q_cache_arr_13__19)
                        , .q_arr_13__18 (q_cache_arr_13__18), .q_arr_13__17 (
                        q_cache_arr_13__17), .q_arr_13__16 (q_cache_arr_13__16)
                        , .q_arr_13__15 (q_cache_arr_13__15), .q_arr_13__14 (
                        q_cache_arr_13__14), .q_arr_13__13 (q_cache_arr_13__13)
                        , .q_arr_13__12 (q_cache_arr_13__12), .q_arr_13__11 (
                        q_cache_arr_13__11), .q_arr_13__10 (q_cache_arr_13__10)
                        , .q_arr_13__9 (q_cache_arr_13__9), .q_arr_13__8 (
                        q_cache_arr_13__8), .q_arr_13__7 (q_cache_arr_13__7), .q_arr_13__6 (
                        q_cache_arr_13__6), .q_arr_13__5 (q_cache_arr_13__5), .q_arr_13__4 (
                        q_cache_arr_13__4), .q_arr_13__3 (q_cache_arr_13__3), .q_arr_13__2 (
                        q_cache_arr_13__2), .q_arr_13__1 (q_cache_arr_13__1), .q_arr_13__0 (
                        q_cache_arr_13__0), .q_arr_14__31 (q_cache_arr_14__31), 
                        .q_arr_14__30 (q_cache_arr_14__30), .q_arr_14__29 (
                        q_cache_arr_14__29), .q_arr_14__28 (q_cache_arr_14__28)
                        , .q_arr_14__27 (q_cache_arr_14__27), .q_arr_14__26 (
                        q_cache_arr_14__26), .q_arr_14__25 (q_cache_arr_14__25)
                        , .q_arr_14__24 (q_cache_arr_14__24), .q_arr_14__23 (
                        q_cache_arr_14__23), .q_arr_14__22 (q_cache_arr_14__22)
                        , .q_arr_14__21 (q_cache_arr_14__21), .q_arr_14__20 (
                        q_cache_arr_14__20), .q_arr_14__19 (q_cache_arr_14__19)
                        , .q_arr_14__18 (q_cache_arr_14__18), .q_arr_14__17 (
                        q_cache_arr_14__17), .q_arr_14__16 (q_cache_arr_14__16)
                        , .q_arr_14__15 (q_cache_arr_14__15), .q_arr_14__14 (
                        q_cache_arr_14__14), .q_arr_14__13 (q_cache_arr_14__13)
                        , .q_arr_14__12 (q_cache_arr_14__12), .q_arr_14__11 (
                        q_cache_arr_14__11), .q_arr_14__10 (q_cache_arr_14__10)
                        , .q_arr_14__9 (q_cache_arr_14__9), .q_arr_14__8 (
                        q_cache_arr_14__8), .q_arr_14__7 (q_cache_arr_14__7), .q_arr_14__6 (
                        q_cache_arr_14__6), .q_arr_14__5 (q_cache_arr_14__5), .q_arr_14__4 (
                        q_cache_arr_14__4), .q_arr_14__3 (q_cache_arr_14__3), .q_arr_14__2 (
                        q_cache_arr_14__2), .q_arr_14__1 (q_cache_arr_14__1), .q_arr_14__0 (
                        q_cache_arr_14__0), .q_arr_15__31 (q_cache_arr_15__31), 
                        .q_arr_15__30 (q_cache_arr_15__30), .q_arr_15__29 (
                        q_cache_arr_15__29), .q_arr_15__28 (q_cache_arr_15__28)
                        , .q_arr_15__27 (q_cache_arr_15__27), .q_arr_15__26 (
                        q_cache_arr_15__26), .q_arr_15__25 (q_cache_arr_15__25)
                        , .q_arr_15__24 (q_cache_arr_15__24), .q_arr_15__23 (
                        q_cache_arr_15__23), .q_arr_15__22 (q_cache_arr_15__22)
                        , .q_arr_15__21 (q_cache_arr_15__21), .q_arr_15__20 (
                        q_cache_arr_15__20), .q_arr_15__19 (q_cache_arr_15__19)
                        , .q_arr_15__18 (q_cache_arr_15__18), .q_arr_15__17 (
                        q_cache_arr_15__17), .q_arr_15__16 (q_cache_arr_15__16)
                        , .q_arr_15__15 (q_cache_arr_15__15), .q_arr_15__14 (
                        q_cache_arr_15__14), .q_arr_15__13 (q_cache_arr_15__13)
                        , .q_arr_15__12 (q_cache_arr_15__12), .q_arr_15__11 (
                        q_cache_arr_15__11), .q_arr_15__10 (q_cache_arr_15__10)
                        , .q_arr_15__9 (q_cache_arr_15__9), .q_arr_15__8 (
                        q_cache_arr_15__8), .q_arr_15__7 (q_cache_arr_15__7), .q_arr_15__6 (
                        q_cache_arr_15__6), .q_arr_15__5 (q_cache_arr_15__5), .q_arr_15__4 (
                        q_cache_arr_15__4), .q_arr_15__3 (q_cache_arr_15__3), .q_arr_15__2 (
                        q_cache_arr_15__2), .q_arr_15__1 (q_cache_arr_15__1), .q_arr_15__0 (
                        q_cache_arr_15__0), .q_arr_16__31 (q_cache_arr_16__31), 
                        .q_arr_16__30 (q_cache_arr_16__30), .q_arr_16__29 (
                        q_cache_arr_16__29), .q_arr_16__28 (q_cache_arr_16__28)
                        , .q_arr_16__27 (q_cache_arr_16__27), .q_arr_16__26 (
                        q_cache_arr_16__26), .q_arr_16__25 (q_cache_arr_16__25)
                        , .q_arr_16__24 (q_cache_arr_16__24), .q_arr_16__23 (
                        q_cache_arr_16__23), .q_arr_16__22 (q_cache_arr_16__22)
                        , .q_arr_16__21 (q_cache_arr_16__21), .q_arr_16__20 (
                        q_cache_arr_16__20), .q_arr_16__19 (q_cache_arr_16__19)
                        , .q_arr_16__18 (q_cache_arr_16__18), .q_arr_16__17 (
                        q_cache_arr_16__17), .q_arr_16__16 (q_cache_arr_16__16)
                        , .q_arr_16__15 (q_cache_arr_16__15), .q_arr_16__14 (
                        q_cache_arr_16__14), .q_arr_16__13 (q_cache_arr_16__13)
                        , .q_arr_16__12 (q_cache_arr_16__12), .q_arr_16__11 (
                        q_cache_arr_16__11), .q_arr_16__10 (q_cache_arr_16__10)
                        , .q_arr_16__9 (q_cache_arr_16__9), .q_arr_16__8 (
                        q_cache_arr_16__8), .q_arr_16__7 (q_cache_arr_16__7), .q_arr_16__6 (
                        q_cache_arr_16__6), .q_arr_16__5 (q_cache_arr_16__5), .q_arr_16__4 (
                        q_cache_arr_16__4), .q_arr_16__3 (q_cache_arr_16__3), .q_arr_16__2 (
                        q_cache_arr_16__2), .q_arr_16__1 (q_cache_arr_16__1), .q_arr_16__0 (
                        q_cache_arr_16__0), .q_arr_17__31 (q_cache_arr_17__31), 
                        .q_arr_17__30 (q_cache_arr_17__30), .q_arr_17__29 (
                        q_cache_arr_17__29), .q_arr_17__28 (q_cache_arr_17__28)
                        , .q_arr_17__27 (q_cache_arr_17__27), .q_arr_17__26 (
                        q_cache_arr_17__26), .q_arr_17__25 (q_cache_arr_17__25)
                        , .q_arr_17__24 (q_cache_arr_17__24), .q_arr_17__23 (
                        q_cache_arr_17__23), .q_arr_17__22 (q_cache_arr_17__22)
                        , .q_arr_17__21 (q_cache_arr_17__21), .q_arr_17__20 (
                        q_cache_arr_17__20), .q_arr_17__19 (q_cache_arr_17__19)
                        , .q_arr_17__18 (q_cache_arr_17__18), .q_arr_17__17 (
                        q_cache_arr_17__17), .q_arr_17__16 (q_cache_arr_17__16)
                        , .q_arr_17__15 (q_cache_arr_17__15), .q_arr_17__14 (
                        q_cache_arr_17__14), .q_arr_17__13 (q_cache_arr_17__13)
                        , .q_arr_17__12 (q_cache_arr_17__12), .q_arr_17__11 (
                        q_cache_arr_17__11), .q_arr_17__10 (q_cache_arr_17__10)
                        , .q_arr_17__9 (q_cache_arr_17__9), .q_arr_17__8 (
                        q_cache_arr_17__8), .q_arr_17__7 (q_cache_arr_17__7), .q_arr_17__6 (
                        q_cache_arr_17__6), .q_arr_17__5 (q_cache_arr_17__5), .q_arr_17__4 (
                        q_cache_arr_17__4), .q_arr_17__3 (q_cache_arr_17__3), .q_arr_17__2 (
                        q_cache_arr_17__2), .q_arr_17__1 (q_cache_arr_17__1), .q_arr_17__0 (
                        q_cache_arr_17__0), .q_arr_18__31 (q_cache_arr_18__31), 
                        .q_arr_18__30 (q_cache_arr_18__30), .q_arr_18__29 (
                        q_cache_arr_18__29), .q_arr_18__28 (q_cache_arr_18__28)
                        , .q_arr_18__27 (q_cache_arr_18__27), .q_arr_18__26 (
                        q_cache_arr_18__26), .q_arr_18__25 (q_cache_arr_18__25)
                        , .q_arr_18__24 (q_cache_arr_18__24), .q_arr_18__23 (
                        q_cache_arr_18__23), .q_arr_18__22 (q_cache_arr_18__22)
                        , .q_arr_18__21 (q_cache_arr_18__21), .q_arr_18__20 (
                        q_cache_arr_18__20), .q_arr_18__19 (q_cache_arr_18__19)
                        , .q_arr_18__18 (q_cache_arr_18__18), .q_arr_18__17 (
                        q_cache_arr_18__17), .q_arr_18__16 (q_cache_arr_18__16)
                        , .q_arr_18__15 (q_cache_arr_18__15), .q_arr_18__14 (
                        q_cache_arr_18__14), .q_arr_18__13 (q_cache_arr_18__13)
                        , .q_arr_18__12 (q_cache_arr_18__12), .q_arr_18__11 (
                        q_cache_arr_18__11), .q_arr_18__10 (q_cache_arr_18__10)
                        , .q_arr_18__9 (q_cache_arr_18__9), .q_arr_18__8 (
                        q_cache_arr_18__8), .q_arr_18__7 (q_cache_arr_18__7), .q_arr_18__6 (
                        q_cache_arr_18__6), .q_arr_18__5 (q_cache_arr_18__5), .q_arr_18__4 (
                        q_cache_arr_18__4), .q_arr_18__3 (q_cache_arr_18__3), .q_arr_18__2 (
                        q_cache_arr_18__2), .q_arr_18__1 (q_cache_arr_18__1), .q_arr_18__0 (
                        q_cache_arr_18__0), .q_arr_19__31 (q_cache_arr_19__31), 
                        .q_arr_19__30 (q_cache_arr_19__30), .q_arr_19__29 (
                        q_cache_arr_19__29), .q_arr_19__28 (q_cache_arr_19__28)
                        , .q_arr_19__27 (q_cache_arr_19__27), .q_arr_19__26 (
                        q_cache_arr_19__26), .q_arr_19__25 (q_cache_arr_19__25)
                        , .q_arr_19__24 (q_cache_arr_19__24), .q_arr_19__23 (
                        q_cache_arr_19__23), .q_arr_19__22 (q_cache_arr_19__22)
                        , .q_arr_19__21 (q_cache_arr_19__21), .q_arr_19__20 (
                        q_cache_arr_19__20), .q_arr_19__19 (q_cache_arr_19__19)
                        , .q_arr_19__18 (q_cache_arr_19__18), .q_arr_19__17 (
                        q_cache_arr_19__17), .q_arr_19__16 (q_cache_arr_19__16)
                        , .q_arr_19__15 (q_cache_arr_19__15), .q_arr_19__14 (
                        q_cache_arr_19__14), .q_arr_19__13 (q_cache_arr_19__13)
                        , .q_arr_19__12 (q_cache_arr_19__12), .q_arr_19__11 (
                        q_cache_arr_19__11), .q_arr_19__10 (q_cache_arr_19__10)
                        , .q_arr_19__9 (q_cache_arr_19__9), .q_arr_19__8 (
                        q_cache_arr_19__8), .q_arr_19__7 (q_cache_arr_19__7), .q_arr_19__6 (
                        q_cache_arr_19__6), .q_arr_19__5 (q_cache_arr_19__5), .q_arr_19__4 (
                        q_cache_arr_19__4), .q_arr_19__3 (q_cache_arr_19__3), .q_arr_19__2 (
                        q_cache_arr_19__2), .q_arr_19__1 (q_cache_arr_19__1), .q_arr_19__0 (
                        q_cache_arr_19__0), .q_arr_20__31 (q_cache_arr_20__31), 
                        .q_arr_20__30 (q_cache_arr_20__30), .q_arr_20__29 (
                        q_cache_arr_20__29), .q_arr_20__28 (q_cache_arr_20__28)
                        , .q_arr_20__27 (q_cache_arr_20__27), .q_arr_20__26 (
                        q_cache_arr_20__26), .q_arr_20__25 (q_cache_arr_20__25)
                        , .q_arr_20__24 (q_cache_arr_20__24), .q_arr_20__23 (
                        q_cache_arr_20__23), .q_arr_20__22 (q_cache_arr_20__22)
                        , .q_arr_20__21 (q_cache_arr_20__21), .q_arr_20__20 (
                        q_cache_arr_20__20), .q_arr_20__19 (q_cache_arr_20__19)
                        , .q_arr_20__18 (q_cache_arr_20__18), .q_arr_20__17 (
                        q_cache_arr_20__17), .q_arr_20__16 (q_cache_arr_20__16)
                        , .q_arr_20__15 (q_cache_arr_20__15), .q_arr_20__14 (
                        q_cache_arr_20__14), .q_arr_20__13 (q_cache_arr_20__13)
                        , .q_arr_20__12 (q_cache_arr_20__12), .q_arr_20__11 (
                        q_cache_arr_20__11), .q_arr_20__10 (q_cache_arr_20__10)
                        , .q_arr_20__9 (q_cache_arr_20__9), .q_arr_20__8 (
                        q_cache_arr_20__8), .q_arr_20__7 (q_cache_arr_20__7), .q_arr_20__6 (
                        q_cache_arr_20__6), .q_arr_20__5 (q_cache_arr_20__5), .q_arr_20__4 (
                        q_cache_arr_20__4), .q_arr_20__3 (q_cache_arr_20__3), .q_arr_20__2 (
                        q_cache_arr_20__2), .q_arr_20__1 (q_cache_arr_20__1), .q_arr_20__0 (
                        q_cache_arr_20__0), .q_arr_21__31 (q_cache_arr_21__31), 
                        .q_arr_21__30 (q_cache_arr_21__30), .q_arr_21__29 (
                        q_cache_arr_21__29), .q_arr_21__28 (q_cache_arr_21__28)
                        , .q_arr_21__27 (q_cache_arr_21__27), .q_arr_21__26 (
                        q_cache_arr_21__26), .q_arr_21__25 (q_cache_arr_21__25)
                        , .q_arr_21__24 (q_cache_arr_21__24), .q_arr_21__23 (
                        q_cache_arr_21__23), .q_arr_21__22 (q_cache_arr_21__22)
                        , .q_arr_21__21 (q_cache_arr_21__21), .q_arr_21__20 (
                        q_cache_arr_21__20), .q_arr_21__19 (q_cache_arr_21__19)
                        , .q_arr_21__18 (q_cache_arr_21__18), .q_arr_21__17 (
                        q_cache_arr_21__17), .q_arr_21__16 (q_cache_arr_21__16)
                        , .q_arr_21__15 (q_cache_arr_21__15), .q_arr_21__14 (
                        q_cache_arr_21__14), .q_arr_21__13 (q_cache_arr_21__13)
                        , .q_arr_21__12 (q_cache_arr_21__12), .q_arr_21__11 (
                        q_cache_arr_21__11), .q_arr_21__10 (q_cache_arr_21__10)
                        , .q_arr_21__9 (q_cache_arr_21__9), .q_arr_21__8 (
                        q_cache_arr_21__8), .q_arr_21__7 (q_cache_arr_21__7), .q_arr_21__6 (
                        q_cache_arr_21__6), .q_arr_21__5 (q_cache_arr_21__5), .q_arr_21__4 (
                        q_cache_arr_21__4), .q_arr_21__3 (q_cache_arr_21__3), .q_arr_21__2 (
                        q_cache_arr_21__2), .q_arr_21__1 (q_cache_arr_21__1), .q_arr_21__0 (
                        q_cache_arr_21__0), .q_arr_22__31 (q_cache_arr_22__31), 
                        .q_arr_22__30 (q_cache_arr_22__30), .q_arr_22__29 (
                        q_cache_arr_22__29), .q_arr_22__28 (q_cache_arr_22__28)
                        , .q_arr_22__27 (q_cache_arr_22__27), .q_arr_22__26 (
                        q_cache_arr_22__26), .q_arr_22__25 (q_cache_arr_22__25)
                        , .q_arr_22__24 (q_cache_arr_22__24), .q_arr_22__23 (
                        q_cache_arr_22__23), .q_arr_22__22 (q_cache_arr_22__22)
                        , .q_arr_22__21 (q_cache_arr_22__21), .q_arr_22__20 (
                        q_cache_arr_22__20), .q_arr_22__19 (q_cache_arr_22__19)
                        , .q_arr_22__18 (q_cache_arr_22__18), .q_arr_22__17 (
                        q_cache_arr_22__17), .q_arr_22__16 (q_cache_arr_22__16)
                        , .q_arr_22__15 (q_cache_arr_22__15), .q_arr_22__14 (
                        q_cache_arr_22__14), .q_arr_22__13 (q_cache_arr_22__13)
                        , .q_arr_22__12 (q_cache_arr_22__12), .q_arr_22__11 (
                        q_cache_arr_22__11), .q_arr_22__10 (q_cache_arr_22__10)
                        , .q_arr_22__9 (q_cache_arr_22__9), .q_arr_22__8 (
                        q_cache_arr_22__8), .q_arr_22__7 (q_cache_arr_22__7), .q_arr_22__6 (
                        q_cache_arr_22__6), .q_arr_22__5 (q_cache_arr_22__5), .q_arr_22__4 (
                        q_cache_arr_22__4), .q_arr_22__3 (q_cache_arr_22__3), .q_arr_22__2 (
                        q_cache_arr_22__2), .q_arr_22__1 (q_cache_arr_22__1), .q_arr_22__0 (
                        q_cache_arr_22__0), .q_arr_23__31 (q_cache_arr_23__31), 
                        .q_arr_23__30 (q_cache_arr_23__30), .q_arr_23__29 (
                        q_cache_arr_23__29), .q_arr_23__28 (q_cache_arr_23__28)
                        , .q_arr_23__27 (q_cache_arr_23__27), .q_arr_23__26 (
                        q_cache_arr_23__26), .q_arr_23__25 (q_cache_arr_23__25)
                        , .q_arr_23__24 (q_cache_arr_23__24), .q_arr_23__23 (
                        q_cache_arr_23__23), .q_arr_23__22 (q_cache_arr_23__22)
                        , .q_arr_23__21 (q_cache_arr_23__21), .q_arr_23__20 (
                        q_cache_arr_23__20), .q_arr_23__19 (q_cache_arr_23__19)
                        , .q_arr_23__18 (q_cache_arr_23__18), .q_arr_23__17 (
                        q_cache_arr_23__17), .q_arr_23__16 (q_cache_arr_23__16)
                        , .q_arr_23__15 (q_cache_arr_23__15), .q_arr_23__14 (
                        q_cache_arr_23__14), .q_arr_23__13 (q_cache_arr_23__13)
                        , .q_arr_23__12 (q_cache_arr_23__12), .q_arr_23__11 (
                        q_cache_arr_23__11), .q_arr_23__10 (q_cache_arr_23__10)
                        , .q_arr_23__9 (q_cache_arr_23__9), .q_arr_23__8 (
                        q_cache_arr_23__8), .q_arr_23__7 (q_cache_arr_23__7), .q_arr_23__6 (
                        q_cache_arr_23__6), .q_arr_23__5 (q_cache_arr_23__5), .q_arr_23__4 (
                        q_cache_arr_23__4), .q_arr_23__3 (q_cache_arr_23__3), .q_arr_23__2 (
                        q_cache_arr_23__2), .q_arr_23__1 (q_cache_arr_23__1), .q_arr_23__0 (
                        q_cache_arr_23__0), .q_arr_24__31 (q_cache_arr_24__31), 
                        .q_arr_24__30 (q_cache_arr_24__30), .q_arr_24__29 (
                        q_cache_arr_24__29), .q_arr_24__28 (q_cache_arr_24__28)
                        , .q_arr_24__27 (q_cache_arr_24__27), .q_arr_24__26 (
                        q_cache_arr_24__26), .q_arr_24__25 (q_cache_arr_24__25)
                        , .q_arr_24__24 (q_cache_arr_24__24), .q_arr_24__23 (
                        q_cache_arr_24__23), .q_arr_24__22 (q_cache_arr_24__22)
                        , .q_arr_24__21 (q_cache_arr_24__21), .q_arr_24__20 (
                        q_cache_arr_24__20), .q_arr_24__19 (q_cache_arr_24__19)
                        , .q_arr_24__18 (q_cache_arr_24__18), .q_arr_24__17 (
                        q_cache_arr_24__17), .q_arr_24__16 (q_cache_arr_24__16)
                        , .q_arr_24__15 (q_cache_arr_24__15), .q_arr_24__14 (
                        q_cache_arr_24__14), .q_arr_24__13 (q_cache_arr_24__13)
                        , .q_arr_24__12 (q_cache_arr_24__12), .q_arr_24__11 (
                        q_cache_arr_24__11), .q_arr_24__10 (q_cache_arr_24__10)
                        , .q_arr_24__9 (q_cache_arr_24__9), .q_arr_24__8 (
                        q_cache_arr_24__8), .q_arr_24__7 (q_cache_arr_24__7), .q_arr_24__6 (
                        q_cache_arr_24__6), .q_arr_24__5 (q_cache_arr_24__5), .q_arr_24__4 (
                        q_cache_arr_24__4), .q_arr_24__3 (q_cache_arr_24__3), .q_arr_24__2 (
                        q_cache_arr_24__2), .q_arr_24__1 (q_cache_arr_24__1), .q_arr_24__0 (
                        q_cache_arr_24__0), .output1_init ({output1_init_q_15,
                        output1_init_q_14,output1_init_q_13,output1_init_q_12,
                        output1_init_q_11,output1_init_q_10,output1_init_q_9,
                        output1_init_q_8,output1_init_q_7,output1_init_q_6,
                        output1_init_q_5,output1_init_q_4,output1_init_q_3,
                        output1_init_q_2,output1_init_q_1,output1_init_q_0}), .output2_init (
                        {output2_init_q_15,output2_init_q_14,output2_init_q_13,
                        output2_init_q_12,output2_init_q_11,output2_init_q_10,
                        output2_init_q_9,output2_init_q_8,output2_init_q_7,
                        output2_init_q_6,output2_init_q_5,output2_init_q_4,
                        output2_init_q_3,output2_init_q_2,output2_init_q_1,
                        output2_init_q_0}), .filter_size (nx1119), .operation (
                        operation_q), .compute_relu (compute_relu_q), .clk (clk)
                        , .en (comp_pipe_en), .reset (comp_pipe_rst), .buffer_ready (
                        buffer_ready_tmp), .semi_ready (semi_ready), .ready (
                        ready_tmp)) ;
    Queue_5_unfolded2 gen_img_window_gen_queues_0_queuei (.d ({
                      img_data_col_0[15],img_data_col_0[14],img_data_col_0[13],
                      img_data_col_0[12],img_data_col_0[11],img_data_col_0[10],
                      img_data_col_0[9],img_data_col_0[8],img_data_col_0[7],
                      img_data_col_0[6],img_data_col_0[5],img_data_col_0[4],
                      img_data_col_0[3],img_data_col_0[2],img_data_col_0[1],
                      img_data_col_0[0]}), .q_0__15 (img_data_0__15), .q_0__14 (
                      img_data_0__14), .q_0__13 (img_data_0__13), .q_0__12 (
                      img_data_0__12), .q_0__11 (img_data_0__11), .q_0__10 (
                      img_data_0__10), .q_0__9 (img_data_0__9), .q_0__8 (
                      img_data_0__8), .q_0__7 (img_data_0__7), .q_0__6 (
                      img_data_0__6), .q_0__5 (img_data_0__5), .q_0__4 (
                      img_data_0__4), .q_0__3 (img_data_0__3), .q_0__2 (
                      img_data_0__2), .q_0__1 (img_data_0__1), .q_0__0 (
                      img_data_0__0), .q_1__15 (img_data_1__15), .q_1__14 (
                      img_data_1__14), .q_1__13 (img_data_1__13), .q_1__12 (
                      img_data_1__12), .q_1__11 (img_data_1__11), .q_1__10 (
                      img_data_1__10), .q_1__9 (img_data_1__9), .q_1__8 (
                      img_data_1__8), .q_1__7 (img_data_1__7), .q_1__6 (
                      img_data_1__6), .q_1__5 (img_data_1__5), .q_1__4 (
                      img_data_1__4), .q_1__3 (img_data_1__3), .q_1__2 (
                      img_data_1__2), .q_1__1 (img_data_1__1), .q_1__0 (
                      img_data_1__0), .q_2__15 (img_data_2__15), .q_2__14 (
                      img_data_2__14), .q_2__13 (img_data_2__13), .q_2__12 (
                      img_data_2__12), .q_2__11 (img_data_2__11), .q_2__10 (
                      img_data_2__10), .q_2__9 (img_data_2__9), .q_2__8 (
                      img_data_2__8), .q_2__7 (img_data_2__7), .q_2__6 (
                      img_data_2__6), .q_2__5 (img_data_2__5), .q_2__4 (
                      img_data_2__4), .q_2__3 (img_data_2__3), .q_2__2 (
                      img_data_2__2), .q_2__1 (img_data_2__1), .q_2__0 (
                      img_data_2__0), .q_3__15 (img_data_3__15), .q_3__14 (
                      img_data_3__14), .q_3__13 (img_data_3__13), .q_3__12 (
                      img_data_3__12), .q_3__11 (img_data_3__11), .q_3__10 (
                      img_data_3__10), .q_3__9 (img_data_3__9), .q_3__8 (
                      img_data_3__8), .q_3__7 (img_data_3__7), .q_3__6 (
                      img_data_3__6), .q_3__5 (img_data_3__5), .q_3__4 (
                      img_data_3__4), .q_3__3 (img_data_3__3), .q_3__2 (
                      img_data_3__2), .q_3__1 (img_data_3__1), .q_3__0 (
                      img_data_3__0), .q_4__15 (img_data_4__15), .q_4__14 (
                      img_data_4__14), .q_4__13 (img_data_4__13), .q_4__12 (
                      img_data_4__12), .q_4__11 (img_data_4__11), .q_4__10 (
                      img_data_4__10), .q_4__9 (img_data_4__9), .q_4__8 (
                      img_data_4__8), .q_4__7 (img_data_4__7), .q_4__6 (
                      img_data_4__6), .q_4__5 (img_data_4__5), .q_4__4 (
                      img_data_4__4), .q_4__3 (img_data_4__3), .q_4__2 (
                      img_data_4__2), .q_4__1 (img_data_4__1), .q_4__0 (
                      img_data_4__0), .clk (nx1181), .load (nx1177), .reset (
                      buffer_ready)) ;
    Queue_5_unfolded2 gen_img_window_gen_queues_1_queuei (.d ({
                      img_data_col_1[15],img_data_col_1[14],img_data_col_1[13],
                      img_data_col_1[12],img_data_col_1[11],img_data_col_1[10],
                      img_data_col_1[9],img_data_col_1[8],img_data_col_1[7],
                      img_data_col_1[6],img_data_col_1[5],img_data_col_1[4],
                      img_data_col_1[3],img_data_col_1[2],img_data_col_1[1],
                      img_data_col_1[0]}), .q_0__15 (img_data_5__15), .q_0__14 (
                      img_data_5__14), .q_0__13 (img_data_5__13), .q_0__12 (
                      img_data_5__12), .q_0__11 (img_data_5__11), .q_0__10 (
                      img_data_5__10), .q_0__9 (img_data_5__9), .q_0__8 (
                      img_data_5__8), .q_0__7 (img_data_5__7), .q_0__6 (
                      img_data_5__6), .q_0__5 (img_data_5__5), .q_0__4 (
                      img_data_5__4), .q_0__3 (img_data_5__3), .q_0__2 (
                      img_data_5__2), .q_0__1 (img_data_5__1), .q_0__0 (
                      img_data_5__0), .q_1__15 (img_data_6__15), .q_1__14 (
                      img_data_6__14), .q_1__13 (img_data_6__13), .q_1__12 (
                      img_data_6__12), .q_1__11 (img_data_6__11), .q_1__10 (
                      img_data_6__10), .q_1__9 (img_data_6__9), .q_1__8 (
                      img_data_6__8), .q_1__7 (img_data_6__7), .q_1__6 (
                      img_data_6__6), .q_1__5 (img_data_6__5), .q_1__4 (
                      img_data_6__4), .q_1__3 (img_data_6__3), .q_1__2 (
                      img_data_6__2), .q_1__1 (img_data_6__1), .q_1__0 (
                      img_data_6__0), .q_2__15 (img_data_7__15), .q_2__14 (
                      img_data_7__14), .q_2__13 (img_data_7__13), .q_2__12 (
                      img_data_7__12), .q_2__11 (img_data_7__11), .q_2__10 (
                      img_data_7__10), .q_2__9 (img_data_7__9), .q_2__8 (
                      img_data_7__8), .q_2__7 (img_data_7__7), .q_2__6 (
                      img_data_7__6), .q_2__5 (img_data_7__5), .q_2__4 (
                      img_data_7__4), .q_2__3 (img_data_7__3), .q_2__2 (
                      img_data_7__2), .q_2__1 (img_data_7__1), .q_2__0 (
                      img_data_7__0), .q_3__15 (img_data_8__15), .q_3__14 (
                      img_data_8__14), .q_3__13 (img_data_8__13), .q_3__12 (
                      img_data_8__12), .q_3__11 (img_data_8__11), .q_3__10 (
                      img_data_8__10), .q_3__9 (img_data_8__9), .q_3__8 (
                      img_data_8__8), .q_3__7 (img_data_8__7), .q_3__6 (
                      img_data_8__6), .q_3__5 (img_data_8__5), .q_3__4 (
                      img_data_8__4), .q_3__3 (img_data_8__3), .q_3__2 (
                      img_data_8__2), .q_3__1 (img_data_8__1), .q_3__0 (
                      img_data_8__0), .q_4__15 (img_data_9__15), .q_4__14 (
                      img_data_9__14), .q_4__13 (img_data_9__13), .q_4__12 (
                      img_data_9__12), .q_4__11 (img_data_9__11), .q_4__10 (
                      img_data_9__10), .q_4__9 (img_data_9__9), .q_4__8 (
                      img_data_9__8), .q_4__7 (img_data_9__7), .q_4__6 (
                      img_data_9__6), .q_4__5 (img_data_9__5), .q_4__4 (
                      img_data_9__4), .q_4__3 (img_data_9__3), .q_4__2 (
                      img_data_9__2), .q_4__1 (img_data_9__1), .q_4__0 (
                      img_data_9__0), .clk (nx1181), .load (nx1177), .reset (
                      buffer_ready)) ;
    Queue_5_unfolded2 gen_img_window_gen_queues_2_queuei (.d ({
                      img_data_col_2[15],img_data_col_2[14],img_data_col_2[13],
                      img_data_col_2[12],img_data_col_2[11],img_data_col_2[10],
                      img_data_col_2[9],img_data_col_2[8],img_data_col_2[7],
                      img_data_col_2[6],img_data_col_2[5],img_data_col_2[4],
                      img_data_col_2[3],img_data_col_2[2],img_data_col_2[1],
                      img_data_col_2[0]}), .q_0__15 (img_data_10__15), .q_0__14 (
                      img_data_10__14), .q_0__13 (img_data_10__13), .q_0__12 (
                      img_data_10__12), .q_0__11 (img_data_10__11), .q_0__10 (
                      img_data_10__10), .q_0__9 (img_data_10__9), .q_0__8 (
                      img_data_10__8), .q_0__7 (img_data_10__7), .q_0__6 (
                      img_data_10__6), .q_0__5 (img_data_10__5), .q_0__4 (
                      img_data_10__4), .q_0__3 (img_data_10__3), .q_0__2 (
                      img_data_10__2), .q_0__1 (img_data_10__1), .q_0__0 (
                      img_data_10__0), .q_1__15 (img_data_11__15), .q_1__14 (
                      img_data_11__14), .q_1__13 (img_data_11__13), .q_1__12 (
                      img_data_11__12), .q_1__11 (img_data_11__11), .q_1__10 (
                      img_data_11__10), .q_1__9 (img_data_11__9), .q_1__8 (
                      img_data_11__8), .q_1__7 (img_data_11__7), .q_1__6 (
                      img_data_11__6), .q_1__5 (img_data_11__5), .q_1__4 (
                      img_data_11__4), .q_1__3 (img_data_11__3), .q_1__2 (
                      img_data_11__2), .q_1__1 (img_data_11__1), .q_1__0 (
                      img_data_11__0), .q_2__15 (img_data_12__15), .q_2__14 (
                      img_data_12__14), .q_2__13 (img_data_12__13), .q_2__12 (
                      img_data_12__12), .q_2__11 (img_data_12__11), .q_2__10 (
                      img_data_12__10), .q_2__9 (img_data_12__9), .q_2__8 (
                      img_data_12__8), .q_2__7 (img_data_12__7), .q_2__6 (
                      img_data_12__6), .q_2__5 (img_data_12__5), .q_2__4 (
                      img_data_12__4), .q_2__3 (img_data_12__3), .q_2__2 (
                      img_data_12__2), .q_2__1 (img_data_12__1), .q_2__0 (
                      img_data_12__0), .q_3__15 (img_data_13__15), .q_3__14 (
                      img_data_13__14), .q_3__13 (img_data_13__13), .q_3__12 (
                      img_data_13__12), .q_3__11 (img_data_13__11), .q_3__10 (
                      img_data_13__10), .q_3__9 (img_data_13__9), .q_3__8 (
                      img_data_13__8), .q_3__7 (img_data_13__7), .q_3__6 (
                      img_data_13__6), .q_3__5 (img_data_13__5), .q_3__4 (
                      img_data_13__4), .q_3__3 (img_data_13__3), .q_3__2 (
                      img_data_13__2), .q_3__1 (img_data_13__1), .q_3__0 (
                      img_data_13__0), .q_4__15 (img_data_14__15), .q_4__14 (
                      img_data_14__14), .q_4__13 (img_data_14__13), .q_4__12 (
                      img_data_14__12), .q_4__11 (img_data_14__11), .q_4__10 (
                      img_data_14__10), .q_4__9 (img_data_14__9), .q_4__8 (
                      img_data_14__8), .q_4__7 (img_data_14__7), .q_4__6 (
                      img_data_14__6), .q_4__5 (img_data_14__5), .q_4__4 (
                      img_data_14__4), .q_4__3 (img_data_14__3), .q_4__2 (
                      img_data_14__2), .q_4__1 (img_data_14__1), .q_4__0 (
                      img_data_14__0), .clk (nx1181), .load (nx1177), .reset (
                      buffer_ready)) ;
    Queue_5_unfolded2 gen_img_window_gen_queues_3_queuei (.d ({
                      img_data_col_3[15],img_data_col_3[14],img_data_col_3[13],
                      img_data_col_3[12],img_data_col_3[11],img_data_col_3[10],
                      img_data_col_3[9],img_data_col_3[8],img_data_col_3[7],
                      img_data_col_3[6],img_data_col_3[5],img_data_col_3[4],
                      img_data_col_3[3],img_data_col_3[2],img_data_col_3[1],
                      img_data_col_3[0]}), .q_0__15 (img_data_15__15), .q_0__14 (
                      img_data_15__14), .q_0__13 (img_data_15__13), .q_0__12 (
                      img_data_15__12), .q_0__11 (img_data_15__11), .q_0__10 (
                      img_data_15__10), .q_0__9 (img_data_15__9), .q_0__8 (
                      img_data_15__8), .q_0__7 (img_data_15__7), .q_0__6 (
                      img_data_15__6), .q_0__5 (img_data_15__5), .q_0__4 (
                      img_data_15__4), .q_0__3 (img_data_15__3), .q_0__2 (
                      img_data_15__2), .q_0__1 (img_data_15__1), .q_0__0 (
                      img_data_15__0), .q_1__15 (img_data_16__15), .q_1__14 (
                      img_data_16__14), .q_1__13 (img_data_16__13), .q_1__12 (
                      img_data_16__12), .q_1__11 (img_data_16__11), .q_1__10 (
                      img_data_16__10), .q_1__9 (img_data_16__9), .q_1__8 (
                      img_data_16__8), .q_1__7 (img_data_16__7), .q_1__6 (
                      img_data_16__6), .q_1__5 (img_data_16__5), .q_1__4 (
                      img_data_16__4), .q_1__3 (img_data_16__3), .q_1__2 (
                      img_data_16__2), .q_1__1 (img_data_16__1), .q_1__0 (
                      img_data_16__0), .q_2__15 (img_data_17__15), .q_2__14 (
                      img_data_17__14), .q_2__13 (img_data_17__13), .q_2__12 (
                      img_data_17__12), .q_2__11 (img_data_17__11), .q_2__10 (
                      img_data_17__10), .q_2__9 (img_data_17__9), .q_2__8 (
                      img_data_17__8), .q_2__7 (img_data_17__7), .q_2__6 (
                      img_data_17__6), .q_2__5 (img_data_17__5), .q_2__4 (
                      img_data_17__4), .q_2__3 (img_data_17__3), .q_2__2 (
                      img_data_17__2), .q_2__1 (img_data_17__1), .q_2__0 (
                      img_data_17__0), .q_3__15 (img_data_18__15), .q_3__14 (
                      img_data_18__14), .q_3__13 (img_data_18__13), .q_3__12 (
                      img_data_18__12), .q_3__11 (img_data_18__11), .q_3__10 (
                      img_data_18__10), .q_3__9 (img_data_18__9), .q_3__8 (
                      img_data_18__8), .q_3__7 (img_data_18__7), .q_3__6 (
                      img_data_18__6), .q_3__5 (img_data_18__5), .q_3__4 (
                      img_data_18__4), .q_3__3 (img_data_18__3), .q_3__2 (
                      img_data_18__2), .q_3__1 (img_data_18__1), .q_3__0 (
                      img_data_18__0), .q_4__15 (img_data_19__15), .q_4__14 (
                      img_data_19__14), .q_4__13 (img_data_19__13), .q_4__12 (
                      img_data_19__12), .q_4__11 (img_data_19__11), .q_4__10 (
                      img_data_19__10), .q_4__9 (img_data_19__9), .q_4__8 (
                      img_data_19__8), .q_4__7 (img_data_19__7), .q_4__6 (
                      img_data_19__6), .q_4__5 (img_data_19__5), .q_4__4 (
                      img_data_19__4), .q_4__3 (img_data_19__3), .q_4__2 (
                      img_data_19__2), .q_4__1 (img_data_19__1), .q_4__0 (
                      img_data_19__0), .clk (nx1183), .load (nx1179), .reset (
                      buffer_ready)) ;
    Queue_5_unfolded2 gen_img_window_gen_queues_4_queuei (.d ({
                      img_data_col_4[15],img_data_col_4[14],img_data_col_4[13],
                      img_data_col_4[12],img_data_col_4[11],img_data_col_4[10],
                      img_data_col_4[9],img_data_col_4[8],img_data_col_4[7],
                      img_data_col_4[6],img_data_col_4[5],img_data_col_4[4],
                      img_data_col_4[3],img_data_col_4[2],img_data_col_4[1],
                      img_data_col_4[0]}), .q_0__15 (img_data_20__15), .q_0__14 (
                      img_data_20__14), .q_0__13 (img_data_20__13), .q_0__12 (
                      img_data_20__12), .q_0__11 (img_data_20__11), .q_0__10 (
                      img_data_20__10), .q_0__9 (img_data_20__9), .q_0__8 (
                      img_data_20__8), .q_0__7 (img_data_20__7), .q_0__6 (
                      img_data_20__6), .q_0__5 (img_data_20__5), .q_0__4 (
                      img_data_20__4), .q_0__3 (img_data_20__3), .q_0__2 (
                      img_data_20__2), .q_0__1 (img_data_20__1), .q_0__0 (
                      img_data_20__0), .q_1__15 (img_data_21__15), .q_1__14 (
                      img_data_21__14), .q_1__13 (img_data_21__13), .q_1__12 (
                      img_data_21__12), .q_1__11 (img_data_21__11), .q_1__10 (
                      img_data_21__10), .q_1__9 (img_data_21__9), .q_1__8 (
                      img_data_21__8), .q_1__7 (img_data_21__7), .q_1__6 (
                      img_data_21__6), .q_1__5 (img_data_21__5), .q_1__4 (
                      img_data_21__4), .q_1__3 (img_data_21__3), .q_1__2 (
                      img_data_21__2), .q_1__1 (img_data_21__1), .q_1__0 (
                      img_data_21__0), .q_2__15 (img_data_22__15), .q_2__14 (
                      img_data_22__14), .q_2__13 (img_data_22__13), .q_2__12 (
                      img_data_22__12), .q_2__11 (img_data_22__11), .q_2__10 (
                      img_data_22__10), .q_2__9 (img_data_22__9), .q_2__8 (
                      img_data_22__8), .q_2__7 (img_data_22__7), .q_2__6 (
                      img_data_22__6), .q_2__5 (img_data_22__5), .q_2__4 (
                      img_data_22__4), .q_2__3 (img_data_22__3), .q_2__2 (
                      img_data_22__2), .q_2__1 (img_data_22__1), .q_2__0 (
                      img_data_22__0), .q_3__15 (img_data_23__15), .q_3__14 (
                      img_data_23__14), .q_3__13 (img_data_23__13), .q_3__12 (
                      img_data_23__12), .q_3__11 (img_data_23__11), .q_3__10 (
                      img_data_23__10), .q_3__9 (img_data_23__9), .q_3__8 (
                      img_data_23__8), .q_3__7 (img_data_23__7), .q_3__6 (
                      img_data_23__6), .q_3__5 (img_data_23__5), .q_3__4 (
                      img_data_23__4), .q_3__3 (img_data_23__3), .q_3__2 (
                      img_data_23__2), .q_3__1 (img_data_23__1), .q_3__0 (
                      img_data_23__0), .q_4__15 (img_data_24__15), .q_4__14 (
                      img_data_24__14), .q_4__13 (img_data_24__13), .q_4__12 (
                      img_data_24__12), .q_4__11 (img_data_24__11), .q_4__10 (
                      img_data_24__10), .q_4__9 (img_data_24__9), .q_4__8 (
                      img_data_24__8), .q_4__7 (img_data_24__7), .q_4__6 (
                      img_data_24__6), .q_4__5 (img_data_24__5), .q_4__4 (
                      img_data_24__4), .q_4__3 (img_data_24__3), .q_4__2 (
                      img_data_24__2), .q_4__1 (img_data_24__1), .q_4__0 (
                      img_data_24__0), .clk (nx1183), .load (nx1179), .reset (
                      buffer_ready)) ;
    Queue_25 gen_filter_window_queuei (.d ({filter_data_word[15],
             filter_data_word[14],filter_data_word[13],filter_data_word[12],
             filter_data_word[11],filter_data_word[10],filter_data_word[9],
             filter_data_word[8],filter_data_word[7],filter_data_word[6],
             filter_data_word[5],filter_data_word[4],filter_data_word[3],
             filter_data_word[2],filter_data_word[1],filter_data_word[0]}), .q_0__15 (
             filter_data_0__15), .q_0__14 (filter_data_0__14), .q_0__13 (
             filter_data_0__13), .q_0__12 (filter_data_0__12), .q_0__11 (
             filter_data_0__11), .q_0__10 (filter_data_0__10), .q_0__9 (
             filter_data_0__9), .q_0__8 (filter_data_0__8), .q_0__7 (
             filter_data_0__7), .q_0__6 (filter_data_0__6), .q_0__5 (
             filter_data_0__5), .q_0__4 (filter_data_0__4), .q_0__3 (
             filter_data_0__3), .q_0__2 (filter_data_0__2), .q_0__1 (
             filter_data_0__1), .q_0__0 (filter_data_0__0), .q_1__15 (
             filter_data_1__15), .q_1__14 (filter_data_1__14), .q_1__13 (
             filter_data_1__13), .q_1__12 (filter_data_1__12), .q_1__11 (
             filter_data_1__11), .q_1__10 (filter_data_1__10), .q_1__9 (
             filter_data_1__9), .q_1__8 (filter_data_1__8), .q_1__7 (
             filter_data_1__7), .q_1__6 (filter_data_1__6), .q_1__5 (
             filter_data_1__5), .q_1__4 (filter_data_1__4), .q_1__3 (
             filter_data_1__3), .q_1__2 (filter_data_1__2), .q_1__1 (
             filter_data_1__1), .q_1__0 (filter_data_1__0), .q_2__15 (
             filter_data_2__15), .q_2__14 (filter_data_2__14), .q_2__13 (
             filter_data_2__13), .q_2__12 (filter_data_2__12), .q_2__11 (
             filter_data_2__11), .q_2__10 (filter_data_2__10), .q_2__9 (
             filter_data_2__9), .q_2__8 (filter_data_2__8), .q_2__7 (
             filter_data_2__7), .q_2__6 (filter_data_2__6), .q_2__5 (
             filter_data_2__5), .q_2__4 (filter_data_2__4), .q_2__3 (
             filter_data_2__3), .q_2__2 (filter_data_2__2), .q_2__1 (
             filter_data_2__1), .q_2__0 (filter_data_2__0), .q_3__15 (
             filter_data_3__15), .q_3__14 (filter_data_3__14), .q_3__13 (
             filter_data_3__13), .q_3__12 (filter_data_3__12), .q_3__11 (
             filter_data_3__11), .q_3__10 (filter_data_3__10), .q_3__9 (
             filter_data_3__9), .q_3__8 (filter_data_3__8), .q_3__7 (
             filter_data_3__7), .q_3__6 (filter_data_3__6), .q_3__5 (
             filter_data_3__5), .q_3__4 (filter_data_3__4), .q_3__3 (
             filter_data_3__3), .q_3__2 (filter_data_3__2), .q_3__1 (
             filter_data_3__1), .q_3__0 (filter_data_3__0), .q_4__15 (
             filter_data_4__15), .q_4__14 (filter_data_4__14), .q_4__13 (
             filter_data_4__13), .q_4__12 (filter_data_4__12), .q_4__11 (
             filter_data_4__11), .q_4__10 (filter_data_4__10), .q_4__9 (
             filter_data_4__9), .q_4__8 (filter_data_4__8), .q_4__7 (
             filter_data_4__7), .q_4__6 (filter_data_4__6), .q_4__5 (
             filter_data_4__5), .q_4__4 (filter_data_4__4), .q_4__3 (
             filter_data_4__3), .q_4__2 (filter_data_4__2), .q_4__1 (
             filter_data_4__1), .q_4__0 (filter_data_4__0), .q_5__15 (
             filter_data_5__15), .q_5__14 (filter_data_5__14), .q_5__13 (
             filter_data_5__13), .q_5__12 (filter_data_5__12), .q_5__11 (
             filter_data_5__11), .q_5__10 (filter_data_5__10), .q_5__9 (
             filter_data_5__9), .q_5__8 (filter_data_5__8), .q_5__7 (
             filter_data_5__7), .q_5__6 (filter_data_5__6), .q_5__5 (
             filter_data_5__5), .q_5__4 (filter_data_5__4), .q_5__3 (
             filter_data_5__3), .q_5__2 (filter_data_5__2), .q_5__1 (
             filter_data_5__1), .q_5__0 (filter_data_5__0), .q_6__15 (
             filter_data_6__15), .q_6__14 (filter_data_6__14), .q_6__13 (
             filter_data_6__13), .q_6__12 (filter_data_6__12), .q_6__11 (
             filter_data_6__11), .q_6__10 (filter_data_6__10), .q_6__9 (
             filter_data_6__9), .q_6__8 (filter_data_6__8), .q_6__7 (
             filter_data_6__7), .q_6__6 (filter_data_6__6), .q_6__5 (
             filter_data_6__5), .q_6__4 (filter_data_6__4), .q_6__3 (
             filter_data_6__3), .q_6__2 (filter_data_6__2), .q_6__1 (
             filter_data_6__1), .q_6__0 (filter_data_6__0), .q_7__15 (
             filter_data_7__15), .q_7__14 (filter_data_7__14), .q_7__13 (
             filter_data_7__13), .q_7__12 (filter_data_7__12), .q_7__11 (
             filter_data_7__11), .q_7__10 (filter_data_7__10), .q_7__9 (
             filter_data_7__9), .q_7__8 (filter_data_7__8), .q_7__7 (
             filter_data_7__7), .q_7__6 (filter_data_7__6), .q_7__5 (
             filter_data_7__5), .q_7__4 (filter_data_7__4), .q_7__3 (
             filter_data_7__3), .q_7__2 (filter_data_7__2), .q_7__1 (
             filter_data_7__1), .q_7__0 (filter_data_7__0), .q_8__15 (
             filter_data_8__15), .q_8__14 (filter_data_8__14), .q_8__13 (
             filter_data_8__13), .q_8__12 (filter_data_8__12), .q_8__11 (
             filter_data_8__11), .q_8__10 (filter_data_8__10), .q_8__9 (
             filter_data_8__9), .q_8__8 (filter_data_8__8), .q_8__7 (
             filter_data_8__7), .q_8__6 (filter_data_8__6), .q_8__5 (
             filter_data_8__5), .q_8__4 (filter_data_8__4), .q_8__3 (
             filter_data_8__3), .q_8__2 (filter_data_8__2), .q_8__1 (
             filter_data_8__1), .q_8__0 (filter_data_8__0), .q_9__15 (
             filter_data_9__15), .q_9__14 (filter_data_9__14), .q_9__13 (
             filter_data_9__13), .q_9__12 (filter_data_9__12), .q_9__11 (
             filter_data_9__11), .q_9__10 (filter_data_9__10), .q_9__9 (
             filter_data_9__9), .q_9__8 (filter_data_9__8), .q_9__7 (
             filter_data_9__7), .q_9__6 (filter_data_9__6), .q_9__5 (
             filter_data_9__5), .q_9__4 (filter_data_9__4), .q_9__3 (
             filter_data_9__3), .q_9__2 (filter_data_9__2), .q_9__1 (
             filter_data_9__1), .q_9__0 (filter_data_9__0), .q_10__15 (
             filter_data_10__15), .q_10__14 (filter_data_10__14), .q_10__13 (
             filter_data_10__13), .q_10__12 (filter_data_10__12), .q_10__11 (
             filter_data_10__11), .q_10__10 (filter_data_10__10), .q_10__9 (
             filter_data_10__9), .q_10__8 (filter_data_10__8), .q_10__7 (
             filter_data_10__7), .q_10__6 (filter_data_10__6), .q_10__5 (
             filter_data_10__5), .q_10__4 (filter_data_10__4), .q_10__3 (
             filter_data_10__3), .q_10__2 (filter_data_10__2), .q_10__1 (
             filter_data_10__1), .q_10__0 (filter_data_10__0), .q_11__15 (
             filter_data_11__15), .q_11__14 (filter_data_11__14), .q_11__13 (
             filter_data_11__13), .q_11__12 (filter_data_11__12), .q_11__11 (
             filter_data_11__11), .q_11__10 (filter_data_11__10), .q_11__9 (
             filter_data_11__9), .q_11__8 (filter_data_11__8), .q_11__7 (
             filter_data_11__7), .q_11__6 (filter_data_11__6), .q_11__5 (
             filter_data_11__5), .q_11__4 (filter_data_11__4), .q_11__3 (
             filter_data_11__3), .q_11__2 (filter_data_11__2), .q_11__1 (
             filter_data_11__1), .q_11__0 (filter_data_11__0), .q_12__15 (
             filter_data_12__15), .q_12__14 (filter_data_12__14), .q_12__13 (
             filter_data_12__13), .q_12__12 (filter_data_12__12), .q_12__11 (
             filter_data_12__11), .q_12__10 (filter_data_12__10), .q_12__9 (
             filter_data_12__9), .q_12__8 (filter_data_12__8), .q_12__7 (
             filter_data_12__7), .q_12__6 (filter_data_12__6), .q_12__5 (
             filter_data_12__5), .q_12__4 (filter_data_12__4), .q_12__3 (
             filter_data_12__3), .q_12__2 (filter_data_12__2), .q_12__1 (
             filter_data_12__1), .q_12__0 (filter_data_12__0), .q_13__15 (
             filter_data_13__15), .q_13__14 (filter_data_13__14), .q_13__13 (
             filter_data_13__13), .q_13__12 (filter_data_13__12), .q_13__11 (
             filter_data_13__11), .q_13__10 (filter_data_13__10), .q_13__9 (
             filter_data_13__9), .q_13__8 (filter_data_13__8), .q_13__7 (
             filter_data_13__7), .q_13__6 (filter_data_13__6), .q_13__5 (
             filter_data_13__5), .q_13__4 (filter_data_13__4), .q_13__3 (
             filter_data_13__3), .q_13__2 (filter_data_13__2), .q_13__1 (
             filter_data_13__1), .q_13__0 (filter_data_13__0), .q_14__15 (
             filter_data_14__15), .q_14__14 (filter_data_14__14), .q_14__13 (
             filter_data_14__13), .q_14__12 (filter_data_14__12), .q_14__11 (
             filter_data_14__11), .q_14__10 (filter_data_14__10), .q_14__9 (
             filter_data_14__9), .q_14__8 (filter_data_14__8), .q_14__7 (
             filter_data_14__7), .q_14__6 (filter_data_14__6), .q_14__5 (
             filter_data_14__5), .q_14__4 (filter_data_14__4), .q_14__3 (
             filter_data_14__3), .q_14__2 (filter_data_14__2), .q_14__1 (
             filter_data_14__1), .q_14__0 (filter_data_14__0), .q_15__15 (
             filter_data_15__15), .q_15__14 (filter_data_15__14), .q_15__13 (
             filter_data_15__13), .q_15__12 (filter_data_15__12), .q_15__11 (
             filter_data_15__11), .q_15__10 (filter_data_15__10), .q_15__9 (
             filter_data_15__9), .q_15__8 (filter_data_15__8), .q_15__7 (
             filter_data_15__7), .q_15__6 (filter_data_15__6), .q_15__5 (
             filter_data_15__5), .q_15__4 (filter_data_15__4), .q_15__3 (
             filter_data_15__3), .q_15__2 (filter_data_15__2), .q_15__1 (
             filter_data_15__1), .q_15__0 (filter_data_15__0), .q_16__15 (
             filter_data_16__15), .q_16__14 (filter_data_16__14), .q_16__13 (
             filter_data_16__13), .q_16__12 (filter_data_16__12), .q_16__11 (
             filter_data_16__11), .q_16__10 (filter_data_16__10), .q_16__9 (
             filter_data_16__9), .q_16__8 (filter_data_16__8), .q_16__7 (
             filter_data_16__7), .q_16__6 (filter_data_16__6), .q_16__5 (
             filter_data_16__5), .q_16__4 (filter_data_16__4), .q_16__3 (
             filter_data_16__3), .q_16__2 (filter_data_16__2), .q_16__1 (
             filter_data_16__1), .q_16__0 (filter_data_16__0), .q_17__15 (
             filter_data_17__15), .q_17__14 (filter_data_17__14), .q_17__13 (
             filter_data_17__13), .q_17__12 (filter_data_17__12), .q_17__11 (
             filter_data_17__11), .q_17__10 (filter_data_17__10), .q_17__9 (
             filter_data_17__9), .q_17__8 (filter_data_17__8), .q_17__7 (
             filter_data_17__7), .q_17__6 (filter_data_17__6), .q_17__5 (
             filter_data_17__5), .q_17__4 (filter_data_17__4), .q_17__3 (
             filter_data_17__3), .q_17__2 (filter_data_17__2), .q_17__1 (
             filter_data_17__1), .q_17__0 (filter_data_17__0), .q_18__15 (
             filter_data_18__15), .q_18__14 (filter_data_18__14), .q_18__13 (
             filter_data_18__13), .q_18__12 (filter_data_18__12), .q_18__11 (
             filter_data_18__11), .q_18__10 (filter_data_18__10), .q_18__9 (
             filter_data_18__9), .q_18__8 (filter_data_18__8), .q_18__7 (
             filter_data_18__7), .q_18__6 (filter_data_18__6), .q_18__5 (
             filter_data_18__5), .q_18__4 (filter_data_18__4), .q_18__3 (
             filter_data_18__3), .q_18__2 (filter_data_18__2), .q_18__1 (
             filter_data_18__1), .q_18__0 (filter_data_18__0), .q_19__15 (
             filter_data_19__15), .q_19__14 (filter_data_19__14), .q_19__13 (
             filter_data_19__13), .q_19__12 (filter_data_19__12), .q_19__11 (
             filter_data_19__11), .q_19__10 (filter_data_19__10), .q_19__9 (
             filter_data_19__9), .q_19__8 (filter_data_19__8), .q_19__7 (
             filter_data_19__7), .q_19__6 (filter_data_19__6), .q_19__5 (
             filter_data_19__5), .q_19__4 (filter_data_19__4), .q_19__3 (
             filter_data_19__3), .q_19__2 (filter_data_19__2), .q_19__1 (
             filter_data_19__1), .q_19__0 (filter_data_19__0), .q_20__15 (
             filter_data_20__15), .q_20__14 (filter_data_20__14), .q_20__13 (
             filter_data_20__13), .q_20__12 (filter_data_20__12), .q_20__11 (
             filter_data_20__11), .q_20__10 (filter_data_20__10), .q_20__9 (
             filter_data_20__9), .q_20__8 (filter_data_20__8), .q_20__7 (
             filter_data_20__7), .q_20__6 (filter_data_20__6), .q_20__5 (
             filter_data_20__5), .q_20__4 (filter_data_20__4), .q_20__3 (
             filter_data_20__3), .q_20__2 (filter_data_20__2), .q_20__1 (
             filter_data_20__1), .q_20__0 (filter_data_20__0), .q_21__15 (
             filter_data_21__15), .q_21__14 (filter_data_21__14), .q_21__13 (
             filter_data_21__13), .q_21__12 (filter_data_21__12), .q_21__11 (
             filter_data_21__11), .q_21__10 (filter_data_21__10), .q_21__9 (
             filter_data_21__9), .q_21__8 (filter_data_21__8), .q_21__7 (
             filter_data_21__7), .q_21__6 (filter_data_21__6), .q_21__5 (
             filter_data_21__5), .q_21__4 (filter_data_21__4), .q_21__3 (
             filter_data_21__3), .q_21__2 (filter_data_21__2), .q_21__1 (
             filter_data_21__1), .q_21__0 (filter_data_21__0), .q_22__15 (
             filter_data_22__15), .q_22__14 (filter_data_22__14), .q_22__13 (
             filter_data_22__13), .q_22__12 (filter_data_22__12), .q_22__11 (
             filter_data_22__11), .q_22__10 (filter_data_22__10), .q_22__9 (
             filter_data_22__9), .q_22__8 (filter_data_22__8), .q_22__7 (
             filter_data_22__7), .q_22__6 (filter_data_22__6), .q_22__5 (
             filter_data_22__5), .q_22__4 (filter_data_22__4), .q_22__3 (
             filter_data_22__3), .q_22__2 (filter_data_22__2), .q_22__1 (
             filter_data_22__1), .q_22__0 (filter_data_22__0), .q_23__15 (
             filter_data_23__15), .q_23__14 (filter_data_23__14), .q_23__13 (
             filter_data_23__13), .q_23__12 (filter_data_23__12), .q_23__11 (
             filter_data_23__11), .q_23__10 (filter_data_23__10), .q_23__9 (
             filter_data_23__9), .q_23__8 (filter_data_23__8), .q_23__7 (
             filter_data_23__7), .q_23__6 (filter_data_23__6), .q_23__5 (
             filter_data_23__5), .q_23__4 (filter_data_23__4), .q_23__3 (
             filter_data_23__3), .q_23__2 (filter_data_23__2), .q_23__1 (
             filter_data_23__1), .q_23__0 (filter_data_23__0), .q_24__15 (
             filter_data_24__15), .q_24__14 (filter_data_24__14), .q_24__13 (
             filter_data_24__13), .q_24__12 (filter_data_24__12), .q_24__11 (
             filter_data_24__11), .q_24__10 (filter_data_24__10), .q_24__9 (
             filter_data_24__9), .q_24__8 (filter_data_24__8), .q_24__7 (
             filter_data_24__7), .q_24__6 (filter_data_24__6), .q_24__5 (
             filter_data_24__5), .q_24__4 (filter_data_24__4), .q_24__3 (
             filter_data_24__3), .q_24__2 (filter_data_24__2), .q_24__1 (
             filter_data_24__1), .q_24__0 (filter_data_24__0), .clk (nx1181), .load (
             filter_load_tmp), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_0_gen_regi (.d ({d_cache_arr_0__31,
           d_cache_arr_0__30,d_cache_arr_0__29,d_cache_arr_0__28,
           d_cache_arr_0__27,d_cache_arr_0__26,d_cache_arr_0__25,
           d_cache_arr_0__24,d_cache_arr_0__23,d_cache_arr_0__22,
           d_cache_arr_0__21,d_cache_arr_0__20,d_cache_arr_0__19,
           d_cache_arr_0__18,d_cache_arr_0__17,d_cache_arr_0__16,
           d_cache_arr_0__15,d_cache_arr_0__14,d_cache_arr_0__13,
           d_cache_arr_0__12,d_cache_arr_0__11,d_cache_arr_0__10,
           d_cache_arr_0__9,d_cache_arr_0__8,d_cache_arr_0__7,d_cache_arr_0__6,
           d_cache_arr_0__5,d_cache_arr_0__4,d_cache_arr_0__3,d_cache_arr_0__2,
           d_cache_arr_0__1,d_cache_arr_0__0}), .q ({q_cache_arr_0__31,
           q_cache_arr_0__30,q_cache_arr_0__29,q_cache_arr_0__28,
           q_cache_arr_0__27,q_cache_arr_0__26,q_cache_arr_0__25,
           q_cache_arr_0__24,q_cache_arr_0__23,q_cache_arr_0__22,
           q_cache_arr_0__21,q_cache_arr_0__20,q_cache_arr_0__19,
           q_cache_arr_0__18,q_cache_arr_0__17,q_cache_arr_0__16,
           q_cache_arr_0__15,q_cache_arr_0__14,q_cache_arr_0__13,
           q_cache_arr_0__12,q_cache_arr_0__11,q_cache_arr_0__10,
           q_cache_arr_0__9,q_cache_arr_0__8,q_cache_arr_0__7,q_cache_arr_0__6,
           q_cache_arr_0__5,q_cache_arr_0__4,q_cache_arr_0__3,q_cache_arr_0__2,
           q_cache_arr_0__1,q_cache_arr_0__0}), .rst_data ({buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready}), .clk (clk), .load (nx1109), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_1_gen_regi (.d ({d_cache_arr_1__31,
           d_cache_arr_1__30,d_cache_arr_1__29,d_cache_arr_1__28,
           d_cache_arr_1__27,d_cache_arr_1__26,d_cache_arr_1__25,
           d_cache_arr_1__24,d_cache_arr_1__23,d_cache_arr_1__22,
           d_cache_arr_1__21,d_cache_arr_1__20,d_cache_arr_1__19,
           d_cache_arr_1__18,d_cache_arr_1__17,d_cache_arr_1__16,
           d_cache_arr_1__15,d_cache_arr_1__14,d_cache_arr_1__13,
           d_cache_arr_1__12,d_cache_arr_1__11,d_cache_arr_1__10,
           d_cache_arr_1__9,d_cache_arr_1__8,d_cache_arr_1__7,d_cache_arr_1__6,
           d_cache_arr_1__5,d_cache_arr_1__4,d_cache_arr_1__3,d_cache_arr_1__2,
           d_cache_arr_1__1,d_cache_arr_1__0}), .q ({q_cache_arr_1__31,
           q_cache_arr_1__30,q_cache_arr_1__29,q_cache_arr_1__28,
           q_cache_arr_1__27,q_cache_arr_1__26,q_cache_arr_1__25,
           q_cache_arr_1__24,q_cache_arr_1__23,q_cache_arr_1__22,
           q_cache_arr_1__21,q_cache_arr_1__20,q_cache_arr_1__19,
           q_cache_arr_1__18,q_cache_arr_1__17,q_cache_arr_1__16,
           q_cache_arr_1__15,q_cache_arr_1__14,q_cache_arr_1__13,
           q_cache_arr_1__12,q_cache_arr_1__11,q_cache_arr_1__10,
           q_cache_arr_1__9,q_cache_arr_1__8,q_cache_arr_1__7,q_cache_arr_1__6,
           q_cache_arr_1__5,q_cache_arr_1__4,q_cache_arr_1__3,q_cache_arr_1__2,
           q_cache_arr_1__1,q_cache_arr_1__0}), .rst_data ({buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready}), .clk (clk), .load (nx1109), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_2_gen_regi (.d ({d_cache_arr_2__31,
           d_cache_arr_2__30,d_cache_arr_2__29,d_cache_arr_2__28,
           d_cache_arr_2__27,d_cache_arr_2__26,d_cache_arr_2__25,
           d_cache_arr_2__24,d_cache_arr_2__23,d_cache_arr_2__22,
           d_cache_arr_2__21,d_cache_arr_2__20,d_cache_arr_2__19,
           d_cache_arr_2__18,d_cache_arr_2__17,d_cache_arr_2__16,
           d_cache_arr_2__15,d_cache_arr_2__14,d_cache_arr_2__13,
           d_cache_arr_2__12,d_cache_arr_2__11,d_cache_arr_2__10,
           d_cache_arr_2__9,d_cache_arr_2__8,d_cache_arr_2__7,d_cache_arr_2__6,
           d_cache_arr_2__5,d_cache_arr_2__4,d_cache_arr_2__3,d_cache_arr_2__2,
           d_cache_arr_2__1,d_cache_arr_2__0}), .q ({q_cache_arr_2__31,
           q_cache_arr_2__30,q_cache_arr_2__29,q_cache_arr_2__28,
           q_cache_arr_2__27,q_cache_arr_2__26,q_cache_arr_2__25,
           q_cache_arr_2__24,q_cache_arr_2__23,q_cache_arr_2__22,
           q_cache_arr_2__21,q_cache_arr_2__20,q_cache_arr_2__19,
           q_cache_arr_2__18,q_cache_arr_2__17,q_cache_arr_2__16,
           q_cache_arr_2__15,q_cache_arr_2__14,q_cache_arr_2__13,
           q_cache_arr_2__12,q_cache_arr_2__11,q_cache_arr_2__10,
           q_cache_arr_2__9,q_cache_arr_2__8,q_cache_arr_2__7,q_cache_arr_2__6,
           q_cache_arr_2__5,q_cache_arr_2__4,q_cache_arr_2__3,q_cache_arr_2__2,
           q_cache_arr_2__1,q_cache_arr_2__0}), .rst_data ({buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready}), .clk (clk), .load (nx1109), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_3_gen_regi (.d ({d_cache_arr_3__31,
           d_cache_arr_3__30,d_cache_arr_3__29,d_cache_arr_3__28,
           d_cache_arr_3__27,d_cache_arr_3__26,d_cache_arr_3__25,
           d_cache_arr_3__24,d_cache_arr_3__23,d_cache_arr_3__22,
           d_cache_arr_3__21,d_cache_arr_3__20,d_cache_arr_3__19,
           d_cache_arr_3__18,d_cache_arr_3__17,d_cache_arr_3__16,
           d_cache_arr_3__15,d_cache_arr_3__14,d_cache_arr_3__13,
           d_cache_arr_3__12,d_cache_arr_3__11,d_cache_arr_3__10,
           d_cache_arr_3__9,d_cache_arr_3__8,d_cache_arr_3__7,d_cache_arr_3__6,
           d_cache_arr_3__5,d_cache_arr_3__4,d_cache_arr_3__3,d_cache_arr_3__2,
           d_cache_arr_3__1,d_cache_arr_3__0}), .q ({q_cache_arr_3__31,
           q_cache_arr_3__30,q_cache_arr_3__29,q_cache_arr_3__28,
           q_cache_arr_3__27,q_cache_arr_3__26,q_cache_arr_3__25,
           q_cache_arr_3__24,q_cache_arr_3__23,q_cache_arr_3__22,
           q_cache_arr_3__21,q_cache_arr_3__20,q_cache_arr_3__19,
           q_cache_arr_3__18,q_cache_arr_3__17,q_cache_arr_3__16,
           q_cache_arr_3__15,q_cache_arr_3__14,q_cache_arr_3__13,
           q_cache_arr_3__12,q_cache_arr_3__11,q_cache_arr_3__10,
           q_cache_arr_3__9,q_cache_arr_3__8,q_cache_arr_3__7,q_cache_arr_3__6,
           q_cache_arr_3__5,q_cache_arr_3__4,q_cache_arr_3__3,q_cache_arr_3__2,
           q_cache_arr_3__1,q_cache_arr_3__0}), .rst_data ({buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready}), .clk (clk), .load (nx1109), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_4_gen_regi (.d ({d_cache_arr_4__31,
           d_cache_arr_4__30,d_cache_arr_4__29,d_cache_arr_4__28,
           d_cache_arr_4__27,d_cache_arr_4__26,d_cache_arr_4__25,
           d_cache_arr_4__24,d_cache_arr_4__23,d_cache_arr_4__22,
           d_cache_arr_4__21,d_cache_arr_4__20,d_cache_arr_4__19,
           d_cache_arr_4__18,d_cache_arr_4__17,d_cache_arr_4__16,
           d_cache_arr_4__15,d_cache_arr_4__14,d_cache_arr_4__13,
           d_cache_arr_4__12,d_cache_arr_4__11,d_cache_arr_4__10,
           d_cache_arr_4__9,d_cache_arr_4__8,d_cache_arr_4__7,d_cache_arr_4__6,
           d_cache_arr_4__5,d_cache_arr_4__4,d_cache_arr_4__3,d_cache_arr_4__2,
           d_cache_arr_4__1,d_cache_arr_4__0}), .q ({q_cache_arr_4__31,
           q_cache_arr_4__30,q_cache_arr_4__29,q_cache_arr_4__28,
           q_cache_arr_4__27,q_cache_arr_4__26,q_cache_arr_4__25,
           q_cache_arr_4__24,q_cache_arr_4__23,q_cache_arr_4__22,
           q_cache_arr_4__21,q_cache_arr_4__20,q_cache_arr_4__19,
           q_cache_arr_4__18,q_cache_arr_4__17,q_cache_arr_4__16,
           q_cache_arr_4__15,q_cache_arr_4__14,q_cache_arr_4__13,
           q_cache_arr_4__12,q_cache_arr_4__11,q_cache_arr_4__10,
           q_cache_arr_4__9,q_cache_arr_4__8,q_cache_arr_4__7,q_cache_arr_4__6,
           q_cache_arr_4__5,q_cache_arr_4__4,q_cache_arr_4__3,q_cache_arr_4__2,
           q_cache_arr_4__1,q_cache_arr_4__0}), .rst_data ({buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready}), .clk (clk), .load (nx1109), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_5_gen_regi (.d ({d_cache_arr_5__31,
           d_cache_arr_5__30,d_cache_arr_5__29,d_cache_arr_5__28,
           d_cache_arr_5__27,d_cache_arr_5__26,d_cache_arr_5__25,
           d_cache_arr_5__24,d_cache_arr_5__23,d_cache_arr_5__22,
           d_cache_arr_5__21,d_cache_arr_5__20,d_cache_arr_5__19,
           d_cache_arr_5__18,d_cache_arr_5__17,d_cache_arr_5__16,
           d_cache_arr_5__15,d_cache_arr_5__14,d_cache_arr_5__13,
           d_cache_arr_5__12,d_cache_arr_5__11,d_cache_arr_5__10,
           d_cache_arr_5__9,d_cache_arr_5__8,d_cache_arr_5__7,d_cache_arr_5__6,
           d_cache_arr_5__5,d_cache_arr_5__4,d_cache_arr_5__3,d_cache_arr_5__2,
           d_cache_arr_5__1,d_cache_arr_5__0}), .q ({q_cache_arr_5__31,
           q_cache_arr_5__30,q_cache_arr_5__29,q_cache_arr_5__28,
           q_cache_arr_5__27,q_cache_arr_5__26,q_cache_arr_5__25,
           q_cache_arr_5__24,q_cache_arr_5__23,q_cache_arr_5__22,
           q_cache_arr_5__21,q_cache_arr_5__20,q_cache_arr_5__19,
           q_cache_arr_5__18,q_cache_arr_5__17,q_cache_arr_5__16,
           q_cache_arr_5__15,q_cache_arr_5__14,q_cache_arr_5__13,
           q_cache_arr_5__12,q_cache_arr_5__11,q_cache_arr_5__10,
           q_cache_arr_5__9,q_cache_arr_5__8,q_cache_arr_5__7,q_cache_arr_5__6,
           q_cache_arr_5__5,q_cache_arr_5__4,q_cache_arr_5__3,q_cache_arr_5__2,
           q_cache_arr_5__1,q_cache_arr_5__0}), .rst_data ({buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready}), .clk (clk), .load (nx1109), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_6_gen_regi (.d ({d_cache_arr_6__31,
           d_cache_arr_6__30,d_cache_arr_6__29,d_cache_arr_6__28,
           d_cache_arr_6__27,d_cache_arr_6__26,d_cache_arr_6__25,
           d_cache_arr_6__24,d_cache_arr_6__23,d_cache_arr_6__22,
           d_cache_arr_6__21,d_cache_arr_6__20,d_cache_arr_6__19,
           d_cache_arr_6__18,d_cache_arr_6__17,d_cache_arr_6__16,
           d_cache_arr_6__15,d_cache_arr_6__14,d_cache_arr_6__13,
           d_cache_arr_6__12,d_cache_arr_6__11,d_cache_arr_6__10,
           d_cache_arr_6__9,d_cache_arr_6__8,d_cache_arr_6__7,d_cache_arr_6__6,
           d_cache_arr_6__5,d_cache_arr_6__4,d_cache_arr_6__3,d_cache_arr_6__2,
           d_cache_arr_6__1,d_cache_arr_6__0}), .q ({q_cache_arr_6__31,
           q_cache_arr_6__30,q_cache_arr_6__29,q_cache_arr_6__28,
           q_cache_arr_6__27,q_cache_arr_6__26,q_cache_arr_6__25,
           q_cache_arr_6__24,q_cache_arr_6__23,q_cache_arr_6__22,
           q_cache_arr_6__21,q_cache_arr_6__20,q_cache_arr_6__19,
           q_cache_arr_6__18,q_cache_arr_6__17,q_cache_arr_6__16,
           q_cache_arr_6__15,q_cache_arr_6__14,q_cache_arr_6__13,
           q_cache_arr_6__12,q_cache_arr_6__11,q_cache_arr_6__10,
           q_cache_arr_6__9,q_cache_arr_6__8,q_cache_arr_6__7,q_cache_arr_6__6,
           q_cache_arr_6__5,q_cache_arr_6__4,q_cache_arr_6__3,q_cache_arr_6__2,
           q_cache_arr_6__1,q_cache_arr_6__0}), .rst_data ({buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready}), .clk (clk), .load (nx1109), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_7_gen_regi (.d ({d_cache_arr_7__31,
           d_cache_arr_7__30,d_cache_arr_7__29,d_cache_arr_7__28,
           d_cache_arr_7__27,d_cache_arr_7__26,d_cache_arr_7__25,
           d_cache_arr_7__24,d_cache_arr_7__23,d_cache_arr_7__22,
           d_cache_arr_7__21,d_cache_arr_7__20,d_cache_arr_7__19,
           d_cache_arr_7__18,d_cache_arr_7__17,d_cache_arr_7__16,
           d_cache_arr_7__15,d_cache_arr_7__14,d_cache_arr_7__13,
           d_cache_arr_7__12,d_cache_arr_7__11,d_cache_arr_7__10,
           d_cache_arr_7__9,d_cache_arr_7__8,d_cache_arr_7__7,d_cache_arr_7__6,
           d_cache_arr_7__5,d_cache_arr_7__4,d_cache_arr_7__3,d_cache_arr_7__2,
           d_cache_arr_7__1,d_cache_arr_7__0}), .q ({q_cache_arr_7__31,
           q_cache_arr_7__30,q_cache_arr_7__29,q_cache_arr_7__28,
           q_cache_arr_7__27,q_cache_arr_7__26,q_cache_arr_7__25,
           q_cache_arr_7__24,q_cache_arr_7__23,q_cache_arr_7__22,
           q_cache_arr_7__21,q_cache_arr_7__20,q_cache_arr_7__19,
           q_cache_arr_7__18,q_cache_arr_7__17,q_cache_arr_7__16,
           q_cache_arr_7__15,q_cache_arr_7__14,q_cache_arr_7__13,
           q_cache_arr_7__12,q_cache_arr_7__11,q_cache_arr_7__10,
           q_cache_arr_7__9,q_cache_arr_7__8,q_cache_arr_7__7,q_cache_arr_7__6,
           q_cache_arr_7__5,q_cache_arr_7__4,q_cache_arr_7__3,q_cache_arr_7__2,
           q_cache_arr_7__1,q_cache_arr_7__0}), .rst_data ({buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready}), .clk (clk), .load (nx1111), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_8_gen_regi (.d ({d_cache_arr_8__31,
           d_cache_arr_8__30,d_cache_arr_8__29,d_cache_arr_8__28,
           d_cache_arr_8__27,d_cache_arr_8__26,d_cache_arr_8__25,
           d_cache_arr_8__24,d_cache_arr_8__23,d_cache_arr_8__22,
           d_cache_arr_8__21,d_cache_arr_8__20,d_cache_arr_8__19,
           d_cache_arr_8__18,d_cache_arr_8__17,d_cache_arr_8__16,
           d_cache_arr_8__15,d_cache_arr_8__14,d_cache_arr_8__13,
           d_cache_arr_8__12,d_cache_arr_8__11,d_cache_arr_8__10,
           d_cache_arr_8__9,d_cache_arr_8__8,d_cache_arr_8__7,d_cache_arr_8__6,
           d_cache_arr_8__5,d_cache_arr_8__4,d_cache_arr_8__3,d_cache_arr_8__2,
           d_cache_arr_8__1,d_cache_arr_8__0}), .q ({q_cache_arr_8__31,
           q_cache_arr_8__30,q_cache_arr_8__29,q_cache_arr_8__28,
           q_cache_arr_8__27,q_cache_arr_8__26,q_cache_arr_8__25,
           q_cache_arr_8__24,q_cache_arr_8__23,q_cache_arr_8__22,
           q_cache_arr_8__21,q_cache_arr_8__20,q_cache_arr_8__19,
           q_cache_arr_8__18,q_cache_arr_8__17,q_cache_arr_8__16,
           q_cache_arr_8__15,q_cache_arr_8__14,q_cache_arr_8__13,
           q_cache_arr_8__12,q_cache_arr_8__11,q_cache_arr_8__10,
           q_cache_arr_8__9,q_cache_arr_8__8,q_cache_arr_8__7,q_cache_arr_8__6,
           q_cache_arr_8__5,q_cache_arr_8__4,q_cache_arr_8__3,q_cache_arr_8__2,
           q_cache_arr_8__1,q_cache_arr_8__0}), .rst_data ({buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready}), .clk (clk), .load (nx1111), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_9_gen_regi (.d ({d_cache_arr_9__31,
           d_cache_arr_9__30,d_cache_arr_9__29,d_cache_arr_9__28,
           d_cache_arr_9__27,d_cache_arr_9__26,d_cache_arr_9__25,
           d_cache_arr_9__24,d_cache_arr_9__23,d_cache_arr_9__22,
           d_cache_arr_9__21,d_cache_arr_9__20,d_cache_arr_9__19,
           d_cache_arr_9__18,d_cache_arr_9__17,d_cache_arr_9__16,
           d_cache_arr_9__15,d_cache_arr_9__14,d_cache_arr_9__13,
           d_cache_arr_9__12,d_cache_arr_9__11,d_cache_arr_9__10,
           d_cache_arr_9__9,d_cache_arr_9__8,d_cache_arr_9__7,d_cache_arr_9__6,
           d_cache_arr_9__5,d_cache_arr_9__4,d_cache_arr_9__3,d_cache_arr_9__2,
           d_cache_arr_9__1,d_cache_arr_9__0}), .q ({q_cache_arr_9__31,
           q_cache_arr_9__30,q_cache_arr_9__29,q_cache_arr_9__28,
           q_cache_arr_9__27,q_cache_arr_9__26,q_cache_arr_9__25,
           q_cache_arr_9__24,q_cache_arr_9__23,q_cache_arr_9__22,
           q_cache_arr_9__21,q_cache_arr_9__20,q_cache_arr_9__19,
           q_cache_arr_9__18,q_cache_arr_9__17,q_cache_arr_9__16,
           q_cache_arr_9__15,q_cache_arr_9__14,q_cache_arr_9__13,
           q_cache_arr_9__12,q_cache_arr_9__11,q_cache_arr_9__10,
           q_cache_arr_9__9,q_cache_arr_9__8,q_cache_arr_9__7,q_cache_arr_9__6,
           q_cache_arr_9__5,q_cache_arr_9__4,q_cache_arr_9__3,q_cache_arr_9__2,
           q_cache_arr_9__1,q_cache_arr_9__0}), .rst_data ({buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready}), .clk (clk), .load (nx1111), .reset (filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_10_gen_regi (.d ({d_cache_arr_10__31,
           d_cache_arr_10__30,d_cache_arr_10__29,d_cache_arr_10__28,
           d_cache_arr_10__27,d_cache_arr_10__26,d_cache_arr_10__25,
           d_cache_arr_10__24,d_cache_arr_10__23,d_cache_arr_10__22,
           d_cache_arr_10__21,d_cache_arr_10__20,d_cache_arr_10__19,
           d_cache_arr_10__18,d_cache_arr_10__17,d_cache_arr_10__16,
           d_cache_arr_10__15,d_cache_arr_10__14,d_cache_arr_10__13,
           d_cache_arr_10__12,d_cache_arr_10__11,d_cache_arr_10__10,
           d_cache_arr_10__9,d_cache_arr_10__8,d_cache_arr_10__7,
           d_cache_arr_10__6,d_cache_arr_10__5,d_cache_arr_10__4,
           d_cache_arr_10__3,d_cache_arr_10__2,d_cache_arr_10__1,
           d_cache_arr_10__0}), .q ({q_cache_arr_10__31,q_cache_arr_10__30,
           q_cache_arr_10__29,q_cache_arr_10__28,q_cache_arr_10__27,
           q_cache_arr_10__26,q_cache_arr_10__25,q_cache_arr_10__24,
           q_cache_arr_10__23,q_cache_arr_10__22,q_cache_arr_10__21,
           q_cache_arr_10__20,q_cache_arr_10__19,q_cache_arr_10__18,
           q_cache_arr_10__17,q_cache_arr_10__16,q_cache_arr_10__15,
           q_cache_arr_10__14,q_cache_arr_10__13,q_cache_arr_10__12,
           q_cache_arr_10__11,q_cache_arr_10__10,q_cache_arr_10__9,
           q_cache_arr_10__8,q_cache_arr_10__7,q_cache_arr_10__6,
           q_cache_arr_10__5,q_cache_arr_10__4,q_cache_arr_10__3,
           q_cache_arr_10__2,q_cache_arr_10__1,q_cache_arr_10__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1111), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_11_gen_regi (.d ({d_cache_arr_11__31,
           d_cache_arr_11__30,d_cache_arr_11__29,d_cache_arr_11__28,
           d_cache_arr_11__27,d_cache_arr_11__26,d_cache_arr_11__25,
           d_cache_arr_11__24,d_cache_arr_11__23,d_cache_arr_11__22,
           d_cache_arr_11__21,d_cache_arr_11__20,d_cache_arr_11__19,
           d_cache_arr_11__18,d_cache_arr_11__17,d_cache_arr_11__16,
           d_cache_arr_11__15,d_cache_arr_11__14,d_cache_arr_11__13,
           d_cache_arr_11__12,d_cache_arr_11__11,d_cache_arr_11__10,
           d_cache_arr_11__9,d_cache_arr_11__8,d_cache_arr_11__7,
           d_cache_arr_11__6,d_cache_arr_11__5,d_cache_arr_11__4,
           d_cache_arr_11__3,d_cache_arr_11__2,d_cache_arr_11__1,
           d_cache_arr_11__0}), .q ({q_cache_arr_11__31,q_cache_arr_11__30,
           q_cache_arr_11__29,q_cache_arr_11__28,q_cache_arr_11__27,
           q_cache_arr_11__26,q_cache_arr_11__25,q_cache_arr_11__24,
           q_cache_arr_11__23,q_cache_arr_11__22,q_cache_arr_11__21,
           q_cache_arr_11__20,q_cache_arr_11__19,q_cache_arr_11__18,
           q_cache_arr_11__17,q_cache_arr_11__16,q_cache_arr_11__15,
           q_cache_arr_11__14,q_cache_arr_11__13,q_cache_arr_11__12,
           q_cache_arr_11__11,q_cache_arr_11__10,q_cache_arr_11__9,
           q_cache_arr_11__8,q_cache_arr_11__7,q_cache_arr_11__6,
           q_cache_arr_11__5,q_cache_arr_11__4,q_cache_arr_11__3,
           q_cache_arr_11__2,q_cache_arr_11__1,q_cache_arr_11__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1111), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_12_gen_regi (.d ({d_cache_arr_12__31,
           d_cache_arr_12__30,d_cache_arr_12__29,d_cache_arr_12__28,
           d_cache_arr_12__27,d_cache_arr_12__26,d_cache_arr_12__25,
           d_cache_arr_12__24,d_cache_arr_12__23,d_cache_arr_12__22,
           d_cache_arr_12__21,d_cache_arr_12__20,d_cache_arr_12__19,
           d_cache_arr_12__18,d_cache_arr_12__17,d_cache_arr_12__16,
           d_cache_arr_12__15,d_cache_arr_12__14,d_cache_arr_12__13,
           d_cache_arr_12__12,d_cache_arr_12__11,d_cache_arr_12__10,
           d_cache_arr_12__9,d_cache_arr_12__8,d_cache_arr_12__7,
           d_cache_arr_12__6,d_cache_arr_12__5,d_cache_arr_12__4,
           d_cache_arr_12__3,d_cache_arr_12__2,d_cache_arr_12__1,
           d_cache_arr_12__0}), .q ({q_cache_arr_12__31,q_cache_arr_12__30,
           q_cache_arr_12__29,q_cache_arr_12__28,q_cache_arr_12__27,
           q_cache_arr_12__26,q_cache_arr_12__25,q_cache_arr_12__24,
           q_cache_arr_12__23,q_cache_arr_12__22,q_cache_arr_12__21,
           q_cache_arr_12__20,q_cache_arr_12__19,q_cache_arr_12__18,
           q_cache_arr_12__17,q_cache_arr_12__16,q_cache_arr_12__15,
           q_cache_arr_12__14,q_cache_arr_12__13,q_cache_arr_12__12,
           q_cache_arr_12__11,q_cache_arr_12__10,q_cache_arr_12__9,
           q_cache_arr_12__8,q_cache_arr_12__7,q_cache_arr_12__6,
           q_cache_arr_12__5,q_cache_arr_12__4,q_cache_arr_12__3,
           q_cache_arr_12__2,q_cache_arr_12__1,q_cache_arr_12__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1111), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_13_gen_regi (.d ({d_cache_arr_13__31,
           d_cache_arr_13__30,d_cache_arr_13__29,d_cache_arr_13__28,
           d_cache_arr_13__27,d_cache_arr_13__26,d_cache_arr_13__25,
           d_cache_arr_13__24,d_cache_arr_13__23,d_cache_arr_13__22,
           d_cache_arr_13__21,d_cache_arr_13__20,d_cache_arr_13__19,
           d_cache_arr_13__18,d_cache_arr_13__17,d_cache_arr_13__16,
           d_cache_arr_13__15,d_cache_arr_13__14,d_cache_arr_13__13,
           d_cache_arr_13__12,d_cache_arr_13__11,d_cache_arr_13__10,
           d_cache_arr_13__9,d_cache_arr_13__8,d_cache_arr_13__7,
           d_cache_arr_13__6,d_cache_arr_13__5,d_cache_arr_13__4,
           d_cache_arr_13__3,d_cache_arr_13__2,d_cache_arr_13__1,
           d_cache_arr_13__0}), .q ({q_cache_arr_13__31,q_cache_arr_13__30,
           q_cache_arr_13__29,q_cache_arr_13__28,q_cache_arr_13__27,
           q_cache_arr_13__26,q_cache_arr_13__25,q_cache_arr_13__24,
           q_cache_arr_13__23,q_cache_arr_13__22,q_cache_arr_13__21,
           q_cache_arr_13__20,q_cache_arr_13__19,q_cache_arr_13__18,
           q_cache_arr_13__17,q_cache_arr_13__16,q_cache_arr_13__15,
           q_cache_arr_13__14,q_cache_arr_13__13,q_cache_arr_13__12,
           q_cache_arr_13__11,q_cache_arr_13__10,q_cache_arr_13__9,
           q_cache_arr_13__8,q_cache_arr_13__7,q_cache_arr_13__6,
           q_cache_arr_13__5,q_cache_arr_13__4,q_cache_arr_13__3,
           q_cache_arr_13__2,q_cache_arr_13__1,q_cache_arr_13__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1111), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_14_gen_regi (.d ({d_cache_arr_14__31,
           d_cache_arr_14__30,d_cache_arr_14__29,d_cache_arr_14__28,
           d_cache_arr_14__27,d_cache_arr_14__26,d_cache_arr_14__25,
           d_cache_arr_14__24,d_cache_arr_14__23,d_cache_arr_14__22,
           d_cache_arr_14__21,d_cache_arr_14__20,d_cache_arr_14__19,
           d_cache_arr_14__18,d_cache_arr_14__17,d_cache_arr_14__16,
           d_cache_arr_14__15,d_cache_arr_14__14,d_cache_arr_14__13,
           d_cache_arr_14__12,d_cache_arr_14__11,d_cache_arr_14__10,
           d_cache_arr_14__9,d_cache_arr_14__8,d_cache_arr_14__7,
           d_cache_arr_14__6,d_cache_arr_14__5,d_cache_arr_14__4,
           d_cache_arr_14__3,d_cache_arr_14__2,d_cache_arr_14__1,
           d_cache_arr_14__0}), .q ({q_cache_arr_14__31,q_cache_arr_14__30,
           q_cache_arr_14__29,q_cache_arr_14__28,q_cache_arr_14__27,
           q_cache_arr_14__26,q_cache_arr_14__25,q_cache_arr_14__24,
           q_cache_arr_14__23,q_cache_arr_14__22,q_cache_arr_14__21,
           q_cache_arr_14__20,q_cache_arr_14__19,q_cache_arr_14__18,
           q_cache_arr_14__17,q_cache_arr_14__16,q_cache_arr_14__15,
           q_cache_arr_14__14,q_cache_arr_14__13,q_cache_arr_14__12,
           q_cache_arr_14__11,q_cache_arr_14__10,q_cache_arr_14__9,
           q_cache_arr_14__8,q_cache_arr_14__7,q_cache_arr_14__6,
           q_cache_arr_14__5,q_cache_arr_14__4,q_cache_arr_14__3,
           q_cache_arr_14__2,q_cache_arr_14__1,q_cache_arr_14__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1113), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_15_gen_regi (.d ({d_cache_arr_15__31,
           d_cache_arr_15__30,d_cache_arr_15__29,d_cache_arr_15__28,
           d_cache_arr_15__27,d_cache_arr_15__26,d_cache_arr_15__25,
           d_cache_arr_15__24,d_cache_arr_15__23,d_cache_arr_15__22,
           d_cache_arr_15__21,d_cache_arr_15__20,d_cache_arr_15__19,
           d_cache_arr_15__18,d_cache_arr_15__17,d_cache_arr_15__16,
           d_cache_arr_15__15,d_cache_arr_15__14,d_cache_arr_15__13,
           d_cache_arr_15__12,d_cache_arr_15__11,d_cache_arr_15__10,
           d_cache_arr_15__9,d_cache_arr_15__8,d_cache_arr_15__7,
           d_cache_arr_15__6,d_cache_arr_15__5,d_cache_arr_15__4,
           d_cache_arr_15__3,d_cache_arr_15__2,d_cache_arr_15__1,
           d_cache_arr_15__0}), .q ({q_cache_arr_15__31,q_cache_arr_15__30,
           q_cache_arr_15__29,q_cache_arr_15__28,q_cache_arr_15__27,
           q_cache_arr_15__26,q_cache_arr_15__25,q_cache_arr_15__24,
           q_cache_arr_15__23,q_cache_arr_15__22,q_cache_arr_15__21,
           q_cache_arr_15__20,q_cache_arr_15__19,q_cache_arr_15__18,
           q_cache_arr_15__17,q_cache_arr_15__16,q_cache_arr_15__15,
           q_cache_arr_15__14,q_cache_arr_15__13,q_cache_arr_15__12,
           q_cache_arr_15__11,q_cache_arr_15__10,q_cache_arr_15__9,
           q_cache_arr_15__8,q_cache_arr_15__7,q_cache_arr_15__6,
           q_cache_arr_15__5,q_cache_arr_15__4,q_cache_arr_15__3,
           q_cache_arr_15__2,q_cache_arr_15__1,q_cache_arr_15__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1113), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_16_gen_regi (.d ({d_cache_arr_16__31,
           d_cache_arr_16__30,d_cache_arr_16__29,d_cache_arr_16__28,
           d_cache_arr_16__27,d_cache_arr_16__26,d_cache_arr_16__25,
           d_cache_arr_16__24,d_cache_arr_16__23,d_cache_arr_16__22,
           d_cache_arr_16__21,d_cache_arr_16__20,d_cache_arr_16__19,
           d_cache_arr_16__18,d_cache_arr_16__17,d_cache_arr_16__16,
           d_cache_arr_16__15,d_cache_arr_16__14,d_cache_arr_16__13,
           d_cache_arr_16__12,d_cache_arr_16__11,d_cache_arr_16__10,
           d_cache_arr_16__9,d_cache_arr_16__8,d_cache_arr_16__7,
           d_cache_arr_16__6,d_cache_arr_16__5,d_cache_arr_16__4,
           d_cache_arr_16__3,d_cache_arr_16__2,d_cache_arr_16__1,
           d_cache_arr_16__0}), .q ({q_cache_arr_16__31,q_cache_arr_16__30,
           q_cache_arr_16__29,q_cache_arr_16__28,q_cache_arr_16__27,
           q_cache_arr_16__26,q_cache_arr_16__25,q_cache_arr_16__24,
           q_cache_arr_16__23,q_cache_arr_16__22,q_cache_arr_16__21,
           q_cache_arr_16__20,q_cache_arr_16__19,q_cache_arr_16__18,
           q_cache_arr_16__17,q_cache_arr_16__16,q_cache_arr_16__15,
           q_cache_arr_16__14,q_cache_arr_16__13,q_cache_arr_16__12,
           q_cache_arr_16__11,q_cache_arr_16__10,q_cache_arr_16__9,
           q_cache_arr_16__8,q_cache_arr_16__7,q_cache_arr_16__6,
           q_cache_arr_16__5,q_cache_arr_16__4,q_cache_arr_16__3,
           q_cache_arr_16__2,q_cache_arr_16__1,q_cache_arr_16__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1113), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_17_gen_regi (.d ({d_cache_arr_17__31,
           d_cache_arr_17__30,d_cache_arr_17__29,d_cache_arr_17__28,
           d_cache_arr_17__27,d_cache_arr_17__26,d_cache_arr_17__25,
           d_cache_arr_17__24,d_cache_arr_17__23,d_cache_arr_17__22,
           d_cache_arr_17__21,d_cache_arr_17__20,d_cache_arr_17__19,
           d_cache_arr_17__18,d_cache_arr_17__17,d_cache_arr_17__16,
           d_cache_arr_17__15,d_cache_arr_17__14,d_cache_arr_17__13,
           d_cache_arr_17__12,d_cache_arr_17__11,d_cache_arr_17__10,
           d_cache_arr_17__9,d_cache_arr_17__8,d_cache_arr_17__7,
           d_cache_arr_17__6,d_cache_arr_17__5,d_cache_arr_17__4,
           d_cache_arr_17__3,d_cache_arr_17__2,d_cache_arr_17__1,
           d_cache_arr_17__0}), .q ({q_cache_arr_17__31,q_cache_arr_17__30,
           q_cache_arr_17__29,q_cache_arr_17__28,q_cache_arr_17__27,
           q_cache_arr_17__26,q_cache_arr_17__25,q_cache_arr_17__24,
           q_cache_arr_17__23,q_cache_arr_17__22,q_cache_arr_17__21,
           q_cache_arr_17__20,q_cache_arr_17__19,q_cache_arr_17__18,
           q_cache_arr_17__17,q_cache_arr_17__16,q_cache_arr_17__15,
           q_cache_arr_17__14,q_cache_arr_17__13,q_cache_arr_17__12,
           q_cache_arr_17__11,q_cache_arr_17__10,q_cache_arr_17__9,
           q_cache_arr_17__8,q_cache_arr_17__7,q_cache_arr_17__6,
           q_cache_arr_17__5,q_cache_arr_17__4,q_cache_arr_17__3,
           q_cache_arr_17__2,q_cache_arr_17__1,q_cache_arr_17__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1113), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_18_gen_regi (.d ({d_cache_arr_18__31,
           d_cache_arr_18__30,d_cache_arr_18__29,d_cache_arr_18__28,
           d_cache_arr_18__27,d_cache_arr_18__26,d_cache_arr_18__25,
           d_cache_arr_18__24,d_cache_arr_18__23,d_cache_arr_18__22,
           d_cache_arr_18__21,d_cache_arr_18__20,d_cache_arr_18__19,
           d_cache_arr_18__18,d_cache_arr_18__17,d_cache_arr_18__16,
           d_cache_arr_18__15,d_cache_arr_18__14,d_cache_arr_18__13,
           d_cache_arr_18__12,d_cache_arr_18__11,d_cache_arr_18__10,
           d_cache_arr_18__9,d_cache_arr_18__8,d_cache_arr_18__7,
           d_cache_arr_18__6,d_cache_arr_18__5,d_cache_arr_18__4,
           d_cache_arr_18__3,d_cache_arr_18__2,d_cache_arr_18__1,
           d_cache_arr_18__0}), .q ({q_cache_arr_18__31,q_cache_arr_18__30,
           q_cache_arr_18__29,q_cache_arr_18__28,q_cache_arr_18__27,
           q_cache_arr_18__26,q_cache_arr_18__25,q_cache_arr_18__24,
           q_cache_arr_18__23,q_cache_arr_18__22,q_cache_arr_18__21,
           q_cache_arr_18__20,q_cache_arr_18__19,q_cache_arr_18__18,
           q_cache_arr_18__17,q_cache_arr_18__16,q_cache_arr_18__15,
           q_cache_arr_18__14,q_cache_arr_18__13,q_cache_arr_18__12,
           q_cache_arr_18__11,q_cache_arr_18__10,q_cache_arr_18__9,
           q_cache_arr_18__8,q_cache_arr_18__7,q_cache_arr_18__6,
           q_cache_arr_18__5,q_cache_arr_18__4,q_cache_arr_18__3,
           q_cache_arr_18__2,q_cache_arr_18__1,q_cache_arr_18__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1113), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_19_gen_regi (.d ({d_cache_arr_19__31,
           d_cache_arr_19__30,d_cache_arr_19__29,d_cache_arr_19__28,
           d_cache_arr_19__27,d_cache_arr_19__26,d_cache_arr_19__25,
           d_cache_arr_19__24,d_cache_arr_19__23,d_cache_arr_19__22,
           d_cache_arr_19__21,d_cache_arr_19__20,d_cache_arr_19__19,
           d_cache_arr_19__18,d_cache_arr_19__17,d_cache_arr_19__16,
           d_cache_arr_19__15,d_cache_arr_19__14,d_cache_arr_19__13,
           d_cache_arr_19__12,d_cache_arr_19__11,d_cache_arr_19__10,
           d_cache_arr_19__9,d_cache_arr_19__8,d_cache_arr_19__7,
           d_cache_arr_19__6,d_cache_arr_19__5,d_cache_arr_19__4,
           d_cache_arr_19__3,d_cache_arr_19__2,d_cache_arr_19__1,
           d_cache_arr_19__0}), .q ({q_cache_arr_19__31,q_cache_arr_19__30,
           q_cache_arr_19__29,q_cache_arr_19__28,q_cache_arr_19__27,
           q_cache_arr_19__26,q_cache_arr_19__25,q_cache_arr_19__24,
           q_cache_arr_19__23,q_cache_arr_19__22,q_cache_arr_19__21,
           q_cache_arr_19__20,q_cache_arr_19__19,q_cache_arr_19__18,
           q_cache_arr_19__17,q_cache_arr_19__16,q_cache_arr_19__15,
           q_cache_arr_19__14,q_cache_arr_19__13,q_cache_arr_19__12,
           q_cache_arr_19__11,q_cache_arr_19__10,q_cache_arr_19__9,
           q_cache_arr_19__8,q_cache_arr_19__7,q_cache_arr_19__6,
           q_cache_arr_19__5,q_cache_arr_19__4,q_cache_arr_19__3,
           q_cache_arr_19__2,q_cache_arr_19__1,q_cache_arr_19__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1113), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_20_gen_regi (.d ({d_cache_arr_20__31,
           d_cache_arr_20__30,d_cache_arr_20__29,d_cache_arr_20__28,
           d_cache_arr_20__27,d_cache_arr_20__26,d_cache_arr_20__25,
           d_cache_arr_20__24,d_cache_arr_20__23,d_cache_arr_20__22,
           d_cache_arr_20__21,d_cache_arr_20__20,d_cache_arr_20__19,
           d_cache_arr_20__18,d_cache_arr_20__17,d_cache_arr_20__16,
           d_cache_arr_20__15,d_cache_arr_20__14,d_cache_arr_20__13,
           d_cache_arr_20__12,d_cache_arr_20__11,d_cache_arr_20__10,
           d_cache_arr_20__9,d_cache_arr_20__8,d_cache_arr_20__7,
           d_cache_arr_20__6,d_cache_arr_20__5,d_cache_arr_20__4,
           d_cache_arr_20__3,d_cache_arr_20__2,d_cache_arr_20__1,
           d_cache_arr_20__0}), .q ({q_cache_arr_20__31,q_cache_arr_20__30,
           q_cache_arr_20__29,q_cache_arr_20__28,q_cache_arr_20__27,
           q_cache_arr_20__26,q_cache_arr_20__25,q_cache_arr_20__24,
           q_cache_arr_20__23,q_cache_arr_20__22,q_cache_arr_20__21,
           q_cache_arr_20__20,q_cache_arr_20__19,q_cache_arr_20__18,
           q_cache_arr_20__17,q_cache_arr_20__16,q_cache_arr_20__15,
           q_cache_arr_20__14,q_cache_arr_20__13,q_cache_arr_20__12,
           q_cache_arr_20__11,q_cache_arr_20__10,q_cache_arr_20__9,
           q_cache_arr_20__8,q_cache_arr_20__7,q_cache_arr_20__6,
           q_cache_arr_20__5,q_cache_arr_20__4,q_cache_arr_20__3,
           q_cache_arr_20__2,q_cache_arr_20__1,q_cache_arr_20__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1113), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_21_gen_regi (.d ({d_cache_arr_21__31,
           d_cache_arr_21__30,d_cache_arr_21__29,d_cache_arr_21__28,
           d_cache_arr_21__27,d_cache_arr_21__26,d_cache_arr_21__25,
           d_cache_arr_21__24,d_cache_arr_21__23,d_cache_arr_21__22,
           d_cache_arr_21__21,d_cache_arr_21__20,d_cache_arr_21__19,
           d_cache_arr_21__18,d_cache_arr_21__17,d_cache_arr_21__16,
           d_cache_arr_21__15,d_cache_arr_21__14,d_cache_arr_21__13,
           d_cache_arr_21__12,d_cache_arr_21__11,d_cache_arr_21__10,
           d_cache_arr_21__9,d_cache_arr_21__8,d_cache_arr_21__7,
           d_cache_arr_21__6,d_cache_arr_21__5,d_cache_arr_21__4,
           d_cache_arr_21__3,d_cache_arr_21__2,d_cache_arr_21__1,
           d_cache_arr_21__0}), .q ({q_cache_arr_21__31,q_cache_arr_21__30,
           q_cache_arr_21__29,q_cache_arr_21__28,q_cache_arr_21__27,
           q_cache_arr_21__26,q_cache_arr_21__25,q_cache_arr_21__24,
           q_cache_arr_21__23,q_cache_arr_21__22,q_cache_arr_21__21,
           q_cache_arr_21__20,q_cache_arr_21__19,q_cache_arr_21__18,
           q_cache_arr_21__17,q_cache_arr_21__16,q_cache_arr_21__15,
           q_cache_arr_21__14,q_cache_arr_21__13,q_cache_arr_21__12,
           q_cache_arr_21__11,q_cache_arr_21__10,q_cache_arr_21__9,
           q_cache_arr_21__8,q_cache_arr_21__7,q_cache_arr_21__6,
           q_cache_arr_21__5,q_cache_arr_21__4,q_cache_arr_21__3,
           q_cache_arr_21__2,q_cache_arr_21__1,q_cache_arr_21__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1115), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_22_gen_regi (.d ({d_cache_arr_22__31,
           d_cache_arr_22__30,d_cache_arr_22__29,d_cache_arr_22__28,
           d_cache_arr_22__27,d_cache_arr_22__26,d_cache_arr_22__25,
           d_cache_arr_22__24,d_cache_arr_22__23,d_cache_arr_22__22,
           d_cache_arr_22__21,d_cache_arr_22__20,d_cache_arr_22__19,
           d_cache_arr_22__18,d_cache_arr_22__17,d_cache_arr_22__16,
           d_cache_arr_22__15,d_cache_arr_22__14,d_cache_arr_22__13,
           d_cache_arr_22__12,d_cache_arr_22__11,d_cache_arr_22__10,
           d_cache_arr_22__9,d_cache_arr_22__8,d_cache_arr_22__7,
           d_cache_arr_22__6,d_cache_arr_22__5,d_cache_arr_22__4,
           d_cache_arr_22__3,d_cache_arr_22__2,d_cache_arr_22__1,
           d_cache_arr_22__0}), .q ({q_cache_arr_22__31,q_cache_arr_22__30,
           q_cache_arr_22__29,q_cache_arr_22__28,q_cache_arr_22__27,
           q_cache_arr_22__26,q_cache_arr_22__25,q_cache_arr_22__24,
           q_cache_arr_22__23,q_cache_arr_22__22,q_cache_arr_22__21,
           q_cache_arr_22__20,q_cache_arr_22__19,q_cache_arr_22__18,
           q_cache_arr_22__17,q_cache_arr_22__16,q_cache_arr_22__15,
           q_cache_arr_22__14,q_cache_arr_22__13,q_cache_arr_22__12,
           q_cache_arr_22__11,q_cache_arr_22__10,q_cache_arr_22__9,
           q_cache_arr_22__8,q_cache_arr_22__7,q_cache_arr_22__6,
           q_cache_arr_22__5,q_cache_arr_22__4,q_cache_arr_22__3,
           q_cache_arr_22__2,q_cache_arr_22__1,q_cache_arr_22__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1115), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_23_gen_regi (.d ({d_cache_arr_23__31,
           d_cache_arr_23__30,d_cache_arr_23__29,d_cache_arr_23__28,
           d_cache_arr_23__27,d_cache_arr_23__26,d_cache_arr_23__25,
           d_cache_arr_23__24,d_cache_arr_23__23,d_cache_arr_23__22,
           d_cache_arr_23__21,d_cache_arr_23__20,d_cache_arr_23__19,
           d_cache_arr_23__18,d_cache_arr_23__17,d_cache_arr_23__16,
           d_cache_arr_23__15,d_cache_arr_23__14,d_cache_arr_23__13,
           d_cache_arr_23__12,d_cache_arr_23__11,d_cache_arr_23__10,
           d_cache_arr_23__9,d_cache_arr_23__8,d_cache_arr_23__7,
           d_cache_arr_23__6,d_cache_arr_23__5,d_cache_arr_23__4,
           d_cache_arr_23__3,d_cache_arr_23__2,d_cache_arr_23__1,
           d_cache_arr_23__0}), .q ({q_cache_arr_23__31,q_cache_arr_23__30,
           q_cache_arr_23__29,q_cache_arr_23__28,q_cache_arr_23__27,
           q_cache_arr_23__26,q_cache_arr_23__25,q_cache_arr_23__24,
           q_cache_arr_23__23,q_cache_arr_23__22,q_cache_arr_23__21,
           q_cache_arr_23__20,q_cache_arr_23__19,q_cache_arr_23__18,
           q_cache_arr_23__17,q_cache_arr_23__16,q_cache_arr_23__15,
           q_cache_arr_23__14,q_cache_arr_23__13,q_cache_arr_23__12,
           q_cache_arr_23__11,q_cache_arr_23__10,q_cache_arr_23__9,
           q_cache_arr_23__8,q_cache_arr_23__7,q_cache_arr_23__6,
           q_cache_arr_23__5,q_cache_arr_23__4,q_cache_arr_23__3,
           q_cache_arr_23__2,q_cache_arr_23__1,q_cache_arr_23__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1115), .reset (
           filter_reset)) ;
    Reg_32 gen_comp_cache_gen_regs_24_gen_regi (.d ({d_cache_arr_24__31,
           d_cache_arr_24__30,d_cache_arr_24__29,d_cache_arr_24__28,
           d_cache_arr_24__27,d_cache_arr_24__26,d_cache_arr_24__25,
           d_cache_arr_24__24,d_cache_arr_24__23,d_cache_arr_24__22,
           d_cache_arr_24__21,d_cache_arr_24__20,d_cache_arr_24__19,
           d_cache_arr_24__18,d_cache_arr_24__17,d_cache_arr_24__16,
           d_cache_arr_24__15,d_cache_arr_24__14,d_cache_arr_24__13,
           d_cache_arr_24__12,d_cache_arr_24__11,d_cache_arr_24__10,
           d_cache_arr_24__9,d_cache_arr_24__8,d_cache_arr_24__7,
           d_cache_arr_24__6,d_cache_arr_24__5,d_cache_arr_24__4,
           d_cache_arr_24__3,d_cache_arr_24__2,d_cache_arr_24__1,
           d_cache_arr_24__0}), .q ({q_cache_arr_24__31,q_cache_arr_24__30,
           q_cache_arr_24__29,q_cache_arr_24__28,q_cache_arr_24__27,
           q_cache_arr_24__26,q_cache_arr_24__25,q_cache_arr_24__24,
           q_cache_arr_24__23,q_cache_arr_24__22,q_cache_arr_24__21,
           q_cache_arr_24__20,q_cache_arr_24__19,q_cache_arr_24__18,
           q_cache_arr_24__17,q_cache_arr_24__16,q_cache_arr_24__15,
           q_cache_arr_24__14,q_cache_arr_24__13,q_cache_arr_24__12,
           q_cache_arr_24__11,q_cache_arr_24__10,q_cache_arr_24__9,
           q_cache_arr_24__8,q_cache_arr_24__7,q_cache_arr_24__6,
           q_cache_arr_24__5,q_cache_arr_24__4,q_cache_arr_24__3,
           q_cache_arr_24__2,q_cache_arr_24__1,q_cache_arr_24__0}), .rst_data ({
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready,buffer_ready,buffer_ready,buffer_ready,
           buffer_ready,buffer_ready}), .clk (clk), .load (nx1115), .reset (
           filter_reset)) ;
    fake_gnd ix48 (.Y (buffer_ready)) ;
    dffs_ni reg_compute_relu_q (.Q (compute_relu_q), .QB (\$dummy [0]), .D (
            nx541), .CLK (nx1137), .S (filter_reset)) ;
    nand02 ix876 (.Y (nx875), .A0 (start), .A1 (ready)) ;
    dffs_ni reg_ready_q (.Q (ready), .QB (\$dummy [1]), .D (nx10), .CLK (nx1183)
            , .S (filter_reset)) ;
    inv01 ix11 (.Y (nx10), .A (nx879)) ;
    oai21 ix880 (.Y (nx879), .A0 (ready), .A1 (ready_tmp), .B0 (nx1151)) ;
    dffr reg_operation_q (.Q (operation_q), .QB (\$dummy [2]), .D (nx531), .CLK (
         nx1137), .R (filter_reset)) ;
    dffr reg_filter_size_q (.Q (filter_size_q), .QB (\$dummy [3]), .D (nx521), .CLK (
         nx1137), .R (filter_reset)) ;
    dffr reg_output2_init_q_0 (.Q (output2_init_q_0), .QB (\$dummy [4]), .D (
         nx361), .CLK (nx1137), .R (filter_reset)) ;
    dffr reg_output2_init_q_1 (.Q (output2_init_q_1), .QB (\$dummy [5]), .D (
         nx371), .CLK (nx1137), .R (filter_reset)) ;
    dffr reg_output2_init_q_2 (.Q (output2_init_q_2), .QB (\$dummy [6]), .D (
         nx381), .CLK (nx1137), .R (filter_reset)) ;
    dffr reg_output2_init_q_3 (.Q (output2_init_q_3), .QB (\$dummy [7]), .D (
         nx391), .CLK (nx1137), .R (filter_reset)) ;
    dffr reg_output2_init_q_4 (.Q (output2_init_q_4), .QB (\$dummy [8]), .D (
         nx401), .CLK (nx1139), .R (filter_reset)) ;
    dffr reg_output2_init_q_5 (.Q (output2_init_q_5), .QB (\$dummy [9]), .D (
         nx411), .CLK (nx1139), .R (filter_reset)) ;
    dffr reg_output2_init_q_6 (.Q (output2_init_q_6), .QB (\$dummy [10]), .D (
         nx421), .CLK (nx1139), .R (filter_reset)) ;
    dffr reg_output2_init_q_7 (.Q (output2_init_q_7), .QB (\$dummy [11]), .D (
         nx431), .CLK (nx1139), .R (filter_reset)) ;
    dffr reg_output2_init_q_8 (.Q (output2_init_q_8), .QB (\$dummy [12]), .D (
         nx441), .CLK (nx1139), .R (filter_reset)) ;
    dffr reg_output2_init_q_9 (.Q (output2_init_q_9), .QB (\$dummy [13]), .D (
         nx451), .CLK (nx1139), .R (filter_reset)) ;
    dffr reg_output2_init_q_10 (.Q (output2_init_q_10), .QB (\$dummy [14]), .D (
         nx461), .CLK (nx1139), .R (filter_reset)) ;
    dffr reg_output2_init_q_11 (.Q (output2_init_q_11), .QB (\$dummy [15]), .D (
         nx471), .CLK (nx1141), .R (filter_reset)) ;
    dffr reg_output2_init_q_12 (.Q (output2_init_q_12), .QB (\$dummy [16]), .D (
         nx481), .CLK (nx1141), .R (filter_reset)) ;
    dffr reg_output2_init_q_13 (.Q (output2_init_q_13), .QB (\$dummy [17]), .D (
         nx491), .CLK (nx1141), .R (filter_reset)) ;
    dffr reg_output2_init_q_14 (.Q (output2_init_q_14), .QB (\$dummy [18]), .D (
         nx501), .CLK (nx1141), .R (filter_reset)) ;
    dffr reg_output2_init_q_15 (.Q (output2_init_q_15), .QB (\$dummy [19]), .D (
         nx511), .CLK (nx1141), .R (filter_reset)) ;
    dffr reg_output1_init_q_0 (.Q (output1_init_q_0), .QB (\$dummy [20]), .D (
         nx201), .CLK (nx1141), .R (filter_reset)) ;
    dffr reg_output1_init_q_1 (.Q (output1_init_q_1), .QB (\$dummy [21]), .D (
         nx211), .CLK (nx1141), .R (filter_reset)) ;
    dffr reg_output1_init_q_2 (.Q (output1_init_q_2), .QB (\$dummy [22]), .D (
         nx221), .CLK (nx1143), .R (filter_reset)) ;
    dffr reg_output1_init_q_3 (.Q (output1_init_q_3), .QB (\$dummy [23]), .D (
         nx231), .CLK (nx1143), .R (filter_reset)) ;
    dffr reg_output1_init_q_4 (.Q (output1_init_q_4), .QB (\$dummy [24]), .D (
         nx241), .CLK (nx1143), .R (filter_reset)) ;
    dffr reg_output1_init_q_5 (.Q (output1_init_q_5), .QB (\$dummy [25]), .D (
         nx251), .CLK (nx1143), .R (filter_reset)) ;
    dffr reg_output1_init_q_6 (.Q (output1_init_q_6), .QB (\$dummy [26]), .D (
         nx261), .CLK (nx1143), .R (filter_reset)) ;
    dffr reg_output1_init_q_7 (.Q (output1_init_q_7), .QB (\$dummy [27]), .D (
         nx271), .CLK (nx1143), .R (filter_reset)) ;
    dffr reg_output1_init_q_8 (.Q (output1_init_q_8), .QB (\$dummy [28]), .D (
         nx281), .CLK (nx1143), .R (filter_reset)) ;
    dffr reg_output1_init_q_9 (.Q (output1_init_q_9), .QB (\$dummy [29]), .D (
         nx291), .CLK (nx1145), .R (filter_reset)) ;
    dffr reg_output1_init_q_10 (.Q (output1_init_q_10), .QB (\$dummy [30]), .D (
         nx301), .CLK (nx1145), .R (filter_reset)) ;
    dffr reg_output1_init_q_11 (.Q (output1_init_q_11), .QB (\$dummy [31]), .D (
         nx311), .CLK (nx1145), .R (filter_reset)) ;
    dffr reg_output1_init_q_12 (.Q (output1_init_q_12), .QB (\$dummy [32]), .D (
         nx321), .CLK (nx1145), .R (filter_reset)) ;
    dffr reg_output1_init_q_13 (.Q (output1_init_q_13), .QB (\$dummy [33]), .D (
         nx331), .CLK (nx1145), .R (filter_reset)) ;
    dffr reg_output1_init_q_14 (.Q (output1_init_q_14), .QB (\$dummy [34]), .D (
         nx341), .CLK (nx1145), .R (filter_reset)) ;
    dffr reg_output1_init_q_15 (.Q (output1_init_q_15), .QB (\$dummy [35]), .D (
         nx351), .CLK (nx1145), .R (filter_reset)) ;
    dffr reg_comp_pipe_en (.Q (comp_pipe_en), .QB (\$dummy [36]), .D (NOT_nx4), 
         .CLK (nx1147), .R (filter_reset)) ;
    nand02 ix987 (.Y (NOT_nx4), .A0 (ready_tmp), .A1 (nx1161)) ;
    dffs_ni reg_comp_pipe_rst (.Q (comp_pipe_rst), .QB (\$dummy [37]), .D (nx4)
            , .CLK (nx1147), .S (filter_reset)) ;
    and02 ix309 (.Y (filter_load_tmp), .A0 (filter_load), .A1 (buffer_ready_dup0
          )) ;
    dffs_ni reg_buffer_ready_q (.Q (buffer_ready_dup0), .QB (\$dummy [38]), .D (
            nx302), .CLK (nx1147), .S (filter_reset)) ;
    inv01 ix303 (.Y (nx302), .A (nx996)) ;
    oai21 ix997 (.Y (nx996), .A0 (buffer_ready_dup0), .A1 (buffer_ready_tmp), .B0 (
          nx1161)) ;
    and02 ix311 (.Y (img_load_tmp), .A0 (img_load), .A1 (buffer_ready_dup0)) ;
    dffr reg_output2_q_0 (.Q (output2[0]), .QB (\$dummy [39]), .D (nx711), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_1 (.Q (output2[1]), .QB (\$dummy [40]), .D (nx721), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_2 (.Q (output2[2]), .QB (\$dummy [41]), .D (nx731), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_3 (.Q (output2[3]), .QB (\$dummy [42]), .D (nx741), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_4 (.Q (output2[4]), .QB (\$dummy [43]), .D (nx751), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_5 (.Q (output2[5]), .QB (\$dummy [44]), .D (nx761), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_6 (.Q (output2[6]), .QB (\$dummy [45]), .D (nx771), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_7 (.Q (output2[7]), .QB (\$dummy [46]), .D (nx781), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_8 (.Q (output2[8]), .QB (\$dummy [47]), .D (nx791), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_9 (.Q (output2[9]), .QB (\$dummy [48]), .D (nx801), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_10 (.Q (output2[10]), .QB (\$dummy [49]), .D (nx811), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_11 (.Q (output2[11]), .QB (\$dummy [50]), .D (nx821), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_12 (.Q (output2[12]), .QB (\$dummy [51]), .D (nx831), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_13 (.Q (output2[13]), .QB (\$dummy [52]), .D (nx841), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_14 (.Q (output2[14]), .QB (\$dummy [53]), .D (nx851), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output2_q_15 (.Q (output2[15]), .QB (\$dummy [54]), .D (nx861), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_0 (.Q (output1[0]), .QB (\$dummy [55]), .D (nx551), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_1 (.Q (output1[1]), .QB (\$dummy [56]), .D (nx561), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_2 (.Q (output1[2]), .QB (\$dummy [57]), .D (nx571), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_3 (.Q (output1[3]), .QB (\$dummy [58]), .D (nx581), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_4 (.Q (output1[4]), .QB (\$dummy [59]), .D (nx591), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_5 (.Q (output1[5]), .QB (\$dummy [60]), .D (nx601), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_6 (.Q (output1[6]), .QB (\$dummy [61]), .D (nx611), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_7 (.Q (output1[7]), .QB (\$dummy [62]), .D (nx621), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_8 (.Q (output1[8]), .QB (\$dummy [63]), .D (nx631), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_9 (.Q (output1[9]), .QB (\$dummy [64]), .D (nx641), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_10 (.Q (output1[10]), .QB (\$dummy [65]), .D (nx651), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_11 (.Q (output1[11]), .QB (\$dummy [66]), .D (nx661), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_12 (.Q (output1[12]), .QB (\$dummy [67]), .D (nx671), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_13 (.Q (output1[13]), .QB (\$dummy [68]), .D (nx681), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_14 (.Q (output1[14]), .QB (\$dummy [69]), .D (nx691), .CLK (
         clk), .R (filter_reset)) ;
    dffr reg_output1_q_15 (.Q (output1[15]), .QB (\$dummy [70]), .D (nx701), .CLK (
         clk), .R (filter_reset)) ;
    inv01 ix5 (.Y (nx4), .A (NOT_nx4)) ;
    buf02 ix1102 (.Y (nx1103), .A (img_data_1__15)) ;
    buf02 ix1104 (.Y (nx1105), .A (img_data_2__15)) ;
    buf02 ix1106 (.Y (nx1107), .A (img_data_6__15)) ;
    inv01 ix1108 (.Y (nx1109), .A (nx1131)) ;
    inv01 ix1110 (.Y (nx1111), .A (nx1131)) ;
    inv01 ix1112 (.Y (nx1113), .A (nx1131)) ;
    inv01 ix1114 (.Y (nx1115), .A (nx1133)) ;
    inv01 ix1116 (.Y (nx1117), .A (filter_size_q)) ;
    inv01 ix1118 (.Y (nx1119), .A (nx1117)) ;
    inv01 ix1120 (.Y (nx1121), .A (nx1117)) ;
    inv02 ix1130 (.Y (nx1131), .A (nx1167)) ;
    inv02 ix1132 (.Y (nx1133), .A (nx1167)) ;
    inv02 ix1136 (.Y (nx1137), .A (clk)) ;
    inv02 ix1138 (.Y (nx1139), .A (clk)) ;
    inv02 ix1140 (.Y (nx1141), .A (clk)) ;
    inv02 ix1142 (.Y (nx1143), .A (clk)) ;
    inv02 ix1144 (.Y (nx1145), .A (clk)) ;
    inv02 ix1146 (.Y (nx1147), .A (clk)) ;
    inv02 ix1150 (.Y (nx1151), .A (nx1185)) ;
    inv02 ix1160 (.Y (nx1161), .A (nx1185)) ;
    mux21_ni ix542 (.Y (nx541), .A0 (compute_relu_q), .A1 (compute_relu), .S0 (
             nx1185)) ;
    mux21_ni ix532 (.Y (nx531), .A0 (operation_q), .A1 (operation), .S0 (nx1185)
             ) ;
    mux21_ni ix522 (.Y (nx521), .A0 (nx1121), .A1 (filter_size), .S0 (nx1185)) ;
    mux21_ni ix362 (.Y (nx361), .A0 (output2_init_q_0), .A1 (output2_init[0]), .S0 (
             nx1185)) ;
    mux21_ni ix372 (.Y (nx371), .A0 (output2_init_q_1), .A1 (output2_init[1]), .S0 (
             nx1185)) ;
    mux21_ni ix382 (.Y (nx381), .A0 (output2_init_q_2), .A1 (output2_init[2]), .S0 (
             nx1187)) ;
    mux21_ni ix392 (.Y (nx391), .A0 (output2_init_q_3), .A1 (output2_init[3]), .S0 (
             nx1187)) ;
    mux21_ni ix402 (.Y (nx401), .A0 (output2_init_q_4), .A1 (output2_init[4]), .S0 (
             nx1187)) ;
    mux21_ni ix412 (.Y (nx411), .A0 (output2_init_q_5), .A1 (output2_init[5]), .S0 (
             nx1187)) ;
    mux21_ni ix422 (.Y (nx421), .A0 (output2_init_q_6), .A1 (output2_init[6]), .S0 (
             nx1187)) ;
    mux21_ni ix432 (.Y (nx431), .A0 (output2_init_q_7), .A1 (output2_init[7]), .S0 (
             nx1187)) ;
    mux21_ni ix442 (.Y (nx441), .A0 (output2_init_q_8), .A1 (output2_init[8]), .S0 (
             nx1187)) ;
    mux21_ni ix452 (.Y (nx451), .A0 (output2_init_q_9), .A1 (output2_init[9]), .S0 (
             nx1189)) ;
    mux21_ni ix462 (.Y (nx461), .A0 (output2_init_q_10), .A1 (output2_init[10])
             , .S0 (nx1189)) ;
    mux21_ni ix472 (.Y (nx471), .A0 (output2_init_q_11), .A1 (output2_init[11])
             , .S0 (nx1189)) ;
    mux21_ni ix482 (.Y (nx481), .A0 (output2_init_q_12), .A1 (output2_init[12])
             , .S0 (nx1189)) ;
    mux21_ni ix492 (.Y (nx491), .A0 (output2_init_q_13), .A1 (output2_init[13])
             , .S0 (nx1189)) ;
    mux21_ni ix502 (.Y (nx501), .A0 (output2_init_q_14), .A1 (output2_init[14])
             , .S0 (nx1189)) ;
    mux21_ni ix512 (.Y (nx511), .A0 (output2_init_q_15), .A1 (output2_init[15])
             , .S0 (nx1189)) ;
    mux21_ni ix202 (.Y (nx201), .A0 (output1_init_q_0), .A1 (output1_init[0]), .S0 (
             nx1191)) ;
    mux21_ni ix212 (.Y (nx211), .A0 (output1_init_q_1), .A1 (output1_init[1]), .S0 (
             nx1191)) ;
    mux21_ni ix222 (.Y (nx221), .A0 (output1_init_q_2), .A1 (output1_init[2]), .S0 (
             nx1191)) ;
    mux21_ni ix232 (.Y (nx231), .A0 (output1_init_q_3), .A1 (output1_init[3]), .S0 (
             nx1191)) ;
    mux21_ni ix242 (.Y (nx241), .A0 (output1_init_q_4), .A1 (output1_init[4]), .S0 (
             nx1191)) ;
    mux21_ni ix252 (.Y (nx251), .A0 (output1_init_q_5), .A1 (output1_init[5]), .S0 (
             nx1191)) ;
    mux21_ni ix262 (.Y (nx261), .A0 (output1_init_q_6), .A1 (output1_init[6]), .S0 (
             nx1191)) ;
    mux21_ni ix272 (.Y (nx271), .A0 (output1_init_q_7), .A1 (output1_init[7]), .S0 (
             nx1193)) ;
    mux21_ni ix282 (.Y (nx281), .A0 (output1_init_q_8), .A1 (output1_init[8]), .S0 (
             nx1193)) ;
    mux21_ni ix292 (.Y (nx291), .A0 (output1_init_q_9), .A1 (output1_init[9]), .S0 (
             nx1193)) ;
    mux21_ni ix302 (.Y (nx301), .A0 (output1_init_q_10), .A1 (output1_init[10])
             , .S0 (nx1193)) ;
    mux21_ni ix312 (.Y (nx311), .A0 (output1_init_q_11), .A1 (output1_init[11])
             , .S0 (nx1193)) ;
    mux21_ni ix322 (.Y (nx321), .A0 (output1_init_q_12), .A1 (output1_init[12])
             , .S0 (nx1193)) ;
    mux21_ni ix332 (.Y (nx331), .A0 (output1_init_q_13), .A1 (output1_init[13])
             , .S0 (nx1193)) ;
    mux21_ni ix342 (.Y (nx341), .A0 (output1_init_q_14), .A1 (output1_init[14])
             , .S0 (nx1195)) ;
    mux21_ni ix352 (.Y (nx351), .A0 (output1_init_q_15), .A1 (output1_init[15])
             , .S0 (nx1195)) ;
    mux21_ni ix712 (.Y (nx711), .A0 (q_cache_arr_1__0), .A1 (output2[0]), .S0 (
             nx1167)) ;
    mux21_ni ix722 (.Y (nx721), .A0 (q_cache_arr_1__1), .A1 (output2[1]), .S0 (
             nx1167)) ;
    mux21_ni ix732 (.Y (nx731), .A0 (q_cache_arr_1__2), .A1 (output2[2]), .S0 (
             nx1167)) ;
    mux21_ni ix742 (.Y (nx741), .A0 (q_cache_arr_1__3), .A1 (output2[3]), .S0 (
             nx1167)) ;
    mux21_ni ix752 (.Y (nx751), .A0 (q_cache_arr_1__4), .A1 (output2[4]), .S0 (
             nx1167)) ;
    mux21_ni ix762 (.Y (nx761), .A0 (q_cache_arr_1__5), .A1 (output2[5]), .S0 (
             nx1169)) ;
    mux21_ni ix772 (.Y (nx771), .A0 (q_cache_arr_1__6), .A1 (output2[6]), .S0 (
             nx1169)) ;
    mux21_ni ix782 (.Y (nx781), .A0 (q_cache_arr_1__7), .A1 (output2[7]), .S0 (
             nx1169)) ;
    mux21_ni ix792 (.Y (nx791), .A0 (q_cache_arr_1__8), .A1 (output2[8]), .S0 (
             nx1169)) ;
    mux21_ni ix802 (.Y (nx801), .A0 (q_cache_arr_1__9), .A1 (output2[9]), .S0 (
             nx1169)) ;
    mux21_ni ix812 (.Y (nx811), .A0 (q_cache_arr_1__10), .A1 (output2[10]), .S0 (
             nx1169)) ;
    mux21_ni ix822 (.Y (nx821), .A0 (q_cache_arr_1__11), .A1 (output2[11]), .S0 (
             nx1169)) ;
    mux21_ni ix832 (.Y (nx831), .A0 (q_cache_arr_1__12), .A1 (output2[12]), .S0 (
             nx1171)) ;
    mux21_ni ix842 (.Y (nx841), .A0 (q_cache_arr_1__13), .A1 (output2[13]), .S0 (
             nx1171)) ;
    mux21_ni ix852 (.Y (nx851), .A0 (q_cache_arr_1__14), .A1 (output2[14]), .S0 (
             nx1171)) ;
    mux21_ni ix862 (.Y (nx861), .A0 (q_cache_arr_1__15), .A1 (output2[15]), .S0 (
             nx1171)) ;
    mux21_ni ix552 (.Y (nx551), .A0 (q_cache_arr_0__0), .A1 (output1[0]), .S0 (
             nx1171)) ;
    mux21_ni ix562 (.Y (nx561), .A0 (q_cache_arr_0__1), .A1 (output1[1]), .S0 (
             nx1171)) ;
    mux21_ni ix572 (.Y (nx571), .A0 (q_cache_arr_0__2), .A1 (output1[2]), .S0 (
             nx1171)) ;
    mux21_ni ix582 (.Y (nx581), .A0 (q_cache_arr_0__3), .A1 (output1[3]), .S0 (
             nx1173)) ;
    mux21_ni ix592 (.Y (nx591), .A0 (q_cache_arr_0__4), .A1 (output1[4]), .S0 (
             nx1173)) ;
    mux21_ni ix602 (.Y (nx601), .A0 (q_cache_arr_0__5), .A1 (output1[5]), .S0 (
             nx1173)) ;
    mux21_ni ix612 (.Y (nx611), .A0 (q_cache_arr_0__6), .A1 (output1[6]), .S0 (
             nx1173)) ;
    mux21_ni ix622 (.Y (nx621), .A0 (q_cache_arr_0__7), .A1 (output1[7]), .S0 (
             nx1173)) ;
    mux21_ni ix632 (.Y (nx631), .A0 (q_cache_arr_0__8), .A1 (output1[8]), .S0 (
             nx1173)) ;
    mux21_ni ix642 (.Y (nx641), .A0 (q_cache_arr_0__9), .A1 (output1[9]), .S0 (
             nx1173)) ;
    mux21_ni ix652 (.Y (nx651), .A0 (q_cache_arr_0__10), .A1 (output1[10]), .S0 (
             nx1175)) ;
    mux21_ni ix662 (.Y (nx661), .A0 (q_cache_arr_0__11), .A1 (output1[11]), .S0 (
             nx1175)) ;
    mux21_ni ix672 (.Y (nx671), .A0 (q_cache_arr_0__12), .A1 (output1[12]), .S0 (
             nx1175)) ;
    mux21_ni ix682 (.Y (nx681), .A0 (q_cache_arr_0__13), .A1 (output1[13]), .S0 (
             nx1175)) ;
    mux21_ni ix692 (.Y (nx691), .A0 (q_cache_arr_0__14), .A1 (output1[14]), .S0 (
             nx1175)) ;
    mux21_ni ix702 (.Y (nx701), .A0 (q_cache_arr_0__15), .A1 (output1[15]), .S0 (
             nx1175)) ;
    inv02 ix1166 (.Y (nx1167), .A (semi_ready)) ;
    inv02 ix1168 (.Y (nx1169), .A (semi_ready)) ;
    inv02 ix1170 (.Y (nx1171), .A (semi_ready)) ;
    inv02 ix1172 (.Y (nx1173), .A (semi_ready)) ;
    inv02 ix1174 (.Y (nx1175), .A (semi_ready)) ;
    buf02 ix1176 (.Y (nx1177), .A (img_load_tmp)) ;
    buf02 ix1178 (.Y (nx1179), .A (img_load_tmp)) ;
    inv02 ix1180 (.Y (nx1181), .A (clk)) ;
    inv02 ix1182 (.Y (nx1183), .A (clk)) ;
    inv02 ix1184 (.Y (nx1185), .A (nx875)) ;
    inv02 ix1186 (.Y (nx1187), .A (nx875)) ;
    inv02 ix1188 (.Y (nx1189), .A (nx875)) ;
    inv02 ix1190 (.Y (nx1191), .A (nx875)) ;
    inv02 ix1192 (.Y (nx1193), .A (nx875)) ;
    inv02 ix1194 (.Y (nx1195), .A (nx875)) ;
endmodule


module Reg_32 ( d, q, rst_data, clk, load, reset ) ;

    input [31:0]d ;
    output [31:0]q ;
    input [31:0]rst_data ;
    input clk ;
    input load ;
    input reset ;

    wire nx114, nx124, nx134, nx144, nx154, nx164, nx174, nx184, nx194, nx204, 
         nx214, nx224, nx234, nx244, nx254, nx264, nx274, nx284, nx294, nx304, 
         nx314, nx324, nx334, nx344, nx354, nx364, nx374, nx384, nx394, nx404, 
         nx414, nx424, nx535, nx537, nx539, nx541, nx543, nx545;
    wire [31:0] \$dummy ;




    dffr reg_q_0 (.Q (q[0]), .QB (\$dummy [0]), .D (nx114), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix115 (.Y (nx114), .A0 (q[0]), .A1 (d[0]), .S0 (nx537)) ;
    dffr reg_q_1 (.Q (q[1]), .QB (\$dummy [1]), .D (nx124), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix125 (.Y (nx124), .A0 (q[1]), .A1 (d[1]), .S0 (nx537)) ;
    dffr reg_q_2 (.Q (q[2]), .QB (\$dummy [2]), .D (nx134), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix135 (.Y (nx134), .A0 (q[2]), .A1 (d[2]), .S0 (nx537)) ;
    dffr reg_q_3 (.Q (q[3]), .QB (\$dummy [3]), .D (nx144), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix145 (.Y (nx144), .A0 (q[3]), .A1 (d[3]), .S0 (nx537)) ;
    dffr reg_q_4 (.Q (q[4]), .QB (\$dummy [4]), .D (nx154), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix155 (.Y (nx154), .A0 (q[4]), .A1 (d[4]), .S0 (nx537)) ;
    dffr reg_q_5 (.Q (q[5]), .QB (\$dummy [5]), .D (nx164), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix165 (.Y (nx164), .A0 (q[5]), .A1 (d[5]), .S0 (nx537)) ;
    dffr reg_q_6 (.Q (q[6]), .QB (\$dummy [6]), .D (nx174), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix175 (.Y (nx174), .A0 (q[6]), .A1 (d[6]), .S0 (nx537)) ;
    dffr reg_q_7 (.Q (q[7]), .QB (\$dummy [7]), .D (nx184), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix185 (.Y (nx184), .A0 (q[7]), .A1 (d[7]), .S0 (nx539)) ;
    dffr reg_q_8 (.Q (q[8]), .QB (\$dummy [8]), .D (nx194), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix195 (.Y (nx194), .A0 (q[8]), .A1 (d[8]), .S0 (nx539)) ;
    dffr reg_q_9 (.Q (q[9]), .QB (\$dummy [9]), .D (nx204), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix205 (.Y (nx204), .A0 (q[9]), .A1 (d[9]), .S0 (nx539)) ;
    dffr reg_q_10 (.Q (q[10]), .QB (\$dummy [10]), .D (nx214), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix215 (.Y (nx214), .A0 (q[10]), .A1 (d[10]), .S0 (nx539)) ;
    dffr reg_q_11 (.Q (q[11]), .QB (\$dummy [11]), .D (nx224), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix225 (.Y (nx224), .A0 (q[11]), .A1 (d[11]), .S0 (nx539)) ;
    dffr reg_q_12 (.Q (q[12]), .QB (\$dummy [12]), .D (nx234), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix235 (.Y (nx234), .A0 (q[12]), .A1 (d[12]), .S0 (nx539)) ;
    dffr reg_q_13 (.Q (q[13]), .QB (\$dummy [13]), .D (nx244), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix245 (.Y (nx244), .A0 (q[13]), .A1 (d[13]), .S0 (nx539)) ;
    dffr reg_q_14 (.Q (q[14]), .QB (\$dummy [14]), .D (nx254), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix255 (.Y (nx254), .A0 (q[14]), .A1 (d[14]), .S0 (nx541)) ;
    dffr reg_q_15 (.Q (q[15]), .QB (\$dummy [15]), .D (nx264), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix265 (.Y (nx264), .A0 (q[15]), .A1 (d[15]), .S0 (nx541)) ;
    dffr reg_q_16 (.Q (q[16]), .QB (\$dummy [16]), .D (nx274), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix275 (.Y (nx274), .A0 (q[16]), .A1 (d[16]), .S0 (nx541)) ;
    dffr reg_q_17 (.Q (q[17]), .QB (\$dummy [17]), .D (nx284), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix285 (.Y (nx284), .A0 (q[17]), .A1 (d[17]), .S0 (nx541)) ;
    dffr reg_q_18 (.Q (q[18]), .QB (\$dummy [18]), .D (nx294), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix295 (.Y (nx294), .A0 (q[18]), .A1 (d[18]), .S0 (nx541)) ;
    dffr reg_q_19 (.Q (q[19]), .QB (\$dummy [19]), .D (nx304), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix305 (.Y (nx304), .A0 (q[19]), .A1 (d[19]), .S0 (nx541)) ;
    dffr reg_q_20 (.Q (q[20]), .QB (\$dummy [20]), .D (nx314), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix315 (.Y (nx314), .A0 (q[20]), .A1 (d[20]), .S0 (nx541)) ;
    dffr reg_q_21 (.Q (q[21]), .QB (\$dummy [21]), .D (nx324), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix325 (.Y (nx324), .A0 (q[21]), .A1 (d[21]), .S0 (nx543)) ;
    dffr reg_q_22 (.Q (q[22]), .QB (\$dummy [22]), .D (nx334), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix335 (.Y (nx334), .A0 (q[22]), .A1 (d[22]), .S0 (nx543)) ;
    dffr reg_q_23 (.Q (q[23]), .QB (\$dummy [23]), .D (nx344), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix345 (.Y (nx344), .A0 (q[23]), .A1 (d[23]), .S0 (nx543)) ;
    dffr reg_q_24 (.Q (q[24]), .QB (\$dummy [24]), .D (nx354), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix355 (.Y (nx354), .A0 (q[24]), .A1 (d[24]), .S0 (nx543)) ;
    dffr reg_q_25 (.Q (q[25]), .QB (\$dummy [25]), .D (nx364), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix365 (.Y (nx364), .A0 (q[25]), .A1 (d[25]), .S0 (nx543)) ;
    dffr reg_q_26 (.Q (q[26]), .QB (\$dummy [26]), .D (nx374), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix375 (.Y (nx374), .A0 (q[26]), .A1 (d[26]), .S0 (nx543)) ;
    dffr reg_q_27 (.Q (q[27]), .QB (\$dummy [27]), .D (nx384), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix385 (.Y (nx384), .A0 (q[27]), .A1 (d[27]), .S0 (nx543)) ;
    dffr reg_q_28 (.Q (q[28]), .QB (\$dummy [28]), .D (nx394), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix395 (.Y (nx394), .A0 (q[28]), .A1 (d[28]), .S0 (nx545)) ;
    dffr reg_q_29 (.Q (q[29]), .QB (\$dummy [29]), .D (nx404), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix405 (.Y (nx404), .A0 (q[29]), .A1 (d[29]), .S0 (nx545)) ;
    dffr reg_q_30 (.Q (q[30]), .QB (\$dummy [30]), .D (nx414), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix415 (.Y (nx414), .A0 (q[30]), .A1 (d[30]), .S0 (nx545)) ;
    dffr reg_q_31 (.Q (q[31]), .QB (\$dummy [31]), .D (nx424), .CLK (clk), .R (
         reset)) ;
    mux21_ni ix425 (.Y (nx424), .A0 (q[31]), .A1 (d[31]), .S0 (nx545)) ;
    inv01 ix534 (.Y (nx535), .A (load)) ;
    inv02 ix536 (.Y (nx537), .A (nx535)) ;
    inv02 ix538 (.Y (nx539), .A (nx535)) ;
    inv02 ix540 (.Y (nx541), .A (nx535)) ;
    inv02 ix542 (.Y (nx543), .A (nx535)) ;
    inv02 ix544 (.Y (nx545), .A (nx535)) ;
endmodule


module Queue_25 ( d, q_0__15, q_0__14, q_0__13, q_0__12, q_0__11, q_0__10, 
                  q_0__9, q_0__8, q_0__7, q_0__6, q_0__5, q_0__4, q_0__3, q_0__2, 
                  q_0__1, q_0__0, q_1__15, q_1__14, q_1__13, q_1__12, q_1__11, 
                  q_1__10, q_1__9, q_1__8, q_1__7, q_1__6, q_1__5, q_1__4, 
                  q_1__3, q_1__2, q_1__1, q_1__0, q_2__15, q_2__14, q_2__13, 
                  q_2__12, q_2__11, q_2__10, q_2__9, q_2__8, q_2__7, q_2__6, 
                  q_2__5, q_2__4, q_2__3, q_2__2, q_2__1, q_2__0, q_3__15, 
                  q_3__14, q_3__13, q_3__12, q_3__11, q_3__10, q_3__9, q_3__8, 
                  q_3__7, q_3__6, q_3__5, q_3__4, q_3__3, q_3__2, q_3__1, q_3__0, 
                  q_4__15, q_4__14, q_4__13, q_4__12, q_4__11, q_4__10, q_4__9, 
                  q_4__8, q_4__7, q_4__6, q_4__5, q_4__4, q_4__3, q_4__2, q_4__1, 
                  q_4__0, q_5__15, q_5__14, q_5__13, q_5__12, q_5__11, q_5__10, 
                  q_5__9, q_5__8, q_5__7, q_5__6, q_5__5, q_5__4, q_5__3, q_5__2, 
                  q_5__1, q_5__0, q_6__15, q_6__14, q_6__13, q_6__12, q_6__11, 
                  q_6__10, q_6__9, q_6__8, q_6__7, q_6__6, q_6__5, q_6__4, 
                  q_6__3, q_6__2, q_6__1, q_6__0, q_7__15, q_7__14, q_7__13, 
                  q_7__12, q_7__11, q_7__10, q_7__9, q_7__8, q_7__7, q_7__6, 
                  q_7__5, q_7__4, q_7__3, q_7__2, q_7__1, q_7__0, q_8__15, 
                  q_8__14, q_8__13, q_8__12, q_8__11, q_8__10, q_8__9, q_8__8, 
                  q_8__7, q_8__6, q_8__5, q_8__4, q_8__3, q_8__2, q_8__1, q_8__0, 
                  q_9__15, q_9__14, q_9__13, q_9__12, q_9__11, q_9__10, q_9__9, 
                  q_9__8, q_9__7, q_9__6, q_9__5, q_9__4, q_9__3, q_9__2, q_9__1, 
                  q_9__0, q_10__15, q_10__14, q_10__13, q_10__12, q_10__11, 
                  q_10__10, q_10__9, q_10__8, q_10__7, q_10__6, q_10__5, q_10__4, 
                  q_10__3, q_10__2, q_10__1, q_10__0, q_11__15, q_11__14, 
                  q_11__13, q_11__12, q_11__11, q_11__10, q_11__9, q_11__8, 
                  q_11__7, q_11__6, q_11__5, q_11__4, q_11__3, q_11__2, q_11__1, 
                  q_11__0, q_12__15, q_12__14, q_12__13, q_12__12, q_12__11, 
                  q_12__10, q_12__9, q_12__8, q_12__7, q_12__6, q_12__5, q_12__4, 
                  q_12__3, q_12__2, q_12__1, q_12__0, q_13__15, q_13__14, 
                  q_13__13, q_13__12, q_13__11, q_13__10, q_13__9, q_13__8, 
                  q_13__7, q_13__6, q_13__5, q_13__4, q_13__3, q_13__2, q_13__1, 
                  q_13__0, q_14__15, q_14__14, q_14__13, q_14__12, q_14__11, 
                  q_14__10, q_14__9, q_14__8, q_14__7, q_14__6, q_14__5, q_14__4, 
                  q_14__3, q_14__2, q_14__1, q_14__0, q_15__15, q_15__14, 
                  q_15__13, q_15__12, q_15__11, q_15__10, q_15__9, q_15__8, 
                  q_15__7, q_15__6, q_15__5, q_15__4, q_15__3, q_15__2, q_15__1, 
                  q_15__0, q_16__15, q_16__14, q_16__13, q_16__12, q_16__11, 
                  q_16__10, q_16__9, q_16__8, q_16__7, q_16__6, q_16__5, q_16__4, 
                  q_16__3, q_16__2, q_16__1, q_16__0, q_17__15, q_17__14, 
                  q_17__13, q_17__12, q_17__11, q_17__10, q_17__9, q_17__8, 
                  q_17__7, q_17__6, q_17__5, q_17__4, q_17__3, q_17__2, q_17__1, 
                  q_17__0, q_18__15, q_18__14, q_18__13, q_18__12, q_18__11, 
                  q_18__10, q_18__9, q_18__8, q_18__7, q_18__6, q_18__5, q_18__4, 
                  q_18__3, q_18__2, q_18__1, q_18__0, q_19__15, q_19__14, 
                  q_19__13, q_19__12, q_19__11, q_19__10, q_19__9, q_19__8, 
                  q_19__7, q_19__6, q_19__5, q_19__4, q_19__3, q_19__2, q_19__1, 
                  q_19__0, q_20__15, q_20__14, q_20__13, q_20__12, q_20__11, 
                  q_20__10, q_20__9, q_20__8, q_20__7, q_20__6, q_20__5, q_20__4, 
                  q_20__3, q_20__2, q_20__1, q_20__0, q_21__15, q_21__14, 
                  q_21__13, q_21__12, q_21__11, q_21__10, q_21__9, q_21__8, 
                  q_21__7, q_21__6, q_21__5, q_21__4, q_21__3, q_21__2, q_21__1, 
                  q_21__0, q_22__15, q_22__14, q_22__13, q_22__12, q_22__11, 
                  q_22__10, q_22__9, q_22__8, q_22__7, q_22__6, q_22__5, q_22__4, 
                  q_22__3, q_22__2, q_22__1, q_22__0, q_23__15, q_23__14, 
                  q_23__13, q_23__12, q_23__11, q_23__10, q_23__9, q_23__8, 
                  q_23__7, q_23__6, q_23__5, q_23__4, q_23__3, q_23__2, q_23__1, 
                  q_23__0, q_24__15, q_24__14, q_24__13, q_24__12, q_24__11, 
                  q_24__10, q_24__9, q_24__8, q_24__7, q_24__6, q_24__5, q_24__4, 
                  q_24__3, q_24__2, q_24__1, q_24__0, clk, load, reset ) ;

    input [15:0]d ;
    output q_0__15 ;
    output q_0__14 ;
    output q_0__13 ;
    output q_0__12 ;
    output q_0__11 ;
    output q_0__10 ;
    output q_0__9 ;
    output q_0__8 ;
    output q_0__7 ;
    output q_0__6 ;
    output q_0__5 ;
    output q_0__4 ;
    output q_0__3 ;
    output q_0__2 ;
    output q_0__1 ;
    output q_0__0 ;
    output q_1__15 ;
    output q_1__14 ;
    output q_1__13 ;
    output q_1__12 ;
    output q_1__11 ;
    output q_1__10 ;
    output q_1__9 ;
    output q_1__8 ;
    output q_1__7 ;
    output q_1__6 ;
    output q_1__5 ;
    output q_1__4 ;
    output q_1__3 ;
    output q_1__2 ;
    output q_1__1 ;
    output q_1__0 ;
    output q_2__15 ;
    output q_2__14 ;
    output q_2__13 ;
    output q_2__12 ;
    output q_2__11 ;
    output q_2__10 ;
    output q_2__9 ;
    output q_2__8 ;
    output q_2__7 ;
    output q_2__6 ;
    output q_2__5 ;
    output q_2__4 ;
    output q_2__3 ;
    output q_2__2 ;
    output q_2__1 ;
    output q_2__0 ;
    output q_3__15 ;
    output q_3__14 ;
    output q_3__13 ;
    output q_3__12 ;
    output q_3__11 ;
    output q_3__10 ;
    output q_3__9 ;
    output q_3__8 ;
    output q_3__7 ;
    output q_3__6 ;
    output q_3__5 ;
    output q_3__4 ;
    output q_3__3 ;
    output q_3__2 ;
    output q_3__1 ;
    output q_3__0 ;
    output q_4__15 ;
    output q_4__14 ;
    output q_4__13 ;
    output q_4__12 ;
    output q_4__11 ;
    output q_4__10 ;
    output q_4__9 ;
    output q_4__8 ;
    output q_4__7 ;
    output q_4__6 ;
    output q_4__5 ;
    output q_4__4 ;
    output q_4__3 ;
    output q_4__2 ;
    output q_4__1 ;
    output q_4__0 ;
    output q_5__15 ;
    output q_5__14 ;
    output q_5__13 ;
    output q_5__12 ;
    output q_5__11 ;
    output q_5__10 ;
    output q_5__9 ;
    output q_5__8 ;
    output q_5__7 ;
    output q_5__6 ;
    output q_5__5 ;
    output q_5__4 ;
    output q_5__3 ;
    output q_5__2 ;
    output q_5__1 ;
    output q_5__0 ;
    output q_6__15 ;
    output q_6__14 ;
    output q_6__13 ;
    output q_6__12 ;
    output q_6__11 ;
    output q_6__10 ;
    output q_6__9 ;
    output q_6__8 ;
    output q_6__7 ;
    output q_6__6 ;
    output q_6__5 ;
    output q_6__4 ;
    output q_6__3 ;
    output q_6__2 ;
    output q_6__1 ;
    output q_6__0 ;
    output q_7__15 ;
    output q_7__14 ;
    output q_7__13 ;
    output q_7__12 ;
    output q_7__11 ;
    output q_7__10 ;
    output q_7__9 ;
    output q_7__8 ;
    output q_7__7 ;
    output q_7__6 ;
    output q_7__5 ;
    output q_7__4 ;
    output q_7__3 ;
    output q_7__2 ;
    output q_7__1 ;
    output q_7__0 ;
    output q_8__15 ;
    output q_8__14 ;
    output q_8__13 ;
    output q_8__12 ;
    output q_8__11 ;
    output q_8__10 ;
    output q_8__9 ;
    output q_8__8 ;
    output q_8__7 ;
    output q_8__6 ;
    output q_8__5 ;
    output q_8__4 ;
    output q_8__3 ;
    output q_8__2 ;
    output q_8__1 ;
    output q_8__0 ;
    output q_9__15 ;
    output q_9__14 ;
    output q_9__13 ;
    output q_9__12 ;
    output q_9__11 ;
    output q_9__10 ;
    output q_9__9 ;
    output q_9__8 ;
    output q_9__7 ;
    output q_9__6 ;
    output q_9__5 ;
    output q_9__4 ;
    output q_9__3 ;
    output q_9__2 ;
    output q_9__1 ;
    output q_9__0 ;
    output q_10__15 ;
    output q_10__14 ;
    output q_10__13 ;
    output q_10__12 ;
    output q_10__11 ;
    output q_10__10 ;
    output q_10__9 ;
    output q_10__8 ;
    output q_10__7 ;
    output q_10__6 ;
    output q_10__5 ;
    output q_10__4 ;
    output q_10__3 ;
    output q_10__2 ;
    output q_10__1 ;
    output q_10__0 ;
    output q_11__15 ;
    output q_11__14 ;
    output q_11__13 ;
    output q_11__12 ;
    output q_11__11 ;
    output q_11__10 ;
    output q_11__9 ;
    output q_11__8 ;
    output q_11__7 ;
    output q_11__6 ;
    output q_11__5 ;
    output q_11__4 ;
    output q_11__3 ;
    output q_11__2 ;
    output q_11__1 ;
    output q_11__0 ;
    output q_12__15 ;
    output q_12__14 ;
    output q_12__13 ;
    output q_12__12 ;
    output q_12__11 ;
    output q_12__10 ;
    output q_12__9 ;
    output q_12__8 ;
    output q_12__7 ;
    output q_12__6 ;
    output q_12__5 ;
    output q_12__4 ;
    output q_12__3 ;
    output q_12__2 ;
    output q_12__1 ;
    output q_12__0 ;
    output q_13__15 ;
    output q_13__14 ;
    output q_13__13 ;
    output q_13__12 ;
    output q_13__11 ;
    output q_13__10 ;
    output q_13__9 ;
    output q_13__8 ;
    output q_13__7 ;
    output q_13__6 ;
    output q_13__5 ;
    output q_13__4 ;
    output q_13__3 ;
    output q_13__2 ;
    output q_13__1 ;
    output q_13__0 ;
    output q_14__15 ;
    output q_14__14 ;
    output q_14__13 ;
    output q_14__12 ;
    output q_14__11 ;
    output q_14__10 ;
    output q_14__9 ;
    output q_14__8 ;
    output q_14__7 ;
    output q_14__6 ;
    output q_14__5 ;
    output q_14__4 ;
    output q_14__3 ;
    output q_14__2 ;
    output q_14__1 ;
    output q_14__0 ;
    output q_15__15 ;
    output q_15__14 ;
    output q_15__13 ;
    output q_15__12 ;
    output q_15__11 ;
    output q_15__10 ;
    output q_15__9 ;
    output q_15__8 ;
    output q_15__7 ;
    output q_15__6 ;
    output q_15__5 ;
    output q_15__4 ;
    output q_15__3 ;
    output q_15__2 ;
    output q_15__1 ;
    output q_15__0 ;
    output q_16__15 ;
    output q_16__14 ;
    output q_16__13 ;
    output q_16__12 ;
    output q_16__11 ;
    output q_16__10 ;
    output q_16__9 ;
    output q_16__8 ;
    output q_16__7 ;
    output q_16__6 ;
    output q_16__5 ;
    output q_16__4 ;
    output q_16__3 ;
    output q_16__2 ;
    output q_16__1 ;
    output q_16__0 ;
    output q_17__15 ;
    output q_17__14 ;
    output q_17__13 ;
    output q_17__12 ;
    output q_17__11 ;
    output q_17__10 ;
    output q_17__9 ;
    output q_17__8 ;
    output q_17__7 ;
    output q_17__6 ;
    output q_17__5 ;
    output q_17__4 ;
    output q_17__3 ;
    output q_17__2 ;
    output q_17__1 ;
    output q_17__0 ;
    output q_18__15 ;
    output q_18__14 ;
    output q_18__13 ;
    output q_18__12 ;
    output q_18__11 ;
    output q_18__10 ;
    output q_18__9 ;
    output q_18__8 ;
    output q_18__7 ;
    output q_18__6 ;
    output q_18__5 ;
    output q_18__4 ;
    output q_18__3 ;
    output q_18__2 ;
    output q_18__1 ;
    output q_18__0 ;
    output q_19__15 ;
    output q_19__14 ;
    output q_19__13 ;
    output q_19__12 ;
    output q_19__11 ;
    output q_19__10 ;
    output q_19__9 ;
    output q_19__8 ;
    output q_19__7 ;
    output q_19__6 ;
    output q_19__5 ;
    output q_19__4 ;
    output q_19__3 ;
    output q_19__2 ;
    output q_19__1 ;
    output q_19__0 ;
    output q_20__15 ;
    output q_20__14 ;
    output q_20__13 ;
    output q_20__12 ;
    output q_20__11 ;
    output q_20__10 ;
    output q_20__9 ;
    output q_20__8 ;
    output q_20__7 ;
    output q_20__6 ;
    output q_20__5 ;
    output q_20__4 ;
    output q_20__3 ;
    output q_20__2 ;
    output q_20__1 ;
    output q_20__0 ;
    output q_21__15 ;
    output q_21__14 ;
    output q_21__13 ;
    output q_21__12 ;
    output q_21__11 ;
    output q_21__10 ;
    output q_21__9 ;
    output q_21__8 ;
    output q_21__7 ;
    output q_21__6 ;
    output q_21__5 ;
    output q_21__4 ;
    output q_21__3 ;
    output q_21__2 ;
    output q_21__1 ;
    output q_21__0 ;
    output q_22__15 ;
    output q_22__14 ;
    output q_22__13 ;
    output q_22__12 ;
    output q_22__11 ;
    output q_22__10 ;
    output q_22__9 ;
    output q_22__8 ;
    output q_22__7 ;
    output q_22__6 ;
    output q_22__5 ;
    output q_22__4 ;
    output q_22__3 ;
    output q_22__2 ;
    output q_22__1 ;
    output q_22__0 ;
    output q_23__15 ;
    output q_23__14 ;
    output q_23__13 ;
    output q_23__12 ;
    output q_23__11 ;
    output q_23__10 ;
    output q_23__9 ;
    output q_23__8 ;
    output q_23__7 ;
    output q_23__6 ;
    output q_23__5 ;
    output q_23__4 ;
    output q_23__3 ;
    output q_23__2 ;
    output q_23__1 ;
    output q_23__0 ;
    output q_24__15 ;
    output q_24__14 ;
    output q_24__13 ;
    output q_24__12 ;
    output q_24__11 ;
    output q_24__10 ;
    output q_24__9 ;
    output q_24__8 ;
    output q_24__7 ;
    output q_24__6 ;
    output q_24__5 ;
    output q_24__4 ;
    output q_24__3 ;
    output q_24__2 ;
    output q_24__1 ;
    output q_24__0 ;
    input clk ;
    input load ;
    input reset ;

    wire nx1733, nx1743, nx1753, nx1763, nx1773, nx1783, nx1793, nx1803, nx1813, 
         nx1823, nx1833, nx1843, nx1853, nx1863, nx1873, nx1883, nx1893, nx1903, 
         nx1913, nx1923, nx1933, nx1943, nx1953, nx1963, nx1973, nx1983, nx1993, 
         nx2003, nx2013, nx2023, nx2033, nx2043, nx2053, nx2063, nx2073, nx2083, 
         nx2093, nx2103, nx2113, nx2123, nx2133, nx2143, nx2153, nx2163, nx2173, 
         nx2183, nx2193, nx2203, nx2213, nx2223, nx2233, nx2243, nx2253, nx2263, 
         nx2273, nx2283, nx2293, nx2303, nx2313, nx2323, nx2333, nx2343, nx2353, 
         nx2363, nx2373, nx2383, nx2393, nx2403, nx2413, nx2423, nx2433, nx2443, 
         nx2453, nx2463, nx2473, nx2483, nx2493, nx2503, nx2513, nx2523, nx2533, 
         nx2543, nx2553, nx2563, nx2573, nx2583, nx2593, nx2603, nx2613, nx2623, 
         nx2633, nx2643, nx2653, nx2663, nx2673, nx2683, nx2693, nx2703, nx2713, 
         nx2723, nx2733, nx2743, nx2753, nx2763, nx2773, nx2783, nx2793, nx2803, 
         nx2813, nx2823, nx2833, nx2843, nx2853, nx2863, nx2873, nx2883, nx2893, 
         nx2903, nx2913, nx2923, nx2933, nx2943, nx2953, nx2963, nx2973, nx2983, 
         nx2993, nx3003, nx3013, nx3023, nx3033, nx3043, nx3053, nx3063, nx3073, 
         nx3083, nx3093, nx3103, nx3113, nx3123, nx3133, nx3143, nx3153, nx3163, 
         nx3173, nx3183, nx3193, nx3203, nx3213, nx3223, nx3233, nx3243, nx3253, 
         nx3263, nx3273, nx3283, nx3293, nx3303, nx3313, nx3323, nx3333, nx3343, 
         nx3353, nx3363, nx3373, nx3383, nx3393, nx3403, nx3413, nx3423, nx3433, 
         nx3443, nx3453, nx3463, nx3473, nx3483, nx3493, nx3503, nx3513, nx3523, 
         nx3533, nx3543, nx3553, nx3563, nx3573, nx3583, nx3593, nx3603, nx3613, 
         nx3623, nx3633, nx3643, nx3653, nx3663, nx3673, nx3683, nx3693, nx3703, 
         nx3713, nx3723, nx3733, nx3743, nx3753, nx3763, nx3773, nx3783, nx3793, 
         nx3803, nx3813, nx3823, nx3833, nx3843, nx3853, nx3863, nx3873, nx3883, 
         nx3893, nx3903, nx3913, nx3923, nx3933, nx3943, nx3953, nx3963, nx3973, 
         nx3983, nx3993, nx4003, nx4013, nx4023, nx4033, nx4043, nx4053, nx4063, 
         nx4073, nx4083, nx4093, nx4103, nx4113, nx4123, nx4133, nx4143, nx4153, 
         nx4163, nx4173, nx4183, nx4193, nx4203, nx4213, nx4223, nx4233, nx4243, 
         nx4253, nx4263, nx4273, nx4283, nx4293, nx4303, nx4313, nx4323, nx4333, 
         nx4343, nx4353, nx4363, nx4373, nx4383, nx4393, nx4403, nx4413, nx4423, 
         nx4433, nx4443, nx4453, nx4463, nx4473, nx4483, nx4493, nx4503, nx4513, 
         nx4523, nx4533, nx4543, nx4553, nx4563, nx4573, nx4583, nx4593, nx4603, 
         nx4613, nx4623, nx4633, nx4643, nx4653, nx4663, nx4673, nx4683, nx4693, 
         nx4703, nx4713, nx4723, nx4733, nx4743, nx4753, nx4763, nx4773, nx4783, 
         nx4793, nx4803, nx4813, nx4823, nx4833, nx4843, nx4853, nx4863, nx4873, 
         nx4883, nx4893, nx4903, nx4913, nx4923, nx4933, nx4943, nx4953, nx4963, 
         nx4973, nx4983, nx4993, nx5003, nx5013, nx5023, nx5033, nx5043, nx5053, 
         nx5063, nx5073, nx5083, nx5093, nx5103, nx5113, nx5123, nx5133, nx5143, 
         nx5153, nx5163, nx5173, nx5183, nx5193, nx5203, nx5213, nx5223, nx5233, 
         nx5243, nx5253, nx5263, nx5273, nx5283, nx5293, nx5303, nx5313, nx5323, 
         nx5333, nx5343, nx5353, nx5363, nx5373, nx5383, nx5393, nx5403, nx5413, 
         nx5423, nx5433, nx5443, nx5453, nx5463, nx5473, nx5483, nx5493, nx5503, 
         nx5513, nx5523, nx5533, nx5543, nx5553, nx5563, nx5573, nx5583, nx5593, 
         nx5603, nx5613, nx5623, nx5633, nx5643, nx5653, nx5663, nx5673, nx5683, 
         nx5693, nx5703, nx5713, nx5723, nx6940, nx6942, nx6944, nx6946, nx6948, 
         nx6950, nx6952, nx6954, nx6956, nx6958, nx6960, nx6962, nx6964, nx6966, 
         nx6968, nx6970, nx6972, nx6974, nx6976, nx6978, nx6980, nx6982, nx6984, 
         nx6986, nx6988, nx6990, nx6992, nx6994, nx6996, nx6998, nx7000, nx7002, 
         nx7004, nx7006, nx7008, nx7010, nx7012, nx7014, nx7016, nx7018, nx7020, 
         nx7022, nx7024, nx7026, nx7028, nx7030, nx7032, nx7034, nx7036, nx7038, 
         nx7040, nx7042, nx7044, nx7046, nx7048, nx7050, nx7052, nx7054, nx7058, 
         nx7060, nx7062, nx7064, nx7066, nx7068, nx7070, nx7072, nx7074, nx7076, 
         nx7078, nx7080, nx7082, nx7084, nx7086, nx7088, nx7090, nx7092, nx7094, 
         nx7096, nx7098, nx7100, nx7102, nx7104, nx7106, nx7108, nx7110, nx7112, 
         nx7114, nx7116, nx7118, nx7120, nx7122, nx7124, nx7126, nx7128, nx7130, 
         nx7132, nx7134, nx7136, nx7138, nx7140, nx7142, nx7144, nx7146, nx7148, 
         nx7150, nx7152, nx7154, nx7156, nx7158, nx7160, nx7162, nx7164, nx7166, 
         nx7168, nx7170, nx7172, nx7174, nx7176, nx7178, nx7180, nx7182, nx7184, 
         nx7186, nx7188, nx7190, nx7192, nx7194, nx7196, nx7198, nx7200, nx7202, 
         nx7204, nx7206, nx7208, nx7214, nx7216, nx7218, nx7220, nx7626, nx7628;
    wire [399:0] \$dummy ;




    dffr gen_regs_24_regi_reg_q_0 (.Q (q_24__0), .QB (\$dummy [0]), .D (nx1973)
         , .CLK (nx7064), .R (reset)) ;
    mux21_ni ix1974 (.Y (nx1973), .A0 (q_24__0), .A1 (q_23__0), .S0 (nx6946)) ;
    dffr gen_regs_23_regi_reg_q_0 (.Q (q_23__0), .QB (\$dummy [1]), .D (nx1963)
         , .CLK (nx7064), .R (reset)) ;
    mux21_ni ix1964 (.Y (nx1963), .A0 (q_23__0), .A1 (q_22__0), .S0 (nx6946)) ;
    dffr gen_regs_22_regi_reg_q_0 (.Q (q_22__0), .QB (\$dummy [2]), .D (nx1953)
         , .CLK (nx7064), .R (reset)) ;
    mux21_ni ix1954 (.Y (nx1953), .A0 (q_22__0), .A1 (q_21__0), .S0 (nx6946)) ;
    dffr gen_regs_21_regi_reg_q_0 (.Q (q_21__0), .QB (\$dummy [3]), .D (nx1943)
         , .CLK (nx7064), .R (reset)) ;
    mux21_ni ix1944 (.Y (nx1943), .A0 (q_21__0), .A1 (q_20__0), .S0 (nx6946)) ;
    dffr gen_regs_20_regi_reg_q_0 (.Q (q_20__0), .QB (\$dummy [4]), .D (nx1933)
         , .CLK (nx7062), .R (reset)) ;
    mux21_ni ix1934 (.Y (nx1933), .A0 (q_20__0), .A1 (q_19__0), .S0 (nx6944)) ;
    dffr gen_regs_19_regi_reg_q_0 (.Q (q_19__0), .QB (\$dummy [5]), .D (nx1923)
         , .CLK (nx7062), .R (reset)) ;
    mux21_ni ix1924 (.Y (nx1923), .A0 (q_19__0), .A1 (q_18__0), .S0 (nx6944)) ;
    dffr gen_regs_18_regi_reg_q_0 (.Q (q_18__0), .QB (\$dummy [6]), .D (nx1913)
         , .CLK (nx7062), .R (reset)) ;
    mux21_ni ix1914 (.Y (nx1913), .A0 (q_18__0), .A1 (q_17__0), .S0 (nx6944)) ;
    dffr gen_regs_17_regi_reg_q_0 (.Q (q_17__0), .QB (\$dummy [7]), .D (nx1903)
         , .CLK (nx7062), .R (reset)) ;
    mux21_ni ix1904 (.Y (nx1903), .A0 (q_17__0), .A1 (q_16__0), .S0 (nx6944)) ;
    dffr gen_regs_16_regi_reg_q_0 (.Q (q_16__0), .QB (\$dummy [8]), .D (nx1893)
         , .CLK (nx7062), .R (reset)) ;
    mux21_ni ix1894 (.Y (nx1893), .A0 (q_16__0), .A1 (q_15__0), .S0 (nx6944)) ;
    dffr gen_regs_15_regi_reg_q_0 (.Q (q_15__0), .QB (\$dummy [9]), .D (nx1883)
         , .CLK (nx7062), .R (reset)) ;
    mux21_ni ix1884 (.Y (nx1883), .A0 (q_15__0), .A1 (q_14__0), .S0 (nx6944)) ;
    dffr gen_regs_14_regi_reg_q_0 (.Q (q_14__0), .QB (\$dummy [10]), .D (nx1873)
         , .CLK (nx7062), .R (reset)) ;
    mux21_ni ix1874 (.Y (nx1873), .A0 (q_14__0), .A1 (q_13__0), .S0 (nx6944)) ;
    dffr gen_regs_13_regi_reg_q_0 (.Q (q_13__0), .QB (\$dummy [11]), .D (nx1863)
         , .CLK (nx7060), .R (reset)) ;
    mux21_ni ix1864 (.Y (nx1863), .A0 (q_13__0), .A1 (q_12__0), .S0 (nx6942)) ;
    dffr gen_regs_12_regi_reg_q_0 (.Q (q_12__0), .QB (\$dummy [12]), .D (nx1853)
         , .CLK (nx7060), .R (reset)) ;
    mux21_ni ix1854 (.Y (nx1853), .A0 (q_12__0), .A1 (q_11__0), .S0 (nx6942)) ;
    dffr gen_regs_11_regi_reg_q_0 (.Q (q_11__0), .QB (\$dummy [13]), .D (nx1843)
         , .CLK (nx7060), .R (reset)) ;
    mux21_ni ix1844 (.Y (nx1843), .A0 (q_11__0), .A1 (q_10__0), .S0 (nx6942)) ;
    dffr gen_regs_10_regi_reg_q_0 (.Q (q_10__0), .QB (\$dummy [14]), .D (nx1833)
         , .CLK (nx7060), .R (reset)) ;
    mux21_ni ix1834 (.Y (nx1833), .A0 (q_10__0), .A1 (q_9__0), .S0 (nx6942)) ;
    dffr gen_regs_9_regi_reg_q_0 (.Q (q_9__0), .QB (\$dummy [15]), .D (nx1823), 
         .CLK (nx7060), .R (reset)) ;
    mux21_ni ix1824 (.Y (nx1823), .A0 (q_9__0), .A1 (q_8__0), .S0 (nx6942)) ;
    dffr gen_regs_8_regi_reg_q_0 (.Q (q_8__0), .QB (\$dummy [16]), .D (nx1813), 
         .CLK (nx7060), .R (reset)) ;
    mux21_ni ix1814 (.Y (nx1813), .A0 (q_8__0), .A1 (q_7__0), .S0 (nx6942)) ;
    dffr gen_regs_7_regi_reg_q_0 (.Q (q_7__0), .QB (\$dummy [17]), .D (nx1803), 
         .CLK (nx7060), .R (reset)) ;
    mux21_ni ix1804 (.Y (nx1803), .A0 (q_7__0), .A1 (q_6__0), .S0 (nx6942)) ;
    dffr gen_regs_6_regi_reg_q_0 (.Q (q_6__0), .QB (\$dummy [18]), .D (nx1793), 
         .CLK (nx7058), .R (reset)) ;
    mux21_ni ix1794 (.Y (nx1793), .A0 (q_6__0), .A1 (q_5__0), .S0 (nx6940)) ;
    dffr gen_regs_5_regi_reg_q_0 (.Q (q_5__0), .QB (\$dummy [19]), .D (nx1783), 
         .CLK (nx7058), .R (reset)) ;
    mux21_ni ix1784 (.Y (nx1783), .A0 (q_5__0), .A1 (q_4__0), .S0 (nx6940)) ;
    dffr gen_regs_4_regi_reg_q_0 (.Q (q_4__0), .QB (\$dummy [20]), .D (nx1773), 
         .CLK (nx7058), .R (reset)) ;
    mux21_ni ix1774 (.Y (nx1773), .A0 (q_4__0), .A1 (q_3__0), .S0 (nx6940)) ;
    dffr gen_regs_3_regi_reg_q_0 (.Q (q_3__0), .QB (\$dummy [21]), .D (nx1763), 
         .CLK (nx7058), .R (reset)) ;
    mux21_ni ix1764 (.Y (nx1763), .A0 (q_3__0), .A1 (q_2__0), .S0 (nx6940)) ;
    dffr gen_regs_2_regi_reg_q_0 (.Q (q_2__0), .QB (\$dummy [22]), .D (nx1753), 
         .CLK (nx7058), .R (reset)) ;
    mux21_ni ix1754 (.Y (nx1753), .A0 (q_2__0), .A1 (q_1__0), .S0 (nx6940)) ;
    dffr gen_regs_1_regi_reg_q_0 (.Q (q_1__0), .QB (\$dummy [23]), .D (nx1743), 
         .CLK (nx7058), .R (reset)) ;
    mux21_ni ix1744 (.Y (nx1743), .A0 (q_1__0), .A1 (q_0__0), .S0 (nx6940)) ;
    dffr reg0_reg_q_0 (.Q (q_0__0), .QB (\$dummy [24]), .D (nx1733), .CLK (
         nx7058), .R (reset)) ;
    mux21_ni ix1734 (.Y (nx1733), .A0 (q_0__0), .A1 (d[0]), .S0 (nx6940)) ;
    dffr gen_regs_24_regi_reg_q_1 (.Q (q_24__1), .QB (\$dummy [25]), .D (nx2223)
         , .CLK (nx7072), .R (reset)) ;
    mux21_ni ix2224 (.Y (nx2223), .A0 (q_24__1), .A1 (q_23__1), .S0 (nx6954)) ;
    dffr gen_regs_23_regi_reg_q_1 (.Q (q_23__1), .QB (\$dummy [26]), .D (nx2213)
         , .CLK (nx7070), .R (reset)) ;
    mux21_ni ix2214 (.Y (nx2213), .A0 (q_23__1), .A1 (q_22__1), .S0 (nx6952)) ;
    dffr gen_regs_22_regi_reg_q_1 (.Q (q_22__1), .QB (\$dummy [27]), .D (nx2203)
         , .CLK (nx7070), .R (reset)) ;
    mux21_ni ix2204 (.Y (nx2203), .A0 (q_22__1), .A1 (q_21__1), .S0 (nx6952)) ;
    dffr gen_regs_21_regi_reg_q_1 (.Q (q_21__1), .QB (\$dummy [28]), .D (nx2193)
         , .CLK (nx7070), .R (reset)) ;
    mux21_ni ix2194 (.Y (nx2193), .A0 (q_21__1), .A1 (q_20__1), .S0 (nx6952)) ;
    dffr gen_regs_20_regi_reg_q_1 (.Q (q_20__1), .QB (\$dummy [29]), .D (nx2183)
         , .CLK (nx7070), .R (reset)) ;
    mux21_ni ix2184 (.Y (nx2183), .A0 (q_20__1), .A1 (q_19__1), .S0 (nx6952)) ;
    dffr gen_regs_19_regi_reg_q_1 (.Q (q_19__1), .QB (\$dummy [30]), .D (nx2173)
         , .CLK (nx7070), .R (reset)) ;
    mux21_ni ix2174 (.Y (nx2173), .A0 (q_19__1), .A1 (q_18__1), .S0 (nx6952)) ;
    dffr gen_regs_18_regi_reg_q_1 (.Q (q_18__1), .QB (\$dummy [31]), .D (nx2163)
         , .CLK (nx7070), .R (reset)) ;
    mux21_ni ix2164 (.Y (nx2163), .A0 (q_18__1), .A1 (q_17__1), .S0 (nx6952)) ;
    dffr gen_regs_17_regi_reg_q_1 (.Q (q_17__1), .QB (\$dummy [32]), .D (nx2153)
         , .CLK (nx7070), .R (reset)) ;
    mux21_ni ix2154 (.Y (nx2153), .A0 (q_17__1), .A1 (q_16__1), .S0 (nx6952)) ;
    dffr gen_regs_16_regi_reg_q_1 (.Q (q_16__1), .QB (\$dummy [33]), .D (nx2143)
         , .CLK (nx7068), .R (reset)) ;
    mux21_ni ix2144 (.Y (nx2143), .A0 (q_16__1), .A1 (q_15__1), .S0 (nx6950)) ;
    dffr gen_regs_15_regi_reg_q_1 (.Q (q_15__1), .QB (\$dummy [34]), .D (nx2133)
         , .CLK (nx7068), .R (reset)) ;
    mux21_ni ix2134 (.Y (nx2133), .A0 (q_15__1), .A1 (q_14__1), .S0 (nx6950)) ;
    dffr gen_regs_14_regi_reg_q_1 (.Q (q_14__1), .QB (\$dummy [35]), .D (nx2123)
         , .CLK (nx7068), .R (reset)) ;
    mux21_ni ix2124 (.Y (nx2123), .A0 (q_14__1), .A1 (q_13__1), .S0 (nx6950)) ;
    dffr gen_regs_13_regi_reg_q_1 (.Q (q_13__1), .QB (\$dummy [36]), .D (nx2113)
         , .CLK (nx7068), .R (reset)) ;
    mux21_ni ix2114 (.Y (nx2113), .A0 (q_13__1), .A1 (q_12__1), .S0 (nx6950)) ;
    dffr gen_regs_12_regi_reg_q_1 (.Q (q_12__1), .QB (\$dummy [37]), .D (nx2103)
         , .CLK (nx7068), .R (reset)) ;
    mux21_ni ix2104 (.Y (nx2103), .A0 (q_12__1), .A1 (q_11__1), .S0 (nx6950)) ;
    dffr gen_regs_11_regi_reg_q_1 (.Q (q_11__1), .QB (\$dummy [38]), .D (nx2093)
         , .CLK (nx7068), .R (reset)) ;
    mux21_ni ix2094 (.Y (nx2093), .A0 (q_11__1), .A1 (q_10__1), .S0 (nx6950)) ;
    dffr gen_regs_10_regi_reg_q_1 (.Q (q_10__1), .QB (\$dummy [39]), .D (nx2083)
         , .CLK (nx7068), .R (reset)) ;
    mux21_ni ix2084 (.Y (nx2083), .A0 (q_10__1), .A1 (q_9__1), .S0 (nx6950)) ;
    dffr gen_regs_9_regi_reg_q_1 (.Q (q_9__1), .QB (\$dummy [40]), .D (nx2073), 
         .CLK (nx7066), .R (reset)) ;
    mux21_ni ix2074 (.Y (nx2073), .A0 (q_9__1), .A1 (q_8__1), .S0 (nx6948)) ;
    dffr gen_regs_8_regi_reg_q_1 (.Q (q_8__1), .QB (\$dummy [41]), .D (nx2063), 
         .CLK (nx7066), .R (reset)) ;
    mux21_ni ix2064 (.Y (nx2063), .A0 (q_8__1), .A1 (q_7__1), .S0 (nx6948)) ;
    dffr gen_regs_7_regi_reg_q_1 (.Q (q_7__1), .QB (\$dummy [42]), .D (nx2053), 
         .CLK (nx7066), .R (reset)) ;
    mux21_ni ix2054 (.Y (nx2053), .A0 (q_7__1), .A1 (q_6__1), .S0 (nx6948)) ;
    dffr gen_regs_6_regi_reg_q_1 (.Q (q_6__1), .QB (\$dummy [43]), .D (nx2043), 
         .CLK (nx7066), .R (reset)) ;
    mux21_ni ix2044 (.Y (nx2043), .A0 (q_6__1), .A1 (q_5__1), .S0 (nx6948)) ;
    dffr gen_regs_5_regi_reg_q_1 (.Q (q_5__1), .QB (\$dummy [44]), .D (nx2033), 
         .CLK (nx7066), .R (reset)) ;
    mux21_ni ix2034 (.Y (nx2033), .A0 (q_5__1), .A1 (q_4__1), .S0 (nx6948)) ;
    dffr gen_regs_4_regi_reg_q_1 (.Q (q_4__1), .QB (\$dummy [45]), .D (nx2023), 
         .CLK (nx7066), .R (reset)) ;
    mux21_ni ix2024 (.Y (nx2023), .A0 (q_4__1), .A1 (q_3__1), .S0 (nx6948)) ;
    dffr gen_regs_3_regi_reg_q_1 (.Q (q_3__1), .QB (\$dummy [46]), .D (nx2013), 
         .CLK (nx7066), .R (reset)) ;
    mux21_ni ix2014 (.Y (nx2013), .A0 (q_3__1), .A1 (q_2__1), .S0 (nx6948)) ;
    dffr gen_regs_2_regi_reg_q_1 (.Q (q_2__1), .QB (\$dummy [47]), .D (nx2003), 
         .CLK (nx7064), .R (reset)) ;
    mux21_ni ix2004 (.Y (nx2003), .A0 (q_2__1), .A1 (q_1__1), .S0 (nx6946)) ;
    dffr gen_regs_1_regi_reg_q_1 (.Q (q_1__1), .QB (\$dummy [48]), .D (nx1993), 
         .CLK (nx7064), .R (reset)) ;
    mux21_ni ix1994 (.Y (nx1993), .A0 (q_1__1), .A1 (q_0__1), .S0 (nx6946)) ;
    dffr reg0_reg_q_1 (.Q (q_0__1), .QB (\$dummy [49]), .D (nx1983), .CLK (
         nx7064), .R (reset)) ;
    mux21_ni ix1984 (.Y (nx1983), .A0 (q_0__1), .A1 (d[1]), .S0 (nx6946)) ;
    dffr gen_regs_24_regi_reg_q_2 (.Q (q_24__2), .QB (\$dummy [50]), .D (nx2473)
         , .CLK (nx7078), .R (reset)) ;
    mux21_ni ix2474 (.Y (nx2473), .A0 (q_24__2), .A1 (q_23__2), .S0 (nx6960)) ;
    dffr gen_regs_23_regi_reg_q_2 (.Q (q_23__2), .QB (\$dummy [51]), .D (nx2463)
         , .CLK (nx7078), .R (reset)) ;
    mux21_ni ix2464 (.Y (nx2463), .A0 (q_23__2), .A1 (q_22__2), .S0 (nx6960)) ;
    dffr gen_regs_22_regi_reg_q_2 (.Q (q_22__2), .QB (\$dummy [52]), .D (nx2453)
         , .CLK (nx7078), .R (reset)) ;
    mux21_ni ix2454 (.Y (nx2453), .A0 (q_22__2), .A1 (q_21__2), .S0 (nx6960)) ;
    dffr gen_regs_21_regi_reg_q_2 (.Q (q_21__2), .QB (\$dummy [53]), .D (nx2443)
         , .CLK (nx7078), .R (reset)) ;
    mux21_ni ix2444 (.Y (nx2443), .A0 (q_21__2), .A1 (q_20__2), .S0 (nx6960)) ;
    dffr gen_regs_20_regi_reg_q_2 (.Q (q_20__2), .QB (\$dummy [54]), .D (nx2433)
         , .CLK (nx7078), .R (reset)) ;
    mux21_ni ix2434 (.Y (nx2433), .A0 (q_20__2), .A1 (q_19__2), .S0 (nx6960)) ;
    dffr gen_regs_19_regi_reg_q_2 (.Q (q_19__2), .QB (\$dummy [55]), .D (nx2423)
         , .CLK (nx7076), .R (reset)) ;
    mux21_ni ix2424 (.Y (nx2423), .A0 (q_19__2), .A1 (q_18__2), .S0 (nx6958)) ;
    dffr gen_regs_18_regi_reg_q_2 (.Q (q_18__2), .QB (\$dummy [56]), .D (nx2413)
         , .CLK (nx7076), .R (reset)) ;
    mux21_ni ix2414 (.Y (nx2413), .A0 (q_18__2), .A1 (q_17__2), .S0 (nx6958)) ;
    dffr gen_regs_17_regi_reg_q_2 (.Q (q_17__2), .QB (\$dummy [57]), .D (nx2403)
         , .CLK (nx7076), .R (reset)) ;
    mux21_ni ix2404 (.Y (nx2403), .A0 (q_17__2), .A1 (q_16__2), .S0 (nx6958)) ;
    dffr gen_regs_16_regi_reg_q_2 (.Q (q_16__2), .QB (\$dummy [58]), .D (nx2393)
         , .CLK (nx7076), .R (reset)) ;
    mux21_ni ix2394 (.Y (nx2393), .A0 (q_16__2), .A1 (q_15__2), .S0 (nx6958)) ;
    dffr gen_regs_15_regi_reg_q_2 (.Q (q_15__2), .QB (\$dummy [59]), .D (nx2383)
         , .CLK (nx7076), .R (reset)) ;
    mux21_ni ix2384 (.Y (nx2383), .A0 (q_15__2), .A1 (q_14__2), .S0 (nx6958)) ;
    dffr gen_regs_14_regi_reg_q_2 (.Q (q_14__2), .QB (\$dummy [60]), .D (nx2373)
         , .CLK (nx7076), .R (reset)) ;
    mux21_ni ix2374 (.Y (nx2373), .A0 (q_14__2), .A1 (q_13__2), .S0 (nx6958)) ;
    dffr gen_regs_13_regi_reg_q_2 (.Q (q_13__2), .QB (\$dummy [61]), .D (nx2363)
         , .CLK (nx7076), .R (reset)) ;
    mux21_ni ix2364 (.Y (nx2363), .A0 (q_13__2), .A1 (q_12__2), .S0 (nx6958)) ;
    dffr gen_regs_12_regi_reg_q_2 (.Q (q_12__2), .QB (\$dummy [62]), .D (nx2353)
         , .CLK (nx7074), .R (reset)) ;
    mux21_ni ix2354 (.Y (nx2353), .A0 (q_12__2), .A1 (q_11__2), .S0 (nx6956)) ;
    dffr gen_regs_11_regi_reg_q_2 (.Q (q_11__2), .QB (\$dummy [63]), .D (nx2343)
         , .CLK (nx7074), .R (reset)) ;
    mux21_ni ix2344 (.Y (nx2343), .A0 (q_11__2), .A1 (q_10__2), .S0 (nx6956)) ;
    dffr gen_regs_10_regi_reg_q_2 (.Q (q_10__2), .QB (\$dummy [64]), .D (nx2333)
         , .CLK (nx7074), .R (reset)) ;
    mux21_ni ix2334 (.Y (nx2333), .A0 (q_10__2), .A1 (q_9__2), .S0 (nx6956)) ;
    dffr gen_regs_9_regi_reg_q_2 (.Q (q_9__2), .QB (\$dummy [65]), .D (nx2323), 
         .CLK (nx7074), .R (reset)) ;
    mux21_ni ix2324 (.Y (nx2323), .A0 (q_9__2), .A1 (q_8__2), .S0 (nx6956)) ;
    dffr gen_regs_8_regi_reg_q_2 (.Q (q_8__2), .QB (\$dummy [66]), .D (nx2313), 
         .CLK (nx7074), .R (reset)) ;
    mux21_ni ix2314 (.Y (nx2313), .A0 (q_8__2), .A1 (q_7__2), .S0 (nx6956)) ;
    dffr gen_regs_7_regi_reg_q_2 (.Q (q_7__2), .QB (\$dummy [67]), .D (nx2303), 
         .CLK (nx7074), .R (reset)) ;
    mux21_ni ix2304 (.Y (nx2303), .A0 (q_7__2), .A1 (q_6__2), .S0 (nx6956)) ;
    dffr gen_regs_6_regi_reg_q_2 (.Q (q_6__2), .QB (\$dummy [68]), .D (nx2293), 
         .CLK (nx7074), .R (reset)) ;
    mux21_ni ix2294 (.Y (nx2293), .A0 (q_6__2), .A1 (q_5__2), .S0 (nx6956)) ;
    dffr gen_regs_5_regi_reg_q_2 (.Q (q_5__2), .QB (\$dummy [69]), .D (nx2283), 
         .CLK (nx7072), .R (reset)) ;
    mux21_ni ix2284 (.Y (nx2283), .A0 (q_5__2), .A1 (q_4__2), .S0 (nx6954)) ;
    dffr gen_regs_4_regi_reg_q_2 (.Q (q_4__2), .QB (\$dummy [70]), .D (nx2273), 
         .CLK (nx7072), .R (reset)) ;
    mux21_ni ix2274 (.Y (nx2273), .A0 (q_4__2), .A1 (q_3__2), .S0 (nx6954)) ;
    dffr gen_regs_3_regi_reg_q_2 (.Q (q_3__2), .QB (\$dummy [71]), .D (nx2263), 
         .CLK (nx7072), .R (reset)) ;
    mux21_ni ix2264 (.Y (nx2263), .A0 (q_3__2), .A1 (q_2__2), .S0 (nx6954)) ;
    dffr gen_regs_2_regi_reg_q_2 (.Q (q_2__2), .QB (\$dummy [72]), .D (nx2253), 
         .CLK (nx7072), .R (reset)) ;
    mux21_ni ix2254 (.Y (nx2253), .A0 (q_2__2), .A1 (q_1__2), .S0 (nx6954)) ;
    dffr gen_regs_1_regi_reg_q_2 (.Q (q_1__2), .QB (\$dummy [73]), .D (nx2243), 
         .CLK (nx7072), .R (reset)) ;
    mux21_ni ix2244 (.Y (nx2243), .A0 (q_1__2), .A1 (q_0__2), .S0 (nx6954)) ;
    dffr reg0_reg_q_2 (.Q (q_0__2), .QB (\$dummy [74]), .D (nx2233), .CLK (
         nx7072), .R (reset)) ;
    mux21_ni ix2234 (.Y (nx2233), .A0 (q_0__2), .A1 (d[2]), .S0 (nx6954)) ;
    dffr gen_regs_24_regi_reg_q_3 (.Q (q_24__3), .QB (\$dummy [75]), .D (nx2723)
         , .CLK (nx7086), .R (reset)) ;
    mux21_ni ix2724 (.Y (nx2723), .A0 (q_24__3), .A1 (q_23__3), .S0 (nx6968)) ;
    dffr gen_regs_23_regi_reg_q_3 (.Q (q_23__3), .QB (\$dummy [76]), .D (nx2713)
         , .CLK (nx7086), .R (reset)) ;
    mux21_ni ix2714 (.Y (nx2713), .A0 (q_23__3), .A1 (q_22__3), .S0 (nx6968)) ;
    dffr gen_regs_22_regi_reg_q_3 (.Q (q_22__3), .QB (\$dummy [77]), .D (nx2703)
         , .CLK (nx7084), .R (reset)) ;
    mux21_ni ix2704 (.Y (nx2703), .A0 (q_22__3), .A1 (q_21__3), .S0 (nx6966)) ;
    dffr gen_regs_21_regi_reg_q_3 (.Q (q_21__3), .QB (\$dummy [78]), .D (nx2693)
         , .CLK (nx7084), .R (reset)) ;
    mux21_ni ix2694 (.Y (nx2693), .A0 (q_21__3), .A1 (q_20__3), .S0 (nx6966)) ;
    dffr gen_regs_20_regi_reg_q_3 (.Q (q_20__3), .QB (\$dummy [79]), .D (nx2683)
         , .CLK (nx7084), .R (reset)) ;
    mux21_ni ix2684 (.Y (nx2683), .A0 (q_20__3), .A1 (q_19__3), .S0 (nx6966)) ;
    dffr gen_regs_19_regi_reg_q_3 (.Q (q_19__3), .QB (\$dummy [80]), .D (nx2673)
         , .CLK (nx7084), .R (reset)) ;
    mux21_ni ix2674 (.Y (nx2673), .A0 (q_19__3), .A1 (q_18__3), .S0 (nx6966)) ;
    dffr gen_regs_18_regi_reg_q_3 (.Q (q_18__3), .QB (\$dummy [81]), .D (nx2663)
         , .CLK (nx7084), .R (reset)) ;
    mux21_ni ix2664 (.Y (nx2663), .A0 (q_18__3), .A1 (q_17__3), .S0 (nx6966)) ;
    dffr gen_regs_17_regi_reg_q_3 (.Q (q_17__3), .QB (\$dummy [82]), .D (nx2653)
         , .CLK (nx7084), .R (reset)) ;
    mux21_ni ix2654 (.Y (nx2653), .A0 (q_17__3), .A1 (q_16__3), .S0 (nx6966)) ;
    dffr gen_regs_16_regi_reg_q_3 (.Q (q_16__3), .QB (\$dummy [83]), .D (nx2643)
         , .CLK (nx7084), .R (reset)) ;
    mux21_ni ix2644 (.Y (nx2643), .A0 (q_16__3), .A1 (q_15__3), .S0 (nx6966)) ;
    dffr gen_regs_15_regi_reg_q_3 (.Q (q_15__3), .QB (\$dummy [84]), .D (nx2633)
         , .CLK (nx7082), .R (reset)) ;
    mux21_ni ix2634 (.Y (nx2633), .A0 (q_15__3), .A1 (q_14__3), .S0 (nx6964)) ;
    dffr gen_regs_14_regi_reg_q_3 (.Q (q_14__3), .QB (\$dummy [85]), .D (nx2623)
         , .CLK (nx7082), .R (reset)) ;
    mux21_ni ix2624 (.Y (nx2623), .A0 (q_14__3), .A1 (q_13__3), .S0 (nx6964)) ;
    dffr gen_regs_13_regi_reg_q_3 (.Q (q_13__3), .QB (\$dummy [86]), .D (nx2613)
         , .CLK (nx7082), .R (reset)) ;
    mux21_ni ix2614 (.Y (nx2613), .A0 (q_13__3), .A1 (q_12__3), .S0 (nx6964)) ;
    dffr gen_regs_12_regi_reg_q_3 (.Q (q_12__3), .QB (\$dummy [87]), .D (nx2603)
         , .CLK (nx7082), .R (reset)) ;
    mux21_ni ix2604 (.Y (nx2603), .A0 (q_12__3), .A1 (q_11__3), .S0 (nx6964)) ;
    dffr gen_regs_11_regi_reg_q_3 (.Q (q_11__3), .QB (\$dummy [88]), .D (nx2593)
         , .CLK (nx7082), .R (reset)) ;
    mux21_ni ix2594 (.Y (nx2593), .A0 (q_11__3), .A1 (q_10__3), .S0 (nx6964)) ;
    dffr gen_regs_10_regi_reg_q_3 (.Q (q_10__3), .QB (\$dummy [89]), .D (nx2583)
         , .CLK (nx7082), .R (reset)) ;
    mux21_ni ix2584 (.Y (nx2583), .A0 (q_10__3), .A1 (q_9__3), .S0 (nx6964)) ;
    dffr gen_regs_9_regi_reg_q_3 (.Q (q_9__3), .QB (\$dummy [90]), .D (nx2573), 
         .CLK (nx7082), .R (reset)) ;
    mux21_ni ix2574 (.Y (nx2573), .A0 (q_9__3), .A1 (q_8__3), .S0 (nx6964)) ;
    dffr gen_regs_8_regi_reg_q_3 (.Q (q_8__3), .QB (\$dummy [91]), .D (nx2563), 
         .CLK (nx7080), .R (reset)) ;
    mux21_ni ix2564 (.Y (nx2563), .A0 (q_8__3), .A1 (q_7__3), .S0 (nx6962)) ;
    dffr gen_regs_7_regi_reg_q_3 (.Q (q_7__3), .QB (\$dummy [92]), .D (nx2553), 
         .CLK (nx7080), .R (reset)) ;
    mux21_ni ix2554 (.Y (nx2553), .A0 (q_7__3), .A1 (q_6__3), .S0 (nx6962)) ;
    dffr gen_regs_6_regi_reg_q_3 (.Q (q_6__3), .QB (\$dummy [93]), .D (nx2543), 
         .CLK (nx7080), .R (reset)) ;
    mux21_ni ix2544 (.Y (nx2543), .A0 (q_6__3), .A1 (q_5__3), .S0 (nx6962)) ;
    dffr gen_regs_5_regi_reg_q_3 (.Q (q_5__3), .QB (\$dummy [94]), .D (nx2533), 
         .CLK (nx7080), .R (reset)) ;
    mux21_ni ix2534 (.Y (nx2533), .A0 (q_5__3), .A1 (q_4__3), .S0 (nx6962)) ;
    dffr gen_regs_4_regi_reg_q_3 (.Q (q_4__3), .QB (\$dummy [95]), .D (nx2523), 
         .CLK (nx7080), .R (reset)) ;
    mux21_ni ix2524 (.Y (nx2523), .A0 (q_4__3), .A1 (q_3__3), .S0 (nx6962)) ;
    dffr gen_regs_3_regi_reg_q_3 (.Q (q_3__3), .QB (\$dummy [96]), .D (nx2513), 
         .CLK (nx7080), .R (reset)) ;
    mux21_ni ix2514 (.Y (nx2513), .A0 (q_3__3), .A1 (q_2__3), .S0 (nx6962)) ;
    dffr gen_regs_2_regi_reg_q_3 (.Q (q_2__3), .QB (\$dummy [97]), .D (nx2503), 
         .CLK (nx7080), .R (reset)) ;
    mux21_ni ix2504 (.Y (nx2503), .A0 (q_2__3), .A1 (q_1__3), .S0 (nx6962)) ;
    dffr gen_regs_1_regi_reg_q_3 (.Q (q_1__3), .QB (\$dummy [98]), .D (nx2493), 
         .CLK (nx7078), .R (reset)) ;
    mux21_ni ix2494 (.Y (nx2493), .A0 (q_1__3), .A1 (q_0__3), .S0 (nx6960)) ;
    dffr reg0_reg_q_3 (.Q (q_0__3), .QB (\$dummy [99]), .D (nx2483), .CLK (
         nx7078), .R (reset)) ;
    mux21_ni ix2484 (.Y (nx2483), .A0 (q_0__3), .A1 (d[3]), .S0 (nx6960)) ;
    dffr gen_regs_24_regi_reg_q_4 (.Q (q_24__4), .QB (\$dummy [100]), .D (nx2973
         ), .CLK (nx7092), .R (reset)) ;
    mux21_ni ix2974 (.Y (nx2973), .A0 (q_24__4), .A1 (q_23__4), .S0 (nx6974)) ;
    dffr gen_regs_23_regi_reg_q_4 (.Q (q_23__4), .QB (\$dummy [101]), .D (nx2963
         ), .CLK (nx7092), .R (reset)) ;
    mux21_ni ix2964 (.Y (nx2963), .A0 (q_23__4), .A1 (q_22__4), .S0 (nx6974)) ;
    dffr gen_regs_22_regi_reg_q_4 (.Q (q_22__4), .QB (\$dummy [102]), .D (nx2953
         ), .CLK (nx7092), .R (reset)) ;
    mux21_ni ix2954 (.Y (nx2953), .A0 (q_22__4), .A1 (q_21__4), .S0 (nx6974)) ;
    dffr gen_regs_21_regi_reg_q_4 (.Q (q_21__4), .QB (\$dummy [103]), .D (nx2943
         ), .CLK (nx7092), .R (reset)) ;
    mux21_ni ix2944 (.Y (nx2943), .A0 (q_21__4), .A1 (q_20__4), .S0 (nx6974)) ;
    dffr gen_regs_20_regi_reg_q_4 (.Q (q_20__4), .QB (\$dummy [104]), .D (nx2933
         ), .CLK (nx7092), .R (reset)) ;
    mux21_ni ix2934 (.Y (nx2933), .A0 (q_20__4), .A1 (q_19__4), .S0 (nx6974)) ;
    dffr gen_regs_19_regi_reg_q_4 (.Q (q_19__4), .QB (\$dummy [105]), .D (nx2923
         ), .CLK (nx7092), .R (reset)) ;
    mux21_ni ix2924 (.Y (nx2923), .A0 (q_19__4), .A1 (q_18__4), .S0 (nx6974)) ;
    dffr gen_regs_18_regi_reg_q_4 (.Q (q_18__4), .QB (\$dummy [106]), .D (nx2913
         ), .CLK (nx7090), .R (reset)) ;
    mux21_ni ix2914 (.Y (nx2913), .A0 (q_18__4), .A1 (q_17__4), .S0 (nx6972)) ;
    dffr gen_regs_17_regi_reg_q_4 (.Q (q_17__4), .QB (\$dummy [107]), .D (nx2903
         ), .CLK (nx7090), .R (reset)) ;
    mux21_ni ix2904 (.Y (nx2903), .A0 (q_17__4), .A1 (q_16__4), .S0 (nx6972)) ;
    dffr gen_regs_16_regi_reg_q_4 (.Q (q_16__4), .QB (\$dummy [108]), .D (nx2893
         ), .CLK (nx7090), .R (reset)) ;
    mux21_ni ix2894 (.Y (nx2893), .A0 (q_16__4), .A1 (q_15__4), .S0 (nx6972)) ;
    dffr gen_regs_15_regi_reg_q_4 (.Q (q_15__4), .QB (\$dummy [109]), .D (nx2883
         ), .CLK (nx7090), .R (reset)) ;
    mux21_ni ix2884 (.Y (nx2883), .A0 (q_15__4), .A1 (q_14__4), .S0 (nx6972)) ;
    dffr gen_regs_14_regi_reg_q_4 (.Q (q_14__4), .QB (\$dummy [110]), .D (nx2873
         ), .CLK (nx7090), .R (reset)) ;
    mux21_ni ix2874 (.Y (nx2873), .A0 (q_14__4), .A1 (q_13__4), .S0 (nx6972)) ;
    dffr gen_regs_13_regi_reg_q_4 (.Q (q_13__4), .QB (\$dummy [111]), .D (nx2863
         ), .CLK (nx7090), .R (reset)) ;
    mux21_ni ix2864 (.Y (nx2863), .A0 (q_13__4), .A1 (q_12__4), .S0 (nx6972)) ;
    dffr gen_regs_12_regi_reg_q_4 (.Q (q_12__4), .QB (\$dummy [112]), .D (nx2853
         ), .CLK (nx7090), .R (reset)) ;
    mux21_ni ix2854 (.Y (nx2853), .A0 (q_12__4), .A1 (q_11__4), .S0 (nx6972)) ;
    dffr gen_regs_11_regi_reg_q_4 (.Q (q_11__4), .QB (\$dummy [113]), .D (nx2843
         ), .CLK (nx7088), .R (reset)) ;
    mux21_ni ix2844 (.Y (nx2843), .A0 (q_11__4), .A1 (q_10__4), .S0 (nx6970)) ;
    dffr gen_regs_10_regi_reg_q_4 (.Q (q_10__4), .QB (\$dummy [114]), .D (nx2833
         ), .CLK (nx7088), .R (reset)) ;
    mux21_ni ix2834 (.Y (nx2833), .A0 (q_10__4), .A1 (q_9__4), .S0 (nx6970)) ;
    dffr gen_regs_9_regi_reg_q_4 (.Q (q_9__4), .QB (\$dummy [115]), .D (nx2823)
         , .CLK (nx7088), .R (reset)) ;
    mux21_ni ix2824 (.Y (nx2823), .A0 (q_9__4), .A1 (q_8__4), .S0 (nx6970)) ;
    dffr gen_regs_8_regi_reg_q_4 (.Q (q_8__4), .QB (\$dummy [116]), .D (nx2813)
         , .CLK (nx7088), .R (reset)) ;
    mux21_ni ix2814 (.Y (nx2813), .A0 (q_8__4), .A1 (q_7__4), .S0 (nx6970)) ;
    dffr gen_regs_7_regi_reg_q_4 (.Q (q_7__4), .QB (\$dummy [117]), .D (nx2803)
         , .CLK (nx7088), .R (reset)) ;
    mux21_ni ix2804 (.Y (nx2803), .A0 (q_7__4), .A1 (q_6__4), .S0 (nx6970)) ;
    dffr gen_regs_6_regi_reg_q_4 (.Q (q_6__4), .QB (\$dummy [118]), .D (nx2793)
         , .CLK (nx7088), .R (reset)) ;
    mux21_ni ix2794 (.Y (nx2793), .A0 (q_6__4), .A1 (q_5__4), .S0 (nx6970)) ;
    dffr gen_regs_5_regi_reg_q_4 (.Q (q_5__4), .QB (\$dummy [119]), .D (nx2783)
         , .CLK (nx7088), .R (reset)) ;
    mux21_ni ix2784 (.Y (nx2783), .A0 (q_5__4), .A1 (q_4__4), .S0 (nx6970)) ;
    dffr gen_regs_4_regi_reg_q_4 (.Q (q_4__4), .QB (\$dummy [120]), .D (nx2773)
         , .CLK (nx7086), .R (reset)) ;
    mux21_ni ix2774 (.Y (nx2773), .A0 (q_4__4), .A1 (q_3__4), .S0 (nx6968)) ;
    dffr gen_regs_3_regi_reg_q_4 (.Q (q_3__4), .QB (\$dummy [121]), .D (nx2763)
         , .CLK (nx7086), .R (reset)) ;
    mux21_ni ix2764 (.Y (nx2763), .A0 (q_3__4), .A1 (q_2__4), .S0 (nx6968)) ;
    dffr gen_regs_2_regi_reg_q_4 (.Q (q_2__4), .QB (\$dummy [122]), .D (nx2753)
         , .CLK (nx7086), .R (reset)) ;
    mux21_ni ix2754 (.Y (nx2753), .A0 (q_2__4), .A1 (q_1__4), .S0 (nx6968)) ;
    dffr gen_regs_1_regi_reg_q_4 (.Q (q_1__4), .QB (\$dummy [123]), .D (nx2743)
         , .CLK (nx7086), .R (reset)) ;
    mux21_ni ix2744 (.Y (nx2743), .A0 (q_1__4), .A1 (q_0__4), .S0 (nx6968)) ;
    dffr reg0_reg_q_4 (.Q (q_0__4), .QB (\$dummy [124]), .D (nx2733), .CLK (
         nx7086), .R (reset)) ;
    mux21_ni ix2734 (.Y (nx2733), .A0 (q_0__4), .A1 (d[4]), .S0 (nx6968)) ;
    dffr gen_regs_24_regi_reg_q_5 (.Q (q_24__5), .QB (\$dummy [125]), .D (nx3223
         ), .CLK (nx7100), .R (reset)) ;
    mux21_ni ix3224 (.Y (nx3223), .A0 (q_24__5), .A1 (q_23__5), .S0 (nx6982)) ;
    dffr gen_regs_23_regi_reg_q_5 (.Q (q_23__5), .QB (\$dummy [126]), .D (nx3213
         ), .CLK (nx7100), .R (reset)) ;
    mux21_ni ix3214 (.Y (nx3213), .A0 (q_23__5), .A1 (q_22__5), .S0 (nx6982)) ;
    dffr gen_regs_22_regi_reg_q_5 (.Q (q_22__5), .QB (\$dummy [127]), .D (nx3203
         ), .CLK (nx7100), .R (reset)) ;
    mux21_ni ix3204 (.Y (nx3203), .A0 (q_22__5), .A1 (q_21__5), .S0 (nx6982)) ;
    dffr gen_regs_21_regi_reg_q_5 (.Q (q_21__5), .QB (\$dummy [128]), .D (nx3193
         ), .CLK (nx7098), .R (reset)) ;
    mux21_ni ix3194 (.Y (nx3193), .A0 (q_21__5), .A1 (q_20__5), .S0 (nx6980)) ;
    dffr gen_regs_20_regi_reg_q_5 (.Q (q_20__5), .QB (\$dummy [129]), .D (nx3183
         ), .CLK (nx7098), .R (reset)) ;
    mux21_ni ix3184 (.Y (nx3183), .A0 (q_20__5), .A1 (q_19__5), .S0 (nx6980)) ;
    dffr gen_regs_19_regi_reg_q_5 (.Q (q_19__5), .QB (\$dummy [130]), .D (nx3173
         ), .CLK (nx7098), .R (reset)) ;
    mux21_ni ix3174 (.Y (nx3173), .A0 (q_19__5), .A1 (q_18__5), .S0 (nx6980)) ;
    dffr gen_regs_18_regi_reg_q_5 (.Q (q_18__5), .QB (\$dummy [131]), .D (nx3163
         ), .CLK (nx7098), .R (reset)) ;
    mux21_ni ix3164 (.Y (nx3163), .A0 (q_18__5), .A1 (q_17__5), .S0 (nx6980)) ;
    dffr gen_regs_17_regi_reg_q_5 (.Q (q_17__5), .QB (\$dummy [132]), .D (nx3153
         ), .CLK (nx7098), .R (reset)) ;
    mux21_ni ix3154 (.Y (nx3153), .A0 (q_17__5), .A1 (q_16__5), .S0 (nx6980)) ;
    dffr gen_regs_16_regi_reg_q_5 (.Q (q_16__5), .QB (\$dummy [133]), .D (nx3143
         ), .CLK (nx7098), .R (reset)) ;
    mux21_ni ix3144 (.Y (nx3143), .A0 (q_16__5), .A1 (q_15__5), .S0 (nx6980)) ;
    dffr gen_regs_15_regi_reg_q_5 (.Q (q_15__5), .QB (\$dummy [134]), .D (nx3133
         ), .CLK (nx7098), .R (reset)) ;
    mux21_ni ix3134 (.Y (nx3133), .A0 (q_15__5), .A1 (q_14__5), .S0 (nx6980)) ;
    dffr gen_regs_14_regi_reg_q_5 (.Q (q_14__5), .QB (\$dummy [135]), .D (nx3123
         ), .CLK (nx7096), .R (reset)) ;
    mux21_ni ix3124 (.Y (nx3123), .A0 (q_14__5), .A1 (q_13__5), .S0 (nx6978)) ;
    dffr gen_regs_13_regi_reg_q_5 (.Q (q_13__5), .QB (\$dummy [136]), .D (nx3113
         ), .CLK (nx7096), .R (reset)) ;
    mux21_ni ix3114 (.Y (nx3113), .A0 (q_13__5), .A1 (q_12__5), .S0 (nx6978)) ;
    dffr gen_regs_12_regi_reg_q_5 (.Q (q_12__5), .QB (\$dummy [137]), .D (nx3103
         ), .CLK (nx7096), .R (reset)) ;
    mux21_ni ix3104 (.Y (nx3103), .A0 (q_12__5), .A1 (q_11__5), .S0 (nx6978)) ;
    dffr gen_regs_11_regi_reg_q_5 (.Q (q_11__5), .QB (\$dummy [138]), .D (nx3093
         ), .CLK (nx7096), .R (reset)) ;
    mux21_ni ix3094 (.Y (nx3093), .A0 (q_11__5), .A1 (q_10__5), .S0 (nx6978)) ;
    dffr gen_regs_10_regi_reg_q_5 (.Q (q_10__5), .QB (\$dummy [139]), .D (nx3083
         ), .CLK (nx7096), .R (reset)) ;
    mux21_ni ix3084 (.Y (nx3083), .A0 (q_10__5), .A1 (q_9__5), .S0 (nx6978)) ;
    dffr gen_regs_9_regi_reg_q_5 (.Q (q_9__5), .QB (\$dummy [140]), .D (nx3073)
         , .CLK (nx7096), .R (reset)) ;
    mux21_ni ix3074 (.Y (nx3073), .A0 (q_9__5), .A1 (q_8__5), .S0 (nx6978)) ;
    dffr gen_regs_8_regi_reg_q_5 (.Q (q_8__5), .QB (\$dummy [141]), .D (nx3063)
         , .CLK (nx7096), .R (reset)) ;
    mux21_ni ix3064 (.Y (nx3063), .A0 (q_8__5), .A1 (q_7__5), .S0 (nx6978)) ;
    dffr gen_regs_7_regi_reg_q_5 (.Q (q_7__5), .QB (\$dummy [142]), .D (nx3053)
         , .CLK (nx7094), .R (reset)) ;
    mux21_ni ix3054 (.Y (nx3053), .A0 (q_7__5), .A1 (q_6__5), .S0 (nx6976)) ;
    dffr gen_regs_6_regi_reg_q_5 (.Q (q_6__5), .QB (\$dummy [143]), .D (nx3043)
         , .CLK (nx7094), .R (reset)) ;
    mux21_ni ix3044 (.Y (nx3043), .A0 (q_6__5), .A1 (q_5__5), .S0 (nx6976)) ;
    dffr gen_regs_5_regi_reg_q_5 (.Q (q_5__5), .QB (\$dummy [144]), .D (nx3033)
         , .CLK (nx7094), .R (reset)) ;
    mux21_ni ix3034 (.Y (nx3033), .A0 (q_5__5), .A1 (q_4__5), .S0 (nx6976)) ;
    dffr gen_regs_4_regi_reg_q_5 (.Q (q_4__5), .QB (\$dummy [145]), .D (nx3023)
         , .CLK (nx7094), .R (reset)) ;
    mux21_ni ix3024 (.Y (nx3023), .A0 (q_4__5), .A1 (q_3__5), .S0 (nx6976)) ;
    dffr gen_regs_3_regi_reg_q_5 (.Q (q_3__5), .QB (\$dummy [146]), .D (nx3013)
         , .CLK (nx7094), .R (reset)) ;
    mux21_ni ix3014 (.Y (nx3013), .A0 (q_3__5), .A1 (q_2__5), .S0 (nx6976)) ;
    dffr gen_regs_2_regi_reg_q_5 (.Q (q_2__5), .QB (\$dummy [147]), .D (nx3003)
         , .CLK (nx7094), .R (reset)) ;
    mux21_ni ix3004 (.Y (nx3003), .A0 (q_2__5), .A1 (q_1__5), .S0 (nx6976)) ;
    dffr gen_regs_1_regi_reg_q_5 (.Q (q_1__5), .QB (\$dummy [148]), .D (nx2993)
         , .CLK (nx7094), .R (reset)) ;
    mux21_ni ix2994 (.Y (nx2993), .A0 (q_1__5), .A1 (q_0__5), .S0 (nx6976)) ;
    dffr reg0_reg_q_5 (.Q (q_0__5), .QB (\$dummy [149]), .D (nx2983), .CLK (
         nx7092), .R (reset)) ;
    mux21_ni ix2984 (.Y (nx2983), .A0 (q_0__5), .A1 (d[5]), .S0 (nx6974)) ;
    dffr gen_regs_24_regi_reg_q_6 (.Q (q_24__6), .QB (\$dummy [150]), .D (nx3473
         ), .CLK (nx7106), .R (reset)) ;
    mux21_ni ix3474 (.Y (nx3473), .A0 (q_24__6), .A1 (q_23__6), .S0 (nx6988)) ;
    dffr gen_regs_23_regi_reg_q_6 (.Q (q_23__6), .QB (\$dummy [151]), .D (nx3463
         ), .CLK (nx7106), .R (reset)) ;
    mux21_ni ix3464 (.Y (nx3463), .A0 (q_23__6), .A1 (q_22__6), .S0 (nx6988)) ;
    dffr gen_regs_22_regi_reg_q_6 (.Q (q_22__6), .QB (\$dummy [152]), .D (nx3453
         ), .CLK (nx7106), .R (reset)) ;
    mux21_ni ix3454 (.Y (nx3453), .A0 (q_22__6), .A1 (q_21__6), .S0 (nx6988)) ;
    dffr gen_regs_21_regi_reg_q_6 (.Q (q_21__6), .QB (\$dummy [153]), .D (nx3443
         ), .CLK (nx7106), .R (reset)) ;
    mux21_ni ix3444 (.Y (nx3443), .A0 (q_21__6), .A1 (q_20__6), .S0 (nx6988)) ;
    dffr gen_regs_20_regi_reg_q_6 (.Q (q_20__6), .QB (\$dummy [154]), .D (nx3433
         ), .CLK (nx7106), .R (reset)) ;
    mux21_ni ix3434 (.Y (nx3433), .A0 (q_20__6), .A1 (q_19__6), .S0 (nx6988)) ;
    dffr gen_regs_19_regi_reg_q_6 (.Q (q_19__6), .QB (\$dummy [155]), .D (nx3423
         ), .CLK (nx7106), .R (reset)) ;
    mux21_ni ix3424 (.Y (nx3423), .A0 (q_19__6), .A1 (q_18__6), .S0 (nx6988)) ;
    dffr gen_regs_18_regi_reg_q_6 (.Q (q_18__6), .QB (\$dummy [156]), .D (nx3413
         ), .CLK (nx7106), .R (reset)) ;
    mux21_ni ix3414 (.Y (nx3413), .A0 (q_18__6), .A1 (q_17__6), .S0 (nx6988)) ;
    dffr gen_regs_17_regi_reg_q_6 (.Q (q_17__6), .QB (\$dummy [157]), .D (nx3403
         ), .CLK (nx7104), .R (reset)) ;
    mux21_ni ix3404 (.Y (nx3403), .A0 (q_17__6), .A1 (q_16__6), .S0 (nx6986)) ;
    dffr gen_regs_16_regi_reg_q_6 (.Q (q_16__6), .QB (\$dummy [158]), .D (nx3393
         ), .CLK (nx7104), .R (reset)) ;
    mux21_ni ix3394 (.Y (nx3393), .A0 (q_16__6), .A1 (q_15__6), .S0 (nx6986)) ;
    dffr gen_regs_15_regi_reg_q_6 (.Q (q_15__6), .QB (\$dummy [159]), .D (nx3383
         ), .CLK (nx7104), .R (reset)) ;
    mux21_ni ix3384 (.Y (nx3383), .A0 (q_15__6), .A1 (q_14__6), .S0 (nx6986)) ;
    dffr gen_regs_14_regi_reg_q_6 (.Q (q_14__6), .QB (\$dummy [160]), .D (nx3373
         ), .CLK (nx7104), .R (reset)) ;
    mux21_ni ix3374 (.Y (nx3373), .A0 (q_14__6), .A1 (q_13__6), .S0 (nx6986)) ;
    dffr gen_regs_13_regi_reg_q_6 (.Q (q_13__6), .QB (\$dummy [161]), .D (nx3363
         ), .CLK (nx7104), .R (reset)) ;
    mux21_ni ix3364 (.Y (nx3363), .A0 (q_13__6), .A1 (q_12__6), .S0 (nx6986)) ;
    dffr gen_regs_12_regi_reg_q_6 (.Q (q_12__6), .QB (\$dummy [162]), .D (nx3353
         ), .CLK (nx7104), .R (reset)) ;
    mux21_ni ix3354 (.Y (nx3353), .A0 (q_12__6), .A1 (q_11__6), .S0 (nx6986)) ;
    dffr gen_regs_11_regi_reg_q_6 (.Q (q_11__6), .QB (\$dummy [163]), .D (nx3343
         ), .CLK (nx7104), .R (reset)) ;
    mux21_ni ix3344 (.Y (nx3343), .A0 (q_11__6), .A1 (q_10__6), .S0 (nx6986)) ;
    dffr gen_regs_10_regi_reg_q_6 (.Q (q_10__6), .QB (\$dummy [164]), .D (nx3333
         ), .CLK (nx7102), .R (reset)) ;
    mux21_ni ix3334 (.Y (nx3333), .A0 (q_10__6), .A1 (q_9__6), .S0 (nx6984)) ;
    dffr gen_regs_9_regi_reg_q_6 (.Q (q_9__6), .QB (\$dummy [165]), .D (nx3323)
         , .CLK (nx7102), .R (reset)) ;
    mux21_ni ix3324 (.Y (nx3323), .A0 (q_9__6), .A1 (q_8__6), .S0 (nx6984)) ;
    dffr gen_regs_8_regi_reg_q_6 (.Q (q_8__6), .QB (\$dummy [166]), .D (nx3313)
         , .CLK (nx7102), .R (reset)) ;
    mux21_ni ix3314 (.Y (nx3313), .A0 (q_8__6), .A1 (q_7__6), .S0 (nx6984)) ;
    dffr gen_regs_7_regi_reg_q_6 (.Q (q_7__6), .QB (\$dummy [167]), .D (nx3303)
         , .CLK (nx7102), .R (reset)) ;
    mux21_ni ix3304 (.Y (nx3303), .A0 (q_7__6), .A1 (q_6__6), .S0 (nx6984)) ;
    dffr gen_regs_6_regi_reg_q_6 (.Q (q_6__6), .QB (\$dummy [168]), .D (nx3293)
         , .CLK (nx7102), .R (reset)) ;
    mux21_ni ix3294 (.Y (nx3293), .A0 (q_6__6), .A1 (q_5__6), .S0 (nx6984)) ;
    dffr gen_regs_5_regi_reg_q_6 (.Q (q_5__6), .QB (\$dummy [169]), .D (nx3283)
         , .CLK (nx7102), .R (reset)) ;
    mux21_ni ix3284 (.Y (nx3283), .A0 (q_5__6), .A1 (q_4__6), .S0 (nx6984)) ;
    dffr gen_regs_4_regi_reg_q_6 (.Q (q_4__6), .QB (\$dummy [170]), .D (nx3273)
         , .CLK (nx7102), .R (reset)) ;
    mux21_ni ix3274 (.Y (nx3273), .A0 (q_4__6), .A1 (q_3__6), .S0 (nx6984)) ;
    dffr gen_regs_3_regi_reg_q_6 (.Q (q_3__6), .QB (\$dummy [171]), .D (nx3263)
         , .CLK (nx7100), .R (reset)) ;
    mux21_ni ix3264 (.Y (nx3263), .A0 (q_3__6), .A1 (q_2__6), .S0 (nx6982)) ;
    dffr gen_regs_2_regi_reg_q_6 (.Q (q_2__6), .QB (\$dummy [172]), .D (nx3253)
         , .CLK (nx7100), .R (reset)) ;
    mux21_ni ix3254 (.Y (nx3253), .A0 (q_2__6), .A1 (q_1__6), .S0 (nx6982)) ;
    dffr gen_regs_1_regi_reg_q_6 (.Q (q_1__6), .QB (\$dummy [173]), .D (nx3243)
         , .CLK (nx7100), .R (reset)) ;
    mux21_ni ix3244 (.Y (nx3243), .A0 (q_1__6), .A1 (q_0__6), .S0 (nx6982)) ;
    dffr reg0_reg_q_6 (.Q (q_0__6), .QB (\$dummy [174]), .D (nx3233), .CLK (
         nx7100), .R (reset)) ;
    mux21_ni ix3234 (.Y (nx3233), .A0 (q_0__6), .A1 (d[6]), .S0 (nx6982)) ;
    dffr gen_regs_24_regi_reg_q_7 (.Q (q_24__7), .QB (\$dummy [175]), .D (nx3723
         ), .CLK (nx7114), .R (reset)) ;
    mux21_ni ix3724 (.Y (nx3723), .A0 (q_24__7), .A1 (q_23__7), .S0 (nx6996)) ;
    dffr gen_regs_23_regi_reg_q_7 (.Q (q_23__7), .QB (\$dummy [176]), .D (nx3713
         ), .CLK (nx7114), .R (reset)) ;
    mux21_ni ix3714 (.Y (nx3713), .A0 (q_23__7), .A1 (q_22__7), .S0 (nx6996)) ;
    dffr gen_regs_22_regi_reg_q_7 (.Q (q_22__7), .QB (\$dummy [177]), .D (nx3703
         ), .CLK (nx7114), .R (reset)) ;
    mux21_ni ix3704 (.Y (nx3703), .A0 (q_22__7), .A1 (q_21__7), .S0 (nx6996)) ;
    dffr gen_regs_21_regi_reg_q_7 (.Q (q_21__7), .QB (\$dummy [178]), .D (nx3693
         ), .CLK (nx7114), .R (reset)) ;
    mux21_ni ix3694 (.Y (nx3693), .A0 (q_21__7), .A1 (q_20__7), .S0 (nx6996)) ;
    dffr gen_regs_20_regi_reg_q_7 (.Q (q_20__7), .QB (\$dummy [179]), .D (nx3683
         ), .CLK (nx7112), .R (reset)) ;
    mux21_ni ix3684 (.Y (nx3683), .A0 (q_20__7), .A1 (q_19__7), .S0 (nx6994)) ;
    dffr gen_regs_19_regi_reg_q_7 (.Q (q_19__7), .QB (\$dummy [180]), .D (nx3673
         ), .CLK (nx7112), .R (reset)) ;
    mux21_ni ix3674 (.Y (nx3673), .A0 (q_19__7), .A1 (q_18__7), .S0 (nx6994)) ;
    dffr gen_regs_18_regi_reg_q_7 (.Q (q_18__7), .QB (\$dummy [181]), .D (nx3663
         ), .CLK (nx7112), .R (reset)) ;
    mux21_ni ix3664 (.Y (nx3663), .A0 (q_18__7), .A1 (q_17__7), .S0 (nx6994)) ;
    dffr gen_regs_17_regi_reg_q_7 (.Q (q_17__7), .QB (\$dummy [182]), .D (nx3653
         ), .CLK (nx7112), .R (reset)) ;
    mux21_ni ix3654 (.Y (nx3653), .A0 (q_17__7), .A1 (q_16__7), .S0 (nx6994)) ;
    dffr gen_regs_16_regi_reg_q_7 (.Q (q_16__7), .QB (\$dummy [183]), .D (nx3643
         ), .CLK (nx7112), .R (reset)) ;
    mux21_ni ix3644 (.Y (nx3643), .A0 (q_16__7), .A1 (q_15__7), .S0 (nx6994)) ;
    dffr gen_regs_15_regi_reg_q_7 (.Q (q_15__7), .QB (\$dummy [184]), .D (nx3633
         ), .CLK (nx7112), .R (reset)) ;
    mux21_ni ix3634 (.Y (nx3633), .A0 (q_15__7), .A1 (q_14__7), .S0 (nx6994)) ;
    dffr gen_regs_14_regi_reg_q_7 (.Q (q_14__7), .QB (\$dummy [185]), .D (nx3623
         ), .CLK (nx7112), .R (reset)) ;
    mux21_ni ix3624 (.Y (nx3623), .A0 (q_14__7), .A1 (q_13__7), .S0 (nx6994)) ;
    dffr gen_regs_13_regi_reg_q_7 (.Q (q_13__7), .QB (\$dummy [186]), .D (nx3613
         ), .CLK (nx7110), .R (reset)) ;
    mux21_ni ix3614 (.Y (nx3613), .A0 (q_13__7), .A1 (q_12__7), .S0 (nx6992)) ;
    dffr gen_regs_12_regi_reg_q_7 (.Q (q_12__7), .QB (\$dummy [187]), .D (nx3603
         ), .CLK (nx7110), .R (reset)) ;
    mux21_ni ix3604 (.Y (nx3603), .A0 (q_12__7), .A1 (q_11__7), .S0 (nx6992)) ;
    dffr gen_regs_11_regi_reg_q_7 (.Q (q_11__7), .QB (\$dummy [188]), .D (nx3593
         ), .CLK (nx7110), .R (reset)) ;
    mux21_ni ix3594 (.Y (nx3593), .A0 (q_11__7), .A1 (q_10__7), .S0 (nx6992)) ;
    dffr gen_regs_10_regi_reg_q_7 (.Q (q_10__7), .QB (\$dummy [189]), .D (nx3583
         ), .CLK (nx7110), .R (reset)) ;
    mux21_ni ix3584 (.Y (nx3583), .A0 (q_10__7), .A1 (q_9__7), .S0 (nx6992)) ;
    dffr gen_regs_9_regi_reg_q_7 (.Q (q_9__7), .QB (\$dummy [190]), .D (nx3573)
         , .CLK (nx7110), .R (reset)) ;
    mux21_ni ix3574 (.Y (nx3573), .A0 (q_9__7), .A1 (q_8__7), .S0 (nx6992)) ;
    dffr gen_regs_8_regi_reg_q_7 (.Q (q_8__7), .QB (\$dummy [191]), .D (nx3563)
         , .CLK (nx7110), .R (reset)) ;
    mux21_ni ix3564 (.Y (nx3563), .A0 (q_8__7), .A1 (q_7__7), .S0 (nx6992)) ;
    dffr gen_regs_7_regi_reg_q_7 (.Q (q_7__7), .QB (\$dummy [192]), .D (nx3553)
         , .CLK (nx7110), .R (reset)) ;
    mux21_ni ix3554 (.Y (nx3553), .A0 (q_7__7), .A1 (q_6__7), .S0 (nx6992)) ;
    dffr gen_regs_6_regi_reg_q_7 (.Q (q_6__7), .QB (\$dummy [193]), .D (nx3543)
         , .CLK (nx7108), .R (reset)) ;
    mux21_ni ix3544 (.Y (nx3543), .A0 (q_6__7), .A1 (q_5__7), .S0 (nx6990)) ;
    dffr gen_regs_5_regi_reg_q_7 (.Q (q_5__7), .QB (\$dummy [194]), .D (nx3533)
         , .CLK (nx7108), .R (reset)) ;
    mux21_ni ix3534 (.Y (nx3533), .A0 (q_5__7), .A1 (q_4__7), .S0 (nx6990)) ;
    dffr gen_regs_4_regi_reg_q_7 (.Q (q_4__7), .QB (\$dummy [195]), .D (nx3523)
         , .CLK (nx7108), .R (reset)) ;
    mux21_ni ix3524 (.Y (nx3523), .A0 (q_4__7), .A1 (q_3__7), .S0 (nx6990)) ;
    dffr gen_regs_3_regi_reg_q_7 (.Q (q_3__7), .QB (\$dummy [196]), .D (nx3513)
         , .CLK (nx7108), .R (reset)) ;
    mux21_ni ix3514 (.Y (nx3513), .A0 (q_3__7), .A1 (q_2__7), .S0 (nx6990)) ;
    dffr gen_regs_2_regi_reg_q_7 (.Q (q_2__7), .QB (\$dummy [197]), .D (nx3503)
         , .CLK (nx7108), .R (reset)) ;
    mux21_ni ix3504 (.Y (nx3503), .A0 (q_2__7), .A1 (q_1__7), .S0 (nx6990)) ;
    dffr gen_regs_1_regi_reg_q_7 (.Q (q_1__7), .QB (\$dummy [198]), .D (nx3493)
         , .CLK (nx7108), .R (reset)) ;
    mux21_ni ix3494 (.Y (nx3493), .A0 (q_1__7), .A1 (q_0__7), .S0 (nx6990)) ;
    dffr reg0_reg_q_7 (.Q (q_0__7), .QB (\$dummy [199]), .D (nx3483), .CLK (
         nx7108), .R (reset)) ;
    mux21_ni ix3484 (.Y (nx3483), .A0 (q_0__7), .A1 (d[7]), .S0 (nx6990)) ;
    dffr gen_regs_24_regi_reg_q_8 (.Q (q_24__8), .QB (\$dummy [200]), .D (nx3973
         ), .CLK (nx7122), .R (reset)) ;
    mux21_ni ix3974 (.Y (nx3973), .A0 (q_24__8), .A1 (q_23__8), .S0 (nx7004)) ;
    dffr gen_regs_23_regi_reg_q_8 (.Q (q_23__8), .QB (\$dummy [201]), .D (nx3963
         ), .CLK (nx7120), .R (reset)) ;
    mux21_ni ix3964 (.Y (nx3963), .A0 (q_23__8), .A1 (q_22__8), .S0 (nx7002)) ;
    dffr gen_regs_22_regi_reg_q_8 (.Q (q_22__8), .QB (\$dummy [202]), .D (nx3953
         ), .CLK (nx7120), .R (reset)) ;
    mux21_ni ix3954 (.Y (nx3953), .A0 (q_22__8), .A1 (q_21__8), .S0 (nx7002)) ;
    dffr gen_regs_21_regi_reg_q_8 (.Q (q_21__8), .QB (\$dummy [203]), .D (nx3943
         ), .CLK (nx7120), .R (reset)) ;
    mux21_ni ix3944 (.Y (nx3943), .A0 (q_21__8), .A1 (q_20__8), .S0 (nx7002)) ;
    dffr gen_regs_20_regi_reg_q_8 (.Q (q_20__8), .QB (\$dummy [204]), .D (nx3933
         ), .CLK (nx7120), .R (reset)) ;
    mux21_ni ix3934 (.Y (nx3933), .A0 (q_20__8), .A1 (q_19__8), .S0 (nx7002)) ;
    dffr gen_regs_19_regi_reg_q_8 (.Q (q_19__8), .QB (\$dummy [205]), .D (nx3923
         ), .CLK (nx7120), .R (reset)) ;
    mux21_ni ix3924 (.Y (nx3923), .A0 (q_19__8), .A1 (q_18__8), .S0 (nx7002)) ;
    dffr gen_regs_18_regi_reg_q_8 (.Q (q_18__8), .QB (\$dummy [206]), .D (nx3913
         ), .CLK (nx7120), .R (reset)) ;
    mux21_ni ix3914 (.Y (nx3913), .A0 (q_18__8), .A1 (q_17__8), .S0 (nx7002)) ;
    dffr gen_regs_17_regi_reg_q_8 (.Q (q_17__8), .QB (\$dummy [207]), .D (nx3903
         ), .CLK (nx7120), .R (reset)) ;
    mux21_ni ix3904 (.Y (nx3903), .A0 (q_17__8), .A1 (q_16__8), .S0 (nx7002)) ;
    dffr gen_regs_16_regi_reg_q_8 (.Q (q_16__8), .QB (\$dummy [208]), .D (nx3893
         ), .CLK (nx7118), .R (reset)) ;
    mux21_ni ix3894 (.Y (nx3893), .A0 (q_16__8), .A1 (q_15__8), .S0 (nx7000)) ;
    dffr gen_regs_15_regi_reg_q_8 (.Q (q_15__8), .QB (\$dummy [209]), .D (nx3883
         ), .CLK (nx7118), .R (reset)) ;
    mux21_ni ix3884 (.Y (nx3883), .A0 (q_15__8), .A1 (q_14__8), .S0 (nx7000)) ;
    dffr gen_regs_14_regi_reg_q_8 (.Q (q_14__8), .QB (\$dummy [210]), .D (nx3873
         ), .CLK (nx7118), .R (reset)) ;
    mux21_ni ix3874 (.Y (nx3873), .A0 (q_14__8), .A1 (q_13__8), .S0 (nx7000)) ;
    dffr gen_regs_13_regi_reg_q_8 (.Q (q_13__8), .QB (\$dummy [211]), .D (nx3863
         ), .CLK (nx7118), .R (reset)) ;
    mux21_ni ix3864 (.Y (nx3863), .A0 (q_13__8), .A1 (q_12__8), .S0 (nx7000)) ;
    dffr gen_regs_12_regi_reg_q_8 (.Q (q_12__8), .QB (\$dummy [212]), .D (nx3853
         ), .CLK (nx7118), .R (reset)) ;
    mux21_ni ix3854 (.Y (nx3853), .A0 (q_12__8), .A1 (q_11__8), .S0 (nx7000)) ;
    dffr gen_regs_11_regi_reg_q_8 (.Q (q_11__8), .QB (\$dummy [213]), .D (nx3843
         ), .CLK (nx7118), .R (reset)) ;
    mux21_ni ix3844 (.Y (nx3843), .A0 (q_11__8), .A1 (q_10__8), .S0 (nx7000)) ;
    dffr gen_regs_10_regi_reg_q_8 (.Q (q_10__8), .QB (\$dummy [214]), .D (nx3833
         ), .CLK (nx7118), .R (reset)) ;
    mux21_ni ix3834 (.Y (nx3833), .A0 (q_10__8), .A1 (q_9__8), .S0 (nx7000)) ;
    dffr gen_regs_9_regi_reg_q_8 (.Q (q_9__8), .QB (\$dummy [215]), .D (nx3823)
         , .CLK (nx7116), .R (reset)) ;
    mux21_ni ix3824 (.Y (nx3823), .A0 (q_9__8), .A1 (q_8__8), .S0 (nx6998)) ;
    dffr gen_regs_8_regi_reg_q_8 (.Q (q_8__8), .QB (\$dummy [216]), .D (nx3813)
         , .CLK (nx7116), .R (reset)) ;
    mux21_ni ix3814 (.Y (nx3813), .A0 (q_8__8), .A1 (q_7__8), .S0 (nx6998)) ;
    dffr gen_regs_7_regi_reg_q_8 (.Q (q_7__8), .QB (\$dummy [217]), .D (nx3803)
         , .CLK (nx7116), .R (reset)) ;
    mux21_ni ix3804 (.Y (nx3803), .A0 (q_7__8), .A1 (q_6__8), .S0 (nx6998)) ;
    dffr gen_regs_6_regi_reg_q_8 (.Q (q_6__8), .QB (\$dummy [218]), .D (nx3793)
         , .CLK (nx7116), .R (reset)) ;
    mux21_ni ix3794 (.Y (nx3793), .A0 (q_6__8), .A1 (q_5__8), .S0 (nx6998)) ;
    dffr gen_regs_5_regi_reg_q_8 (.Q (q_5__8), .QB (\$dummy [219]), .D (nx3783)
         , .CLK (nx7116), .R (reset)) ;
    mux21_ni ix3784 (.Y (nx3783), .A0 (q_5__8), .A1 (q_4__8), .S0 (nx6998)) ;
    dffr gen_regs_4_regi_reg_q_8 (.Q (q_4__8), .QB (\$dummy [220]), .D (nx3773)
         , .CLK (nx7116), .R (reset)) ;
    mux21_ni ix3774 (.Y (nx3773), .A0 (q_4__8), .A1 (q_3__8), .S0 (nx6998)) ;
    dffr gen_regs_3_regi_reg_q_8 (.Q (q_3__8), .QB (\$dummy [221]), .D (nx3763)
         , .CLK (nx7116), .R (reset)) ;
    mux21_ni ix3764 (.Y (nx3763), .A0 (q_3__8), .A1 (q_2__8), .S0 (nx6998)) ;
    dffr gen_regs_2_regi_reg_q_8 (.Q (q_2__8), .QB (\$dummy [222]), .D (nx3753)
         , .CLK (nx7114), .R (reset)) ;
    mux21_ni ix3754 (.Y (nx3753), .A0 (q_2__8), .A1 (q_1__8), .S0 (nx6996)) ;
    dffr gen_regs_1_regi_reg_q_8 (.Q (q_1__8), .QB (\$dummy [223]), .D (nx3743)
         , .CLK (nx7114), .R (reset)) ;
    mux21_ni ix3744 (.Y (nx3743), .A0 (q_1__8), .A1 (q_0__8), .S0 (nx6996)) ;
    dffr reg0_reg_q_8 (.Q (q_0__8), .QB (\$dummy [224]), .D (nx3733), .CLK (
         nx7114), .R (reset)) ;
    mux21_ni ix3734 (.Y (nx3733), .A0 (q_0__8), .A1 (d[8]), .S0 (nx6996)) ;
    dffr gen_regs_24_regi_reg_q_9 (.Q (q_24__9), .QB (\$dummy [225]), .D (nx4223
         ), .CLK (nx7128), .R (reset)) ;
    mux21_ni ix4224 (.Y (nx4223), .A0 (q_24__9), .A1 (q_23__9), .S0 (nx7010)) ;
    dffr gen_regs_23_regi_reg_q_9 (.Q (q_23__9), .QB (\$dummy [226]), .D (nx4213
         ), .CLK (nx7128), .R (reset)) ;
    mux21_ni ix4214 (.Y (nx4213), .A0 (q_23__9), .A1 (q_22__9), .S0 (nx7010)) ;
    dffr gen_regs_22_regi_reg_q_9 (.Q (q_22__9), .QB (\$dummy [227]), .D (nx4203
         ), .CLK (nx7128), .R (reset)) ;
    mux21_ni ix4204 (.Y (nx4203), .A0 (q_22__9), .A1 (q_21__9), .S0 (nx7010)) ;
    dffr gen_regs_21_regi_reg_q_9 (.Q (q_21__9), .QB (\$dummy [228]), .D (nx4193
         ), .CLK (nx7128), .R (reset)) ;
    mux21_ni ix4194 (.Y (nx4193), .A0 (q_21__9), .A1 (q_20__9), .S0 (nx7010)) ;
    dffr gen_regs_20_regi_reg_q_9 (.Q (q_20__9), .QB (\$dummy [229]), .D (nx4183
         ), .CLK (nx7128), .R (reset)) ;
    mux21_ni ix4184 (.Y (nx4183), .A0 (q_20__9), .A1 (q_19__9), .S0 (nx7010)) ;
    dffr gen_regs_19_regi_reg_q_9 (.Q (q_19__9), .QB (\$dummy [230]), .D (nx4173
         ), .CLK (nx7126), .R (reset)) ;
    mux21_ni ix4174 (.Y (nx4173), .A0 (q_19__9), .A1 (q_18__9), .S0 (nx7008)) ;
    dffr gen_regs_18_regi_reg_q_9 (.Q (q_18__9), .QB (\$dummy [231]), .D (nx4163
         ), .CLK (nx7126), .R (reset)) ;
    mux21_ni ix4164 (.Y (nx4163), .A0 (q_18__9), .A1 (q_17__9), .S0 (nx7008)) ;
    dffr gen_regs_17_regi_reg_q_9 (.Q (q_17__9), .QB (\$dummy [232]), .D (nx4153
         ), .CLK (nx7126), .R (reset)) ;
    mux21_ni ix4154 (.Y (nx4153), .A0 (q_17__9), .A1 (q_16__9), .S0 (nx7008)) ;
    dffr gen_regs_16_regi_reg_q_9 (.Q (q_16__9), .QB (\$dummy [233]), .D (nx4143
         ), .CLK (nx7126), .R (reset)) ;
    mux21_ni ix4144 (.Y (nx4143), .A0 (q_16__9), .A1 (q_15__9), .S0 (nx7008)) ;
    dffr gen_regs_15_regi_reg_q_9 (.Q (q_15__9), .QB (\$dummy [234]), .D (nx4133
         ), .CLK (nx7126), .R (reset)) ;
    mux21_ni ix4134 (.Y (nx4133), .A0 (q_15__9), .A1 (q_14__9), .S0 (nx7008)) ;
    dffr gen_regs_14_regi_reg_q_9 (.Q (q_14__9), .QB (\$dummy [235]), .D (nx4123
         ), .CLK (nx7126), .R (reset)) ;
    mux21_ni ix4124 (.Y (nx4123), .A0 (q_14__9), .A1 (q_13__9), .S0 (nx7008)) ;
    dffr gen_regs_13_regi_reg_q_9 (.Q (q_13__9), .QB (\$dummy [236]), .D (nx4113
         ), .CLK (nx7126), .R (reset)) ;
    mux21_ni ix4114 (.Y (nx4113), .A0 (q_13__9), .A1 (q_12__9), .S0 (nx7008)) ;
    dffr gen_regs_12_regi_reg_q_9 (.Q (q_12__9), .QB (\$dummy [237]), .D (nx4103
         ), .CLK (nx7124), .R (reset)) ;
    mux21_ni ix4104 (.Y (nx4103), .A0 (q_12__9), .A1 (q_11__9), .S0 (nx7006)) ;
    dffr gen_regs_11_regi_reg_q_9 (.Q (q_11__9), .QB (\$dummy [238]), .D (nx4093
         ), .CLK (nx7124), .R (reset)) ;
    mux21_ni ix4094 (.Y (nx4093), .A0 (q_11__9), .A1 (q_10__9), .S0 (nx7006)) ;
    dffr gen_regs_10_regi_reg_q_9 (.Q (q_10__9), .QB (\$dummy [239]), .D (nx4083
         ), .CLK (nx7124), .R (reset)) ;
    mux21_ni ix4084 (.Y (nx4083), .A0 (q_10__9), .A1 (q_9__9), .S0 (nx7006)) ;
    dffr gen_regs_9_regi_reg_q_9 (.Q (q_9__9), .QB (\$dummy [240]), .D (nx4073)
         , .CLK (nx7124), .R (reset)) ;
    mux21_ni ix4074 (.Y (nx4073), .A0 (q_9__9), .A1 (q_8__9), .S0 (nx7006)) ;
    dffr gen_regs_8_regi_reg_q_9 (.Q (q_8__9), .QB (\$dummy [241]), .D (nx4063)
         , .CLK (nx7124), .R (reset)) ;
    mux21_ni ix4064 (.Y (nx4063), .A0 (q_8__9), .A1 (q_7__9), .S0 (nx7006)) ;
    dffr gen_regs_7_regi_reg_q_9 (.Q (q_7__9), .QB (\$dummy [242]), .D (nx4053)
         , .CLK (nx7124), .R (reset)) ;
    mux21_ni ix4054 (.Y (nx4053), .A0 (q_7__9), .A1 (q_6__9), .S0 (nx7006)) ;
    dffr gen_regs_6_regi_reg_q_9 (.Q (q_6__9), .QB (\$dummy [243]), .D (nx4043)
         , .CLK (nx7124), .R (reset)) ;
    mux21_ni ix4044 (.Y (nx4043), .A0 (q_6__9), .A1 (q_5__9), .S0 (nx7006)) ;
    dffr gen_regs_5_regi_reg_q_9 (.Q (q_5__9), .QB (\$dummy [244]), .D (nx4033)
         , .CLK (nx7122), .R (reset)) ;
    mux21_ni ix4034 (.Y (nx4033), .A0 (q_5__9), .A1 (q_4__9), .S0 (nx7004)) ;
    dffr gen_regs_4_regi_reg_q_9 (.Q (q_4__9), .QB (\$dummy [245]), .D (nx4023)
         , .CLK (nx7122), .R (reset)) ;
    mux21_ni ix4024 (.Y (nx4023), .A0 (q_4__9), .A1 (q_3__9), .S0 (nx7004)) ;
    dffr gen_regs_3_regi_reg_q_9 (.Q (q_3__9), .QB (\$dummy [246]), .D (nx4013)
         , .CLK (nx7122), .R (reset)) ;
    mux21_ni ix4014 (.Y (nx4013), .A0 (q_3__9), .A1 (q_2__9), .S0 (nx7004)) ;
    dffr gen_regs_2_regi_reg_q_9 (.Q (q_2__9), .QB (\$dummy [247]), .D (nx4003)
         , .CLK (nx7122), .R (reset)) ;
    mux21_ni ix4004 (.Y (nx4003), .A0 (q_2__9), .A1 (q_1__9), .S0 (nx7004)) ;
    dffr gen_regs_1_regi_reg_q_9 (.Q (q_1__9), .QB (\$dummy [248]), .D (nx3993)
         , .CLK (nx7122), .R (reset)) ;
    mux21_ni ix3994 (.Y (nx3993), .A0 (q_1__9), .A1 (q_0__9), .S0 (nx7004)) ;
    dffr reg0_reg_q_9 (.Q (q_0__9), .QB (\$dummy [249]), .D (nx3983), .CLK (
         nx7122), .R (reset)) ;
    mux21_ni ix3984 (.Y (nx3983), .A0 (q_0__9), .A1 (d[9]), .S0 (nx7004)) ;
    dffr gen_regs_24_regi_reg_q_10 (.Q (q_24__10), .QB (\$dummy [250]), .D (
         nx4473), .CLK (nx7136), .R (reset)) ;
    mux21_ni ix4474 (.Y (nx4473), .A0 (q_24__10), .A1 (q_23__10), .S0 (nx7018)
             ) ;
    dffr gen_regs_23_regi_reg_q_10 (.Q (q_23__10), .QB (\$dummy [251]), .D (
         nx4463), .CLK (nx7136), .R (reset)) ;
    mux21_ni ix4464 (.Y (nx4463), .A0 (q_23__10), .A1 (q_22__10), .S0 (nx7018)
             ) ;
    dffr gen_regs_22_regi_reg_q_10 (.Q (q_22__10), .QB (\$dummy [252]), .D (
         nx4453), .CLK (nx7134), .R (reset)) ;
    mux21_ni ix4454 (.Y (nx4453), .A0 (q_22__10), .A1 (q_21__10), .S0 (nx7016)
             ) ;
    dffr gen_regs_21_regi_reg_q_10 (.Q (q_21__10), .QB (\$dummy [253]), .D (
         nx4443), .CLK (nx7134), .R (reset)) ;
    mux21_ni ix4444 (.Y (nx4443), .A0 (q_21__10), .A1 (q_20__10), .S0 (nx7016)
             ) ;
    dffr gen_regs_20_regi_reg_q_10 (.Q (q_20__10), .QB (\$dummy [254]), .D (
         nx4433), .CLK (nx7134), .R (reset)) ;
    mux21_ni ix4434 (.Y (nx4433), .A0 (q_20__10), .A1 (q_19__10), .S0 (nx7016)
             ) ;
    dffr gen_regs_19_regi_reg_q_10 (.Q (q_19__10), .QB (\$dummy [255]), .D (
         nx4423), .CLK (nx7134), .R (reset)) ;
    mux21_ni ix4424 (.Y (nx4423), .A0 (q_19__10), .A1 (q_18__10), .S0 (nx7016)
             ) ;
    dffr gen_regs_18_regi_reg_q_10 (.Q (q_18__10), .QB (\$dummy [256]), .D (
         nx4413), .CLK (nx7134), .R (reset)) ;
    mux21_ni ix4414 (.Y (nx4413), .A0 (q_18__10), .A1 (q_17__10), .S0 (nx7016)
             ) ;
    dffr gen_regs_17_regi_reg_q_10 (.Q (q_17__10), .QB (\$dummy [257]), .D (
         nx4403), .CLK (nx7134), .R (reset)) ;
    mux21_ni ix4404 (.Y (nx4403), .A0 (q_17__10), .A1 (q_16__10), .S0 (nx7016)
             ) ;
    dffr gen_regs_16_regi_reg_q_10 (.Q (q_16__10), .QB (\$dummy [258]), .D (
         nx4393), .CLK (nx7134), .R (reset)) ;
    mux21_ni ix4394 (.Y (nx4393), .A0 (q_16__10), .A1 (q_15__10), .S0 (nx7016)
             ) ;
    dffr gen_regs_15_regi_reg_q_10 (.Q (q_15__10), .QB (\$dummy [259]), .D (
         nx4383), .CLK (nx7132), .R (reset)) ;
    mux21_ni ix4384 (.Y (nx4383), .A0 (q_15__10), .A1 (q_14__10), .S0 (nx7014)
             ) ;
    dffr gen_regs_14_regi_reg_q_10 (.Q (q_14__10), .QB (\$dummy [260]), .D (
         nx4373), .CLK (nx7132), .R (reset)) ;
    mux21_ni ix4374 (.Y (nx4373), .A0 (q_14__10), .A1 (q_13__10), .S0 (nx7014)
             ) ;
    dffr gen_regs_13_regi_reg_q_10 (.Q (q_13__10), .QB (\$dummy [261]), .D (
         nx4363), .CLK (nx7132), .R (reset)) ;
    mux21_ni ix4364 (.Y (nx4363), .A0 (q_13__10), .A1 (q_12__10), .S0 (nx7014)
             ) ;
    dffr gen_regs_12_regi_reg_q_10 (.Q (q_12__10), .QB (\$dummy [262]), .D (
         nx4353), .CLK (nx7132), .R (reset)) ;
    mux21_ni ix4354 (.Y (nx4353), .A0 (q_12__10), .A1 (q_11__10), .S0 (nx7014)
             ) ;
    dffr gen_regs_11_regi_reg_q_10 (.Q (q_11__10), .QB (\$dummy [263]), .D (
         nx4343), .CLK (nx7132), .R (reset)) ;
    mux21_ni ix4344 (.Y (nx4343), .A0 (q_11__10), .A1 (q_10__10), .S0 (nx7014)
             ) ;
    dffr gen_regs_10_regi_reg_q_10 (.Q (q_10__10), .QB (\$dummy [264]), .D (
         nx4333), .CLK (nx7132), .R (reset)) ;
    mux21_ni ix4334 (.Y (nx4333), .A0 (q_10__10), .A1 (q_9__10), .S0 (nx7014)) ;
    dffr gen_regs_9_regi_reg_q_10 (.Q (q_9__10), .QB (\$dummy [265]), .D (nx4323
         ), .CLK (nx7132), .R (reset)) ;
    mux21_ni ix4324 (.Y (nx4323), .A0 (q_9__10), .A1 (q_8__10), .S0 (nx7014)) ;
    dffr gen_regs_8_regi_reg_q_10 (.Q (q_8__10), .QB (\$dummy [266]), .D (nx4313
         ), .CLK (nx7130), .R (reset)) ;
    mux21_ni ix4314 (.Y (nx4313), .A0 (q_8__10), .A1 (q_7__10), .S0 (nx7012)) ;
    dffr gen_regs_7_regi_reg_q_10 (.Q (q_7__10), .QB (\$dummy [267]), .D (nx4303
         ), .CLK (nx7130), .R (reset)) ;
    mux21_ni ix4304 (.Y (nx4303), .A0 (q_7__10), .A1 (q_6__10), .S0 (nx7012)) ;
    dffr gen_regs_6_regi_reg_q_10 (.Q (q_6__10), .QB (\$dummy [268]), .D (nx4293
         ), .CLK (nx7130), .R (reset)) ;
    mux21_ni ix4294 (.Y (nx4293), .A0 (q_6__10), .A1 (q_5__10), .S0 (nx7012)) ;
    dffr gen_regs_5_regi_reg_q_10 (.Q (q_5__10), .QB (\$dummy [269]), .D (nx4283
         ), .CLK (nx7130), .R (reset)) ;
    mux21_ni ix4284 (.Y (nx4283), .A0 (q_5__10), .A1 (q_4__10), .S0 (nx7012)) ;
    dffr gen_regs_4_regi_reg_q_10 (.Q (q_4__10), .QB (\$dummy [270]), .D (nx4273
         ), .CLK (nx7130), .R (reset)) ;
    mux21_ni ix4274 (.Y (nx4273), .A0 (q_4__10), .A1 (q_3__10), .S0 (nx7012)) ;
    dffr gen_regs_3_regi_reg_q_10 (.Q (q_3__10), .QB (\$dummy [271]), .D (nx4263
         ), .CLK (nx7130), .R (reset)) ;
    mux21_ni ix4264 (.Y (nx4263), .A0 (q_3__10), .A1 (q_2__10), .S0 (nx7012)) ;
    dffr gen_regs_2_regi_reg_q_10 (.Q (q_2__10), .QB (\$dummy [272]), .D (nx4253
         ), .CLK (nx7130), .R (reset)) ;
    mux21_ni ix4254 (.Y (nx4253), .A0 (q_2__10), .A1 (q_1__10), .S0 (nx7012)) ;
    dffr gen_regs_1_regi_reg_q_10 (.Q (q_1__10), .QB (\$dummy [273]), .D (nx4243
         ), .CLK (nx7128), .R (reset)) ;
    mux21_ni ix4244 (.Y (nx4243), .A0 (q_1__10), .A1 (q_0__10), .S0 (nx7010)) ;
    dffr reg0_reg_q_10 (.Q (q_0__10), .QB (\$dummy [274]), .D (nx4233), .CLK (
         nx7128), .R (reset)) ;
    mux21_ni ix4234 (.Y (nx4233), .A0 (q_0__10), .A1 (d[10]), .S0 (nx7010)) ;
    dffr gen_regs_24_regi_reg_q_11 (.Q (q_24__11), .QB (\$dummy [275]), .D (
         nx4723), .CLK (nx7142), .R (reset)) ;
    mux21_ni ix4724 (.Y (nx4723), .A0 (q_24__11), .A1 (q_23__11), .S0 (nx7024)
             ) ;
    dffr gen_regs_23_regi_reg_q_11 (.Q (q_23__11), .QB (\$dummy [276]), .D (
         nx4713), .CLK (nx7142), .R (reset)) ;
    mux21_ni ix4714 (.Y (nx4713), .A0 (q_23__11), .A1 (q_22__11), .S0 (nx7024)
             ) ;
    dffr gen_regs_22_regi_reg_q_11 (.Q (q_22__11), .QB (\$dummy [277]), .D (
         nx4703), .CLK (nx7142), .R (reset)) ;
    mux21_ni ix4704 (.Y (nx4703), .A0 (q_22__11), .A1 (q_21__11), .S0 (nx7024)
             ) ;
    dffr gen_regs_21_regi_reg_q_11 (.Q (q_21__11), .QB (\$dummy [278]), .D (
         nx4693), .CLK (nx7142), .R (reset)) ;
    mux21_ni ix4694 (.Y (nx4693), .A0 (q_21__11), .A1 (q_20__11), .S0 (nx7024)
             ) ;
    dffr gen_regs_20_regi_reg_q_11 (.Q (q_20__11), .QB (\$dummy [279]), .D (
         nx4683), .CLK (nx7142), .R (reset)) ;
    mux21_ni ix4684 (.Y (nx4683), .A0 (q_20__11), .A1 (q_19__11), .S0 (nx7024)
             ) ;
    dffr gen_regs_19_regi_reg_q_11 (.Q (q_19__11), .QB (\$dummy [280]), .D (
         nx4673), .CLK (nx7142), .R (reset)) ;
    mux21_ni ix4674 (.Y (nx4673), .A0 (q_19__11), .A1 (q_18__11), .S0 (nx7024)
             ) ;
    dffr gen_regs_18_regi_reg_q_11 (.Q (q_18__11), .QB (\$dummy [281]), .D (
         nx4663), .CLK (nx7140), .R (reset)) ;
    mux21_ni ix4664 (.Y (nx4663), .A0 (q_18__11), .A1 (q_17__11), .S0 (nx7022)
             ) ;
    dffr gen_regs_17_regi_reg_q_11 (.Q (q_17__11), .QB (\$dummy [282]), .D (
         nx4653), .CLK (nx7140), .R (reset)) ;
    mux21_ni ix4654 (.Y (nx4653), .A0 (q_17__11), .A1 (q_16__11), .S0 (nx7022)
             ) ;
    dffr gen_regs_16_regi_reg_q_11 (.Q (q_16__11), .QB (\$dummy [283]), .D (
         nx4643), .CLK (nx7140), .R (reset)) ;
    mux21_ni ix4644 (.Y (nx4643), .A0 (q_16__11), .A1 (q_15__11), .S0 (nx7022)
             ) ;
    dffr gen_regs_15_regi_reg_q_11 (.Q (q_15__11), .QB (\$dummy [284]), .D (
         nx4633), .CLK (nx7140), .R (reset)) ;
    mux21_ni ix4634 (.Y (nx4633), .A0 (q_15__11), .A1 (q_14__11), .S0 (nx7022)
             ) ;
    dffr gen_regs_14_regi_reg_q_11 (.Q (q_14__11), .QB (\$dummy [285]), .D (
         nx4623), .CLK (nx7140), .R (reset)) ;
    mux21_ni ix4624 (.Y (nx4623), .A0 (q_14__11), .A1 (q_13__11), .S0 (nx7022)
             ) ;
    dffr gen_regs_13_regi_reg_q_11 (.Q (q_13__11), .QB (\$dummy [286]), .D (
         nx4613), .CLK (nx7140), .R (reset)) ;
    mux21_ni ix4614 (.Y (nx4613), .A0 (q_13__11), .A1 (q_12__11), .S0 (nx7022)
             ) ;
    dffr gen_regs_12_regi_reg_q_11 (.Q (q_12__11), .QB (\$dummy [287]), .D (
         nx4603), .CLK (nx7140), .R (reset)) ;
    mux21_ni ix4604 (.Y (nx4603), .A0 (q_12__11), .A1 (q_11__11), .S0 (nx7022)
             ) ;
    dffr gen_regs_11_regi_reg_q_11 (.Q (q_11__11), .QB (\$dummy [288]), .D (
         nx4593), .CLK (nx7138), .R (reset)) ;
    mux21_ni ix4594 (.Y (nx4593), .A0 (q_11__11), .A1 (q_10__11), .S0 (nx7020)
             ) ;
    dffr gen_regs_10_regi_reg_q_11 (.Q (q_10__11), .QB (\$dummy [289]), .D (
         nx4583), .CLK (nx7138), .R (reset)) ;
    mux21_ni ix4584 (.Y (nx4583), .A0 (q_10__11), .A1 (q_9__11), .S0 (nx7020)) ;
    dffr gen_regs_9_regi_reg_q_11 (.Q (q_9__11), .QB (\$dummy [290]), .D (nx4573
         ), .CLK (nx7138), .R (reset)) ;
    mux21_ni ix4574 (.Y (nx4573), .A0 (q_9__11), .A1 (q_8__11), .S0 (nx7020)) ;
    dffr gen_regs_8_regi_reg_q_11 (.Q (q_8__11), .QB (\$dummy [291]), .D (nx4563
         ), .CLK (nx7138), .R (reset)) ;
    mux21_ni ix4564 (.Y (nx4563), .A0 (q_8__11), .A1 (q_7__11), .S0 (nx7020)) ;
    dffr gen_regs_7_regi_reg_q_11 (.Q (q_7__11), .QB (\$dummy [292]), .D (nx4553
         ), .CLK (nx7138), .R (reset)) ;
    mux21_ni ix4554 (.Y (nx4553), .A0 (q_7__11), .A1 (q_6__11), .S0 (nx7020)) ;
    dffr gen_regs_6_regi_reg_q_11 (.Q (q_6__11), .QB (\$dummy [293]), .D (nx4543
         ), .CLK (nx7138), .R (reset)) ;
    mux21_ni ix4544 (.Y (nx4543), .A0 (q_6__11), .A1 (q_5__11), .S0 (nx7020)) ;
    dffr gen_regs_5_regi_reg_q_11 (.Q (q_5__11), .QB (\$dummy [294]), .D (nx4533
         ), .CLK (nx7138), .R (reset)) ;
    mux21_ni ix4534 (.Y (nx4533), .A0 (q_5__11), .A1 (q_4__11), .S0 (nx7020)) ;
    dffr gen_regs_4_regi_reg_q_11 (.Q (q_4__11), .QB (\$dummy [295]), .D (nx4523
         ), .CLK (nx7136), .R (reset)) ;
    mux21_ni ix4524 (.Y (nx4523), .A0 (q_4__11), .A1 (q_3__11), .S0 (nx7018)) ;
    dffr gen_regs_3_regi_reg_q_11 (.Q (q_3__11), .QB (\$dummy [296]), .D (nx4513
         ), .CLK (nx7136), .R (reset)) ;
    mux21_ni ix4514 (.Y (nx4513), .A0 (q_3__11), .A1 (q_2__11), .S0 (nx7018)) ;
    dffr gen_regs_2_regi_reg_q_11 (.Q (q_2__11), .QB (\$dummy [297]), .D (nx4503
         ), .CLK (nx7136), .R (reset)) ;
    mux21_ni ix4504 (.Y (nx4503), .A0 (q_2__11), .A1 (q_1__11), .S0 (nx7018)) ;
    dffr gen_regs_1_regi_reg_q_11 (.Q (q_1__11), .QB (\$dummy [298]), .D (nx4493
         ), .CLK (nx7136), .R (reset)) ;
    mux21_ni ix4494 (.Y (nx4493), .A0 (q_1__11), .A1 (q_0__11), .S0 (nx7018)) ;
    dffr reg0_reg_q_11 (.Q (q_0__11), .QB (\$dummy [299]), .D (nx4483), .CLK (
         nx7136), .R (reset)) ;
    mux21_ni ix4484 (.Y (nx4483), .A0 (q_0__11), .A1 (d[11]), .S0 (nx7018)) ;
    dffr gen_regs_24_regi_reg_q_12 (.Q (q_24__12), .QB (\$dummy [300]), .D (
         nx4973), .CLK (nx7150), .R (reset)) ;
    mux21_ni ix4974 (.Y (nx4973), .A0 (q_24__12), .A1 (q_23__12), .S0 (nx7032)
             ) ;
    dffr gen_regs_23_regi_reg_q_12 (.Q (q_23__12), .QB (\$dummy [301]), .D (
         nx4963), .CLK (nx7150), .R (reset)) ;
    mux21_ni ix4964 (.Y (nx4963), .A0 (q_23__12), .A1 (q_22__12), .S0 (nx7032)
             ) ;
    dffr gen_regs_22_regi_reg_q_12 (.Q (q_22__12), .QB (\$dummy [302]), .D (
         nx4953), .CLK (nx7150), .R (reset)) ;
    mux21_ni ix4954 (.Y (nx4953), .A0 (q_22__12), .A1 (q_21__12), .S0 (nx7032)
             ) ;
    dffr gen_regs_21_regi_reg_q_12 (.Q (q_21__12), .QB (\$dummy [303]), .D (
         nx4943), .CLK (nx7148), .R (reset)) ;
    mux21_ni ix4944 (.Y (nx4943), .A0 (q_21__12), .A1 (q_20__12), .S0 (nx7030)
             ) ;
    dffr gen_regs_20_regi_reg_q_12 (.Q (q_20__12), .QB (\$dummy [304]), .D (
         nx4933), .CLK (nx7148), .R (reset)) ;
    mux21_ni ix4934 (.Y (nx4933), .A0 (q_20__12), .A1 (q_19__12), .S0 (nx7030)
             ) ;
    dffr gen_regs_19_regi_reg_q_12 (.Q (q_19__12), .QB (\$dummy [305]), .D (
         nx4923), .CLK (nx7148), .R (reset)) ;
    mux21_ni ix4924 (.Y (nx4923), .A0 (q_19__12), .A1 (q_18__12), .S0 (nx7030)
             ) ;
    dffr gen_regs_18_regi_reg_q_12 (.Q (q_18__12), .QB (\$dummy [306]), .D (
         nx4913), .CLK (nx7148), .R (reset)) ;
    mux21_ni ix4914 (.Y (nx4913), .A0 (q_18__12), .A1 (q_17__12), .S0 (nx7030)
             ) ;
    dffr gen_regs_17_regi_reg_q_12 (.Q (q_17__12), .QB (\$dummy [307]), .D (
         nx4903), .CLK (nx7148), .R (reset)) ;
    mux21_ni ix4904 (.Y (nx4903), .A0 (q_17__12), .A1 (q_16__12), .S0 (nx7030)
             ) ;
    dffr gen_regs_16_regi_reg_q_12 (.Q (q_16__12), .QB (\$dummy [308]), .D (
         nx4893), .CLK (nx7148), .R (reset)) ;
    mux21_ni ix4894 (.Y (nx4893), .A0 (q_16__12), .A1 (q_15__12), .S0 (nx7030)
             ) ;
    dffr gen_regs_15_regi_reg_q_12 (.Q (q_15__12), .QB (\$dummy [309]), .D (
         nx4883), .CLK (nx7148), .R (reset)) ;
    mux21_ni ix4884 (.Y (nx4883), .A0 (q_15__12), .A1 (q_14__12), .S0 (nx7030)
             ) ;
    dffr gen_regs_14_regi_reg_q_12 (.Q (q_14__12), .QB (\$dummy [310]), .D (
         nx4873), .CLK (nx7146), .R (reset)) ;
    mux21_ni ix4874 (.Y (nx4873), .A0 (q_14__12), .A1 (q_13__12), .S0 (nx7028)
             ) ;
    dffr gen_regs_13_regi_reg_q_12 (.Q (q_13__12), .QB (\$dummy [311]), .D (
         nx4863), .CLK (nx7146), .R (reset)) ;
    mux21_ni ix4864 (.Y (nx4863), .A0 (q_13__12), .A1 (q_12__12), .S0 (nx7028)
             ) ;
    dffr gen_regs_12_regi_reg_q_12 (.Q (q_12__12), .QB (\$dummy [312]), .D (
         nx4853), .CLK (nx7146), .R (reset)) ;
    mux21_ni ix4854 (.Y (nx4853), .A0 (q_12__12), .A1 (q_11__12), .S0 (nx7028)
             ) ;
    dffr gen_regs_11_regi_reg_q_12 (.Q (q_11__12), .QB (\$dummy [313]), .D (
         nx4843), .CLK (nx7146), .R (reset)) ;
    mux21_ni ix4844 (.Y (nx4843), .A0 (q_11__12), .A1 (q_10__12), .S0 (nx7028)
             ) ;
    dffr gen_regs_10_regi_reg_q_12 (.Q (q_10__12), .QB (\$dummy [314]), .D (
         nx4833), .CLK (nx7146), .R (reset)) ;
    mux21_ni ix4834 (.Y (nx4833), .A0 (q_10__12), .A1 (q_9__12), .S0 (nx7028)) ;
    dffr gen_regs_9_regi_reg_q_12 (.Q (q_9__12), .QB (\$dummy [315]), .D (nx4823
         ), .CLK (nx7146), .R (reset)) ;
    mux21_ni ix4824 (.Y (nx4823), .A0 (q_9__12), .A1 (q_8__12), .S0 (nx7028)) ;
    dffr gen_regs_8_regi_reg_q_12 (.Q (q_8__12), .QB (\$dummy [316]), .D (nx4813
         ), .CLK (nx7146), .R (reset)) ;
    mux21_ni ix4814 (.Y (nx4813), .A0 (q_8__12), .A1 (q_7__12), .S0 (nx7028)) ;
    dffr gen_regs_7_regi_reg_q_12 (.Q (q_7__12), .QB (\$dummy [317]), .D (nx4803
         ), .CLK (nx7144), .R (reset)) ;
    mux21_ni ix4804 (.Y (nx4803), .A0 (q_7__12), .A1 (q_6__12), .S0 (nx7026)) ;
    dffr gen_regs_6_regi_reg_q_12 (.Q (q_6__12), .QB (\$dummy [318]), .D (nx4793
         ), .CLK (nx7144), .R (reset)) ;
    mux21_ni ix4794 (.Y (nx4793), .A0 (q_6__12), .A1 (q_5__12), .S0 (nx7026)) ;
    dffr gen_regs_5_regi_reg_q_12 (.Q (q_5__12), .QB (\$dummy [319]), .D (nx4783
         ), .CLK (nx7144), .R (reset)) ;
    mux21_ni ix4784 (.Y (nx4783), .A0 (q_5__12), .A1 (q_4__12), .S0 (nx7026)) ;
    dffr gen_regs_4_regi_reg_q_12 (.Q (q_4__12), .QB (\$dummy [320]), .D (nx4773
         ), .CLK (nx7144), .R (reset)) ;
    mux21_ni ix4774 (.Y (nx4773), .A0 (q_4__12), .A1 (q_3__12), .S0 (nx7026)) ;
    dffr gen_regs_3_regi_reg_q_12 (.Q (q_3__12), .QB (\$dummy [321]), .D (nx4763
         ), .CLK (nx7144), .R (reset)) ;
    mux21_ni ix4764 (.Y (nx4763), .A0 (q_3__12), .A1 (q_2__12), .S0 (nx7026)) ;
    dffr gen_regs_2_regi_reg_q_12 (.Q (q_2__12), .QB (\$dummy [322]), .D (nx4753
         ), .CLK (nx7144), .R (reset)) ;
    mux21_ni ix4754 (.Y (nx4753), .A0 (q_2__12), .A1 (q_1__12), .S0 (nx7026)) ;
    dffr gen_regs_1_regi_reg_q_12 (.Q (q_1__12), .QB (\$dummy [323]), .D (nx4743
         ), .CLK (nx7144), .R (reset)) ;
    mux21_ni ix4744 (.Y (nx4743), .A0 (q_1__12), .A1 (q_0__12), .S0 (nx7026)) ;
    dffr reg0_reg_q_12 (.Q (q_0__12), .QB (\$dummy [324]), .D (nx4733), .CLK (
         nx7142), .R (reset)) ;
    mux21_ni ix4734 (.Y (nx4733), .A0 (q_0__12), .A1 (d[12]), .S0 (nx7024)) ;
    dffr gen_regs_24_regi_reg_q_13 (.Q (q_24__13), .QB (\$dummy [325]), .D (
         nx5223), .CLK (nx7156), .R (reset)) ;
    mux21_ni ix5224 (.Y (nx5223), .A0 (q_24__13), .A1 (q_23__13), .S0 (nx7038)
             ) ;
    dffr gen_regs_23_regi_reg_q_13 (.Q (q_23__13), .QB (\$dummy [326]), .D (
         nx5213), .CLK (nx7156), .R (reset)) ;
    mux21_ni ix5214 (.Y (nx5213), .A0 (q_23__13), .A1 (q_22__13), .S0 (nx7038)
             ) ;
    dffr gen_regs_22_regi_reg_q_13 (.Q (q_22__13), .QB (\$dummy [327]), .D (
         nx5203), .CLK (nx7156), .R (reset)) ;
    mux21_ni ix5204 (.Y (nx5203), .A0 (q_22__13), .A1 (q_21__13), .S0 (nx7038)
             ) ;
    dffr gen_regs_21_regi_reg_q_13 (.Q (q_21__13), .QB (\$dummy [328]), .D (
         nx5193), .CLK (nx7156), .R (reset)) ;
    mux21_ni ix5194 (.Y (nx5193), .A0 (q_21__13), .A1 (q_20__13), .S0 (nx7038)
             ) ;
    dffr gen_regs_20_regi_reg_q_13 (.Q (q_20__13), .QB (\$dummy [329]), .D (
         nx5183), .CLK (nx7156), .R (reset)) ;
    mux21_ni ix5184 (.Y (nx5183), .A0 (q_20__13), .A1 (q_19__13), .S0 (nx7038)
             ) ;
    dffr gen_regs_19_regi_reg_q_13 (.Q (q_19__13), .QB (\$dummy [330]), .D (
         nx5173), .CLK (nx7156), .R (reset)) ;
    mux21_ni ix5174 (.Y (nx5173), .A0 (q_19__13), .A1 (q_18__13), .S0 (nx7038)
             ) ;
    dffr gen_regs_18_regi_reg_q_13 (.Q (q_18__13), .QB (\$dummy [331]), .D (
         nx5163), .CLK (nx7156), .R (reset)) ;
    mux21_ni ix5164 (.Y (nx5163), .A0 (q_18__13), .A1 (q_17__13), .S0 (nx7038)
             ) ;
    dffr gen_regs_17_regi_reg_q_13 (.Q (q_17__13), .QB (\$dummy [332]), .D (
         nx5153), .CLK (nx7154), .R (reset)) ;
    mux21_ni ix5154 (.Y (nx5153), .A0 (q_17__13), .A1 (q_16__13), .S0 (nx7036)
             ) ;
    dffr gen_regs_16_regi_reg_q_13 (.Q (q_16__13), .QB (\$dummy [333]), .D (
         nx5143), .CLK (nx7154), .R (reset)) ;
    mux21_ni ix5144 (.Y (nx5143), .A0 (q_16__13), .A1 (q_15__13), .S0 (nx7036)
             ) ;
    dffr gen_regs_15_regi_reg_q_13 (.Q (q_15__13), .QB (\$dummy [334]), .D (
         nx5133), .CLK (nx7154), .R (reset)) ;
    mux21_ni ix5134 (.Y (nx5133), .A0 (q_15__13), .A1 (q_14__13), .S0 (nx7036)
             ) ;
    dffr gen_regs_14_regi_reg_q_13 (.Q (q_14__13), .QB (\$dummy [335]), .D (
         nx5123), .CLK (nx7154), .R (reset)) ;
    mux21_ni ix5124 (.Y (nx5123), .A0 (q_14__13), .A1 (q_13__13), .S0 (nx7036)
             ) ;
    dffr gen_regs_13_regi_reg_q_13 (.Q (q_13__13), .QB (\$dummy [336]), .D (
         nx5113), .CLK (nx7154), .R (reset)) ;
    mux21_ni ix5114 (.Y (nx5113), .A0 (q_13__13), .A1 (q_12__13), .S0 (nx7036)
             ) ;
    dffr gen_regs_12_regi_reg_q_13 (.Q (q_12__13), .QB (\$dummy [337]), .D (
         nx5103), .CLK (nx7154), .R (reset)) ;
    mux21_ni ix5104 (.Y (nx5103), .A0 (q_12__13), .A1 (q_11__13), .S0 (nx7036)
             ) ;
    dffr gen_regs_11_regi_reg_q_13 (.Q (q_11__13), .QB (\$dummy [338]), .D (
         nx5093), .CLK (nx7154), .R (reset)) ;
    mux21_ni ix5094 (.Y (nx5093), .A0 (q_11__13), .A1 (q_10__13), .S0 (nx7036)
             ) ;
    dffr gen_regs_10_regi_reg_q_13 (.Q (q_10__13), .QB (\$dummy [339]), .D (
         nx5083), .CLK (nx7152), .R (reset)) ;
    mux21_ni ix5084 (.Y (nx5083), .A0 (q_10__13), .A1 (q_9__13), .S0 (nx7034)) ;
    dffr gen_regs_9_regi_reg_q_13 (.Q (q_9__13), .QB (\$dummy [340]), .D (nx5073
         ), .CLK (nx7152), .R (reset)) ;
    mux21_ni ix5074 (.Y (nx5073), .A0 (q_9__13), .A1 (q_8__13), .S0 (nx7034)) ;
    dffr gen_regs_8_regi_reg_q_13 (.Q (q_8__13), .QB (\$dummy [341]), .D (nx5063
         ), .CLK (nx7152), .R (reset)) ;
    mux21_ni ix5064 (.Y (nx5063), .A0 (q_8__13), .A1 (q_7__13), .S0 (nx7034)) ;
    dffr gen_regs_7_regi_reg_q_13 (.Q (q_7__13), .QB (\$dummy [342]), .D (nx5053
         ), .CLK (nx7152), .R (reset)) ;
    mux21_ni ix5054 (.Y (nx5053), .A0 (q_7__13), .A1 (q_6__13), .S0 (nx7034)) ;
    dffr gen_regs_6_regi_reg_q_13 (.Q (q_6__13), .QB (\$dummy [343]), .D (nx5043
         ), .CLK (nx7152), .R (reset)) ;
    mux21_ni ix5044 (.Y (nx5043), .A0 (q_6__13), .A1 (q_5__13), .S0 (nx7034)) ;
    dffr gen_regs_5_regi_reg_q_13 (.Q (q_5__13), .QB (\$dummy [344]), .D (nx5033
         ), .CLK (nx7152), .R (reset)) ;
    mux21_ni ix5034 (.Y (nx5033), .A0 (q_5__13), .A1 (q_4__13), .S0 (nx7034)) ;
    dffr gen_regs_4_regi_reg_q_13 (.Q (q_4__13), .QB (\$dummy [345]), .D (nx5023
         ), .CLK (nx7152), .R (reset)) ;
    mux21_ni ix5024 (.Y (nx5023), .A0 (q_4__13), .A1 (q_3__13), .S0 (nx7034)) ;
    dffr gen_regs_3_regi_reg_q_13 (.Q (q_3__13), .QB (\$dummy [346]), .D (nx5013
         ), .CLK (nx7150), .R (reset)) ;
    mux21_ni ix5014 (.Y (nx5013), .A0 (q_3__13), .A1 (q_2__13), .S0 (nx7032)) ;
    dffr gen_regs_2_regi_reg_q_13 (.Q (q_2__13), .QB (\$dummy [347]), .D (nx5003
         ), .CLK (nx7150), .R (reset)) ;
    mux21_ni ix5004 (.Y (nx5003), .A0 (q_2__13), .A1 (q_1__13), .S0 (nx7032)) ;
    dffr gen_regs_1_regi_reg_q_13 (.Q (q_1__13), .QB (\$dummy [348]), .D (nx4993
         ), .CLK (nx7150), .R (reset)) ;
    mux21_ni ix4994 (.Y (nx4993), .A0 (q_1__13), .A1 (q_0__13), .S0 (nx7032)) ;
    dffr reg0_reg_q_13 (.Q (q_0__13), .QB (\$dummy [349]), .D (nx4983), .CLK (
         nx7150), .R (reset)) ;
    mux21_ni ix4984 (.Y (nx4983), .A0 (q_0__13), .A1 (d[13]), .S0 (nx7032)) ;
    dffr gen_regs_24_regi_reg_q_14 (.Q (q_24__14), .QB (\$dummy [350]), .D (
         nx5473), .CLK (nx7164), .R (reset)) ;
    mux21_ni ix5474 (.Y (nx5473), .A0 (q_24__14), .A1 (q_23__14), .S0 (nx7046)
             ) ;
    dffr gen_regs_23_regi_reg_q_14 (.Q (q_23__14), .QB (\$dummy [351]), .D (
         nx5463), .CLK (nx7164), .R (reset)) ;
    mux21_ni ix5464 (.Y (nx5463), .A0 (q_23__14), .A1 (q_22__14), .S0 (nx7046)
             ) ;
    dffr gen_regs_22_regi_reg_q_14 (.Q (q_22__14), .QB (\$dummy [352]), .D (
         nx5453), .CLK (nx7164), .R (reset)) ;
    mux21_ni ix5454 (.Y (nx5453), .A0 (q_22__14), .A1 (q_21__14), .S0 (nx7046)
             ) ;
    dffr gen_regs_21_regi_reg_q_14 (.Q (q_21__14), .QB (\$dummy [353]), .D (
         nx5443), .CLK (nx7164), .R (reset)) ;
    mux21_ni ix5444 (.Y (nx5443), .A0 (q_21__14), .A1 (q_20__14), .S0 (nx7046)
             ) ;
    dffr gen_regs_20_regi_reg_q_14 (.Q (q_20__14), .QB (\$dummy [354]), .D (
         nx5433), .CLK (nx7162), .R (reset)) ;
    mux21_ni ix5434 (.Y (nx5433), .A0 (q_20__14), .A1 (q_19__14), .S0 (nx7044)
             ) ;
    dffr gen_regs_19_regi_reg_q_14 (.Q (q_19__14), .QB (\$dummy [355]), .D (
         nx5423), .CLK (nx7162), .R (reset)) ;
    mux21_ni ix5424 (.Y (nx5423), .A0 (q_19__14), .A1 (q_18__14), .S0 (nx7044)
             ) ;
    dffr gen_regs_18_regi_reg_q_14 (.Q (q_18__14), .QB (\$dummy [356]), .D (
         nx5413), .CLK (nx7162), .R (reset)) ;
    mux21_ni ix5414 (.Y (nx5413), .A0 (q_18__14), .A1 (q_17__14), .S0 (nx7044)
             ) ;
    dffr gen_regs_17_regi_reg_q_14 (.Q (q_17__14), .QB (\$dummy [357]), .D (
         nx5403), .CLK (nx7162), .R (reset)) ;
    mux21_ni ix5404 (.Y (nx5403), .A0 (q_17__14), .A1 (q_16__14), .S0 (nx7044)
             ) ;
    dffr gen_regs_16_regi_reg_q_14 (.Q (q_16__14), .QB (\$dummy [358]), .D (
         nx5393), .CLK (nx7162), .R (reset)) ;
    mux21_ni ix5394 (.Y (nx5393), .A0 (q_16__14), .A1 (q_15__14), .S0 (nx7044)
             ) ;
    dffr gen_regs_15_regi_reg_q_14 (.Q (q_15__14), .QB (\$dummy [359]), .D (
         nx5383), .CLK (nx7162), .R (reset)) ;
    mux21_ni ix5384 (.Y (nx5383), .A0 (q_15__14), .A1 (q_14__14), .S0 (nx7044)
             ) ;
    dffr gen_regs_14_regi_reg_q_14 (.Q (q_14__14), .QB (\$dummy [360]), .D (
         nx5373), .CLK (nx7162), .R (reset)) ;
    mux21_ni ix5374 (.Y (nx5373), .A0 (q_14__14), .A1 (q_13__14), .S0 (nx7044)
             ) ;
    dffr gen_regs_13_regi_reg_q_14 (.Q (q_13__14), .QB (\$dummy [361]), .D (
         nx5363), .CLK (nx7160), .R (reset)) ;
    mux21_ni ix5364 (.Y (nx5363), .A0 (q_13__14), .A1 (q_12__14), .S0 (nx7042)
             ) ;
    dffr gen_regs_12_regi_reg_q_14 (.Q (q_12__14), .QB (\$dummy [362]), .D (
         nx5353), .CLK (nx7160), .R (reset)) ;
    mux21_ni ix5354 (.Y (nx5353), .A0 (q_12__14), .A1 (q_11__14), .S0 (nx7042)
             ) ;
    dffr gen_regs_11_regi_reg_q_14 (.Q (q_11__14), .QB (\$dummy [363]), .D (
         nx5343), .CLK (nx7160), .R (reset)) ;
    mux21_ni ix5344 (.Y (nx5343), .A0 (q_11__14), .A1 (q_10__14), .S0 (nx7042)
             ) ;
    dffr gen_regs_10_regi_reg_q_14 (.Q (q_10__14), .QB (\$dummy [364]), .D (
         nx5333), .CLK (nx7160), .R (reset)) ;
    mux21_ni ix5334 (.Y (nx5333), .A0 (q_10__14), .A1 (q_9__14), .S0 (nx7042)) ;
    dffr gen_regs_9_regi_reg_q_14 (.Q (q_9__14), .QB (\$dummy [365]), .D (nx5323
         ), .CLK (nx7160), .R (reset)) ;
    mux21_ni ix5324 (.Y (nx5323), .A0 (q_9__14), .A1 (q_8__14), .S0 (nx7042)) ;
    dffr gen_regs_8_regi_reg_q_14 (.Q (q_8__14), .QB (\$dummy [366]), .D (nx5313
         ), .CLK (nx7160), .R (reset)) ;
    mux21_ni ix5314 (.Y (nx5313), .A0 (q_8__14), .A1 (q_7__14), .S0 (nx7042)) ;
    dffr gen_regs_7_regi_reg_q_14 (.Q (q_7__14), .QB (\$dummy [367]), .D (nx5303
         ), .CLK (nx7160), .R (reset)) ;
    mux21_ni ix5304 (.Y (nx5303), .A0 (q_7__14), .A1 (q_6__14), .S0 (nx7042)) ;
    dffr gen_regs_6_regi_reg_q_14 (.Q (q_6__14), .QB (\$dummy [368]), .D (nx5293
         ), .CLK (nx7158), .R (reset)) ;
    mux21_ni ix5294 (.Y (nx5293), .A0 (q_6__14), .A1 (q_5__14), .S0 (nx7040)) ;
    dffr gen_regs_5_regi_reg_q_14 (.Q (q_5__14), .QB (\$dummy [369]), .D (nx5283
         ), .CLK (nx7158), .R (reset)) ;
    mux21_ni ix5284 (.Y (nx5283), .A0 (q_5__14), .A1 (q_4__14), .S0 (nx7040)) ;
    dffr gen_regs_4_regi_reg_q_14 (.Q (q_4__14), .QB (\$dummy [370]), .D (nx5273
         ), .CLK (nx7158), .R (reset)) ;
    mux21_ni ix5274 (.Y (nx5273), .A0 (q_4__14), .A1 (q_3__14), .S0 (nx7040)) ;
    dffr gen_regs_3_regi_reg_q_14 (.Q (q_3__14), .QB (\$dummy [371]), .D (nx5263
         ), .CLK (nx7158), .R (reset)) ;
    mux21_ni ix5264 (.Y (nx5263), .A0 (q_3__14), .A1 (q_2__14), .S0 (nx7040)) ;
    dffr gen_regs_2_regi_reg_q_14 (.Q (q_2__14), .QB (\$dummy [372]), .D (nx5253
         ), .CLK (nx7158), .R (reset)) ;
    mux21_ni ix5254 (.Y (nx5253), .A0 (q_2__14), .A1 (q_1__14), .S0 (nx7040)) ;
    dffr gen_regs_1_regi_reg_q_14 (.Q (q_1__14), .QB (\$dummy [373]), .D (nx5243
         ), .CLK (nx7158), .R (reset)) ;
    mux21_ni ix5244 (.Y (nx5243), .A0 (q_1__14), .A1 (q_0__14), .S0 (nx7040)) ;
    dffr reg0_reg_q_14 (.Q (q_0__14), .QB (\$dummy [374]), .D (nx5233), .CLK (
         nx7158), .R (reset)) ;
    mux21_ni ix5234 (.Y (nx5233), .A0 (q_0__14), .A1 (d[14]), .S0 (nx7040)) ;
    dffr gen_regs_24_regi_reg_q_15 (.Q (q_24__15), .QB (\$dummy [375]), .D (
         nx5723), .CLK (nx7172), .R (reset)) ;
    mux21_ni ix5724 (.Y (nx5723), .A0 (q_24__15), .A1 (q_23__15), .S0 (nx7054)
             ) ;
    dffr gen_regs_23_regi_reg_q_15 (.Q (q_23__15), .QB (\$dummy [376]), .D (
         nx5713), .CLK (nx7170), .R (reset)) ;
    mux21_ni ix5714 (.Y (nx5713), .A0 (q_23__15), .A1 (q_22__15), .S0 (nx7052)
             ) ;
    dffr gen_regs_22_regi_reg_q_15 (.Q (q_22__15), .QB (\$dummy [377]), .D (
         nx5703), .CLK (nx7170), .R (reset)) ;
    mux21_ni ix5704 (.Y (nx5703), .A0 (q_22__15), .A1 (q_21__15), .S0 (nx7052)
             ) ;
    dffr gen_regs_21_regi_reg_q_15 (.Q (q_21__15), .QB (\$dummy [378]), .D (
         nx5693), .CLK (nx7170), .R (reset)) ;
    mux21_ni ix5694 (.Y (nx5693), .A0 (q_21__15), .A1 (q_20__15), .S0 (nx7052)
             ) ;
    dffr gen_regs_20_regi_reg_q_15 (.Q (q_20__15), .QB (\$dummy [379]), .D (
         nx5683), .CLK (nx7170), .R (reset)) ;
    mux21_ni ix5684 (.Y (nx5683), .A0 (q_20__15), .A1 (q_19__15), .S0 (nx7052)
             ) ;
    dffr gen_regs_19_regi_reg_q_15 (.Q (q_19__15), .QB (\$dummy [380]), .D (
         nx5673), .CLK (nx7170), .R (reset)) ;
    mux21_ni ix5674 (.Y (nx5673), .A0 (q_19__15), .A1 (q_18__15), .S0 (nx7052)
             ) ;
    dffr gen_regs_18_regi_reg_q_15 (.Q (q_18__15), .QB (\$dummy [381]), .D (
         nx5663), .CLK (nx7170), .R (reset)) ;
    mux21_ni ix5664 (.Y (nx5663), .A0 (q_18__15), .A1 (q_17__15), .S0 (nx7052)
             ) ;
    dffr gen_regs_17_regi_reg_q_15 (.Q (q_17__15), .QB (\$dummy [382]), .D (
         nx5653), .CLK (nx7170), .R (reset)) ;
    mux21_ni ix5654 (.Y (nx5653), .A0 (q_17__15), .A1 (q_16__15), .S0 (nx7052)
             ) ;
    dffr gen_regs_16_regi_reg_q_15 (.Q (q_16__15), .QB (\$dummy [383]), .D (
         nx5643), .CLK (nx7168), .R (reset)) ;
    mux21_ni ix5644 (.Y (nx5643), .A0 (q_16__15), .A1 (q_15__15), .S0 (nx7050)
             ) ;
    dffr gen_regs_15_regi_reg_q_15 (.Q (q_15__15), .QB (\$dummy [384]), .D (
         nx5633), .CLK (nx7168), .R (reset)) ;
    mux21_ni ix5634 (.Y (nx5633), .A0 (q_15__15), .A1 (q_14__15), .S0 (nx7050)
             ) ;
    dffr gen_regs_14_regi_reg_q_15 (.Q (q_14__15), .QB (\$dummy [385]), .D (
         nx5623), .CLK (nx7168), .R (reset)) ;
    mux21_ni ix5624 (.Y (nx5623), .A0 (q_14__15), .A1 (q_13__15), .S0 (nx7050)
             ) ;
    dffr gen_regs_13_regi_reg_q_15 (.Q (q_13__15), .QB (\$dummy [386]), .D (
         nx5613), .CLK (nx7168), .R (reset)) ;
    mux21_ni ix5614 (.Y (nx5613), .A0 (q_13__15), .A1 (q_12__15), .S0 (nx7050)
             ) ;
    dffr gen_regs_12_regi_reg_q_15 (.Q (q_12__15), .QB (\$dummy [387]), .D (
         nx5603), .CLK (nx7168), .R (reset)) ;
    mux21_ni ix5604 (.Y (nx5603), .A0 (q_12__15), .A1 (q_11__15), .S0 (nx7050)
             ) ;
    dffr gen_regs_11_regi_reg_q_15 (.Q (q_11__15), .QB (\$dummy [388]), .D (
         nx5593), .CLK (nx7168), .R (reset)) ;
    mux21_ni ix5594 (.Y (nx5593), .A0 (q_11__15), .A1 (q_10__15), .S0 (nx7050)
             ) ;
    dffr gen_regs_10_regi_reg_q_15 (.Q (q_10__15), .QB (\$dummy [389]), .D (
         nx5583), .CLK (nx7168), .R (reset)) ;
    mux21_ni ix5584 (.Y (nx5583), .A0 (q_10__15), .A1 (q_9__15), .S0 (nx7050)) ;
    dffr gen_regs_9_regi_reg_q_15 (.Q (q_9__15), .QB (\$dummy [390]), .D (nx5573
         ), .CLK (nx7166), .R (reset)) ;
    mux21_ni ix5574 (.Y (nx5573), .A0 (q_9__15), .A1 (q_8__15), .S0 (nx7048)) ;
    dffr gen_regs_8_regi_reg_q_15 (.Q (q_8__15), .QB (\$dummy [391]), .D (nx5563
         ), .CLK (nx7166), .R (reset)) ;
    mux21_ni ix5564 (.Y (nx5563), .A0 (q_8__15), .A1 (q_7__15), .S0 (nx7048)) ;
    dffr gen_regs_7_regi_reg_q_15 (.Q (q_7__15), .QB (\$dummy [392]), .D (nx5553
         ), .CLK (nx7166), .R (reset)) ;
    mux21_ni ix5554 (.Y (nx5553), .A0 (q_7__15), .A1 (q_6__15), .S0 (nx7048)) ;
    dffr gen_regs_6_regi_reg_q_15 (.Q (q_6__15), .QB (\$dummy [393]), .D (nx5543
         ), .CLK (nx7166), .R (reset)) ;
    mux21_ni ix5544 (.Y (nx5543), .A0 (q_6__15), .A1 (q_5__15), .S0 (nx7048)) ;
    dffr gen_regs_5_regi_reg_q_15 (.Q (q_5__15), .QB (\$dummy [394]), .D (nx5533
         ), .CLK (nx7166), .R (reset)) ;
    mux21_ni ix5534 (.Y (nx5533), .A0 (q_5__15), .A1 (q_4__15), .S0 (nx7048)) ;
    dffr gen_regs_4_regi_reg_q_15 (.Q (q_4__15), .QB (\$dummy [395]), .D (nx5523
         ), .CLK (nx7166), .R (reset)) ;
    mux21_ni ix5524 (.Y (nx5523), .A0 (q_4__15), .A1 (q_3__15), .S0 (nx7048)) ;
    dffr gen_regs_3_regi_reg_q_15 (.Q (q_3__15), .QB (\$dummy [396]), .D (nx5513
         ), .CLK (nx7166), .R (reset)) ;
    mux21_ni ix5514 (.Y (nx5513), .A0 (q_3__15), .A1 (q_2__15), .S0 (nx7048)) ;
    dffr gen_regs_2_regi_reg_q_15 (.Q (q_2__15), .QB (\$dummy [397]), .D (nx5503
         ), .CLK (nx7164), .R (reset)) ;
    mux21_ni ix5504 (.Y (nx5503), .A0 (q_2__15), .A1 (q_1__15), .S0 (nx7046)) ;
    dffr gen_regs_1_regi_reg_q_15 (.Q (q_1__15), .QB (\$dummy [398]), .D (nx5493
         ), .CLK (nx7164), .R (reset)) ;
    mux21_ni ix5494 (.Y (nx5493), .A0 (q_1__15), .A1 (q_0__15), .S0 (nx7046)) ;
    dffr reg0_reg_q_15 (.Q (q_0__15), .QB (\$dummy [399]), .D (nx5483), .CLK (
         nx7164), .R (reset)) ;
    mux21_ni ix5484 (.Y (nx5483), .A0 (q_0__15), .A1 (d[15]), .S0 (nx7046)) ;
    inv02 ix6939 (.Y (nx6940), .A (nx7626)) ;
    inv02 ix6941 (.Y (nx6942), .A (nx7626)) ;
    inv02 ix6943 (.Y (nx6944), .A (nx7626)) ;
    inv02 ix6945 (.Y (nx6946), .A (nx7626)) ;
    inv02 ix6947 (.Y (nx6948), .A (nx7626)) ;
    inv02 ix6949 (.Y (nx6950), .A (nx7626)) ;
    inv02 ix6951 (.Y (nx6952), .A (nx7174)) ;
    inv02 ix6953 (.Y (nx6954), .A (nx7176)) ;
    inv02 ix6955 (.Y (nx6956), .A (nx7176)) ;
    inv02 ix6957 (.Y (nx6958), .A (nx7176)) ;
    inv02 ix6959 (.Y (nx6960), .A (nx7176)) ;
    inv02 ix6961 (.Y (nx6962), .A (nx7176)) ;
    inv02 ix6963 (.Y (nx6964), .A (nx7176)) ;
    inv02 ix6965 (.Y (nx6966), .A (nx7176)) ;
    inv02 ix6967 (.Y (nx6968), .A (nx7178)) ;
    inv02 ix6969 (.Y (nx6970), .A (nx7178)) ;
    inv02 ix6971 (.Y (nx6972), .A (nx7178)) ;
    inv02 ix6973 (.Y (nx6974), .A (nx7178)) ;
    inv02 ix6975 (.Y (nx6976), .A (nx7178)) ;
    inv02 ix6977 (.Y (nx6978), .A (nx7178)) ;
    inv02 ix6979 (.Y (nx6980), .A (nx7178)) ;
    inv02 ix6981 (.Y (nx6982), .A (nx7180)) ;
    inv02 ix6983 (.Y (nx6984), .A (nx7180)) ;
    inv02 ix6985 (.Y (nx6986), .A (nx7180)) ;
    inv02 ix6987 (.Y (nx6988), .A (nx7180)) ;
    inv02 ix6989 (.Y (nx6990), .A (nx7180)) ;
    inv02 ix6991 (.Y (nx6992), .A (nx7180)) ;
    inv02 ix6993 (.Y (nx6994), .A (nx7180)) ;
    inv02 ix6995 (.Y (nx6996), .A (nx7182)) ;
    inv02 ix6997 (.Y (nx6998), .A (nx7182)) ;
    inv02 ix6999 (.Y (nx7000), .A (nx7182)) ;
    inv02 ix7001 (.Y (nx7002), .A (nx7182)) ;
    inv02 ix7003 (.Y (nx7004), .A (nx7182)) ;
    inv02 ix7005 (.Y (nx7006), .A (nx7182)) ;
    inv02 ix7007 (.Y (nx7008), .A (nx7182)) ;
    inv02 ix7009 (.Y (nx7010), .A (nx7184)) ;
    inv02 ix7011 (.Y (nx7012), .A (nx7184)) ;
    inv02 ix7013 (.Y (nx7014), .A (nx7184)) ;
    inv02 ix7015 (.Y (nx7016), .A (nx7184)) ;
    inv02 ix7017 (.Y (nx7018), .A (nx7184)) ;
    inv02 ix7019 (.Y (nx7020), .A (nx7184)) ;
    inv02 ix7021 (.Y (nx7022), .A (nx7184)) ;
    inv02 ix7023 (.Y (nx7024), .A (nx7186)) ;
    inv02 ix7025 (.Y (nx7026), .A (nx7186)) ;
    inv02 ix7027 (.Y (nx7028), .A (nx7186)) ;
    inv02 ix7029 (.Y (nx7030), .A (nx7186)) ;
    inv02 ix7031 (.Y (nx7032), .A (nx7186)) ;
    inv02 ix7033 (.Y (nx7034), .A (nx7186)) ;
    inv02 ix7035 (.Y (nx7036), .A (nx7186)) ;
    inv02 ix7037 (.Y (nx7038), .A (nx7188)) ;
    inv02 ix7039 (.Y (nx7040), .A (nx7188)) ;
    inv02 ix7041 (.Y (nx7042), .A (nx7188)) ;
    inv02 ix7043 (.Y (nx7044), .A (nx7188)) ;
    inv02 ix7045 (.Y (nx7046), .A (nx7188)) ;
    inv02 ix7047 (.Y (nx7048), .A (nx7188)) ;
    inv02 ix7049 (.Y (nx7050), .A (nx7188)) ;
    inv02 ix7051 (.Y (nx7052), .A (nx7190)) ;
    inv02 ix7053 (.Y (nx7054), .A (nx7190)) ;
    inv02 ix7057 (.Y (nx7058), .A (nx7628)) ;
    inv02 ix7059 (.Y (nx7060), .A (nx7628)) ;
    inv02 ix7061 (.Y (nx7062), .A (nx7628)) ;
    inv02 ix7063 (.Y (nx7064), .A (nx7628)) ;
    inv02 ix7065 (.Y (nx7066), .A (nx7628)) ;
    inv02 ix7067 (.Y (nx7068), .A (nx7628)) ;
    inv02 ix7069 (.Y (nx7070), .A (nx7192)) ;
    inv02 ix7071 (.Y (nx7072), .A (nx7194)) ;
    inv02 ix7073 (.Y (nx7074), .A (nx7194)) ;
    inv02 ix7075 (.Y (nx7076), .A (nx7194)) ;
    inv02 ix7077 (.Y (nx7078), .A (nx7194)) ;
    inv02 ix7079 (.Y (nx7080), .A (nx7194)) ;
    inv02 ix7081 (.Y (nx7082), .A (nx7194)) ;
    inv02 ix7083 (.Y (nx7084), .A (nx7194)) ;
    inv02 ix7085 (.Y (nx7086), .A (nx7196)) ;
    inv02 ix7087 (.Y (nx7088), .A (nx7196)) ;
    inv02 ix7089 (.Y (nx7090), .A (nx7196)) ;
    inv02 ix7091 (.Y (nx7092), .A (nx7196)) ;
    inv02 ix7093 (.Y (nx7094), .A (nx7196)) ;
    inv02 ix7095 (.Y (nx7096), .A (nx7196)) ;
    inv02 ix7097 (.Y (nx7098), .A (nx7196)) ;
    inv02 ix7099 (.Y (nx7100), .A (nx7198)) ;
    inv02 ix7101 (.Y (nx7102), .A (nx7198)) ;
    inv02 ix7103 (.Y (nx7104), .A (nx7198)) ;
    inv02 ix7105 (.Y (nx7106), .A (nx7198)) ;
    inv02 ix7107 (.Y (nx7108), .A (nx7198)) ;
    inv02 ix7109 (.Y (nx7110), .A (nx7198)) ;
    inv02 ix7111 (.Y (nx7112), .A (nx7198)) ;
    inv02 ix7113 (.Y (nx7114), .A (nx7200)) ;
    inv02 ix7115 (.Y (nx7116), .A (nx7200)) ;
    inv02 ix7117 (.Y (nx7118), .A (nx7200)) ;
    inv02 ix7119 (.Y (nx7120), .A (nx7200)) ;
    inv02 ix7121 (.Y (nx7122), .A (nx7200)) ;
    inv02 ix7123 (.Y (nx7124), .A (nx7200)) ;
    inv02 ix7125 (.Y (nx7126), .A (nx7200)) ;
    inv02 ix7127 (.Y (nx7128), .A (nx7202)) ;
    inv02 ix7129 (.Y (nx7130), .A (nx7202)) ;
    inv02 ix7131 (.Y (nx7132), .A (nx7202)) ;
    inv02 ix7133 (.Y (nx7134), .A (nx7202)) ;
    inv02 ix7135 (.Y (nx7136), .A (nx7202)) ;
    inv02 ix7137 (.Y (nx7138), .A (nx7202)) ;
    inv02 ix7139 (.Y (nx7140), .A (nx7202)) ;
    inv02 ix7141 (.Y (nx7142), .A (nx7204)) ;
    inv02 ix7143 (.Y (nx7144), .A (nx7204)) ;
    inv02 ix7145 (.Y (nx7146), .A (nx7204)) ;
    inv02 ix7147 (.Y (nx7148), .A (nx7204)) ;
    inv02 ix7149 (.Y (nx7150), .A (nx7204)) ;
    inv02 ix7151 (.Y (nx7152), .A (nx7204)) ;
    inv02 ix7153 (.Y (nx7154), .A (nx7204)) ;
    inv02 ix7155 (.Y (nx7156), .A (nx7206)) ;
    inv02 ix7157 (.Y (nx7158), .A (nx7206)) ;
    inv02 ix7159 (.Y (nx7160), .A (nx7206)) ;
    inv02 ix7161 (.Y (nx7162), .A (nx7206)) ;
    inv02 ix7163 (.Y (nx7164), .A (nx7206)) ;
    inv02 ix7165 (.Y (nx7166), .A (nx7206)) ;
    inv02 ix7167 (.Y (nx7168), .A (nx7206)) ;
    inv02 ix7169 (.Y (nx7170), .A (nx7208)) ;
    inv02 ix7171 (.Y (nx7172), .A (nx7208)) ;
    inv02 ix7173 (.Y (nx7174), .A (load)) ;
    inv02 ix7175 (.Y (nx7176), .A (nx7214)) ;
    inv02 ix7177 (.Y (nx7178), .A (nx7214)) ;
    inv02 ix7179 (.Y (nx7180), .A (nx7214)) ;
    inv02 ix7181 (.Y (nx7182), .A (nx7214)) ;
    inv02 ix7183 (.Y (nx7184), .A (nx7214)) ;
    inv02 ix7185 (.Y (nx7186), .A (nx7216)) ;
    inv02 ix7187 (.Y (nx7188), .A (nx7216)) ;
    inv02 ix7189 (.Y (nx7190), .A (nx7216)) ;
    inv02 ix7191 (.Y (nx7192), .A (clk)) ;
    inv02 ix7193 (.Y (nx7194), .A (nx7218)) ;
    inv02 ix7195 (.Y (nx7196), .A (nx7218)) ;
    inv02 ix7197 (.Y (nx7198), .A (nx7218)) ;
    inv02 ix7199 (.Y (nx7200), .A (nx7218)) ;
    inv02 ix7201 (.Y (nx7202), .A (nx7218)) ;
    inv02 ix7203 (.Y (nx7204), .A (nx7220)) ;
    inv02 ix7205 (.Y (nx7206), .A (nx7220)) ;
    inv02 ix7207 (.Y (nx7208), .A (nx7220)) ;
    inv01 ix7213 (.Y (nx7214), .A (nx7626)) ;
    inv01 ix7215 (.Y (nx7216), .A (nx7174)) ;
    inv01 ix7217 (.Y (nx7218), .A (nx7628)) ;
    inv01 ix7219 (.Y (nx7220), .A (nx7192)) ;
    inv02 ix7625 (.Y (nx7626), .A (load)) ;
    inv02 ix7627 (.Y (nx7628), .A (clk)) ;
endmodule


module Queue_5_unfolded2 ( d, q_0__15, q_0__14, q_0__13, q_0__12, q_0__11, 
                           q_0__10, q_0__9, q_0__8, q_0__7, q_0__6, q_0__5, 
                           q_0__4, q_0__3, q_0__2, q_0__1, q_0__0, q_1__15, 
                           q_1__14, q_1__13, q_1__12, q_1__11, q_1__10, q_1__9, 
                           q_1__8, q_1__7, q_1__6, q_1__5, q_1__4, q_1__3, 
                           q_1__2, q_1__1, q_1__0, q_2__15, q_2__14, q_2__13, 
                           q_2__12, q_2__11, q_2__10, q_2__9, q_2__8, q_2__7, 
                           q_2__6, q_2__5, q_2__4, q_2__3, q_2__2, q_2__1, 
                           q_2__0, q_3__15, q_3__14, q_3__13, q_3__12, q_3__11, 
                           q_3__10, q_3__9, q_3__8, q_3__7, q_3__6, q_3__5, 
                           q_3__4, q_3__3, q_3__2, q_3__1, q_3__0, q_4__15, 
                           q_4__14, q_4__13, q_4__12, q_4__11, q_4__10, q_4__9, 
                           q_4__8, q_4__7, q_4__6, q_4__5, q_4__4, q_4__3, 
                           q_4__2, q_4__1, q_4__0, clk, load, reset ) ;

    input [15:0]d ;
    output q_0__15 ;
    output q_0__14 ;
    output q_0__13 ;
    output q_0__12 ;
    output q_0__11 ;
    output q_0__10 ;
    output q_0__9 ;
    output q_0__8 ;
    output q_0__7 ;
    output q_0__6 ;
    output q_0__5 ;
    output q_0__4 ;
    output q_0__3 ;
    output q_0__2 ;
    output q_0__1 ;
    output q_0__0 ;
    output q_1__15 ;
    output q_1__14 ;
    output q_1__13 ;
    output q_1__12 ;
    output q_1__11 ;
    output q_1__10 ;
    output q_1__9 ;
    output q_1__8 ;
    output q_1__7 ;
    output q_1__6 ;
    output q_1__5 ;
    output q_1__4 ;
    output q_1__3 ;
    output q_1__2 ;
    output q_1__1 ;
    output q_1__0 ;
    output q_2__15 ;
    output q_2__14 ;
    output q_2__13 ;
    output q_2__12 ;
    output q_2__11 ;
    output q_2__10 ;
    output q_2__9 ;
    output q_2__8 ;
    output q_2__7 ;
    output q_2__6 ;
    output q_2__5 ;
    output q_2__4 ;
    output q_2__3 ;
    output q_2__2 ;
    output q_2__1 ;
    output q_2__0 ;
    output q_3__15 ;
    output q_3__14 ;
    output q_3__13 ;
    output q_3__12 ;
    output q_3__11 ;
    output q_3__10 ;
    output q_3__9 ;
    output q_3__8 ;
    output q_3__7 ;
    output q_3__6 ;
    output q_3__5 ;
    output q_3__4 ;
    output q_3__3 ;
    output q_3__2 ;
    output q_3__1 ;
    output q_3__0 ;
    output q_4__15 ;
    output q_4__14 ;
    output q_4__13 ;
    output q_4__12 ;
    output q_4__11 ;
    output q_4__10 ;
    output q_4__9 ;
    output q_4__8 ;
    output q_4__7 ;
    output q_4__6 ;
    output q_4__5 ;
    output q_4__4 ;
    output q_4__3 ;
    output q_4__2 ;
    output q_4__1 ;
    output q_4__0 ;
    input clk ;
    input load ;
    input reset ;

    wire nx240, nx250, nx260, nx270, nx280, nx290, nx300, nx310, nx320, nx330, 
         nx340, nx350, nx360, nx370, nx380, nx390, nx400, nx410, nx420, nx430, 
         nx440, nx450, nx460, nx470, nx480, nx490, nx500, nx510, nx520, nx530, 
         nx540, nx550, nx560, nx570, nx580, nx590, nx600, nx610, nx620, nx630, 
         nx640, nx650, nx660, nx670, nx680, nx690, nx700, nx710, nx720, nx730, 
         nx740, nx750, nx760, nx770, nx780, nx790, nx800, nx810, nx820, nx830, 
         nx840, nx850, nx860, nx870, nx880, nx890, nx900, nx910, nx920, nx930, 
         nx940, nx950, nx960, nx970, nx980, nx990, nx1000, nx1010, nx1020, 
         nx1030, nx1287, nx1289, nx1291, nx1293, nx1295, nx1297, nx1299, nx1301, 
         nx1303, nx1305, nx1307, nx1309, nx1313, nx1315, nx1317, nx1319, nx1321, 
         nx1323, nx1325, nx1327, nx1329, nx1331, nx1333, nx1335, nx1337, nx1339, 
         nx1341, nx1343;
    wire [79:0] \$dummy ;




    dff gen_regs_4_regi_reg_q_0 (.Q (q_4__0), .QB (\$dummy [0]), .D (nx280), .CLK (
        nx1313)) ;
    mux21_ni ix281 (.Y (nx280), .A0 (q_4__0), .A1 (q_3__0), .S0 (nx1287)) ;
    dff gen_regs_3_regi_reg_q_0 (.Q (q_3__0), .QB (\$dummy [1]), .D (nx270), .CLK (
        nx1313)) ;
    mux21_ni ix271 (.Y (nx270), .A0 (q_3__0), .A1 (q_2__0), .S0 (nx1287)) ;
    dff gen_regs_2_regi_reg_q_0 (.Q (q_2__0), .QB (\$dummy [2]), .D (nx260), .CLK (
        nx1313)) ;
    mux21_ni ix261 (.Y (nx260), .A0 (q_2__0), .A1 (q_1__0), .S0 (nx1287)) ;
    dff gen_regs_1_regi_reg_q_0 (.Q (q_1__0), .QB (\$dummy [3]), .D (nx250), .CLK (
        nx1313)) ;
    mux21_ni ix251 (.Y (nx250), .A0 (q_1__0), .A1 (q_0__0), .S0 (nx1287)) ;
    dff reg0_reg_q_0 (.Q (q_0__0), .QB (\$dummy [4]), .D (nx240), .CLK (nx1313)
        ) ;
    mux21_ni ix241 (.Y (nx240), .A0 (q_0__0), .A1 (d[0]), .S0 (nx1287)) ;
    dff gen_regs_4_regi_reg_q_1 (.Q (q_4__1), .QB (\$dummy [5]), .D (nx330), .CLK (
        nx1315)) ;
    mux21_ni ix331 (.Y (nx330), .A0 (q_4__1), .A1 (q_3__1), .S0 (nx1289)) ;
    dff gen_regs_3_regi_reg_q_1 (.Q (q_3__1), .QB (\$dummy [6]), .D (nx320), .CLK (
        nx1315)) ;
    mux21_ni ix321 (.Y (nx320), .A0 (q_3__1), .A1 (q_2__1), .S0 (nx1289)) ;
    dff gen_regs_2_regi_reg_q_1 (.Q (q_2__1), .QB (\$dummy [7]), .D (nx310), .CLK (
        nx1315)) ;
    mux21_ni ix311 (.Y (nx310), .A0 (q_2__1), .A1 (q_1__1), .S0 (nx1289)) ;
    dff gen_regs_1_regi_reg_q_1 (.Q (q_1__1), .QB (\$dummy [8]), .D (nx300), .CLK (
        nx1313)) ;
    mux21_ni ix301 (.Y (nx300), .A0 (q_1__1), .A1 (q_0__1), .S0 (nx1287)) ;
    dff reg0_reg_q_1 (.Q (q_0__1), .QB (\$dummy [9]), .D (nx290), .CLK (nx1313)
        ) ;
    mux21_ni ix291 (.Y (nx290), .A0 (q_0__1), .A1 (d[1]), .S0 (nx1287)) ;
    dff gen_regs_4_regi_reg_q_2 (.Q (q_4__2), .QB (\$dummy [10]), .D (nx380), .CLK (
        nx1317)) ;
    mux21_ni ix381 (.Y (nx380), .A0 (q_4__2), .A1 (q_3__2), .S0 (nx1291)) ;
    dff gen_regs_3_regi_reg_q_2 (.Q (q_3__2), .QB (\$dummy [11]), .D (nx370), .CLK (
        nx1315)) ;
    mux21_ni ix371 (.Y (nx370), .A0 (q_3__2), .A1 (q_2__2), .S0 (nx1289)) ;
    dff gen_regs_2_regi_reg_q_2 (.Q (q_2__2), .QB (\$dummy [12]), .D (nx360), .CLK (
        nx1315)) ;
    mux21_ni ix361 (.Y (nx360), .A0 (q_2__2), .A1 (q_1__2), .S0 (nx1289)) ;
    dff gen_regs_1_regi_reg_q_2 (.Q (q_1__2), .QB (\$dummy [13]), .D (nx350), .CLK (
        nx1315)) ;
    mux21_ni ix351 (.Y (nx350), .A0 (q_1__2), .A1 (q_0__2), .S0 (nx1289)) ;
    dff reg0_reg_q_2 (.Q (q_0__2), .QB (\$dummy [14]), .D (nx340), .CLK (nx1315)
        ) ;
    mux21_ni ix341 (.Y (nx340), .A0 (q_0__2), .A1 (d[2]), .S0 (nx1289)) ;
    dff gen_regs_4_regi_reg_q_3 (.Q (q_4__3), .QB (\$dummy [15]), .D (nx430), .CLK (
        nx1317)) ;
    mux21_ni ix431 (.Y (nx430), .A0 (q_4__3), .A1 (q_3__3), .S0 (nx1291)) ;
    dff gen_regs_3_regi_reg_q_3 (.Q (q_3__3), .QB (\$dummy [16]), .D (nx420), .CLK (
        nx1317)) ;
    mux21_ni ix421 (.Y (nx420), .A0 (q_3__3), .A1 (q_2__3), .S0 (nx1291)) ;
    dff gen_regs_2_regi_reg_q_3 (.Q (q_2__3), .QB (\$dummy [17]), .D (nx410), .CLK (
        nx1317)) ;
    mux21_ni ix411 (.Y (nx410), .A0 (q_2__3), .A1 (q_1__3), .S0 (nx1291)) ;
    dff gen_regs_1_regi_reg_q_3 (.Q (q_1__3), .QB (\$dummy [18]), .D (nx400), .CLK (
        nx1317)) ;
    mux21_ni ix401 (.Y (nx400), .A0 (q_1__3), .A1 (q_0__3), .S0 (nx1291)) ;
    dff reg0_reg_q_3 (.Q (q_0__3), .QB (\$dummy [19]), .D (nx390), .CLK (nx1317)
        ) ;
    mux21_ni ix391 (.Y (nx390), .A0 (q_0__3), .A1 (d[3]), .S0 (nx1291)) ;
    dff gen_regs_4_regi_reg_q_4 (.Q (q_4__4), .QB (\$dummy [20]), .D (nx480), .CLK (
        nx1319)) ;
    mux21_ni ix481 (.Y (nx480), .A0 (q_4__4), .A1 (q_3__4), .S0 (nx1293)) ;
    dff gen_regs_3_regi_reg_q_4 (.Q (q_3__4), .QB (\$dummy [21]), .D (nx470), .CLK (
        nx1319)) ;
    mux21_ni ix471 (.Y (nx470), .A0 (q_3__4), .A1 (q_2__4), .S0 (nx1293)) ;
    dff gen_regs_2_regi_reg_q_4 (.Q (q_2__4), .QB (\$dummy [22]), .D (nx460), .CLK (
        nx1319)) ;
    mux21_ni ix461 (.Y (nx460), .A0 (q_2__4), .A1 (q_1__4), .S0 (nx1293)) ;
    dff gen_regs_1_regi_reg_q_4 (.Q (q_1__4), .QB (\$dummy [23]), .D (nx450), .CLK (
        nx1319)) ;
    mux21_ni ix451 (.Y (nx450), .A0 (q_1__4), .A1 (q_0__4), .S0 (nx1293)) ;
    dff reg0_reg_q_4 (.Q (q_0__4), .QB (\$dummy [24]), .D (nx440), .CLK (nx1317)
        ) ;
    mux21_ni ix441 (.Y (nx440), .A0 (q_0__4), .A1 (d[4]), .S0 (nx1291)) ;
    dff gen_regs_4_regi_reg_q_5 (.Q (q_4__5), .QB (\$dummy [25]), .D (nx530), .CLK (
        nx1321)) ;
    mux21_ni ix531 (.Y (nx530), .A0 (q_4__5), .A1 (q_3__5), .S0 (nx1295)) ;
    dff gen_regs_3_regi_reg_q_5 (.Q (q_3__5), .QB (\$dummy [26]), .D (nx520), .CLK (
        nx1321)) ;
    mux21_ni ix521 (.Y (nx520), .A0 (q_3__5), .A1 (q_2__5), .S0 (nx1295)) ;
    dff gen_regs_2_regi_reg_q_5 (.Q (q_2__5), .QB (\$dummy [27]), .D (nx510), .CLK (
        nx1319)) ;
    mux21_ni ix511 (.Y (nx510), .A0 (q_2__5), .A1 (q_1__5), .S0 (nx1293)) ;
    dff gen_regs_1_regi_reg_q_5 (.Q (q_1__5), .QB (\$dummy [28]), .D (nx500), .CLK (
        nx1319)) ;
    mux21_ni ix501 (.Y (nx500), .A0 (q_1__5), .A1 (q_0__5), .S0 (nx1293)) ;
    dff reg0_reg_q_5 (.Q (q_0__5), .QB (\$dummy [29]), .D (nx490), .CLK (nx1319)
        ) ;
    mux21_ni ix491 (.Y (nx490), .A0 (q_0__5), .A1 (d[5]), .S0 (nx1293)) ;
    dff gen_regs_4_regi_reg_q_6 (.Q (q_4__6), .QB (\$dummy [30]), .D (nx580), .CLK (
        nx1321)) ;
    mux21_ni ix581 (.Y (nx580), .A0 (q_4__6), .A1 (q_3__6), .S0 (nx1295)) ;
    dff gen_regs_3_regi_reg_q_6 (.Q (q_3__6), .QB (\$dummy [31]), .D (nx570), .CLK (
        nx1321)) ;
    mux21_ni ix571 (.Y (nx570), .A0 (q_3__6), .A1 (q_2__6), .S0 (nx1295)) ;
    dff gen_regs_2_regi_reg_q_6 (.Q (q_2__6), .QB (\$dummy [32]), .D (nx560), .CLK (
        nx1321)) ;
    mux21_ni ix561 (.Y (nx560), .A0 (q_2__6), .A1 (q_1__6), .S0 (nx1295)) ;
    dff gen_regs_1_regi_reg_q_6 (.Q (q_1__6), .QB (\$dummy [33]), .D (nx550), .CLK (
        nx1321)) ;
    mux21_ni ix551 (.Y (nx550), .A0 (q_1__6), .A1 (q_0__6), .S0 (nx1295)) ;
    dff reg0_reg_q_6 (.Q (q_0__6), .QB (\$dummy [34]), .D (nx540), .CLK (nx1321)
        ) ;
    mux21_ni ix541 (.Y (nx540), .A0 (q_0__6), .A1 (d[6]), .S0 (nx1295)) ;
    dff gen_regs_4_regi_reg_q_7 (.Q (q_4__7), .QB (\$dummy [35]), .D (nx630), .CLK (
        nx1323)) ;
    mux21_ni ix631 (.Y (nx630), .A0 (q_4__7), .A1 (q_3__7), .S0 (nx1297)) ;
    dff gen_regs_3_regi_reg_q_7 (.Q (q_3__7), .QB (\$dummy [36]), .D (nx620), .CLK (
        nx1323)) ;
    mux21_ni ix621 (.Y (nx620), .A0 (q_3__7), .A1 (q_2__7), .S0 (nx1297)) ;
    dff gen_regs_2_regi_reg_q_7 (.Q (q_2__7), .QB (\$dummy [37]), .D (nx610), .CLK (
        nx1323)) ;
    mux21_ni ix611 (.Y (nx610), .A0 (q_2__7), .A1 (q_1__7), .S0 (nx1297)) ;
    dff gen_regs_1_regi_reg_q_7 (.Q (q_1__7), .QB (\$dummy [38]), .D (nx600), .CLK (
        nx1323)) ;
    mux21_ni ix601 (.Y (nx600), .A0 (q_1__7), .A1 (q_0__7), .S0 (nx1297)) ;
    dff reg0_reg_q_7 (.Q (q_0__7), .QB (\$dummy [39]), .D (nx590), .CLK (nx1323)
        ) ;
    mux21_ni ix591 (.Y (nx590), .A0 (q_0__7), .A1 (d[7]), .S0 (nx1297)) ;
    dff gen_regs_4_regi_reg_q_8 (.Q (q_4__8), .QB (\$dummy [40]), .D (nx680), .CLK (
        nx1325)) ;
    mux21_ni ix681 (.Y (nx680), .A0 (q_4__8), .A1 (q_3__8), .S0 (nx1299)) ;
    dff gen_regs_3_regi_reg_q_8 (.Q (q_3__8), .QB (\$dummy [41]), .D (nx670), .CLK (
        nx1325)) ;
    mux21_ni ix671 (.Y (nx670), .A0 (q_3__8), .A1 (q_2__8), .S0 (nx1299)) ;
    dff gen_regs_2_regi_reg_q_8 (.Q (q_2__8), .QB (\$dummy [42]), .D (nx660), .CLK (
        nx1325)) ;
    mux21_ni ix661 (.Y (nx660), .A0 (q_2__8), .A1 (q_1__8), .S0 (nx1299)) ;
    dff gen_regs_1_regi_reg_q_8 (.Q (q_1__8), .QB (\$dummy [43]), .D (nx650), .CLK (
        nx1323)) ;
    mux21_ni ix651 (.Y (nx650), .A0 (q_1__8), .A1 (q_0__8), .S0 (nx1297)) ;
    dff reg0_reg_q_8 (.Q (q_0__8), .QB (\$dummy [44]), .D (nx640), .CLK (nx1323)
        ) ;
    mux21_ni ix641 (.Y (nx640), .A0 (q_0__8), .A1 (d[8]), .S0 (nx1297)) ;
    dff gen_regs_4_regi_reg_q_9 (.Q (q_4__9), .QB (\$dummy [45]), .D (nx730), .CLK (
        nx1327)) ;
    mux21_ni ix731 (.Y (nx730), .A0 (q_4__9), .A1 (q_3__9), .S0 (nx1301)) ;
    dff gen_regs_3_regi_reg_q_9 (.Q (q_3__9), .QB (\$dummy [46]), .D (nx720), .CLK (
        nx1325)) ;
    mux21_ni ix721 (.Y (nx720), .A0 (q_3__9), .A1 (q_2__9), .S0 (nx1299)) ;
    dff gen_regs_2_regi_reg_q_9 (.Q (q_2__9), .QB (\$dummy [47]), .D (nx710), .CLK (
        nx1325)) ;
    mux21_ni ix711 (.Y (nx710), .A0 (q_2__9), .A1 (q_1__9), .S0 (nx1299)) ;
    dff gen_regs_1_regi_reg_q_9 (.Q (q_1__9), .QB (\$dummy [48]), .D (nx700), .CLK (
        nx1325)) ;
    mux21_ni ix701 (.Y (nx700), .A0 (q_1__9), .A1 (q_0__9), .S0 (nx1299)) ;
    dff reg0_reg_q_9 (.Q (q_0__9), .QB (\$dummy [49]), .D (nx690), .CLK (nx1325)
        ) ;
    mux21_ni ix691 (.Y (nx690), .A0 (q_0__9), .A1 (d[9]), .S0 (nx1299)) ;
    dff gen_regs_4_regi_reg_q_10 (.Q (q_4__10), .QB (\$dummy [50]), .D (nx780), 
        .CLK (nx1327)) ;
    mux21_ni ix781 (.Y (nx780), .A0 (q_4__10), .A1 (q_3__10), .S0 (nx1301)) ;
    dff gen_regs_3_regi_reg_q_10 (.Q (q_3__10), .QB (\$dummy [51]), .D (nx770), 
        .CLK (nx1327)) ;
    mux21_ni ix771 (.Y (nx770), .A0 (q_3__10), .A1 (q_2__10), .S0 (nx1301)) ;
    dff gen_regs_2_regi_reg_q_10 (.Q (q_2__10), .QB (\$dummy [52]), .D (nx760), 
        .CLK (nx1327)) ;
    mux21_ni ix761 (.Y (nx760), .A0 (q_2__10), .A1 (q_1__10), .S0 (nx1301)) ;
    dff gen_regs_1_regi_reg_q_10 (.Q (q_1__10), .QB (\$dummy [53]), .D (nx750), 
        .CLK (nx1327)) ;
    mux21_ni ix751 (.Y (nx750), .A0 (q_1__10), .A1 (q_0__10), .S0 (nx1301)) ;
    dff reg0_reg_q_10 (.Q (q_0__10), .QB (\$dummy [54]), .D (nx740), .CLK (
        nx1327)) ;
    mux21_ni ix741 (.Y (nx740), .A0 (q_0__10), .A1 (d[10]), .S0 (nx1301)) ;
    dff gen_regs_4_regi_reg_q_11 (.Q (q_4__11), .QB (\$dummy [55]), .D (nx830), 
        .CLK (nx1329)) ;
    mux21_ni ix831 (.Y (nx830), .A0 (q_4__11), .A1 (q_3__11), .S0 (nx1303)) ;
    dff gen_regs_3_regi_reg_q_11 (.Q (q_3__11), .QB (\$dummy [56]), .D (nx820), 
        .CLK (nx1329)) ;
    mux21_ni ix821 (.Y (nx820), .A0 (q_3__11), .A1 (q_2__11), .S0 (nx1303)) ;
    dff gen_regs_2_regi_reg_q_11 (.Q (q_2__11), .QB (\$dummy [57]), .D (nx810), 
        .CLK (nx1329)) ;
    mux21_ni ix811 (.Y (nx810), .A0 (q_2__11), .A1 (q_1__11), .S0 (nx1303)) ;
    dff gen_regs_1_regi_reg_q_11 (.Q (q_1__11), .QB (\$dummy [58]), .D (nx800), 
        .CLK (nx1329)) ;
    mux21_ni ix801 (.Y (nx800), .A0 (q_1__11), .A1 (q_0__11), .S0 (nx1303)) ;
    dff reg0_reg_q_11 (.Q (q_0__11), .QB (\$dummy [59]), .D (nx790), .CLK (
        nx1327)) ;
    mux21_ni ix791 (.Y (nx790), .A0 (q_0__11), .A1 (d[11]), .S0 (nx1301)) ;
    dff gen_regs_4_regi_reg_q_12 (.Q (q_4__12), .QB (\$dummy [60]), .D (nx880), 
        .CLK (nx1331)) ;
    mux21_ni ix881 (.Y (nx880), .A0 (q_4__12), .A1 (q_3__12), .S0 (nx1305)) ;
    dff gen_regs_3_regi_reg_q_12 (.Q (q_3__12), .QB (\$dummy [61]), .D (nx870), 
        .CLK (nx1331)) ;
    mux21_ni ix871 (.Y (nx870), .A0 (q_3__12), .A1 (q_2__12), .S0 (nx1305)) ;
    dff gen_regs_2_regi_reg_q_12 (.Q (q_2__12), .QB (\$dummy [62]), .D (nx860), 
        .CLK (nx1329)) ;
    mux21_ni ix861 (.Y (nx860), .A0 (q_2__12), .A1 (q_1__12), .S0 (nx1303)) ;
    dff gen_regs_1_regi_reg_q_12 (.Q (q_1__12), .QB (\$dummy [63]), .D (nx850), 
        .CLK (nx1329)) ;
    mux21_ni ix851 (.Y (nx850), .A0 (q_1__12), .A1 (q_0__12), .S0 (nx1303)) ;
    dff reg0_reg_q_12 (.Q (q_0__12), .QB (\$dummy [64]), .D (nx840), .CLK (
        nx1329)) ;
    mux21_ni ix841 (.Y (nx840), .A0 (q_0__12), .A1 (d[12]), .S0 (nx1303)) ;
    dff gen_regs_4_regi_reg_q_13 (.Q (q_4__13), .QB (\$dummy [65]), .D (nx930), 
        .CLK (nx1331)) ;
    mux21_ni ix931 (.Y (nx930), .A0 (q_4__13), .A1 (q_3__13), .S0 (nx1305)) ;
    dff gen_regs_3_regi_reg_q_13 (.Q (q_3__13), .QB (\$dummy [66]), .D (nx920), 
        .CLK (nx1331)) ;
    mux21_ni ix921 (.Y (nx920), .A0 (q_3__13), .A1 (q_2__13), .S0 (nx1305)) ;
    dff gen_regs_2_regi_reg_q_13 (.Q (q_2__13), .QB (\$dummy [67]), .D (nx910), 
        .CLK (nx1331)) ;
    mux21_ni ix911 (.Y (nx910), .A0 (q_2__13), .A1 (q_1__13), .S0 (nx1305)) ;
    dff gen_regs_1_regi_reg_q_13 (.Q (q_1__13), .QB (\$dummy [68]), .D (nx900), 
        .CLK (nx1331)) ;
    mux21_ni ix901 (.Y (nx900), .A0 (q_1__13), .A1 (q_0__13), .S0 (nx1305)) ;
    dff reg0_reg_q_13 (.Q (q_0__13), .QB (\$dummy [69]), .D (nx890), .CLK (
        nx1331)) ;
    mux21_ni ix891 (.Y (nx890), .A0 (q_0__13), .A1 (d[13]), .S0 (nx1305)) ;
    dff gen_regs_4_regi_reg_q_14 (.Q (q_4__14), .QB (\$dummy [70]), .D (nx980), 
        .CLK (nx1333)) ;
    mux21_ni ix981 (.Y (nx980), .A0 (q_4__14), .A1 (q_3__14), .S0 (nx1307)) ;
    dff gen_regs_3_regi_reg_q_14 (.Q (q_3__14), .QB (\$dummy [71]), .D (nx970), 
        .CLK (nx1333)) ;
    mux21_ni ix971 (.Y (nx970), .A0 (q_3__14), .A1 (q_2__14), .S0 (nx1307)) ;
    dff gen_regs_2_regi_reg_q_14 (.Q (q_2__14), .QB (\$dummy [72]), .D (nx960), 
        .CLK (nx1333)) ;
    mux21_ni ix961 (.Y (nx960), .A0 (q_2__14), .A1 (q_1__14), .S0 (nx1307)) ;
    dff gen_regs_1_regi_reg_q_14 (.Q (q_1__14), .QB (\$dummy [73]), .D (nx950), 
        .CLK (nx1333)) ;
    mux21_ni ix951 (.Y (nx950), .A0 (q_1__14), .A1 (q_0__14), .S0 (nx1307)) ;
    dff reg0_reg_q_14 (.Q (q_0__14), .QB (\$dummy [74]), .D (nx940), .CLK (
        nx1333)) ;
    mux21_ni ix941 (.Y (nx940), .A0 (q_0__14), .A1 (d[14]), .S0 (nx1307)) ;
    dff gen_regs_4_regi_reg_q_15 (.Q (q_4__15), .QB (\$dummy [75]), .D (nx1030)
        , .CLK (nx1335)) ;
    mux21_ni ix1031 (.Y (nx1030), .A0 (q_4__15), .A1 (q_3__15), .S0 (nx1309)) ;
    dff gen_regs_3_regi_reg_q_15 (.Q (q_3__15), .QB (\$dummy [76]), .D (nx1020)
        , .CLK (nx1335)) ;
    mux21_ni ix1021 (.Y (nx1020), .A0 (q_3__15), .A1 (q_2__15), .S0 (nx1309)) ;
    dff gen_regs_2_regi_reg_q_15 (.Q (q_2__15), .QB (\$dummy [77]), .D (nx1010)
        , .CLK (nx1335)) ;
    mux21_ni ix1011 (.Y (nx1010), .A0 (q_2__15), .A1 (q_1__15), .S0 (nx1309)) ;
    dff gen_regs_1_regi_reg_q_15 (.Q (q_1__15), .QB (\$dummy [78]), .D (nx1000)
        , .CLK (nx1333)) ;
    mux21_ni ix1001 (.Y (nx1000), .A0 (q_1__15), .A1 (q_0__15), .S0 (nx1307)) ;
    dff reg0_reg_q_15 (.Q (q_0__15), .QB (\$dummy [79]), .D (nx990), .CLK (
        nx1333)) ;
    mux21_ni ix991 (.Y (nx990), .A0 (q_0__15), .A1 (d[15]), .S0 (nx1307)) ;
    inv02 ix1286 (.Y (nx1287), .A (nx1337)) ;
    inv02 ix1288 (.Y (nx1289), .A (nx1337)) ;
    inv02 ix1290 (.Y (nx1291), .A (nx1337)) ;
    inv02 ix1292 (.Y (nx1293), .A (nx1337)) ;
    inv02 ix1294 (.Y (nx1295), .A (nx1337)) ;
    inv02 ix1296 (.Y (nx1297), .A (nx1337)) ;
    inv02 ix1298 (.Y (nx1299), .A (nx1337)) ;
    inv02 ix1300 (.Y (nx1301), .A (nx1339)) ;
    inv02 ix1302 (.Y (nx1303), .A (nx1339)) ;
    inv02 ix1304 (.Y (nx1305), .A (nx1339)) ;
    inv02 ix1306 (.Y (nx1307), .A (nx1339)) ;
    inv02 ix1308 (.Y (nx1309), .A (nx1339)) ;
    inv02 ix1312 (.Y (nx1313), .A (nx1341)) ;
    inv02 ix1314 (.Y (nx1315), .A (nx1341)) ;
    inv02 ix1316 (.Y (nx1317), .A (nx1341)) ;
    inv02 ix1318 (.Y (nx1319), .A (nx1341)) ;
    inv02 ix1320 (.Y (nx1321), .A (nx1341)) ;
    inv02 ix1322 (.Y (nx1323), .A (nx1341)) ;
    inv02 ix1324 (.Y (nx1325), .A (nx1341)) ;
    inv02 ix1326 (.Y (nx1327), .A (nx1343)) ;
    inv02 ix1328 (.Y (nx1329), .A (nx1343)) ;
    inv02 ix1330 (.Y (nx1331), .A (nx1343)) ;
    inv02 ix1332 (.Y (nx1333), .A (nx1343)) ;
    inv02 ix1334 (.Y (nx1335), .A (nx1343)) ;
    inv02 ix1336 (.Y (nx1337), .A (load)) ;
    inv02 ix1338 (.Y (nx1339), .A (load)) ;
    inv02 ix1340 (.Y (nx1341), .A (clk)) ;
    inv02 ix1342 (.Y (nx1343), .A (clk)) ;
endmodule


module ComputationPipeline ( img_data_0__15, img_data_0__14, img_data_0__13, 
                             img_data_0__12, img_data_0__11, img_data_0__10, 
                             img_data_0__9, img_data_0__8, img_data_0__7, 
                             img_data_0__6, img_data_0__5, img_data_0__4, 
                             img_data_0__3, img_data_0__2, img_data_0__1, 
                             img_data_0__0, img_data_1__15, img_data_1__14, 
                             img_data_1__13, img_data_1__12, img_data_1__11, 
                             img_data_1__10, img_data_1__9, img_data_1__8, 
                             img_data_1__7, img_data_1__6, img_data_1__5, 
                             img_data_1__4, img_data_1__3, img_data_1__2, 
                             img_data_1__1, img_data_1__0, img_data_2__15, 
                             img_data_2__14, img_data_2__13, img_data_2__12, 
                             img_data_2__11, img_data_2__10, img_data_2__9, 
                             img_data_2__8, img_data_2__7, img_data_2__6, 
                             img_data_2__5, img_data_2__4, img_data_2__3, 
                             img_data_2__2, img_data_2__1, img_data_2__0, 
                             img_data_3__15, img_data_3__14, img_data_3__13, 
                             img_data_3__12, img_data_3__11, img_data_3__10, 
                             img_data_3__9, img_data_3__8, img_data_3__7, 
                             img_data_3__6, img_data_3__5, img_data_3__4, 
                             img_data_3__3, img_data_3__2, img_data_3__1, 
                             img_data_3__0, img_data_4__15, img_data_4__14, 
                             img_data_4__13, img_data_4__12, img_data_4__11, 
                             img_data_4__10, img_data_4__9, img_data_4__8, 
                             img_data_4__7, img_data_4__6, img_data_4__5, 
                             img_data_4__4, img_data_4__3, img_data_4__2, 
                             img_data_4__1, img_data_4__0, img_data_5__15, 
                             img_data_5__14, img_data_5__13, img_data_5__12, 
                             img_data_5__11, img_data_5__10, img_data_5__9, 
                             img_data_5__8, img_data_5__7, img_data_5__6, 
                             img_data_5__5, img_data_5__4, img_data_5__3, 
                             img_data_5__2, img_data_5__1, img_data_5__0, 
                             img_data_6__15, img_data_6__14, img_data_6__13, 
                             img_data_6__12, img_data_6__11, img_data_6__10, 
                             img_data_6__9, img_data_6__8, img_data_6__7, 
                             img_data_6__6, img_data_6__5, img_data_6__4, 
                             img_data_6__3, img_data_6__2, img_data_6__1, 
                             img_data_6__0, img_data_7__15, img_data_7__14, 
                             img_data_7__13, img_data_7__12, img_data_7__11, 
                             img_data_7__10, img_data_7__9, img_data_7__8, 
                             img_data_7__7, img_data_7__6, img_data_7__5, 
                             img_data_7__4, img_data_7__3, img_data_7__2, 
                             img_data_7__1, img_data_7__0, img_data_8__15, 
                             img_data_8__14, img_data_8__13, img_data_8__12, 
                             img_data_8__11, img_data_8__10, img_data_8__9, 
                             img_data_8__8, img_data_8__7, img_data_8__6, 
                             img_data_8__5, img_data_8__4, img_data_8__3, 
                             img_data_8__2, img_data_8__1, img_data_8__0, 
                             img_data_9__15, img_data_9__14, img_data_9__13, 
                             img_data_9__12, img_data_9__11, img_data_9__10, 
                             img_data_9__9, img_data_9__8, img_data_9__7, 
                             img_data_9__6, img_data_9__5, img_data_9__4, 
                             img_data_9__3, img_data_9__2, img_data_9__1, 
                             img_data_9__0, img_data_10__15, img_data_10__14, 
                             img_data_10__13, img_data_10__12, img_data_10__11, 
                             img_data_10__10, img_data_10__9, img_data_10__8, 
                             img_data_10__7, img_data_10__6, img_data_10__5, 
                             img_data_10__4, img_data_10__3, img_data_10__2, 
                             img_data_10__1, img_data_10__0, img_data_11__15, 
                             img_data_11__14, img_data_11__13, img_data_11__12, 
                             img_data_11__11, img_data_11__10, img_data_11__9, 
                             img_data_11__8, img_data_11__7, img_data_11__6, 
                             img_data_11__5, img_data_11__4, img_data_11__3, 
                             img_data_11__2, img_data_11__1, img_data_11__0, 
                             img_data_12__15, img_data_12__14, img_data_12__13, 
                             img_data_12__12, img_data_12__11, img_data_12__10, 
                             img_data_12__9, img_data_12__8, img_data_12__7, 
                             img_data_12__6, img_data_12__5, img_data_12__4, 
                             img_data_12__3, img_data_12__2, img_data_12__1, 
                             img_data_12__0, img_data_13__15, img_data_13__14, 
                             img_data_13__13, img_data_13__12, img_data_13__11, 
                             img_data_13__10, img_data_13__9, img_data_13__8, 
                             img_data_13__7, img_data_13__6, img_data_13__5, 
                             img_data_13__4, img_data_13__3, img_data_13__2, 
                             img_data_13__1, img_data_13__0, img_data_14__15, 
                             img_data_14__14, img_data_14__13, img_data_14__12, 
                             img_data_14__11, img_data_14__10, img_data_14__9, 
                             img_data_14__8, img_data_14__7, img_data_14__6, 
                             img_data_14__5, img_data_14__4, img_data_14__3, 
                             img_data_14__2, img_data_14__1, img_data_14__0, 
                             img_data_15__15, img_data_15__14, img_data_15__13, 
                             img_data_15__12, img_data_15__11, img_data_15__10, 
                             img_data_15__9, img_data_15__8, img_data_15__7, 
                             img_data_15__6, img_data_15__5, img_data_15__4, 
                             img_data_15__3, img_data_15__2, img_data_15__1, 
                             img_data_15__0, img_data_16__15, img_data_16__14, 
                             img_data_16__13, img_data_16__12, img_data_16__11, 
                             img_data_16__10, img_data_16__9, img_data_16__8, 
                             img_data_16__7, img_data_16__6, img_data_16__5, 
                             img_data_16__4, img_data_16__3, img_data_16__2, 
                             img_data_16__1, img_data_16__0, img_data_17__15, 
                             img_data_17__14, img_data_17__13, img_data_17__12, 
                             img_data_17__11, img_data_17__10, img_data_17__9, 
                             img_data_17__8, img_data_17__7, img_data_17__6, 
                             img_data_17__5, img_data_17__4, img_data_17__3, 
                             img_data_17__2, img_data_17__1, img_data_17__0, 
                             img_data_18__15, img_data_18__14, img_data_18__13, 
                             img_data_18__12, img_data_18__11, img_data_18__10, 
                             img_data_18__9, img_data_18__8, img_data_18__7, 
                             img_data_18__6, img_data_18__5, img_data_18__4, 
                             img_data_18__3, img_data_18__2, img_data_18__1, 
                             img_data_18__0, img_data_19__15, img_data_19__14, 
                             img_data_19__13, img_data_19__12, img_data_19__11, 
                             img_data_19__10, img_data_19__9, img_data_19__8, 
                             img_data_19__7, img_data_19__6, img_data_19__5, 
                             img_data_19__4, img_data_19__3, img_data_19__2, 
                             img_data_19__1, img_data_19__0, img_data_20__15, 
                             img_data_20__14, img_data_20__13, img_data_20__12, 
                             img_data_20__11, img_data_20__10, img_data_20__9, 
                             img_data_20__8, img_data_20__7, img_data_20__6, 
                             img_data_20__5, img_data_20__4, img_data_20__3, 
                             img_data_20__2, img_data_20__1, img_data_20__0, 
                             img_data_21__15, img_data_21__14, img_data_21__13, 
                             img_data_21__12, img_data_21__11, img_data_21__10, 
                             img_data_21__9, img_data_21__8, img_data_21__7, 
                             img_data_21__6, img_data_21__5, img_data_21__4, 
                             img_data_21__3, img_data_21__2, img_data_21__1, 
                             img_data_21__0, img_data_22__15, img_data_22__14, 
                             img_data_22__13, img_data_22__12, img_data_22__11, 
                             img_data_22__10, img_data_22__9, img_data_22__8, 
                             img_data_22__7, img_data_22__6, img_data_22__5, 
                             img_data_22__4, img_data_22__3, img_data_22__2, 
                             img_data_22__1, img_data_22__0, img_data_23__15, 
                             img_data_23__14, img_data_23__13, img_data_23__12, 
                             img_data_23__11, img_data_23__10, img_data_23__9, 
                             img_data_23__8, img_data_23__7, img_data_23__6, 
                             img_data_23__5, img_data_23__4, img_data_23__3, 
                             img_data_23__2, img_data_23__1, img_data_23__0, 
                             img_data_24__15, img_data_24__14, img_data_24__13, 
                             img_data_24__12, img_data_24__11, img_data_24__10, 
                             img_data_24__9, img_data_24__8, img_data_24__7, 
                             img_data_24__6, img_data_24__5, img_data_24__4, 
                             img_data_24__3, img_data_24__2, img_data_24__1, 
                             img_data_24__0, filter_data_0__15, 
                             filter_data_0__14, filter_data_0__13, 
                             filter_data_0__12, filter_data_0__11, 
                             filter_data_0__10, filter_data_0__9, 
                             filter_data_0__8, filter_data_0__7, 
                             filter_data_0__6, filter_data_0__5, 
                             filter_data_0__4, filter_data_0__3, 
                             filter_data_0__2, filter_data_0__1, 
                             filter_data_0__0, filter_data_1__15, 
                             filter_data_1__14, filter_data_1__13, 
                             filter_data_1__12, filter_data_1__11, 
                             filter_data_1__10, filter_data_1__9, 
                             filter_data_1__8, filter_data_1__7, 
                             filter_data_1__6, filter_data_1__5, 
                             filter_data_1__4, filter_data_1__3, 
                             filter_data_1__2, filter_data_1__1, 
                             filter_data_1__0, filter_data_2__15, 
                             filter_data_2__14, filter_data_2__13, 
                             filter_data_2__12, filter_data_2__11, 
                             filter_data_2__10, filter_data_2__9, 
                             filter_data_2__8, filter_data_2__7, 
                             filter_data_2__6, filter_data_2__5, 
                             filter_data_2__4, filter_data_2__3, 
                             filter_data_2__2, filter_data_2__1, 
                             filter_data_2__0, filter_data_3__15, 
                             filter_data_3__14, filter_data_3__13, 
                             filter_data_3__12, filter_data_3__11, 
                             filter_data_3__10, filter_data_3__9, 
                             filter_data_3__8, filter_data_3__7, 
                             filter_data_3__6, filter_data_3__5, 
                             filter_data_3__4, filter_data_3__3, 
                             filter_data_3__2, filter_data_3__1, 
                             filter_data_3__0, filter_data_4__15, 
                             filter_data_4__14, filter_data_4__13, 
                             filter_data_4__12, filter_data_4__11, 
                             filter_data_4__10, filter_data_4__9, 
                             filter_data_4__8, filter_data_4__7, 
                             filter_data_4__6, filter_data_4__5, 
                             filter_data_4__4, filter_data_4__3, 
                             filter_data_4__2, filter_data_4__1, 
                             filter_data_4__0, filter_data_5__15, 
                             filter_data_5__14, filter_data_5__13, 
                             filter_data_5__12, filter_data_5__11, 
                             filter_data_5__10, filter_data_5__9, 
                             filter_data_5__8, filter_data_5__7, 
                             filter_data_5__6, filter_data_5__5, 
                             filter_data_5__4, filter_data_5__3, 
                             filter_data_5__2, filter_data_5__1, 
                             filter_data_5__0, filter_data_6__15, 
                             filter_data_6__14, filter_data_6__13, 
                             filter_data_6__12, filter_data_6__11, 
                             filter_data_6__10, filter_data_6__9, 
                             filter_data_6__8, filter_data_6__7, 
                             filter_data_6__6, filter_data_6__5, 
                             filter_data_6__4, filter_data_6__3, 
                             filter_data_6__2, filter_data_6__1, 
                             filter_data_6__0, filter_data_7__15, 
                             filter_data_7__14, filter_data_7__13, 
                             filter_data_7__12, filter_data_7__11, 
                             filter_data_7__10, filter_data_7__9, 
                             filter_data_7__8, filter_data_7__7, 
                             filter_data_7__6, filter_data_7__5, 
                             filter_data_7__4, filter_data_7__3, 
                             filter_data_7__2, filter_data_7__1, 
                             filter_data_7__0, filter_data_8__15, 
                             filter_data_8__14, filter_data_8__13, 
                             filter_data_8__12, filter_data_8__11, 
                             filter_data_8__10, filter_data_8__9, 
                             filter_data_8__8, filter_data_8__7, 
                             filter_data_8__6, filter_data_8__5, 
                             filter_data_8__4, filter_data_8__3, 
                             filter_data_8__2, filter_data_8__1, 
                             filter_data_8__0, filter_data_9__15, 
                             filter_data_9__14, filter_data_9__13, 
                             filter_data_9__12, filter_data_9__11, 
                             filter_data_9__10, filter_data_9__9, 
                             filter_data_9__8, filter_data_9__7, 
                             filter_data_9__6, filter_data_9__5, 
                             filter_data_9__4, filter_data_9__3, 
                             filter_data_9__2, filter_data_9__1, 
                             filter_data_9__0, filter_data_10__15, 
                             filter_data_10__14, filter_data_10__13, 
                             filter_data_10__12, filter_data_10__11, 
                             filter_data_10__10, filter_data_10__9, 
                             filter_data_10__8, filter_data_10__7, 
                             filter_data_10__6, filter_data_10__5, 
                             filter_data_10__4, filter_data_10__3, 
                             filter_data_10__2, filter_data_10__1, 
                             filter_data_10__0, filter_data_11__15, 
                             filter_data_11__14, filter_data_11__13, 
                             filter_data_11__12, filter_data_11__11, 
                             filter_data_11__10, filter_data_11__9, 
                             filter_data_11__8, filter_data_11__7, 
                             filter_data_11__6, filter_data_11__5, 
                             filter_data_11__4, filter_data_11__3, 
                             filter_data_11__2, filter_data_11__1, 
                             filter_data_11__0, filter_data_12__15, 
                             filter_data_12__14, filter_data_12__13, 
                             filter_data_12__12, filter_data_12__11, 
                             filter_data_12__10, filter_data_12__9, 
                             filter_data_12__8, filter_data_12__7, 
                             filter_data_12__6, filter_data_12__5, 
                             filter_data_12__4, filter_data_12__3, 
                             filter_data_12__2, filter_data_12__1, 
                             filter_data_12__0, filter_data_13__15, 
                             filter_data_13__14, filter_data_13__13, 
                             filter_data_13__12, filter_data_13__11, 
                             filter_data_13__10, filter_data_13__9, 
                             filter_data_13__8, filter_data_13__7, 
                             filter_data_13__6, filter_data_13__5, 
                             filter_data_13__4, filter_data_13__3, 
                             filter_data_13__2, filter_data_13__1, 
                             filter_data_13__0, filter_data_14__15, 
                             filter_data_14__14, filter_data_14__13, 
                             filter_data_14__12, filter_data_14__11, 
                             filter_data_14__10, filter_data_14__9, 
                             filter_data_14__8, filter_data_14__7, 
                             filter_data_14__6, filter_data_14__5, 
                             filter_data_14__4, filter_data_14__3, 
                             filter_data_14__2, filter_data_14__1, 
                             filter_data_14__0, filter_data_15__15, 
                             filter_data_15__14, filter_data_15__13, 
                             filter_data_15__12, filter_data_15__11, 
                             filter_data_15__10, filter_data_15__9, 
                             filter_data_15__8, filter_data_15__7, 
                             filter_data_15__6, filter_data_15__5, 
                             filter_data_15__4, filter_data_15__3, 
                             filter_data_15__2, filter_data_15__1, 
                             filter_data_15__0, filter_data_16__15, 
                             filter_data_16__14, filter_data_16__13, 
                             filter_data_16__12, filter_data_16__11, 
                             filter_data_16__10, filter_data_16__9, 
                             filter_data_16__8, filter_data_16__7, 
                             filter_data_16__6, filter_data_16__5, 
                             filter_data_16__4, filter_data_16__3, 
                             filter_data_16__2, filter_data_16__1, 
                             filter_data_16__0, filter_data_17__15, 
                             filter_data_17__14, filter_data_17__13, 
                             filter_data_17__12, filter_data_17__11, 
                             filter_data_17__10, filter_data_17__9, 
                             filter_data_17__8, filter_data_17__7, 
                             filter_data_17__6, filter_data_17__5, 
                             filter_data_17__4, filter_data_17__3, 
                             filter_data_17__2, filter_data_17__1, 
                             filter_data_17__0, filter_data_18__15, 
                             filter_data_18__14, filter_data_18__13, 
                             filter_data_18__12, filter_data_18__11, 
                             filter_data_18__10, filter_data_18__9, 
                             filter_data_18__8, filter_data_18__7, 
                             filter_data_18__6, filter_data_18__5, 
                             filter_data_18__4, filter_data_18__3, 
                             filter_data_18__2, filter_data_18__1, 
                             filter_data_18__0, filter_data_19__15, 
                             filter_data_19__14, filter_data_19__13, 
                             filter_data_19__12, filter_data_19__11, 
                             filter_data_19__10, filter_data_19__9, 
                             filter_data_19__8, filter_data_19__7, 
                             filter_data_19__6, filter_data_19__5, 
                             filter_data_19__4, filter_data_19__3, 
                             filter_data_19__2, filter_data_19__1, 
                             filter_data_19__0, filter_data_20__15, 
                             filter_data_20__14, filter_data_20__13, 
                             filter_data_20__12, filter_data_20__11, 
                             filter_data_20__10, filter_data_20__9, 
                             filter_data_20__8, filter_data_20__7, 
                             filter_data_20__6, filter_data_20__5, 
                             filter_data_20__4, filter_data_20__3, 
                             filter_data_20__2, filter_data_20__1, 
                             filter_data_20__0, filter_data_21__15, 
                             filter_data_21__14, filter_data_21__13, 
                             filter_data_21__12, filter_data_21__11, 
                             filter_data_21__10, filter_data_21__9, 
                             filter_data_21__8, filter_data_21__7, 
                             filter_data_21__6, filter_data_21__5, 
                             filter_data_21__4, filter_data_21__3, 
                             filter_data_21__2, filter_data_21__1, 
                             filter_data_21__0, filter_data_22__15, 
                             filter_data_22__14, filter_data_22__13, 
                             filter_data_22__12, filter_data_22__11, 
                             filter_data_22__10, filter_data_22__9, 
                             filter_data_22__8, filter_data_22__7, 
                             filter_data_22__6, filter_data_22__5, 
                             filter_data_22__4, filter_data_22__3, 
                             filter_data_22__2, filter_data_22__1, 
                             filter_data_22__0, filter_data_23__15, 
                             filter_data_23__14, filter_data_23__13, 
                             filter_data_23__12, filter_data_23__11, 
                             filter_data_23__10, filter_data_23__9, 
                             filter_data_23__8, filter_data_23__7, 
                             filter_data_23__6, filter_data_23__5, 
                             filter_data_23__4, filter_data_23__3, 
                             filter_data_23__2, filter_data_23__1, 
                             filter_data_23__0, filter_data_24__15, 
                             filter_data_24__14, filter_data_24__13, 
                             filter_data_24__12, filter_data_24__11, 
                             filter_data_24__10, filter_data_24__9, 
                             filter_data_24__8, filter_data_24__7, 
                             filter_data_24__6, filter_data_24__5, 
                             filter_data_24__4, filter_data_24__3, 
                             filter_data_24__2, filter_data_24__1, 
                             filter_data_24__0, d_arr_0__31, d_arr_0__30, 
                             d_arr_0__29, d_arr_0__28, d_arr_0__27, d_arr_0__26, 
                             d_arr_0__25, d_arr_0__24, d_arr_0__23, d_arr_0__22, 
                             d_arr_0__21, d_arr_0__20, d_arr_0__19, d_arr_0__18, 
                             d_arr_0__17, d_arr_0__16, d_arr_0__15, d_arr_0__14, 
                             d_arr_0__13, d_arr_0__12, d_arr_0__11, d_arr_0__10, 
                             d_arr_0__9, d_arr_0__8, d_arr_0__7, d_arr_0__6, 
                             d_arr_0__5, d_arr_0__4, d_arr_0__3, d_arr_0__2, 
                             d_arr_0__1, d_arr_0__0, d_arr_1__31, d_arr_1__30, 
                             d_arr_1__29, d_arr_1__28, d_arr_1__27, d_arr_1__26, 
                             d_arr_1__25, d_arr_1__24, d_arr_1__23, d_arr_1__22, 
                             d_arr_1__21, d_arr_1__20, d_arr_1__19, d_arr_1__18, 
                             d_arr_1__17, d_arr_1__16, d_arr_1__15, d_arr_1__14, 
                             d_arr_1__13, d_arr_1__12, d_arr_1__11, d_arr_1__10, 
                             d_arr_1__9, d_arr_1__8, d_arr_1__7, d_arr_1__6, 
                             d_arr_1__5, d_arr_1__4, d_arr_1__3, d_arr_1__2, 
                             d_arr_1__1, d_arr_1__0, d_arr_2__31, d_arr_2__30, 
                             d_arr_2__29, d_arr_2__28, d_arr_2__27, d_arr_2__26, 
                             d_arr_2__25, d_arr_2__24, d_arr_2__23, d_arr_2__22, 
                             d_arr_2__21, d_arr_2__20, d_arr_2__19, d_arr_2__18, 
                             d_arr_2__17, d_arr_2__16, d_arr_2__15, d_arr_2__14, 
                             d_arr_2__13, d_arr_2__12, d_arr_2__11, d_arr_2__10, 
                             d_arr_2__9, d_arr_2__8, d_arr_2__7, d_arr_2__6, 
                             d_arr_2__5, d_arr_2__4, d_arr_2__3, d_arr_2__2, 
                             d_arr_2__1, d_arr_2__0, d_arr_3__31, d_arr_3__30, 
                             d_arr_3__29, d_arr_3__28, d_arr_3__27, d_arr_3__26, 
                             d_arr_3__25, d_arr_3__24, d_arr_3__23, d_arr_3__22, 
                             d_arr_3__21, d_arr_3__20, d_arr_3__19, d_arr_3__18, 
                             d_arr_3__17, d_arr_3__16, d_arr_3__15, d_arr_3__14, 
                             d_arr_3__13, d_arr_3__12, d_arr_3__11, d_arr_3__10, 
                             d_arr_3__9, d_arr_3__8, d_arr_3__7, d_arr_3__6, 
                             d_arr_3__5, d_arr_3__4, d_arr_3__3, d_arr_3__2, 
                             d_arr_3__1, d_arr_3__0, d_arr_4__31, d_arr_4__30, 
                             d_arr_4__29, d_arr_4__28, d_arr_4__27, d_arr_4__26, 
                             d_arr_4__25, d_arr_4__24, d_arr_4__23, d_arr_4__22, 
                             d_arr_4__21, d_arr_4__20, d_arr_4__19, d_arr_4__18, 
                             d_arr_4__17, d_arr_4__16, d_arr_4__15, d_arr_4__14, 
                             d_arr_4__13, d_arr_4__12, d_arr_4__11, d_arr_4__10, 
                             d_arr_4__9, d_arr_4__8, d_arr_4__7, d_arr_4__6, 
                             d_arr_4__5, d_arr_4__4, d_arr_4__3, d_arr_4__2, 
                             d_arr_4__1, d_arr_4__0, d_arr_5__31, d_arr_5__30, 
                             d_arr_5__29, d_arr_5__28, d_arr_5__27, d_arr_5__26, 
                             d_arr_5__25, d_arr_5__24, d_arr_5__23, d_arr_5__22, 
                             d_arr_5__21, d_arr_5__20, d_arr_5__19, d_arr_5__18, 
                             d_arr_5__17, d_arr_5__16, d_arr_5__15, d_arr_5__14, 
                             d_arr_5__13, d_arr_5__12, d_arr_5__11, d_arr_5__10, 
                             d_arr_5__9, d_arr_5__8, d_arr_5__7, d_arr_5__6, 
                             d_arr_5__5, d_arr_5__4, d_arr_5__3, d_arr_5__2, 
                             d_arr_5__1, d_arr_5__0, d_arr_6__31, d_arr_6__30, 
                             d_arr_6__29, d_arr_6__28, d_arr_6__27, d_arr_6__26, 
                             d_arr_6__25, d_arr_6__24, d_arr_6__23, d_arr_6__22, 
                             d_arr_6__21, d_arr_6__20, d_arr_6__19, d_arr_6__18, 
                             d_arr_6__17, d_arr_6__16, d_arr_6__15, d_arr_6__14, 
                             d_arr_6__13, d_arr_6__12, d_arr_6__11, d_arr_6__10, 
                             d_arr_6__9, d_arr_6__8, d_arr_6__7, d_arr_6__6, 
                             d_arr_6__5, d_arr_6__4, d_arr_6__3, d_arr_6__2, 
                             d_arr_6__1, d_arr_6__0, d_arr_7__31, d_arr_7__30, 
                             d_arr_7__29, d_arr_7__28, d_arr_7__27, d_arr_7__26, 
                             d_arr_7__25, d_arr_7__24, d_arr_7__23, d_arr_7__22, 
                             d_arr_7__21, d_arr_7__20, d_arr_7__19, d_arr_7__18, 
                             d_arr_7__17, d_arr_7__16, d_arr_7__15, d_arr_7__14, 
                             d_arr_7__13, d_arr_7__12, d_arr_7__11, d_arr_7__10, 
                             d_arr_7__9, d_arr_7__8, d_arr_7__7, d_arr_7__6, 
                             d_arr_7__5, d_arr_7__4, d_arr_7__3, d_arr_7__2, 
                             d_arr_7__1, d_arr_7__0, d_arr_8__31, d_arr_8__30, 
                             d_arr_8__29, d_arr_8__28, d_arr_8__27, d_arr_8__26, 
                             d_arr_8__25, d_arr_8__24, d_arr_8__23, d_arr_8__22, 
                             d_arr_8__21, d_arr_8__20, d_arr_8__19, d_arr_8__18, 
                             d_arr_8__17, d_arr_8__16, d_arr_8__15, d_arr_8__14, 
                             d_arr_8__13, d_arr_8__12, d_arr_8__11, d_arr_8__10, 
                             d_arr_8__9, d_arr_8__8, d_arr_8__7, d_arr_8__6, 
                             d_arr_8__5, d_arr_8__4, d_arr_8__3, d_arr_8__2, 
                             d_arr_8__1, d_arr_8__0, d_arr_9__31, d_arr_9__30, 
                             d_arr_9__29, d_arr_9__28, d_arr_9__27, d_arr_9__26, 
                             d_arr_9__25, d_arr_9__24, d_arr_9__23, d_arr_9__22, 
                             d_arr_9__21, d_arr_9__20, d_arr_9__19, d_arr_9__18, 
                             d_arr_9__17, d_arr_9__16, d_arr_9__15, d_arr_9__14, 
                             d_arr_9__13, d_arr_9__12, d_arr_9__11, d_arr_9__10, 
                             d_arr_9__9, d_arr_9__8, d_arr_9__7, d_arr_9__6, 
                             d_arr_9__5, d_arr_9__4, d_arr_9__3, d_arr_9__2, 
                             d_arr_9__1, d_arr_9__0, d_arr_10__31, d_arr_10__30, 
                             d_arr_10__29, d_arr_10__28, d_arr_10__27, 
                             d_arr_10__26, d_arr_10__25, d_arr_10__24, 
                             d_arr_10__23, d_arr_10__22, d_arr_10__21, 
                             d_arr_10__20, d_arr_10__19, d_arr_10__18, 
                             d_arr_10__17, d_arr_10__16, d_arr_10__15, 
                             d_arr_10__14, d_arr_10__13, d_arr_10__12, 
                             d_arr_10__11, d_arr_10__10, d_arr_10__9, 
                             d_arr_10__8, d_arr_10__7, d_arr_10__6, d_arr_10__5, 
                             d_arr_10__4, d_arr_10__3, d_arr_10__2, d_arr_10__1, 
                             d_arr_10__0, d_arr_11__31, d_arr_11__30, 
                             d_arr_11__29, d_arr_11__28, d_arr_11__27, 
                             d_arr_11__26, d_arr_11__25, d_arr_11__24, 
                             d_arr_11__23, d_arr_11__22, d_arr_11__21, 
                             d_arr_11__20, d_arr_11__19, d_arr_11__18, 
                             d_arr_11__17, d_arr_11__16, d_arr_11__15, 
                             d_arr_11__14, d_arr_11__13, d_arr_11__12, 
                             d_arr_11__11, d_arr_11__10, d_arr_11__9, 
                             d_arr_11__8, d_arr_11__7, d_arr_11__6, d_arr_11__5, 
                             d_arr_11__4, d_arr_11__3, d_arr_11__2, d_arr_11__1, 
                             d_arr_11__0, d_arr_12__31, d_arr_12__30, 
                             d_arr_12__29, d_arr_12__28, d_arr_12__27, 
                             d_arr_12__26, d_arr_12__25, d_arr_12__24, 
                             d_arr_12__23, d_arr_12__22, d_arr_12__21, 
                             d_arr_12__20, d_arr_12__19, d_arr_12__18, 
                             d_arr_12__17, d_arr_12__16, d_arr_12__15, 
                             d_arr_12__14, d_arr_12__13, d_arr_12__12, 
                             d_arr_12__11, d_arr_12__10, d_arr_12__9, 
                             d_arr_12__8, d_arr_12__7, d_arr_12__6, d_arr_12__5, 
                             d_arr_12__4, d_arr_12__3, d_arr_12__2, d_arr_12__1, 
                             d_arr_12__0, d_arr_13__31, d_arr_13__30, 
                             d_arr_13__29, d_arr_13__28, d_arr_13__27, 
                             d_arr_13__26, d_arr_13__25, d_arr_13__24, 
                             d_arr_13__23, d_arr_13__22, d_arr_13__21, 
                             d_arr_13__20, d_arr_13__19, d_arr_13__18, 
                             d_arr_13__17, d_arr_13__16, d_arr_13__15, 
                             d_arr_13__14, d_arr_13__13, d_arr_13__12, 
                             d_arr_13__11, d_arr_13__10, d_arr_13__9, 
                             d_arr_13__8, d_arr_13__7, d_arr_13__6, d_arr_13__5, 
                             d_arr_13__4, d_arr_13__3, d_arr_13__2, d_arr_13__1, 
                             d_arr_13__0, d_arr_14__31, d_arr_14__30, 
                             d_arr_14__29, d_arr_14__28, d_arr_14__27, 
                             d_arr_14__26, d_arr_14__25, d_arr_14__24, 
                             d_arr_14__23, d_arr_14__22, d_arr_14__21, 
                             d_arr_14__20, d_arr_14__19, d_arr_14__18, 
                             d_arr_14__17, d_arr_14__16, d_arr_14__15, 
                             d_arr_14__14, d_arr_14__13, d_arr_14__12, 
                             d_arr_14__11, d_arr_14__10, d_arr_14__9, 
                             d_arr_14__8, d_arr_14__7, d_arr_14__6, d_arr_14__5, 
                             d_arr_14__4, d_arr_14__3, d_arr_14__2, d_arr_14__1, 
                             d_arr_14__0, d_arr_15__31, d_arr_15__30, 
                             d_arr_15__29, d_arr_15__28, d_arr_15__27, 
                             d_arr_15__26, d_arr_15__25, d_arr_15__24, 
                             d_arr_15__23, d_arr_15__22, d_arr_15__21, 
                             d_arr_15__20, d_arr_15__19, d_arr_15__18, 
                             d_arr_15__17, d_arr_15__16, d_arr_15__15, 
                             d_arr_15__14, d_arr_15__13, d_arr_15__12, 
                             d_arr_15__11, d_arr_15__10, d_arr_15__9, 
                             d_arr_15__8, d_arr_15__7, d_arr_15__6, d_arr_15__5, 
                             d_arr_15__4, d_arr_15__3, d_arr_15__2, d_arr_15__1, 
                             d_arr_15__0, d_arr_16__31, d_arr_16__30, 
                             d_arr_16__29, d_arr_16__28, d_arr_16__27, 
                             d_arr_16__26, d_arr_16__25, d_arr_16__24, 
                             d_arr_16__23, d_arr_16__22, d_arr_16__21, 
                             d_arr_16__20, d_arr_16__19, d_arr_16__18, 
                             d_arr_16__17, d_arr_16__16, d_arr_16__15, 
                             d_arr_16__14, d_arr_16__13, d_arr_16__12, 
                             d_arr_16__11, d_arr_16__10, d_arr_16__9, 
                             d_arr_16__8, d_arr_16__7, d_arr_16__6, d_arr_16__5, 
                             d_arr_16__4, d_arr_16__3, d_arr_16__2, d_arr_16__1, 
                             d_arr_16__0, d_arr_17__31, d_arr_17__30, 
                             d_arr_17__29, d_arr_17__28, d_arr_17__27, 
                             d_arr_17__26, d_arr_17__25, d_arr_17__24, 
                             d_arr_17__23, d_arr_17__22, d_arr_17__21, 
                             d_arr_17__20, d_arr_17__19, d_arr_17__18, 
                             d_arr_17__17, d_arr_17__16, d_arr_17__15, 
                             d_arr_17__14, d_arr_17__13, d_arr_17__12, 
                             d_arr_17__11, d_arr_17__10, d_arr_17__9, 
                             d_arr_17__8, d_arr_17__7, d_arr_17__6, d_arr_17__5, 
                             d_arr_17__4, d_arr_17__3, d_arr_17__2, d_arr_17__1, 
                             d_arr_17__0, d_arr_18__31, d_arr_18__30, 
                             d_arr_18__29, d_arr_18__28, d_arr_18__27, 
                             d_arr_18__26, d_arr_18__25, d_arr_18__24, 
                             d_arr_18__23, d_arr_18__22, d_arr_18__21, 
                             d_arr_18__20, d_arr_18__19, d_arr_18__18, 
                             d_arr_18__17, d_arr_18__16, d_arr_18__15, 
                             d_arr_18__14, d_arr_18__13, d_arr_18__12, 
                             d_arr_18__11, d_arr_18__10, d_arr_18__9, 
                             d_arr_18__8, d_arr_18__7, d_arr_18__6, d_arr_18__5, 
                             d_arr_18__4, d_arr_18__3, d_arr_18__2, d_arr_18__1, 
                             d_arr_18__0, d_arr_19__31, d_arr_19__30, 
                             d_arr_19__29, d_arr_19__28, d_arr_19__27, 
                             d_arr_19__26, d_arr_19__25, d_arr_19__24, 
                             d_arr_19__23, d_arr_19__22, d_arr_19__21, 
                             d_arr_19__20, d_arr_19__19, d_arr_19__18, 
                             d_arr_19__17, d_arr_19__16, d_arr_19__15, 
                             d_arr_19__14, d_arr_19__13, d_arr_19__12, 
                             d_arr_19__11, d_arr_19__10, d_arr_19__9, 
                             d_arr_19__8, d_arr_19__7, d_arr_19__6, d_arr_19__5, 
                             d_arr_19__4, d_arr_19__3, d_arr_19__2, d_arr_19__1, 
                             d_arr_19__0, d_arr_20__31, d_arr_20__30, 
                             d_arr_20__29, d_arr_20__28, d_arr_20__27, 
                             d_arr_20__26, d_arr_20__25, d_arr_20__24, 
                             d_arr_20__23, d_arr_20__22, d_arr_20__21, 
                             d_arr_20__20, d_arr_20__19, d_arr_20__18, 
                             d_arr_20__17, d_arr_20__16, d_arr_20__15, 
                             d_arr_20__14, d_arr_20__13, d_arr_20__12, 
                             d_arr_20__11, d_arr_20__10, d_arr_20__9, 
                             d_arr_20__8, d_arr_20__7, d_arr_20__6, d_arr_20__5, 
                             d_arr_20__4, d_arr_20__3, d_arr_20__2, d_arr_20__1, 
                             d_arr_20__0, d_arr_21__31, d_arr_21__30, 
                             d_arr_21__29, d_arr_21__28, d_arr_21__27, 
                             d_arr_21__26, d_arr_21__25, d_arr_21__24, 
                             d_arr_21__23, d_arr_21__22, d_arr_21__21, 
                             d_arr_21__20, d_arr_21__19, d_arr_21__18, 
                             d_arr_21__17, d_arr_21__16, d_arr_21__15, 
                             d_arr_21__14, d_arr_21__13, d_arr_21__12, 
                             d_arr_21__11, d_arr_21__10, d_arr_21__9, 
                             d_arr_21__8, d_arr_21__7, d_arr_21__6, d_arr_21__5, 
                             d_arr_21__4, d_arr_21__3, d_arr_21__2, d_arr_21__1, 
                             d_arr_21__0, d_arr_22__31, d_arr_22__30, 
                             d_arr_22__29, d_arr_22__28, d_arr_22__27, 
                             d_arr_22__26, d_arr_22__25, d_arr_22__24, 
                             d_arr_22__23, d_arr_22__22, d_arr_22__21, 
                             d_arr_22__20, d_arr_22__19, d_arr_22__18, 
                             d_arr_22__17, d_arr_22__16, d_arr_22__15, 
                             d_arr_22__14, d_arr_22__13, d_arr_22__12, 
                             d_arr_22__11, d_arr_22__10, d_arr_22__9, 
                             d_arr_22__8, d_arr_22__7, d_arr_22__6, d_arr_22__5, 
                             d_arr_22__4, d_arr_22__3, d_arr_22__2, d_arr_22__1, 
                             d_arr_22__0, d_arr_23__31, d_arr_23__30, 
                             d_arr_23__29, d_arr_23__28, d_arr_23__27, 
                             d_arr_23__26, d_arr_23__25, d_arr_23__24, 
                             d_arr_23__23, d_arr_23__22, d_arr_23__21, 
                             d_arr_23__20, d_arr_23__19, d_arr_23__18, 
                             d_arr_23__17, d_arr_23__16, d_arr_23__15, 
                             d_arr_23__14, d_arr_23__13, d_arr_23__12, 
                             d_arr_23__11, d_arr_23__10, d_arr_23__9, 
                             d_arr_23__8, d_arr_23__7, d_arr_23__6, d_arr_23__5, 
                             d_arr_23__4, d_arr_23__3, d_arr_23__2, d_arr_23__1, 
                             d_arr_23__0, d_arr_24__31, d_arr_24__30, 
                             d_arr_24__29, d_arr_24__28, d_arr_24__27, 
                             d_arr_24__26, d_arr_24__25, d_arr_24__24, 
                             d_arr_24__23, d_arr_24__22, d_arr_24__21, 
                             d_arr_24__20, d_arr_24__19, d_arr_24__18, 
                             d_arr_24__17, d_arr_24__16, d_arr_24__15, 
                             d_arr_24__14, d_arr_24__13, d_arr_24__12, 
                             d_arr_24__11, d_arr_24__10, d_arr_24__9, 
                             d_arr_24__8, d_arr_24__7, d_arr_24__6, d_arr_24__5, 
                             d_arr_24__4, d_arr_24__3, d_arr_24__2, d_arr_24__1, 
                             d_arr_24__0, q_arr_0__31, q_arr_0__30, q_arr_0__29, 
                             q_arr_0__28, q_arr_0__27, q_arr_0__26, q_arr_0__25, 
                             q_arr_0__24, q_arr_0__23, q_arr_0__22, q_arr_0__21, 
                             q_arr_0__20, q_arr_0__19, q_arr_0__18, q_arr_0__17, 
                             q_arr_0__16, q_arr_0__15, q_arr_0__14, q_arr_0__13, 
                             q_arr_0__12, q_arr_0__11, q_arr_0__10, q_arr_0__9, 
                             q_arr_0__8, q_arr_0__7, q_arr_0__6, q_arr_0__5, 
                             q_arr_0__4, q_arr_0__3, q_arr_0__2, q_arr_0__1, 
                             q_arr_0__0, q_arr_1__31, q_arr_1__30, q_arr_1__29, 
                             q_arr_1__28, q_arr_1__27, q_arr_1__26, q_arr_1__25, 
                             q_arr_1__24, q_arr_1__23, q_arr_1__22, q_arr_1__21, 
                             q_arr_1__20, q_arr_1__19, q_arr_1__18, q_arr_1__17, 
                             q_arr_1__16, q_arr_1__15, q_arr_1__14, q_arr_1__13, 
                             q_arr_1__12, q_arr_1__11, q_arr_1__10, q_arr_1__9, 
                             q_arr_1__8, q_arr_1__7, q_arr_1__6, q_arr_1__5, 
                             q_arr_1__4, q_arr_1__3, q_arr_1__2, q_arr_1__1, 
                             q_arr_1__0, q_arr_2__31, q_arr_2__30, q_arr_2__29, 
                             q_arr_2__28, q_arr_2__27, q_arr_2__26, q_arr_2__25, 
                             q_arr_2__24, q_arr_2__23, q_arr_2__22, q_arr_2__21, 
                             q_arr_2__20, q_arr_2__19, q_arr_2__18, q_arr_2__17, 
                             q_arr_2__16, q_arr_2__15, q_arr_2__14, q_arr_2__13, 
                             q_arr_2__12, q_arr_2__11, q_arr_2__10, q_arr_2__9, 
                             q_arr_2__8, q_arr_2__7, q_arr_2__6, q_arr_2__5, 
                             q_arr_2__4, q_arr_2__3, q_arr_2__2, q_arr_2__1, 
                             q_arr_2__0, q_arr_3__31, q_arr_3__30, q_arr_3__29, 
                             q_arr_3__28, q_arr_3__27, q_arr_3__26, q_arr_3__25, 
                             q_arr_3__24, q_arr_3__23, q_arr_3__22, q_arr_3__21, 
                             q_arr_3__20, q_arr_3__19, q_arr_3__18, q_arr_3__17, 
                             q_arr_3__16, q_arr_3__15, q_arr_3__14, q_arr_3__13, 
                             q_arr_3__12, q_arr_3__11, q_arr_3__10, q_arr_3__9, 
                             q_arr_3__8, q_arr_3__7, q_arr_3__6, q_arr_3__5, 
                             q_arr_3__4, q_arr_3__3, q_arr_3__2, q_arr_3__1, 
                             q_arr_3__0, q_arr_4__31, q_arr_4__30, q_arr_4__29, 
                             q_arr_4__28, q_arr_4__27, q_arr_4__26, q_arr_4__25, 
                             q_arr_4__24, q_arr_4__23, q_arr_4__22, q_arr_4__21, 
                             q_arr_4__20, q_arr_4__19, q_arr_4__18, q_arr_4__17, 
                             q_arr_4__16, q_arr_4__15, q_arr_4__14, q_arr_4__13, 
                             q_arr_4__12, q_arr_4__11, q_arr_4__10, q_arr_4__9, 
                             q_arr_4__8, q_arr_4__7, q_arr_4__6, q_arr_4__5, 
                             q_arr_4__4, q_arr_4__3, q_arr_4__2, q_arr_4__1, 
                             q_arr_4__0, q_arr_5__31, q_arr_5__30, q_arr_5__29, 
                             q_arr_5__28, q_arr_5__27, q_arr_5__26, q_arr_5__25, 
                             q_arr_5__24, q_arr_5__23, q_arr_5__22, q_arr_5__21, 
                             q_arr_5__20, q_arr_5__19, q_arr_5__18, q_arr_5__17, 
                             q_arr_5__16, q_arr_5__15, q_arr_5__14, q_arr_5__13, 
                             q_arr_5__12, q_arr_5__11, q_arr_5__10, q_arr_5__9, 
                             q_arr_5__8, q_arr_5__7, q_arr_5__6, q_arr_5__5, 
                             q_arr_5__4, q_arr_5__3, q_arr_5__2, q_arr_5__1, 
                             q_arr_5__0, q_arr_6__31, q_arr_6__30, q_arr_6__29, 
                             q_arr_6__28, q_arr_6__27, q_arr_6__26, q_arr_6__25, 
                             q_arr_6__24, q_arr_6__23, q_arr_6__22, q_arr_6__21, 
                             q_arr_6__20, q_arr_6__19, q_arr_6__18, q_arr_6__17, 
                             q_arr_6__16, q_arr_6__15, q_arr_6__14, q_arr_6__13, 
                             q_arr_6__12, q_arr_6__11, q_arr_6__10, q_arr_6__9, 
                             q_arr_6__8, q_arr_6__7, q_arr_6__6, q_arr_6__5, 
                             q_arr_6__4, q_arr_6__3, q_arr_6__2, q_arr_6__1, 
                             q_arr_6__0, q_arr_7__31, q_arr_7__30, q_arr_7__29, 
                             q_arr_7__28, q_arr_7__27, q_arr_7__26, q_arr_7__25, 
                             q_arr_7__24, q_arr_7__23, q_arr_7__22, q_arr_7__21, 
                             q_arr_7__20, q_arr_7__19, q_arr_7__18, q_arr_7__17, 
                             q_arr_7__16, q_arr_7__15, q_arr_7__14, q_arr_7__13, 
                             q_arr_7__12, q_arr_7__11, q_arr_7__10, q_arr_7__9, 
                             q_arr_7__8, q_arr_7__7, q_arr_7__6, q_arr_7__5, 
                             q_arr_7__4, q_arr_7__3, q_arr_7__2, q_arr_7__1, 
                             q_arr_7__0, q_arr_8__31, q_arr_8__30, q_arr_8__29, 
                             q_arr_8__28, q_arr_8__27, q_arr_8__26, q_arr_8__25, 
                             q_arr_8__24, q_arr_8__23, q_arr_8__22, q_arr_8__21, 
                             q_arr_8__20, q_arr_8__19, q_arr_8__18, q_arr_8__17, 
                             q_arr_8__16, q_arr_8__15, q_arr_8__14, q_arr_8__13, 
                             q_arr_8__12, q_arr_8__11, q_arr_8__10, q_arr_8__9, 
                             q_arr_8__8, q_arr_8__7, q_arr_8__6, q_arr_8__5, 
                             q_arr_8__4, q_arr_8__3, q_arr_8__2, q_arr_8__1, 
                             q_arr_8__0, q_arr_9__31, q_arr_9__30, q_arr_9__29, 
                             q_arr_9__28, q_arr_9__27, q_arr_9__26, q_arr_9__25, 
                             q_arr_9__24, q_arr_9__23, q_arr_9__22, q_arr_9__21, 
                             q_arr_9__20, q_arr_9__19, q_arr_9__18, q_arr_9__17, 
                             q_arr_9__16, q_arr_9__15, q_arr_9__14, q_arr_9__13, 
                             q_arr_9__12, q_arr_9__11, q_arr_9__10, q_arr_9__9, 
                             q_arr_9__8, q_arr_9__7, q_arr_9__6, q_arr_9__5, 
                             q_arr_9__4, q_arr_9__3, q_arr_9__2, q_arr_9__1, 
                             q_arr_9__0, q_arr_10__31, q_arr_10__30, 
                             q_arr_10__29, q_arr_10__28, q_arr_10__27, 
                             q_arr_10__26, q_arr_10__25, q_arr_10__24, 
                             q_arr_10__23, q_arr_10__22, q_arr_10__21, 
                             q_arr_10__20, q_arr_10__19, q_arr_10__18, 
                             q_arr_10__17, q_arr_10__16, q_arr_10__15, 
                             q_arr_10__14, q_arr_10__13, q_arr_10__12, 
                             q_arr_10__11, q_arr_10__10, q_arr_10__9, 
                             q_arr_10__8, q_arr_10__7, q_arr_10__6, q_arr_10__5, 
                             q_arr_10__4, q_arr_10__3, q_arr_10__2, q_arr_10__1, 
                             q_arr_10__0, q_arr_11__31, q_arr_11__30, 
                             q_arr_11__29, q_arr_11__28, q_arr_11__27, 
                             q_arr_11__26, q_arr_11__25, q_arr_11__24, 
                             q_arr_11__23, q_arr_11__22, q_arr_11__21, 
                             q_arr_11__20, q_arr_11__19, q_arr_11__18, 
                             q_arr_11__17, q_arr_11__16, q_arr_11__15, 
                             q_arr_11__14, q_arr_11__13, q_arr_11__12, 
                             q_arr_11__11, q_arr_11__10, q_arr_11__9, 
                             q_arr_11__8, q_arr_11__7, q_arr_11__6, q_arr_11__5, 
                             q_arr_11__4, q_arr_11__3, q_arr_11__2, q_arr_11__1, 
                             q_arr_11__0, q_arr_12__31, q_arr_12__30, 
                             q_arr_12__29, q_arr_12__28, q_arr_12__27, 
                             q_arr_12__26, q_arr_12__25, q_arr_12__24, 
                             q_arr_12__23, q_arr_12__22, q_arr_12__21, 
                             q_arr_12__20, q_arr_12__19, q_arr_12__18, 
                             q_arr_12__17, q_arr_12__16, q_arr_12__15, 
                             q_arr_12__14, q_arr_12__13, q_arr_12__12, 
                             q_arr_12__11, q_arr_12__10, q_arr_12__9, 
                             q_arr_12__8, q_arr_12__7, q_arr_12__6, q_arr_12__5, 
                             q_arr_12__4, q_arr_12__3, q_arr_12__2, q_arr_12__1, 
                             q_arr_12__0, q_arr_13__31, q_arr_13__30, 
                             q_arr_13__29, q_arr_13__28, q_arr_13__27, 
                             q_arr_13__26, q_arr_13__25, q_arr_13__24, 
                             q_arr_13__23, q_arr_13__22, q_arr_13__21, 
                             q_arr_13__20, q_arr_13__19, q_arr_13__18, 
                             q_arr_13__17, q_arr_13__16, q_arr_13__15, 
                             q_arr_13__14, q_arr_13__13, q_arr_13__12, 
                             q_arr_13__11, q_arr_13__10, q_arr_13__9, 
                             q_arr_13__8, q_arr_13__7, q_arr_13__6, q_arr_13__5, 
                             q_arr_13__4, q_arr_13__3, q_arr_13__2, q_arr_13__1, 
                             q_arr_13__0, q_arr_14__31, q_arr_14__30, 
                             q_arr_14__29, q_arr_14__28, q_arr_14__27, 
                             q_arr_14__26, q_arr_14__25, q_arr_14__24, 
                             q_arr_14__23, q_arr_14__22, q_arr_14__21, 
                             q_arr_14__20, q_arr_14__19, q_arr_14__18, 
                             q_arr_14__17, q_arr_14__16, q_arr_14__15, 
                             q_arr_14__14, q_arr_14__13, q_arr_14__12, 
                             q_arr_14__11, q_arr_14__10, q_arr_14__9, 
                             q_arr_14__8, q_arr_14__7, q_arr_14__6, q_arr_14__5, 
                             q_arr_14__4, q_arr_14__3, q_arr_14__2, q_arr_14__1, 
                             q_arr_14__0, q_arr_15__31, q_arr_15__30, 
                             q_arr_15__29, q_arr_15__28, q_arr_15__27, 
                             q_arr_15__26, q_arr_15__25, q_arr_15__24, 
                             q_arr_15__23, q_arr_15__22, q_arr_15__21, 
                             q_arr_15__20, q_arr_15__19, q_arr_15__18, 
                             q_arr_15__17, q_arr_15__16, q_arr_15__15, 
                             q_arr_15__14, q_arr_15__13, q_arr_15__12, 
                             q_arr_15__11, q_arr_15__10, q_arr_15__9, 
                             q_arr_15__8, q_arr_15__7, q_arr_15__6, q_arr_15__5, 
                             q_arr_15__4, q_arr_15__3, q_arr_15__2, q_arr_15__1, 
                             q_arr_15__0, q_arr_16__31, q_arr_16__30, 
                             q_arr_16__29, q_arr_16__28, q_arr_16__27, 
                             q_arr_16__26, q_arr_16__25, q_arr_16__24, 
                             q_arr_16__23, q_arr_16__22, q_arr_16__21, 
                             q_arr_16__20, q_arr_16__19, q_arr_16__18, 
                             q_arr_16__17, q_arr_16__16, q_arr_16__15, 
                             q_arr_16__14, q_arr_16__13, q_arr_16__12, 
                             q_arr_16__11, q_arr_16__10, q_arr_16__9, 
                             q_arr_16__8, q_arr_16__7, q_arr_16__6, q_arr_16__5, 
                             q_arr_16__4, q_arr_16__3, q_arr_16__2, q_arr_16__1, 
                             q_arr_16__0, q_arr_17__31, q_arr_17__30, 
                             q_arr_17__29, q_arr_17__28, q_arr_17__27, 
                             q_arr_17__26, q_arr_17__25, q_arr_17__24, 
                             q_arr_17__23, q_arr_17__22, q_arr_17__21, 
                             q_arr_17__20, q_arr_17__19, q_arr_17__18, 
                             q_arr_17__17, q_arr_17__16, q_arr_17__15, 
                             q_arr_17__14, q_arr_17__13, q_arr_17__12, 
                             q_arr_17__11, q_arr_17__10, q_arr_17__9, 
                             q_arr_17__8, q_arr_17__7, q_arr_17__6, q_arr_17__5, 
                             q_arr_17__4, q_arr_17__3, q_arr_17__2, q_arr_17__1, 
                             q_arr_17__0, q_arr_18__31, q_arr_18__30, 
                             q_arr_18__29, q_arr_18__28, q_arr_18__27, 
                             q_arr_18__26, q_arr_18__25, q_arr_18__24, 
                             q_arr_18__23, q_arr_18__22, q_arr_18__21, 
                             q_arr_18__20, q_arr_18__19, q_arr_18__18, 
                             q_arr_18__17, q_arr_18__16, q_arr_18__15, 
                             q_arr_18__14, q_arr_18__13, q_arr_18__12, 
                             q_arr_18__11, q_arr_18__10, q_arr_18__9, 
                             q_arr_18__8, q_arr_18__7, q_arr_18__6, q_arr_18__5, 
                             q_arr_18__4, q_arr_18__3, q_arr_18__2, q_arr_18__1, 
                             q_arr_18__0, q_arr_19__31, q_arr_19__30, 
                             q_arr_19__29, q_arr_19__28, q_arr_19__27, 
                             q_arr_19__26, q_arr_19__25, q_arr_19__24, 
                             q_arr_19__23, q_arr_19__22, q_arr_19__21, 
                             q_arr_19__20, q_arr_19__19, q_arr_19__18, 
                             q_arr_19__17, q_arr_19__16, q_arr_19__15, 
                             q_arr_19__14, q_arr_19__13, q_arr_19__12, 
                             q_arr_19__11, q_arr_19__10, q_arr_19__9, 
                             q_arr_19__8, q_arr_19__7, q_arr_19__6, q_arr_19__5, 
                             q_arr_19__4, q_arr_19__3, q_arr_19__2, q_arr_19__1, 
                             q_arr_19__0, q_arr_20__31, q_arr_20__30, 
                             q_arr_20__29, q_arr_20__28, q_arr_20__27, 
                             q_arr_20__26, q_arr_20__25, q_arr_20__24, 
                             q_arr_20__23, q_arr_20__22, q_arr_20__21, 
                             q_arr_20__20, q_arr_20__19, q_arr_20__18, 
                             q_arr_20__17, q_arr_20__16, q_arr_20__15, 
                             q_arr_20__14, q_arr_20__13, q_arr_20__12, 
                             q_arr_20__11, q_arr_20__10, q_arr_20__9, 
                             q_arr_20__8, q_arr_20__7, q_arr_20__6, q_arr_20__5, 
                             q_arr_20__4, q_arr_20__3, q_arr_20__2, q_arr_20__1, 
                             q_arr_20__0, q_arr_21__31, q_arr_21__30, 
                             q_arr_21__29, q_arr_21__28, q_arr_21__27, 
                             q_arr_21__26, q_arr_21__25, q_arr_21__24, 
                             q_arr_21__23, q_arr_21__22, q_arr_21__21, 
                             q_arr_21__20, q_arr_21__19, q_arr_21__18, 
                             q_arr_21__17, q_arr_21__16, q_arr_21__15, 
                             q_arr_21__14, q_arr_21__13, q_arr_21__12, 
                             q_arr_21__11, q_arr_21__10, q_arr_21__9, 
                             q_arr_21__8, q_arr_21__7, q_arr_21__6, q_arr_21__5, 
                             q_arr_21__4, q_arr_21__3, q_arr_21__2, q_arr_21__1, 
                             q_arr_21__0, q_arr_22__31, q_arr_22__30, 
                             q_arr_22__29, q_arr_22__28, q_arr_22__27, 
                             q_arr_22__26, q_arr_22__25, q_arr_22__24, 
                             q_arr_22__23, q_arr_22__22, q_arr_22__21, 
                             q_arr_22__20, q_arr_22__19, q_arr_22__18, 
                             q_arr_22__17, q_arr_22__16, q_arr_22__15, 
                             q_arr_22__14, q_arr_22__13, q_arr_22__12, 
                             q_arr_22__11, q_arr_22__10, q_arr_22__9, 
                             q_arr_22__8, q_arr_22__7, q_arr_22__6, q_arr_22__5, 
                             q_arr_22__4, q_arr_22__3, q_arr_22__2, q_arr_22__1, 
                             q_arr_22__0, q_arr_23__31, q_arr_23__30, 
                             q_arr_23__29, q_arr_23__28, q_arr_23__27, 
                             q_arr_23__26, q_arr_23__25, q_arr_23__24, 
                             q_arr_23__23, q_arr_23__22, q_arr_23__21, 
                             q_arr_23__20, q_arr_23__19, q_arr_23__18, 
                             q_arr_23__17, q_arr_23__16, q_arr_23__15, 
                             q_arr_23__14, q_arr_23__13, q_arr_23__12, 
                             q_arr_23__11, q_arr_23__10, q_arr_23__9, 
                             q_arr_23__8, q_arr_23__7, q_arr_23__6, q_arr_23__5, 
                             q_arr_23__4, q_arr_23__3, q_arr_23__2, q_arr_23__1, 
                             q_arr_23__0, q_arr_24__31, q_arr_24__30, 
                             q_arr_24__29, q_arr_24__28, q_arr_24__27, 
                             q_arr_24__26, q_arr_24__25, q_arr_24__24, 
                             q_arr_24__23, q_arr_24__22, q_arr_24__21, 
                             q_arr_24__20, q_arr_24__19, q_arr_24__18, 
                             q_arr_24__17, q_arr_24__16, q_arr_24__15, 
                             q_arr_24__14, q_arr_24__13, q_arr_24__12, 
                             q_arr_24__11, q_arr_24__10, q_arr_24__9, 
                             q_arr_24__8, q_arr_24__7, q_arr_24__6, q_arr_24__5, 
                             q_arr_24__4, q_arr_24__3, q_arr_24__2, q_arr_24__1, 
                             q_arr_24__0, output1_init, output2_init, 
                             filter_size, operation, compute_relu, clk, en, 
                             reset, buffer_ready, semi_ready, ready ) ;

    input img_data_0__15 ;
    input img_data_0__14 ;
    input img_data_0__13 ;
    input img_data_0__12 ;
    input img_data_0__11 ;
    input img_data_0__10 ;
    input img_data_0__9 ;
    input img_data_0__8 ;
    input img_data_0__7 ;
    input img_data_0__6 ;
    input img_data_0__5 ;
    input img_data_0__4 ;
    input img_data_0__3 ;
    input img_data_0__2 ;
    input img_data_0__1 ;
    input img_data_0__0 ;
    input img_data_1__15 ;
    input img_data_1__14 ;
    input img_data_1__13 ;
    input img_data_1__12 ;
    input img_data_1__11 ;
    input img_data_1__10 ;
    input img_data_1__9 ;
    input img_data_1__8 ;
    input img_data_1__7 ;
    input img_data_1__6 ;
    input img_data_1__5 ;
    input img_data_1__4 ;
    input img_data_1__3 ;
    input img_data_1__2 ;
    input img_data_1__1 ;
    input img_data_1__0 ;
    input img_data_2__15 ;
    input img_data_2__14 ;
    input img_data_2__13 ;
    input img_data_2__12 ;
    input img_data_2__11 ;
    input img_data_2__10 ;
    input img_data_2__9 ;
    input img_data_2__8 ;
    input img_data_2__7 ;
    input img_data_2__6 ;
    input img_data_2__5 ;
    input img_data_2__4 ;
    input img_data_2__3 ;
    input img_data_2__2 ;
    input img_data_2__1 ;
    input img_data_2__0 ;
    input img_data_3__15 ;
    input img_data_3__14 ;
    input img_data_3__13 ;
    input img_data_3__12 ;
    input img_data_3__11 ;
    input img_data_3__10 ;
    input img_data_3__9 ;
    input img_data_3__8 ;
    input img_data_3__7 ;
    input img_data_3__6 ;
    input img_data_3__5 ;
    input img_data_3__4 ;
    input img_data_3__3 ;
    input img_data_3__2 ;
    input img_data_3__1 ;
    input img_data_3__0 ;
    input img_data_4__15 ;
    input img_data_4__14 ;
    input img_data_4__13 ;
    input img_data_4__12 ;
    input img_data_4__11 ;
    input img_data_4__10 ;
    input img_data_4__9 ;
    input img_data_4__8 ;
    input img_data_4__7 ;
    input img_data_4__6 ;
    input img_data_4__5 ;
    input img_data_4__4 ;
    input img_data_4__3 ;
    input img_data_4__2 ;
    input img_data_4__1 ;
    input img_data_4__0 ;
    input img_data_5__15 ;
    input img_data_5__14 ;
    input img_data_5__13 ;
    input img_data_5__12 ;
    input img_data_5__11 ;
    input img_data_5__10 ;
    input img_data_5__9 ;
    input img_data_5__8 ;
    input img_data_5__7 ;
    input img_data_5__6 ;
    input img_data_5__5 ;
    input img_data_5__4 ;
    input img_data_5__3 ;
    input img_data_5__2 ;
    input img_data_5__1 ;
    input img_data_5__0 ;
    input img_data_6__15 ;
    input img_data_6__14 ;
    input img_data_6__13 ;
    input img_data_6__12 ;
    input img_data_6__11 ;
    input img_data_6__10 ;
    input img_data_6__9 ;
    input img_data_6__8 ;
    input img_data_6__7 ;
    input img_data_6__6 ;
    input img_data_6__5 ;
    input img_data_6__4 ;
    input img_data_6__3 ;
    input img_data_6__2 ;
    input img_data_6__1 ;
    input img_data_6__0 ;
    input img_data_7__15 ;
    input img_data_7__14 ;
    input img_data_7__13 ;
    input img_data_7__12 ;
    input img_data_7__11 ;
    input img_data_7__10 ;
    input img_data_7__9 ;
    input img_data_7__8 ;
    input img_data_7__7 ;
    input img_data_7__6 ;
    input img_data_7__5 ;
    input img_data_7__4 ;
    input img_data_7__3 ;
    input img_data_7__2 ;
    input img_data_7__1 ;
    input img_data_7__0 ;
    input img_data_8__15 ;
    input img_data_8__14 ;
    input img_data_8__13 ;
    input img_data_8__12 ;
    input img_data_8__11 ;
    input img_data_8__10 ;
    input img_data_8__9 ;
    input img_data_8__8 ;
    input img_data_8__7 ;
    input img_data_8__6 ;
    input img_data_8__5 ;
    input img_data_8__4 ;
    input img_data_8__3 ;
    input img_data_8__2 ;
    input img_data_8__1 ;
    input img_data_8__0 ;
    input img_data_9__15 ;
    input img_data_9__14 ;
    input img_data_9__13 ;
    input img_data_9__12 ;
    input img_data_9__11 ;
    input img_data_9__10 ;
    input img_data_9__9 ;
    input img_data_9__8 ;
    input img_data_9__7 ;
    input img_data_9__6 ;
    input img_data_9__5 ;
    input img_data_9__4 ;
    input img_data_9__3 ;
    input img_data_9__2 ;
    input img_data_9__1 ;
    input img_data_9__0 ;
    input img_data_10__15 ;
    input img_data_10__14 ;
    input img_data_10__13 ;
    input img_data_10__12 ;
    input img_data_10__11 ;
    input img_data_10__10 ;
    input img_data_10__9 ;
    input img_data_10__8 ;
    input img_data_10__7 ;
    input img_data_10__6 ;
    input img_data_10__5 ;
    input img_data_10__4 ;
    input img_data_10__3 ;
    input img_data_10__2 ;
    input img_data_10__1 ;
    input img_data_10__0 ;
    input img_data_11__15 ;
    input img_data_11__14 ;
    input img_data_11__13 ;
    input img_data_11__12 ;
    input img_data_11__11 ;
    input img_data_11__10 ;
    input img_data_11__9 ;
    input img_data_11__8 ;
    input img_data_11__7 ;
    input img_data_11__6 ;
    input img_data_11__5 ;
    input img_data_11__4 ;
    input img_data_11__3 ;
    input img_data_11__2 ;
    input img_data_11__1 ;
    input img_data_11__0 ;
    input img_data_12__15 ;
    input img_data_12__14 ;
    input img_data_12__13 ;
    input img_data_12__12 ;
    input img_data_12__11 ;
    input img_data_12__10 ;
    input img_data_12__9 ;
    input img_data_12__8 ;
    input img_data_12__7 ;
    input img_data_12__6 ;
    input img_data_12__5 ;
    input img_data_12__4 ;
    input img_data_12__3 ;
    input img_data_12__2 ;
    input img_data_12__1 ;
    input img_data_12__0 ;
    input img_data_13__15 ;
    input img_data_13__14 ;
    input img_data_13__13 ;
    input img_data_13__12 ;
    input img_data_13__11 ;
    input img_data_13__10 ;
    input img_data_13__9 ;
    input img_data_13__8 ;
    input img_data_13__7 ;
    input img_data_13__6 ;
    input img_data_13__5 ;
    input img_data_13__4 ;
    input img_data_13__3 ;
    input img_data_13__2 ;
    input img_data_13__1 ;
    input img_data_13__0 ;
    input img_data_14__15 ;
    input img_data_14__14 ;
    input img_data_14__13 ;
    input img_data_14__12 ;
    input img_data_14__11 ;
    input img_data_14__10 ;
    input img_data_14__9 ;
    input img_data_14__8 ;
    input img_data_14__7 ;
    input img_data_14__6 ;
    input img_data_14__5 ;
    input img_data_14__4 ;
    input img_data_14__3 ;
    input img_data_14__2 ;
    input img_data_14__1 ;
    input img_data_14__0 ;
    input img_data_15__15 ;
    input img_data_15__14 ;
    input img_data_15__13 ;
    input img_data_15__12 ;
    input img_data_15__11 ;
    input img_data_15__10 ;
    input img_data_15__9 ;
    input img_data_15__8 ;
    input img_data_15__7 ;
    input img_data_15__6 ;
    input img_data_15__5 ;
    input img_data_15__4 ;
    input img_data_15__3 ;
    input img_data_15__2 ;
    input img_data_15__1 ;
    input img_data_15__0 ;
    input img_data_16__15 ;
    input img_data_16__14 ;
    input img_data_16__13 ;
    input img_data_16__12 ;
    input img_data_16__11 ;
    input img_data_16__10 ;
    input img_data_16__9 ;
    input img_data_16__8 ;
    input img_data_16__7 ;
    input img_data_16__6 ;
    input img_data_16__5 ;
    input img_data_16__4 ;
    input img_data_16__3 ;
    input img_data_16__2 ;
    input img_data_16__1 ;
    input img_data_16__0 ;
    input img_data_17__15 ;
    input img_data_17__14 ;
    input img_data_17__13 ;
    input img_data_17__12 ;
    input img_data_17__11 ;
    input img_data_17__10 ;
    input img_data_17__9 ;
    input img_data_17__8 ;
    input img_data_17__7 ;
    input img_data_17__6 ;
    input img_data_17__5 ;
    input img_data_17__4 ;
    input img_data_17__3 ;
    input img_data_17__2 ;
    input img_data_17__1 ;
    input img_data_17__0 ;
    input img_data_18__15 ;
    input img_data_18__14 ;
    input img_data_18__13 ;
    input img_data_18__12 ;
    input img_data_18__11 ;
    input img_data_18__10 ;
    input img_data_18__9 ;
    input img_data_18__8 ;
    input img_data_18__7 ;
    input img_data_18__6 ;
    input img_data_18__5 ;
    input img_data_18__4 ;
    input img_data_18__3 ;
    input img_data_18__2 ;
    input img_data_18__1 ;
    input img_data_18__0 ;
    input img_data_19__15 ;
    input img_data_19__14 ;
    input img_data_19__13 ;
    input img_data_19__12 ;
    input img_data_19__11 ;
    input img_data_19__10 ;
    input img_data_19__9 ;
    input img_data_19__8 ;
    input img_data_19__7 ;
    input img_data_19__6 ;
    input img_data_19__5 ;
    input img_data_19__4 ;
    input img_data_19__3 ;
    input img_data_19__2 ;
    input img_data_19__1 ;
    input img_data_19__0 ;
    input img_data_20__15 ;
    input img_data_20__14 ;
    input img_data_20__13 ;
    input img_data_20__12 ;
    input img_data_20__11 ;
    input img_data_20__10 ;
    input img_data_20__9 ;
    input img_data_20__8 ;
    input img_data_20__7 ;
    input img_data_20__6 ;
    input img_data_20__5 ;
    input img_data_20__4 ;
    input img_data_20__3 ;
    input img_data_20__2 ;
    input img_data_20__1 ;
    input img_data_20__0 ;
    input img_data_21__15 ;
    input img_data_21__14 ;
    input img_data_21__13 ;
    input img_data_21__12 ;
    input img_data_21__11 ;
    input img_data_21__10 ;
    input img_data_21__9 ;
    input img_data_21__8 ;
    input img_data_21__7 ;
    input img_data_21__6 ;
    input img_data_21__5 ;
    input img_data_21__4 ;
    input img_data_21__3 ;
    input img_data_21__2 ;
    input img_data_21__1 ;
    input img_data_21__0 ;
    input img_data_22__15 ;
    input img_data_22__14 ;
    input img_data_22__13 ;
    input img_data_22__12 ;
    input img_data_22__11 ;
    input img_data_22__10 ;
    input img_data_22__9 ;
    input img_data_22__8 ;
    input img_data_22__7 ;
    input img_data_22__6 ;
    input img_data_22__5 ;
    input img_data_22__4 ;
    input img_data_22__3 ;
    input img_data_22__2 ;
    input img_data_22__1 ;
    input img_data_22__0 ;
    input img_data_23__15 ;
    input img_data_23__14 ;
    input img_data_23__13 ;
    input img_data_23__12 ;
    input img_data_23__11 ;
    input img_data_23__10 ;
    input img_data_23__9 ;
    input img_data_23__8 ;
    input img_data_23__7 ;
    input img_data_23__6 ;
    input img_data_23__5 ;
    input img_data_23__4 ;
    input img_data_23__3 ;
    input img_data_23__2 ;
    input img_data_23__1 ;
    input img_data_23__0 ;
    input img_data_24__15 ;
    input img_data_24__14 ;
    input img_data_24__13 ;
    input img_data_24__12 ;
    input img_data_24__11 ;
    input img_data_24__10 ;
    input img_data_24__9 ;
    input img_data_24__8 ;
    input img_data_24__7 ;
    input img_data_24__6 ;
    input img_data_24__5 ;
    input img_data_24__4 ;
    input img_data_24__3 ;
    input img_data_24__2 ;
    input img_data_24__1 ;
    input img_data_24__0 ;
    input filter_data_0__15 ;
    input filter_data_0__14 ;
    input filter_data_0__13 ;
    input filter_data_0__12 ;
    input filter_data_0__11 ;
    input filter_data_0__10 ;
    input filter_data_0__9 ;
    input filter_data_0__8 ;
    input filter_data_0__7 ;
    input filter_data_0__6 ;
    input filter_data_0__5 ;
    input filter_data_0__4 ;
    input filter_data_0__3 ;
    input filter_data_0__2 ;
    input filter_data_0__1 ;
    input filter_data_0__0 ;
    input filter_data_1__15 ;
    input filter_data_1__14 ;
    input filter_data_1__13 ;
    input filter_data_1__12 ;
    input filter_data_1__11 ;
    input filter_data_1__10 ;
    input filter_data_1__9 ;
    input filter_data_1__8 ;
    input filter_data_1__7 ;
    input filter_data_1__6 ;
    input filter_data_1__5 ;
    input filter_data_1__4 ;
    input filter_data_1__3 ;
    input filter_data_1__2 ;
    input filter_data_1__1 ;
    input filter_data_1__0 ;
    input filter_data_2__15 ;
    input filter_data_2__14 ;
    input filter_data_2__13 ;
    input filter_data_2__12 ;
    input filter_data_2__11 ;
    input filter_data_2__10 ;
    input filter_data_2__9 ;
    input filter_data_2__8 ;
    input filter_data_2__7 ;
    input filter_data_2__6 ;
    input filter_data_2__5 ;
    input filter_data_2__4 ;
    input filter_data_2__3 ;
    input filter_data_2__2 ;
    input filter_data_2__1 ;
    input filter_data_2__0 ;
    input filter_data_3__15 ;
    input filter_data_3__14 ;
    input filter_data_3__13 ;
    input filter_data_3__12 ;
    input filter_data_3__11 ;
    input filter_data_3__10 ;
    input filter_data_3__9 ;
    input filter_data_3__8 ;
    input filter_data_3__7 ;
    input filter_data_3__6 ;
    input filter_data_3__5 ;
    input filter_data_3__4 ;
    input filter_data_3__3 ;
    input filter_data_3__2 ;
    input filter_data_3__1 ;
    input filter_data_3__0 ;
    input filter_data_4__15 ;
    input filter_data_4__14 ;
    input filter_data_4__13 ;
    input filter_data_4__12 ;
    input filter_data_4__11 ;
    input filter_data_4__10 ;
    input filter_data_4__9 ;
    input filter_data_4__8 ;
    input filter_data_4__7 ;
    input filter_data_4__6 ;
    input filter_data_4__5 ;
    input filter_data_4__4 ;
    input filter_data_4__3 ;
    input filter_data_4__2 ;
    input filter_data_4__1 ;
    input filter_data_4__0 ;
    input filter_data_5__15 ;
    input filter_data_5__14 ;
    input filter_data_5__13 ;
    input filter_data_5__12 ;
    input filter_data_5__11 ;
    input filter_data_5__10 ;
    input filter_data_5__9 ;
    input filter_data_5__8 ;
    input filter_data_5__7 ;
    input filter_data_5__6 ;
    input filter_data_5__5 ;
    input filter_data_5__4 ;
    input filter_data_5__3 ;
    input filter_data_5__2 ;
    input filter_data_5__1 ;
    input filter_data_5__0 ;
    input filter_data_6__15 ;
    input filter_data_6__14 ;
    input filter_data_6__13 ;
    input filter_data_6__12 ;
    input filter_data_6__11 ;
    input filter_data_6__10 ;
    input filter_data_6__9 ;
    input filter_data_6__8 ;
    input filter_data_6__7 ;
    input filter_data_6__6 ;
    input filter_data_6__5 ;
    input filter_data_6__4 ;
    input filter_data_6__3 ;
    input filter_data_6__2 ;
    input filter_data_6__1 ;
    input filter_data_6__0 ;
    input filter_data_7__15 ;
    input filter_data_7__14 ;
    input filter_data_7__13 ;
    input filter_data_7__12 ;
    input filter_data_7__11 ;
    input filter_data_7__10 ;
    input filter_data_7__9 ;
    input filter_data_7__8 ;
    input filter_data_7__7 ;
    input filter_data_7__6 ;
    input filter_data_7__5 ;
    input filter_data_7__4 ;
    input filter_data_7__3 ;
    input filter_data_7__2 ;
    input filter_data_7__1 ;
    input filter_data_7__0 ;
    input filter_data_8__15 ;
    input filter_data_8__14 ;
    input filter_data_8__13 ;
    input filter_data_8__12 ;
    input filter_data_8__11 ;
    input filter_data_8__10 ;
    input filter_data_8__9 ;
    input filter_data_8__8 ;
    input filter_data_8__7 ;
    input filter_data_8__6 ;
    input filter_data_8__5 ;
    input filter_data_8__4 ;
    input filter_data_8__3 ;
    input filter_data_8__2 ;
    input filter_data_8__1 ;
    input filter_data_8__0 ;
    input filter_data_9__15 ;
    input filter_data_9__14 ;
    input filter_data_9__13 ;
    input filter_data_9__12 ;
    input filter_data_9__11 ;
    input filter_data_9__10 ;
    input filter_data_9__9 ;
    input filter_data_9__8 ;
    input filter_data_9__7 ;
    input filter_data_9__6 ;
    input filter_data_9__5 ;
    input filter_data_9__4 ;
    input filter_data_9__3 ;
    input filter_data_9__2 ;
    input filter_data_9__1 ;
    input filter_data_9__0 ;
    input filter_data_10__15 ;
    input filter_data_10__14 ;
    input filter_data_10__13 ;
    input filter_data_10__12 ;
    input filter_data_10__11 ;
    input filter_data_10__10 ;
    input filter_data_10__9 ;
    input filter_data_10__8 ;
    input filter_data_10__7 ;
    input filter_data_10__6 ;
    input filter_data_10__5 ;
    input filter_data_10__4 ;
    input filter_data_10__3 ;
    input filter_data_10__2 ;
    input filter_data_10__1 ;
    input filter_data_10__0 ;
    input filter_data_11__15 ;
    input filter_data_11__14 ;
    input filter_data_11__13 ;
    input filter_data_11__12 ;
    input filter_data_11__11 ;
    input filter_data_11__10 ;
    input filter_data_11__9 ;
    input filter_data_11__8 ;
    input filter_data_11__7 ;
    input filter_data_11__6 ;
    input filter_data_11__5 ;
    input filter_data_11__4 ;
    input filter_data_11__3 ;
    input filter_data_11__2 ;
    input filter_data_11__1 ;
    input filter_data_11__0 ;
    input filter_data_12__15 ;
    input filter_data_12__14 ;
    input filter_data_12__13 ;
    input filter_data_12__12 ;
    input filter_data_12__11 ;
    input filter_data_12__10 ;
    input filter_data_12__9 ;
    input filter_data_12__8 ;
    input filter_data_12__7 ;
    input filter_data_12__6 ;
    input filter_data_12__5 ;
    input filter_data_12__4 ;
    input filter_data_12__3 ;
    input filter_data_12__2 ;
    input filter_data_12__1 ;
    input filter_data_12__0 ;
    input filter_data_13__15 ;
    input filter_data_13__14 ;
    input filter_data_13__13 ;
    input filter_data_13__12 ;
    input filter_data_13__11 ;
    input filter_data_13__10 ;
    input filter_data_13__9 ;
    input filter_data_13__8 ;
    input filter_data_13__7 ;
    input filter_data_13__6 ;
    input filter_data_13__5 ;
    input filter_data_13__4 ;
    input filter_data_13__3 ;
    input filter_data_13__2 ;
    input filter_data_13__1 ;
    input filter_data_13__0 ;
    input filter_data_14__15 ;
    input filter_data_14__14 ;
    input filter_data_14__13 ;
    input filter_data_14__12 ;
    input filter_data_14__11 ;
    input filter_data_14__10 ;
    input filter_data_14__9 ;
    input filter_data_14__8 ;
    input filter_data_14__7 ;
    input filter_data_14__6 ;
    input filter_data_14__5 ;
    input filter_data_14__4 ;
    input filter_data_14__3 ;
    input filter_data_14__2 ;
    input filter_data_14__1 ;
    input filter_data_14__0 ;
    input filter_data_15__15 ;
    input filter_data_15__14 ;
    input filter_data_15__13 ;
    input filter_data_15__12 ;
    input filter_data_15__11 ;
    input filter_data_15__10 ;
    input filter_data_15__9 ;
    input filter_data_15__8 ;
    input filter_data_15__7 ;
    input filter_data_15__6 ;
    input filter_data_15__5 ;
    input filter_data_15__4 ;
    input filter_data_15__3 ;
    input filter_data_15__2 ;
    input filter_data_15__1 ;
    input filter_data_15__0 ;
    input filter_data_16__15 ;
    input filter_data_16__14 ;
    input filter_data_16__13 ;
    input filter_data_16__12 ;
    input filter_data_16__11 ;
    input filter_data_16__10 ;
    input filter_data_16__9 ;
    input filter_data_16__8 ;
    input filter_data_16__7 ;
    input filter_data_16__6 ;
    input filter_data_16__5 ;
    input filter_data_16__4 ;
    input filter_data_16__3 ;
    input filter_data_16__2 ;
    input filter_data_16__1 ;
    input filter_data_16__0 ;
    input filter_data_17__15 ;
    input filter_data_17__14 ;
    input filter_data_17__13 ;
    input filter_data_17__12 ;
    input filter_data_17__11 ;
    input filter_data_17__10 ;
    input filter_data_17__9 ;
    input filter_data_17__8 ;
    input filter_data_17__7 ;
    input filter_data_17__6 ;
    input filter_data_17__5 ;
    input filter_data_17__4 ;
    input filter_data_17__3 ;
    input filter_data_17__2 ;
    input filter_data_17__1 ;
    input filter_data_17__0 ;
    input filter_data_18__15 ;
    input filter_data_18__14 ;
    input filter_data_18__13 ;
    input filter_data_18__12 ;
    input filter_data_18__11 ;
    input filter_data_18__10 ;
    input filter_data_18__9 ;
    input filter_data_18__8 ;
    input filter_data_18__7 ;
    input filter_data_18__6 ;
    input filter_data_18__5 ;
    input filter_data_18__4 ;
    input filter_data_18__3 ;
    input filter_data_18__2 ;
    input filter_data_18__1 ;
    input filter_data_18__0 ;
    input filter_data_19__15 ;
    input filter_data_19__14 ;
    input filter_data_19__13 ;
    input filter_data_19__12 ;
    input filter_data_19__11 ;
    input filter_data_19__10 ;
    input filter_data_19__9 ;
    input filter_data_19__8 ;
    input filter_data_19__7 ;
    input filter_data_19__6 ;
    input filter_data_19__5 ;
    input filter_data_19__4 ;
    input filter_data_19__3 ;
    input filter_data_19__2 ;
    input filter_data_19__1 ;
    input filter_data_19__0 ;
    input filter_data_20__15 ;
    input filter_data_20__14 ;
    input filter_data_20__13 ;
    input filter_data_20__12 ;
    input filter_data_20__11 ;
    input filter_data_20__10 ;
    input filter_data_20__9 ;
    input filter_data_20__8 ;
    input filter_data_20__7 ;
    input filter_data_20__6 ;
    input filter_data_20__5 ;
    input filter_data_20__4 ;
    input filter_data_20__3 ;
    input filter_data_20__2 ;
    input filter_data_20__1 ;
    input filter_data_20__0 ;
    input filter_data_21__15 ;
    input filter_data_21__14 ;
    input filter_data_21__13 ;
    input filter_data_21__12 ;
    input filter_data_21__11 ;
    input filter_data_21__10 ;
    input filter_data_21__9 ;
    input filter_data_21__8 ;
    input filter_data_21__7 ;
    input filter_data_21__6 ;
    input filter_data_21__5 ;
    input filter_data_21__4 ;
    input filter_data_21__3 ;
    input filter_data_21__2 ;
    input filter_data_21__1 ;
    input filter_data_21__0 ;
    input filter_data_22__15 ;
    input filter_data_22__14 ;
    input filter_data_22__13 ;
    input filter_data_22__12 ;
    input filter_data_22__11 ;
    input filter_data_22__10 ;
    input filter_data_22__9 ;
    input filter_data_22__8 ;
    input filter_data_22__7 ;
    input filter_data_22__6 ;
    input filter_data_22__5 ;
    input filter_data_22__4 ;
    input filter_data_22__3 ;
    input filter_data_22__2 ;
    input filter_data_22__1 ;
    input filter_data_22__0 ;
    input filter_data_23__15 ;
    input filter_data_23__14 ;
    input filter_data_23__13 ;
    input filter_data_23__12 ;
    input filter_data_23__11 ;
    input filter_data_23__10 ;
    input filter_data_23__9 ;
    input filter_data_23__8 ;
    input filter_data_23__7 ;
    input filter_data_23__6 ;
    input filter_data_23__5 ;
    input filter_data_23__4 ;
    input filter_data_23__3 ;
    input filter_data_23__2 ;
    input filter_data_23__1 ;
    input filter_data_23__0 ;
    input filter_data_24__15 ;
    input filter_data_24__14 ;
    input filter_data_24__13 ;
    input filter_data_24__12 ;
    input filter_data_24__11 ;
    input filter_data_24__10 ;
    input filter_data_24__9 ;
    input filter_data_24__8 ;
    input filter_data_24__7 ;
    input filter_data_24__6 ;
    input filter_data_24__5 ;
    input filter_data_24__4 ;
    input filter_data_24__3 ;
    input filter_data_24__2 ;
    input filter_data_24__1 ;
    input filter_data_24__0 ;
    output d_arr_0__31 ;
    output d_arr_0__30 ;
    output d_arr_0__29 ;
    output d_arr_0__28 ;
    output d_arr_0__27 ;
    output d_arr_0__26 ;
    output d_arr_0__25 ;
    output d_arr_0__24 ;
    output d_arr_0__23 ;
    output d_arr_0__22 ;
    output d_arr_0__21 ;
    output d_arr_0__20 ;
    output d_arr_0__19 ;
    output d_arr_0__18 ;
    output d_arr_0__17 ;
    output d_arr_0__16 ;
    output d_arr_0__15 ;
    output d_arr_0__14 ;
    output d_arr_0__13 ;
    output d_arr_0__12 ;
    output d_arr_0__11 ;
    output d_arr_0__10 ;
    output d_arr_0__9 ;
    output d_arr_0__8 ;
    output d_arr_0__7 ;
    output d_arr_0__6 ;
    output d_arr_0__5 ;
    output d_arr_0__4 ;
    output d_arr_0__3 ;
    output d_arr_0__2 ;
    output d_arr_0__1 ;
    output d_arr_0__0 ;
    output d_arr_1__31 ;
    output d_arr_1__30 ;
    output d_arr_1__29 ;
    output d_arr_1__28 ;
    output d_arr_1__27 ;
    output d_arr_1__26 ;
    output d_arr_1__25 ;
    output d_arr_1__24 ;
    output d_arr_1__23 ;
    output d_arr_1__22 ;
    output d_arr_1__21 ;
    output d_arr_1__20 ;
    output d_arr_1__19 ;
    output d_arr_1__18 ;
    output d_arr_1__17 ;
    output d_arr_1__16 ;
    output d_arr_1__15 ;
    output d_arr_1__14 ;
    output d_arr_1__13 ;
    output d_arr_1__12 ;
    output d_arr_1__11 ;
    output d_arr_1__10 ;
    output d_arr_1__9 ;
    output d_arr_1__8 ;
    output d_arr_1__7 ;
    output d_arr_1__6 ;
    output d_arr_1__5 ;
    output d_arr_1__4 ;
    output d_arr_1__3 ;
    output d_arr_1__2 ;
    output d_arr_1__1 ;
    output d_arr_1__0 ;
    output d_arr_2__31 ;
    output d_arr_2__30 ;
    output d_arr_2__29 ;
    output d_arr_2__28 ;
    output d_arr_2__27 ;
    output d_arr_2__26 ;
    output d_arr_2__25 ;
    output d_arr_2__24 ;
    output d_arr_2__23 ;
    output d_arr_2__22 ;
    output d_arr_2__21 ;
    output d_arr_2__20 ;
    output d_arr_2__19 ;
    output d_arr_2__18 ;
    output d_arr_2__17 ;
    output d_arr_2__16 ;
    output d_arr_2__15 ;
    output d_arr_2__14 ;
    output d_arr_2__13 ;
    output d_arr_2__12 ;
    output d_arr_2__11 ;
    output d_arr_2__10 ;
    output d_arr_2__9 ;
    output d_arr_2__8 ;
    output d_arr_2__7 ;
    output d_arr_2__6 ;
    output d_arr_2__5 ;
    output d_arr_2__4 ;
    output d_arr_2__3 ;
    output d_arr_2__2 ;
    output d_arr_2__1 ;
    output d_arr_2__0 ;
    output d_arr_3__31 ;
    output d_arr_3__30 ;
    output d_arr_3__29 ;
    output d_arr_3__28 ;
    output d_arr_3__27 ;
    output d_arr_3__26 ;
    output d_arr_3__25 ;
    output d_arr_3__24 ;
    output d_arr_3__23 ;
    output d_arr_3__22 ;
    output d_arr_3__21 ;
    output d_arr_3__20 ;
    output d_arr_3__19 ;
    output d_arr_3__18 ;
    output d_arr_3__17 ;
    output d_arr_3__16 ;
    output d_arr_3__15 ;
    output d_arr_3__14 ;
    output d_arr_3__13 ;
    output d_arr_3__12 ;
    output d_arr_3__11 ;
    output d_arr_3__10 ;
    output d_arr_3__9 ;
    output d_arr_3__8 ;
    output d_arr_3__7 ;
    output d_arr_3__6 ;
    output d_arr_3__5 ;
    output d_arr_3__4 ;
    output d_arr_3__3 ;
    output d_arr_3__2 ;
    output d_arr_3__1 ;
    output d_arr_3__0 ;
    output d_arr_4__31 ;
    output d_arr_4__30 ;
    output d_arr_4__29 ;
    output d_arr_4__28 ;
    output d_arr_4__27 ;
    output d_arr_4__26 ;
    output d_arr_4__25 ;
    output d_arr_4__24 ;
    output d_arr_4__23 ;
    output d_arr_4__22 ;
    output d_arr_4__21 ;
    output d_arr_4__20 ;
    output d_arr_4__19 ;
    output d_arr_4__18 ;
    output d_arr_4__17 ;
    output d_arr_4__16 ;
    output d_arr_4__15 ;
    output d_arr_4__14 ;
    output d_arr_4__13 ;
    output d_arr_4__12 ;
    output d_arr_4__11 ;
    output d_arr_4__10 ;
    output d_arr_4__9 ;
    output d_arr_4__8 ;
    output d_arr_4__7 ;
    output d_arr_4__6 ;
    output d_arr_4__5 ;
    output d_arr_4__4 ;
    output d_arr_4__3 ;
    output d_arr_4__2 ;
    output d_arr_4__1 ;
    output d_arr_4__0 ;
    output d_arr_5__31 ;
    output d_arr_5__30 ;
    output d_arr_5__29 ;
    output d_arr_5__28 ;
    output d_arr_5__27 ;
    output d_arr_5__26 ;
    output d_arr_5__25 ;
    output d_arr_5__24 ;
    output d_arr_5__23 ;
    output d_arr_5__22 ;
    output d_arr_5__21 ;
    output d_arr_5__20 ;
    output d_arr_5__19 ;
    output d_arr_5__18 ;
    output d_arr_5__17 ;
    output d_arr_5__16 ;
    output d_arr_5__15 ;
    output d_arr_5__14 ;
    output d_arr_5__13 ;
    output d_arr_5__12 ;
    output d_arr_5__11 ;
    output d_arr_5__10 ;
    output d_arr_5__9 ;
    output d_arr_5__8 ;
    output d_arr_5__7 ;
    output d_arr_5__6 ;
    output d_arr_5__5 ;
    output d_arr_5__4 ;
    output d_arr_5__3 ;
    output d_arr_5__2 ;
    output d_arr_5__1 ;
    output d_arr_5__0 ;
    output d_arr_6__31 ;
    output d_arr_6__30 ;
    output d_arr_6__29 ;
    output d_arr_6__28 ;
    output d_arr_6__27 ;
    output d_arr_6__26 ;
    output d_arr_6__25 ;
    output d_arr_6__24 ;
    output d_arr_6__23 ;
    output d_arr_6__22 ;
    output d_arr_6__21 ;
    output d_arr_6__20 ;
    output d_arr_6__19 ;
    output d_arr_6__18 ;
    output d_arr_6__17 ;
    output d_arr_6__16 ;
    output d_arr_6__15 ;
    output d_arr_6__14 ;
    output d_arr_6__13 ;
    output d_arr_6__12 ;
    output d_arr_6__11 ;
    output d_arr_6__10 ;
    output d_arr_6__9 ;
    output d_arr_6__8 ;
    output d_arr_6__7 ;
    output d_arr_6__6 ;
    output d_arr_6__5 ;
    output d_arr_6__4 ;
    output d_arr_6__3 ;
    output d_arr_6__2 ;
    output d_arr_6__1 ;
    output d_arr_6__0 ;
    output d_arr_7__31 ;
    output d_arr_7__30 ;
    output d_arr_7__29 ;
    output d_arr_7__28 ;
    output d_arr_7__27 ;
    output d_arr_7__26 ;
    output d_arr_7__25 ;
    output d_arr_7__24 ;
    output d_arr_7__23 ;
    output d_arr_7__22 ;
    output d_arr_7__21 ;
    output d_arr_7__20 ;
    output d_arr_7__19 ;
    output d_arr_7__18 ;
    output d_arr_7__17 ;
    output d_arr_7__16 ;
    output d_arr_7__15 ;
    output d_arr_7__14 ;
    output d_arr_7__13 ;
    output d_arr_7__12 ;
    output d_arr_7__11 ;
    output d_arr_7__10 ;
    output d_arr_7__9 ;
    output d_arr_7__8 ;
    output d_arr_7__7 ;
    output d_arr_7__6 ;
    output d_arr_7__5 ;
    output d_arr_7__4 ;
    output d_arr_7__3 ;
    output d_arr_7__2 ;
    output d_arr_7__1 ;
    output d_arr_7__0 ;
    output d_arr_8__31 ;
    output d_arr_8__30 ;
    output d_arr_8__29 ;
    output d_arr_8__28 ;
    output d_arr_8__27 ;
    output d_arr_8__26 ;
    output d_arr_8__25 ;
    output d_arr_8__24 ;
    output d_arr_8__23 ;
    output d_arr_8__22 ;
    output d_arr_8__21 ;
    output d_arr_8__20 ;
    output d_arr_8__19 ;
    output d_arr_8__18 ;
    output d_arr_8__17 ;
    output d_arr_8__16 ;
    output d_arr_8__15 ;
    output d_arr_8__14 ;
    output d_arr_8__13 ;
    output d_arr_8__12 ;
    output d_arr_8__11 ;
    output d_arr_8__10 ;
    output d_arr_8__9 ;
    output d_arr_8__8 ;
    output d_arr_8__7 ;
    output d_arr_8__6 ;
    output d_arr_8__5 ;
    output d_arr_8__4 ;
    output d_arr_8__3 ;
    output d_arr_8__2 ;
    output d_arr_8__1 ;
    output d_arr_8__0 ;
    output d_arr_9__31 ;
    output d_arr_9__30 ;
    output d_arr_9__29 ;
    output d_arr_9__28 ;
    output d_arr_9__27 ;
    output d_arr_9__26 ;
    output d_arr_9__25 ;
    output d_arr_9__24 ;
    output d_arr_9__23 ;
    output d_arr_9__22 ;
    output d_arr_9__21 ;
    output d_arr_9__20 ;
    output d_arr_9__19 ;
    output d_arr_9__18 ;
    output d_arr_9__17 ;
    output d_arr_9__16 ;
    output d_arr_9__15 ;
    output d_arr_9__14 ;
    output d_arr_9__13 ;
    output d_arr_9__12 ;
    output d_arr_9__11 ;
    output d_arr_9__10 ;
    output d_arr_9__9 ;
    output d_arr_9__8 ;
    output d_arr_9__7 ;
    output d_arr_9__6 ;
    output d_arr_9__5 ;
    output d_arr_9__4 ;
    output d_arr_9__3 ;
    output d_arr_9__2 ;
    output d_arr_9__1 ;
    output d_arr_9__0 ;
    output d_arr_10__31 ;
    output d_arr_10__30 ;
    output d_arr_10__29 ;
    output d_arr_10__28 ;
    output d_arr_10__27 ;
    output d_arr_10__26 ;
    output d_arr_10__25 ;
    output d_arr_10__24 ;
    output d_arr_10__23 ;
    output d_arr_10__22 ;
    output d_arr_10__21 ;
    output d_arr_10__20 ;
    output d_arr_10__19 ;
    output d_arr_10__18 ;
    output d_arr_10__17 ;
    output d_arr_10__16 ;
    output d_arr_10__15 ;
    output d_arr_10__14 ;
    output d_arr_10__13 ;
    output d_arr_10__12 ;
    output d_arr_10__11 ;
    output d_arr_10__10 ;
    output d_arr_10__9 ;
    output d_arr_10__8 ;
    output d_arr_10__7 ;
    output d_arr_10__6 ;
    output d_arr_10__5 ;
    output d_arr_10__4 ;
    output d_arr_10__3 ;
    output d_arr_10__2 ;
    output d_arr_10__1 ;
    output d_arr_10__0 ;
    output d_arr_11__31 ;
    output d_arr_11__30 ;
    output d_arr_11__29 ;
    output d_arr_11__28 ;
    output d_arr_11__27 ;
    output d_arr_11__26 ;
    output d_arr_11__25 ;
    output d_arr_11__24 ;
    output d_arr_11__23 ;
    output d_arr_11__22 ;
    output d_arr_11__21 ;
    output d_arr_11__20 ;
    output d_arr_11__19 ;
    output d_arr_11__18 ;
    output d_arr_11__17 ;
    output d_arr_11__16 ;
    output d_arr_11__15 ;
    output d_arr_11__14 ;
    output d_arr_11__13 ;
    output d_arr_11__12 ;
    output d_arr_11__11 ;
    output d_arr_11__10 ;
    output d_arr_11__9 ;
    output d_arr_11__8 ;
    output d_arr_11__7 ;
    output d_arr_11__6 ;
    output d_arr_11__5 ;
    output d_arr_11__4 ;
    output d_arr_11__3 ;
    output d_arr_11__2 ;
    output d_arr_11__1 ;
    output d_arr_11__0 ;
    output d_arr_12__31 ;
    output d_arr_12__30 ;
    output d_arr_12__29 ;
    output d_arr_12__28 ;
    output d_arr_12__27 ;
    output d_arr_12__26 ;
    output d_arr_12__25 ;
    output d_arr_12__24 ;
    output d_arr_12__23 ;
    output d_arr_12__22 ;
    output d_arr_12__21 ;
    output d_arr_12__20 ;
    output d_arr_12__19 ;
    output d_arr_12__18 ;
    output d_arr_12__17 ;
    output d_arr_12__16 ;
    output d_arr_12__15 ;
    output d_arr_12__14 ;
    output d_arr_12__13 ;
    output d_arr_12__12 ;
    output d_arr_12__11 ;
    output d_arr_12__10 ;
    output d_arr_12__9 ;
    output d_arr_12__8 ;
    output d_arr_12__7 ;
    output d_arr_12__6 ;
    output d_arr_12__5 ;
    output d_arr_12__4 ;
    output d_arr_12__3 ;
    output d_arr_12__2 ;
    output d_arr_12__1 ;
    output d_arr_12__0 ;
    output d_arr_13__31 ;
    output d_arr_13__30 ;
    output d_arr_13__29 ;
    output d_arr_13__28 ;
    output d_arr_13__27 ;
    output d_arr_13__26 ;
    output d_arr_13__25 ;
    output d_arr_13__24 ;
    output d_arr_13__23 ;
    output d_arr_13__22 ;
    output d_arr_13__21 ;
    output d_arr_13__20 ;
    output d_arr_13__19 ;
    output d_arr_13__18 ;
    output d_arr_13__17 ;
    output d_arr_13__16 ;
    output d_arr_13__15 ;
    output d_arr_13__14 ;
    output d_arr_13__13 ;
    output d_arr_13__12 ;
    output d_arr_13__11 ;
    output d_arr_13__10 ;
    output d_arr_13__9 ;
    output d_arr_13__8 ;
    output d_arr_13__7 ;
    output d_arr_13__6 ;
    output d_arr_13__5 ;
    output d_arr_13__4 ;
    output d_arr_13__3 ;
    output d_arr_13__2 ;
    output d_arr_13__1 ;
    output d_arr_13__0 ;
    output d_arr_14__31 ;
    output d_arr_14__30 ;
    output d_arr_14__29 ;
    output d_arr_14__28 ;
    output d_arr_14__27 ;
    output d_arr_14__26 ;
    output d_arr_14__25 ;
    output d_arr_14__24 ;
    output d_arr_14__23 ;
    output d_arr_14__22 ;
    output d_arr_14__21 ;
    output d_arr_14__20 ;
    output d_arr_14__19 ;
    output d_arr_14__18 ;
    output d_arr_14__17 ;
    output d_arr_14__16 ;
    output d_arr_14__15 ;
    output d_arr_14__14 ;
    output d_arr_14__13 ;
    output d_arr_14__12 ;
    output d_arr_14__11 ;
    output d_arr_14__10 ;
    output d_arr_14__9 ;
    output d_arr_14__8 ;
    output d_arr_14__7 ;
    output d_arr_14__6 ;
    output d_arr_14__5 ;
    output d_arr_14__4 ;
    output d_arr_14__3 ;
    output d_arr_14__2 ;
    output d_arr_14__1 ;
    output d_arr_14__0 ;
    output d_arr_15__31 ;
    output d_arr_15__30 ;
    output d_arr_15__29 ;
    output d_arr_15__28 ;
    output d_arr_15__27 ;
    output d_arr_15__26 ;
    output d_arr_15__25 ;
    output d_arr_15__24 ;
    output d_arr_15__23 ;
    output d_arr_15__22 ;
    output d_arr_15__21 ;
    output d_arr_15__20 ;
    output d_arr_15__19 ;
    output d_arr_15__18 ;
    output d_arr_15__17 ;
    output d_arr_15__16 ;
    output d_arr_15__15 ;
    output d_arr_15__14 ;
    output d_arr_15__13 ;
    output d_arr_15__12 ;
    output d_arr_15__11 ;
    output d_arr_15__10 ;
    output d_arr_15__9 ;
    output d_arr_15__8 ;
    output d_arr_15__7 ;
    output d_arr_15__6 ;
    output d_arr_15__5 ;
    output d_arr_15__4 ;
    output d_arr_15__3 ;
    output d_arr_15__2 ;
    output d_arr_15__1 ;
    output d_arr_15__0 ;
    output d_arr_16__31 ;
    output d_arr_16__30 ;
    output d_arr_16__29 ;
    output d_arr_16__28 ;
    output d_arr_16__27 ;
    output d_arr_16__26 ;
    output d_arr_16__25 ;
    output d_arr_16__24 ;
    output d_arr_16__23 ;
    output d_arr_16__22 ;
    output d_arr_16__21 ;
    output d_arr_16__20 ;
    output d_arr_16__19 ;
    output d_arr_16__18 ;
    output d_arr_16__17 ;
    output d_arr_16__16 ;
    output d_arr_16__15 ;
    output d_arr_16__14 ;
    output d_arr_16__13 ;
    output d_arr_16__12 ;
    output d_arr_16__11 ;
    output d_arr_16__10 ;
    output d_arr_16__9 ;
    output d_arr_16__8 ;
    output d_arr_16__7 ;
    output d_arr_16__6 ;
    output d_arr_16__5 ;
    output d_arr_16__4 ;
    output d_arr_16__3 ;
    output d_arr_16__2 ;
    output d_arr_16__1 ;
    output d_arr_16__0 ;
    output d_arr_17__31 ;
    output d_arr_17__30 ;
    output d_arr_17__29 ;
    output d_arr_17__28 ;
    output d_arr_17__27 ;
    output d_arr_17__26 ;
    output d_arr_17__25 ;
    output d_arr_17__24 ;
    output d_arr_17__23 ;
    output d_arr_17__22 ;
    output d_arr_17__21 ;
    output d_arr_17__20 ;
    output d_arr_17__19 ;
    output d_arr_17__18 ;
    output d_arr_17__17 ;
    output d_arr_17__16 ;
    output d_arr_17__15 ;
    output d_arr_17__14 ;
    output d_arr_17__13 ;
    output d_arr_17__12 ;
    output d_arr_17__11 ;
    output d_arr_17__10 ;
    output d_arr_17__9 ;
    output d_arr_17__8 ;
    output d_arr_17__7 ;
    output d_arr_17__6 ;
    output d_arr_17__5 ;
    output d_arr_17__4 ;
    output d_arr_17__3 ;
    output d_arr_17__2 ;
    output d_arr_17__1 ;
    output d_arr_17__0 ;
    output d_arr_18__31 ;
    output d_arr_18__30 ;
    output d_arr_18__29 ;
    output d_arr_18__28 ;
    output d_arr_18__27 ;
    output d_arr_18__26 ;
    output d_arr_18__25 ;
    output d_arr_18__24 ;
    output d_arr_18__23 ;
    output d_arr_18__22 ;
    output d_arr_18__21 ;
    output d_arr_18__20 ;
    output d_arr_18__19 ;
    output d_arr_18__18 ;
    output d_arr_18__17 ;
    output d_arr_18__16 ;
    output d_arr_18__15 ;
    output d_arr_18__14 ;
    output d_arr_18__13 ;
    output d_arr_18__12 ;
    output d_arr_18__11 ;
    output d_arr_18__10 ;
    output d_arr_18__9 ;
    output d_arr_18__8 ;
    output d_arr_18__7 ;
    output d_arr_18__6 ;
    output d_arr_18__5 ;
    output d_arr_18__4 ;
    output d_arr_18__3 ;
    output d_arr_18__2 ;
    output d_arr_18__1 ;
    output d_arr_18__0 ;
    output d_arr_19__31 ;
    output d_arr_19__30 ;
    output d_arr_19__29 ;
    output d_arr_19__28 ;
    output d_arr_19__27 ;
    output d_arr_19__26 ;
    output d_arr_19__25 ;
    output d_arr_19__24 ;
    output d_arr_19__23 ;
    output d_arr_19__22 ;
    output d_arr_19__21 ;
    output d_arr_19__20 ;
    output d_arr_19__19 ;
    output d_arr_19__18 ;
    output d_arr_19__17 ;
    output d_arr_19__16 ;
    output d_arr_19__15 ;
    output d_arr_19__14 ;
    output d_arr_19__13 ;
    output d_arr_19__12 ;
    output d_arr_19__11 ;
    output d_arr_19__10 ;
    output d_arr_19__9 ;
    output d_arr_19__8 ;
    output d_arr_19__7 ;
    output d_arr_19__6 ;
    output d_arr_19__5 ;
    output d_arr_19__4 ;
    output d_arr_19__3 ;
    output d_arr_19__2 ;
    output d_arr_19__1 ;
    output d_arr_19__0 ;
    output d_arr_20__31 ;
    output d_arr_20__30 ;
    output d_arr_20__29 ;
    output d_arr_20__28 ;
    output d_arr_20__27 ;
    output d_arr_20__26 ;
    output d_arr_20__25 ;
    output d_arr_20__24 ;
    output d_arr_20__23 ;
    output d_arr_20__22 ;
    output d_arr_20__21 ;
    output d_arr_20__20 ;
    output d_arr_20__19 ;
    output d_arr_20__18 ;
    output d_arr_20__17 ;
    output d_arr_20__16 ;
    output d_arr_20__15 ;
    output d_arr_20__14 ;
    output d_arr_20__13 ;
    output d_arr_20__12 ;
    output d_arr_20__11 ;
    output d_arr_20__10 ;
    output d_arr_20__9 ;
    output d_arr_20__8 ;
    output d_arr_20__7 ;
    output d_arr_20__6 ;
    output d_arr_20__5 ;
    output d_arr_20__4 ;
    output d_arr_20__3 ;
    output d_arr_20__2 ;
    output d_arr_20__1 ;
    output d_arr_20__0 ;
    output d_arr_21__31 ;
    output d_arr_21__30 ;
    output d_arr_21__29 ;
    output d_arr_21__28 ;
    output d_arr_21__27 ;
    output d_arr_21__26 ;
    output d_arr_21__25 ;
    output d_arr_21__24 ;
    output d_arr_21__23 ;
    output d_arr_21__22 ;
    output d_arr_21__21 ;
    output d_arr_21__20 ;
    output d_arr_21__19 ;
    output d_arr_21__18 ;
    output d_arr_21__17 ;
    output d_arr_21__16 ;
    output d_arr_21__15 ;
    output d_arr_21__14 ;
    output d_arr_21__13 ;
    output d_arr_21__12 ;
    output d_arr_21__11 ;
    output d_arr_21__10 ;
    output d_arr_21__9 ;
    output d_arr_21__8 ;
    output d_arr_21__7 ;
    output d_arr_21__6 ;
    output d_arr_21__5 ;
    output d_arr_21__4 ;
    output d_arr_21__3 ;
    output d_arr_21__2 ;
    output d_arr_21__1 ;
    output d_arr_21__0 ;
    output d_arr_22__31 ;
    output d_arr_22__30 ;
    output d_arr_22__29 ;
    output d_arr_22__28 ;
    output d_arr_22__27 ;
    output d_arr_22__26 ;
    output d_arr_22__25 ;
    output d_arr_22__24 ;
    output d_arr_22__23 ;
    output d_arr_22__22 ;
    output d_arr_22__21 ;
    output d_arr_22__20 ;
    output d_arr_22__19 ;
    output d_arr_22__18 ;
    output d_arr_22__17 ;
    output d_arr_22__16 ;
    output d_arr_22__15 ;
    output d_arr_22__14 ;
    output d_arr_22__13 ;
    output d_arr_22__12 ;
    output d_arr_22__11 ;
    output d_arr_22__10 ;
    output d_arr_22__9 ;
    output d_arr_22__8 ;
    output d_arr_22__7 ;
    output d_arr_22__6 ;
    output d_arr_22__5 ;
    output d_arr_22__4 ;
    output d_arr_22__3 ;
    output d_arr_22__2 ;
    output d_arr_22__1 ;
    output d_arr_22__0 ;
    output d_arr_23__31 ;
    output d_arr_23__30 ;
    output d_arr_23__29 ;
    output d_arr_23__28 ;
    output d_arr_23__27 ;
    output d_arr_23__26 ;
    output d_arr_23__25 ;
    output d_arr_23__24 ;
    output d_arr_23__23 ;
    output d_arr_23__22 ;
    output d_arr_23__21 ;
    output d_arr_23__20 ;
    output d_arr_23__19 ;
    output d_arr_23__18 ;
    output d_arr_23__17 ;
    output d_arr_23__16 ;
    output d_arr_23__15 ;
    output d_arr_23__14 ;
    output d_arr_23__13 ;
    output d_arr_23__12 ;
    output d_arr_23__11 ;
    output d_arr_23__10 ;
    output d_arr_23__9 ;
    output d_arr_23__8 ;
    output d_arr_23__7 ;
    output d_arr_23__6 ;
    output d_arr_23__5 ;
    output d_arr_23__4 ;
    output d_arr_23__3 ;
    output d_arr_23__2 ;
    output d_arr_23__1 ;
    output d_arr_23__0 ;
    output d_arr_24__31 ;
    output d_arr_24__30 ;
    output d_arr_24__29 ;
    output d_arr_24__28 ;
    output d_arr_24__27 ;
    output d_arr_24__26 ;
    output d_arr_24__25 ;
    output d_arr_24__24 ;
    output d_arr_24__23 ;
    output d_arr_24__22 ;
    output d_arr_24__21 ;
    output d_arr_24__20 ;
    output d_arr_24__19 ;
    output d_arr_24__18 ;
    output d_arr_24__17 ;
    output d_arr_24__16 ;
    output d_arr_24__15 ;
    output d_arr_24__14 ;
    output d_arr_24__13 ;
    output d_arr_24__12 ;
    output d_arr_24__11 ;
    output d_arr_24__10 ;
    output d_arr_24__9 ;
    output d_arr_24__8 ;
    output d_arr_24__7 ;
    output d_arr_24__6 ;
    output d_arr_24__5 ;
    output d_arr_24__4 ;
    output d_arr_24__3 ;
    output d_arr_24__2 ;
    output d_arr_24__1 ;
    output d_arr_24__0 ;
    input q_arr_0__31 ;
    input q_arr_0__30 ;
    input q_arr_0__29 ;
    input q_arr_0__28 ;
    input q_arr_0__27 ;
    input q_arr_0__26 ;
    input q_arr_0__25 ;
    input q_arr_0__24 ;
    input q_arr_0__23 ;
    input q_arr_0__22 ;
    input q_arr_0__21 ;
    input q_arr_0__20 ;
    input q_arr_0__19 ;
    input q_arr_0__18 ;
    input q_arr_0__17 ;
    input q_arr_0__16 ;
    input q_arr_0__15 ;
    input q_arr_0__14 ;
    input q_arr_0__13 ;
    input q_arr_0__12 ;
    input q_arr_0__11 ;
    input q_arr_0__10 ;
    input q_arr_0__9 ;
    input q_arr_0__8 ;
    input q_arr_0__7 ;
    input q_arr_0__6 ;
    input q_arr_0__5 ;
    input q_arr_0__4 ;
    input q_arr_0__3 ;
    input q_arr_0__2 ;
    input q_arr_0__1 ;
    input q_arr_0__0 ;
    input q_arr_1__31 ;
    input q_arr_1__30 ;
    input q_arr_1__29 ;
    input q_arr_1__28 ;
    input q_arr_1__27 ;
    input q_arr_1__26 ;
    input q_arr_1__25 ;
    input q_arr_1__24 ;
    input q_arr_1__23 ;
    input q_arr_1__22 ;
    input q_arr_1__21 ;
    input q_arr_1__20 ;
    input q_arr_1__19 ;
    input q_arr_1__18 ;
    input q_arr_1__17 ;
    input q_arr_1__16 ;
    input q_arr_1__15 ;
    input q_arr_1__14 ;
    input q_arr_1__13 ;
    input q_arr_1__12 ;
    input q_arr_1__11 ;
    input q_arr_1__10 ;
    input q_arr_1__9 ;
    input q_arr_1__8 ;
    input q_arr_1__7 ;
    input q_arr_1__6 ;
    input q_arr_1__5 ;
    input q_arr_1__4 ;
    input q_arr_1__3 ;
    input q_arr_1__2 ;
    input q_arr_1__1 ;
    input q_arr_1__0 ;
    input q_arr_2__31 ;
    input q_arr_2__30 ;
    input q_arr_2__29 ;
    input q_arr_2__28 ;
    input q_arr_2__27 ;
    input q_arr_2__26 ;
    input q_arr_2__25 ;
    input q_arr_2__24 ;
    input q_arr_2__23 ;
    input q_arr_2__22 ;
    input q_arr_2__21 ;
    input q_arr_2__20 ;
    input q_arr_2__19 ;
    input q_arr_2__18 ;
    input q_arr_2__17 ;
    input q_arr_2__16 ;
    input q_arr_2__15 ;
    input q_arr_2__14 ;
    input q_arr_2__13 ;
    input q_arr_2__12 ;
    input q_arr_2__11 ;
    input q_arr_2__10 ;
    input q_arr_2__9 ;
    input q_arr_2__8 ;
    input q_arr_2__7 ;
    input q_arr_2__6 ;
    input q_arr_2__5 ;
    input q_arr_2__4 ;
    input q_arr_2__3 ;
    input q_arr_2__2 ;
    input q_arr_2__1 ;
    input q_arr_2__0 ;
    input q_arr_3__31 ;
    input q_arr_3__30 ;
    input q_arr_3__29 ;
    input q_arr_3__28 ;
    input q_arr_3__27 ;
    input q_arr_3__26 ;
    input q_arr_3__25 ;
    input q_arr_3__24 ;
    input q_arr_3__23 ;
    input q_arr_3__22 ;
    input q_arr_3__21 ;
    input q_arr_3__20 ;
    input q_arr_3__19 ;
    input q_arr_3__18 ;
    input q_arr_3__17 ;
    input q_arr_3__16 ;
    input q_arr_3__15 ;
    input q_arr_3__14 ;
    input q_arr_3__13 ;
    input q_arr_3__12 ;
    input q_arr_3__11 ;
    input q_arr_3__10 ;
    input q_arr_3__9 ;
    input q_arr_3__8 ;
    input q_arr_3__7 ;
    input q_arr_3__6 ;
    input q_arr_3__5 ;
    input q_arr_3__4 ;
    input q_arr_3__3 ;
    input q_arr_3__2 ;
    input q_arr_3__1 ;
    input q_arr_3__0 ;
    input q_arr_4__31 ;
    input q_arr_4__30 ;
    input q_arr_4__29 ;
    input q_arr_4__28 ;
    input q_arr_4__27 ;
    input q_arr_4__26 ;
    input q_arr_4__25 ;
    input q_arr_4__24 ;
    input q_arr_4__23 ;
    input q_arr_4__22 ;
    input q_arr_4__21 ;
    input q_arr_4__20 ;
    input q_arr_4__19 ;
    input q_arr_4__18 ;
    input q_arr_4__17 ;
    input q_arr_4__16 ;
    input q_arr_4__15 ;
    input q_arr_4__14 ;
    input q_arr_4__13 ;
    input q_arr_4__12 ;
    input q_arr_4__11 ;
    input q_arr_4__10 ;
    input q_arr_4__9 ;
    input q_arr_4__8 ;
    input q_arr_4__7 ;
    input q_arr_4__6 ;
    input q_arr_4__5 ;
    input q_arr_4__4 ;
    input q_arr_4__3 ;
    input q_arr_4__2 ;
    input q_arr_4__1 ;
    input q_arr_4__0 ;
    input q_arr_5__31 ;
    input q_arr_5__30 ;
    input q_arr_5__29 ;
    input q_arr_5__28 ;
    input q_arr_5__27 ;
    input q_arr_5__26 ;
    input q_arr_5__25 ;
    input q_arr_5__24 ;
    input q_arr_5__23 ;
    input q_arr_5__22 ;
    input q_arr_5__21 ;
    input q_arr_5__20 ;
    input q_arr_5__19 ;
    input q_arr_5__18 ;
    input q_arr_5__17 ;
    input q_arr_5__16 ;
    input q_arr_5__15 ;
    input q_arr_5__14 ;
    input q_arr_5__13 ;
    input q_arr_5__12 ;
    input q_arr_5__11 ;
    input q_arr_5__10 ;
    input q_arr_5__9 ;
    input q_arr_5__8 ;
    input q_arr_5__7 ;
    input q_arr_5__6 ;
    input q_arr_5__5 ;
    input q_arr_5__4 ;
    input q_arr_5__3 ;
    input q_arr_5__2 ;
    input q_arr_5__1 ;
    input q_arr_5__0 ;
    input q_arr_6__31 ;
    input q_arr_6__30 ;
    input q_arr_6__29 ;
    input q_arr_6__28 ;
    input q_arr_6__27 ;
    input q_arr_6__26 ;
    input q_arr_6__25 ;
    input q_arr_6__24 ;
    input q_arr_6__23 ;
    input q_arr_6__22 ;
    input q_arr_6__21 ;
    input q_arr_6__20 ;
    input q_arr_6__19 ;
    input q_arr_6__18 ;
    input q_arr_6__17 ;
    input q_arr_6__16 ;
    input q_arr_6__15 ;
    input q_arr_6__14 ;
    input q_arr_6__13 ;
    input q_arr_6__12 ;
    input q_arr_6__11 ;
    input q_arr_6__10 ;
    input q_arr_6__9 ;
    input q_arr_6__8 ;
    input q_arr_6__7 ;
    input q_arr_6__6 ;
    input q_arr_6__5 ;
    input q_arr_6__4 ;
    input q_arr_6__3 ;
    input q_arr_6__2 ;
    input q_arr_6__1 ;
    input q_arr_6__0 ;
    input q_arr_7__31 ;
    input q_arr_7__30 ;
    input q_arr_7__29 ;
    input q_arr_7__28 ;
    input q_arr_7__27 ;
    input q_arr_7__26 ;
    input q_arr_7__25 ;
    input q_arr_7__24 ;
    input q_arr_7__23 ;
    input q_arr_7__22 ;
    input q_arr_7__21 ;
    input q_arr_7__20 ;
    input q_arr_7__19 ;
    input q_arr_7__18 ;
    input q_arr_7__17 ;
    input q_arr_7__16 ;
    input q_arr_7__15 ;
    input q_arr_7__14 ;
    input q_arr_7__13 ;
    input q_arr_7__12 ;
    input q_arr_7__11 ;
    input q_arr_7__10 ;
    input q_arr_7__9 ;
    input q_arr_7__8 ;
    input q_arr_7__7 ;
    input q_arr_7__6 ;
    input q_arr_7__5 ;
    input q_arr_7__4 ;
    input q_arr_7__3 ;
    input q_arr_7__2 ;
    input q_arr_7__1 ;
    input q_arr_7__0 ;
    input q_arr_8__31 ;
    input q_arr_8__30 ;
    input q_arr_8__29 ;
    input q_arr_8__28 ;
    input q_arr_8__27 ;
    input q_arr_8__26 ;
    input q_arr_8__25 ;
    input q_arr_8__24 ;
    input q_arr_8__23 ;
    input q_arr_8__22 ;
    input q_arr_8__21 ;
    input q_arr_8__20 ;
    input q_arr_8__19 ;
    input q_arr_8__18 ;
    input q_arr_8__17 ;
    input q_arr_8__16 ;
    input q_arr_8__15 ;
    input q_arr_8__14 ;
    input q_arr_8__13 ;
    input q_arr_8__12 ;
    input q_arr_8__11 ;
    input q_arr_8__10 ;
    input q_arr_8__9 ;
    input q_arr_8__8 ;
    input q_arr_8__7 ;
    input q_arr_8__6 ;
    input q_arr_8__5 ;
    input q_arr_8__4 ;
    input q_arr_8__3 ;
    input q_arr_8__2 ;
    input q_arr_8__1 ;
    input q_arr_8__0 ;
    input q_arr_9__31 ;
    input q_arr_9__30 ;
    input q_arr_9__29 ;
    input q_arr_9__28 ;
    input q_arr_9__27 ;
    input q_arr_9__26 ;
    input q_arr_9__25 ;
    input q_arr_9__24 ;
    input q_arr_9__23 ;
    input q_arr_9__22 ;
    input q_arr_9__21 ;
    input q_arr_9__20 ;
    input q_arr_9__19 ;
    input q_arr_9__18 ;
    input q_arr_9__17 ;
    input q_arr_9__16 ;
    input q_arr_9__15 ;
    input q_arr_9__14 ;
    input q_arr_9__13 ;
    input q_arr_9__12 ;
    input q_arr_9__11 ;
    input q_arr_9__10 ;
    input q_arr_9__9 ;
    input q_arr_9__8 ;
    input q_arr_9__7 ;
    input q_arr_9__6 ;
    input q_arr_9__5 ;
    input q_arr_9__4 ;
    input q_arr_9__3 ;
    input q_arr_9__2 ;
    input q_arr_9__1 ;
    input q_arr_9__0 ;
    input q_arr_10__31 ;
    input q_arr_10__30 ;
    input q_arr_10__29 ;
    input q_arr_10__28 ;
    input q_arr_10__27 ;
    input q_arr_10__26 ;
    input q_arr_10__25 ;
    input q_arr_10__24 ;
    input q_arr_10__23 ;
    input q_arr_10__22 ;
    input q_arr_10__21 ;
    input q_arr_10__20 ;
    input q_arr_10__19 ;
    input q_arr_10__18 ;
    input q_arr_10__17 ;
    input q_arr_10__16 ;
    input q_arr_10__15 ;
    input q_arr_10__14 ;
    input q_arr_10__13 ;
    input q_arr_10__12 ;
    input q_arr_10__11 ;
    input q_arr_10__10 ;
    input q_arr_10__9 ;
    input q_arr_10__8 ;
    input q_arr_10__7 ;
    input q_arr_10__6 ;
    input q_arr_10__5 ;
    input q_arr_10__4 ;
    input q_arr_10__3 ;
    input q_arr_10__2 ;
    input q_arr_10__1 ;
    input q_arr_10__0 ;
    input q_arr_11__31 ;
    input q_arr_11__30 ;
    input q_arr_11__29 ;
    input q_arr_11__28 ;
    input q_arr_11__27 ;
    input q_arr_11__26 ;
    input q_arr_11__25 ;
    input q_arr_11__24 ;
    input q_arr_11__23 ;
    input q_arr_11__22 ;
    input q_arr_11__21 ;
    input q_arr_11__20 ;
    input q_arr_11__19 ;
    input q_arr_11__18 ;
    input q_arr_11__17 ;
    input q_arr_11__16 ;
    input q_arr_11__15 ;
    input q_arr_11__14 ;
    input q_arr_11__13 ;
    input q_arr_11__12 ;
    input q_arr_11__11 ;
    input q_arr_11__10 ;
    input q_arr_11__9 ;
    input q_arr_11__8 ;
    input q_arr_11__7 ;
    input q_arr_11__6 ;
    input q_arr_11__5 ;
    input q_arr_11__4 ;
    input q_arr_11__3 ;
    input q_arr_11__2 ;
    input q_arr_11__1 ;
    input q_arr_11__0 ;
    input q_arr_12__31 ;
    input q_arr_12__30 ;
    input q_arr_12__29 ;
    input q_arr_12__28 ;
    input q_arr_12__27 ;
    input q_arr_12__26 ;
    input q_arr_12__25 ;
    input q_arr_12__24 ;
    input q_arr_12__23 ;
    input q_arr_12__22 ;
    input q_arr_12__21 ;
    input q_arr_12__20 ;
    input q_arr_12__19 ;
    input q_arr_12__18 ;
    input q_arr_12__17 ;
    input q_arr_12__16 ;
    input q_arr_12__15 ;
    input q_arr_12__14 ;
    input q_arr_12__13 ;
    input q_arr_12__12 ;
    input q_arr_12__11 ;
    input q_arr_12__10 ;
    input q_arr_12__9 ;
    input q_arr_12__8 ;
    input q_arr_12__7 ;
    input q_arr_12__6 ;
    input q_arr_12__5 ;
    input q_arr_12__4 ;
    input q_arr_12__3 ;
    input q_arr_12__2 ;
    input q_arr_12__1 ;
    input q_arr_12__0 ;
    input q_arr_13__31 ;
    input q_arr_13__30 ;
    input q_arr_13__29 ;
    input q_arr_13__28 ;
    input q_arr_13__27 ;
    input q_arr_13__26 ;
    input q_arr_13__25 ;
    input q_arr_13__24 ;
    input q_arr_13__23 ;
    input q_arr_13__22 ;
    input q_arr_13__21 ;
    input q_arr_13__20 ;
    input q_arr_13__19 ;
    input q_arr_13__18 ;
    input q_arr_13__17 ;
    input q_arr_13__16 ;
    input q_arr_13__15 ;
    input q_arr_13__14 ;
    input q_arr_13__13 ;
    input q_arr_13__12 ;
    input q_arr_13__11 ;
    input q_arr_13__10 ;
    input q_arr_13__9 ;
    input q_arr_13__8 ;
    input q_arr_13__7 ;
    input q_arr_13__6 ;
    input q_arr_13__5 ;
    input q_arr_13__4 ;
    input q_arr_13__3 ;
    input q_arr_13__2 ;
    input q_arr_13__1 ;
    input q_arr_13__0 ;
    input q_arr_14__31 ;
    input q_arr_14__30 ;
    input q_arr_14__29 ;
    input q_arr_14__28 ;
    input q_arr_14__27 ;
    input q_arr_14__26 ;
    input q_arr_14__25 ;
    input q_arr_14__24 ;
    input q_arr_14__23 ;
    input q_arr_14__22 ;
    input q_arr_14__21 ;
    input q_arr_14__20 ;
    input q_arr_14__19 ;
    input q_arr_14__18 ;
    input q_arr_14__17 ;
    input q_arr_14__16 ;
    input q_arr_14__15 ;
    input q_arr_14__14 ;
    input q_arr_14__13 ;
    input q_arr_14__12 ;
    input q_arr_14__11 ;
    input q_arr_14__10 ;
    input q_arr_14__9 ;
    input q_arr_14__8 ;
    input q_arr_14__7 ;
    input q_arr_14__6 ;
    input q_arr_14__5 ;
    input q_arr_14__4 ;
    input q_arr_14__3 ;
    input q_arr_14__2 ;
    input q_arr_14__1 ;
    input q_arr_14__0 ;
    input q_arr_15__31 ;
    input q_arr_15__30 ;
    input q_arr_15__29 ;
    input q_arr_15__28 ;
    input q_arr_15__27 ;
    input q_arr_15__26 ;
    input q_arr_15__25 ;
    input q_arr_15__24 ;
    input q_arr_15__23 ;
    input q_arr_15__22 ;
    input q_arr_15__21 ;
    input q_arr_15__20 ;
    input q_arr_15__19 ;
    input q_arr_15__18 ;
    input q_arr_15__17 ;
    input q_arr_15__16 ;
    input q_arr_15__15 ;
    input q_arr_15__14 ;
    input q_arr_15__13 ;
    input q_arr_15__12 ;
    input q_arr_15__11 ;
    input q_arr_15__10 ;
    input q_arr_15__9 ;
    input q_arr_15__8 ;
    input q_arr_15__7 ;
    input q_arr_15__6 ;
    input q_arr_15__5 ;
    input q_arr_15__4 ;
    input q_arr_15__3 ;
    input q_arr_15__2 ;
    input q_arr_15__1 ;
    input q_arr_15__0 ;
    input q_arr_16__31 ;
    input q_arr_16__30 ;
    input q_arr_16__29 ;
    input q_arr_16__28 ;
    input q_arr_16__27 ;
    input q_arr_16__26 ;
    input q_arr_16__25 ;
    input q_arr_16__24 ;
    input q_arr_16__23 ;
    input q_arr_16__22 ;
    input q_arr_16__21 ;
    input q_arr_16__20 ;
    input q_arr_16__19 ;
    input q_arr_16__18 ;
    input q_arr_16__17 ;
    input q_arr_16__16 ;
    input q_arr_16__15 ;
    input q_arr_16__14 ;
    input q_arr_16__13 ;
    input q_arr_16__12 ;
    input q_arr_16__11 ;
    input q_arr_16__10 ;
    input q_arr_16__9 ;
    input q_arr_16__8 ;
    input q_arr_16__7 ;
    input q_arr_16__6 ;
    input q_arr_16__5 ;
    input q_arr_16__4 ;
    input q_arr_16__3 ;
    input q_arr_16__2 ;
    input q_arr_16__1 ;
    input q_arr_16__0 ;
    input q_arr_17__31 ;
    input q_arr_17__30 ;
    input q_arr_17__29 ;
    input q_arr_17__28 ;
    input q_arr_17__27 ;
    input q_arr_17__26 ;
    input q_arr_17__25 ;
    input q_arr_17__24 ;
    input q_arr_17__23 ;
    input q_arr_17__22 ;
    input q_arr_17__21 ;
    input q_arr_17__20 ;
    input q_arr_17__19 ;
    input q_arr_17__18 ;
    input q_arr_17__17 ;
    input q_arr_17__16 ;
    input q_arr_17__15 ;
    input q_arr_17__14 ;
    input q_arr_17__13 ;
    input q_arr_17__12 ;
    input q_arr_17__11 ;
    input q_arr_17__10 ;
    input q_arr_17__9 ;
    input q_arr_17__8 ;
    input q_arr_17__7 ;
    input q_arr_17__6 ;
    input q_arr_17__5 ;
    input q_arr_17__4 ;
    input q_arr_17__3 ;
    input q_arr_17__2 ;
    input q_arr_17__1 ;
    input q_arr_17__0 ;
    input q_arr_18__31 ;
    input q_arr_18__30 ;
    input q_arr_18__29 ;
    input q_arr_18__28 ;
    input q_arr_18__27 ;
    input q_arr_18__26 ;
    input q_arr_18__25 ;
    input q_arr_18__24 ;
    input q_arr_18__23 ;
    input q_arr_18__22 ;
    input q_arr_18__21 ;
    input q_arr_18__20 ;
    input q_arr_18__19 ;
    input q_arr_18__18 ;
    input q_arr_18__17 ;
    input q_arr_18__16 ;
    input q_arr_18__15 ;
    input q_arr_18__14 ;
    input q_arr_18__13 ;
    input q_arr_18__12 ;
    input q_arr_18__11 ;
    input q_arr_18__10 ;
    input q_arr_18__9 ;
    input q_arr_18__8 ;
    input q_arr_18__7 ;
    input q_arr_18__6 ;
    input q_arr_18__5 ;
    input q_arr_18__4 ;
    input q_arr_18__3 ;
    input q_arr_18__2 ;
    input q_arr_18__1 ;
    input q_arr_18__0 ;
    input q_arr_19__31 ;
    input q_arr_19__30 ;
    input q_arr_19__29 ;
    input q_arr_19__28 ;
    input q_arr_19__27 ;
    input q_arr_19__26 ;
    input q_arr_19__25 ;
    input q_arr_19__24 ;
    input q_arr_19__23 ;
    input q_arr_19__22 ;
    input q_arr_19__21 ;
    input q_arr_19__20 ;
    input q_arr_19__19 ;
    input q_arr_19__18 ;
    input q_arr_19__17 ;
    input q_arr_19__16 ;
    input q_arr_19__15 ;
    input q_arr_19__14 ;
    input q_arr_19__13 ;
    input q_arr_19__12 ;
    input q_arr_19__11 ;
    input q_arr_19__10 ;
    input q_arr_19__9 ;
    input q_arr_19__8 ;
    input q_arr_19__7 ;
    input q_arr_19__6 ;
    input q_arr_19__5 ;
    input q_arr_19__4 ;
    input q_arr_19__3 ;
    input q_arr_19__2 ;
    input q_arr_19__1 ;
    input q_arr_19__0 ;
    input q_arr_20__31 ;
    input q_arr_20__30 ;
    input q_arr_20__29 ;
    input q_arr_20__28 ;
    input q_arr_20__27 ;
    input q_arr_20__26 ;
    input q_arr_20__25 ;
    input q_arr_20__24 ;
    input q_arr_20__23 ;
    input q_arr_20__22 ;
    input q_arr_20__21 ;
    input q_arr_20__20 ;
    input q_arr_20__19 ;
    input q_arr_20__18 ;
    input q_arr_20__17 ;
    input q_arr_20__16 ;
    input q_arr_20__15 ;
    input q_arr_20__14 ;
    input q_arr_20__13 ;
    input q_arr_20__12 ;
    input q_arr_20__11 ;
    input q_arr_20__10 ;
    input q_arr_20__9 ;
    input q_arr_20__8 ;
    input q_arr_20__7 ;
    input q_arr_20__6 ;
    input q_arr_20__5 ;
    input q_arr_20__4 ;
    input q_arr_20__3 ;
    input q_arr_20__2 ;
    input q_arr_20__1 ;
    input q_arr_20__0 ;
    input q_arr_21__31 ;
    input q_arr_21__30 ;
    input q_arr_21__29 ;
    input q_arr_21__28 ;
    input q_arr_21__27 ;
    input q_arr_21__26 ;
    input q_arr_21__25 ;
    input q_arr_21__24 ;
    input q_arr_21__23 ;
    input q_arr_21__22 ;
    input q_arr_21__21 ;
    input q_arr_21__20 ;
    input q_arr_21__19 ;
    input q_arr_21__18 ;
    input q_arr_21__17 ;
    input q_arr_21__16 ;
    input q_arr_21__15 ;
    input q_arr_21__14 ;
    input q_arr_21__13 ;
    input q_arr_21__12 ;
    input q_arr_21__11 ;
    input q_arr_21__10 ;
    input q_arr_21__9 ;
    input q_arr_21__8 ;
    input q_arr_21__7 ;
    input q_arr_21__6 ;
    input q_arr_21__5 ;
    input q_arr_21__4 ;
    input q_arr_21__3 ;
    input q_arr_21__2 ;
    input q_arr_21__1 ;
    input q_arr_21__0 ;
    input q_arr_22__31 ;
    input q_arr_22__30 ;
    input q_arr_22__29 ;
    input q_arr_22__28 ;
    input q_arr_22__27 ;
    input q_arr_22__26 ;
    input q_arr_22__25 ;
    input q_arr_22__24 ;
    input q_arr_22__23 ;
    input q_arr_22__22 ;
    input q_arr_22__21 ;
    input q_arr_22__20 ;
    input q_arr_22__19 ;
    input q_arr_22__18 ;
    input q_arr_22__17 ;
    input q_arr_22__16 ;
    input q_arr_22__15 ;
    input q_arr_22__14 ;
    input q_arr_22__13 ;
    input q_arr_22__12 ;
    input q_arr_22__11 ;
    input q_arr_22__10 ;
    input q_arr_22__9 ;
    input q_arr_22__8 ;
    input q_arr_22__7 ;
    input q_arr_22__6 ;
    input q_arr_22__5 ;
    input q_arr_22__4 ;
    input q_arr_22__3 ;
    input q_arr_22__2 ;
    input q_arr_22__1 ;
    input q_arr_22__0 ;
    input q_arr_23__31 ;
    input q_arr_23__30 ;
    input q_arr_23__29 ;
    input q_arr_23__28 ;
    input q_arr_23__27 ;
    input q_arr_23__26 ;
    input q_arr_23__25 ;
    input q_arr_23__24 ;
    input q_arr_23__23 ;
    input q_arr_23__22 ;
    input q_arr_23__21 ;
    input q_arr_23__20 ;
    input q_arr_23__19 ;
    input q_arr_23__18 ;
    input q_arr_23__17 ;
    input q_arr_23__16 ;
    input q_arr_23__15 ;
    input q_arr_23__14 ;
    input q_arr_23__13 ;
    input q_arr_23__12 ;
    input q_arr_23__11 ;
    input q_arr_23__10 ;
    input q_arr_23__9 ;
    input q_arr_23__8 ;
    input q_arr_23__7 ;
    input q_arr_23__6 ;
    input q_arr_23__5 ;
    input q_arr_23__4 ;
    input q_arr_23__3 ;
    input q_arr_23__2 ;
    input q_arr_23__1 ;
    input q_arr_23__0 ;
    input q_arr_24__31 ;
    input q_arr_24__30 ;
    input q_arr_24__29 ;
    input q_arr_24__28 ;
    input q_arr_24__27 ;
    input q_arr_24__26 ;
    input q_arr_24__25 ;
    input q_arr_24__24 ;
    input q_arr_24__23 ;
    input q_arr_24__22 ;
    input q_arr_24__21 ;
    input q_arr_24__20 ;
    input q_arr_24__19 ;
    input q_arr_24__18 ;
    input q_arr_24__17 ;
    input q_arr_24__16 ;
    input q_arr_24__15 ;
    input q_arr_24__14 ;
    input q_arr_24__13 ;
    input q_arr_24__12 ;
    input q_arr_24__11 ;
    input q_arr_24__10 ;
    input q_arr_24__9 ;
    input q_arr_24__8 ;
    input q_arr_24__7 ;
    input q_arr_24__6 ;
    input q_arr_24__5 ;
    input q_arr_24__4 ;
    input q_arr_24__3 ;
    input q_arr_24__2 ;
    input q_arr_24__1 ;
    input q_arr_24__0 ;
    input [15:0]output1_init ;
    input [15:0]output2_init ;
    input filter_size ;
    input operation ;
    input compute_relu ;
    input clk ;
    input en ;
    input reset ;
    output buffer_ready ;
    output semi_ready ;
    output ready ;

    wire counter_15, counter_14, counter_13, counter_0, 
         ordered_filter_data_3__15, ordered_filter_data_3__14, 
         ordered_filter_data_3__13, ordered_filter_data_3__12, 
         ordered_filter_data_3__11, ordered_filter_data_3__10, 
         ordered_filter_data_3__9, ordered_filter_data_3__8, 
         ordered_filter_data_3__7, ordered_filter_data_3__6, 
         ordered_filter_data_3__5, ordered_filter_data_3__4, 
         ordered_filter_data_3__3, ordered_filter_data_3__2, 
         ordered_filter_data_3__1, ordered_filter_data_3__0, 
         ordered_filter_data_4__15, ordered_filter_data_4__14, 
         ordered_filter_data_4__13, ordered_filter_data_4__12, 
         ordered_filter_data_4__11, ordered_filter_data_4__10, 
         ordered_filter_data_4__9, ordered_filter_data_4__8, 
         ordered_filter_data_4__7, ordered_filter_data_4__6, 
         ordered_filter_data_4__5, ordered_filter_data_4__4, 
         ordered_filter_data_4__3, ordered_filter_data_4__2, 
         ordered_filter_data_4__1, ordered_filter_data_4__0, 
         ordered_filter_data_5__15, ordered_filter_data_5__14, 
         ordered_filter_data_5__13, ordered_filter_data_5__12, 
         ordered_filter_data_5__11, ordered_filter_data_5__10, 
         ordered_filter_data_5__9, ordered_filter_data_5__8, 
         ordered_filter_data_5__7, ordered_filter_data_5__6, 
         ordered_filter_data_5__5, ordered_filter_data_5__4, 
         ordered_filter_data_5__3, ordered_filter_data_5__2, 
         ordered_filter_data_5__1, ordered_filter_data_5__0, 
         ordered_filter_data_6__15, ordered_filter_data_6__14, 
         ordered_filter_data_6__13, ordered_filter_data_6__12, 
         ordered_filter_data_6__11, ordered_filter_data_6__10, 
         ordered_filter_data_6__9, ordered_filter_data_6__8, 
         ordered_filter_data_6__7, ordered_filter_data_6__6, 
         ordered_filter_data_6__5, ordered_filter_data_6__4, 
         ordered_filter_data_6__3, ordered_filter_data_6__2, 
         ordered_filter_data_6__1, ordered_filter_data_6__0, 
         ordered_filter_data_7__15, ordered_filter_data_7__14, 
         ordered_filter_data_7__13, ordered_filter_data_7__12, 
         ordered_filter_data_7__11, ordered_filter_data_7__10, 
         ordered_filter_data_7__9, ordered_filter_data_7__8, 
         ordered_filter_data_7__7, ordered_filter_data_7__6, 
         ordered_filter_data_7__5, ordered_filter_data_7__4, 
         ordered_filter_data_7__3, ordered_filter_data_7__2, 
         ordered_filter_data_7__1, ordered_filter_data_7__0, 
         ordered_filter_data_8__15, ordered_filter_data_8__14, 
         ordered_filter_data_8__13, ordered_filter_data_8__12, 
         ordered_filter_data_8__11, ordered_filter_data_8__10, 
         ordered_filter_data_8__9, ordered_filter_data_8__8, 
         ordered_filter_data_8__7, ordered_filter_data_8__6, 
         ordered_filter_data_8__5, ordered_filter_data_8__4, 
         ordered_filter_data_8__3, ordered_filter_data_8__2, 
         ordered_filter_data_8__1, ordered_filter_data_8__0, 
         ordered_filter_data_9__15, ordered_filter_data_9__14, 
         ordered_filter_data_9__13, ordered_filter_data_9__12, 
         ordered_filter_data_9__11, ordered_filter_data_9__10, 
         ordered_filter_data_9__9, ordered_filter_data_9__8, 
         ordered_filter_data_9__7, ordered_filter_data_9__6, 
         ordered_filter_data_9__5, ordered_filter_data_9__4, 
         ordered_filter_data_9__3, ordered_filter_data_9__2, 
         ordered_filter_data_9__1, ordered_filter_data_9__0, 
         ordered_filter_data_10__15, ordered_filter_data_10__14, 
         ordered_filter_data_10__13, ordered_filter_data_10__12, 
         ordered_filter_data_10__11, ordered_filter_data_10__10, 
         ordered_filter_data_10__9, ordered_filter_data_10__8, 
         ordered_filter_data_10__7, ordered_filter_data_10__6, 
         ordered_filter_data_10__5, ordered_filter_data_10__4, 
         ordered_filter_data_10__3, ordered_filter_data_10__2, 
         ordered_filter_data_10__1, ordered_filter_data_10__0, 
         ordered_filter_data_11__15, ordered_filter_data_11__14, 
         ordered_filter_data_11__13, ordered_filter_data_11__12, 
         ordered_filter_data_11__11, ordered_filter_data_11__10, 
         ordered_filter_data_11__9, ordered_filter_data_11__8, 
         ordered_filter_data_11__7, ordered_filter_data_11__6, 
         ordered_filter_data_11__5, ordered_filter_data_11__4, 
         ordered_filter_data_11__3, ordered_filter_data_11__2, 
         ordered_filter_data_11__1, ordered_filter_data_11__0, 
         ordered_filter_data_12__15, ordered_filter_data_12__14, 
         ordered_filter_data_12__13, ordered_filter_data_12__12, 
         ordered_filter_data_12__11, ordered_filter_data_12__10, 
         ordered_filter_data_12__9, ordered_filter_data_12__8, 
         ordered_filter_data_12__7, ordered_filter_data_12__6, 
         ordered_filter_data_12__5, ordered_filter_data_12__4, 
         ordered_filter_data_12__3, ordered_filter_data_12__2, 
         ordered_filter_data_12__1, ordered_filter_data_12__0, 
         ordered_filter_data_13__15, ordered_filter_data_13__14, 
         ordered_filter_data_13__13, ordered_filter_data_13__12, 
         ordered_filter_data_13__11, ordered_filter_data_13__10, 
         ordered_filter_data_13__9, ordered_filter_data_13__8, 
         ordered_filter_data_13__7, ordered_filter_data_13__6, 
         ordered_filter_data_13__5, ordered_filter_data_13__4, 
         ordered_filter_data_13__3, ordered_filter_data_13__2, 
         ordered_filter_data_13__1, ordered_filter_data_13__0, 
         ordered_filter_data_14__15, ordered_filter_data_14__14, 
         ordered_filter_data_14__13, ordered_filter_data_14__12, 
         ordered_filter_data_14__11, ordered_filter_data_14__10, 
         ordered_filter_data_14__9, ordered_filter_data_14__8, 
         ordered_filter_data_14__7, ordered_filter_data_14__6, 
         ordered_filter_data_14__5, ordered_filter_data_14__4, 
         ordered_filter_data_14__3, ordered_filter_data_14__2, 
         ordered_filter_data_14__1, ordered_filter_data_14__0, 
         ordered_filter_data_15__15, ordered_filter_data_15__14, 
         ordered_filter_data_15__13, ordered_filter_data_15__12, 
         ordered_filter_data_15__11, ordered_filter_data_15__10, 
         ordered_filter_data_15__9, ordered_filter_data_15__8, 
         ordered_filter_data_15__7, ordered_filter_data_15__6, 
         ordered_filter_data_15__5, ordered_filter_data_15__4, 
         ordered_filter_data_15__3, ordered_filter_data_15__2, 
         ordered_filter_data_15__1, ordered_filter_data_15__0, 
         ordered_filter_data_16__15, ordered_filter_data_16__14, 
         ordered_filter_data_16__13, ordered_filter_data_16__12, 
         ordered_filter_data_16__11, ordered_filter_data_16__10, 
         ordered_filter_data_16__9, ordered_filter_data_16__8, 
         ordered_filter_data_16__7, ordered_filter_data_16__6, 
         ordered_filter_data_16__5, ordered_filter_data_16__4, 
         ordered_filter_data_16__3, ordered_filter_data_16__2, 
         ordered_filter_data_16__1, ordered_filter_data_16__0, 
         ordered_filter_data_17__15, ordered_filter_data_17__14, 
         ordered_filter_data_17__13, ordered_filter_data_17__12, 
         ordered_filter_data_17__11, ordered_filter_data_17__10, 
         ordered_filter_data_17__9, ordered_filter_data_17__8, 
         ordered_filter_data_17__7, ordered_filter_data_17__6, 
         ordered_filter_data_17__5, ordered_filter_data_17__4, 
         ordered_filter_data_17__3, ordered_filter_data_17__2, 
         ordered_filter_data_17__1, ordered_filter_data_17__0, 
         ordered_img_data_9__31, ordered_img_data_9__14, ordered_img_data_9__13, 
         ordered_img_data_9__12, ordered_img_data_9__11, ordered_img_data_9__10, 
         ordered_img_data_9__9, ordered_img_data_9__8, ordered_img_data_9__7, 
         ordered_img_data_9__6, ordered_img_data_9__5, ordered_img_data_9__4, 
         ordered_img_data_9__3, ordered_img_data_9__2, ordered_img_data_9__1, 
         ordered_img_data_9__0, ordered_img_data_10__31, ordered_img_data_10__14, 
         ordered_img_data_10__13, ordered_img_data_10__12, 
         ordered_img_data_10__11, ordered_img_data_10__10, 
         ordered_img_data_10__9, ordered_img_data_10__8, ordered_img_data_10__7, 
         ordered_img_data_10__6, ordered_img_data_10__5, ordered_img_data_10__4, 
         ordered_img_data_10__3, ordered_img_data_10__2, ordered_img_data_10__1, 
         ordered_img_data_10__0, ordered_img_data_11__31, 
         ordered_img_data_11__14, ordered_img_data_11__13, 
         ordered_img_data_11__12, ordered_img_data_11__11, 
         ordered_img_data_11__10, ordered_img_data_11__9, ordered_img_data_11__8, 
         ordered_img_data_11__7, ordered_img_data_11__6, ordered_img_data_11__5, 
         ordered_img_data_11__4, ordered_img_data_11__3, ordered_img_data_11__2, 
         ordered_img_data_11__1, ordered_img_data_11__0, ordered_img_data_12__31, 
         ordered_img_data_12__14, ordered_img_data_12__13, 
         ordered_img_data_12__12, ordered_img_data_12__11, 
         ordered_img_data_12__10, ordered_img_data_12__9, ordered_img_data_12__8, 
         ordered_img_data_12__7, ordered_img_data_12__6, ordered_img_data_12__5, 
         ordered_img_data_12__4, ordered_img_data_12__3, ordered_img_data_12__2, 
         ordered_img_data_12__1, ordered_img_data_12__0, ordered_img_data_13__31, 
         ordered_img_data_13__14, ordered_img_data_13__13, 
         ordered_img_data_13__12, ordered_img_data_13__11, 
         ordered_img_data_13__10, ordered_img_data_13__9, ordered_img_data_13__8, 
         ordered_img_data_13__7, ordered_img_data_13__6, ordered_img_data_13__5, 
         ordered_img_data_13__4, ordered_img_data_13__3, ordered_img_data_13__2, 
         ordered_img_data_13__1, ordered_img_data_13__0, ordered_img_data_14__31, 
         ordered_img_data_14__14, ordered_img_data_14__13, 
         ordered_img_data_14__12, ordered_img_data_14__11, 
         ordered_img_data_14__10, ordered_img_data_14__9, ordered_img_data_14__8, 
         ordered_img_data_14__7, ordered_img_data_14__6, ordered_img_data_14__5, 
         ordered_img_data_14__4, ordered_img_data_14__3, ordered_img_data_14__2, 
         ordered_img_data_14__1, ordered_img_data_14__0, ordered_img_data_15__31, 
         ordered_img_data_15__14, ordered_img_data_15__13, 
         ordered_img_data_15__12, ordered_img_data_15__11, 
         ordered_img_data_15__10, ordered_img_data_15__9, ordered_img_data_15__8, 
         ordered_img_data_15__7, ordered_img_data_15__6, ordered_img_data_15__5, 
         ordered_img_data_15__4, ordered_img_data_15__3, ordered_img_data_15__2, 
         ordered_img_data_15__1, ordered_img_data_15__0, ordered_img_data_16__31, 
         ordered_img_data_16__14, ordered_img_data_16__13, 
         ordered_img_data_16__12, ordered_img_data_16__11, 
         ordered_img_data_16__10, ordered_img_data_16__9, ordered_img_data_16__8, 
         ordered_img_data_16__7, ordered_img_data_16__6, ordered_img_data_16__5, 
         ordered_img_data_16__4, ordered_img_data_16__3, ordered_img_data_16__2, 
         ordered_img_data_16__1, ordered_img_data_16__0, ordered_img_data_17__31, 
         ordered_img_data_17__14, ordered_img_data_17__13, 
         ordered_img_data_17__12, ordered_img_data_17__11, 
         ordered_img_data_17__10, ordered_img_data_17__9, ordered_img_data_17__8, 
         ordered_img_data_17__7, ordered_img_data_17__6, ordered_img_data_17__5, 
         ordered_img_data_17__4, ordered_img_data_17__3, ordered_img_data_17__2, 
         ordered_img_data_17__1, ordered_img_data_17__0, d_arr_mul_0__31, 
         d_arr_mul_0__30, d_arr_mul_0__29, d_arr_mul_0__28, d_arr_mul_0__27, 
         d_arr_mul_0__26, d_arr_mul_0__25, d_arr_mul_0__24, d_arr_mul_0__23, 
         d_arr_mul_0__22, d_arr_mul_0__21, d_arr_mul_0__20, d_arr_mul_0__19, 
         d_arr_mul_0__18, d_arr_mul_0__17, d_arr_mul_0__16, d_arr_mul_0__15, 
         d_arr_mul_0__14, d_arr_mul_0__13, d_arr_mul_0__12, d_arr_mul_0__11, 
         d_arr_mul_0__10, d_arr_mul_0__9, d_arr_mul_0__8, d_arr_mul_0__7, 
         d_arr_mul_0__6, d_arr_mul_0__5, d_arr_mul_0__4, d_arr_mul_0__3, 
         d_arr_mul_0__2, d_arr_mul_0__1, d_arr_mul_0__0, d_arr_mul_1__31, 
         d_arr_mul_1__30, d_arr_mul_1__29, d_arr_mul_1__28, d_arr_mul_1__27, 
         d_arr_mul_1__26, d_arr_mul_1__25, d_arr_mul_1__24, d_arr_mul_1__23, 
         d_arr_mul_1__22, d_arr_mul_1__21, d_arr_mul_1__20, d_arr_mul_1__19, 
         d_arr_mul_1__18, d_arr_mul_1__17, d_arr_mul_1__16, d_arr_mul_1__15, 
         d_arr_mul_1__14, d_arr_mul_1__13, d_arr_mul_1__12, d_arr_mul_1__11, 
         d_arr_mul_1__10, d_arr_mul_1__9, d_arr_mul_1__8, d_arr_mul_1__7, 
         d_arr_mul_1__6, d_arr_mul_1__5, d_arr_mul_1__4, d_arr_mul_1__3, 
         d_arr_mul_1__2, d_arr_mul_1__1, d_arr_mul_1__0, d_arr_mul_2__31, 
         d_arr_mul_2__30, d_arr_mul_2__29, d_arr_mul_2__28, d_arr_mul_2__27, 
         d_arr_mul_2__26, d_arr_mul_2__25, d_arr_mul_2__24, d_arr_mul_2__23, 
         d_arr_mul_2__22, d_arr_mul_2__21, d_arr_mul_2__20, d_arr_mul_2__19, 
         d_arr_mul_2__18, d_arr_mul_2__17, d_arr_mul_2__16, d_arr_mul_2__15, 
         d_arr_mul_2__14, d_arr_mul_2__13, d_arr_mul_2__12, d_arr_mul_2__11, 
         d_arr_mul_2__10, d_arr_mul_2__9, d_arr_mul_2__8, d_arr_mul_2__7, 
         d_arr_mul_2__6, d_arr_mul_2__5, d_arr_mul_2__4, d_arr_mul_2__3, 
         d_arr_mul_2__2, d_arr_mul_2__1, d_arr_mul_2__0, d_arr_mul_3__31, 
         d_arr_mul_3__30, d_arr_mul_3__29, d_arr_mul_3__28, d_arr_mul_3__27, 
         d_arr_mul_3__26, d_arr_mul_3__25, d_arr_mul_3__24, d_arr_mul_3__23, 
         d_arr_mul_3__22, d_arr_mul_3__21, d_arr_mul_3__20, d_arr_mul_3__19, 
         d_arr_mul_3__18, d_arr_mul_3__17, d_arr_mul_3__16, d_arr_mul_3__15, 
         d_arr_mul_3__14, d_arr_mul_3__13, d_arr_mul_3__12, d_arr_mul_3__11, 
         d_arr_mul_3__10, d_arr_mul_3__9, d_arr_mul_3__8, d_arr_mul_3__7, 
         d_arr_mul_3__6, d_arr_mul_3__5, d_arr_mul_3__4, d_arr_mul_3__3, 
         d_arr_mul_3__2, d_arr_mul_3__1, d_arr_mul_3__0, d_arr_mul_4__31, 
         d_arr_mul_4__30, d_arr_mul_4__29, d_arr_mul_4__28, d_arr_mul_4__27, 
         d_arr_mul_4__26, d_arr_mul_4__25, d_arr_mul_4__24, d_arr_mul_4__23, 
         d_arr_mul_4__22, d_arr_mul_4__21, d_arr_mul_4__20, d_arr_mul_4__19, 
         d_arr_mul_4__18, d_arr_mul_4__17, d_arr_mul_4__16, d_arr_mul_4__15, 
         d_arr_mul_4__14, d_arr_mul_4__13, d_arr_mul_4__12, d_arr_mul_4__11, 
         d_arr_mul_4__10, d_arr_mul_4__9, d_arr_mul_4__8, d_arr_mul_4__7, 
         d_arr_mul_4__6, d_arr_mul_4__5, d_arr_mul_4__4, d_arr_mul_4__3, 
         d_arr_mul_4__2, d_arr_mul_4__1, d_arr_mul_4__0, d_arr_mul_5__31, 
         d_arr_mul_5__30, d_arr_mul_5__29, d_arr_mul_5__28, d_arr_mul_5__27, 
         d_arr_mul_5__26, d_arr_mul_5__25, d_arr_mul_5__24, d_arr_mul_5__23, 
         d_arr_mul_5__22, d_arr_mul_5__21, d_arr_mul_5__20, d_arr_mul_5__19, 
         d_arr_mul_5__18, d_arr_mul_5__17, d_arr_mul_5__16, d_arr_mul_5__15, 
         d_arr_mul_5__14, d_arr_mul_5__13, d_arr_mul_5__12, d_arr_mul_5__11, 
         d_arr_mul_5__10, d_arr_mul_5__9, d_arr_mul_5__8, d_arr_mul_5__7, 
         d_arr_mul_5__6, d_arr_mul_5__5, d_arr_mul_5__4, d_arr_mul_5__3, 
         d_arr_mul_5__2, d_arr_mul_5__1, d_arr_mul_5__0, d_arr_mul_6__31, 
         d_arr_mul_6__30, d_arr_mul_6__29, d_arr_mul_6__28, d_arr_mul_6__27, 
         d_arr_mul_6__26, d_arr_mul_6__25, d_arr_mul_6__24, d_arr_mul_6__23, 
         d_arr_mul_6__22, d_arr_mul_6__21, d_arr_mul_6__20, d_arr_mul_6__19, 
         d_arr_mul_6__18, d_arr_mul_6__17, d_arr_mul_6__16, d_arr_mul_6__15, 
         d_arr_mul_6__14, d_arr_mul_6__13, d_arr_mul_6__12, d_arr_mul_6__11, 
         d_arr_mul_6__10, d_arr_mul_6__9, d_arr_mul_6__8, d_arr_mul_6__7, 
         d_arr_mul_6__6, d_arr_mul_6__5, d_arr_mul_6__4, d_arr_mul_6__3, 
         d_arr_mul_6__2, d_arr_mul_6__1, d_arr_mul_6__0, d_arr_mul_7__31, 
         d_arr_mul_7__30, d_arr_mul_7__29, d_arr_mul_7__28, d_arr_mul_7__27, 
         d_arr_mul_7__26, d_arr_mul_7__25, d_arr_mul_7__24, d_arr_mul_7__23, 
         d_arr_mul_7__22, d_arr_mul_7__21, d_arr_mul_7__20, d_arr_mul_7__19, 
         d_arr_mul_7__18, d_arr_mul_7__17, d_arr_mul_7__16, d_arr_mul_7__15, 
         d_arr_mul_7__14, d_arr_mul_7__13, d_arr_mul_7__12, d_arr_mul_7__11, 
         d_arr_mul_7__10, d_arr_mul_7__9, d_arr_mul_7__8, d_arr_mul_7__7, 
         d_arr_mul_7__6, d_arr_mul_7__5, d_arr_mul_7__4, d_arr_mul_7__3, 
         d_arr_mul_7__2, d_arr_mul_7__1, d_arr_mul_7__0, d_arr_mul_8__31, 
         d_arr_mul_8__30, d_arr_mul_8__29, d_arr_mul_8__28, d_arr_mul_8__27, 
         d_arr_mul_8__26, d_arr_mul_8__25, d_arr_mul_8__24, d_arr_mul_8__23, 
         d_arr_mul_8__22, d_arr_mul_8__21, d_arr_mul_8__20, d_arr_mul_8__19, 
         d_arr_mul_8__18, d_arr_mul_8__17, d_arr_mul_8__16, d_arr_mul_8__15, 
         d_arr_mul_8__14, d_arr_mul_8__13, d_arr_mul_8__12, d_arr_mul_8__11, 
         d_arr_mul_8__10, d_arr_mul_8__9, d_arr_mul_8__8, d_arr_mul_8__7, 
         d_arr_mul_8__6, d_arr_mul_8__5, d_arr_mul_8__4, d_arr_mul_8__3, 
         d_arr_mul_8__2, d_arr_mul_8__1, d_arr_mul_8__0, d_arr_mul_9__31, 
         d_arr_mul_9__30, d_arr_mul_9__29, d_arr_mul_9__28, d_arr_mul_9__27, 
         d_arr_mul_9__26, d_arr_mul_9__25, d_arr_mul_9__24, d_arr_mul_9__23, 
         d_arr_mul_9__22, d_arr_mul_9__21, d_arr_mul_9__20, d_arr_mul_9__19, 
         d_arr_mul_9__18, d_arr_mul_9__17, d_arr_mul_9__16, d_arr_mul_9__15, 
         d_arr_mul_9__14, d_arr_mul_9__13, d_arr_mul_9__12, d_arr_mul_9__11, 
         d_arr_mul_9__10, d_arr_mul_9__9, d_arr_mul_9__8, d_arr_mul_9__7, 
         d_arr_mul_9__6, d_arr_mul_9__5, d_arr_mul_9__4, d_arr_mul_9__3, 
         d_arr_mul_9__2, d_arr_mul_9__1, d_arr_mul_9__0, d_arr_mul_10__31, 
         d_arr_mul_10__30, d_arr_mul_10__29, d_arr_mul_10__28, d_arr_mul_10__27, 
         d_arr_mul_10__26, d_arr_mul_10__25, d_arr_mul_10__24, d_arr_mul_10__23, 
         d_arr_mul_10__22, d_arr_mul_10__21, d_arr_mul_10__20, d_arr_mul_10__19, 
         d_arr_mul_10__18, d_arr_mul_10__17, d_arr_mul_10__16, d_arr_mul_10__15, 
         d_arr_mul_10__14, d_arr_mul_10__13, d_arr_mul_10__12, d_arr_mul_10__11, 
         d_arr_mul_10__10, d_arr_mul_10__9, d_arr_mul_10__8, d_arr_mul_10__7, 
         d_arr_mul_10__6, d_arr_mul_10__5, d_arr_mul_10__4, d_arr_mul_10__3, 
         d_arr_mul_10__2, d_arr_mul_10__1, d_arr_mul_10__0, d_arr_mul_11__31, 
         d_arr_mul_11__30, d_arr_mul_11__29, d_arr_mul_11__28, d_arr_mul_11__27, 
         d_arr_mul_11__26, d_arr_mul_11__25, d_arr_mul_11__24, d_arr_mul_11__23, 
         d_arr_mul_11__22, d_arr_mul_11__21, d_arr_mul_11__20, d_arr_mul_11__19, 
         d_arr_mul_11__18, d_arr_mul_11__17, d_arr_mul_11__16, d_arr_mul_11__15, 
         d_arr_mul_11__14, d_arr_mul_11__13, d_arr_mul_11__12, d_arr_mul_11__11, 
         d_arr_mul_11__10, d_arr_mul_11__9, d_arr_mul_11__8, d_arr_mul_11__7, 
         d_arr_mul_11__6, d_arr_mul_11__5, d_arr_mul_11__4, d_arr_mul_11__3, 
         d_arr_mul_11__2, d_arr_mul_11__1, d_arr_mul_11__0, d_arr_mul_12__31, 
         d_arr_mul_12__30, d_arr_mul_12__29, d_arr_mul_12__28, d_arr_mul_12__27, 
         d_arr_mul_12__26, d_arr_mul_12__25, d_arr_mul_12__24, d_arr_mul_12__23, 
         d_arr_mul_12__22, d_arr_mul_12__21, d_arr_mul_12__20, d_arr_mul_12__19, 
         d_arr_mul_12__18, d_arr_mul_12__17, d_arr_mul_12__16, d_arr_mul_12__15, 
         d_arr_mul_12__14, d_arr_mul_12__13, d_arr_mul_12__12, d_arr_mul_12__11, 
         d_arr_mul_12__10, d_arr_mul_12__9, d_arr_mul_12__8, d_arr_mul_12__7, 
         d_arr_mul_12__6, d_arr_mul_12__5, d_arr_mul_12__4, d_arr_mul_12__3, 
         d_arr_mul_12__2, d_arr_mul_12__1, d_arr_mul_12__0, d_arr_mul_13__31, 
         d_arr_mul_13__30, d_arr_mul_13__29, d_arr_mul_13__28, d_arr_mul_13__27, 
         d_arr_mul_13__26, d_arr_mul_13__25, d_arr_mul_13__24, d_arr_mul_13__23, 
         d_arr_mul_13__22, d_arr_mul_13__21, d_arr_mul_13__20, d_arr_mul_13__19, 
         d_arr_mul_13__18, d_arr_mul_13__17, d_arr_mul_13__16, d_arr_mul_13__15, 
         d_arr_mul_13__14, d_arr_mul_13__13, d_arr_mul_13__12, d_arr_mul_13__11, 
         d_arr_mul_13__10, d_arr_mul_13__9, d_arr_mul_13__8, d_arr_mul_13__7, 
         d_arr_mul_13__6, d_arr_mul_13__5, d_arr_mul_13__4, d_arr_mul_13__3, 
         d_arr_mul_13__2, d_arr_mul_13__1, d_arr_mul_13__0, d_arr_mul_14__31, 
         d_arr_mul_14__30, d_arr_mul_14__29, d_arr_mul_14__28, d_arr_mul_14__27, 
         d_arr_mul_14__26, d_arr_mul_14__25, d_arr_mul_14__24, d_arr_mul_14__23, 
         d_arr_mul_14__22, d_arr_mul_14__21, d_arr_mul_14__20, d_arr_mul_14__19, 
         d_arr_mul_14__18, d_arr_mul_14__17, d_arr_mul_14__16, d_arr_mul_14__15, 
         d_arr_mul_14__14, d_arr_mul_14__13, d_arr_mul_14__12, d_arr_mul_14__11, 
         d_arr_mul_14__10, d_arr_mul_14__9, d_arr_mul_14__8, d_arr_mul_14__7, 
         d_arr_mul_14__6, d_arr_mul_14__5, d_arr_mul_14__4, d_arr_mul_14__3, 
         d_arr_mul_14__2, d_arr_mul_14__1, d_arr_mul_14__0, d_arr_mul_15__31, 
         d_arr_mul_15__30, d_arr_mul_15__29, d_arr_mul_15__28, d_arr_mul_15__27, 
         d_arr_mul_15__26, d_arr_mul_15__25, d_arr_mul_15__24, d_arr_mul_15__23, 
         d_arr_mul_15__22, d_arr_mul_15__21, d_arr_mul_15__20, d_arr_mul_15__19, 
         d_arr_mul_15__18, d_arr_mul_15__17, d_arr_mul_15__16, d_arr_mul_15__15, 
         d_arr_mul_15__14, d_arr_mul_15__13, d_arr_mul_15__12, d_arr_mul_15__11, 
         d_arr_mul_15__10, d_arr_mul_15__9, d_arr_mul_15__8, d_arr_mul_15__7, 
         d_arr_mul_15__6, d_arr_mul_15__5, d_arr_mul_15__4, d_arr_mul_15__3, 
         d_arr_mul_15__2, d_arr_mul_15__1, d_arr_mul_15__0, d_arr_mul_16__31, 
         d_arr_mul_16__30, d_arr_mul_16__29, d_arr_mul_16__28, d_arr_mul_16__27, 
         d_arr_mul_16__26, d_arr_mul_16__25, d_arr_mul_16__24, d_arr_mul_16__23, 
         d_arr_mul_16__22, d_arr_mul_16__21, d_arr_mul_16__20, d_arr_mul_16__19, 
         d_arr_mul_16__18, d_arr_mul_16__17, d_arr_mul_16__16, d_arr_mul_16__15, 
         d_arr_mul_16__14, d_arr_mul_16__13, d_arr_mul_16__12, d_arr_mul_16__11, 
         d_arr_mul_16__10, d_arr_mul_16__9, d_arr_mul_16__8, d_arr_mul_16__7, 
         d_arr_mul_16__6, d_arr_mul_16__5, d_arr_mul_16__4, d_arr_mul_16__3, 
         d_arr_mul_16__2, d_arr_mul_16__1, d_arr_mul_16__0, d_arr_mul_17__31, 
         d_arr_mul_17__30, d_arr_mul_17__29, d_arr_mul_17__28, d_arr_mul_17__27, 
         d_arr_mul_17__26, d_arr_mul_17__25, d_arr_mul_17__24, d_arr_mul_17__23, 
         d_arr_mul_17__22, d_arr_mul_17__21, d_arr_mul_17__20, d_arr_mul_17__19, 
         d_arr_mul_17__18, d_arr_mul_17__17, d_arr_mul_17__16, d_arr_mul_17__15, 
         d_arr_mul_17__14, d_arr_mul_17__13, d_arr_mul_17__12, d_arr_mul_17__11, 
         d_arr_mul_17__10, d_arr_mul_17__9, d_arr_mul_17__8, d_arr_mul_17__7, 
         d_arr_mul_17__6, d_arr_mul_17__5, d_arr_mul_17__4, d_arr_mul_17__3, 
         d_arr_mul_17__2, d_arr_mul_17__1, d_arr_mul_17__0, d_arr_mul_18__31, 
         d_arr_mul_18__30, d_arr_mul_18__29, d_arr_mul_18__28, d_arr_mul_18__27, 
         d_arr_mul_18__26, d_arr_mul_18__25, d_arr_mul_18__24, d_arr_mul_18__23, 
         d_arr_mul_18__22, d_arr_mul_18__21, d_arr_mul_18__20, d_arr_mul_18__19, 
         d_arr_mul_18__18, d_arr_mul_18__17, d_arr_mul_18__16, d_arr_mul_18__15, 
         d_arr_mul_18__14, d_arr_mul_18__13, d_arr_mul_18__12, d_arr_mul_18__11, 
         d_arr_mul_18__10, d_arr_mul_18__9, d_arr_mul_18__8, d_arr_mul_18__7, 
         d_arr_mul_18__6, d_arr_mul_18__5, d_arr_mul_18__4, d_arr_mul_18__3, 
         d_arr_mul_18__2, d_arr_mul_18__1, d_arr_mul_18__0, d_arr_mul_19__31, 
         d_arr_mul_19__30, d_arr_mul_19__29, d_arr_mul_19__28, d_arr_mul_19__27, 
         d_arr_mul_19__26, d_arr_mul_19__25, d_arr_mul_19__24, d_arr_mul_19__23, 
         d_arr_mul_19__22, d_arr_mul_19__21, d_arr_mul_19__20, d_arr_mul_19__19, 
         d_arr_mul_19__18, d_arr_mul_19__17, d_arr_mul_19__16, d_arr_mul_19__15, 
         d_arr_mul_19__14, d_arr_mul_19__13, d_arr_mul_19__12, d_arr_mul_19__11, 
         d_arr_mul_19__10, d_arr_mul_19__9, d_arr_mul_19__8, d_arr_mul_19__7, 
         d_arr_mul_19__6, d_arr_mul_19__5, d_arr_mul_19__4, d_arr_mul_19__3, 
         d_arr_mul_19__2, d_arr_mul_19__1, d_arr_mul_19__0, d_arr_mul_20__31, 
         d_arr_mul_20__30, d_arr_mul_20__29, d_arr_mul_20__28, d_arr_mul_20__27, 
         d_arr_mul_20__26, d_arr_mul_20__25, d_arr_mul_20__24, d_arr_mul_20__23, 
         d_arr_mul_20__22, d_arr_mul_20__21, d_arr_mul_20__20, d_arr_mul_20__19, 
         d_arr_mul_20__18, d_arr_mul_20__17, d_arr_mul_20__16, d_arr_mul_20__15, 
         d_arr_mul_20__14, d_arr_mul_20__13, d_arr_mul_20__12, d_arr_mul_20__11, 
         d_arr_mul_20__10, d_arr_mul_20__9, d_arr_mul_20__8, d_arr_mul_20__7, 
         d_arr_mul_20__6, d_arr_mul_20__5, d_arr_mul_20__4, d_arr_mul_20__3, 
         d_arr_mul_20__2, d_arr_mul_20__1, d_arr_mul_20__0, d_arr_mul_21__31, 
         d_arr_mul_21__30, d_arr_mul_21__29, d_arr_mul_21__28, d_arr_mul_21__27, 
         d_arr_mul_21__26, d_arr_mul_21__25, d_arr_mul_21__24, d_arr_mul_21__23, 
         d_arr_mul_21__22, d_arr_mul_21__21, d_arr_mul_21__20, d_arr_mul_21__19, 
         d_arr_mul_21__18, d_arr_mul_21__17, d_arr_mul_21__16, d_arr_mul_21__15, 
         d_arr_mul_21__14, d_arr_mul_21__13, d_arr_mul_21__12, d_arr_mul_21__11, 
         d_arr_mul_21__10, d_arr_mul_21__9, d_arr_mul_21__8, d_arr_mul_21__7, 
         d_arr_mul_21__6, d_arr_mul_21__5, d_arr_mul_21__4, d_arr_mul_21__3, 
         d_arr_mul_21__2, d_arr_mul_21__1, d_arr_mul_21__0, d_arr_mul_22__31, 
         d_arr_mul_22__30, d_arr_mul_22__29, d_arr_mul_22__28, d_arr_mul_22__27, 
         d_arr_mul_22__26, d_arr_mul_22__25, d_arr_mul_22__24, d_arr_mul_22__23, 
         d_arr_mul_22__22, d_arr_mul_22__21, d_arr_mul_22__20, d_arr_mul_22__19, 
         d_arr_mul_22__18, d_arr_mul_22__17, d_arr_mul_22__16, d_arr_mul_22__15, 
         d_arr_mul_22__14, d_arr_mul_22__13, d_arr_mul_22__12, d_arr_mul_22__11, 
         d_arr_mul_22__10, d_arr_mul_22__9, d_arr_mul_22__8, d_arr_mul_22__7, 
         d_arr_mul_22__6, d_arr_mul_22__5, d_arr_mul_22__4, d_arr_mul_22__3, 
         d_arr_mul_22__2, d_arr_mul_22__1, d_arr_mul_22__0, d_arr_mul_23__31, 
         d_arr_mul_23__30, d_arr_mul_23__29, d_arr_mul_23__28, d_arr_mul_23__27, 
         d_arr_mul_23__26, d_arr_mul_23__25, d_arr_mul_23__24, d_arr_mul_23__23, 
         d_arr_mul_23__22, d_arr_mul_23__21, d_arr_mul_23__20, d_arr_mul_23__19, 
         d_arr_mul_23__18, d_arr_mul_23__17, d_arr_mul_23__16, d_arr_mul_23__15, 
         d_arr_mul_23__14, d_arr_mul_23__13, d_arr_mul_23__12, d_arr_mul_23__11, 
         d_arr_mul_23__10, d_arr_mul_23__9, d_arr_mul_23__8, d_arr_mul_23__7, 
         d_arr_mul_23__6, d_arr_mul_23__5, d_arr_mul_23__4, d_arr_mul_23__3, 
         d_arr_mul_23__2, d_arr_mul_23__1, d_arr_mul_23__0, d_arr_mul_24__31, 
         d_arr_mul_24__30, d_arr_mul_24__29, d_arr_mul_24__28, d_arr_mul_24__27, 
         d_arr_mul_24__26, d_arr_mul_24__25, d_arr_mul_24__24, d_arr_mul_24__23, 
         d_arr_mul_24__22, d_arr_mul_24__21, d_arr_mul_24__20, d_arr_mul_24__19, 
         d_arr_mul_24__18, d_arr_mul_24__17, d_arr_mul_24__16, d_arr_mul_24__15, 
         d_arr_mul_24__14, d_arr_mul_24__13, d_arr_mul_24__12, d_arr_mul_24__11, 
         d_arr_mul_24__10, d_arr_mul_24__9, d_arr_mul_24__8, d_arr_mul_24__7, 
         d_arr_mul_24__6, d_arr_mul_24__5, d_arr_mul_24__4, d_arr_mul_24__3, 
         d_arr_mul_24__2, d_arr_mul_24__1, d_arr_mul_24__0, d_arr_add_0__31, 
         d_arr_add_0__30, d_arr_add_0__29, d_arr_add_0__28, d_arr_add_0__27, 
         d_arr_add_0__26, d_arr_add_0__25, d_arr_add_0__24, d_arr_add_0__23, 
         d_arr_add_0__22, d_arr_add_0__21, d_arr_add_0__20, d_arr_add_0__19, 
         d_arr_add_0__18, d_arr_add_0__17, d_arr_add_0__16, d_arr_add_0__15, 
         d_arr_add_0__14, d_arr_add_0__13, d_arr_add_0__12, d_arr_add_0__11, 
         d_arr_add_0__10, d_arr_add_0__9, d_arr_add_0__8, d_arr_add_0__7, 
         d_arr_add_0__6, d_arr_add_0__5, d_arr_add_0__4, d_arr_add_0__3, 
         d_arr_add_0__2, d_arr_add_0__1, d_arr_add_0__0, d_arr_add_1__31, 
         d_arr_add_1__30, d_arr_add_1__29, d_arr_add_1__28, d_arr_add_1__27, 
         d_arr_add_1__26, d_arr_add_1__25, d_arr_add_1__24, d_arr_add_1__23, 
         d_arr_add_1__22, d_arr_add_1__21, d_arr_add_1__20, d_arr_add_1__19, 
         d_arr_add_1__18, d_arr_add_1__17, d_arr_add_1__16, d_arr_add_1__15, 
         d_arr_add_1__14, d_arr_add_1__13, d_arr_add_1__12, d_arr_add_1__11, 
         d_arr_add_1__10, d_arr_add_1__9, d_arr_add_1__8, d_arr_add_1__7, 
         d_arr_add_1__6, d_arr_add_1__5, d_arr_add_1__4, d_arr_add_1__3, 
         d_arr_add_1__2, d_arr_add_1__1, d_arr_add_1__0, d_arr_add_2__31, 
         d_arr_add_2__30, d_arr_add_2__29, d_arr_add_2__28, d_arr_add_2__27, 
         d_arr_add_2__26, d_arr_add_2__25, d_arr_add_2__24, d_arr_add_2__23, 
         d_arr_add_2__22, d_arr_add_2__21, d_arr_add_2__20, d_arr_add_2__19, 
         d_arr_add_2__18, d_arr_add_2__17, d_arr_add_2__16, d_arr_add_2__15, 
         d_arr_add_2__14, d_arr_add_2__13, d_arr_add_2__12, d_arr_add_2__11, 
         d_arr_add_2__10, d_arr_add_2__9, d_arr_add_2__8, d_arr_add_2__7, 
         d_arr_add_2__6, d_arr_add_2__5, d_arr_add_2__4, d_arr_add_2__3, 
         d_arr_add_2__2, d_arr_add_2__1, d_arr_add_2__0, d_arr_add_3__31, 
         d_arr_add_3__30, d_arr_add_3__29, d_arr_add_3__28, d_arr_add_3__27, 
         d_arr_add_3__26, d_arr_add_3__25, d_arr_add_3__24, d_arr_add_3__23, 
         d_arr_add_3__22, d_arr_add_3__21, d_arr_add_3__20, d_arr_add_3__19, 
         d_arr_add_3__18, d_arr_add_3__17, d_arr_add_3__16, d_arr_add_3__15, 
         d_arr_add_3__14, d_arr_add_3__13, d_arr_add_3__12, d_arr_add_3__11, 
         d_arr_add_3__10, d_arr_add_3__9, d_arr_add_3__8, d_arr_add_3__7, 
         d_arr_add_3__6, d_arr_add_3__5, d_arr_add_3__4, d_arr_add_3__3, 
         d_arr_add_3__2, d_arr_add_3__1, d_arr_add_3__0, d_arr_add_9__31, 
         d_arr_add_9__30, d_arr_add_9__29, d_arr_add_9__28, d_arr_add_9__27, 
         d_arr_add_9__26, d_arr_add_9__25, d_arr_add_9__24, d_arr_add_9__23, 
         d_arr_add_9__22, d_arr_add_9__21, d_arr_add_9__20, d_arr_add_9__19, 
         d_arr_add_9__18, d_arr_add_9__17, d_arr_add_9__16, d_arr_add_9__15, 
         d_arr_add_9__14, d_arr_add_9__13, d_arr_add_9__12, d_arr_add_9__11, 
         d_arr_add_9__10, d_arr_add_9__9, d_arr_add_9__8, d_arr_add_9__7, 
         d_arr_add_9__6, d_arr_add_9__5, d_arr_add_9__4, d_arr_add_9__3, 
         d_arr_add_9__2, d_arr_add_9__1, d_arr_add_9__0, d_arr_add_10__31, 
         d_arr_add_10__30, d_arr_add_10__29, d_arr_add_10__28, d_arr_add_10__27, 
         d_arr_add_10__26, d_arr_add_10__25, d_arr_add_10__24, d_arr_add_10__23, 
         d_arr_add_10__22, d_arr_add_10__21, d_arr_add_10__20, d_arr_add_10__19, 
         d_arr_add_10__18, d_arr_add_10__17, d_arr_add_10__16, d_arr_add_10__15, 
         d_arr_add_10__14, d_arr_add_10__13, d_arr_add_10__12, d_arr_add_10__11, 
         d_arr_add_10__10, d_arr_add_10__9, d_arr_add_10__8, d_arr_add_10__7, 
         d_arr_add_10__6, d_arr_add_10__5, d_arr_add_10__4, d_arr_add_10__3, 
         d_arr_add_10__2, d_arr_add_10__1, d_arr_add_10__0, d_arr_add_11__31, 
         d_arr_add_11__30, d_arr_add_11__29, d_arr_add_11__28, d_arr_add_11__27, 
         d_arr_add_11__26, d_arr_add_11__25, d_arr_add_11__24, d_arr_add_11__23, 
         d_arr_add_11__22, d_arr_add_11__21, d_arr_add_11__20, d_arr_add_11__19, 
         d_arr_add_11__18, d_arr_add_11__17, d_arr_add_11__16, d_arr_add_11__15, 
         d_arr_add_11__14, d_arr_add_11__13, d_arr_add_11__12, d_arr_add_11__11, 
         d_arr_add_11__10, d_arr_add_11__9, d_arr_add_11__8, d_arr_add_11__7, 
         d_arr_add_11__6, d_arr_add_11__5, d_arr_add_11__4, d_arr_add_11__3, 
         d_arr_add_11__2, d_arr_add_11__1, d_arr_add_11__0, d_arr_add_12__31, 
         d_arr_add_12__30, d_arr_add_12__29, d_arr_add_12__28, d_arr_add_12__27, 
         d_arr_add_12__26, d_arr_add_12__25, d_arr_add_12__24, d_arr_add_12__23, 
         d_arr_add_12__22, d_arr_add_12__21, d_arr_add_12__20, d_arr_add_12__19, 
         d_arr_add_12__18, d_arr_add_12__17, d_arr_add_12__16, d_arr_add_12__15, 
         d_arr_add_12__14, d_arr_add_12__13, d_arr_add_12__12, d_arr_add_12__11, 
         d_arr_add_12__10, d_arr_add_12__9, d_arr_add_12__8, d_arr_add_12__7, 
         d_arr_add_12__6, d_arr_add_12__5, d_arr_add_12__4, d_arr_add_12__3, 
         d_arr_add_12__2, d_arr_add_12__1, d_arr_add_12__0, d_arr_add_18__31, 
         d_arr_add_18__30, d_arr_add_18__29, d_arr_add_18__28, d_arr_add_18__27, 
         d_arr_add_18__26, d_arr_add_18__25, d_arr_add_18__24, d_arr_add_18__23, 
         d_arr_add_18__22, d_arr_add_18__21, d_arr_add_18__20, d_arr_add_18__19, 
         d_arr_add_18__18, d_arr_add_18__17, d_arr_add_18__16, d_arr_add_18__15, 
         d_arr_add_18__14, d_arr_add_18__13, d_arr_add_18__12, d_arr_add_18__11, 
         d_arr_add_18__10, d_arr_add_18__9, d_arr_add_18__8, d_arr_add_18__7, 
         d_arr_add_18__6, d_arr_add_18__5, d_arr_add_18__4, d_arr_add_18__3, 
         d_arr_add_18__2, d_arr_add_18__1, d_arr_add_18__0, d_arr_add_19__31, 
         d_arr_add_19__30, d_arr_add_19__29, d_arr_add_19__28, d_arr_add_19__27, 
         d_arr_add_19__26, d_arr_add_19__25, d_arr_add_19__24, d_arr_add_19__23, 
         d_arr_add_19__22, d_arr_add_19__21, d_arr_add_19__20, d_arr_add_19__19, 
         d_arr_add_19__18, d_arr_add_19__17, d_arr_add_19__16, d_arr_add_19__15, 
         d_arr_add_19__14, d_arr_add_19__13, d_arr_add_19__12, d_arr_add_19__11, 
         d_arr_add_19__10, d_arr_add_19__9, d_arr_add_19__8, d_arr_add_19__7, 
         d_arr_add_19__6, d_arr_add_19__5, d_arr_add_19__4, d_arr_add_19__3, 
         d_arr_add_19__2, d_arr_add_19__1, d_arr_add_19__0, d_arr_add_20__31, 
         d_arr_add_20__30, d_arr_add_20__29, d_arr_add_20__28, d_arr_add_20__27, 
         d_arr_add_20__26, d_arr_add_20__25, d_arr_add_20__24, d_arr_add_20__23, 
         d_arr_add_20__22, d_arr_add_20__21, d_arr_add_20__20, d_arr_add_20__19, 
         d_arr_add_20__18, d_arr_add_20__17, d_arr_add_20__16, d_arr_add_20__15, 
         d_arr_add_20__14, d_arr_add_20__13, d_arr_add_20__12, d_arr_add_20__11, 
         d_arr_add_20__10, d_arr_add_20__9, d_arr_add_20__8, d_arr_add_20__7, 
         d_arr_add_20__6, d_arr_add_20__5, d_arr_add_20__4, d_arr_add_20__3, 
         d_arr_add_20__2, d_arr_add_20__1, d_arr_add_20__0, d_arr_merge1_0__31, 
         d_arr_merge1_0__30, d_arr_merge1_0__29, d_arr_merge1_0__28, 
         d_arr_merge1_0__27, d_arr_merge1_0__26, d_arr_merge1_0__25, 
         d_arr_merge1_0__24, d_arr_merge1_0__23, d_arr_merge1_0__22, 
         d_arr_merge1_0__21, d_arr_merge1_0__20, d_arr_merge1_0__19, 
         d_arr_merge1_0__18, d_arr_merge1_0__17, d_arr_merge1_0__16, 
         d_arr_merge1_0__15, d_arr_merge1_0__14, d_arr_merge1_0__13, 
         d_arr_merge1_0__12, d_arr_merge1_0__11, d_arr_merge1_0__10, 
         d_arr_merge1_0__9, d_arr_merge1_0__8, d_arr_merge1_0__7, 
         d_arr_merge1_0__6, d_arr_merge1_0__5, d_arr_merge1_0__4, 
         d_arr_merge1_0__3, d_arr_merge1_0__2, d_arr_merge1_0__1, 
         d_arr_merge1_0__0, d_arr_merge1_1__31, d_arr_merge1_1__30, 
         d_arr_merge1_1__29, d_arr_merge1_1__28, d_arr_merge1_1__27, 
         d_arr_merge1_1__26, d_arr_merge1_1__25, d_arr_merge1_1__24, 
         d_arr_merge1_1__23, d_arr_merge1_1__22, d_arr_merge1_1__21, 
         d_arr_merge1_1__20, d_arr_merge1_1__19, d_arr_merge1_1__18, 
         d_arr_merge1_1__17, d_arr_merge1_1__16, d_arr_merge1_1__15, 
         d_arr_merge1_1__14, d_arr_merge1_1__13, d_arr_merge1_1__12, 
         d_arr_merge1_1__11, d_arr_merge1_1__10, d_arr_merge1_1__9, 
         d_arr_merge1_1__8, d_arr_merge1_1__7, d_arr_merge1_1__6, 
         d_arr_merge1_1__5, d_arr_merge1_1__4, d_arr_merge1_1__3, 
         d_arr_merge1_1__2, d_arr_merge1_1__1, d_arr_merge1_1__0, 
         d_arr_merge2_0__31, d_arr_merge2_0__26, d_arr_merge2_0__25, 
         d_arr_merge2_0__24, d_arr_merge2_0__23, d_arr_merge2_0__22, 
         d_arr_merge2_0__21, d_arr_merge2_0__20, d_arr_merge2_0__19, 
         d_arr_merge2_0__18, d_arr_merge2_0__17, d_arr_merge2_0__16, 
         d_arr_merge2_0__15, d_arr_merge2_0__14, d_arr_merge2_0__13, 
         d_arr_merge2_0__12, d_arr_merge2_0__11, d_arr_merge2_0__10, 
         d_arr_merge2_0__9, d_arr_merge2_0__8, d_arr_merge2_0__7, 
         d_arr_merge2_0__6, d_arr_merge2_0__5, d_arr_merge2_0__4, 
         d_arr_merge2_0__3, d_arr_merge2_0__2, d_arr_merge2_0__1, 
         d_arr_merge2_0__0, d_arr_merge2_1__31, d_arr_merge2_1__26, 
         d_arr_merge2_1__25, d_arr_merge2_1__24, d_arr_merge2_1__23, 
         d_arr_merge2_1__22, d_arr_merge2_1__21, d_arr_merge2_1__20, 
         d_arr_merge2_1__19, d_arr_merge2_1__18, d_arr_merge2_1__17, 
         d_arr_merge2_1__16, d_arr_merge2_1__15, d_arr_merge2_1__14, 
         d_arr_merge2_1__13, d_arr_merge2_1__12, d_arr_merge2_1__11, 
         d_arr_merge2_1__10, d_arr_merge2_1__9, d_arr_merge2_1__8, 
         d_arr_merge2_1__7, d_arr_merge2_1__6, d_arr_merge2_1__5, 
         d_arr_merge2_1__4, d_arr_merge2_1__3, d_arr_merge2_1__2, 
         d_arr_merge2_1__1, d_arr_merge2_1__0, d_arr_relu_0__31, 
         d_arr_relu_0__30, d_arr_relu_0__29, d_arr_relu_0__28, d_arr_relu_0__27, 
         d_arr_relu_0__26, d_arr_relu_0__25, d_arr_relu_0__24, d_arr_relu_0__23, 
         d_arr_relu_0__22, d_arr_relu_0__21, d_arr_relu_0__20, d_arr_relu_0__19, 
         d_arr_relu_0__18, d_arr_relu_0__17, d_arr_relu_0__16, d_arr_relu_0__14, 
         d_arr_relu_0__13, d_arr_relu_0__12, d_arr_relu_0__11, d_arr_relu_0__10, 
         d_arr_relu_0__9, d_arr_relu_0__8, d_arr_relu_0__7, d_arr_relu_0__6, 
         d_arr_relu_0__5, d_arr_relu_0__4, d_arr_relu_0__3, d_arr_relu_0__2, 
         d_arr_relu_0__1, d_arr_relu_0__0, d_arr_relu_1__31, d_arr_relu_1__30, 
         d_arr_relu_1__29, d_arr_relu_1__28, d_arr_relu_1__27, d_arr_relu_1__26, 
         d_arr_relu_1__25, d_arr_relu_1__24, d_arr_relu_1__23, d_arr_relu_1__22, 
         d_arr_relu_1__21, d_arr_relu_1__20, d_arr_relu_1__19, d_arr_relu_1__18, 
         d_arr_relu_1__17, d_arr_relu_1__16, d_arr_relu_1__14, d_arr_relu_1__13, 
         d_arr_relu_1__12, d_arr_relu_1__11, d_arr_relu_1__10, d_arr_relu_1__9, 
         d_arr_relu_1__8, d_arr_relu_1__7, d_arr_relu_1__6, d_arr_relu_1__5, 
         d_arr_relu_1__4, d_arr_relu_1__3, d_arr_relu_1__2, d_arr_relu_1__1, 
         d_arr_relu_1__0, sel_mul, sel_add, GND0, counter_12, counter_11, 
         counter_10, counter_9, counter_7, counter_6, counter_5, counter_4, 
         counter_3, counter_2, counter_1, nx20, nx92, nx194, nx16101, nx16115, 
         nx16125, nx16135, nx16145, nx16155, nx16165, nx16175, nx16185, nx16195, 
         nx16205, nx16215, nx16225, nx16235, nx16245, nx16255, nx16265, nx16276, 
         nx16278, nx16281, nx16285, nx16289, nx16293, nx16295, nx16299, nx16301, 
         nx16306, nx16309, nx16313, nx16315, nx16319, nx16321, nx16325, nx16327, 
         nx16331, nx16333, nx16337, nx16339, nx16343, nx16345, nx16349, nx16351, 
         nx16353, nx16361, nx16363, nx16366, nx16371, nx16373, nx16375, nx16380, 
         nx16382, nx16386, nx16388, nx16390, nx16399, nx16401, nx16403, nx16405, 
         nx16407, nx16409, nx16411, nx16413, nx16415, nx16417, nx16419, nx16421, 
         nx16423, nx16425, nx16427, nx16429, nx16431, nx16433, nx16435, nx16437, 
         nx16439, nx16441, nx16443, nx16445, nx16447, nx16449, nx16451, nx16453, 
         nx16455, nx16457, nx16459, nx16461, nx16463, nx16465, nx16467, nx16469, 
         nx16471, nx16473, nx16475, nx16477, nx16479, nx16481, nx16483, nx16485, 
         nx16487, nx16489, nx16491, nx16497, nx16499, nx16501, nx16503, nx16505, 
         nx16507, nx16509, nx16511, nx16513, nx16515, nx16517, nx16519, nx16521, 
         nx16523, nx16525, nx16527, nx16529, nx16531, nx16533, nx16535, nx16537, 
         nx16539, nx16541, nx16543, nx16545, nx16547, nx16549, nx16551, nx16553, 
         nx16555, nx16557, nx16559, nx16561, nx16563, nx16565, nx16567, nx16569, 
         nx16571, nx16573, nx16575, nx16577, nx16579, nx16581, nx16583, nx16585, 
         nx16587, nx16589, nx16591, nx16593, nx16595, nx16597, nx16599, nx16601, 
         nx16603, nx16605, nx16607, nx16609, nx16611, nx16613, nx16615, nx16617, 
         nx16619, nx16621, nx16623, nx16625, nx16627, nx16629, nx16631, nx16633, 
         nx16635, nx16637, nx16639, nx16641, nx16643, nx16645, nx16651, nx16653, 
         nx16659, nx16661, nx16663, nx16665, nx16667, nx19388, nx19390, nx19396, 
         nx19398, nx19400, nx19402, nx19404, nx19406, nx19408, nx19410, nx19412, 
         nx19414, nx19416, nx19418, nx19420, nx19422, nx19424, nx19426, nx19428, 
         nx19430, nx19432, nx19434, nx19436, nx19438, nx19440, nx19442, nx19444, 
         nx19446, nx19448, nx19450, nx19452, nx19454, nx19456, nx19458, nx19460, 
         nx19462, nx19464, nx19466, nx19468, nx19470, nx19472, nx19474, nx19476, 
         nx19478, nx19480, nx19482, nx19484, nx19486, nx19488, nx19490, nx19492, 
         nx19494;
    wire [2714:0] \$dummy ;




    CacheMuxer cache_muxer_gen (.d_arr_mux_0__31 (img_data_0__15), .d_arr_mux_0__30 (
               GND0), .d_arr_mux_0__29 (GND0), .d_arr_mux_0__28 (GND0), .d_arr_mux_0__27 (
               GND0), .d_arr_mux_0__26 (GND0), .d_arr_mux_0__25 (GND0), .d_arr_mux_0__24 (
               GND0), .d_arr_mux_0__23 (GND0), .d_arr_mux_0__22 (GND0), .d_arr_mux_0__21 (
               GND0), .d_arr_mux_0__20 (GND0), .d_arr_mux_0__19 (GND0), .d_arr_mux_0__18 (
               GND0), .d_arr_mux_0__17 (GND0), .d_arr_mux_0__16 (GND0), .d_arr_mux_0__15 (
               GND0), .d_arr_mux_0__14 (nx19396), .d_arr_mux_0__13 (
               img_data_0__13), .d_arr_mux_0__12 (img_data_0__12), .d_arr_mux_0__11 (
               img_data_0__11), .d_arr_mux_0__10 (img_data_0__10), .d_arr_mux_0__9 (
               img_data_0__9), .d_arr_mux_0__8 (img_data_0__8), .d_arr_mux_0__7 (
               img_data_0__7), .d_arr_mux_0__6 (img_data_0__6), .d_arr_mux_0__5 (
               img_data_0__5), .d_arr_mux_0__4 (img_data_0__4), .d_arr_mux_0__3 (
               img_data_0__3), .d_arr_mux_0__2 (img_data_0__2), .d_arr_mux_0__1 (
               img_data_0__1), .d_arr_mux_0__0 (img_data_0__0), .d_arr_mux_1__31 (
               img_data_1__15), .d_arr_mux_1__30 (GND0), .d_arr_mux_1__29 (GND0)
               , .d_arr_mux_1__28 (GND0), .d_arr_mux_1__27 (GND0), .d_arr_mux_1__26 (
               GND0), .d_arr_mux_1__25 (GND0), .d_arr_mux_1__24 (GND0), .d_arr_mux_1__23 (
               GND0), .d_arr_mux_1__22 (GND0), .d_arr_mux_1__21 (GND0), .d_arr_mux_1__20 (
               GND0), .d_arr_mux_1__19 (GND0), .d_arr_mux_1__18 (GND0), .d_arr_mux_1__17 (
               GND0), .d_arr_mux_1__16 (GND0), .d_arr_mux_1__15 (GND0), .d_arr_mux_1__14 (
               nx19398), .d_arr_mux_1__13 (img_data_1__13), .d_arr_mux_1__12 (
               img_data_1__12), .d_arr_mux_1__11 (img_data_1__11), .d_arr_mux_1__10 (
               nx19402), .d_arr_mux_1__9 (img_data_1__9), .d_arr_mux_1__8 (
               img_data_1__8), .d_arr_mux_1__7 (img_data_1__7), .d_arr_mux_1__6 (
               img_data_1__6), .d_arr_mux_1__5 (img_data_1__5), .d_arr_mux_1__4 (
               img_data_1__4), .d_arr_mux_1__3 (img_data_1__3), .d_arr_mux_1__2 (
               img_data_1__2), .d_arr_mux_1__1 (img_data_1__1), .d_arr_mux_1__0 (
               img_data_1__0), .d_arr_mux_2__31 (img_data_2__15), .d_arr_mux_2__30 (
               GND0), .d_arr_mux_2__29 (GND0), .d_arr_mux_2__28 (GND0), .d_arr_mux_2__27 (
               GND0), .d_arr_mux_2__26 (GND0), .d_arr_mux_2__25 (GND0), .d_arr_mux_2__24 (
               GND0), .d_arr_mux_2__23 (GND0), .d_arr_mux_2__22 (GND0), .d_arr_mux_2__21 (
               GND0), .d_arr_mux_2__20 (GND0), .d_arr_mux_2__19 (GND0), .d_arr_mux_2__18 (
               GND0), .d_arr_mux_2__17 (GND0), .d_arr_mux_2__16 (GND0), .d_arr_mux_2__15 (
               GND0), .d_arr_mux_2__14 (nx19404), .d_arr_mux_2__13 (
               img_data_2__13), .d_arr_mux_2__12 (img_data_2__12), .d_arr_mux_2__11 (
               img_data_2__11), .d_arr_mux_2__10 (nx19408), .d_arr_mux_2__9 (
               img_data_2__9), .d_arr_mux_2__8 (img_data_2__8), .d_arr_mux_2__7 (
               img_data_2__7), .d_arr_mux_2__6 (img_data_2__6), .d_arr_mux_2__5 (
               img_data_2__5), .d_arr_mux_2__4 (img_data_2__4), .d_arr_mux_2__3 (
               img_data_2__3), .d_arr_mux_2__2 (img_data_2__2), .d_arr_mux_2__1 (
               img_data_2__1), .d_arr_mux_2__0 (img_data_2__0), .d_arr_mux_3__31 (
               img_data_5__15), .d_arr_mux_3__30 (GND0), .d_arr_mux_3__29 (GND0)
               , .d_arr_mux_3__28 (GND0), .d_arr_mux_3__27 (GND0), .d_arr_mux_3__26 (
               GND0), .d_arr_mux_3__25 (GND0), .d_arr_mux_3__24 (GND0), .d_arr_mux_3__23 (
               GND0), .d_arr_mux_3__22 (GND0), .d_arr_mux_3__21 (GND0), .d_arr_mux_3__20 (
               GND0), .d_arr_mux_3__19 (GND0), .d_arr_mux_3__18 (GND0), .d_arr_mux_3__17 (
               GND0), .d_arr_mux_3__16 (GND0), .d_arr_mux_3__15 (GND0), .d_arr_mux_3__14 (
               nx19410), .d_arr_mux_3__13 (img_data_5__13), .d_arr_mux_3__12 (
               img_data_5__12), .d_arr_mux_3__11 (img_data_5__11), .d_arr_mux_3__10 (
               img_data_5__10), .d_arr_mux_3__9 (img_data_5__9), .d_arr_mux_3__8 (
               img_data_5__8), .d_arr_mux_3__7 (img_data_5__7), .d_arr_mux_3__6 (
               img_data_5__6), .d_arr_mux_3__5 (img_data_5__5), .d_arr_mux_3__4 (
               img_data_5__4), .d_arr_mux_3__3 (img_data_5__3), .d_arr_mux_3__2 (
               img_data_5__2), .d_arr_mux_3__1 (img_data_5__1), .d_arr_mux_3__0 (
               img_data_5__0), .d_arr_mux_4__31 (img_data_6__15), .d_arr_mux_4__30 (
               GND0), .d_arr_mux_4__29 (GND0), .d_arr_mux_4__28 (GND0), .d_arr_mux_4__27 (
               GND0), .d_arr_mux_4__26 (GND0), .d_arr_mux_4__25 (GND0), .d_arr_mux_4__24 (
               GND0), .d_arr_mux_4__23 (GND0), .d_arr_mux_4__22 (GND0), .d_arr_mux_4__21 (
               GND0), .d_arr_mux_4__20 (GND0), .d_arr_mux_4__19 (GND0), .d_arr_mux_4__18 (
               GND0), .d_arr_mux_4__17 (GND0), .d_arr_mux_4__16 (GND0), .d_arr_mux_4__15 (
               GND0), .d_arr_mux_4__14 (nx19412), .d_arr_mux_4__13 (
               img_data_6__13), .d_arr_mux_4__12 (img_data_6__12), .d_arr_mux_4__11 (
               img_data_6__11), .d_arr_mux_4__10 (nx19416), .d_arr_mux_4__9 (
               img_data_6__9), .d_arr_mux_4__8 (img_data_6__8), .d_arr_mux_4__7 (
               img_data_6__7), .d_arr_mux_4__6 (img_data_6__6), .d_arr_mux_4__5 (
               img_data_6__5), .d_arr_mux_4__4 (img_data_6__4), .d_arr_mux_4__3 (
               img_data_6__3), .d_arr_mux_4__2 (img_data_6__2), .d_arr_mux_4__1 (
               img_data_6__1), .d_arr_mux_4__0 (img_data_6__0), .d_arr_mux_5__31 (
               nx16659), .d_arr_mux_5__30 (GND0), .d_arr_mux_5__29 (GND0), .d_arr_mux_5__28 (
               GND0), .d_arr_mux_5__27 (GND0), .d_arr_mux_5__26 (GND0), .d_arr_mux_5__25 (
               GND0), .d_arr_mux_5__24 (GND0), .d_arr_mux_5__23 (GND0), .d_arr_mux_5__22 (
               GND0), .d_arr_mux_5__21 (GND0), .d_arr_mux_5__20 (GND0), .d_arr_mux_5__19 (
               GND0), .d_arr_mux_5__18 (GND0), .d_arr_mux_5__17 (GND0), .d_arr_mux_5__16 (
               GND0), .d_arr_mux_5__15 (GND0), .d_arr_mux_5__14 (nx19418), .d_arr_mux_5__13 (
               img_data_7__13), .d_arr_mux_5__12 (img_data_7__12), .d_arr_mux_5__11 (
               img_data_7__11), .d_arr_mux_5__10 (nx19422), .d_arr_mux_5__9 (
               img_data_7__9), .d_arr_mux_5__8 (img_data_7__8), .d_arr_mux_5__7 (
               img_data_7__7), .d_arr_mux_5__6 (img_data_7__6), .d_arr_mux_5__5 (
               img_data_7__5), .d_arr_mux_5__4 (img_data_7__4), .d_arr_mux_5__3 (
               img_data_7__3), .d_arr_mux_5__2 (img_data_7__2), .d_arr_mux_5__1 (
               img_data_7__1), .d_arr_mux_5__0 (img_data_7__0), .d_arr_mux_6__31 (
               img_data_10__15), .d_arr_mux_6__30 (GND0), .d_arr_mux_6__29 (GND0
               ), .d_arr_mux_6__28 (GND0), .d_arr_mux_6__27 (GND0), .d_arr_mux_6__26 (
               GND0), .d_arr_mux_6__25 (GND0), .d_arr_mux_6__24 (GND0), .d_arr_mux_6__23 (
               GND0), .d_arr_mux_6__22 (GND0), .d_arr_mux_6__21 (GND0), .d_arr_mux_6__20 (
               GND0), .d_arr_mux_6__19 (GND0), .d_arr_mux_6__18 (GND0), .d_arr_mux_6__17 (
               GND0), .d_arr_mux_6__16 (GND0), .d_arr_mux_6__15 (GND0), .d_arr_mux_6__14 (
               nx19424), .d_arr_mux_6__13 (img_data_10__13), .d_arr_mux_6__12 (
               img_data_10__12), .d_arr_mux_6__11 (img_data_10__11), .d_arr_mux_6__10 (
               img_data_10__10), .d_arr_mux_6__9 (img_data_10__9), .d_arr_mux_6__8 (
               img_data_10__8), .d_arr_mux_6__7 (img_data_10__7), .d_arr_mux_6__6 (
               img_data_10__6), .d_arr_mux_6__5 (img_data_10__5), .d_arr_mux_6__4 (
               img_data_10__4), .d_arr_mux_6__3 (img_data_10__3), .d_arr_mux_6__2 (
               img_data_10__2), .d_arr_mux_6__1 (img_data_10__1), .d_arr_mux_6__0 (
               img_data_10__0), .d_arr_mux_7__31 (nx16661), .d_arr_mux_7__30 (
               GND0), .d_arr_mux_7__29 (GND0), .d_arr_mux_7__28 (GND0), .d_arr_mux_7__27 (
               GND0), .d_arr_mux_7__26 (GND0), .d_arr_mux_7__25 (GND0), .d_arr_mux_7__24 (
               GND0), .d_arr_mux_7__23 (GND0), .d_arr_mux_7__22 (GND0), .d_arr_mux_7__21 (
               GND0), .d_arr_mux_7__20 (GND0), .d_arr_mux_7__19 (GND0), .d_arr_mux_7__18 (
               GND0), .d_arr_mux_7__17 (GND0), .d_arr_mux_7__16 (GND0), .d_arr_mux_7__15 (
               GND0), .d_arr_mux_7__14 (nx19426), .d_arr_mux_7__13 (
               img_data_11__13), .d_arr_mux_7__12 (img_data_11__12), .d_arr_mux_7__11 (
               img_data_11__11), .d_arr_mux_7__10 (nx19430), .d_arr_mux_7__9 (
               img_data_11__9), .d_arr_mux_7__8 (img_data_11__8), .d_arr_mux_7__7 (
               img_data_11__7), .d_arr_mux_7__6 (img_data_11__6), .d_arr_mux_7__5 (
               img_data_11__5), .d_arr_mux_7__4 (img_data_11__4), .d_arr_mux_7__3 (
               img_data_11__3), .d_arr_mux_7__2 (img_data_11__2), .d_arr_mux_7__1 (
               img_data_11__1), .d_arr_mux_7__0 (img_data_11__0), .d_arr_mux_8__31 (
               nx16663), .d_arr_mux_8__30 (GND0), .d_arr_mux_8__29 (GND0), .d_arr_mux_8__28 (
               GND0), .d_arr_mux_8__27 (GND0), .d_arr_mux_8__26 (GND0), .d_arr_mux_8__25 (
               GND0), .d_arr_mux_8__24 (GND0), .d_arr_mux_8__23 (GND0), .d_arr_mux_8__22 (
               GND0), .d_arr_mux_8__21 (GND0), .d_arr_mux_8__20 (GND0), .d_arr_mux_8__19 (
               GND0), .d_arr_mux_8__18 (GND0), .d_arr_mux_8__17 (GND0), .d_arr_mux_8__16 (
               GND0), .d_arr_mux_8__15 (GND0), .d_arr_mux_8__14 (nx19432), .d_arr_mux_8__13 (
               img_data_12__13), .d_arr_mux_8__12 (img_data_12__12), .d_arr_mux_8__11 (
               img_data_12__11), .d_arr_mux_8__10 (nx19436), .d_arr_mux_8__9 (
               img_data_12__9), .d_arr_mux_8__8 (img_data_12__8), .d_arr_mux_8__7 (
               img_data_12__7), .d_arr_mux_8__6 (img_data_12__6), .d_arr_mux_8__5 (
               img_data_12__5), .d_arr_mux_8__4 (img_data_12__4), .d_arr_mux_8__3 (
               img_data_12__3), .d_arr_mux_8__2 (img_data_12__2), .d_arr_mux_8__1 (
               img_data_12__1), .d_arr_mux_8__0 (img_data_12__0), .d_arr_mux_9__31 (
               nx16401), .d_arr_mux_9__30 (nx16401), .d_arr_mux_9__29 (nx16401)
               , .d_arr_mux_9__28 (nx16401), .d_arr_mux_9__27 (nx16401), .d_arr_mux_9__26 (
               nx16401), .d_arr_mux_9__25 (nx16401), .d_arr_mux_9__24 (nx16403)
               , .d_arr_mux_9__23 (nx16403), .d_arr_mux_9__22 (nx16403), .d_arr_mux_9__21 (
               nx16403), .d_arr_mux_9__20 (nx16403), .d_arr_mux_9__19 (nx16403)
               , .d_arr_mux_9__18 (nx16403), .d_arr_mux_9__17 (nx16405), .d_arr_mux_9__16 (
               nx16405), .d_arr_mux_9__15 (nx16405), .d_arr_mux_9__14 (
               ordered_img_data_9__14), .d_arr_mux_9__13 (ordered_img_data_9__13
               ), .d_arr_mux_9__12 (ordered_img_data_9__12), .d_arr_mux_9__11 (
               ordered_img_data_9__11), .d_arr_mux_9__10 (ordered_img_data_9__10
               ), .d_arr_mux_9__9 (ordered_img_data_9__9), .d_arr_mux_9__8 (
               ordered_img_data_9__8), .d_arr_mux_9__7 (ordered_img_data_9__7), 
               .d_arr_mux_9__6 (ordered_img_data_9__6), .d_arr_mux_9__5 (
               ordered_img_data_9__5), .d_arr_mux_9__4 (ordered_img_data_9__4), 
               .d_arr_mux_9__3 (ordered_img_data_9__3), .d_arr_mux_9__2 (
               ordered_img_data_9__2), .d_arr_mux_9__1 (ordered_img_data_9__1), 
               .d_arr_mux_9__0 (ordered_img_data_9__0), .d_arr_mux_10__31 (
               nx16409), .d_arr_mux_10__30 (nx16409), .d_arr_mux_10__29 (nx16409
               ), .d_arr_mux_10__28 (nx16409), .d_arr_mux_10__27 (nx16409), .d_arr_mux_10__26 (
               nx16409), .d_arr_mux_10__25 (nx16409), .d_arr_mux_10__24 (nx16411
               ), .d_arr_mux_10__23 (nx16411), .d_arr_mux_10__22 (nx16411), .d_arr_mux_10__21 (
               nx16411), .d_arr_mux_10__20 (nx16411), .d_arr_mux_10__19 (nx16411
               ), .d_arr_mux_10__18 (nx16411), .d_arr_mux_10__17 (nx16413), .d_arr_mux_10__16 (
               nx16413), .d_arr_mux_10__15 (nx16413), .d_arr_mux_10__14 (
               ordered_img_data_10__14), .d_arr_mux_10__13 (
               ordered_img_data_10__13), .d_arr_mux_10__12 (
               ordered_img_data_10__12), .d_arr_mux_10__11 (
               ordered_img_data_10__11), .d_arr_mux_10__10 (
               ordered_img_data_10__10), .d_arr_mux_10__9 (
               ordered_img_data_10__9), .d_arr_mux_10__8 (ordered_img_data_10__8
               ), .d_arr_mux_10__7 (ordered_img_data_10__7), .d_arr_mux_10__6 (
               ordered_img_data_10__6), .d_arr_mux_10__5 (ordered_img_data_10__5
               ), .d_arr_mux_10__4 (ordered_img_data_10__4), .d_arr_mux_10__3 (
               ordered_img_data_10__3), .d_arr_mux_10__2 (ordered_img_data_10__2
               ), .d_arr_mux_10__1 (ordered_img_data_10__1), .d_arr_mux_10__0 (
               ordered_img_data_10__0), .d_arr_mux_11__31 (nx16417), .d_arr_mux_11__30 (
               nx16417), .d_arr_mux_11__29 (nx16417), .d_arr_mux_11__28 (nx16417
               ), .d_arr_mux_11__27 (nx16417), .d_arr_mux_11__26 (nx16417), .d_arr_mux_11__25 (
               nx16417), .d_arr_mux_11__24 (nx16419), .d_arr_mux_11__23 (nx16419
               ), .d_arr_mux_11__22 (nx16419), .d_arr_mux_11__21 (nx16419), .d_arr_mux_11__20 (
               nx16419), .d_arr_mux_11__19 (nx16419), .d_arr_mux_11__18 (nx16419
               ), .d_arr_mux_11__17 (nx16421), .d_arr_mux_11__16 (nx16421), .d_arr_mux_11__15 (
               nx16421), .d_arr_mux_11__14 (ordered_img_data_11__14), .d_arr_mux_11__13 (
               ordered_img_data_11__13), .d_arr_mux_11__12 (
               ordered_img_data_11__12), .d_arr_mux_11__11 (
               ordered_img_data_11__11), .d_arr_mux_11__10 (
               ordered_img_data_11__10), .d_arr_mux_11__9 (
               ordered_img_data_11__9), .d_arr_mux_11__8 (ordered_img_data_11__8
               ), .d_arr_mux_11__7 (ordered_img_data_11__7), .d_arr_mux_11__6 (
               ordered_img_data_11__6), .d_arr_mux_11__5 (ordered_img_data_11__5
               ), .d_arr_mux_11__4 (ordered_img_data_11__4), .d_arr_mux_11__3 (
               ordered_img_data_11__3), .d_arr_mux_11__2 (ordered_img_data_11__2
               ), .d_arr_mux_11__1 (ordered_img_data_11__1), .d_arr_mux_11__0 (
               ordered_img_data_11__0), .d_arr_mux_12__31 (nx16425), .d_arr_mux_12__30 (
               nx16425), .d_arr_mux_12__29 (nx16425), .d_arr_mux_12__28 (nx16425
               ), .d_arr_mux_12__27 (nx16425), .d_arr_mux_12__26 (nx16425), .d_arr_mux_12__25 (
               nx16425), .d_arr_mux_12__24 (nx16427), .d_arr_mux_12__23 (nx16427
               ), .d_arr_mux_12__22 (nx16427), .d_arr_mux_12__21 (nx16427), .d_arr_mux_12__20 (
               nx16427), .d_arr_mux_12__19 (nx16427), .d_arr_mux_12__18 (nx16427
               ), .d_arr_mux_12__17 (nx16429), .d_arr_mux_12__16 (nx16429), .d_arr_mux_12__15 (
               nx16429), .d_arr_mux_12__14 (ordered_img_data_12__14), .d_arr_mux_12__13 (
               ordered_img_data_12__13), .d_arr_mux_12__12 (
               ordered_img_data_12__12), .d_arr_mux_12__11 (
               ordered_img_data_12__11), .d_arr_mux_12__10 (
               ordered_img_data_12__10), .d_arr_mux_12__9 (
               ordered_img_data_12__9), .d_arr_mux_12__8 (ordered_img_data_12__8
               ), .d_arr_mux_12__7 (ordered_img_data_12__7), .d_arr_mux_12__6 (
               ordered_img_data_12__6), .d_arr_mux_12__5 (ordered_img_data_12__5
               ), .d_arr_mux_12__4 (ordered_img_data_12__4), .d_arr_mux_12__3 (
               ordered_img_data_12__3), .d_arr_mux_12__2 (ordered_img_data_12__2
               ), .d_arr_mux_12__1 (ordered_img_data_12__1), .d_arr_mux_12__0 (
               ordered_img_data_12__0), .d_arr_mux_13__31 (nx16433), .d_arr_mux_13__30 (
               nx16433), .d_arr_mux_13__29 (nx16433), .d_arr_mux_13__28 (nx16433
               ), .d_arr_mux_13__27 (nx16433), .d_arr_mux_13__26 (nx16433), .d_arr_mux_13__25 (
               nx16433), .d_arr_mux_13__24 (nx16435), .d_arr_mux_13__23 (nx16435
               ), .d_arr_mux_13__22 (nx16435), .d_arr_mux_13__21 (nx16435), .d_arr_mux_13__20 (
               nx16435), .d_arr_mux_13__19 (nx16435), .d_arr_mux_13__18 (nx16435
               ), .d_arr_mux_13__17 (nx16437), .d_arr_mux_13__16 (nx16437), .d_arr_mux_13__15 (
               nx16437), .d_arr_mux_13__14 (ordered_img_data_13__14), .d_arr_mux_13__13 (
               ordered_img_data_13__13), .d_arr_mux_13__12 (
               ordered_img_data_13__12), .d_arr_mux_13__11 (
               ordered_img_data_13__11), .d_arr_mux_13__10 (
               ordered_img_data_13__10), .d_arr_mux_13__9 (
               ordered_img_data_13__9), .d_arr_mux_13__8 (ordered_img_data_13__8
               ), .d_arr_mux_13__7 (ordered_img_data_13__7), .d_arr_mux_13__6 (
               ordered_img_data_13__6), .d_arr_mux_13__5 (ordered_img_data_13__5
               ), .d_arr_mux_13__4 (ordered_img_data_13__4), .d_arr_mux_13__3 (
               ordered_img_data_13__3), .d_arr_mux_13__2 (ordered_img_data_13__2
               ), .d_arr_mux_13__1 (ordered_img_data_13__1), .d_arr_mux_13__0 (
               ordered_img_data_13__0), .d_arr_mux_14__31 (nx16441), .d_arr_mux_14__30 (
               nx16441), .d_arr_mux_14__29 (nx16441), .d_arr_mux_14__28 (nx16441
               ), .d_arr_mux_14__27 (nx16441), .d_arr_mux_14__26 (nx16441), .d_arr_mux_14__25 (
               nx16441), .d_arr_mux_14__24 (nx16443), .d_arr_mux_14__23 (nx16443
               ), .d_arr_mux_14__22 (nx16443), .d_arr_mux_14__21 (nx16443), .d_arr_mux_14__20 (
               nx16443), .d_arr_mux_14__19 (nx16443), .d_arr_mux_14__18 (nx16443
               ), .d_arr_mux_14__17 (nx16445), .d_arr_mux_14__16 (nx16445), .d_arr_mux_14__15 (
               nx16445), .d_arr_mux_14__14 (ordered_img_data_14__14), .d_arr_mux_14__13 (
               ordered_img_data_14__13), .d_arr_mux_14__12 (
               ordered_img_data_14__12), .d_arr_mux_14__11 (
               ordered_img_data_14__11), .d_arr_mux_14__10 (
               ordered_img_data_14__10), .d_arr_mux_14__9 (
               ordered_img_data_14__9), .d_arr_mux_14__8 (ordered_img_data_14__8
               ), .d_arr_mux_14__7 (ordered_img_data_14__7), .d_arr_mux_14__6 (
               ordered_img_data_14__6), .d_arr_mux_14__5 (ordered_img_data_14__5
               ), .d_arr_mux_14__4 (ordered_img_data_14__4), .d_arr_mux_14__3 (
               ordered_img_data_14__3), .d_arr_mux_14__2 (ordered_img_data_14__2
               ), .d_arr_mux_14__1 (ordered_img_data_14__1), .d_arr_mux_14__0 (
               ordered_img_data_14__0), .d_arr_mux_15__31 (nx16449), .d_arr_mux_15__30 (
               nx16449), .d_arr_mux_15__29 (nx16449), .d_arr_mux_15__28 (nx16449
               ), .d_arr_mux_15__27 (nx16449), .d_arr_mux_15__26 (nx16449), .d_arr_mux_15__25 (
               nx16449), .d_arr_mux_15__24 (nx16451), .d_arr_mux_15__23 (nx16451
               ), .d_arr_mux_15__22 (nx16451), .d_arr_mux_15__21 (nx16451), .d_arr_mux_15__20 (
               nx16451), .d_arr_mux_15__19 (nx16451), .d_arr_mux_15__18 (nx16451
               ), .d_arr_mux_15__17 (nx16453), .d_arr_mux_15__16 (nx16453), .d_arr_mux_15__15 (
               nx16453), .d_arr_mux_15__14 (ordered_img_data_15__14), .d_arr_mux_15__13 (
               ordered_img_data_15__13), .d_arr_mux_15__12 (
               ordered_img_data_15__12), .d_arr_mux_15__11 (
               ordered_img_data_15__11), .d_arr_mux_15__10 (
               ordered_img_data_15__10), .d_arr_mux_15__9 (
               ordered_img_data_15__9), .d_arr_mux_15__8 (ordered_img_data_15__8
               ), .d_arr_mux_15__7 (ordered_img_data_15__7), .d_arr_mux_15__6 (
               ordered_img_data_15__6), .d_arr_mux_15__5 (ordered_img_data_15__5
               ), .d_arr_mux_15__4 (ordered_img_data_15__4), .d_arr_mux_15__3 (
               ordered_img_data_15__3), .d_arr_mux_15__2 (ordered_img_data_15__2
               ), .d_arr_mux_15__1 (ordered_img_data_15__1), .d_arr_mux_15__0 (
               ordered_img_data_15__0), .d_arr_mux_16__31 (nx16457), .d_arr_mux_16__30 (
               nx16457), .d_arr_mux_16__29 (nx16457), .d_arr_mux_16__28 (nx16457
               ), .d_arr_mux_16__27 (nx16457), .d_arr_mux_16__26 (nx16457), .d_arr_mux_16__25 (
               nx16457), .d_arr_mux_16__24 (nx16459), .d_arr_mux_16__23 (nx16459
               ), .d_arr_mux_16__22 (nx16459), .d_arr_mux_16__21 (nx16459), .d_arr_mux_16__20 (
               nx16459), .d_arr_mux_16__19 (nx16459), .d_arr_mux_16__18 (nx16459
               ), .d_arr_mux_16__17 (nx16461), .d_arr_mux_16__16 (nx16461), .d_arr_mux_16__15 (
               nx16461), .d_arr_mux_16__14 (ordered_img_data_16__14), .d_arr_mux_16__13 (
               ordered_img_data_16__13), .d_arr_mux_16__12 (
               ordered_img_data_16__12), .d_arr_mux_16__11 (
               ordered_img_data_16__11), .d_arr_mux_16__10 (
               ordered_img_data_16__10), .d_arr_mux_16__9 (
               ordered_img_data_16__9), .d_arr_mux_16__8 (ordered_img_data_16__8
               ), .d_arr_mux_16__7 (ordered_img_data_16__7), .d_arr_mux_16__6 (
               ordered_img_data_16__6), .d_arr_mux_16__5 (ordered_img_data_16__5
               ), .d_arr_mux_16__4 (ordered_img_data_16__4), .d_arr_mux_16__3 (
               ordered_img_data_16__3), .d_arr_mux_16__2 (ordered_img_data_16__2
               ), .d_arr_mux_16__1 (ordered_img_data_16__1), .d_arr_mux_16__0 (
               ordered_img_data_16__0), .d_arr_mux_17__31 (nx16465), .d_arr_mux_17__30 (
               nx16465), .d_arr_mux_17__29 (nx16465), .d_arr_mux_17__28 (nx16465
               ), .d_arr_mux_17__27 (nx16465), .d_arr_mux_17__26 (nx16465), .d_arr_mux_17__25 (
               nx16465), .d_arr_mux_17__24 (nx16467), .d_arr_mux_17__23 (nx16467
               ), .d_arr_mux_17__22 (nx16467), .d_arr_mux_17__21 (nx16467), .d_arr_mux_17__20 (
               nx16467), .d_arr_mux_17__19 (nx16467), .d_arr_mux_17__18 (nx16467
               ), .d_arr_mux_17__17 (nx16469), .d_arr_mux_17__16 (nx16469), .d_arr_mux_17__15 (
               nx16469), .d_arr_mux_17__14 (ordered_img_data_17__14), .d_arr_mux_17__13 (
               ordered_img_data_17__13), .d_arr_mux_17__12 (
               ordered_img_data_17__12), .d_arr_mux_17__11 (
               ordered_img_data_17__11), .d_arr_mux_17__10 (
               ordered_img_data_17__10), .d_arr_mux_17__9 (
               ordered_img_data_17__9), .d_arr_mux_17__8 (ordered_img_data_17__8
               ), .d_arr_mux_17__7 (ordered_img_data_17__7), .d_arr_mux_17__6 (
               ordered_img_data_17__6), .d_arr_mux_17__5 (ordered_img_data_17__5
               ), .d_arr_mux_17__4 (ordered_img_data_17__4), .d_arr_mux_17__3 (
               ordered_img_data_17__3), .d_arr_mux_17__2 (ordered_img_data_17__2
               ), .d_arr_mux_17__1 (ordered_img_data_17__1), .d_arr_mux_17__0 (
               ordered_img_data_17__0), .d_arr_mux_18__31 (img_data_18__15), .d_arr_mux_18__30 (
               GND0), .d_arr_mux_18__29 (GND0), .d_arr_mux_18__28 (GND0), .d_arr_mux_18__27 (
               GND0), .d_arr_mux_18__26 (GND0), .d_arr_mux_18__25 (GND0), .d_arr_mux_18__24 (
               GND0), .d_arr_mux_18__23 (GND0), .d_arr_mux_18__22 (GND0), .d_arr_mux_18__21 (
               GND0), .d_arr_mux_18__20 (GND0), .d_arr_mux_18__19 (GND0), .d_arr_mux_18__18 (
               GND0), .d_arr_mux_18__17 (GND0), .d_arr_mux_18__16 (GND0), .d_arr_mux_18__15 (
               GND0), .d_arr_mux_18__14 (nx19438), .d_arr_mux_18__13 (
               img_data_18__13), .d_arr_mux_18__12 (img_data_18__12), .d_arr_mux_18__11 (
               img_data_18__11), .d_arr_mux_18__10 (img_data_18__10), .d_arr_mux_18__9 (
               img_data_18__9), .d_arr_mux_18__8 (img_data_18__8), .d_arr_mux_18__7 (
               img_data_18__7), .d_arr_mux_18__6 (img_data_18__6), .d_arr_mux_18__5 (
               img_data_18__5), .d_arr_mux_18__4 (img_data_18__4), .d_arr_mux_18__3 (
               img_data_18__3), .d_arr_mux_18__2 (img_data_18__2), .d_arr_mux_18__1 (
               img_data_18__1), .d_arr_mux_18__0 (img_data_18__0), .d_arr_mux_19__31 (
               img_data_19__15), .d_arr_mux_19__30 (GND0), .d_arr_mux_19__29 (
               GND0), .d_arr_mux_19__28 (GND0), .d_arr_mux_19__27 (GND0), .d_arr_mux_19__26 (
               GND0), .d_arr_mux_19__25 (GND0), .d_arr_mux_19__24 (GND0), .d_arr_mux_19__23 (
               GND0), .d_arr_mux_19__22 (GND0), .d_arr_mux_19__21 (GND0), .d_arr_mux_19__20 (
               GND0), .d_arr_mux_19__19 (GND0), .d_arr_mux_19__18 (GND0), .d_arr_mux_19__17 (
               GND0), .d_arr_mux_19__16 (GND0), .d_arr_mux_19__15 (GND0), .d_arr_mux_19__14 (
               img_data_19__14), .d_arr_mux_19__13 (img_data_19__13), .d_arr_mux_19__12 (
               img_data_19__12), .d_arr_mux_19__11 (img_data_19__11), .d_arr_mux_19__10 (
               img_data_19__10), .d_arr_mux_19__9 (img_data_19__9), .d_arr_mux_19__8 (
               img_data_19__8), .d_arr_mux_19__7 (img_data_19__7), .d_arr_mux_19__6 (
               img_data_19__6), .d_arr_mux_19__5 (img_data_19__5), .d_arr_mux_19__4 (
               img_data_19__4), .d_arr_mux_19__3 (img_data_19__3), .d_arr_mux_19__2 (
               img_data_19__2), .d_arr_mux_19__1 (img_data_19__1), .d_arr_mux_19__0 (
               img_data_19__0), .d_arr_mux_20__31 (img_data_20__15), .d_arr_mux_20__30 (
               GND0), .d_arr_mux_20__29 (GND0), .d_arr_mux_20__28 (GND0), .d_arr_mux_20__27 (
               GND0), .d_arr_mux_20__26 (GND0), .d_arr_mux_20__25 (GND0), .d_arr_mux_20__24 (
               GND0), .d_arr_mux_20__23 (GND0), .d_arr_mux_20__22 (GND0), .d_arr_mux_20__21 (
               GND0), .d_arr_mux_20__20 (GND0), .d_arr_mux_20__19 (GND0), .d_arr_mux_20__18 (
               GND0), .d_arr_mux_20__17 (GND0), .d_arr_mux_20__16 (GND0), .d_arr_mux_20__15 (
               GND0), .d_arr_mux_20__14 (nx19440), .d_arr_mux_20__13 (
               img_data_20__13), .d_arr_mux_20__12 (img_data_20__12), .d_arr_mux_20__11 (
               img_data_20__11), .d_arr_mux_20__10 (img_data_20__10), .d_arr_mux_20__9 (
               img_data_20__9), .d_arr_mux_20__8 (img_data_20__8), .d_arr_mux_20__7 (
               img_data_20__7), .d_arr_mux_20__6 (img_data_20__6), .d_arr_mux_20__5 (
               img_data_20__5), .d_arr_mux_20__4 (img_data_20__4), .d_arr_mux_20__3 (
               img_data_20__3), .d_arr_mux_20__2 (img_data_20__2), .d_arr_mux_20__1 (
               img_data_20__1), .d_arr_mux_20__0 (img_data_20__0), .d_arr_mux_21__31 (
               img_data_21__15), .d_arr_mux_21__30 (GND0), .d_arr_mux_21__29 (
               GND0), .d_arr_mux_21__28 (GND0), .d_arr_mux_21__27 (GND0), .d_arr_mux_21__26 (
               GND0), .d_arr_mux_21__25 (GND0), .d_arr_mux_21__24 (GND0), .d_arr_mux_21__23 (
               GND0), .d_arr_mux_21__22 (GND0), .d_arr_mux_21__21 (GND0), .d_arr_mux_21__20 (
               GND0), .d_arr_mux_21__19 (GND0), .d_arr_mux_21__18 (GND0), .d_arr_mux_21__17 (
               GND0), .d_arr_mux_21__16 (GND0), .d_arr_mux_21__15 (GND0), .d_arr_mux_21__14 (
               nx19442), .d_arr_mux_21__13 (img_data_21__13), .d_arr_mux_21__12 (
               img_data_21__12), .d_arr_mux_21__11 (img_data_21__11), .d_arr_mux_21__10 (
               img_data_21__10), .d_arr_mux_21__9 (img_data_21__9), .d_arr_mux_21__8 (
               img_data_21__8), .d_arr_mux_21__7 (img_data_21__7), .d_arr_mux_21__6 (
               img_data_21__6), .d_arr_mux_21__5 (img_data_21__5), .d_arr_mux_21__4 (
               img_data_21__4), .d_arr_mux_21__3 (img_data_21__3), .d_arr_mux_21__2 (
               img_data_21__2), .d_arr_mux_21__1 (img_data_21__1), .d_arr_mux_21__0 (
               img_data_21__0), .d_arr_mux_22__31 (img_data_22__15), .d_arr_mux_22__30 (
               GND0), .d_arr_mux_22__29 (GND0), .d_arr_mux_22__28 (GND0), .d_arr_mux_22__27 (
               GND0), .d_arr_mux_22__26 (GND0), .d_arr_mux_22__25 (GND0), .d_arr_mux_22__24 (
               GND0), .d_arr_mux_22__23 (GND0), .d_arr_mux_22__22 (GND0), .d_arr_mux_22__21 (
               GND0), .d_arr_mux_22__20 (GND0), .d_arr_mux_22__19 (GND0), .d_arr_mux_22__18 (
               GND0), .d_arr_mux_22__17 (GND0), .d_arr_mux_22__16 (GND0), .d_arr_mux_22__15 (
               GND0), .d_arr_mux_22__14 (nx19444), .d_arr_mux_22__13 (
               img_data_22__13), .d_arr_mux_22__12 (img_data_22__12), .d_arr_mux_22__11 (
               img_data_22__11), .d_arr_mux_22__10 (img_data_22__10), .d_arr_mux_22__9 (
               img_data_22__9), .d_arr_mux_22__8 (img_data_22__8), .d_arr_mux_22__7 (
               img_data_22__7), .d_arr_mux_22__6 (img_data_22__6), .d_arr_mux_22__5 (
               img_data_22__5), .d_arr_mux_22__4 (img_data_22__4), .d_arr_mux_22__3 (
               img_data_22__3), .d_arr_mux_22__2 (img_data_22__2), .d_arr_mux_22__1 (
               img_data_22__1), .d_arr_mux_22__0 (img_data_22__0), .d_arr_mux_23__31 (
               img_data_23__15), .d_arr_mux_23__30 (GND0), .d_arr_mux_23__29 (
               GND0), .d_arr_mux_23__28 (GND0), .d_arr_mux_23__27 (GND0), .d_arr_mux_23__26 (
               GND0), .d_arr_mux_23__25 (GND0), .d_arr_mux_23__24 (GND0), .d_arr_mux_23__23 (
               GND0), .d_arr_mux_23__22 (GND0), .d_arr_mux_23__21 (GND0), .d_arr_mux_23__20 (
               GND0), .d_arr_mux_23__19 (GND0), .d_arr_mux_23__18 (GND0), .d_arr_mux_23__17 (
               GND0), .d_arr_mux_23__16 (GND0), .d_arr_mux_23__15 (GND0), .d_arr_mux_23__14 (
               nx19446), .d_arr_mux_23__13 (img_data_23__13), .d_arr_mux_23__12 (
               img_data_23__12), .d_arr_mux_23__11 (img_data_23__11), .d_arr_mux_23__10 (
               img_data_23__10), .d_arr_mux_23__9 (img_data_23__9), .d_arr_mux_23__8 (
               img_data_23__8), .d_arr_mux_23__7 (img_data_23__7), .d_arr_mux_23__6 (
               img_data_23__6), .d_arr_mux_23__5 (img_data_23__5), .d_arr_mux_23__4 (
               img_data_23__4), .d_arr_mux_23__3 (img_data_23__3), .d_arr_mux_23__2 (
               img_data_23__2), .d_arr_mux_23__1 (img_data_23__1), .d_arr_mux_23__0 (
               img_data_23__0), .d_arr_mux_24__31 (img_data_24__15), .d_arr_mux_24__30 (
               GND0), .d_arr_mux_24__29 (GND0), .d_arr_mux_24__28 (GND0), .d_arr_mux_24__27 (
               GND0), .d_arr_mux_24__26 (GND0), .d_arr_mux_24__25 (GND0), .d_arr_mux_24__24 (
               GND0), .d_arr_mux_24__23 (GND0), .d_arr_mux_24__22 (GND0), .d_arr_mux_24__21 (
               GND0), .d_arr_mux_24__20 (GND0), .d_arr_mux_24__19 (GND0), .d_arr_mux_24__18 (
               GND0), .d_arr_mux_24__17 (GND0), .d_arr_mux_24__16 (GND0), .d_arr_mux_24__15 (
               GND0), .d_arr_mux_24__14 (img_data_24__14), .d_arr_mux_24__13 (
               img_data_24__13), .d_arr_mux_24__12 (img_data_24__12), .d_arr_mux_24__11 (
               img_data_24__11), .d_arr_mux_24__10 (img_data_24__10), .d_arr_mux_24__9 (
               img_data_24__9), .d_arr_mux_24__8 (img_data_24__8), .d_arr_mux_24__7 (
               img_data_24__7), .d_arr_mux_24__6 (img_data_24__6), .d_arr_mux_24__5 (
               img_data_24__5), .d_arr_mux_24__4 (img_data_24__4), .d_arr_mux_24__3 (
               img_data_24__3), .d_arr_mux_24__2 (img_data_24__2), .d_arr_mux_24__1 (
               img_data_24__1), .d_arr_mux_24__0 (img_data_24__0), .d_arr_mul_0__31 (
               d_arr_mul_0__31), .d_arr_mul_0__30 (d_arr_mul_0__30), .d_arr_mul_0__29 (
               d_arr_mul_0__29), .d_arr_mul_0__28 (d_arr_mul_0__28), .d_arr_mul_0__27 (
               d_arr_mul_0__27), .d_arr_mul_0__26 (d_arr_mul_0__26), .d_arr_mul_0__25 (
               d_arr_mul_0__25), .d_arr_mul_0__24 (d_arr_mul_0__24), .d_arr_mul_0__23 (
               d_arr_mul_0__23), .d_arr_mul_0__22 (d_arr_mul_0__22), .d_arr_mul_0__21 (
               d_arr_mul_0__21), .d_arr_mul_0__20 (d_arr_mul_0__20), .d_arr_mul_0__19 (
               d_arr_mul_0__19), .d_arr_mul_0__18 (d_arr_mul_0__18), .d_arr_mul_0__17 (
               d_arr_mul_0__17), .d_arr_mul_0__16 (d_arr_mul_0__16), .d_arr_mul_0__15 (
               d_arr_mul_0__15), .d_arr_mul_0__14 (d_arr_mul_0__14), .d_arr_mul_0__13 (
               d_arr_mul_0__13), .d_arr_mul_0__12 (d_arr_mul_0__12), .d_arr_mul_0__11 (
               d_arr_mul_0__11), .d_arr_mul_0__10 (d_arr_mul_0__10), .d_arr_mul_0__9 (
               d_arr_mul_0__9), .d_arr_mul_0__8 (d_arr_mul_0__8), .d_arr_mul_0__7 (
               d_arr_mul_0__7), .d_arr_mul_0__6 (d_arr_mul_0__6), .d_arr_mul_0__5 (
               d_arr_mul_0__5), .d_arr_mul_0__4 (d_arr_mul_0__4), .d_arr_mul_0__3 (
               d_arr_mul_0__3), .d_arr_mul_0__2 (d_arr_mul_0__2), .d_arr_mul_0__1 (
               d_arr_mul_0__1), .d_arr_mul_0__0 (d_arr_mul_0__0), .d_arr_mul_1__31 (
               d_arr_mul_1__31), .d_arr_mul_1__30 (d_arr_mul_1__30), .d_arr_mul_1__29 (
               d_arr_mul_1__29), .d_arr_mul_1__28 (d_arr_mul_1__28), .d_arr_mul_1__27 (
               d_arr_mul_1__27), .d_arr_mul_1__26 (d_arr_mul_1__26), .d_arr_mul_1__25 (
               d_arr_mul_1__25), .d_arr_mul_1__24 (d_arr_mul_1__24), .d_arr_mul_1__23 (
               d_arr_mul_1__23), .d_arr_mul_1__22 (d_arr_mul_1__22), .d_arr_mul_1__21 (
               d_arr_mul_1__21), .d_arr_mul_1__20 (d_arr_mul_1__20), .d_arr_mul_1__19 (
               d_arr_mul_1__19), .d_arr_mul_1__18 (d_arr_mul_1__18), .d_arr_mul_1__17 (
               d_arr_mul_1__17), .d_arr_mul_1__16 (d_arr_mul_1__16), .d_arr_mul_1__15 (
               d_arr_mul_1__15), .d_arr_mul_1__14 (d_arr_mul_1__14), .d_arr_mul_1__13 (
               d_arr_mul_1__13), .d_arr_mul_1__12 (d_arr_mul_1__12), .d_arr_mul_1__11 (
               d_arr_mul_1__11), .d_arr_mul_1__10 (d_arr_mul_1__10), .d_arr_mul_1__9 (
               d_arr_mul_1__9), .d_arr_mul_1__8 (d_arr_mul_1__8), .d_arr_mul_1__7 (
               d_arr_mul_1__7), .d_arr_mul_1__6 (d_arr_mul_1__6), .d_arr_mul_1__5 (
               d_arr_mul_1__5), .d_arr_mul_1__4 (d_arr_mul_1__4), .d_arr_mul_1__3 (
               d_arr_mul_1__3), .d_arr_mul_1__2 (d_arr_mul_1__2), .d_arr_mul_1__1 (
               d_arr_mul_1__1), .d_arr_mul_1__0 (d_arr_mul_1__0), .d_arr_mul_2__31 (
               d_arr_mul_2__31), .d_arr_mul_2__30 (d_arr_mul_2__30), .d_arr_mul_2__29 (
               d_arr_mul_2__29), .d_arr_mul_2__28 (d_arr_mul_2__28), .d_arr_mul_2__27 (
               d_arr_mul_2__27), .d_arr_mul_2__26 (d_arr_mul_2__26), .d_arr_mul_2__25 (
               d_arr_mul_2__25), .d_arr_mul_2__24 (d_arr_mul_2__24), .d_arr_mul_2__23 (
               d_arr_mul_2__23), .d_arr_mul_2__22 (d_arr_mul_2__22), .d_arr_mul_2__21 (
               d_arr_mul_2__21), .d_arr_mul_2__20 (d_arr_mul_2__20), .d_arr_mul_2__19 (
               d_arr_mul_2__19), .d_arr_mul_2__18 (d_arr_mul_2__18), .d_arr_mul_2__17 (
               d_arr_mul_2__17), .d_arr_mul_2__16 (d_arr_mul_2__16), .d_arr_mul_2__15 (
               d_arr_mul_2__15), .d_arr_mul_2__14 (d_arr_mul_2__14), .d_arr_mul_2__13 (
               d_arr_mul_2__13), .d_arr_mul_2__12 (d_arr_mul_2__12), .d_arr_mul_2__11 (
               d_arr_mul_2__11), .d_arr_mul_2__10 (d_arr_mul_2__10), .d_arr_mul_2__9 (
               d_arr_mul_2__9), .d_arr_mul_2__8 (d_arr_mul_2__8), .d_arr_mul_2__7 (
               d_arr_mul_2__7), .d_arr_mul_2__6 (d_arr_mul_2__6), .d_arr_mul_2__5 (
               d_arr_mul_2__5), .d_arr_mul_2__4 (d_arr_mul_2__4), .d_arr_mul_2__3 (
               d_arr_mul_2__3), .d_arr_mul_2__2 (d_arr_mul_2__2), .d_arr_mul_2__1 (
               d_arr_mul_2__1), .d_arr_mul_2__0 (d_arr_mul_2__0), .d_arr_mul_3__31 (
               d_arr_mul_3__31), .d_arr_mul_3__30 (d_arr_mul_3__30), .d_arr_mul_3__29 (
               d_arr_mul_3__29), .d_arr_mul_3__28 (d_arr_mul_3__28), .d_arr_mul_3__27 (
               d_arr_mul_3__27), .d_arr_mul_3__26 (d_arr_mul_3__26), .d_arr_mul_3__25 (
               d_arr_mul_3__25), .d_arr_mul_3__24 (d_arr_mul_3__24), .d_arr_mul_3__23 (
               d_arr_mul_3__23), .d_arr_mul_3__22 (d_arr_mul_3__22), .d_arr_mul_3__21 (
               d_arr_mul_3__21), .d_arr_mul_3__20 (d_arr_mul_3__20), .d_arr_mul_3__19 (
               d_arr_mul_3__19), .d_arr_mul_3__18 (d_arr_mul_3__18), .d_arr_mul_3__17 (
               d_arr_mul_3__17), .d_arr_mul_3__16 (d_arr_mul_3__16), .d_arr_mul_3__15 (
               d_arr_mul_3__15), .d_arr_mul_3__14 (d_arr_mul_3__14), .d_arr_mul_3__13 (
               d_arr_mul_3__13), .d_arr_mul_3__12 (d_arr_mul_3__12), .d_arr_mul_3__11 (
               d_arr_mul_3__11), .d_arr_mul_3__10 (d_arr_mul_3__10), .d_arr_mul_3__9 (
               d_arr_mul_3__9), .d_arr_mul_3__8 (d_arr_mul_3__8), .d_arr_mul_3__7 (
               d_arr_mul_3__7), .d_arr_mul_3__6 (d_arr_mul_3__6), .d_arr_mul_3__5 (
               d_arr_mul_3__5), .d_arr_mul_3__4 (d_arr_mul_3__4), .d_arr_mul_3__3 (
               d_arr_mul_3__3), .d_arr_mul_3__2 (d_arr_mul_3__2), .d_arr_mul_3__1 (
               d_arr_mul_3__1), .d_arr_mul_3__0 (d_arr_mul_3__0), .d_arr_mul_4__31 (
               d_arr_mul_4__31), .d_arr_mul_4__30 (d_arr_mul_4__30), .d_arr_mul_4__29 (
               d_arr_mul_4__29), .d_arr_mul_4__28 (d_arr_mul_4__28), .d_arr_mul_4__27 (
               d_arr_mul_4__27), .d_arr_mul_4__26 (d_arr_mul_4__26), .d_arr_mul_4__25 (
               d_arr_mul_4__25), .d_arr_mul_4__24 (d_arr_mul_4__24), .d_arr_mul_4__23 (
               d_arr_mul_4__23), .d_arr_mul_4__22 (d_arr_mul_4__22), .d_arr_mul_4__21 (
               d_arr_mul_4__21), .d_arr_mul_4__20 (d_arr_mul_4__20), .d_arr_mul_4__19 (
               d_arr_mul_4__19), .d_arr_mul_4__18 (d_arr_mul_4__18), .d_arr_mul_4__17 (
               d_arr_mul_4__17), .d_arr_mul_4__16 (d_arr_mul_4__16), .d_arr_mul_4__15 (
               d_arr_mul_4__15), .d_arr_mul_4__14 (d_arr_mul_4__14), .d_arr_mul_4__13 (
               d_arr_mul_4__13), .d_arr_mul_4__12 (d_arr_mul_4__12), .d_arr_mul_4__11 (
               d_arr_mul_4__11), .d_arr_mul_4__10 (d_arr_mul_4__10), .d_arr_mul_4__9 (
               d_arr_mul_4__9), .d_arr_mul_4__8 (d_arr_mul_4__8), .d_arr_mul_4__7 (
               d_arr_mul_4__7), .d_arr_mul_4__6 (d_arr_mul_4__6), .d_arr_mul_4__5 (
               d_arr_mul_4__5), .d_arr_mul_4__4 (d_arr_mul_4__4), .d_arr_mul_4__3 (
               d_arr_mul_4__3), .d_arr_mul_4__2 (d_arr_mul_4__2), .d_arr_mul_4__1 (
               d_arr_mul_4__1), .d_arr_mul_4__0 (d_arr_mul_4__0), .d_arr_mul_5__31 (
               d_arr_mul_5__31), .d_arr_mul_5__30 (d_arr_mul_5__30), .d_arr_mul_5__29 (
               d_arr_mul_5__29), .d_arr_mul_5__28 (d_arr_mul_5__28), .d_arr_mul_5__27 (
               d_arr_mul_5__27), .d_arr_mul_5__26 (d_arr_mul_5__26), .d_arr_mul_5__25 (
               d_arr_mul_5__25), .d_arr_mul_5__24 (d_arr_mul_5__24), .d_arr_mul_5__23 (
               d_arr_mul_5__23), .d_arr_mul_5__22 (d_arr_mul_5__22), .d_arr_mul_5__21 (
               d_arr_mul_5__21), .d_arr_mul_5__20 (d_arr_mul_5__20), .d_arr_mul_5__19 (
               d_arr_mul_5__19), .d_arr_mul_5__18 (d_arr_mul_5__18), .d_arr_mul_5__17 (
               d_arr_mul_5__17), .d_arr_mul_5__16 (d_arr_mul_5__16), .d_arr_mul_5__15 (
               d_arr_mul_5__15), .d_arr_mul_5__14 (d_arr_mul_5__14), .d_arr_mul_5__13 (
               d_arr_mul_5__13), .d_arr_mul_5__12 (d_arr_mul_5__12), .d_arr_mul_5__11 (
               d_arr_mul_5__11), .d_arr_mul_5__10 (d_arr_mul_5__10), .d_arr_mul_5__9 (
               d_arr_mul_5__9), .d_arr_mul_5__8 (d_arr_mul_5__8), .d_arr_mul_5__7 (
               d_arr_mul_5__7), .d_arr_mul_5__6 (d_arr_mul_5__6), .d_arr_mul_5__5 (
               d_arr_mul_5__5), .d_arr_mul_5__4 (d_arr_mul_5__4), .d_arr_mul_5__3 (
               d_arr_mul_5__3), .d_arr_mul_5__2 (d_arr_mul_5__2), .d_arr_mul_5__1 (
               d_arr_mul_5__1), .d_arr_mul_5__0 (d_arr_mul_5__0), .d_arr_mul_6__31 (
               d_arr_mul_6__31), .d_arr_mul_6__30 (d_arr_mul_6__30), .d_arr_mul_6__29 (
               d_arr_mul_6__29), .d_arr_mul_6__28 (d_arr_mul_6__28), .d_arr_mul_6__27 (
               d_arr_mul_6__27), .d_arr_mul_6__26 (d_arr_mul_6__26), .d_arr_mul_6__25 (
               d_arr_mul_6__25), .d_arr_mul_6__24 (d_arr_mul_6__24), .d_arr_mul_6__23 (
               d_arr_mul_6__23), .d_arr_mul_6__22 (d_arr_mul_6__22), .d_arr_mul_6__21 (
               d_arr_mul_6__21), .d_arr_mul_6__20 (d_arr_mul_6__20), .d_arr_mul_6__19 (
               d_arr_mul_6__19), .d_arr_mul_6__18 (d_arr_mul_6__18), .d_arr_mul_6__17 (
               d_arr_mul_6__17), .d_arr_mul_6__16 (d_arr_mul_6__16), .d_arr_mul_6__15 (
               d_arr_mul_6__15), .d_arr_mul_6__14 (d_arr_mul_6__14), .d_arr_mul_6__13 (
               d_arr_mul_6__13), .d_arr_mul_6__12 (d_arr_mul_6__12), .d_arr_mul_6__11 (
               d_arr_mul_6__11), .d_arr_mul_6__10 (d_arr_mul_6__10), .d_arr_mul_6__9 (
               d_arr_mul_6__9), .d_arr_mul_6__8 (d_arr_mul_6__8), .d_arr_mul_6__7 (
               d_arr_mul_6__7), .d_arr_mul_6__6 (d_arr_mul_6__6), .d_arr_mul_6__5 (
               d_arr_mul_6__5), .d_arr_mul_6__4 (d_arr_mul_6__4), .d_arr_mul_6__3 (
               d_arr_mul_6__3), .d_arr_mul_6__2 (d_arr_mul_6__2), .d_arr_mul_6__1 (
               d_arr_mul_6__1), .d_arr_mul_6__0 (d_arr_mul_6__0), .d_arr_mul_7__31 (
               d_arr_mul_7__31), .d_arr_mul_7__30 (d_arr_mul_7__30), .d_arr_mul_7__29 (
               d_arr_mul_7__29), .d_arr_mul_7__28 (d_arr_mul_7__28), .d_arr_mul_7__27 (
               d_arr_mul_7__27), .d_arr_mul_7__26 (d_arr_mul_7__26), .d_arr_mul_7__25 (
               d_arr_mul_7__25), .d_arr_mul_7__24 (d_arr_mul_7__24), .d_arr_mul_7__23 (
               d_arr_mul_7__23), .d_arr_mul_7__22 (d_arr_mul_7__22), .d_arr_mul_7__21 (
               d_arr_mul_7__21), .d_arr_mul_7__20 (d_arr_mul_7__20), .d_arr_mul_7__19 (
               d_arr_mul_7__19), .d_arr_mul_7__18 (d_arr_mul_7__18), .d_arr_mul_7__17 (
               d_arr_mul_7__17), .d_arr_mul_7__16 (d_arr_mul_7__16), .d_arr_mul_7__15 (
               d_arr_mul_7__15), .d_arr_mul_7__14 (d_arr_mul_7__14), .d_arr_mul_7__13 (
               d_arr_mul_7__13), .d_arr_mul_7__12 (d_arr_mul_7__12), .d_arr_mul_7__11 (
               d_arr_mul_7__11), .d_arr_mul_7__10 (d_arr_mul_7__10), .d_arr_mul_7__9 (
               d_arr_mul_7__9), .d_arr_mul_7__8 (d_arr_mul_7__8), .d_arr_mul_7__7 (
               d_arr_mul_7__7), .d_arr_mul_7__6 (d_arr_mul_7__6), .d_arr_mul_7__5 (
               d_arr_mul_7__5), .d_arr_mul_7__4 (d_arr_mul_7__4), .d_arr_mul_7__3 (
               d_arr_mul_7__3), .d_arr_mul_7__2 (d_arr_mul_7__2), .d_arr_mul_7__1 (
               d_arr_mul_7__1), .d_arr_mul_7__0 (d_arr_mul_7__0), .d_arr_mul_8__31 (
               d_arr_mul_8__31), .d_arr_mul_8__30 (d_arr_mul_8__30), .d_arr_mul_8__29 (
               d_arr_mul_8__29), .d_arr_mul_8__28 (d_arr_mul_8__28), .d_arr_mul_8__27 (
               d_arr_mul_8__27), .d_arr_mul_8__26 (d_arr_mul_8__26), .d_arr_mul_8__25 (
               d_arr_mul_8__25), .d_arr_mul_8__24 (d_arr_mul_8__24), .d_arr_mul_8__23 (
               d_arr_mul_8__23), .d_arr_mul_8__22 (d_arr_mul_8__22), .d_arr_mul_8__21 (
               d_arr_mul_8__21), .d_arr_mul_8__20 (d_arr_mul_8__20), .d_arr_mul_8__19 (
               d_arr_mul_8__19), .d_arr_mul_8__18 (d_arr_mul_8__18), .d_arr_mul_8__17 (
               d_arr_mul_8__17), .d_arr_mul_8__16 (d_arr_mul_8__16), .d_arr_mul_8__15 (
               d_arr_mul_8__15), .d_arr_mul_8__14 (d_arr_mul_8__14), .d_arr_mul_8__13 (
               d_arr_mul_8__13), .d_arr_mul_8__12 (d_arr_mul_8__12), .d_arr_mul_8__11 (
               d_arr_mul_8__11), .d_arr_mul_8__10 (d_arr_mul_8__10), .d_arr_mul_8__9 (
               d_arr_mul_8__9), .d_arr_mul_8__8 (d_arr_mul_8__8), .d_arr_mul_8__7 (
               d_arr_mul_8__7), .d_arr_mul_8__6 (d_arr_mul_8__6), .d_arr_mul_8__5 (
               d_arr_mul_8__5), .d_arr_mul_8__4 (d_arr_mul_8__4), .d_arr_mul_8__3 (
               d_arr_mul_8__3), .d_arr_mul_8__2 (d_arr_mul_8__2), .d_arr_mul_8__1 (
               d_arr_mul_8__1), .d_arr_mul_8__0 (d_arr_mul_8__0), .d_arr_mul_9__31 (
               d_arr_mul_9__31), .d_arr_mul_9__30 (d_arr_mul_9__30), .d_arr_mul_9__29 (
               d_arr_mul_9__29), .d_arr_mul_9__28 (d_arr_mul_9__28), .d_arr_mul_9__27 (
               d_arr_mul_9__27), .d_arr_mul_9__26 (d_arr_mul_9__26), .d_arr_mul_9__25 (
               d_arr_mul_9__25), .d_arr_mul_9__24 (d_arr_mul_9__24), .d_arr_mul_9__23 (
               d_arr_mul_9__23), .d_arr_mul_9__22 (d_arr_mul_9__22), .d_arr_mul_9__21 (
               d_arr_mul_9__21), .d_arr_mul_9__20 (d_arr_mul_9__20), .d_arr_mul_9__19 (
               d_arr_mul_9__19), .d_arr_mul_9__18 (d_arr_mul_9__18), .d_arr_mul_9__17 (
               d_arr_mul_9__17), .d_arr_mul_9__16 (d_arr_mul_9__16), .d_arr_mul_9__15 (
               d_arr_mul_9__15), .d_arr_mul_9__14 (d_arr_mul_9__14), .d_arr_mul_9__13 (
               d_arr_mul_9__13), .d_arr_mul_9__12 (d_arr_mul_9__12), .d_arr_mul_9__11 (
               d_arr_mul_9__11), .d_arr_mul_9__10 (d_arr_mul_9__10), .d_arr_mul_9__9 (
               d_arr_mul_9__9), .d_arr_mul_9__8 (d_arr_mul_9__8), .d_arr_mul_9__7 (
               d_arr_mul_9__7), .d_arr_mul_9__6 (d_arr_mul_9__6), .d_arr_mul_9__5 (
               d_arr_mul_9__5), .d_arr_mul_9__4 (d_arr_mul_9__4), .d_arr_mul_9__3 (
               d_arr_mul_9__3), .d_arr_mul_9__2 (d_arr_mul_9__2), .d_arr_mul_9__1 (
               d_arr_mul_9__1), .d_arr_mul_9__0 (d_arr_mul_9__0), .d_arr_mul_10__31 (
               d_arr_mul_10__31), .d_arr_mul_10__30 (d_arr_mul_10__30), .d_arr_mul_10__29 (
               d_arr_mul_10__29), .d_arr_mul_10__28 (d_arr_mul_10__28), .d_arr_mul_10__27 (
               d_arr_mul_10__27), .d_arr_mul_10__26 (d_arr_mul_10__26), .d_arr_mul_10__25 (
               d_arr_mul_10__25), .d_arr_mul_10__24 (d_arr_mul_10__24), .d_arr_mul_10__23 (
               d_arr_mul_10__23), .d_arr_mul_10__22 (d_arr_mul_10__22), .d_arr_mul_10__21 (
               d_arr_mul_10__21), .d_arr_mul_10__20 (d_arr_mul_10__20), .d_arr_mul_10__19 (
               d_arr_mul_10__19), .d_arr_mul_10__18 (d_arr_mul_10__18), .d_arr_mul_10__17 (
               d_arr_mul_10__17), .d_arr_mul_10__16 (d_arr_mul_10__16), .d_arr_mul_10__15 (
               d_arr_mul_10__15), .d_arr_mul_10__14 (d_arr_mul_10__14), .d_arr_mul_10__13 (
               d_arr_mul_10__13), .d_arr_mul_10__12 (d_arr_mul_10__12), .d_arr_mul_10__11 (
               d_arr_mul_10__11), .d_arr_mul_10__10 (d_arr_mul_10__10), .d_arr_mul_10__9 (
               d_arr_mul_10__9), .d_arr_mul_10__8 (d_arr_mul_10__8), .d_arr_mul_10__7 (
               d_arr_mul_10__7), .d_arr_mul_10__6 (d_arr_mul_10__6), .d_arr_mul_10__5 (
               d_arr_mul_10__5), .d_arr_mul_10__4 (d_arr_mul_10__4), .d_arr_mul_10__3 (
               d_arr_mul_10__3), .d_arr_mul_10__2 (d_arr_mul_10__2), .d_arr_mul_10__1 (
               d_arr_mul_10__1), .d_arr_mul_10__0 (d_arr_mul_10__0), .d_arr_mul_11__31 (
               d_arr_mul_11__31), .d_arr_mul_11__30 (d_arr_mul_11__30), .d_arr_mul_11__29 (
               d_arr_mul_11__29), .d_arr_mul_11__28 (d_arr_mul_11__28), .d_arr_mul_11__27 (
               d_arr_mul_11__27), .d_arr_mul_11__26 (d_arr_mul_11__26), .d_arr_mul_11__25 (
               d_arr_mul_11__25), .d_arr_mul_11__24 (d_arr_mul_11__24), .d_arr_mul_11__23 (
               d_arr_mul_11__23), .d_arr_mul_11__22 (d_arr_mul_11__22), .d_arr_mul_11__21 (
               d_arr_mul_11__21), .d_arr_mul_11__20 (d_arr_mul_11__20), .d_arr_mul_11__19 (
               d_arr_mul_11__19), .d_arr_mul_11__18 (d_arr_mul_11__18), .d_arr_mul_11__17 (
               d_arr_mul_11__17), .d_arr_mul_11__16 (d_arr_mul_11__16), .d_arr_mul_11__15 (
               d_arr_mul_11__15), .d_arr_mul_11__14 (d_arr_mul_11__14), .d_arr_mul_11__13 (
               d_arr_mul_11__13), .d_arr_mul_11__12 (d_arr_mul_11__12), .d_arr_mul_11__11 (
               d_arr_mul_11__11), .d_arr_mul_11__10 (d_arr_mul_11__10), .d_arr_mul_11__9 (
               d_arr_mul_11__9), .d_arr_mul_11__8 (d_arr_mul_11__8), .d_arr_mul_11__7 (
               d_arr_mul_11__7), .d_arr_mul_11__6 (d_arr_mul_11__6), .d_arr_mul_11__5 (
               d_arr_mul_11__5), .d_arr_mul_11__4 (d_arr_mul_11__4), .d_arr_mul_11__3 (
               d_arr_mul_11__3), .d_arr_mul_11__2 (d_arr_mul_11__2), .d_arr_mul_11__1 (
               d_arr_mul_11__1), .d_arr_mul_11__0 (d_arr_mul_11__0), .d_arr_mul_12__31 (
               d_arr_mul_12__31), .d_arr_mul_12__30 (d_arr_mul_12__30), .d_arr_mul_12__29 (
               d_arr_mul_12__29), .d_arr_mul_12__28 (d_arr_mul_12__28), .d_arr_mul_12__27 (
               d_arr_mul_12__27), .d_arr_mul_12__26 (d_arr_mul_12__26), .d_arr_mul_12__25 (
               d_arr_mul_12__25), .d_arr_mul_12__24 (d_arr_mul_12__24), .d_arr_mul_12__23 (
               d_arr_mul_12__23), .d_arr_mul_12__22 (d_arr_mul_12__22), .d_arr_mul_12__21 (
               d_arr_mul_12__21), .d_arr_mul_12__20 (d_arr_mul_12__20), .d_arr_mul_12__19 (
               d_arr_mul_12__19), .d_arr_mul_12__18 (d_arr_mul_12__18), .d_arr_mul_12__17 (
               d_arr_mul_12__17), .d_arr_mul_12__16 (d_arr_mul_12__16), .d_arr_mul_12__15 (
               d_arr_mul_12__15), .d_arr_mul_12__14 (d_arr_mul_12__14), .d_arr_mul_12__13 (
               d_arr_mul_12__13), .d_arr_mul_12__12 (d_arr_mul_12__12), .d_arr_mul_12__11 (
               d_arr_mul_12__11), .d_arr_mul_12__10 (d_arr_mul_12__10), .d_arr_mul_12__9 (
               d_arr_mul_12__9), .d_arr_mul_12__8 (d_arr_mul_12__8), .d_arr_mul_12__7 (
               d_arr_mul_12__7), .d_arr_mul_12__6 (d_arr_mul_12__6), .d_arr_mul_12__5 (
               d_arr_mul_12__5), .d_arr_mul_12__4 (d_arr_mul_12__4), .d_arr_mul_12__3 (
               d_arr_mul_12__3), .d_arr_mul_12__2 (d_arr_mul_12__2), .d_arr_mul_12__1 (
               d_arr_mul_12__1), .d_arr_mul_12__0 (d_arr_mul_12__0), .d_arr_mul_13__31 (
               d_arr_mul_13__31), .d_arr_mul_13__30 (d_arr_mul_13__30), .d_arr_mul_13__29 (
               d_arr_mul_13__29), .d_arr_mul_13__28 (d_arr_mul_13__28), .d_arr_mul_13__27 (
               d_arr_mul_13__27), .d_arr_mul_13__26 (d_arr_mul_13__26), .d_arr_mul_13__25 (
               d_arr_mul_13__25), .d_arr_mul_13__24 (d_arr_mul_13__24), .d_arr_mul_13__23 (
               d_arr_mul_13__23), .d_arr_mul_13__22 (d_arr_mul_13__22), .d_arr_mul_13__21 (
               d_arr_mul_13__21), .d_arr_mul_13__20 (d_arr_mul_13__20), .d_arr_mul_13__19 (
               d_arr_mul_13__19), .d_arr_mul_13__18 (d_arr_mul_13__18), .d_arr_mul_13__17 (
               d_arr_mul_13__17), .d_arr_mul_13__16 (d_arr_mul_13__16), .d_arr_mul_13__15 (
               d_arr_mul_13__15), .d_arr_mul_13__14 (d_arr_mul_13__14), .d_arr_mul_13__13 (
               d_arr_mul_13__13), .d_arr_mul_13__12 (d_arr_mul_13__12), .d_arr_mul_13__11 (
               d_arr_mul_13__11), .d_arr_mul_13__10 (d_arr_mul_13__10), .d_arr_mul_13__9 (
               d_arr_mul_13__9), .d_arr_mul_13__8 (d_arr_mul_13__8), .d_arr_mul_13__7 (
               d_arr_mul_13__7), .d_arr_mul_13__6 (d_arr_mul_13__6), .d_arr_mul_13__5 (
               d_arr_mul_13__5), .d_arr_mul_13__4 (d_arr_mul_13__4), .d_arr_mul_13__3 (
               d_arr_mul_13__3), .d_arr_mul_13__2 (d_arr_mul_13__2), .d_arr_mul_13__1 (
               d_arr_mul_13__1), .d_arr_mul_13__0 (d_arr_mul_13__0), .d_arr_mul_14__31 (
               d_arr_mul_14__31), .d_arr_mul_14__30 (d_arr_mul_14__30), .d_arr_mul_14__29 (
               d_arr_mul_14__29), .d_arr_mul_14__28 (d_arr_mul_14__28), .d_arr_mul_14__27 (
               d_arr_mul_14__27), .d_arr_mul_14__26 (d_arr_mul_14__26), .d_arr_mul_14__25 (
               d_arr_mul_14__25), .d_arr_mul_14__24 (d_arr_mul_14__24), .d_arr_mul_14__23 (
               d_arr_mul_14__23), .d_arr_mul_14__22 (d_arr_mul_14__22), .d_arr_mul_14__21 (
               d_arr_mul_14__21), .d_arr_mul_14__20 (d_arr_mul_14__20), .d_arr_mul_14__19 (
               d_arr_mul_14__19), .d_arr_mul_14__18 (d_arr_mul_14__18), .d_arr_mul_14__17 (
               d_arr_mul_14__17), .d_arr_mul_14__16 (d_arr_mul_14__16), .d_arr_mul_14__15 (
               d_arr_mul_14__15), .d_arr_mul_14__14 (d_arr_mul_14__14), .d_arr_mul_14__13 (
               d_arr_mul_14__13), .d_arr_mul_14__12 (d_arr_mul_14__12), .d_arr_mul_14__11 (
               d_arr_mul_14__11), .d_arr_mul_14__10 (d_arr_mul_14__10), .d_arr_mul_14__9 (
               d_arr_mul_14__9), .d_arr_mul_14__8 (d_arr_mul_14__8), .d_arr_mul_14__7 (
               d_arr_mul_14__7), .d_arr_mul_14__6 (d_arr_mul_14__6), .d_arr_mul_14__5 (
               d_arr_mul_14__5), .d_arr_mul_14__4 (d_arr_mul_14__4), .d_arr_mul_14__3 (
               d_arr_mul_14__3), .d_arr_mul_14__2 (d_arr_mul_14__2), .d_arr_mul_14__1 (
               d_arr_mul_14__1), .d_arr_mul_14__0 (d_arr_mul_14__0), .d_arr_mul_15__31 (
               d_arr_mul_15__31), .d_arr_mul_15__30 (d_arr_mul_15__30), .d_arr_mul_15__29 (
               d_arr_mul_15__29), .d_arr_mul_15__28 (d_arr_mul_15__28), .d_arr_mul_15__27 (
               d_arr_mul_15__27), .d_arr_mul_15__26 (d_arr_mul_15__26), .d_arr_mul_15__25 (
               d_arr_mul_15__25), .d_arr_mul_15__24 (d_arr_mul_15__24), .d_arr_mul_15__23 (
               d_arr_mul_15__23), .d_arr_mul_15__22 (d_arr_mul_15__22), .d_arr_mul_15__21 (
               d_arr_mul_15__21), .d_arr_mul_15__20 (d_arr_mul_15__20), .d_arr_mul_15__19 (
               d_arr_mul_15__19), .d_arr_mul_15__18 (d_arr_mul_15__18), .d_arr_mul_15__17 (
               d_arr_mul_15__17), .d_arr_mul_15__16 (d_arr_mul_15__16), .d_arr_mul_15__15 (
               d_arr_mul_15__15), .d_arr_mul_15__14 (d_arr_mul_15__14), .d_arr_mul_15__13 (
               d_arr_mul_15__13), .d_arr_mul_15__12 (d_arr_mul_15__12), .d_arr_mul_15__11 (
               d_arr_mul_15__11), .d_arr_mul_15__10 (d_arr_mul_15__10), .d_arr_mul_15__9 (
               d_arr_mul_15__9), .d_arr_mul_15__8 (d_arr_mul_15__8), .d_arr_mul_15__7 (
               d_arr_mul_15__7), .d_arr_mul_15__6 (d_arr_mul_15__6), .d_arr_mul_15__5 (
               d_arr_mul_15__5), .d_arr_mul_15__4 (d_arr_mul_15__4), .d_arr_mul_15__3 (
               d_arr_mul_15__3), .d_arr_mul_15__2 (d_arr_mul_15__2), .d_arr_mul_15__1 (
               d_arr_mul_15__1), .d_arr_mul_15__0 (d_arr_mul_15__0), .d_arr_mul_16__31 (
               d_arr_mul_16__31), .d_arr_mul_16__30 (d_arr_mul_16__30), .d_arr_mul_16__29 (
               d_arr_mul_16__29), .d_arr_mul_16__28 (d_arr_mul_16__28), .d_arr_mul_16__27 (
               d_arr_mul_16__27), .d_arr_mul_16__26 (d_arr_mul_16__26), .d_arr_mul_16__25 (
               d_arr_mul_16__25), .d_arr_mul_16__24 (d_arr_mul_16__24), .d_arr_mul_16__23 (
               d_arr_mul_16__23), .d_arr_mul_16__22 (d_arr_mul_16__22), .d_arr_mul_16__21 (
               d_arr_mul_16__21), .d_arr_mul_16__20 (d_arr_mul_16__20), .d_arr_mul_16__19 (
               d_arr_mul_16__19), .d_arr_mul_16__18 (d_arr_mul_16__18), .d_arr_mul_16__17 (
               d_arr_mul_16__17), .d_arr_mul_16__16 (d_arr_mul_16__16), .d_arr_mul_16__15 (
               d_arr_mul_16__15), .d_arr_mul_16__14 (d_arr_mul_16__14), .d_arr_mul_16__13 (
               d_arr_mul_16__13), .d_arr_mul_16__12 (d_arr_mul_16__12), .d_arr_mul_16__11 (
               d_arr_mul_16__11), .d_arr_mul_16__10 (d_arr_mul_16__10), .d_arr_mul_16__9 (
               d_arr_mul_16__9), .d_arr_mul_16__8 (d_arr_mul_16__8), .d_arr_mul_16__7 (
               d_arr_mul_16__7), .d_arr_mul_16__6 (d_arr_mul_16__6), .d_arr_mul_16__5 (
               d_arr_mul_16__5), .d_arr_mul_16__4 (d_arr_mul_16__4), .d_arr_mul_16__3 (
               d_arr_mul_16__3), .d_arr_mul_16__2 (d_arr_mul_16__2), .d_arr_mul_16__1 (
               d_arr_mul_16__1), .d_arr_mul_16__0 (d_arr_mul_16__0), .d_arr_mul_17__31 (
               d_arr_mul_17__31), .d_arr_mul_17__30 (d_arr_mul_17__30), .d_arr_mul_17__29 (
               d_arr_mul_17__29), .d_arr_mul_17__28 (d_arr_mul_17__28), .d_arr_mul_17__27 (
               d_arr_mul_17__27), .d_arr_mul_17__26 (d_arr_mul_17__26), .d_arr_mul_17__25 (
               d_arr_mul_17__25), .d_arr_mul_17__24 (d_arr_mul_17__24), .d_arr_mul_17__23 (
               d_arr_mul_17__23), .d_arr_mul_17__22 (d_arr_mul_17__22), .d_arr_mul_17__21 (
               d_arr_mul_17__21), .d_arr_mul_17__20 (d_arr_mul_17__20), .d_arr_mul_17__19 (
               d_arr_mul_17__19), .d_arr_mul_17__18 (d_arr_mul_17__18), .d_arr_mul_17__17 (
               d_arr_mul_17__17), .d_arr_mul_17__16 (d_arr_mul_17__16), .d_arr_mul_17__15 (
               d_arr_mul_17__15), .d_arr_mul_17__14 (d_arr_mul_17__14), .d_arr_mul_17__13 (
               d_arr_mul_17__13), .d_arr_mul_17__12 (d_arr_mul_17__12), .d_arr_mul_17__11 (
               d_arr_mul_17__11), .d_arr_mul_17__10 (d_arr_mul_17__10), .d_arr_mul_17__9 (
               d_arr_mul_17__9), .d_arr_mul_17__8 (d_arr_mul_17__8), .d_arr_mul_17__7 (
               d_arr_mul_17__7), .d_arr_mul_17__6 (d_arr_mul_17__6), .d_arr_mul_17__5 (
               d_arr_mul_17__5), .d_arr_mul_17__4 (d_arr_mul_17__4), .d_arr_mul_17__3 (
               d_arr_mul_17__3), .d_arr_mul_17__2 (d_arr_mul_17__2), .d_arr_mul_17__1 (
               d_arr_mul_17__1), .d_arr_mul_17__0 (d_arr_mul_17__0), .d_arr_mul_18__31 (
               d_arr_mul_18__31), .d_arr_mul_18__30 (d_arr_mul_18__30), .d_arr_mul_18__29 (
               d_arr_mul_18__29), .d_arr_mul_18__28 (d_arr_mul_18__28), .d_arr_mul_18__27 (
               d_arr_mul_18__27), .d_arr_mul_18__26 (d_arr_mul_18__26), .d_arr_mul_18__25 (
               d_arr_mul_18__25), .d_arr_mul_18__24 (d_arr_mul_18__24), .d_arr_mul_18__23 (
               d_arr_mul_18__23), .d_arr_mul_18__22 (d_arr_mul_18__22), .d_arr_mul_18__21 (
               d_arr_mul_18__21), .d_arr_mul_18__20 (d_arr_mul_18__20), .d_arr_mul_18__19 (
               d_arr_mul_18__19), .d_arr_mul_18__18 (d_arr_mul_18__18), .d_arr_mul_18__17 (
               d_arr_mul_18__17), .d_arr_mul_18__16 (d_arr_mul_18__16), .d_arr_mul_18__15 (
               d_arr_mul_18__15), .d_arr_mul_18__14 (d_arr_mul_18__14), .d_arr_mul_18__13 (
               d_arr_mul_18__13), .d_arr_mul_18__12 (d_arr_mul_18__12), .d_arr_mul_18__11 (
               d_arr_mul_18__11), .d_arr_mul_18__10 (d_arr_mul_18__10), .d_arr_mul_18__9 (
               d_arr_mul_18__9), .d_arr_mul_18__8 (d_arr_mul_18__8), .d_arr_mul_18__7 (
               d_arr_mul_18__7), .d_arr_mul_18__6 (d_arr_mul_18__6), .d_arr_mul_18__5 (
               d_arr_mul_18__5), .d_arr_mul_18__4 (d_arr_mul_18__4), .d_arr_mul_18__3 (
               d_arr_mul_18__3), .d_arr_mul_18__2 (d_arr_mul_18__2), .d_arr_mul_18__1 (
               d_arr_mul_18__1), .d_arr_mul_18__0 (d_arr_mul_18__0), .d_arr_mul_19__31 (
               d_arr_mul_19__31), .d_arr_mul_19__30 (d_arr_mul_19__30), .d_arr_mul_19__29 (
               d_arr_mul_19__29), .d_arr_mul_19__28 (d_arr_mul_19__28), .d_arr_mul_19__27 (
               d_arr_mul_19__27), .d_arr_mul_19__26 (d_arr_mul_19__26), .d_arr_mul_19__25 (
               d_arr_mul_19__25), .d_arr_mul_19__24 (d_arr_mul_19__24), .d_arr_mul_19__23 (
               d_arr_mul_19__23), .d_arr_mul_19__22 (d_arr_mul_19__22), .d_arr_mul_19__21 (
               d_arr_mul_19__21), .d_arr_mul_19__20 (d_arr_mul_19__20), .d_arr_mul_19__19 (
               d_arr_mul_19__19), .d_arr_mul_19__18 (d_arr_mul_19__18), .d_arr_mul_19__17 (
               d_arr_mul_19__17), .d_arr_mul_19__16 (d_arr_mul_19__16), .d_arr_mul_19__15 (
               d_arr_mul_19__15), .d_arr_mul_19__14 (d_arr_mul_19__14), .d_arr_mul_19__13 (
               d_arr_mul_19__13), .d_arr_mul_19__12 (d_arr_mul_19__12), .d_arr_mul_19__11 (
               d_arr_mul_19__11), .d_arr_mul_19__10 (d_arr_mul_19__10), .d_arr_mul_19__9 (
               d_arr_mul_19__9), .d_arr_mul_19__8 (d_arr_mul_19__8), .d_arr_mul_19__7 (
               d_arr_mul_19__7), .d_arr_mul_19__6 (d_arr_mul_19__6), .d_arr_mul_19__5 (
               d_arr_mul_19__5), .d_arr_mul_19__4 (d_arr_mul_19__4), .d_arr_mul_19__3 (
               d_arr_mul_19__3), .d_arr_mul_19__2 (d_arr_mul_19__2), .d_arr_mul_19__1 (
               d_arr_mul_19__1), .d_arr_mul_19__0 (d_arr_mul_19__0), .d_arr_mul_20__31 (
               d_arr_mul_20__31), .d_arr_mul_20__30 (d_arr_mul_20__30), .d_arr_mul_20__29 (
               d_arr_mul_20__29), .d_arr_mul_20__28 (d_arr_mul_20__28), .d_arr_mul_20__27 (
               d_arr_mul_20__27), .d_arr_mul_20__26 (d_arr_mul_20__26), .d_arr_mul_20__25 (
               d_arr_mul_20__25), .d_arr_mul_20__24 (d_arr_mul_20__24), .d_arr_mul_20__23 (
               d_arr_mul_20__23), .d_arr_mul_20__22 (d_arr_mul_20__22), .d_arr_mul_20__21 (
               d_arr_mul_20__21), .d_arr_mul_20__20 (d_arr_mul_20__20), .d_arr_mul_20__19 (
               d_arr_mul_20__19), .d_arr_mul_20__18 (d_arr_mul_20__18), .d_arr_mul_20__17 (
               d_arr_mul_20__17), .d_arr_mul_20__16 (d_arr_mul_20__16), .d_arr_mul_20__15 (
               d_arr_mul_20__15), .d_arr_mul_20__14 (d_arr_mul_20__14), .d_arr_mul_20__13 (
               d_arr_mul_20__13), .d_arr_mul_20__12 (d_arr_mul_20__12), .d_arr_mul_20__11 (
               d_arr_mul_20__11), .d_arr_mul_20__10 (d_arr_mul_20__10), .d_arr_mul_20__9 (
               d_arr_mul_20__9), .d_arr_mul_20__8 (d_arr_mul_20__8), .d_arr_mul_20__7 (
               d_arr_mul_20__7), .d_arr_mul_20__6 (d_arr_mul_20__6), .d_arr_mul_20__5 (
               d_arr_mul_20__5), .d_arr_mul_20__4 (d_arr_mul_20__4), .d_arr_mul_20__3 (
               d_arr_mul_20__3), .d_arr_mul_20__2 (d_arr_mul_20__2), .d_arr_mul_20__1 (
               d_arr_mul_20__1), .d_arr_mul_20__0 (d_arr_mul_20__0), .d_arr_mul_21__31 (
               d_arr_mul_21__31), .d_arr_mul_21__30 (d_arr_mul_21__30), .d_arr_mul_21__29 (
               d_arr_mul_21__29), .d_arr_mul_21__28 (d_arr_mul_21__28), .d_arr_mul_21__27 (
               d_arr_mul_21__27), .d_arr_mul_21__26 (d_arr_mul_21__26), .d_arr_mul_21__25 (
               d_arr_mul_21__25), .d_arr_mul_21__24 (d_arr_mul_21__24), .d_arr_mul_21__23 (
               d_arr_mul_21__23), .d_arr_mul_21__22 (d_arr_mul_21__22), .d_arr_mul_21__21 (
               d_arr_mul_21__21), .d_arr_mul_21__20 (d_arr_mul_21__20), .d_arr_mul_21__19 (
               d_arr_mul_21__19), .d_arr_mul_21__18 (d_arr_mul_21__18), .d_arr_mul_21__17 (
               d_arr_mul_21__17), .d_arr_mul_21__16 (d_arr_mul_21__16), .d_arr_mul_21__15 (
               d_arr_mul_21__15), .d_arr_mul_21__14 (d_arr_mul_21__14), .d_arr_mul_21__13 (
               d_arr_mul_21__13), .d_arr_mul_21__12 (d_arr_mul_21__12), .d_arr_mul_21__11 (
               d_arr_mul_21__11), .d_arr_mul_21__10 (d_arr_mul_21__10), .d_arr_mul_21__9 (
               d_arr_mul_21__9), .d_arr_mul_21__8 (d_arr_mul_21__8), .d_arr_mul_21__7 (
               d_arr_mul_21__7), .d_arr_mul_21__6 (d_arr_mul_21__6), .d_arr_mul_21__5 (
               d_arr_mul_21__5), .d_arr_mul_21__4 (d_arr_mul_21__4), .d_arr_mul_21__3 (
               d_arr_mul_21__3), .d_arr_mul_21__2 (d_arr_mul_21__2), .d_arr_mul_21__1 (
               d_arr_mul_21__1), .d_arr_mul_21__0 (d_arr_mul_21__0), .d_arr_mul_22__31 (
               d_arr_mul_22__31), .d_arr_mul_22__30 (d_arr_mul_22__30), .d_arr_mul_22__29 (
               d_arr_mul_22__29), .d_arr_mul_22__28 (d_arr_mul_22__28), .d_arr_mul_22__27 (
               d_arr_mul_22__27), .d_arr_mul_22__26 (d_arr_mul_22__26), .d_arr_mul_22__25 (
               d_arr_mul_22__25), .d_arr_mul_22__24 (d_arr_mul_22__24), .d_arr_mul_22__23 (
               d_arr_mul_22__23), .d_arr_mul_22__22 (d_arr_mul_22__22), .d_arr_mul_22__21 (
               d_arr_mul_22__21), .d_arr_mul_22__20 (d_arr_mul_22__20), .d_arr_mul_22__19 (
               d_arr_mul_22__19), .d_arr_mul_22__18 (d_arr_mul_22__18), .d_arr_mul_22__17 (
               d_arr_mul_22__17), .d_arr_mul_22__16 (d_arr_mul_22__16), .d_arr_mul_22__15 (
               d_arr_mul_22__15), .d_arr_mul_22__14 (d_arr_mul_22__14), .d_arr_mul_22__13 (
               d_arr_mul_22__13), .d_arr_mul_22__12 (d_arr_mul_22__12), .d_arr_mul_22__11 (
               d_arr_mul_22__11), .d_arr_mul_22__10 (d_arr_mul_22__10), .d_arr_mul_22__9 (
               d_arr_mul_22__9), .d_arr_mul_22__8 (d_arr_mul_22__8), .d_arr_mul_22__7 (
               d_arr_mul_22__7), .d_arr_mul_22__6 (d_arr_mul_22__6), .d_arr_mul_22__5 (
               d_arr_mul_22__5), .d_arr_mul_22__4 (d_arr_mul_22__4), .d_arr_mul_22__3 (
               d_arr_mul_22__3), .d_arr_mul_22__2 (d_arr_mul_22__2), .d_arr_mul_22__1 (
               d_arr_mul_22__1), .d_arr_mul_22__0 (d_arr_mul_22__0), .d_arr_mul_23__31 (
               d_arr_mul_23__31), .d_arr_mul_23__30 (d_arr_mul_23__30), .d_arr_mul_23__29 (
               d_arr_mul_23__29), .d_arr_mul_23__28 (d_arr_mul_23__28), .d_arr_mul_23__27 (
               d_arr_mul_23__27), .d_arr_mul_23__26 (d_arr_mul_23__26), .d_arr_mul_23__25 (
               d_arr_mul_23__25), .d_arr_mul_23__24 (d_arr_mul_23__24), .d_arr_mul_23__23 (
               d_arr_mul_23__23), .d_arr_mul_23__22 (d_arr_mul_23__22), .d_arr_mul_23__21 (
               d_arr_mul_23__21), .d_arr_mul_23__20 (d_arr_mul_23__20), .d_arr_mul_23__19 (
               d_arr_mul_23__19), .d_arr_mul_23__18 (d_arr_mul_23__18), .d_arr_mul_23__17 (
               d_arr_mul_23__17), .d_arr_mul_23__16 (d_arr_mul_23__16), .d_arr_mul_23__15 (
               d_arr_mul_23__15), .d_arr_mul_23__14 (d_arr_mul_23__14), .d_arr_mul_23__13 (
               d_arr_mul_23__13), .d_arr_mul_23__12 (d_arr_mul_23__12), .d_arr_mul_23__11 (
               d_arr_mul_23__11), .d_arr_mul_23__10 (d_arr_mul_23__10), .d_arr_mul_23__9 (
               d_arr_mul_23__9), .d_arr_mul_23__8 (d_arr_mul_23__8), .d_arr_mul_23__7 (
               d_arr_mul_23__7), .d_arr_mul_23__6 (d_arr_mul_23__6), .d_arr_mul_23__5 (
               d_arr_mul_23__5), .d_arr_mul_23__4 (d_arr_mul_23__4), .d_arr_mul_23__3 (
               d_arr_mul_23__3), .d_arr_mul_23__2 (d_arr_mul_23__2), .d_arr_mul_23__1 (
               d_arr_mul_23__1), .d_arr_mul_23__0 (d_arr_mul_23__0), .d_arr_mul_24__31 (
               d_arr_mul_24__31), .d_arr_mul_24__30 (d_arr_mul_24__30), .d_arr_mul_24__29 (
               d_arr_mul_24__29), .d_arr_mul_24__28 (d_arr_mul_24__28), .d_arr_mul_24__27 (
               d_arr_mul_24__27), .d_arr_mul_24__26 (d_arr_mul_24__26), .d_arr_mul_24__25 (
               d_arr_mul_24__25), .d_arr_mul_24__24 (d_arr_mul_24__24), .d_arr_mul_24__23 (
               d_arr_mul_24__23), .d_arr_mul_24__22 (d_arr_mul_24__22), .d_arr_mul_24__21 (
               d_arr_mul_24__21), .d_arr_mul_24__20 (d_arr_mul_24__20), .d_arr_mul_24__19 (
               d_arr_mul_24__19), .d_arr_mul_24__18 (d_arr_mul_24__18), .d_arr_mul_24__17 (
               d_arr_mul_24__17), .d_arr_mul_24__16 (d_arr_mul_24__16), .d_arr_mul_24__15 (
               d_arr_mul_24__15), .d_arr_mul_24__14 (d_arr_mul_24__14), .d_arr_mul_24__13 (
               d_arr_mul_24__13), .d_arr_mul_24__12 (d_arr_mul_24__12), .d_arr_mul_24__11 (
               d_arr_mul_24__11), .d_arr_mul_24__10 (d_arr_mul_24__10), .d_arr_mul_24__9 (
               d_arr_mul_24__9), .d_arr_mul_24__8 (d_arr_mul_24__8), .d_arr_mul_24__7 (
               d_arr_mul_24__7), .d_arr_mul_24__6 (d_arr_mul_24__6), .d_arr_mul_24__5 (
               d_arr_mul_24__5), .d_arr_mul_24__4 (d_arr_mul_24__4), .d_arr_mul_24__3 (
               d_arr_mul_24__3), .d_arr_mul_24__2 (d_arr_mul_24__2), .d_arr_mul_24__1 (
               d_arr_mul_24__1), .d_arr_mul_24__0 (d_arr_mul_24__0), .d_arr_add_0__31 (
               d_arr_add_0__31), .d_arr_add_0__30 (d_arr_add_0__30), .d_arr_add_0__29 (
               d_arr_add_0__29), .d_arr_add_0__28 (d_arr_add_0__28), .d_arr_add_0__27 (
               d_arr_add_0__27), .d_arr_add_0__26 (d_arr_add_0__26), .d_arr_add_0__25 (
               d_arr_add_0__25), .d_arr_add_0__24 (d_arr_add_0__24), .d_arr_add_0__23 (
               d_arr_add_0__23), .d_arr_add_0__22 (d_arr_add_0__22), .d_arr_add_0__21 (
               d_arr_add_0__21), .d_arr_add_0__20 (d_arr_add_0__20), .d_arr_add_0__19 (
               d_arr_add_0__19), .d_arr_add_0__18 (d_arr_add_0__18), .d_arr_add_0__17 (
               d_arr_add_0__17), .d_arr_add_0__16 (d_arr_add_0__16), .d_arr_add_0__15 (
               d_arr_add_0__15), .d_arr_add_0__14 (d_arr_add_0__14), .d_arr_add_0__13 (
               d_arr_add_0__13), .d_arr_add_0__12 (d_arr_add_0__12), .d_arr_add_0__11 (
               d_arr_add_0__11), .d_arr_add_0__10 (d_arr_add_0__10), .d_arr_add_0__9 (
               d_arr_add_0__9), .d_arr_add_0__8 (d_arr_add_0__8), .d_arr_add_0__7 (
               d_arr_add_0__7), .d_arr_add_0__6 (d_arr_add_0__6), .d_arr_add_0__5 (
               d_arr_add_0__5), .d_arr_add_0__4 (d_arr_add_0__4), .d_arr_add_0__3 (
               d_arr_add_0__3), .d_arr_add_0__2 (d_arr_add_0__2), .d_arr_add_0__1 (
               d_arr_add_0__1), .d_arr_add_0__0 (d_arr_add_0__0), .d_arr_add_1__31 (
               d_arr_add_1__31), .d_arr_add_1__30 (d_arr_add_1__30), .d_arr_add_1__29 (
               d_arr_add_1__29), .d_arr_add_1__28 (d_arr_add_1__28), .d_arr_add_1__27 (
               d_arr_add_1__27), .d_arr_add_1__26 (d_arr_add_1__26), .d_arr_add_1__25 (
               d_arr_add_1__25), .d_arr_add_1__24 (d_arr_add_1__24), .d_arr_add_1__23 (
               d_arr_add_1__23), .d_arr_add_1__22 (d_arr_add_1__22), .d_arr_add_1__21 (
               d_arr_add_1__21), .d_arr_add_1__20 (d_arr_add_1__20), .d_arr_add_1__19 (
               d_arr_add_1__19), .d_arr_add_1__18 (d_arr_add_1__18), .d_arr_add_1__17 (
               d_arr_add_1__17), .d_arr_add_1__16 (d_arr_add_1__16), .d_arr_add_1__15 (
               d_arr_add_1__15), .d_arr_add_1__14 (d_arr_add_1__14), .d_arr_add_1__13 (
               d_arr_add_1__13), .d_arr_add_1__12 (d_arr_add_1__12), .d_arr_add_1__11 (
               d_arr_add_1__11), .d_arr_add_1__10 (d_arr_add_1__10), .d_arr_add_1__9 (
               d_arr_add_1__9), .d_arr_add_1__8 (d_arr_add_1__8), .d_arr_add_1__7 (
               d_arr_add_1__7), .d_arr_add_1__6 (d_arr_add_1__6), .d_arr_add_1__5 (
               d_arr_add_1__5), .d_arr_add_1__4 (d_arr_add_1__4), .d_arr_add_1__3 (
               d_arr_add_1__3), .d_arr_add_1__2 (d_arr_add_1__2), .d_arr_add_1__1 (
               d_arr_add_1__1), .d_arr_add_1__0 (d_arr_add_1__0), .d_arr_add_2__31 (
               d_arr_add_2__31), .d_arr_add_2__30 (d_arr_add_2__30), .d_arr_add_2__29 (
               d_arr_add_2__29), .d_arr_add_2__28 (d_arr_add_2__28), .d_arr_add_2__27 (
               d_arr_add_2__27), .d_arr_add_2__26 (d_arr_add_2__26), .d_arr_add_2__25 (
               d_arr_add_2__25), .d_arr_add_2__24 (d_arr_add_2__24), .d_arr_add_2__23 (
               d_arr_add_2__23), .d_arr_add_2__22 (d_arr_add_2__22), .d_arr_add_2__21 (
               d_arr_add_2__21), .d_arr_add_2__20 (d_arr_add_2__20), .d_arr_add_2__19 (
               d_arr_add_2__19), .d_arr_add_2__18 (d_arr_add_2__18), .d_arr_add_2__17 (
               d_arr_add_2__17), .d_arr_add_2__16 (d_arr_add_2__16), .d_arr_add_2__15 (
               d_arr_add_2__15), .d_arr_add_2__14 (d_arr_add_2__14), .d_arr_add_2__13 (
               d_arr_add_2__13), .d_arr_add_2__12 (d_arr_add_2__12), .d_arr_add_2__11 (
               d_arr_add_2__11), .d_arr_add_2__10 (d_arr_add_2__10), .d_arr_add_2__9 (
               d_arr_add_2__9), .d_arr_add_2__8 (d_arr_add_2__8), .d_arr_add_2__7 (
               d_arr_add_2__7), .d_arr_add_2__6 (d_arr_add_2__6), .d_arr_add_2__5 (
               d_arr_add_2__5), .d_arr_add_2__4 (d_arr_add_2__4), .d_arr_add_2__3 (
               d_arr_add_2__3), .d_arr_add_2__2 (d_arr_add_2__2), .d_arr_add_2__1 (
               d_arr_add_2__1), .d_arr_add_2__0 (d_arr_add_2__0), .d_arr_add_3__31 (
               d_arr_add_3__31), .d_arr_add_3__30 (d_arr_add_3__30), .d_arr_add_3__29 (
               d_arr_add_3__29), .d_arr_add_3__28 (d_arr_add_3__28), .d_arr_add_3__27 (
               d_arr_add_3__27), .d_arr_add_3__26 (d_arr_add_3__26), .d_arr_add_3__25 (
               d_arr_add_3__25), .d_arr_add_3__24 (d_arr_add_3__24), .d_arr_add_3__23 (
               d_arr_add_3__23), .d_arr_add_3__22 (d_arr_add_3__22), .d_arr_add_3__21 (
               d_arr_add_3__21), .d_arr_add_3__20 (d_arr_add_3__20), .d_arr_add_3__19 (
               d_arr_add_3__19), .d_arr_add_3__18 (d_arr_add_3__18), .d_arr_add_3__17 (
               d_arr_add_3__17), .d_arr_add_3__16 (d_arr_add_3__16), .d_arr_add_3__15 (
               d_arr_add_3__15), .d_arr_add_3__14 (d_arr_add_3__14), .d_arr_add_3__13 (
               d_arr_add_3__13), .d_arr_add_3__12 (d_arr_add_3__12), .d_arr_add_3__11 (
               d_arr_add_3__11), .d_arr_add_3__10 (d_arr_add_3__10), .d_arr_add_3__9 (
               d_arr_add_3__9), .d_arr_add_3__8 (d_arr_add_3__8), .d_arr_add_3__7 (
               d_arr_add_3__7), .d_arr_add_3__6 (d_arr_add_3__6), .d_arr_add_3__5 (
               d_arr_add_3__5), .d_arr_add_3__4 (d_arr_add_3__4), .d_arr_add_3__3 (
               d_arr_add_3__3), .d_arr_add_3__2 (d_arr_add_3__2), .d_arr_add_3__1 (
               d_arr_add_3__1), .d_arr_add_3__0 (d_arr_add_3__0), .d_arr_add_4__31 (
               q_arr_8__31), .d_arr_add_4__30 (q_arr_8__30), .d_arr_add_4__29 (
               q_arr_8__29), .d_arr_add_4__28 (q_arr_8__28), .d_arr_add_4__27 (
               q_arr_8__27), .d_arr_add_4__26 (q_arr_8__26), .d_arr_add_4__25 (
               q_arr_8__25), .d_arr_add_4__24 (q_arr_8__24), .d_arr_add_4__23 (
               q_arr_8__23), .d_arr_add_4__22 (q_arr_8__22), .d_arr_add_4__21 (
               q_arr_8__21), .d_arr_add_4__20 (q_arr_8__20), .d_arr_add_4__19 (
               q_arr_8__19), .d_arr_add_4__18 (q_arr_8__18), .d_arr_add_4__17 (
               q_arr_8__17), .d_arr_add_4__16 (q_arr_8__16), .d_arr_add_4__15 (
               q_arr_8__15), .d_arr_add_4__14 (q_arr_8__14), .d_arr_add_4__13 (
               q_arr_8__13), .d_arr_add_4__12 (q_arr_8__12), .d_arr_add_4__11 (
               q_arr_8__11), .d_arr_add_4__10 (q_arr_8__10), .d_arr_add_4__9 (
               q_arr_8__9), .d_arr_add_4__8 (q_arr_8__8), .d_arr_add_4__7 (
               q_arr_8__7), .d_arr_add_4__6 (q_arr_8__6), .d_arr_add_4__5 (
               q_arr_8__5), .d_arr_add_4__4 (q_arr_8__4), .d_arr_add_4__3 (
               q_arr_8__3), .d_arr_add_4__2 (q_arr_8__2), .d_arr_add_4__1 (
               q_arr_8__1), .d_arr_add_4__0 (q_arr_8__0), .d_arr_add_5__31 (GND0
               ), .d_arr_add_5__30 (GND0), .d_arr_add_5__29 (GND0), .d_arr_add_5__28 (
               GND0), .d_arr_add_5__27 (GND0), .d_arr_add_5__26 (GND0), .d_arr_add_5__25 (
               GND0), .d_arr_add_5__24 (GND0), .d_arr_add_5__23 (GND0), .d_arr_add_5__22 (
               GND0), .d_arr_add_5__21 (GND0), .d_arr_add_5__20 (GND0), .d_arr_add_5__19 (
               GND0), .d_arr_add_5__18 (GND0), .d_arr_add_5__17 (GND0), .d_arr_add_5__16 (
               GND0), .d_arr_add_5__15 (GND0), .d_arr_add_5__14 (GND0), .d_arr_add_5__13 (
               GND0), .d_arr_add_5__12 (GND0), .d_arr_add_5__11 (GND0), .d_arr_add_5__10 (
               GND0), .d_arr_add_5__9 (GND0), .d_arr_add_5__8 (GND0), .d_arr_add_5__7 (
               GND0), .d_arr_add_5__6 (GND0), .d_arr_add_5__5 (GND0), .d_arr_add_5__4 (
               GND0), .d_arr_add_5__3 (GND0), .d_arr_add_5__2 (GND0), .d_arr_add_5__1 (
               GND0), .d_arr_add_5__0 (GND0), .d_arr_add_6__31 (GND0), .d_arr_add_6__30 (
               GND0), .d_arr_add_6__29 (GND0), .d_arr_add_6__28 (GND0), .d_arr_add_6__27 (
               GND0), .d_arr_add_6__26 (GND0), .d_arr_add_6__25 (GND0), .d_arr_add_6__24 (
               GND0), .d_arr_add_6__23 (GND0), .d_arr_add_6__22 (GND0), .d_arr_add_6__21 (
               GND0), .d_arr_add_6__20 (GND0), .d_arr_add_6__19 (GND0), .d_arr_add_6__18 (
               GND0), .d_arr_add_6__17 (GND0), .d_arr_add_6__16 (GND0), .d_arr_add_6__15 (
               GND0), .d_arr_add_6__14 (GND0), .d_arr_add_6__13 (GND0), .d_arr_add_6__12 (
               GND0), .d_arr_add_6__11 (GND0), .d_arr_add_6__10 (GND0), .d_arr_add_6__9 (
               GND0), .d_arr_add_6__8 (GND0), .d_arr_add_6__7 (GND0), .d_arr_add_6__6 (
               GND0), .d_arr_add_6__5 (GND0), .d_arr_add_6__4 (GND0), .d_arr_add_6__3 (
               GND0), .d_arr_add_6__2 (GND0), .d_arr_add_6__1 (GND0), .d_arr_add_6__0 (
               GND0), .d_arr_add_7__31 (GND0), .d_arr_add_7__30 (GND0), .d_arr_add_7__29 (
               GND0), .d_arr_add_7__28 (GND0), .d_arr_add_7__27 (GND0), .d_arr_add_7__26 (
               GND0), .d_arr_add_7__25 (GND0), .d_arr_add_7__24 (GND0), .d_arr_add_7__23 (
               GND0), .d_arr_add_7__22 (GND0), .d_arr_add_7__21 (GND0), .d_arr_add_7__20 (
               GND0), .d_arr_add_7__19 (GND0), .d_arr_add_7__18 (GND0), .d_arr_add_7__17 (
               GND0), .d_arr_add_7__16 (GND0), .d_arr_add_7__15 (GND0), .d_arr_add_7__14 (
               GND0), .d_arr_add_7__13 (GND0), .d_arr_add_7__12 (GND0), .d_arr_add_7__11 (
               GND0), .d_arr_add_7__10 (GND0), .d_arr_add_7__9 (GND0), .d_arr_add_7__8 (
               GND0), .d_arr_add_7__7 (GND0), .d_arr_add_7__6 (GND0), .d_arr_add_7__5 (
               GND0), .d_arr_add_7__4 (GND0), .d_arr_add_7__3 (GND0), .d_arr_add_7__2 (
               GND0), .d_arr_add_7__1 (GND0), .d_arr_add_7__0 (GND0), .d_arr_add_8__31 (
               GND0), .d_arr_add_8__30 (GND0), .d_arr_add_8__29 (GND0), .d_arr_add_8__28 (
               GND0), .d_arr_add_8__27 (GND0), .d_arr_add_8__26 (GND0), .d_arr_add_8__25 (
               GND0), .d_arr_add_8__24 (GND0), .d_arr_add_8__23 (GND0), .d_arr_add_8__22 (
               GND0), .d_arr_add_8__21 (GND0), .d_arr_add_8__20 (GND0), .d_arr_add_8__19 (
               GND0), .d_arr_add_8__18 (GND0), .d_arr_add_8__17 (GND0), .d_arr_add_8__16 (
               GND0), .d_arr_add_8__15 (GND0), .d_arr_add_8__14 (GND0), .d_arr_add_8__13 (
               GND0), .d_arr_add_8__12 (GND0), .d_arr_add_8__11 (GND0), .d_arr_add_8__10 (
               GND0), .d_arr_add_8__9 (GND0), .d_arr_add_8__8 (GND0), .d_arr_add_8__7 (
               GND0), .d_arr_add_8__6 (GND0), .d_arr_add_8__5 (GND0), .d_arr_add_8__4 (
               GND0), .d_arr_add_8__3 (GND0), .d_arr_add_8__2 (GND0), .d_arr_add_8__1 (
               GND0), .d_arr_add_8__0 (GND0), .d_arr_add_9__31 (d_arr_add_9__31)
               , .d_arr_add_9__30 (d_arr_add_9__30), .d_arr_add_9__29 (
               d_arr_add_9__29), .d_arr_add_9__28 (d_arr_add_9__28), .d_arr_add_9__27 (
               d_arr_add_9__27), .d_arr_add_9__26 (d_arr_add_9__26), .d_arr_add_9__25 (
               d_arr_add_9__25), .d_arr_add_9__24 (d_arr_add_9__24), .d_arr_add_9__23 (
               d_arr_add_9__23), .d_arr_add_9__22 (d_arr_add_9__22), .d_arr_add_9__21 (
               d_arr_add_9__21), .d_arr_add_9__20 (d_arr_add_9__20), .d_arr_add_9__19 (
               d_arr_add_9__19), .d_arr_add_9__18 (d_arr_add_9__18), .d_arr_add_9__17 (
               d_arr_add_9__17), .d_arr_add_9__16 (d_arr_add_9__16), .d_arr_add_9__15 (
               d_arr_add_9__15), .d_arr_add_9__14 (d_arr_add_9__14), .d_arr_add_9__13 (
               d_arr_add_9__13), .d_arr_add_9__12 (d_arr_add_9__12), .d_arr_add_9__11 (
               d_arr_add_9__11), .d_arr_add_9__10 (d_arr_add_9__10), .d_arr_add_9__9 (
               d_arr_add_9__9), .d_arr_add_9__8 (d_arr_add_9__8), .d_arr_add_9__7 (
               d_arr_add_9__7), .d_arr_add_9__6 (d_arr_add_9__6), .d_arr_add_9__5 (
               d_arr_add_9__5), .d_arr_add_9__4 (d_arr_add_9__4), .d_arr_add_9__3 (
               d_arr_add_9__3), .d_arr_add_9__2 (d_arr_add_9__2), .d_arr_add_9__1 (
               d_arr_add_9__1), .d_arr_add_9__0 (d_arr_add_9__0), .d_arr_add_10__31 (
               d_arr_add_10__31), .d_arr_add_10__30 (d_arr_add_10__30), .d_arr_add_10__29 (
               d_arr_add_10__29), .d_arr_add_10__28 (d_arr_add_10__28), .d_arr_add_10__27 (
               d_arr_add_10__27), .d_arr_add_10__26 (d_arr_add_10__26), .d_arr_add_10__25 (
               d_arr_add_10__25), .d_arr_add_10__24 (d_arr_add_10__24), .d_arr_add_10__23 (
               d_arr_add_10__23), .d_arr_add_10__22 (d_arr_add_10__22), .d_arr_add_10__21 (
               d_arr_add_10__21), .d_arr_add_10__20 (d_arr_add_10__20), .d_arr_add_10__19 (
               d_arr_add_10__19), .d_arr_add_10__18 (d_arr_add_10__18), .d_arr_add_10__17 (
               d_arr_add_10__17), .d_arr_add_10__16 (d_arr_add_10__16), .d_arr_add_10__15 (
               d_arr_add_10__15), .d_arr_add_10__14 (d_arr_add_10__14), .d_arr_add_10__13 (
               d_arr_add_10__13), .d_arr_add_10__12 (d_arr_add_10__12), .d_arr_add_10__11 (
               d_arr_add_10__11), .d_arr_add_10__10 (d_arr_add_10__10), .d_arr_add_10__9 (
               d_arr_add_10__9), .d_arr_add_10__8 (d_arr_add_10__8), .d_arr_add_10__7 (
               d_arr_add_10__7), .d_arr_add_10__6 (d_arr_add_10__6), .d_arr_add_10__5 (
               d_arr_add_10__5), .d_arr_add_10__4 (d_arr_add_10__4), .d_arr_add_10__3 (
               d_arr_add_10__3), .d_arr_add_10__2 (d_arr_add_10__2), .d_arr_add_10__1 (
               d_arr_add_10__1), .d_arr_add_10__0 (d_arr_add_10__0), .d_arr_add_11__31 (
               d_arr_add_11__31), .d_arr_add_11__30 (d_arr_add_11__30), .d_arr_add_11__29 (
               d_arr_add_11__29), .d_arr_add_11__28 (d_arr_add_11__28), .d_arr_add_11__27 (
               d_arr_add_11__27), .d_arr_add_11__26 (d_arr_add_11__26), .d_arr_add_11__25 (
               d_arr_add_11__25), .d_arr_add_11__24 (d_arr_add_11__24), .d_arr_add_11__23 (
               d_arr_add_11__23), .d_arr_add_11__22 (d_arr_add_11__22), .d_arr_add_11__21 (
               d_arr_add_11__21), .d_arr_add_11__20 (d_arr_add_11__20), .d_arr_add_11__19 (
               d_arr_add_11__19), .d_arr_add_11__18 (d_arr_add_11__18), .d_arr_add_11__17 (
               d_arr_add_11__17), .d_arr_add_11__16 (d_arr_add_11__16), .d_arr_add_11__15 (
               d_arr_add_11__15), .d_arr_add_11__14 (d_arr_add_11__14), .d_arr_add_11__13 (
               d_arr_add_11__13), .d_arr_add_11__12 (d_arr_add_11__12), .d_arr_add_11__11 (
               d_arr_add_11__11), .d_arr_add_11__10 (d_arr_add_11__10), .d_arr_add_11__9 (
               d_arr_add_11__9), .d_arr_add_11__8 (d_arr_add_11__8), .d_arr_add_11__7 (
               d_arr_add_11__7), .d_arr_add_11__6 (d_arr_add_11__6), .d_arr_add_11__5 (
               d_arr_add_11__5), .d_arr_add_11__4 (d_arr_add_11__4), .d_arr_add_11__3 (
               d_arr_add_11__3), .d_arr_add_11__2 (d_arr_add_11__2), .d_arr_add_11__1 (
               d_arr_add_11__1), .d_arr_add_11__0 (d_arr_add_11__0), .d_arr_add_12__31 (
               d_arr_add_12__31), .d_arr_add_12__30 (d_arr_add_12__30), .d_arr_add_12__29 (
               d_arr_add_12__29), .d_arr_add_12__28 (d_arr_add_12__28), .d_arr_add_12__27 (
               d_arr_add_12__27), .d_arr_add_12__26 (d_arr_add_12__26), .d_arr_add_12__25 (
               d_arr_add_12__25), .d_arr_add_12__24 (d_arr_add_12__24), .d_arr_add_12__23 (
               d_arr_add_12__23), .d_arr_add_12__22 (d_arr_add_12__22), .d_arr_add_12__21 (
               d_arr_add_12__21), .d_arr_add_12__20 (d_arr_add_12__20), .d_arr_add_12__19 (
               d_arr_add_12__19), .d_arr_add_12__18 (d_arr_add_12__18), .d_arr_add_12__17 (
               d_arr_add_12__17), .d_arr_add_12__16 (d_arr_add_12__16), .d_arr_add_12__15 (
               d_arr_add_12__15), .d_arr_add_12__14 (d_arr_add_12__14), .d_arr_add_12__13 (
               d_arr_add_12__13), .d_arr_add_12__12 (d_arr_add_12__12), .d_arr_add_12__11 (
               d_arr_add_12__11), .d_arr_add_12__10 (d_arr_add_12__10), .d_arr_add_12__9 (
               d_arr_add_12__9), .d_arr_add_12__8 (d_arr_add_12__8), .d_arr_add_12__7 (
               d_arr_add_12__7), .d_arr_add_12__6 (d_arr_add_12__6), .d_arr_add_12__5 (
               d_arr_add_12__5), .d_arr_add_12__4 (d_arr_add_12__4), .d_arr_add_12__3 (
               d_arr_add_12__3), .d_arr_add_12__2 (d_arr_add_12__2), .d_arr_add_12__1 (
               d_arr_add_12__1), .d_arr_add_12__0 (d_arr_add_12__0), .d_arr_add_13__31 (
               q_arr_17__31), .d_arr_add_13__30 (q_arr_17__30), .d_arr_add_13__29 (
               q_arr_17__29), .d_arr_add_13__28 (q_arr_17__28), .d_arr_add_13__27 (
               q_arr_17__27), .d_arr_add_13__26 (q_arr_17__26), .d_arr_add_13__25 (
               q_arr_17__25), .d_arr_add_13__24 (q_arr_17__24), .d_arr_add_13__23 (
               q_arr_17__23), .d_arr_add_13__22 (q_arr_17__22), .d_arr_add_13__21 (
               q_arr_17__21), .d_arr_add_13__20 (q_arr_17__20), .d_arr_add_13__19 (
               q_arr_17__19), .d_arr_add_13__18 (q_arr_17__18), .d_arr_add_13__17 (
               q_arr_17__17), .d_arr_add_13__16 (q_arr_17__16), .d_arr_add_13__15 (
               q_arr_17__15), .d_arr_add_13__14 (q_arr_17__14), .d_arr_add_13__13 (
               q_arr_17__13), .d_arr_add_13__12 (q_arr_17__12), .d_arr_add_13__11 (
               q_arr_17__11), .d_arr_add_13__10 (q_arr_17__10), .d_arr_add_13__9 (
               q_arr_17__9), .d_arr_add_13__8 (q_arr_17__8), .d_arr_add_13__7 (
               q_arr_17__7), .d_arr_add_13__6 (q_arr_17__6), .d_arr_add_13__5 (
               q_arr_17__5), .d_arr_add_13__4 (q_arr_17__4), .d_arr_add_13__3 (
               q_arr_17__3), .d_arr_add_13__2 (q_arr_17__2), .d_arr_add_13__1 (
               q_arr_17__1), .d_arr_add_13__0 (q_arr_17__0), .d_arr_add_14__31 (
               GND0), .d_arr_add_14__30 (GND0), .d_arr_add_14__29 (GND0), .d_arr_add_14__28 (
               GND0), .d_arr_add_14__27 (GND0), .d_arr_add_14__26 (GND0), .d_arr_add_14__25 (
               GND0), .d_arr_add_14__24 (GND0), .d_arr_add_14__23 (GND0), .d_arr_add_14__22 (
               GND0), .d_arr_add_14__21 (GND0), .d_arr_add_14__20 (GND0), .d_arr_add_14__19 (
               GND0), .d_arr_add_14__18 (GND0), .d_arr_add_14__17 (GND0), .d_arr_add_14__16 (
               GND0), .d_arr_add_14__15 (GND0), .d_arr_add_14__14 (GND0), .d_arr_add_14__13 (
               GND0), .d_arr_add_14__12 (GND0), .d_arr_add_14__11 (GND0), .d_arr_add_14__10 (
               GND0), .d_arr_add_14__9 (GND0), .d_arr_add_14__8 (GND0), .d_arr_add_14__7 (
               GND0), .d_arr_add_14__6 (GND0), .d_arr_add_14__5 (GND0), .d_arr_add_14__4 (
               GND0), .d_arr_add_14__3 (GND0), .d_arr_add_14__2 (GND0), .d_arr_add_14__1 (
               GND0), .d_arr_add_14__0 (GND0), .d_arr_add_15__31 (GND0), .d_arr_add_15__30 (
               GND0), .d_arr_add_15__29 (GND0), .d_arr_add_15__28 (GND0), .d_arr_add_15__27 (
               GND0), .d_arr_add_15__26 (GND0), .d_arr_add_15__25 (GND0), .d_arr_add_15__24 (
               GND0), .d_arr_add_15__23 (GND0), .d_arr_add_15__22 (GND0), .d_arr_add_15__21 (
               GND0), .d_arr_add_15__20 (GND0), .d_arr_add_15__19 (GND0), .d_arr_add_15__18 (
               GND0), .d_arr_add_15__17 (GND0), .d_arr_add_15__16 (GND0), .d_arr_add_15__15 (
               GND0), .d_arr_add_15__14 (GND0), .d_arr_add_15__13 (GND0), .d_arr_add_15__12 (
               GND0), .d_arr_add_15__11 (GND0), .d_arr_add_15__10 (GND0), .d_arr_add_15__9 (
               GND0), .d_arr_add_15__8 (GND0), .d_arr_add_15__7 (GND0), .d_arr_add_15__6 (
               GND0), .d_arr_add_15__5 (GND0), .d_arr_add_15__4 (GND0), .d_arr_add_15__3 (
               GND0), .d_arr_add_15__2 (GND0), .d_arr_add_15__1 (GND0), .d_arr_add_15__0 (
               GND0), .d_arr_add_16__31 (GND0), .d_arr_add_16__30 (GND0), .d_arr_add_16__29 (
               GND0), .d_arr_add_16__28 (GND0), .d_arr_add_16__27 (GND0), .d_arr_add_16__26 (
               GND0), .d_arr_add_16__25 (GND0), .d_arr_add_16__24 (GND0), .d_arr_add_16__23 (
               GND0), .d_arr_add_16__22 (GND0), .d_arr_add_16__21 (GND0), .d_arr_add_16__20 (
               GND0), .d_arr_add_16__19 (GND0), .d_arr_add_16__18 (GND0), .d_arr_add_16__17 (
               GND0), .d_arr_add_16__16 (GND0), .d_arr_add_16__15 (GND0), .d_arr_add_16__14 (
               GND0), .d_arr_add_16__13 (GND0), .d_arr_add_16__12 (GND0), .d_arr_add_16__11 (
               GND0), .d_arr_add_16__10 (GND0), .d_arr_add_16__9 (GND0), .d_arr_add_16__8 (
               GND0), .d_arr_add_16__7 (GND0), .d_arr_add_16__6 (GND0), .d_arr_add_16__5 (
               GND0), .d_arr_add_16__4 (GND0), .d_arr_add_16__3 (GND0), .d_arr_add_16__2 (
               GND0), .d_arr_add_16__1 (GND0), .d_arr_add_16__0 (GND0), .d_arr_add_17__31 (
               GND0), .d_arr_add_17__30 (GND0), .d_arr_add_17__29 (GND0), .d_arr_add_17__28 (
               GND0), .d_arr_add_17__27 (GND0), .d_arr_add_17__26 (GND0), .d_arr_add_17__25 (
               GND0), .d_arr_add_17__24 (GND0), .d_arr_add_17__23 (GND0), .d_arr_add_17__22 (
               GND0), .d_arr_add_17__21 (GND0), .d_arr_add_17__20 (GND0), .d_arr_add_17__19 (
               GND0), .d_arr_add_17__18 (GND0), .d_arr_add_17__17 (GND0), .d_arr_add_17__16 (
               GND0), .d_arr_add_17__15 (GND0), .d_arr_add_17__14 (GND0), .d_arr_add_17__13 (
               GND0), .d_arr_add_17__12 (GND0), .d_arr_add_17__11 (GND0), .d_arr_add_17__10 (
               GND0), .d_arr_add_17__9 (GND0), .d_arr_add_17__8 (GND0), .d_arr_add_17__7 (
               GND0), .d_arr_add_17__6 (GND0), .d_arr_add_17__5 (GND0), .d_arr_add_17__4 (
               GND0), .d_arr_add_17__3 (GND0), .d_arr_add_17__2 (GND0), .d_arr_add_17__1 (
               GND0), .d_arr_add_17__0 (GND0), .d_arr_add_18__31 (
               d_arr_add_18__31), .d_arr_add_18__30 (d_arr_add_18__30), .d_arr_add_18__29 (
               d_arr_add_18__29), .d_arr_add_18__28 (d_arr_add_18__28), .d_arr_add_18__27 (
               d_arr_add_18__27), .d_arr_add_18__26 (d_arr_add_18__26), .d_arr_add_18__25 (
               d_arr_add_18__25), .d_arr_add_18__24 (d_arr_add_18__24), .d_arr_add_18__23 (
               d_arr_add_18__23), .d_arr_add_18__22 (d_arr_add_18__22), .d_arr_add_18__21 (
               d_arr_add_18__21), .d_arr_add_18__20 (d_arr_add_18__20), .d_arr_add_18__19 (
               d_arr_add_18__19), .d_arr_add_18__18 (d_arr_add_18__18), .d_arr_add_18__17 (
               d_arr_add_18__17), .d_arr_add_18__16 (d_arr_add_18__16), .d_arr_add_18__15 (
               d_arr_add_18__15), .d_arr_add_18__14 (d_arr_add_18__14), .d_arr_add_18__13 (
               d_arr_add_18__13), .d_arr_add_18__12 (d_arr_add_18__12), .d_arr_add_18__11 (
               d_arr_add_18__11), .d_arr_add_18__10 (d_arr_add_18__10), .d_arr_add_18__9 (
               d_arr_add_18__9), .d_arr_add_18__8 (d_arr_add_18__8), .d_arr_add_18__7 (
               d_arr_add_18__7), .d_arr_add_18__6 (d_arr_add_18__6), .d_arr_add_18__5 (
               d_arr_add_18__5), .d_arr_add_18__4 (d_arr_add_18__4), .d_arr_add_18__3 (
               d_arr_add_18__3), .d_arr_add_18__2 (d_arr_add_18__2), .d_arr_add_18__1 (
               d_arr_add_18__1), .d_arr_add_18__0 (d_arr_add_18__0), .d_arr_add_19__31 (
               d_arr_add_19__31), .d_arr_add_19__30 (d_arr_add_19__30), .d_arr_add_19__29 (
               d_arr_add_19__29), .d_arr_add_19__28 (d_arr_add_19__28), .d_arr_add_19__27 (
               d_arr_add_19__27), .d_arr_add_19__26 (d_arr_add_19__26), .d_arr_add_19__25 (
               d_arr_add_19__25), .d_arr_add_19__24 (d_arr_add_19__24), .d_arr_add_19__23 (
               d_arr_add_19__23), .d_arr_add_19__22 (d_arr_add_19__22), .d_arr_add_19__21 (
               d_arr_add_19__21), .d_arr_add_19__20 (d_arr_add_19__20), .d_arr_add_19__19 (
               d_arr_add_19__19), .d_arr_add_19__18 (d_arr_add_19__18), .d_arr_add_19__17 (
               d_arr_add_19__17), .d_arr_add_19__16 (d_arr_add_19__16), .d_arr_add_19__15 (
               d_arr_add_19__15), .d_arr_add_19__14 (d_arr_add_19__14), .d_arr_add_19__13 (
               d_arr_add_19__13), .d_arr_add_19__12 (d_arr_add_19__12), .d_arr_add_19__11 (
               d_arr_add_19__11), .d_arr_add_19__10 (d_arr_add_19__10), .d_arr_add_19__9 (
               d_arr_add_19__9), .d_arr_add_19__8 (d_arr_add_19__8), .d_arr_add_19__7 (
               d_arr_add_19__7), .d_arr_add_19__6 (d_arr_add_19__6), .d_arr_add_19__5 (
               d_arr_add_19__5), .d_arr_add_19__4 (d_arr_add_19__4), .d_arr_add_19__3 (
               d_arr_add_19__3), .d_arr_add_19__2 (d_arr_add_19__2), .d_arr_add_19__1 (
               d_arr_add_19__1), .d_arr_add_19__0 (d_arr_add_19__0), .d_arr_add_20__31 (
               d_arr_add_20__31), .d_arr_add_20__30 (d_arr_add_20__30), .d_arr_add_20__29 (
               d_arr_add_20__29), .d_arr_add_20__28 (d_arr_add_20__28), .d_arr_add_20__27 (
               d_arr_add_20__27), .d_arr_add_20__26 (d_arr_add_20__26), .d_arr_add_20__25 (
               d_arr_add_20__25), .d_arr_add_20__24 (d_arr_add_20__24), .d_arr_add_20__23 (
               d_arr_add_20__23), .d_arr_add_20__22 (d_arr_add_20__22), .d_arr_add_20__21 (
               d_arr_add_20__21), .d_arr_add_20__20 (d_arr_add_20__20), .d_arr_add_20__19 (
               d_arr_add_20__19), .d_arr_add_20__18 (d_arr_add_20__18), .d_arr_add_20__17 (
               d_arr_add_20__17), .d_arr_add_20__16 (d_arr_add_20__16), .d_arr_add_20__15 (
               d_arr_add_20__15), .d_arr_add_20__14 (d_arr_add_20__14), .d_arr_add_20__13 (
               d_arr_add_20__13), .d_arr_add_20__12 (d_arr_add_20__12), .d_arr_add_20__11 (
               d_arr_add_20__11), .d_arr_add_20__10 (d_arr_add_20__10), .d_arr_add_20__9 (
               d_arr_add_20__9), .d_arr_add_20__8 (d_arr_add_20__8), .d_arr_add_20__7 (
               d_arr_add_20__7), .d_arr_add_20__6 (d_arr_add_20__6), .d_arr_add_20__5 (
               d_arr_add_20__5), .d_arr_add_20__4 (d_arr_add_20__4), .d_arr_add_20__3 (
               d_arr_add_20__3), .d_arr_add_20__2 (d_arr_add_20__2), .d_arr_add_20__1 (
               d_arr_add_20__1), .d_arr_add_20__0 (d_arr_add_20__0), .d_arr_add_21__31 (
               q_arr_24__31), .d_arr_add_21__30 (q_arr_24__30), .d_arr_add_21__29 (
               q_arr_24__29), .d_arr_add_21__28 (q_arr_24__28), .d_arr_add_21__27 (
               q_arr_24__27), .d_arr_add_21__26 (q_arr_24__26), .d_arr_add_21__25 (
               q_arr_24__25), .d_arr_add_21__24 (q_arr_24__24), .d_arr_add_21__23 (
               q_arr_24__23), .d_arr_add_21__22 (q_arr_24__22), .d_arr_add_21__21 (
               q_arr_24__21), .d_arr_add_21__20 (q_arr_24__20), .d_arr_add_21__19 (
               q_arr_24__19), .d_arr_add_21__18 (q_arr_24__18), .d_arr_add_21__17 (
               q_arr_24__17), .d_arr_add_21__16 (q_arr_24__16), .d_arr_add_21__15 (
               q_arr_24__15), .d_arr_add_21__14 (q_arr_24__14), .d_arr_add_21__13 (
               q_arr_24__13), .d_arr_add_21__12 (q_arr_24__12), .d_arr_add_21__11 (
               q_arr_24__11), .d_arr_add_21__10 (q_arr_24__10), .d_arr_add_21__9 (
               q_arr_24__9), .d_arr_add_21__8 (q_arr_24__8), .d_arr_add_21__7 (
               q_arr_24__7), .d_arr_add_21__6 (q_arr_24__6), .d_arr_add_21__5 (
               q_arr_24__5), .d_arr_add_21__4 (q_arr_24__4), .d_arr_add_21__3 (
               q_arr_24__3), .d_arr_add_21__2 (q_arr_24__2), .d_arr_add_21__1 (
               q_arr_24__1), .d_arr_add_21__0 (q_arr_24__0), .d_arr_add_22__31 (
               GND0), .d_arr_add_22__30 (GND0), .d_arr_add_22__29 (GND0), .d_arr_add_22__28 (
               GND0), .d_arr_add_22__27 (GND0), .d_arr_add_22__26 (GND0), .d_arr_add_22__25 (
               GND0), .d_arr_add_22__24 (GND0), .d_arr_add_22__23 (GND0), .d_arr_add_22__22 (
               GND0), .d_arr_add_22__21 (GND0), .d_arr_add_22__20 (GND0), .d_arr_add_22__19 (
               GND0), .d_arr_add_22__18 (GND0), .d_arr_add_22__17 (GND0), .d_arr_add_22__16 (
               GND0), .d_arr_add_22__15 (GND0), .d_arr_add_22__14 (GND0), .d_arr_add_22__13 (
               GND0), .d_arr_add_22__12 (GND0), .d_arr_add_22__11 (GND0), .d_arr_add_22__10 (
               GND0), .d_arr_add_22__9 (GND0), .d_arr_add_22__8 (GND0), .d_arr_add_22__7 (
               GND0), .d_arr_add_22__6 (GND0), .d_arr_add_22__5 (GND0), .d_arr_add_22__4 (
               GND0), .d_arr_add_22__3 (GND0), .d_arr_add_22__2 (GND0), .d_arr_add_22__1 (
               GND0), .d_arr_add_22__0 (GND0), .d_arr_add_23__31 (GND0), .d_arr_add_23__30 (
               GND0), .d_arr_add_23__29 (GND0), .d_arr_add_23__28 (GND0), .d_arr_add_23__27 (
               GND0), .d_arr_add_23__26 (GND0), .d_arr_add_23__25 (GND0), .d_arr_add_23__24 (
               GND0), .d_arr_add_23__23 (GND0), .d_arr_add_23__22 (GND0), .d_arr_add_23__21 (
               GND0), .d_arr_add_23__20 (GND0), .d_arr_add_23__19 (GND0), .d_arr_add_23__18 (
               GND0), .d_arr_add_23__17 (GND0), .d_arr_add_23__16 (GND0), .d_arr_add_23__15 (
               GND0), .d_arr_add_23__14 (GND0), .d_arr_add_23__13 (GND0), .d_arr_add_23__12 (
               GND0), .d_arr_add_23__11 (GND0), .d_arr_add_23__10 (GND0), .d_arr_add_23__9 (
               GND0), .d_arr_add_23__8 (GND0), .d_arr_add_23__7 (GND0), .d_arr_add_23__6 (
               GND0), .d_arr_add_23__5 (GND0), .d_arr_add_23__4 (GND0), .d_arr_add_23__3 (
               GND0), .d_arr_add_23__2 (GND0), .d_arr_add_23__1 (GND0), .d_arr_add_23__0 (
               GND0), .d_arr_add_24__31 (GND0), .d_arr_add_24__30 (GND0), .d_arr_add_24__29 (
               GND0), .d_arr_add_24__28 (GND0), .d_arr_add_24__27 (GND0), .d_arr_add_24__26 (
               GND0), .d_arr_add_24__25 (GND0), .d_arr_add_24__24 (GND0), .d_arr_add_24__23 (
               GND0), .d_arr_add_24__22 (GND0), .d_arr_add_24__21 (GND0), .d_arr_add_24__20 (
               GND0), .d_arr_add_24__19 (GND0), .d_arr_add_24__18 (GND0), .d_arr_add_24__17 (
               GND0), .d_arr_add_24__16 (GND0), .d_arr_add_24__15 (GND0), .d_arr_add_24__14 (
               GND0), .d_arr_add_24__13 (GND0), .d_arr_add_24__12 (GND0), .d_arr_add_24__11 (
               GND0), .d_arr_add_24__10 (GND0), .d_arr_add_24__9 (GND0), .d_arr_add_24__8 (
               GND0), .d_arr_add_24__7 (GND0), .d_arr_add_24__6 (GND0), .d_arr_add_24__5 (
               GND0), .d_arr_add_24__4 (GND0), .d_arr_add_24__3 (GND0), .d_arr_add_24__2 (
               GND0), .d_arr_add_24__1 (GND0), .d_arr_add_24__0 (GND0), .d_arr_merge1_0__31 (
               d_arr_merge1_0__31), .d_arr_merge1_0__30 (d_arr_merge1_0__30), .d_arr_merge1_0__29 (
               d_arr_merge1_0__29), .d_arr_merge1_0__28 (d_arr_merge1_0__28), .d_arr_merge1_0__27 (
               d_arr_merge1_0__27), .d_arr_merge1_0__26 (d_arr_merge1_0__26), .d_arr_merge1_0__25 (
               d_arr_merge1_0__25), .d_arr_merge1_0__24 (d_arr_merge1_0__24), .d_arr_merge1_0__23 (
               d_arr_merge1_0__23), .d_arr_merge1_0__22 (d_arr_merge1_0__22), .d_arr_merge1_0__21 (
               d_arr_merge1_0__21), .d_arr_merge1_0__20 (d_arr_merge1_0__20), .d_arr_merge1_0__19 (
               d_arr_merge1_0__19), .d_arr_merge1_0__18 (d_arr_merge1_0__18), .d_arr_merge1_0__17 (
               d_arr_merge1_0__17), .d_arr_merge1_0__16 (d_arr_merge1_0__16), .d_arr_merge1_0__15 (
               d_arr_merge1_0__15), .d_arr_merge1_0__14 (d_arr_merge1_0__14), .d_arr_merge1_0__13 (
               d_arr_merge1_0__13), .d_arr_merge1_0__12 (d_arr_merge1_0__12), .d_arr_merge1_0__11 (
               d_arr_merge1_0__11), .d_arr_merge1_0__10 (d_arr_merge1_0__10), .d_arr_merge1_0__9 (
               d_arr_merge1_0__9), .d_arr_merge1_0__8 (d_arr_merge1_0__8), .d_arr_merge1_0__7 (
               d_arr_merge1_0__7), .d_arr_merge1_0__6 (d_arr_merge1_0__6), .d_arr_merge1_0__5 (
               d_arr_merge1_0__5), .d_arr_merge1_0__4 (d_arr_merge1_0__4), .d_arr_merge1_0__3 (
               d_arr_merge1_0__3), .d_arr_merge1_0__2 (d_arr_merge1_0__2), .d_arr_merge1_0__1 (
               d_arr_merge1_0__1), .d_arr_merge1_0__0 (d_arr_merge1_0__0), .d_arr_merge1_1__31 (
               d_arr_merge1_1__31), .d_arr_merge1_1__30 (d_arr_merge1_1__30), .d_arr_merge1_1__29 (
               d_arr_merge1_1__29), .d_arr_merge1_1__28 (d_arr_merge1_1__28), .d_arr_merge1_1__27 (
               d_arr_merge1_1__27), .d_arr_merge1_1__26 (d_arr_merge1_1__26), .d_arr_merge1_1__25 (
               d_arr_merge1_1__25), .d_arr_merge1_1__24 (d_arr_merge1_1__24), .d_arr_merge1_1__23 (
               d_arr_merge1_1__23), .d_arr_merge1_1__22 (d_arr_merge1_1__22), .d_arr_merge1_1__21 (
               d_arr_merge1_1__21), .d_arr_merge1_1__20 (d_arr_merge1_1__20), .d_arr_merge1_1__19 (
               d_arr_merge1_1__19), .d_arr_merge1_1__18 (d_arr_merge1_1__18), .d_arr_merge1_1__17 (
               d_arr_merge1_1__17), .d_arr_merge1_1__16 (d_arr_merge1_1__16), .d_arr_merge1_1__15 (
               d_arr_merge1_1__15), .d_arr_merge1_1__14 (d_arr_merge1_1__14), .d_arr_merge1_1__13 (
               d_arr_merge1_1__13), .d_arr_merge1_1__12 (d_arr_merge1_1__12), .d_arr_merge1_1__11 (
               d_arr_merge1_1__11), .d_arr_merge1_1__10 (d_arr_merge1_1__10), .d_arr_merge1_1__9 (
               d_arr_merge1_1__9), .d_arr_merge1_1__8 (d_arr_merge1_1__8), .d_arr_merge1_1__7 (
               d_arr_merge1_1__7), .d_arr_merge1_1__6 (d_arr_merge1_1__6), .d_arr_merge1_1__5 (
               d_arr_merge1_1__5), .d_arr_merge1_1__4 (d_arr_merge1_1__4), .d_arr_merge1_1__3 (
               d_arr_merge1_1__3), .d_arr_merge1_1__2 (d_arr_merge1_1__2), .d_arr_merge1_1__1 (
               d_arr_merge1_1__1), .d_arr_merge1_1__0 (d_arr_merge1_1__0), .d_arr_merge1_2__31 (
               GND0), .d_arr_merge1_2__30 (GND0), .d_arr_merge1_2__29 (GND0), .d_arr_merge1_2__28 (
               GND0), .d_arr_merge1_2__27 (GND0), .d_arr_merge1_2__26 (GND0), .d_arr_merge1_2__25 (
               GND0), .d_arr_merge1_2__24 (GND0), .d_arr_merge1_2__23 (GND0), .d_arr_merge1_2__22 (
               GND0), .d_arr_merge1_2__21 (GND0), .d_arr_merge1_2__20 (GND0), .d_arr_merge1_2__19 (
               GND0), .d_arr_merge1_2__18 (GND0), .d_arr_merge1_2__17 (GND0), .d_arr_merge1_2__16 (
               GND0), .d_arr_merge1_2__15 (GND0), .d_arr_merge1_2__14 (GND0), .d_arr_merge1_2__13 (
               GND0), .d_arr_merge1_2__12 (GND0), .d_arr_merge1_2__11 (GND0), .d_arr_merge1_2__10 (
               GND0), .d_arr_merge1_2__9 (GND0), .d_arr_merge1_2__8 (GND0), .d_arr_merge1_2__7 (
               GND0), .d_arr_merge1_2__6 (GND0), .d_arr_merge1_2__5 (GND0), .d_arr_merge1_2__4 (
               GND0), .d_arr_merge1_2__3 (GND0), .d_arr_merge1_2__2 (GND0), .d_arr_merge1_2__1 (
               GND0), .d_arr_merge1_2__0 (GND0), .d_arr_merge1_3__31 (GND0), .d_arr_merge1_3__30 (
               GND0), .d_arr_merge1_3__29 (GND0), .d_arr_merge1_3__28 (GND0), .d_arr_merge1_3__27 (
               GND0), .d_arr_merge1_3__26 (GND0), .d_arr_merge1_3__25 (GND0), .d_arr_merge1_3__24 (
               GND0), .d_arr_merge1_3__23 (GND0), .d_arr_merge1_3__22 (GND0), .d_arr_merge1_3__21 (
               GND0), .d_arr_merge1_3__20 (GND0), .d_arr_merge1_3__19 (GND0), .d_arr_merge1_3__18 (
               GND0), .d_arr_merge1_3__17 (GND0), .d_arr_merge1_3__16 (GND0), .d_arr_merge1_3__15 (
               GND0), .d_arr_merge1_3__14 (GND0), .d_arr_merge1_3__13 (GND0), .d_arr_merge1_3__12 (
               GND0), .d_arr_merge1_3__11 (GND0), .d_arr_merge1_3__10 (GND0), .d_arr_merge1_3__9 (
               GND0), .d_arr_merge1_3__8 (GND0), .d_arr_merge1_3__7 (GND0), .d_arr_merge1_3__6 (
               GND0), .d_arr_merge1_3__5 (GND0), .d_arr_merge1_3__4 (GND0), .d_arr_merge1_3__3 (
               GND0), .d_arr_merge1_3__2 (GND0), .d_arr_merge1_3__1 (GND0), .d_arr_merge1_3__0 (
               GND0), .d_arr_merge1_4__31 (GND0), .d_arr_merge1_4__30 (GND0), .d_arr_merge1_4__29 (
               GND0), .d_arr_merge1_4__28 (GND0), .d_arr_merge1_4__27 (GND0), .d_arr_merge1_4__26 (
               GND0), .d_arr_merge1_4__25 (GND0), .d_arr_merge1_4__24 (GND0), .d_arr_merge1_4__23 (
               GND0), .d_arr_merge1_4__22 (GND0), .d_arr_merge1_4__21 (GND0), .d_arr_merge1_4__20 (
               GND0), .d_arr_merge1_4__19 (GND0), .d_arr_merge1_4__18 (GND0), .d_arr_merge1_4__17 (
               GND0), .d_arr_merge1_4__16 (GND0), .d_arr_merge1_4__15 (GND0), .d_arr_merge1_4__14 (
               GND0), .d_arr_merge1_4__13 (GND0), .d_arr_merge1_4__12 (GND0), .d_arr_merge1_4__11 (
               GND0), .d_arr_merge1_4__10 (GND0), .d_arr_merge1_4__9 (GND0), .d_arr_merge1_4__8 (
               GND0), .d_arr_merge1_4__7 (GND0), .d_arr_merge1_4__6 (GND0), .d_arr_merge1_4__5 (
               GND0), .d_arr_merge1_4__4 (GND0), .d_arr_merge1_4__3 (GND0), .d_arr_merge1_4__2 (
               GND0), .d_arr_merge1_4__1 (GND0), .d_arr_merge1_4__0 (GND0), .d_arr_merge1_5__31 (
               GND0), .d_arr_merge1_5__30 (GND0), .d_arr_merge1_5__29 (GND0), .d_arr_merge1_5__28 (
               GND0), .d_arr_merge1_5__27 (GND0), .d_arr_merge1_5__26 (GND0), .d_arr_merge1_5__25 (
               GND0), .d_arr_merge1_5__24 (GND0), .d_arr_merge1_5__23 (GND0), .d_arr_merge1_5__22 (
               GND0), .d_arr_merge1_5__21 (GND0), .d_arr_merge1_5__20 (GND0), .d_arr_merge1_5__19 (
               GND0), .d_arr_merge1_5__18 (GND0), .d_arr_merge1_5__17 (GND0), .d_arr_merge1_5__16 (
               GND0), .d_arr_merge1_5__15 (GND0), .d_arr_merge1_5__14 (GND0), .d_arr_merge1_5__13 (
               GND0), .d_arr_merge1_5__12 (GND0), .d_arr_merge1_5__11 (GND0), .d_arr_merge1_5__10 (
               GND0), .d_arr_merge1_5__9 (GND0), .d_arr_merge1_5__8 (GND0), .d_arr_merge1_5__7 (
               GND0), .d_arr_merge1_5__6 (GND0), .d_arr_merge1_5__5 (GND0), .d_arr_merge1_5__4 (
               GND0), .d_arr_merge1_5__3 (GND0), .d_arr_merge1_5__2 (GND0), .d_arr_merge1_5__1 (
               GND0), .d_arr_merge1_5__0 (GND0), .d_arr_merge1_6__31 (GND0), .d_arr_merge1_6__30 (
               GND0), .d_arr_merge1_6__29 (GND0), .d_arr_merge1_6__28 (GND0), .d_arr_merge1_6__27 (
               GND0), .d_arr_merge1_6__26 (GND0), .d_arr_merge1_6__25 (GND0), .d_arr_merge1_6__24 (
               GND0), .d_arr_merge1_6__23 (GND0), .d_arr_merge1_6__22 (GND0), .d_arr_merge1_6__21 (
               GND0), .d_arr_merge1_6__20 (GND0), .d_arr_merge1_6__19 (GND0), .d_arr_merge1_6__18 (
               GND0), .d_arr_merge1_6__17 (GND0), .d_arr_merge1_6__16 (GND0), .d_arr_merge1_6__15 (
               GND0), .d_arr_merge1_6__14 (GND0), .d_arr_merge1_6__13 (GND0), .d_arr_merge1_6__12 (
               GND0), .d_arr_merge1_6__11 (GND0), .d_arr_merge1_6__10 (GND0), .d_arr_merge1_6__9 (
               GND0), .d_arr_merge1_6__8 (GND0), .d_arr_merge1_6__7 (GND0), .d_arr_merge1_6__6 (
               GND0), .d_arr_merge1_6__5 (GND0), .d_arr_merge1_6__4 (GND0), .d_arr_merge1_6__3 (
               GND0), .d_arr_merge1_6__2 (GND0), .d_arr_merge1_6__1 (GND0), .d_arr_merge1_6__0 (
               GND0), .d_arr_merge1_7__31 (GND0), .d_arr_merge1_7__30 (GND0), .d_arr_merge1_7__29 (
               GND0), .d_arr_merge1_7__28 (GND0), .d_arr_merge1_7__27 (GND0), .d_arr_merge1_7__26 (
               GND0), .d_arr_merge1_7__25 (GND0), .d_arr_merge1_7__24 (GND0), .d_arr_merge1_7__23 (
               GND0), .d_arr_merge1_7__22 (GND0), .d_arr_merge1_7__21 (GND0), .d_arr_merge1_7__20 (
               GND0), .d_arr_merge1_7__19 (GND0), .d_arr_merge1_7__18 (GND0), .d_arr_merge1_7__17 (
               GND0), .d_arr_merge1_7__16 (GND0), .d_arr_merge1_7__15 (GND0), .d_arr_merge1_7__14 (
               GND0), .d_arr_merge1_7__13 (GND0), .d_arr_merge1_7__12 (GND0), .d_arr_merge1_7__11 (
               GND0), .d_arr_merge1_7__10 (GND0), .d_arr_merge1_7__9 (GND0), .d_arr_merge1_7__8 (
               GND0), .d_arr_merge1_7__7 (GND0), .d_arr_merge1_7__6 (GND0), .d_arr_merge1_7__5 (
               GND0), .d_arr_merge1_7__4 (GND0), .d_arr_merge1_7__3 (GND0), .d_arr_merge1_7__2 (
               GND0), .d_arr_merge1_7__1 (GND0), .d_arr_merge1_7__0 (GND0), .d_arr_merge1_8__31 (
               GND0), .d_arr_merge1_8__30 (GND0), .d_arr_merge1_8__29 (GND0), .d_arr_merge1_8__28 (
               GND0), .d_arr_merge1_8__27 (GND0), .d_arr_merge1_8__26 (GND0), .d_arr_merge1_8__25 (
               GND0), .d_arr_merge1_8__24 (GND0), .d_arr_merge1_8__23 (GND0), .d_arr_merge1_8__22 (
               GND0), .d_arr_merge1_8__21 (GND0), .d_arr_merge1_8__20 (GND0), .d_arr_merge1_8__19 (
               GND0), .d_arr_merge1_8__18 (GND0), .d_arr_merge1_8__17 (GND0), .d_arr_merge1_8__16 (
               GND0), .d_arr_merge1_8__15 (GND0), .d_arr_merge1_8__14 (GND0), .d_arr_merge1_8__13 (
               GND0), .d_arr_merge1_8__12 (GND0), .d_arr_merge1_8__11 (GND0), .d_arr_merge1_8__10 (
               GND0), .d_arr_merge1_8__9 (GND0), .d_arr_merge1_8__8 (GND0), .d_arr_merge1_8__7 (
               GND0), .d_arr_merge1_8__6 (GND0), .d_arr_merge1_8__5 (GND0), .d_arr_merge1_8__4 (
               GND0), .d_arr_merge1_8__3 (GND0), .d_arr_merge1_8__2 (GND0), .d_arr_merge1_8__1 (
               GND0), .d_arr_merge1_8__0 (GND0), .d_arr_merge1_9__31 (GND0), .d_arr_merge1_9__30 (
               GND0), .d_arr_merge1_9__29 (GND0), .d_arr_merge1_9__28 (GND0), .d_arr_merge1_9__27 (
               GND0), .d_arr_merge1_9__26 (GND0), .d_arr_merge1_9__25 (GND0), .d_arr_merge1_9__24 (
               GND0), .d_arr_merge1_9__23 (GND0), .d_arr_merge1_9__22 (GND0), .d_arr_merge1_9__21 (
               GND0), .d_arr_merge1_9__20 (GND0), .d_arr_merge1_9__19 (GND0), .d_arr_merge1_9__18 (
               GND0), .d_arr_merge1_9__17 (GND0), .d_arr_merge1_9__16 (GND0), .d_arr_merge1_9__15 (
               GND0), .d_arr_merge1_9__14 (GND0), .d_arr_merge1_9__13 (GND0), .d_arr_merge1_9__12 (
               GND0), .d_arr_merge1_9__11 (GND0), .d_arr_merge1_9__10 (GND0), .d_arr_merge1_9__9 (
               GND0), .d_arr_merge1_9__8 (GND0), .d_arr_merge1_9__7 (GND0), .d_arr_merge1_9__6 (
               GND0), .d_arr_merge1_9__5 (GND0), .d_arr_merge1_9__4 (GND0), .d_arr_merge1_9__3 (
               GND0), .d_arr_merge1_9__2 (GND0), .d_arr_merge1_9__1 (GND0), .d_arr_merge1_9__0 (
               GND0), .d_arr_merge1_10__31 (GND0), .d_arr_merge1_10__30 (GND0), 
               .d_arr_merge1_10__29 (GND0), .d_arr_merge1_10__28 (GND0), .d_arr_merge1_10__27 (
               GND0), .d_arr_merge1_10__26 (GND0), .d_arr_merge1_10__25 (GND0), 
               .d_arr_merge1_10__24 (GND0), .d_arr_merge1_10__23 (GND0), .d_arr_merge1_10__22 (
               GND0), .d_arr_merge1_10__21 (GND0), .d_arr_merge1_10__20 (GND0), 
               .d_arr_merge1_10__19 (GND0), .d_arr_merge1_10__18 (GND0), .d_arr_merge1_10__17 (
               GND0), .d_arr_merge1_10__16 (GND0), .d_arr_merge1_10__15 (GND0), 
               .d_arr_merge1_10__14 (GND0), .d_arr_merge1_10__13 (GND0), .d_arr_merge1_10__12 (
               GND0), .d_arr_merge1_10__11 (GND0), .d_arr_merge1_10__10 (GND0), 
               .d_arr_merge1_10__9 (GND0), .d_arr_merge1_10__8 (GND0), .d_arr_merge1_10__7 (
               GND0), .d_arr_merge1_10__6 (GND0), .d_arr_merge1_10__5 (GND0), .d_arr_merge1_10__4 (
               GND0), .d_arr_merge1_10__3 (GND0), .d_arr_merge1_10__2 (GND0), .d_arr_merge1_10__1 (
               GND0), .d_arr_merge1_10__0 (GND0), .d_arr_merge1_11__31 (GND0), .d_arr_merge1_11__30 (
               GND0), .d_arr_merge1_11__29 (GND0), .d_arr_merge1_11__28 (GND0), 
               .d_arr_merge1_11__27 (GND0), .d_arr_merge1_11__26 (GND0), .d_arr_merge1_11__25 (
               GND0), .d_arr_merge1_11__24 (GND0), .d_arr_merge1_11__23 (GND0), 
               .d_arr_merge1_11__22 (GND0), .d_arr_merge1_11__21 (GND0), .d_arr_merge1_11__20 (
               GND0), .d_arr_merge1_11__19 (GND0), .d_arr_merge1_11__18 (GND0), 
               .d_arr_merge1_11__17 (GND0), .d_arr_merge1_11__16 (GND0), .d_arr_merge1_11__15 (
               GND0), .d_arr_merge1_11__14 (GND0), .d_arr_merge1_11__13 (GND0), 
               .d_arr_merge1_11__12 (GND0), .d_arr_merge1_11__11 (GND0), .d_arr_merge1_11__10 (
               GND0), .d_arr_merge1_11__9 (GND0), .d_arr_merge1_11__8 (GND0), .d_arr_merge1_11__7 (
               GND0), .d_arr_merge1_11__6 (GND0), .d_arr_merge1_11__5 (GND0), .d_arr_merge1_11__4 (
               GND0), .d_arr_merge1_11__3 (GND0), .d_arr_merge1_11__2 (GND0), .d_arr_merge1_11__1 (
               GND0), .d_arr_merge1_11__0 (GND0), .d_arr_merge1_12__31 (GND0), .d_arr_merge1_12__30 (
               GND0), .d_arr_merge1_12__29 (GND0), .d_arr_merge1_12__28 (GND0), 
               .d_arr_merge1_12__27 (GND0), .d_arr_merge1_12__26 (GND0), .d_arr_merge1_12__25 (
               GND0), .d_arr_merge1_12__24 (GND0), .d_arr_merge1_12__23 (GND0), 
               .d_arr_merge1_12__22 (GND0), .d_arr_merge1_12__21 (GND0), .d_arr_merge1_12__20 (
               GND0), .d_arr_merge1_12__19 (GND0), .d_arr_merge1_12__18 (GND0), 
               .d_arr_merge1_12__17 (GND0), .d_arr_merge1_12__16 (GND0), .d_arr_merge1_12__15 (
               GND0), .d_arr_merge1_12__14 (GND0), .d_arr_merge1_12__13 (GND0), 
               .d_arr_merge1_12__12 (GND0), .d_arr_merge1_12__11 (GND0), .d_arr_merge1_12__10 (
               GND0), .d_arr_merge1_12__9 (GND0), .d_arr_merge1_12__8 (GND0), .d_arr_merge1_12__7 (
               GND0), .d_arr_merge1_12__6 (GND0), .d_arr_merge1_12__5 (GND0), .d_arr_merge1_12__4 (
               GND0), .d_arr_merge1_12__3 (GND0), .d_arr_merge1_12__2 (GND0), .d_arr_merge1_12__1 (
               GND0), .d_arr_merge1_12__0 (GND0), .d_arr_merge1_13__31 (GND0), .d_arr_merge1_13__30 (
               GND0), .d_arr_merge1_13__29 (GND0), .d_arr_merge1_13__28 (GND0), 
               .d_arr_merge1_13__27 (GND0), .d_arr_merge1_13__26 (GND0), .d_arr_merge1_13__25 (
               GND0), .d_arr_merge1_13__24 (GND0), .d_arr_merge1_13__23 (GND0), 
               .d_arr_merge1_13__22 (GND0), .d_arr_merge1_13__21 (GND0), .d_arr_merge1_13__20 (
               GND0), .d_arr_merge1_13__19 (GND0), .d_arr_merge1_13__18 (GND0), 
               .d_arr_merge1_13__17 (GND0), .d_arr_merge1_13__16 (GND0), .d_arr_merge1_13__15 (
               GND0), .d_arr_merge1_13__14 (GND0), .d_arr_merge1_13__13 (GND0), 
               .d_arr_merge1_13__12 (GND0), .d_arr_merge1_13__11 (GND0), .d_arr_merge1_13__10 (
               GND0), .d_arr_merge1_13__9 (GND0), .d_arr_merge1_13__8 (GND0), .d_arr_merge1_13__7 (
               GND0), .d_arr_merge1_13__6 (GND0), .d_arr_merge1_13__5 (GND0), .d_arr_merge1_13__4 (
               GND0), .d_arr_merge1_13__3 (GND0), .d_arr_merge1_13__2 (GND0), .d_arr_merge1_13__1 (
               GND0), .d_arr_merge1_13__0 (GND0), .d_arr_merge1_14__31 (GND0), .d_arr_merge1_14__30 (
               GND0), .d_arr_merge1_14__29 (GND0), .d_arr_merge1_14__28 (GND0), 
               .d_arr_merge1_14__27 (GND0), .d_arr_merge1_14__26 (GND0), .d_arr_merge1_14__25 (
               GND0), .d_arr_merge1_14__24 (GND0), .d_arr_merge1_14__23 (GND0), 
               .d_arr_merge1_14__22 (GND0), .d_arr_merge1_14__21 (GND0), .d_arr_merge1_14__20 (
               GND0), .d_arr_merge1_14__19 (GND0), .d_arr_merge1_14__18 (GND0), 
               .d_arr_merge1_14__17 (GND0), .d_arr_merge1_14__16 (GND0), .d_arr_merge1_14__15 (
               GND0), .d_arr_merge1_14__14 (GND0), .d_arr_merge1_14__13 (GND0), 
               .d_arr_merge1_14__12 (GND0), .d_arr_merge1_14__11 (GND0), .d_arr_merge1_14__10 (
               GND0), .d_arr_merge1_14__9 (GND0), .d_arr_merge1_14__8 (GND0), .d_arr_merge1_14__7 (
               GND0), .d_arr_merge1_14__6 (GND0), .d_arr_merge1_14__5 (GND0), .d_arr_merge1_14__4 (
               GND0), .d_arr_merge1_14__3 (GND0), .d_arr_merge1_14__2 (GND0), .d_arr_merge1_14__1 (
               GND0), .d_arr_merge1_14__0 (GND0), .d_arr_merge1_15__31 (GND0), .d_arr_merge1_15__30 (
               GND0), .d_arr_merge1_15__29 (GND0), .d_arr_merge1_15__28 (GND0), 
               .d_arr_merge1_15__27 (GND0), .d_arr_merge1_15__26 (GND0), .d_arr_merge1_15__25 (
               GND0), .d_arr_merge1_15__24 (GND0), .d_arr_merge1_15__23 (GND0), 
               .d_arr_merge1_15__22 (GND0), .d_arr_merge1_15__21 (GND0), .d_arr_merge1_15__20 (
               GND0), .d_arr_merge1_15__19 (GND0), .d_arr_merge1_15__18 (GND0), 
               .d_arr_merge1_15__17 (GND0), .d_arr_merge1_15__16 (GND0), .d_arr_merge1_15__15 (
               GND0), .d_arr_merge1_15__14 (GND0), .d_arr_merge1_15__13 (GND0), 
               .d_arr_merge1_15__12 (GND0), .d_arr_merge1_15__11 (GND0), .d_arr_merge1_15__10 (
               GND0), .d_arr_merge1_15__9 (GND0), .d_arr_merge1_15__8 (GND0), .d_arr_merge1_15__7 (
               GND0), .d_arr_merge1_15__6 (GND0), .d_arr_merge1_15__5 (GND0), .d_arr_merge1_15__4 (
               GND0), .d_arr_merge1_15__3 (GND0), .d_arr_merge1_15__2 (GND0), .d_arr_merge1_15__1 (
               GND0), .d_arr_merge1_15__0 (GND0), .d_arr_merge1_16__31 (GND0), .d_arr_merge1_16__30 (
               GND0), .d_arr_merge1_16__29 (GND0), .d_arr_merge1_16__28 (GND0), 
               .d_arr_merge1_16__27 (GND0), .d_arr_merge1_16__26 (GND0), .d_arr_merge1_16__25 (
               GND0), .d_arr_merge1_16__24 (GND0), .d_arr_merge1_16__23 (GND0), 
               .d_arr_merge1_16__22 (GND0), .d_arr_merge1_16__21 (GND0), .d_arr_merge1_16__20 (
               GND0), .d_arr_merge1_16__19 (GND0), .d_arr_merge1_16__18 (GND0), 
               .d_arr_merge1_16__17 (GND0), .d_arr_merge1_16__16 (GND0), .d_arr_merge1_16__15 (
               GND0), .d_arr_merge1_16__14 (GND0), .d_arr_merge1_16__13 (GND0), 
               .d_arr_merge1_16__12 (GND0), .d_arr_merge1_16__11 (GND0), .d_arr_merge1_16__10 (
               GND0), .d_arr_merge1_16__9 (GND0), .d_arr_merge1_16__8 (GND0), .d_arr_merge1_16__7 (
               GND0), .d_arr_merge1_16__6 (GND0), .d_arr_merge1_16__5 (GND0), .d_arr_merge1_16__4 (
               GND0), .d_arr_merge1_16__3 (GND0), .d_arr_merge1_16__2 (GND0), .d_arr_merge1_16__1 (
               GND0), .d_arr_merge1_16__0 (GND0), .d_arr_merge1_17__31 (GND0), .d_arr_merge1_17__30 (
               GND0), .d_arr_merge1_17__29 (GND0), .d_arr_merge1_17__28 (GND0), 
               .d_arr_merge1_17__27 (GND0), .d_arr_merge1_17__26 (GND0), .d_arr_merge1_17__25 (
               GND0), .d_arr_merge1_17__24 (GND0), .d_arr_merge1_17__23 (GND0), 
               .d_arr_merge1_17__22 (GND0), .d_arr_merge1_17__21 (GND0), .d_arr_merge1_17__20 (
               GND0), .d_arr_merge1_17__19 (GND0), .d_arr_merge1_17__18 (GND0), 
               .d_arr_merge1_17__17 (GND0), .d_arr_merge1_17__16 (GND0), .d_arr_merge1_17__15 (
               GND0), .d_arr_merge1_17__14 (GND0), .d_arr_merge1_17__13 (GND0), 
               .d_arr_merge1_17__12 (GND0), .d_arr_merge1_17__11 (GND0), .d_arr_merge1_17__10 (
               GND0), .d_arr_merge1_17__9 (GND0), .d_arr_merge1_17__8 (GND0), .d_arr_merge1_17__7 (
               GND0), .d_arr_merge1_17__6 (GND0), .d_arr_merge1_17__5 (GND0), .d_arr_merge1_17__4 (
               GND0), .d_arr_merge1_17__3 (GND0), .d_arr_merge1_17__2 (GND0), .d_arr_merge1_17__1 (
               GND0), .d_arr_merge1_17__0 (GND0), .d_arr_merge1_18__31 (GND0), .d_arr_merge1_18__30 (
               GND0), .d_arr_merge1_18__29 (GND0), .d_arr_merge1_18__28 (GND0), 
               .d_arr_merge1_18__27 (GND0), .d_arr_merge1_18__26 (GND0), .d_arr_merge1_18__25 (
               GND0), .d_arr_merge1_18__24 (GND0), .d_arr_merge1_18__23 (GND0), 
               .d_arr_merge1_18__22 (GND0), .d_arr_merge1_18__21 (GND0), .d_arr_merge1_18__20 (
               GND0), .d_arr_merge1_18__19 (GND0), .d_arr_merge1_18__18 (GND0), 
               .d_arr_merge1_18__17 (GND0), .d_arr_merge1_18__16 (GND0), .d_arr_merge1_18__15 (
               GND0), .d_arr_merge1_18__14 (GND0), .d_arr_merge1_18__13 (GND0), 
               .d_arr_merge1_18__12 (GND0), .d_arr_merge1_18__11 (GND0), .d_arr_merge1_18__10 (
               GND0), .d_arr_merge1_18__9 (GND0), .d_arr_merge1_18__8 (GND0), .d_arr_merge1_18__7 (
               GND0), .d_arr_merge1_18__6 (GND0), .d_arr_merge1_18__5 (GND0), .d_arr_merge1_18__4 (
               GND0), .d_arr_merge1_18__3 (GND0), .d_arr_merge1_18__2 (GND0), .d_arr_merge1_18__1 (
               GND0), .d_arr_merge1_18__0 (GND0), .d_arr_merge1_19__31 (GND0), .d_arr_merge1_19__30 (
               GND0), .d_arr_merge1_19__29 (GND0), .d_arr_merge1_19__28 (GND0), 
               .d_arr_merge1_19__27 (GND0), .d_arr_merge1_19__26 (GND0), .d_arr_merge1_19__25 (
               GND0), .d_arr_merge1_19__24 (GND0), .d_arr_merge1_19__23 (GND0), 
               .d_arr_merge1_19__22 (GND0), .d_arr_merge1_19__21 (GND0), .d_arr_merge1_19__20 (
               GND0), .d_arr_merge1_19__19 (GND0), .d_arr_merge1_19__18 (GND0), 
               .d_arr_merge1_19__17 (GND0), .d_arr_merge1_19__16 (GND0), .d_arr_merge1_19__15 (
               GND0), .d_arr_merge1_19__14 (GND0), .d_arr_merge1_19__13 (GND0), 
               .d_arr_merge1_19__12 (GND0), .d_arr_merge1_19__11 (GND0), .d_arr_merge1_19__10 (
               GND0), .d_arr_merge1_19__9 (GND0), .d_arr_merge1_19__8 (GND0), .d_arr_merge1_19__7 (
               GND0), .d_arr_merge1_19__6 (GND0), .d_arr_merge1_19__5 (GND0), .d_arr_merge1_19__4 (
               GND0), .d_arr_merge1_19__3 (GND0), .d_arr_merge1_19__2 (GND0), .d_arr_merge1_19__1 (
               GND0), .d_arr_merge1_19__0 (GND0), .d_arr_merge1_20__31 (GND0), .d_arr_merge1_20__30 (
               GND0), .d_arr_merge1_20__29 (GND0), .d_arr_merge1_20__28 (GND0), 
               .d_arr_merge1_20__27 (GND0), .d_arr_merge1_20__26 (GND0), .d_arr_merge1_20__25 (
               GND0), .d_arr_merge1_20__24 (GND0), .d_arr_merge1_20__23 (GND0), 
               .d_arr_merge1_20__22 (GND0), .d_arr_merge1_20__21 (GND0), .d_arr_merge1_20__20 (
               GND0), .d_arr_merge1_20__19 (GND0), .d_arr_merge1_20__18 (GND0), 
               .d_arr_merge1_20__17 (GND0), .d_arr_merge1_20__16 (GND0), .d_arr_merge1_20__15 (
               GND0), .d_arr_merge1_20__14 (GND0), .d_arr_merge1_20__13 (GND0), 
               .d_arr_merge1_20__12 (GND0), .d_arr_merge1_20__11 (GND0), .d_arr_merge1_20__10 (
               GND0), .d_arr_merge1_20__9 (GND0), .d_arr_merge1_20__8 (GND0), .d_arr_merge1_20__7 (
               GND0), .d_arr_merge1_20__6 (GND0), .d_arr_merge1_20__5 (GND0), .d_arr_merge1_20__4 (
               GND0), .d_arr_merge1_20__3 (GND0), .d_arr_merge1_20__2 (GND0), .d_arr_merge1_20__1 (
               GND0), .d_arr_merge1_20__0 (GND0), .d_arr_merge1_21__31 (GND0), .d_arr_merge1_21__30 (
               GND0), .d_arr_merge1_21__29 (GND0), .d_arr_merge1_21__28 (GND0), 
               .d_arr_merge1_21__27 (GND0), .d_arr_merge1_21__26 (GND0), .d_arr_merge1_21__25 (
               GND0), .d_arr_merge1_21__24 (GND0), .d_arr_merge1_21__23 (GND0), 
               .d_arr_merge1_21__22 (GND0), .d_arr_merge1_21__21 (GND0), .d_arr_merge1_21__20 (
               GND0), .d_arr_merge1_21__19 (GND0), .d_arr_merge1_21__18 (GND0), 
               .d_arr_merge1_21__17 (GND0), .d_arr_merge1_21__16 (GND0), .d_arr_merge1_21__15 (
               GND0), .d_arr_merge1_21__14 (GND0), .d_arr_merge1_21__13 (GND0), 
               .d_arr_merge1_21__12 (GND0), .d_arr_merge1_21__11 (GND0), .d_arr_merge1_21__10 (
               GND0), .d_arr_merge1_21__9 (GND0), .d_arr_merge1_21__8 (GND0), .d_arr_merge1_21__7 (
               GND0), .d_arr_merge1_21__6 (GND0), .d_arr_merge1_21__5 (GND0), .d_arr_merge1_21__4 (
               GND0), .d_arr_merge1_21__3 (GND0), .d_arr_merge1_21__2 (GND0), .d_arr_merge1_21__1 (
               GND0), .d_arr_merge1_21__0 (GND0), .d_arr_merge1_22__31 (GND0), .d_arr_merge1_22__30 (
               GND0), .d_arr_merge1_22__29 (GND0), .d_arr_merge1_22__28 (GND0), 
               .d_arr_merge1_22__27 (GND0), .d_arr_merge1_22__26 (GND0), .d_arr_merge1_22__25 (
               GND0), .d_arr_merge1_22__24 (GND0), .d_arr_merge1_22__23 (GND0), 
               .d_arr_merge1_22__22 (GND0), .d_arr_merge1_22__21 (GND0), .d_arr_merge1_22__20 (
               GND0), .d_arr_merge1_22__19 (GND0), .d_arr_merge1_22__18 (GND0), 
               .d_arr_merge1_22__17 (GND0), .d_arr_merge1_22__16 (GND0), .d_arr_merge1_22__15 (
               GND0), .d_arr_merge1_22__14 (GND0), .d_arr_merge1_22__13 (GND0), 
               .d_arr_merge1_22__12 (GND0), .d_arr_merge1_22__11 (GND0), .d_arr_merge1_22__10 (
               GND0), .d_arr_merge1_22__9 (GND0), .d_arr_merge1_22__8 (GND0), .d_arr_merge1_22__7 (
               GND0), .d_arr_merge1_22__6 (GND0), .d_arr_merge1_22__5 (GND0), .d_arr_merge1_22__4 (
               GND0), .d_arr_merge1_22__3 (GND0), .d_arr_merge1_22__2 (GND0), .d_arr_merge1_22__1 (
               GND0), .d_arr_merge1_22__0 (GND0), .d_arr_merge1_23__31 (GND0), .d_arr_merge1_23__30 (
               GND0), .d_arr_merge1_23__29 (GND0), .d_arr_merge1_23__28 (GND0), 
               .d_arr_merge1_23__27 (GND0), .d_arr_merge1_23__26 (GND0), .d_arr_merge1_23__25 (
               GND0), .d_arr_merge1_23__24 (GND0), .d_arr_merge1_23__23 (GND0), 
               .d_arr_merge1_23__22 (GND0), .d_arr_merge1_23__21 (GND0), .d_arr_merge1_23__20 (
               GND0), .d_arr_merge1_23__19 (GND0), .d_arr_merge1_23__18 (GND0), 
               .d_arr_merge1_23__17 (GND0), .d_arr_merge1_23__16 (GND0), .d_arr_merge1_23__15 (
               GND0), .d_arr_merge1_23__14 (GND0), .d_arr_merge1_23__13 (GND0), 
               .d_arr_merge1_23__12 (GND0), .d_arr_merge1_23__11 (GND0), .d_arr_merge1_23__10 (
               GND0), .d_arr_merge1_23__9 (GND0), .d_arr_merge1_23__8 (GND0), .d_arr_merge1_23__7 (
               GND0), .d_arr_merge1_23__6 (GND0), .d_arr_merge1_23__5 (GND0), .d_arr_merge1_23__4 (
               GND0), .d_arr_merge1_23__3 (GND0), .d_arr_merge1_23__2 (GND0), .d_arr_merge1_23__1 (
               GND0), .d_arr_merge1_23__0 (GND0), .d_arr_merge1_24__31 (GND0), .d_arr_merge1_24__30 (
               GND0), .d_arr_merge1_24__29 (GND0), .d_arr_merge1_24__28 (GND0), 
               .d_arr_merge1_24__27 (GND0), .d_arr_merge1_24__26 (GND0), .d_arr_merge1_24__25 (
               GND0), .d_arr_merge1_24__24 (GND0), .d_arr_merge1_24__23 (GND0), 
               .d_arr_merge1_24__22 (GND0), .d_arr_merge1_24__21 (GND0), .d_arr_merge1_24__20 (
               GND0), .d_arr_merge1_24__19 (GND0), .d_arr_merge1_24__18 (GND0), 
               .d_arr_merge1_24__17 (GND0), .d_arr_merge1_24__16 (GND0), .d_arr_merge1_24__15 (
               GND0), .d_arr_merge1_24__14 (GND0), .d_arr_merge1_24__13 (GND0), 
               .d_arr_merge1_24__12 (GND0), .d_arr_merge1_24__11 (GND0), .d_arr_merge1_24__10 (
               GND0), .d_arr_merge1_24__9 (GND0), .d_arr_merge1_24__8 (GND0), .d_arr_merge1_24__7 (
               GND0), .d_arr_merge1_24__6 (GND0), .d_arr_merge1_24__5 (GND0), .d_arr_merge1_24__4 (
               GND0), .d_arr_merge1_24__3 (GND0), .d_arr_merge1_24__2 (GND0), .d_arr_merge1_24__1 (
               GND0), .d_arr_merge1_24__0 (GND0), .d_arr_merge2_0__31 (
               d_arr_merge2_0__31), .d_arr_merge2_0__30 (d_arr_merge2_0__31), .d_arr_merge2_0__29 (
               d_arr_merge2_0__31), .d_arr_merge2_0__28 (d_arr_merge2_0__31), .d_arr_merge2_0__27 (
               d_arr_merge2_0__31), .d_arr_merge2_0__26 (d_arr_merge2_0__26), .d_arr_merge2_0__25 (
               d_arr_merge2_0__25), .d_arr_merge2_0__24 (d_arr_merge2_0__24), .d_arr_merge2_0__23 (
               d_arr_merge2_0__23), .d_arr_merge2_0__22 (d_arr_merge2_0__22), .d_arr_merge2_0__21 (
               d_arr_merge2_0__21), .d_arr_merge2_0__20 (d_arr_merge2_0__20), .d_arr_merge2_0__19 (
               d_arr_merge2_0__19), .d_arr_merge2_0__18 (d_arr_merge2_0__18), .d_arr_merge2_0__17 (
               d_arr_merge2_0__17), .d_arr_merge2_0__16 (d_arr_merge2_0__16), .d_arr_merge2_0__15 (
               d_arr_merge2_0__15), .d_arr_merge2_0__14 (d_arr_merge2_0__14), .d_arr_merge2_0__13 (
               d_arr_merge2_0__13), .d_arr_merge2_0__12 (d_arr_merge2_0__12), .d_arr_merge2_0__11 (
               d_arr_merge2_0__11), .d_arr_merge2_0__10 (d_arr_merge2_0__10), .d_arr_merge2_0__9 (
               d_arr_merge2_0__9), .d_arr_merge2_0__8 (d_arr_merge2_0__8), .d_arr_merge2_0__7 (
               d_arr_merge2_0__7), .d_arr_merge2_0__6 (d_arr_merge2_0__6), .d_arr_merge2_0__5 (
               d_arr_merge2_0__5), .d_arr_merge2_0__4 (d_arr_merge2_0__4), .d_arr_merge2_0__3 (
               d_arr_merge2_0__3), .d_arr_merge2_0__2 (d_arr_merge2_0__2), .d_arr_merge2_0__1 (
               d_arr_merge2_0__1), .d_arr_merge2_0__0 (d_arr_merge2_0__0), .d_arr_merge2_1__31 (
               d_arr_merge2_1__31), .d_arr_merge2_1__30 (d_arr_merge2_1__31), .d_arr_merge2_1__29 (
               d_arr_merge2_1__31), .d_arr_merge2_1__28 (d_arr_merge2_1__31), .d_arr_merge2_1__27 (
               d_arr_merge2_1__31), .d_arr_merge2_1__26 (d_arr_merge2_1__26), .d_arr_merge2_1__25 (
               d_arr_merge2_1__25), .d_arr_merge2_1__24 (d_arr_merge2_1__24), .d_arr_merge2_1__23 (
               d_arr_merge2_1__23), .d_arr_merge2_1__22 (d_arr_merge2_1__22), .d_arr_merge2_1__21 (
               d_arr_merge2_1__21), .d_arr_merge2_1__20 (d_arr_merge2_1__20), .d_arr_merge2_1__19 (
               d_arr_merge2_1__19), .d_arr_merge2_1__18 (d_arr_merge2_1__18), .d_arr_merge2_1__17 (
               d_arr_merge2_1__17), .d_arr_merge2_1__16 (d_arr_merge2_1__16), .d_arr_merge2_1__15 (
               d_arr_merge2_1__15), .d_arr_merge2_1__14 (d_arr_merge2_1__14), .d_arr_merge2_1__13 (
               d_arr_merge2_1__13), .d_arr_merge2_1__12 (d_arr_merge2_1__12), .d_arr_merge2_1__11 (
               d_arr_merge2_1__11), .d_arr_merge2_1__10 (d_arr_merge2_1__10), .d_arr_merge2_1__9 (
               d_arr_merge2_1__9), .d_arr_merge2_1__8 (d_arr_merge2_1__8), .d_arr_merge2_1__7 (
               d_arr_merge2_1__7), .d_arr_merge2_1__6 (d_arr_merge2_1__6), .d_arr_merge2_1__5 (
               d_arr_merge2_1__5), .d_arr_merge2_1__4 (d_arr_merge2_1__4), .d_arr_merge2_1__3 (
               d_arr_merge2_1__3), .d_arr_merge2_1__2 (d_arr_merge2_1__2), .d_arr_merge2_1__1 (
               d_arr_merge2_1__1), .d_arr_merge2_1__0 (d_arr_merge2_1__0), .d_arr_merge2_2__31 (
               GND0), .d_arr_merge2_2__30 (GND0), .d_arr_merge2_2__29 (GND0), .d_arr_merge2_2__28 (
               GND0), .d_arr_merge2_2__27 (GND0), .d_arr_merge2_2__26 (GND0), .d_arr_merge2_2__25 (
               GND0), .d_arr_merge2_2__24 (GND0), .d_arr_merge2_2__23 (GND0), .d_arr_merge2_2__22 (
               GND0), .d_arr_merge2_2__21 (GND0), .d_arr_merge2_2__20 (GND0), .d_arr_merge2_2__19 (
               GND0), .d_arr_merge2_2__18 (GND0), .d_arr_merge2_2__17 (GND0), .d_arr_merge2_2__16 (
               GND0), .d_arr_merge2_2__15 (GND0), .d_arr_merge2_2__14 (GND0), .d_arr_merge2_2__13 (
               GND0), .d_arr_merge2_2__12 (GND0), .d_arr_merge2_2__11 (GND0), .d_arr_merge2_2__10 (
               GND0), .d_arr_merge2_2__9 (GND0), .d_arr_merge2_2__8 (GND0), .d_arr_merge2_2__7 (
               GND0), .d_arr_merge2_2__6 (GND0), .d_arr_merge2_2__5 (GND0), .d_arr_merge2_2__4 (
               GND0), .d_arr_merge2_2__3 (GND0), .d_arr_merge2_2__2 (GND0), .d_arr_merge2_2__1 (
               GND0), .d_arr_merge2_2__0 (GND0), .d_arr_merge2_3__31 (GND0), .d_arr_merge2_3__30 (
               GND0), .d_arr_merge2_3__29 (GND0), .d_arr_merge2_3__28 (GND0), .d_arr_merge2_3__27 (
               GND0), .d_arr_merge2_3__26 (GND0), .d_arr_merge2_3__25 (GND0), .d_arr_merge2_3__24 (
               GND0), .d_arr_merge2_3__23 (GND0), .d_arr_merge2_3__22 (GND0), .d_arr_merge2_3__21 (
               GND0), .d_arr_merge2_3__20 (GND0), .d_arr_merge2_3__19 (GND0), .d_arr_merge2_3__18 (
               GND0), .d_arr_merge2_3__17 (GND0), .d_arr_merge2_3__16 (GND0), .d_arr_merge2_3__15 (
               GND0), .d_arr_merge2_3__14 (GND0), .d_arr_merge2_3__13 (GND0), .d_arr_merge2_3__12 (
               GND0), .d_arr_merge2_3__11 (GND0), .d_arr_merge2_3__10 (GND0), .d_arr_merge2_3__9 (
               GND0), .d_arr_merge2_3__8 (GND0), .d_arr_merge2_3__7 (GND0), .d_arr_merge2_3__6 (
               GND0), .d_arr_merge2_3__5 (GND0), .d_arr_merge2_3__4 (GND0), .d_arr_merge2_3__3 (
               GND0), .d_arr_merge2_3__2 (GND0), .d_arr_merge2_3__1 (GND0), .d_arr_merge2_3__0 (
               GND0), .d_arr_merge2_4__31 (GND0), .d_arr_merge2_4__30 (GND0), .d_arr_merge2_4__29 (
               GND0), .d_arr_merge2_4__28 (GND0), .d_arr_merge2_4__27 (GND0), .d_arr_merge2_4__26 (
               GND0), .d_arr_merge2_4__25 (GND0), .d_arr_merge2_4__24 (GND0), .d_arr_merge2_4__23 (
               GND0), .d_arr_merge2_4__22 (GND0), .d_arr_merge2_4__21 (GND0), .d_arr_merge2_4__20 (
               GND0), .d_arr_merge2_4__19 (GND0), .d_arr_merge2_4__18 (GND0), .d_arr_merge2_4__17 (
               GND0), .d_arr_merge2_4__16 (GND0), .d_arr_merge2_4__15 (GND0), .d_arr_merge2_4__14 (
               GND0), .d_arr_merge2_4__13 (GND0), .d_arr_merge2_4__12 (GND0), .d_arr_merge2_4__11 (
               GND0), .d_arr_merge2_4__10 (GND0), .d_arr_merge2_4__9 (GND0), .d_arr_merge2_4__8 (
               GND0), .d_arr_merge2_4__7 (GND0), .d_arr_merge2_4__6 (GND0), .d_arr_merge2_4__5 (
               GND0), .d_arr_merge2_4__4 (GND0), .d_arr_merge2_4__3 (GND0), .d_arr_merge2_4__2 (
               GND0), .d_arr_merge2_4__1 (GND0), .d_arr_merge2_4__0 (GND0), .d_arr_merge2_5__31 (
               GND0), .d_arr_merge2_5__30 (GND0), .d_arr_merge2_5__29 (GND0), .d_arr_merge2_5__28 (
               GND0), .d_arr_merge2_5__27 (GND0), .d_arr_merge2_5__26 (GND0), .d_arr_merge2_5__25 (
               GND0), .d_arr_merge2_5__24 (GND0), .d_arr_merge2_5__23 (GND0), .d_arr_merge2_5__22 (
               GND0), .d_arr_merge2_5__21 (GND0), .d_arr_merge2_5__20 (GND0), .d_arr_merge2_5__19 (
               GND0), .d_arr_merge2_5__18 (GND0), .d_arr_merge2_5__17 (GND0), .d_arr_merge2_5__16 (
               GND0), .d_arr_merge2_5__15 (GND0), .d_arr_merge2_5__14 (GND0), .d_arr_merge2_5__13 (
               GND0), .d_arr_merge2_5__12 (GND0), .d_arr_merge2_5__11 (GND0), .d_arr_merge2_5__10 (
               GND0), .d_arr_merge2_5__9 (GND0), .d_arr_merge2_5__8 (GND0), .d_arr_merge2_5__7 (
               GND0), .d_arr_merge2_5__6 (GND0), .d_arr_merge2_5__5 (GND0), .d_arr_merge2_5__4 (
               GND0), .d_arr_merge2_5__3 (GND0), .d_arr_merge2_5__2 (GND0), .d_arr_merge2_5__1 (
               GND0), .d_arr_merge2_5__0 (GND0), .d_arr_merge2_6__31 (GND0), .d_arr_merge2_6__30 (
               GND0), .d_arr_merge2_6__29 (GND0), .d_arr_merge2_6__28 (GND0), .d_arr_merge2_6__27 (
               GND0), .d_arr_merge2_6__26 (GND0), .d_arr_merge2_6__25 (GND0), .d_arr_merge2_6__24 (
               GND0), .d_arr_merge2_6__23 (GND0), .d_arr_merge2_6__22 (GND0), .d_arr_merge2_6__21 (
               GND0), .d_arr_merge2_6__20 (GND0), .d_arr_merge2_6__19 (GND0), .d_arr_merge2_6__18 (
               GND0), .d_arr_merge2_6__17 (GND0), .d_arr_merge2_6__16 (GND0), .d_arr_merge2_6__15 (
               GND0), .d_arr_merge2_6__14 (GND0), .d_arr_merge2_6__13 (GND0), .d_arr_merge2_6__12 (
               GND0), .d_arr_merge2_6__11 (GND0), .d_arr_merge2_6__10 (GND0), .d_arr_merge2_6__9 (
               GND0), .d_arr_merge2_6__8 (GND0), .d_arr_merge2_6__7 (GND0), .d_arr_merge2_6__6 (
               GND0), .d_arr_merge2_6__5 (GND0), .d_arr_merge2_6__4 (GND0), .d_arr_merge2_6__3 (
               GND0), .d_arr_merge2_6__2 (GND0), .d_arr_merge2_6__1 (GND0), .d_arr_merge2_6__0 (
               GND0), .d_arr_merge2_7__31 (GND0), .d_arr_merge2_7__30 (GND0), .d_arr_merge2_7__29 (
               GND0), .d_arr_merge2_7__28 (GND0), .d_arr_merge2_7__27 (GND0), .d_arr_merge2_7__26 (
               GND0), .d_arr_merge2_7__25 (GND0), .d_arr_merge2_7__24 (GND0), .d_arr_merge2_7__23 (
               GND0), .d_arr_merge2_7__22 (GND0), .d_arr_merge2_7__21 (GND0), .d_arr_merge2_7__20 (
               GND0), .d_arr_merge2_7__19 (GND0), .d_arr_merge2_7__18 (GND0), .d_arr_merge2_7__17 (
               GND0), .d_arr_merge2_7__16 (GND0), .d_arr_merge2_7__15 (GND0), .d_arr_merge2_7__14 (
               GND0), .d_arr_merge2_7__13 (GND0), .d_arr_merge2_7__12 (GND0), .d_arr_merge2_7__11 (
               GND0), .d_arr_merge2_7__10 (GND0), .d_arr_merge2_7__9 (GND0), .d_arr_merge2_7__8 (
               GND0), .d_arr_merge2_7__7 (GND0), .d_arr_merge2_7__6 (GND0), .d_arr_merge2_7__5 (
               GND0), .d_arr_merge2_7__4 (GND0), .d_arr_merge2_7__3 (GND0), .d_arr_merge2_7__2 (
               GND0), .d_arr_merge2_7__1 (GND0), .d_arr_merge2_7__0 (GND0), .d_arr_merge2_8__31 (
               GND0), .d_arr_merge2_8__30 (GND0), .d_arr_merge2_8__29 (GND0), .d_arr_merge2_8__28 (
               GND0), .d_arr_merge2_8__27 (GND0), .d_arr_merge2_8__26 (GND0), .d_arr_merge2_8__25 (
               GND0), .d_arr_merge2_8__24 (GND0), .d_arr_merge2_8__23 (GND0), .d_arr_merge2_8__22 (
               GND0), .d_arr_merge2_8__21 (GND0), .d_arr_merge2_8__20 (GND0), .d_arr_merge2_8__19 (
               GND0), .d_arr_merge2_8__18 (GND0), .d_arr_merge2_8__17 (GND0), .d_arr_merge2_8__16 (
               GND0), .d_arr_merge2_8__15 (GND0), .d_arr_merge2_8__14 (GND0), .d_arr_merge2_8__13 (
               GND0), .d_arr_merge2_8__12 (GND0), .d_arr_merge2_8__11 (GND0), .d_arr_merge2_8__10 (
               GND0), .d_arr_merge2_8__9 (GND0), .d_arr_merge2_8__8 (GND0), .d_arr_merge2_8__7 (
               GND0), .d_arr_merge2_8__6 (GND0), .d_arr_merge2_8__5 (GND0), .d_arr_merge2_8__4 (
               GND0), .d_arr_merge2_8__3 (GND0), .d_arr_merge2_8__2 (GND0), .d_arr_merge2_8__1 (
               GND0), .d_arr_merge2_8__0 (GND0), .d_arr_merge2_9__31 (GND0), .d_arr_merge2_9__30 (
               GND0), .d_arr_merge2_9__29 (GND0), .d_arr_merge2_9__28 (GND0), .d_arr_merge2_9__27 (
               GND0), .d_arr_merge2_9__26 (GND0), .d_arr_merge2_9__25 (GND0), .d_arr_merge2_9__24 (
               GND0), .d_arr_merge2_9__23 (GND0), .d_arr_merge2_9__22 (GND0), .d_arr_merge2_9__21 (
               GND0), .d_arr_merge2_9__20 (GND0), .d_arr_merge2_9__19 (GND0), .d_arr_merge2_9__18 (
               GND0), .d_arr_merge2_9__17 (GND0), .d_arr_merge2_9__16 (GND0), .d_arr_merge2_9__15 (
               GND0), .d_arr_merge2_9__14 (GND0), .d_arr_merge2_9__13 (GND0), .d_arr_merge2_9__12 (
               GND0), .d_arr_merge2_9__11 (GND0), .d_arr_merge2_9__10 (GND0), .d_arr_merge2_9__9 (
               GND0), .d_arr_merge2_9__8 (GND0), .d_arr_merge2_9__7 (GND0), .d_arr_merge2_9__6 (
               GND0), .d_arr_merge2_9__5 (GND0), .d_arr_merge2_9__4 (GND0), .d_arr_merge2_9__3 (
               GND0), .d_arr_merge2_9__2 (GND0), .d_arr_merge2_9__1 (GND0), .d_arr_merge2_9__0 (
               GND0), .d_arr_merge2_10__31 (GND0), .d_arr_merge2_10__30 (GND0), 
               .d_arr_merge2_10__29 (GND0), .d_arr_merge2_10__28 (GND0), .d_arr_merge2_10__27 (
               GND0), .d_arr_merge2_10__26 (GND0), .d_arr_merge2_10__25 (GND0), 
               .d_arr_merge2_10__24 (GND0), .d_arr_merge2_10__23 (GND0), .d_arr_merge2_10__22 (
               GND0), .d_arr_merge2_10__21 (GND0), .d_arr_merge2_10__20 (GND0), 
               .d_arr_merge2_10__19 (GND0), .d_arr_merge2_10__18 (GND0), .d_arr_merge2_10__17 (
               GND0), .d_arr_merge2_10__16 (GND0), .d_arr_merge2_10__15 (GND0), 
               .d_arr_merge2_10__14 (GND0), .d_arr_merge2_10__13 (GND0), .d_arr_merge2_10__12 (
               GND0), .d_arr_merge2_10__11 (GND0), .d_arr_merge2_10__10 (GND0), 
               .d_arr_merge2_10__9 (GND0), .d_arr_merge2_10__8 (GND0), .d_arr_merge2_10__7 (
               GND0), .d_arr_merge2_10__6 (GND0), .d_arr_merge2_10__5 (GND0), .d_arr_merge2_10__4 (
               GND0), .d_arr_merge2_10__3 (GND0), .d_arr_merge2_10__2 (GND0), .d_arr_merge2_10__1 (
               GND0), .d_arr_merge2_10__0 (GND0), .d_arr_merge2_11__31 (GND0), .d_arr_merge2_11__30 (
               GND0), .d_arr_merge2_11__29 (GND0), .d_arr_merge2_11__28 (GND0), 
               .d_arr_merge2_11__27 (GND0), .d_arr_merge2_11__26 (GND0), .d_arr_merge2_11__25 (
               GND0), .d_arr_merge2_11__24 (GND0), .d_arr_merge2_11__23 (GND0), 
               .d_arr_merge2_11__22 (GND0), .d_arr_merge2_11__21 (GND0), .d_arr_merge2_11__20 (
               GND0), .d_arr_merge2_11__19 (GND0), .d_arr_merge2_11__18 (GND0), 
               .d_arr_merge2_11__17 (GND0), .d_arr_merge2_11__16 (GND0), .d_arr_merge2_11__15 (
               GND0), .d_arr_merge2_11__14 (GND0), .d_arr_merge2_11__13 (GND0), 
               .d_arr_merge2_11__12 (GND0), .d_arr_merge2_11__11 (GND0), .d_arr_merge2_11__10 (
               GND0), .d_arr_merge2_11__9 (GND0), .d_arr_merge2_11__8 (GND0), .d_arr_merge2_11__7 (
               GND0), .d_arr_merge2_11__6 (GND0), .d_arr_merge2_11__5 (GND0), .d_arr_merge2_11__4 (
               GND0), .d_arr_merge2_11__3 (GND0), .d_arr_merge2_11__2 (GND0), .d_arr_merge2_11__1 (
               GND0), .d_arr_merge2_11__0 (GND0), .d_arr_merge2_12__31 (GND0), .d_arr_merge2_12__30 (
               GND0), .d_arr_merge2_12__29 (GND0), .d_arr_merge2_12__28 (GND0), 
               .d_arr_merge2_12__27 (GND0), .d_arr_merge2_12__26 (GND0), .d_arr_merge2_12__25 (
               GND0), .d_arr_merge2_12__24 (GND0), .d_arr_merge2_12__23 (GND0), 
               .d_arr_merge2_12__22 (GND0), .d_arr_merge2_12__21 (GND0), .d_arr_merge2_12__20 (
               GND0), .d_arr_merge2_12__19 (GND0), .d_arr_merge2_12__18 (GND0), 
               .d_arr_merge2_12__17 (GND0), .d_arr_merge2_12__16 (GND0), .d_arr_merge2_12__15 (
               GND0), .d_arr_merge2_12__14 (GND0), .d_arr_merge2_12__13 (GND0), 
               .d_arr_merge2_12__12 (GND0), .d_arr_merge2_12__11 (GND0), .d_arr_merge2_12__10 (
               GND0), .d_arr_merge2_12__9 (GND0), .d_arr_merge2_12__8 (GND0), .d_arr_merge2_12__7 (
               GND0), .d_arr_merge2_12__6 (GND0), .d_arr_merge2_12__5 (GND0), .d_arr_merge2_12__4 (
               GND0), .d_arr_merge2_12__3 (GND0), .d_arr_merge2_12__2 (GND0), .d_arr_merge2_12__1 (
               GND0), .d_arr_merge2_12__0 (GND0), .d_arr_merge2_13__31 (GND0), .d_arr_merge2_13__30 (
               GND0), .d_arr_merge2_13__29 (GND0), .d_arr_merge2_13__28 (GND0), 
               .d_arr_merge2_13__27 (GND0), .d_arr_merge2_13__26 (GND0), .d_arr_merge2_13__25 (
               GND0), .d_arr_merge2_13__24 (GND0), .d_arr_merge2_13__23 (GND0), 
               .d_arr_merge2_13__22 (GND0), .d_arr_merge2_13__21 (GND0), .d_arr_merge2_13__20 (
               GND0), .d_arr_merge2_13__19 (GND0), .d_arr_merge2_13__18 (GND0), 
               .d_arr_merge2_13__17 (GND0), .d_arr_merge2_13__16 (GND0), .d_arr_merge2_13__15 (
               GND0), .d_arr_merge2_13__14 (GND0), .d_arr_merge2_13__13 (GND0), 
               .d_arr_merge2_13__12 (GND0), .d_arr_merge2_13__11 (GND0), .d_arr_merge2_13__10 (
               GND0), .d_arr_merge2_13__9 (GND0), .d_arr_merge2_13__8 (GND0), .d_arr_merge2_13__7 (
               GND0), .d_arr_merge2_13__6 (GND0), .d_arr_merge2_13__5 (GND0), .d_arr_merge2_13__4 (
               GND0), .d_arr_merge2_13__3 (GND0), .d_arr_merge2_13__2 (GND0), .d_arr_merge2_13__1 (
               GND0), .d_arr_merge2_13__0 (GND0), .d_arr_merge2_14__31 (GND0), .d_arr_merge2_14__30 (
               GND0), .d_arr_merge2_14__29 (GND0), .d_arr_merge2_14__28 (GND0), 
               .d_arr_merge2_14__27 (GND0), .d_arr_merge2_14__26 (GND0), .d_arr_merge2_14__25 (
               GND0), .d_arr_merge2_14__24 (GND0), .d_arr_merge2_14__23 (GND0), 
               .d_arr_merge2_14__22 (GND0), .d_arr_merge2_14__21 (GND0), .d_arr_merge2_14__20 (
               GND0), .d_arr_merge2_14__19 (GND0), .d_arr_merge2_14__18 (GND0), 
               .d_arr_merge2_14__17 (GND0), .d_arr_merge2_14__16 (GND0), .d_arr_merge2_14__15 (
               GND0), .d_arr_merge2_14__14 (GND0), .d_arr_merge2_14__13 (GND0), 
               .d_arr_merge2_14__12 (GND0), .d_arr_merge2_14__11 (GND0), .d_arr_merge2_14__10 (
               GND0), .d_arr_merge2_14__9 (GND0), .d_arr_merge2_14__8 (GND0), .d_arr_merge2_14__7 (
               GND0), .d_arr_merge2_14__6 (GND0), .d_arr_merge2_14__5 (GND0), .d_arr_merge2_14__4 (
               GND0), .d_arr_merge2_14__3 (GND0), .d_arr_merge2_14__2 (GND0), .d_arr_merge2_14__1 (
               GND0), .d_arr_merge2_14__0 (GND0), .d_arr_merge2_15__31 (GND0), .d_arr_merge2_15__30 (
               GND0), .d_arr_merge2_15__29 (GND0), .d_arr_merge2_15__28 (GND0), 
               .d_arr_merge2_15__27 (GND0), .d_arr_merge2_15__26 (GND0), .d_arr_merge2_15__25 (
               GND0), .d_arr_merge2_15__24 (GND0), .d_arr_merge2_15__23 (GND0), 
               .d_arr_merge2_15__22 (GND0), .d_arr_merge2_15__21 (GND0), .d_arr_merge2_15__20 (
               GND0), .d_arr_merge2_15__19 (GND0), .d_arr_merge2_15__18 (GND0), 
               .d_arr_merge2_15__17 (GND0), .d_arr_merge2_15__16 (GND0), .d_arr_merge2_15__15 (
               GND0), .d_arr_merge2_15__14 (GND0), .d_arr_merge2_15__13 (GND0), 
               .d_arr_merge2_15__12 (GND0), .d_arr_merge2_15__11 (GND0), .d_arr_merge2_15__10 (
               GND0), .d_arr_merge2_15__9 (GND0), .d_arr_merge2_15__8 (GND0), .d_arr_merge2_15__7 (
               GND0), .d_arr_merge2_15__6 (GND0), .d_arr_merge2_15__5 (GND0), .d_arr_merge2_15__4 (
               GND0), .d_arr_merge2_15__3 (GND0), .d_arr_merge2_15__2 (GND0), .d_arr_merge2_15__1 (
               GND0), .d_arr_merge2_15__0 (GND0), .d_arr_merge2_16__31 (GND0), .d_arr_merge2_16__30 (
               GND0), .d_arr_merge2_16__29 (GND0), .d_arr_merge2_16__28 (GND0), 
               .d_arr_merge2_16__27 (GND0), .d_arr_merge2_16__26 (GND0), .d_arr_merge2_16__25 (
               GND0), .d_arr_merge2_16__24 (GND0), .d_arr_merge2_16__23 (GND0), 
               .d_arr_merge2_16__22 (GND0), .d_arr_merge2_16__21 (GND0), .d_arr_merge2_16__20 (
               GND0), .d_arr_merge2_16__19 (GND0), .d_arr_merge2_16__18 (GND0), 
               .d_arr_merge2_16__17 (GND0), .d_arr_merge2_16__16 (GND0), .d_arr_merge2_16__15 (
               GND0), .d_arr_merge2_16__14 (GND0), .d_arr_merge2_16__13 (GND0), 
               .d_arr_merge2_16__12 (GND0), .d_arr_merge2_16__11 (GND0), .d_arr_merge2_16__10 (
               GND0), .d_arr_merge2_16__9 (GND0), .d_arr_merge2_16__8 (GND0), .d_arr_merge2_16__7 (
               GND0), .d_arr_merge2_16__6 (GND0), .d_arr_merge2_16__5 (GND0), .d_arr_merge2_16__4 (
               GND0), .d_arr_merge2_16__3 (GND0), .d_arr_merge2_16__2 (GND0), .d_arr_merge2_16__1 (
               GND0), .d_arr_merge2_16__0 (GND0), .d_arr_merge2_17__31 (GND0), .d_arr_merge2_17__30 (
               GND0), .d_arr_merge2_17__29 (GND0), .d_arr_merge2_17__28 (GND0), 
               .d_arr_merge2_17__27 (GND0), .d_arr_merge2_17__26 (GND0), .d_arr_merge2_17__25 (
               GND0), .d_arr_merge2_17__24 (GND0), .d_arr_merge2_17__23 (GND0), 
               .d_arr_merge2_17__22 (GND0), .d_arr_merge2_17__21 (GND0), .d_arr_merge2_17__20 (
               GND0), .d_arr_merge2_17__19 (GND0), .d_arr_merge2_17__18 (GND0), 
               .d_arr_merge2_17__17 (GND0), .d_arr_merge2_17__16 (GND0), .d_arr_merge2_17__15 (
               GND0), .d_arr_merge2_17__14 (GND0), .d_arr_merge2_17__13 (GND0), 
               .d_arr_merge2_17__12 (GND0), .d_arr_merge2_17__11 (GND0), .d_arr_merge2_17__10 (
               GND0), .d_arr_merge2_17__9 (GND0), .d_arr_merge2_17__8 (GND0), .d_arr_merge2_17__7 (
               GND0), .d_arr_merge2_17__6 (GND0), .d_arr_merge2_17__5 (GND0), .d_arr_merge2_17__4 (
               GND0), .d_arr_merge2_17__3 (GND0), .d_arr_merge2_17__2 (GND0), .d_arr_merge2_17__1 (
               GND0), .d_arr_merge2_17__0 (GND0), .d_arr_merge2_18__31 (GND0), .d_arr_merge2_18__30 (
               GND0), .d_arr_merge2_18__29 (GND0), .d_arr_merge2_18__28 (GND0), 
               .d_arr_merge2_18__27 (GND0), .d_arr_merge2_18__26 (GND0), .d_arr_merge2_18__25 (
               GND0), .d_arr_merge2_18__24 (GND0), .d_arr_merge2_18__23 (GND0), 
               .d_arr_merge2_18__22 (GND0), .d_arr_merge2_18__21 (GND0), .d_arr_merge2_18__20 (
               GND0), .d_arr_merge2_18__19 (GND0), .d_arr_merge2_18__18 (GND0), 
               .d_arr_merge2_18__17 (GND0), .d_arr_merge2_18__16 (GND0), .d_arr_merge2_18__15 (
               GND0), .d_arr_merge2_18__14 (GND0), .d_arr_merge2_18__13 (GND0), 
               .d_arr_merge2_18__12 (GND0), .d_arr_merge2_18__11 (GND0), .d_arr_merge2_18__10 (
               GND0), .d_arr_merge2_18__9 (GND0), .d_arr_merge2_18__8 (GND0), .d_arr_merge2_18__7 (
               GND0), .d_arr_merge2_18__6 (GND0), .d_arr_merge2_18__5 (GND0), .d_arr_merge2_18__4 (
               GND0), .d_arr_merge2_18__3 (GND0), .d_arr_merge2_18__2 (GND0), .d_arr_merge2_18__1 (
               GND0), .d_arr_merge2_18__0 (GND0), .d_arr_merge2_19__31 (GND0), .d_arr_merge2_19__30 (
               GND0), .d_arr_merge2_19__29 (GND0), .d_arr_merge2_19__28 (GND0), 
               .d_arr_merge2_19__27 (GND0), .d_arr_merge2_19__26 (GND0), .d_arr_merge2_19__25 (
               GND0), .d_arr_merge2_19__24 (GND0), .d_arr_merge2_19__23 (GND0), 
               .d_arr_merge2_19__22 (GND0), .d_arr_merge2_19__21 (GND0), .d_arr_merge2_19__20 (
               GND0), .d_arr_merge2_19__19 (GND0), .d_arr_merge2_19__18 (GND0), 
               .d_arr_merge2_19__17 (GND0), .d_arr_merge2_19__16 (GND0), .d_arr_merge2_19__15 (
               GND0), .d_arr_merge2_19__14 (GND0), .d_arr_merge2_19__13 (GND0), 
               .d_arr_merge2_19__12 (GND0), .d_arr_merge2_19__11 (GND0), .d_arr_merge2_19__10 (
               GND0), .d_arr_merge2_19__9 (GND0), .d_arr_merge2_19__8 (GND0), .d_arr_merge2_19__7 (
               GND0), .d_arr_merge2_19__6 (GND0), .d_arr_merge2_19__5 (GND0), .d_arr_merge2_19__4 (
               GND0), .d_arr_merge2_19__3 (GND0), .d_arr_merge2_19__2 (GND0), .d_arr_merge2_19__1 (
               GND0), .d_arr_merge2_19__0 (GND0), .d_arr_merge2_20__31 (GND0), .d_arr_merge2_20__30 (
               GND0), .d_arr_merge2_20__29 (GND0), .d_arr_merge2_20__28 (GND0), 
               .d_arr_merge2_20__27 (GND0), .d_arr_merge2_20__26 (GND0), .d_arr_merge2_20__25 (
               GND0), .d_arr_merge2_20__24 (GND0), .d_arr_merge2_20__23 (GND0), 
               .d_arr_merge2_20__22 (GND0), .d_arr_merge2_20__21 (GND0), .d_arr_merge2_20__20 (
               GND0), .d_arr_merge2_20__19 (GND0), .d_arr_merge2_20__18 (GND0), 
               .d_arr_merge2_20__17 (GND0), .d_arr_merge2_20__16 (GND0), .d_arr_merge2_20__15 (
               GND0), .d_arr_merge2_20__14 (GND0), .d_arr_merge2_20__13 (GND0), 
               .d_arr_merge2_20__12 (GND0), .d_arr_merge2_20__11 (GND0), .d_arr_merge2_20__10 (
               GND0), .d_arr_merge2_20__9 (GND0), .d_arr_merge2_20__8 (GND0), .d_arr_merge2_20__7 (
               GND0), .d_arr_merge2_20__6 (GND0), .d_arr_merge2_20__5 (GND0), .d_arr_merge2_20__4 (
               GND0), .d_arr_merge2_20__3 (GND0), .d_arr_merge2_20__2 (GND0), .d_arr_merge2_20__1 (
               GND0), .d_arr_merge2_20__0 (GND0), .d_arr_merge2_21__31 (GND0), .d_arr_merge2_21__30 (
               GND0), .d_arr_merge2_21__29 (GND0), .d_arr_merge2_21__28 (GND0), 
               .d_arr_merge2_21__27 (GND0), .d_arr_merge2_21__26 (GND0), .d_arr_merge2_21__25 (
               GND0), .d_arr_merge2_21__24 (GND0), .d_arr_merge2_21__23 (GND0), 
               .d_arr_merge2_21__22 (GND0), .d_arr_merge2_21__21 (GND0), .d_arr_merge2_21__20 (
               GND0), .d_arr_merge2_21__19 (GND0), .d_arr_merge2_21__18 (GND0), 
               .d_arr_merge2_21__17 (GND0), .d_arr_merge2_21__16 (GND0), .d_arr_merge2_21__15 (
               GND0), .d_arr_merge2_21__14 (GND0), .d_arr_merge2_21__13 (GND0), 
               .d_arr_merge2_21__12 (GND0), .d_arr_merge2_21__11 (GND0), .d_arr_merge2_21__10 (
               GND0), .d_arr_merge2_21__9 (GND0), .d_arr_merge2_21__8 (GND0), .d_arr_merge2_21__7 (
               GND0), .d_arr_merge2_21__6 (GND0), .d_arr_merge2_21__5 (GND0), .d_arr_merge2_21__4 (
               GND0), .d_arr_merge2_21__3 (GND0), .d_arr_merge2_21__2 (GND0), .d_arr_merge2_21__1 (
               GND0), .d_arr_merge2_21__0 (GND0), .d_arr_merge2_22__31 (GND0), .d_arr_merge2_22__30 (
               GND0), .d_arr_merge2_22__29 (GND0), .d_arr_merge2_22__28 (GND0), 
               .d_arr_merge2_22__27 (GND0), .d_arr_merge2_22__26 (GND0), .d_arr_merge2_22__25 (
               GND0), .d_arr_merge2_22__24 (GND0), .d_arr_merge2_22__23 (GND0), 
               .d_arr_merge2_22__22 (GND0), .d_arr_merge2_22__21 (GND0), .d_arr_merge2_22__20 (
               GND0), .d_arr_merge2_22__19 (GND0), .d_arr_merge2_22__18 (GND0), 
               .d_arr_merge2_22__17 (GND0), .d_arr_merge2_22__16 (GND0), .d_arr_merge2_22__15 (
               GND0), .d_arr_merge2_22__14 (GND0), .d_arr_merge2_22__13 (GND0), 
               .d_arr_merge2_22__12 (GND0), .d_arr_merge2_22__11 (GND0), .d_arr_merge2_22__10 (
               GND0), .d_arr_merge2_22__9 (GND0), .d_arr_merge2_22__8 (GND0), .d_arr_merge2_22__7 (
               GND0), .d_arr_merge2_22__6 (GND0), .d_arr_merge2_22__5 (GND0), .d_arr_merge2_22__4 (
               GND0), .d_arr_merge2_22__3 (GND0), .d_arr_merge2_22__2 (GND0), .d_arr_merge2_22__1 (
               GND0), .d_arr_merge2_22__0 (GND0), .d_arr_merge2_23__31 (GND0), .d_arr_merge2_23__30 (
               GND0), .d_arr_merge2_23__29 (GND0), .d_arr_merge2_23__28 (GND0), 
               .d_arr_merge2_23__27 (GND0), .d_arr_merge2_23__26 (GND0), .d_arr_merge2_23__25 (
               GND0), .d_arr_merge2_23__24 (GND0), .d_arr_merge2_23__23 (GND0), 
               .d_arr_merge2_23__22 (GND0), .d_arr_merge2_23__21 (GND0), .d_arr_merge2_23__20 (
               GND0), .d_arr_merge2_23__19 (GND0), .d_arr_merge2_23__18 (GND0), 
               .d_arr_merge2_23__17 (GND0), .d_arr_merge2_23__16 (GND0), .d_arr_merge2_23__15 (
               GND0), .d_arr_merge2_23__14 (GND0), .d_arr_merge2_23__13 (GND0), 
               .d_arr_merge2_23__12 (GND0), .d_arr_merge2_23__11 (GND0), .d_arr_merge2_23__10 (
               GND0), .d_arr_merge2_23__9 (GND0), .d_arr_merge2_23__8 (GND0), .d_arr_merge2_23__7 (
               GND0), .d_arr_merge2_23__6 (GND0), .d_arr_merge2_23__5 (GND0), .d_arr_merge2_23__4 (
               GND0), .d_arr_merge2_23__3 (GND0), .d_arr_merge2_23__2 (GND0), .d_arr_merge2_23__1 (
               GND0), .d_arr_merge2_23__0 (GND0), .d_arr_merge2_24__31 (GND0), .d_arr_merge2_24__30 (
               GND0), .d_arr_merge2_24__29 (GND0), .d_arr_merge2_24__28 (GND0), 
               .d_arr_merge2_24__27 (GND0), .d_arr_merge2_24__26 (GND0), .d_arr_merge2_24__25 (
               GND0), .d_arr_merge2_24__24 (GND0), .d_arr_merge2_24__23 (GND0), 
               .d_arr_merge2_24__22 (GND0), .d_arr_merge2_24__21 (GND0), .d_arr_merge2_24__20 (
               GND0), .d_arr_merge2_24__19 (GND0), .d_arr_merge2_24__18 (GND0), 
               .d_arr_merge2_24__17 (GND0), .d_arr_merge2_24__16 (GND0), .d_arr_merge2_24__15 (
               GND0), .d_arr_merge2_24__14 (GND0), .d_arr_merge2_24__13 (GND0), 
               .d_arr_merge2_24__12 (GND0), .d_arr_merge2_24__11 (GND0), .d_arr_merge2_24__10 (
               GND0), .d_arr_merge2_24__9 (GND0), .d_arr_merge2_24__8 (GND0), .d_arr_merge2_24__7 (
               GND0), .d_arr_merge2_24__6 (GND0), .d_arr_merge2_24__5 (GND0), .d_arr_merge2_24__4 (
               GND0), .d_arr_merge2_24__3 (GND0), .d_arr_merge2_24__2 (GND0), .d_arr_merge2_24__1 (
               GND0), .d_arr_merge2_24__0 (GND0), .d_arr_relu_0__31 (
               d_arr_relu_0__31), .d_arr_relu_0__30 (d_arr_relu_0__30), .d_arr_relu_0__29 (
               d_arr_relu_0__29), .d_arr_relu_0__28 (d_arr_relu_0__28), .d_arr_relu_0__27 (
               d_arr_relu_0__27), .d_arr_relu_0__26 (d_arr_relu_0__26), .d_arr_relu_0__25 (
               d_arr_relu_0__25), .d_arr_relu_0__24 (d_arr_relu_0__24), .d_arr_relu_0__23 (
               d_arr_relu_0__23), .d_arr_relu_0__22 (d_arr_relu_0__22), .d_arr_relu_0__21 (
               d_arr_relu_0__21), .d_arr_relu_0__20 (d_arr_relu_0__20), .d_arr_relu_0__19 (
               d_arr_relu_0__19), .d_arr_relu_0__18 (d_arr_relu_0__18), .d_arr_relu_0__17 (
               d_arr_relu_0__17), .d_arr_relu_0__16 (d_arr_relu_0__16), .d_arr_relu_0__15 (
               GND0), .d_arr_relu_0__14 (d_arr_relu_0__14), .d_arr_relu_0__13 (
               d_arr_relu_0__13), .d_arr_relu_0__12 (d_arr_relu_0__12), .d_arr_relu_0__11 (
               d_arr_relu_0__11), .d_arr_relu_0__10 (d_arr_relu_0__10), .d_arr_relu_0__9 (
               d_arr_relu_0__9), .d_arr_relu_0__8 (d_arr_relu_0__8), .d_arr_relu_0__7 (
               d_arr_relu_0__7), .d_arr_relu_0__6 (d_arr_relu_0__6), .d_arr_relu_0__5 (
               d_arr_relu_0__5), .d_arr_relu_0__4 (d_arr_relu_0__4), .d_arr_relu_0__3 (
               d_arr_relu_0__3), .d_arr_relu_0__2 (d_arr_relu_0__2), .d_arr_relu_0__1 (
               d_arr_relu_0__1), .d_arr_relu_0__0 (d_arr_relu_0__0), .d_arr_relu_1__31 (
               d_arr_relu_1__31), .d_arr_relu_1__30 (d_arr_relu_1__30), .d_arr_relu_1__29 (
               d_arr_relu_1__29), .d_arr_relu_1__28 (d_arr_relu_1__28), .d_arr_relu_1__27 (
               d_arr_relu_1__27), .d_arr_relu_1__26 (d_arr_relu_1__26), .d_arr_relu_1__25 (
               d_arr_relu_1__25), .d_arr_relu_1__24 (d_arr_relu_1__24), .d_arr_relu_1__23 (
               d_arr_relu_1__23), .d_arr_relu_1__22 (d_arr_relu_1__22), .d_arr_relu_1__21 (
               d_arr_relu_1__21), .d_arr_relu_1__20 (d_arr_relu_1__20), .d_arr_relu_1__19 (
               d_arr_relu_1__19), .d_arr_relu_1__18 (d_arr_relu_1__18), .d_arr_relu_1__17 (
               d_arr_relu_1__17), .d_arr_relu_1__16 (d_arr_relu_1__16), .d_arr_relu_1__15 (
               GND0), .d_arr_relu_1__14 (d_arr_relu_1__14), .d_arr_relu_1__13 (
               d_arr_relu_1__13), .d_arr_relu_1__12 (d_arr_relu_1__12), .d_arr_relu_1__11 (
               d_arr_relu_1__11), .d_arr_relu_1__10 (d_arr_relu_1__10), .d_arr_relu_1__9 (
               d_arr_relu_1__9), .d_arr_relu_1__8 (d_arr_relu_1__8), .d_arr_relu_1__7 (
               d_arr_relu_1__7), .d_arr_relu_1__6 (d_arr_relu_1__6), .d_arr_relu_1__5 (
               d_arr_relu_1__5), .d_arr_relu_1__4 (d_arr_relu_1__4), .d_arr_relu_1__3 (
               d_arr_relu_1__3), .d_arr_relu_1__2 (d_arr_relu_1__2), .d_arr_relu_1__1 (
               d_arr_relu_1__1), .d_arr_relu_1__0 (d_arr_relu_1__0), .d_arr_relu_2__31 (
               GND0), .d_arr_relu_2__30 (GND0), .d_arr_relu_2__29 (GND0), .d_arr_relu_2__28 (
               GND0), .d_arr_relu_2__27 (GND0), .d_arr_relu_2__26 (GND0), .d_arr_relu_2__25 (
               GND0), .d_arr_relu_2__24 (GND0), .d_arr_relu_2__23 (GND0), .d_arr_relu_2__22 (
               GND0), .d_arr_relu_2__21 (GND0), .d_arr_relu_2__20 (GND0), .d_arr_relu_2__19 (
               GND0), .d_arr_relu_2__18 (GND0), .d_arr_relu_2__17 (GND0), .d_arr_relu_2__16 (
               GND0), .d_arr_relu_2__15 (GND0), .d_arr_relu_2__14 (GND0), .d_arr_relu_2__13 (
               GND0), .d_arr_relu_2__12 (GND0), .d_arr_relu_2__11 (GND0), .d_arr_relu_2__10 (
               GND0), .d_arr_relu_2__9 (GND0), .d_arr_relu_2__8 (GND0), .d_arr_relu_2__7 (
               GND0), .d_arr_relu_2__6 (GND0), .d_arr_relu_2__5 (GND0), .d_arr_relu_2__4 (
               GND0), .d_arr_relu_2__3 (GND0), .d_arr_relu_2__2 (GND0), .d_arr_relu_2__1 (
               GND0), .d_arr_relu_2__0 (GND0), .d_arr_relu_3__31 (GND0), .d_arr_relu_3__30 (
               GND0), .d_arr_relu_3__29 (GND0), .d_arr_relu_3__28 (GND0), .d_arr_relu_3__27 (
               GND0), .d_arr_relu_3__26 (GND0), .d_arr_relu_3__25 (GND0), .d_arr_relu_3__24 (
               GND0), .d_arr_relu_3__23 (GND0), .d_arr_relu_3__22 (GND0), .d_arr_relu_3__21 (
               GND0), .d_arr_relu_3__20 (GND0), .d_arr_relu_3__19 (GND0), .d_arr_relu_3__18 (
               GND0), .d_arr_relu_3__17 (GND0), .d_arr_relu_3__16 (GND0), .d_arr_relu_3__15 (
               GND0), .d_arr_relu_3__14 (GND0), .d_arr_relu_3__13 (GND0), .d_arr_relu_3__12 (
               GND0), .d_arr_relu_3__11 (GND0), .d_arr_relu_3__10 (GND0), .d_arr_relu_3__9 (
               GND0), .d_arr_relu_3__8 (GND0), .d_arr_relu_3__7 (GND0), .d_arr_relu_3__6 (
               GND0), .d_arr_relu_3__5 (GND0), .d_arr_relu_3__4 (GND0), .d_arr_relu_3__3 (
               GND0), .d_arr_relu_3__2 (GND0), .d_arr_relu_3__1 (GND0), .d_arr_relu_3__0 (
               GND0), .d_arr_relu_4__31 (GND0), .d_arr_relu_4__30 (GND0), .d_arr_relu_4__29 (
               GND0), .d_arr_relu_4__28 (GND0), .d_arr_relu_4__27 (GND0), .d_arr_relu_4__26 (
               GND0), .d_arr_relu_4__25 (GND0), .d_arr_relu_4__24 (GND0), .d_arr_relu_4__23 (
               GND0), .d_arr_relu_4__22 (GND0), .d_arr_relu_4__21 (GND0), .d_arr_relu_4__20 (
               GND0), .d_arr_relu_4__19 (GND0), .d_arr_relu_4__18 (GND0), .d_arr_relu_4__17 (
               GND0), .d_arr_relu_4__16 (GND0), .d_arr_relu_4__15 (GND0), .d_arr_relu_4__14 (
               GND0), .d_arr_relu_4__13 (GND0), .d_arr_relu_4__12 (GND0), .d_arr_relu_4__11 (
               GND0), .d_arr_relu_4__10 (GND0), .d_arr_relu_4__9 (GND0), .d_arr_relu_4__8 (
               GND0), .d_arr_relu_4__7 (GND0), .d_arr_relu_4__6 (GND0), .d_arr_relu_4__5 (
               GND0), .d_arr_relu_4__4 (GND0), .d_arr_relu_4__3 (GND0), .d_arr_relu_4__2 (
               GND0), .d_arr_relu_4__1 (GND0), .d_arr_relu_4__0 (GND0), .d_arr_relu_5__31 (
               GND0), .d_arr_relu_5__30 (GND0), .d_arr_relu_5__29 (GND0), .d_arr_relu_5__28 (
               GND0), .d_arr_relu_5__27 (GND0), .d_arr_relu_5__26 (GND0), .d_arr_relu_5__25 (
               GND0), .d_arr_relu_5__24 (GND0), .d_arr_relu_5__23 (GND0), .d_arr_relu_5__22 (
               GND0), .d_arr_relu_5__21 (GND0), .d_arr_relu_5__20 (GND0), .d_arr_relu_5__19 (
               GND0), .d_arr_relu_5__18 (GND0), .d_arr_relu_5__17 (GND0), .d_arr_relu_5__16 (
               GND0), .d_arr_relu_5__15 (GND0), .d_arr_relu_5__14 (GND0), .d_arr_relu_5__13 (
               GND0), .d_arr_relu_5__12 (GND0), .d_arr_relu_5__11 (GND0), .d_arr_relu_5__10 (
               GND0), .d_arr_relu_5__9 (GND0), .d_arr_relu_5__8 (GND0), .d_arr_relu_5__7 (
               GND0), .d_arr_relu_5__6 (GND0), .d_arr_relu_5__5 (GND0), .d_arr_relu_5__4 (
               GND0), .d_arr_relu_5__3 (GND0), .d_arr_relu_5__2 (GND0), .d_arr_relu_5__1 (
               GND0), .d_arr_relu_5__0 (GND0), .d_arr_relu_6__31 (GND0), .d_arr_relu_6__30 (
               GND0), .d_arr_relu_6__29 (GND0), .d_arr_relu_6__28 (GND0), .d_arr_relu_6__27 (
               GND0), .d_arr_relu_6__26 (GND0), .d_arr_relu_6__25 (GND0), .d_arr_relu_6__24 (
               GND0), .d_arr_relu_6__23 (GND0), .d_arr_relu_6__22 (GND0), .d_arr_relu_6__21 (
               GND0), .d_arr_relu_6__20 (GND0), .d_arr_relu_6__19 (GND0), .d_arr_relu_6__18 (
               GND0), .d_arr_relu_6__17 (GND0), .d_arr_relu_6__16 (GND0), .d_arr_relu_6__15 (
               GND0), .d_arr_relu_6__14 (GND0), .d_arr_relu_6__13 (GND0), .d_arr_relu_6__12 (
               GND0), .d_arr_relu_6__11 (GND0), .d_arr_relu_6__10 (GND0), .d_arr_relu_6__9 (
               GND0), .d_arr_relu_6__8 (GND0), .d_arr_relu_6__7 (GND0), .d_arr_relu_6__6 (
               GND0), .d_arr_relu_6__5 (GND0), .d_arr_relu_6__4 (GND0), .d_arr_relu_6__3 (
               GND0), .d_arr_relu_6__2 (GND0), .d_arr_relu_6__1 (GND0), .d_arr_relu_6__0 (
               GND0), .d_arr_relu_7__31 (GND0), .d_arr_relu_7__30 (GND0), .d_arr_relu_7__29 (
               GND0), .d_arr_relu_7__28 (GND0), .d_arr_relu_7__27 (GND0), .d_arr_relu_7__26 (
               GND0), .d_arr_relu_7__25 (GND0), .d_arr_relu_7__24 (GND0), .d_arr_relu_7__23 (
               GND0), .d_arr_relu_7__22 (GND0), .d_arr_relu_7__21 (GND0), .d_arr_relu_7__20 (
               GND0), .d_arr_relu_7__19 (GND0), .d_arr_relu_7__18 (GND0), .d_arr_relu_7__17 (
               GND0), .d_arr_relu_7__16 (GND0), .d_arr_relu_7__15 (GND0), .d_arr_relu_7__14 (
               GND0), .d_arr_relu_7__13 (GND0), .d_arr_relu_7__12 (GND0), .d_arr_relu_7__11 (
               GND0), .d_arr_relu_7__10 (GND0), .d_arr_relu_7__9 (GND0), .d_arr_relu_7__8 (
               GND0), .d_arr_relu_7__7 (GND0), .d_arr_relu_7__6 (GND0), .d_arr_relu_7__5 (
               GND0), .d_arr_relu_7__4 (GND0), .d_arr_relu_7__3 (GND0), .d_arr_relu_7__2 (
               GND0), .d_arr_relu_7__1 (GND0), .d_arr_relu_7__0 (GND0), .d_arr_relu_8__31 (
               GND0), .d_arr_relu_8__30 (GND0), .d_arr_relu_8__29 (GND0), .d_arr_relu_8__28 (
               GND0), .d_arr_relu_8__27 (GND0), .d_arr_relu_8__26 (GND0), .d_arr_relu_8__25 (
               GND0), .d_arr_relu_8__24 (GND0), .d_arr_relu_8__23 (GND0), .d_arr_relu_8__22 (
               GND0), .d_arr_relu_8__21 (GND0), .d_arr_relu_8__20 (GND0), .d_arr_relu_8__19 (
               GND0), .d_arr_relu_8__18 (GND0), .d_arr_relu_8__17 (GND0), .d_arr_relu_8__16 (
               GND0), .d_arr_relu_8__15 (GND0), .d_arr_relu_8__14 (GND0), .d_arr_relu_8__13 (
               GND0), .d_arr_relu_8__12 (GND0), .d_arr_relu_8__11 (GND0), .d_arr_relu_8__10 (
               GND0), .d_arr_relu_8__9 (GND0), .d_arr_relu_8__8 (GND0), .d_arr_relu_8__7 (
               GND0), .d_arr_relu_8__6 (GND0), .d_arr_relu_8__5 (GND0), .d_arr_relu_8__4 (
               GND0), .d_arr_relu_8__3 (GND0), .d_arr_relu_8__2 (GND0), .d_arr_relu_8__1 (
               GND0), .d_arr_relu_8__0 (GND0), .d_arr_relu_9__31 (GND0), .d_arr_relu_9__30 (
               GND0), .d_arr_relu_9__29 (GND0), .d_arr_relu_9__28 (GND0), .d_arr_relu_9__27 (
               GND0), .d_arr_relu_9__26 (GND0), .d_arr_relu_9__25 (GND0), .d_arr_relu_9__24 (
               GND0), .d_arr_relu_9__23 (GND0), .d_arr_relu_9__22 (GND0), .d_arr_relu_9__21 (
               GND0), .d_arr_relu_9__20 (GND0), .d_arr_relu_9__19 (GND0), .d_arr_relu_9__18 (
               GND0), .d_arr_relu_9__17 (GND0), .d_arr_relu_9__16 (GND0), .d_arr_relu_9__15 (
               GND0), .d_arr_relu_9__14 (GND0), .d_arr_relu_9__13 (GND0), .d_arr_relu_9__12 (
               GND0), .d_arr_relu_9__11 (GND0), .d_arr_relu_9__10 (GND0), .d_arr_relu_9__9 (
               GND0), .d_arr_relu_9__8 (GND0), .d_arr_relu_9__7 (GND0), .d_arr_relu_9__6 (
               GND0), .d_arr_relu_9__5 (GND0), .d_arr_relu_9__4 (GND0), .d_arr_relu_9__3 (
               GND0), .d_arr_relu_9__2 (GND0), .d_arr_relu_9__1 (GND0), .d_arr_relu_9__0 (
               GND0), .d_arr_relu_10__31 (GND0), .d_arr_relu_10__30 (GND0), .d_arr_relu_10__29 (
               GND0), .d_arr_relu_10__28 (GND0), .d_arr_relu_10__27 (GND0), .d_arr_relu_10__26 (
               GND0), .d_arr_relu_10__25 (GND0), .d_arr_relu_10__24 (GND0), .d_arr_relu_10__23 (
               GND0), .d_arr_relu_10__22 (GND0), .d_arr_relu_10__21 (GND0), .d_arr_relu_10__20 (
               GND0), .d_arr_relu_10__19 (GND0), .d_arr_relu_10__18 (GND0), .d_arr_relu_10__17 (
               GND0), .d_arr_relu_10__16 (GND0), .d_arr_relu_10__15 (GND0), .d_arr_relu_10__14 (
               GND0), .d_arr_relu_10__13 (GND0), .d_arr_relu_10__12 (GND0), .d_arr_relu_10__11 (
               GND0), .d_arr_relu_10__10 (GND0), .d_arr_relu_10__9 (GND0), .d_arr_relu_10__8 (
               GND0), .d_arr_relu_10__7 (GND0), .d_arr_relu_10__6 (GND0), .d_arr_relu_10__5 (
               GND0), .d_arr_relu_10__4 (GND0), .d_arr_relu_10__3 (GND0), .d_arr_relu_10__2 (
               GND0), .d_arr_relu_10__1 (GND0), .d_arr_relu_10__0 (GND0), .d_arr_relu_11__31 (
               GND0), .d_arr_relu_11__30 (GND0), .d_arr_relu_11__29 (GND0), .d_arr_relu_11__28 (
               GND0), .d_arr_relu_11__27 (GND0), .d_arr_relu_11__26 (GND0), .d_arr_relu_11__25 (
               GND0), .d_arr_relu_11__24 (GND0), .d_arr_relu_11__23 (GND0), .d_arr_relu_11__22 (
               GND0), .d_arr_relu_11__21 (GND0), .d_arr_relu_11__20 (GND0), .d_arr_relu_11__19 (
               GND0), .d_arr_relu_11__18 (GND0), .d_arr_relu_11__17 (GND0), .d_arr_relu_11__16 (
               GND0), .d_arr_relu_11__15 (GND0), .d_arr_relu_11__14 (GND0), .d_arr_relu_11__13 (
               GND0), .d_arr_relu_11__12 (GND0), .d_arr_relu_11__11 (GND0), .d_arr_relu_11__10 (
               GND0), .d_arr_relu_11__9 (GND0), .d_arr_relu_11__8 (GND0), .d_arr_relu_11__7 (
               GND0), .d_arr_relu_11__6 (GND0), .d_arr_relu_11__5 (GND0), .d_arr_relu_11__4 (
               GND0), .d_arr_relu_11__3 (GND0), .d_arr_relu_11__2 (GND0), .d_arr_relu_11__1 (
               GND0), .d_arr_relu_11__0 (GND0), .d_arr_relu_12__31 (GND0), .d_arr_relu_12__30 (
               GND0), .d_arr_relu_12__29 (GND0), .d_arr_relu_12__28 (GND0), .d_arr_relu_12__27 (
               GND0), .d_arr_relu_12__26 (GND0), .d_arr_relu_12__25 (GND0), .d_arr_relu_12__24 (
               GND0), .d_arr_relu_12__23 (GND0), .d_arr_relu_12__22 (GND0), .d_arr_relu_12__21 (
               GND0), .d_arr_relu_12__20 (GND0), .d_arr_relu_12__19 (GND0), .d_arr_relu_12__18 (
               GND0), .d_arr_relu_12__17 (GND0), .d_arr_relu_12__16 (GND0), .d_arr_relu_12__15 (
               GND0), .d_arr_relu_12__14 (GND0), .d_arr_relu_12__13 (GND0), .d_arr_relu_12__12 (
               GND0), .d_arr_relu_12__11 (GND0), .d_arr_relu_12__10 (GND0), .d_arr_relu_12__9 (
               GND0), .d_arr_relu_12__8 (GND0), .d_arr_relu_12__7 (GND0), .d_arr_relu_12__6 (
               GND0), .d_arr_relu_12__5 (GND0), .d_arr_relu_12__4 (GND0), .d_arr_relu_12__3 (
               GND0), .d_arr_relu_12__2 (GND0), .d_arr_relu_12__1 (GND0), .d_arr_relu_12__0 (
               GND0), .d_arr_relu_13__31 (GND0), .d_arr_relu_13__30 (GND0), .d_arr_relu_13__29 (
               GND0), .d_arr_relu_13__28 (GND0), .d_arr_relu_13__27 (GND0), .d_arr_relu_13__26 (
               GND0), .d_arr_relu_13__25 (GND0), .d_arr_relu_13__24 (GND0), .d_arr_relu_13__23 (
               GND0), .d_arr_relu_13__22 (GND0), .d_arr_relu_13__21 (GND0), .d_arr_relu_13__20 (
               GND0), .d_arr_relu_13__19 (GND0), .d_arr_relu_13__18 (GND0), .d_arr_relu_13__17 (
               GND0), .d_arr_relu_13__16 (GND0), .d_arr_relu_13__15 (GND0), .d_arr_relu_13__14 (
               GND0), .d_arr_relu_13__13 (GND0), .d_arr_relu_13__12 (GND0), .d_arr_relu_13__11 (
               GND0), .d_arr_relu_13__10 (GND0), .d_arr_relu_13__9 (GND0), .d_arr_relu_13__8 (
               GND0), .d_arr_relu_13__7 (GND0), .d_arr_relu_13__6 (GND0), .d_arr_relu_13__5 (
               GND0), .d_arr_relu_13__4 (GND0), .d_arr_relu_13__3 (GND0), .d_arr_relu_13__2 (
               GND0), .d_arr_relu_13__1 (GND0), .d_arr_relu_13__0 (GND0), .d_arr_relu_14__31 (
               GND0), .d_arr_relu_14__30 (GND0), .d_arr_relu_14__29 (GND0), .d_arr_relu_14__28 (
               GND0), .d_arr_relu_14__27 (GND0), .d_arr_relu_14__26 (GND0), .d_arr_relu_14__25 (
               GND0), .d_arr_relu_14__24 (GND0), .d_arr_relu_14__23 (GND0), .d_arr_relu_14__22 (
               GND0), .d_arr_relu_14__21 (GND0), .d_arr_relu_14__20 (GND0), .d_arr_relu_14__19 (
               GND0), .d_arr_relu_14__18 (GND0), .d_arr_relu_14__17 (GND0), .d_arr_relu_14__16 (
               GND0), .d_arr_relu_14__15 (GND0), .d_arr_relu_14__14 (GND0), .d_arr_relu_14__13 (
               GND0), .d_arr_relu_14__12 (GND0), .d_arr_relu_14__11 (GND0), .d_arr_relu_14__10 (
               GND0), .d_arr_relu_14__9 (GND0), .d_arr_relu_14__8 (GND0), .d_arr_relu_14__7 (
               GND0), .d_arr_relu_14__6 (GND0), .d_arr_relu_14__5 (GND0), .d_arr_relu_14__4 (
               GND0), .d_arr_relu_14__3 (GND0), .d_arr_relu_14__2 (GND0), .d_arr_relu_14__1 (
               GND0), .d_arr_relu_14__0 (GND0), .d_arr_relu_15__31 (GND0), .d_arr_relu_15__30 (
               GND0), .d_arr_relu_15__29 (GND0), .d_arr_relu_15__28 (GND0), .d_arr_relu_15__27 (
               GND0), .d_arr_relu_15__26 (GND0), .d_arr_relu_15__25 (GND0), .d_arr_relu_15__24 (
               GND0), .d_arr_relu_15__23 (GND0), .d_arr_relu_15__22 (GND0), .d_arr_relu_15__21 (
               GND0), .d_arr_relu_15__20 (GND0), .d_arr_relu_15__19 (GND0), .d_arr_relu_15__18 (
               GND0), .d_arr_relu_15__17 (GND0), .d_arr_relu_15__16 (GND0), .d_arr_relu_15__15 (
               GND0), .d_arr_relu_15__14 (GND0), .d_arr_relu_15__13 (GND0), .d_arr_relu_15__12 (
               GND0), .d_arr_relu_15__11 (GND0), .d_arr_relu_15__10 (GND0), .d_arr_relu_15__9 (
               GND0), .d_arr_relu_15__8 (GND0), .d_arr_relu_15__7 (GND0), .d_arr_relu_15__6 (
               GND0), .d_arr_relu_15__5 (GND0), .d_arr_relu_15__4 (GND0), .d_arr_relu_15__3 (
               GND0), .d_arr_relu_15__2 (GND0), .d_arr_relu_15__1 (GND0), .d_arr_relu_15__0 (
               GND0), .d_arr_relu_16__31 (GND0), .d_arr_relu_16__30 (GND0), .d_arr_relu_16__29 (
               GND0), .d_arr_relu_16__28 (GND0), .d_arr_relu_16__27 (GND0), .d_arr_relu_16__26 (
               GND0), .d_arr_relu_16__25 (GND0), .d_arr_relu_16__24 (GND0), .d_arr_relu_16__23 (
               GND0), .d_arr_relu_16__22 (GND0), .d_arr_relu_16__21 (GND0), .d_arr_relu_16__20 (
               GND0), .d_arr_relu_16__19 (GND0), .d_arr_relu_16__18 (GND0), .d_arr_relu_16__17 (
               GND0), .d_arr_relu_16__16 (GND0), .d_arr_relu_16__15 (GND0), .d_arr_relu_16__14 (
               GND0), .d_arr_relu_16__13 (GND0), .d_arr_relu_16__12 (GND0), .d_arr_relu_16__11 (
               GND0), .d_arr_relu_16__10 (GND0), .d_arr_relu_16__9 (GND0), .d_arr_relu_16__8 (
               GND0), .d_arr_relu_16__7 (GND0), .d_arr_relu_16__6 (GND0), .d_arr_relu_16__5 (
               GND0), .d_arr_relu_16__4 (GND0), .d_arr_relu_16__3 (GND0), .d_arr_relu_16__2 (
               GND0), .d_arr_relu_16__1 (GND0), .d_arr_relu_16__0 (GND0), .d_arr_relu_17__31 (
               GND0), .d_arr_relu_17__30 (GND0), .d_arr_relu_17__29 (GND0), .d_arr_relu_17__28 (
               GND0), .d_arr_relu_17__27 (GND0), .d_arr_relu_17__26 (GND0), .d_arr_relu_17__25 (
               GND0), .d_arr_relu_17__24 (GND0), .d_arr_relu_17__23 (GND0), .d_arr_relu_17__22 (
               GND0), .d_arr_relu_17__21 (GND0), .d_arr_relu_17__20 (GND0), .d_arr_relu_17__19 (
               GND0), .d_arr_relu_17__18 (GND0), .d_arr_relu_17__17 (GND0), .d_arr_relu_17__16 (
               GND0), .d_arr_relu_17__15 (GND0), .d_arr_relu_17__14 (GND0), .d_arr_relu_17__13 (
               GND0), .d_arr_relu_17__12 (GND0), .d_arr_relu_17__11 (GND0), .d_arr_relu_17__10 (
               GND0), .d_arr_relu_17__9 (GND0), .d_arr_relu_17__8 (GND0), .d_arr_relu_17__7 (
               GND0), .d_arr_relu_17__6 (GND0), .d_arr_relu_17__5 (GND0), .d_arr_relu_17__4 (
               GND0), .d_arr_relu_17__3 (GND0), .d_arr_relu_17__2 (GND0), .d_arr_relu_17__1 (
               GND0), .d_arr_relu_17__0 (GND0), .d_arr_relu_18__31 (GND0), .d_arr_relu_18__30 (
               GND0), .d_arr_relu_18__29 (GND0), .d_arr_relu_18__28 (GND0), .d_arr_relu_18__27 (
               GND0), .d_arr_relu_18__26 (GND0), .d_arr_relu_18__25 (GND0), .d_arr_relu_18__24 (
               GND0), .d_arr_relu_18__23 (GND0), .d_arr_relu_18__22 (GND0), .d_arr_relu_18__21 (
               GND0), .d_arr_relu_18__20 (GND0), .d_arr_relu_18__19 (GND0), .d_arr_relu_18__18 (
               GND0), .d_arr_relu_18__17 (GND0), .d_arr_relu_18__16 (GND0), .d_arr_relu_18__15 (
               GND0), .d_arr_relu_18__14 (GND0), .d_arr_relu_18__13 (GND0), .d_arr_relu_18__12 (
               GND0), .d_arr_relu_18__11 (GND0), .d_arr_relu_18__10 (GND0), .d_arr_relu_18__9 (
               GND0), .d_arr_relu_18__8 (GND0), .d_arr_relu_18__7 (GND0), .d_arr_relu_18__6 (
               GND0), .d_arr_relu_18__5 (GND0), .d_arr_relu_18__4 (GND0), .d_arr_relu_18__3 (
               GND0), .d_arr_relu_18__2 (GND0), .d_arr_relu_18__1 (GND0), .d_arr_relu_18__0 (
               GND0), .d_arr_relu_19__31 (GND0), .d_arr_relu_19__30 (GND0), .d_arr_relu_19__29 (
               GND0), .d_arr_relu_19__28 (GND0), .d_arr_relu_19__27 (GND0), .d_arr_relu_19__26 (
               GND0), .d_arr_relu_19__25 (GND0), .d_arr_relu_19__24 (GND0), .d_arr_relu_19__23 (
               GND0), .d_arr_relu_19__22 (GND0), .d_arr_relu_19__21 (GND0), .d_arr_relu_19__20 (
               GND0), .d_arr_relu_19__19 (GND0), .d_arr_relu_19__18 (GND0), .d_arr_relu_19__17 (
               GND0), .d_arr_relu_19__16 (GND0), .d_arr_relu_19__15 (GND0), .d_arr_relu_19__14 (
               GND0), .d_arr_relu_19__13 (GND0), .d_arr_relu_19__12 (GND0), .d_arr_relu_19__11 (
               GND0), .d_arr_relu_19__10 (GND0), .d_arr_relu_19__9 (GND0), .d_arr_relu_19__8 (
               GND0), .d_arr_relu_19__7 (GND0), .d_arr_relu_19__6 (GND0), .d_arr_relu_19__5 (
               GND0), .d_arr_relu_19__4 (GND0), .d_arr_relu_19__3 (GND0), .d_arr_relu_19__2 (
               GND0), .d_arr_relu_19__1 (GND0), .d_arr_relu_19__0 (GND0), .d_arr_relu_20__31 (
               GND0), .d_arr_relu_20__30 (GND0), .d_arr_relu_20__29 (GND0), .d_arr_relu_20__28 (
               GND0), .d_arr_relu_20__27 (GND0), .d_arr_relu_20__26 (GND0), .d_arr_relu_20__25 (
               GND0), .d_arr_relu_20__24 (GND0), .d_arr_relu_20__23 (GND0), .d_arr_relu_20__22 (
               GND0), .d_arr_relu_20__21 (GND0), .d_arr_relu_20__20 (GND0), .d_arr_relu_20__19 (
               GND0), .d_arr_relu_20__18 (GND0), .d_arr_relu_20__17 (GND0), .d_arr_relu_20__16 (
               GND0), .d_arr_relu_20__15 (GND0), .d_arr_relu_20__14 (GND0), .d_arr_relu_20__13 (
               GND0), .d_arr_relu_20__12 (GND0), .d_arr_relu_20__11 (GND0), .d_arr_relu_20__10 (
               GND0), .d_arr_relu_20__9 (GND0), .d_arr_relu_20__8 (GND0), .d_arr_relu_20__7 (
               GND0), .d_arr_relu_20__6 (GND0), .d_arr_relu_20__5 (GND0), .d_arr_relu_20__4 (
               GND0), .d_arr_relu_20__3 (GND0), .d_arr_relu_20__2 (GND0), .d_arr_relu_20__1 (
               GND0), .d_arr_relu_20__0 (GND0), .d_arr_relu_21__31 (GND0), .d_arr_relu_21__30 (
               GND0), .d_arr_relu_21__29 (GND0), .d_arr_relu_21__28 (GND0), .d_arr_relu_21__27 (
               GND0), .d_arr_relu_21__26 (GND0), .d_arr_relu_21__25 (GND0), .d_arr_relu_21__24 (
               GND0), .d_arr_relu_21__23 (GND0), .d_arr_relu_21__22 (GND0), .d_arr_relu_21__21 (
               GND0), .d_arr_relu_21__20 (GND0), .d_arr_relu_21__19 (GND0), .d_arr_relu_21__18 (
               GND0), .d_arr_relu_21__17 (GND0), .d_arr_relu_21__16 (GND0), .d_arr_relu_21__15 (
               GND0), .d_arr_relu_21__14 (GND0), .d_arr_relu_21__13 (GND0), .d_arr_relu_21__12 (
               GND0), .d_arr_relu_21__11 (GND0), .d_arr_relu_21__10 (GND0), .d_arr_relu_21__9 (
               GND0), .d_arr_relu_21__8 (GND0), .d_arr_relu_21__7 (GND0), .d_arr_relu_21__6 (
               GND0), .d_arr_relu_21__5 (GND0), .d_arr_relu_21__4 (GND0), .d_arr_relu_21__3 (
               GND0), .d_arr_relu_21__2 (GND0), .d_arr_relu_21__1 (GND0), .d_arr_relu_21__0 (
               GND0), .d_arr_relu_22__31 (GND0), .d_arr_relu_22__30 (GND0), .d_arr_relu_22__29 (
               GND0), .d_arr_relu_22__28 (GND0), .d_arr_relu_22__27 (GND0), .d_arr_relu_22__26 (
               GND0), .d_arr_relu_22__25 (GND0), .d_arr_relu_22__24 (GND0), .d_arr_relu_22__23 (
               GND0), .d_arr_relu_22__22 (GND0), .d_arr_relu_22__21 (GND0), .d_arr_relu_22__20 (
               GND0), .d_arr_relu_22__19 (GND0), .d_arr_relu_22__18 (GND0), .d_arr_relu_22__17 (
               GND0), .d_arr_relu_22__16 (GND0), .d_arr_relu_22__15 (GND0), .d_arr_relu_22__14 (
               GND0), .d_arr_relu_22__13 (GND0), .d_arr_relu_22__12 (GND0), .d_arr_relu_22__11 (
               GND0), .d_arr_relu_22__10 (GND0), .d_arr_relu_22__9 (GND0), .d_arr_relu_22__8 (
               GND0), .d_arr_relu_22__7 (GND0), .d_arr_relu_22__6 (GND0), .d_arr_relu_22__5 (
               GND0), .d_arr_relu_22__4 (GND0), .d_arr_relu_22__3 (GND0), .d_arr_relu_22__2 (
               GND0), .d_arr_relu_22__1 (GND0), .d_arr_relu_22__0 (GND0), .d_arr_relu_23__31 (
               GND0), .d_arr_relu_23__30 (GND0), .d_arr_relu_23__29 (GND0), .d_arr_relu_23__28 (
               GND0), .d_arr_relu_23__27 (GND0), .d_arr_relu_23__26 (GND0), .d_arr_relu_23__25 (
               GND0), .d_arr_relu_23__24 (GND0), .d_arr_relu_23__23 (GND0), .d_arr_relu_23__22 (
               GND0), .d_arr_relu_23__21 (GND0), .d_arr_relu_23__20 (GND0), .d_arr_relu_23__19 (
               GND0), .d_arr_relu_23__18 (GND0), .d_arr_relu_23__17 (GND0), .d_arr_relu_23__16 (
               GND0), .d_arr_relu_23__15 (GND0), .d_arr_relu_23__14 (GND0), .d_arr_relu_23__13 (
               GND0), .d_arr_relu_23__12 (GND0), .d_arr_relu_23__11 (GND0), .d_arr_relu_23__10 (
               GND0), .d_arr_relu_23__9 (GND0), .d_arr_relu_23__8 (GND0), .d_arr_relu_23__7 (
               GND0), .d_arr_relu_23__6 (GND0), .d_arr_relu_23__5 (GND0), .d_arr_relu_23__4 (
               GND0), .d_arr_relu_23__3 (GND0), .d_arr_relu_23__2 (GND0), .d_arr_relu_23__1 (
               GND0), .d_arr_relu_23__0 (GND0), .d_arr_relu_24__31 (GND0), .d_arr_relu_24__30 (
               GND0), .d_arr_relu_24__29 (GND0), .d_arr_relu_24__28 (GND0), .d_arr_relu_24__27 (
               GND0), .d_arr_relu_24__26 (GND0), .d_arr_relu_24__25 (GND0), .d_arr_relu_24__24 (
               GND0), .d_arr_relu_24__23 (GND0), .d_arr_relu_24__22 (GND0), .d_arr_relu_24__21 (
               GND0), .d_arr_relu_24__20 (GND0), .d_arr_relu_24__19 (GND0), .d_arr_relu_24__18 (
               GND0), .d_arr_relu_24__17 (GND0), .d_arr_relu_24__16 (GND0), .d_arr_relu_24__15 (
               GND0), .d_arr_relu_24__14 (GND0), .d_arr_relu_24__13 (GND0), .d_arr_relu_24__12 (
               GND0), .d_arr_relu_24__11 (GND0), .d_arr_relu_24__10 (GND0), .d_arr_relu_24__9 (
               GND0), .d_arr_relu_24__8 (GND0), .d_arr_relu_24__7 (GND0), .d_arr_relu_24__6 (
               GND0), .d_arr_relu_24__5 (GND0), .d_arr_relu_24__4 (GND0), .d_arr_relu_24__3 (
               GND0), .d_arr_relu_24__2 (GND0), .d_arr_relu_24__1 (GND0), .d_arr_relu_24__0 (
               GND0), .sel_mux (counter_0), .sel_mul (nx16627), .sel_add (
               sel_add), .sel_merge1 (counter_13), .sel_merge2 (counter_14), .sel_relu (
               counter_15), .d_arr_0__31 (d_arr_0__31), .d_arr_0__30 (
               d_arr_0__30), .d_arr_0__29 (d_arr_0__29), .d_arr_0__28 (
               d_arr_0__28), .d_arr_0__27 (d_arr_0__27), .d_arr_0__26 (
               d_arr_0__26), .d_arr_0__25 (d_arr_0__25), .d_arr_0__24 (
               d_arr_0__24), .d_arr_0__23 (d_arr_0__23), .d_arr_0__22 (
               d_arr_0__22), .d_arr_0__21 (d_arr_0__21), .d_arr_0__20 (
               d_arr_0__20), .d_arr_0__19 (d_arr_0__19), .d_arr_0__18 (
               d_arr_0__18), .d_arr_0__17 (d_arr_0__17), .d_arr_0__16 (
               d_arr_0__16), .d_arr_0__15 (d_arr_0__15), .d_arr_0__14 (
               d_arr_0__14), .d_arr_0__13 (d_arr_0__13), .d_arr_0__12 (
               d_arr_0__12), .d_arr_0__11 (d_arr_0__11), .d_arr_0__10 (
               d_arr_0__10), .d_arr_0__9 (d_arr_0__9), .d_arr_0__8 (d_arr_0__8)
               , .d_arr_0__7 (d_arr_0__7), .d_arr_0__6 (d_arr_0__6), .d_arr_0__5 (
               d_arr_0__5), .d_arr_0__4 (d_arr_0__4), .d_arr_0__3 (d_arr_0__3), 
               .d_arr_0__2 (d_arr_0__2), .d_arr_0__1 (d_arr_0__1), .d_arr_0__0 (
               d_arr_0__0), .d_arr_1__31 (d_arr_1__31), .d_arr_1__30 (
               d_arr_1__30), .d_arr_1__29 (d_arr_1__29), .d_arr_1__28 (
               d_arr_1__28), .d_arr_1__27 (d_arr_1__27), .d_arr_1__26 (
               d_arr_1__26), .d_arr_1__25 (d_arr_1__25), .d_arr_1__24 (
               d_arr_1__24), .d_arr_1__23 (d_arr_1__23), .d_arr_1__22 (
               d_arr_1__22), .d_arr_1__21 (d_arr_1__21), .d_arr_1__20 (
               d_arr_1__20), .d_arr_1__19 (d_arr_1__19), .d_arr_1__18 (
               d_arr_1__18), .d_arr_1__17 (d_arr_1__17), .d_arr_1__16 (
               d_arr_1__16), .d_arr_1__15 (d_arr_1__15), .d_arr_1__14 (
               d_arr_1__14), .d_arr_1__13 (d_arr_1__13), .d_arr_1__12 (
               d_arr_1__12), .d_arr_1__11 (d_arr_1__11), .d_arr_1__10 (
               d_arr_1__10), .d_arr_1__9 (d_arr_1__9), .d_arr_1__8 (d_arr_1__8)
               , .d_arr_1__7 (d_arr_1__7), .d_arr_1__6 (d_arr_1__6), .d_arr_1__5 (
               d_arr_1__5), .d_arr_1__4 (d_arr_1__4), .d_arr_1__3 (d_arr_1__3), 
               .d_arr_1__2 (d_arr_1__2), .d_arr_1__1 (d_arr_1__1), .d_arr_1__0 (
               d_arr_1__0), .d_arr_2__31 (d_arr_2__31), .d_arr_2__30 (
               d_arr_2__30), .d_arr_2__29 (d_arr_2__29), .d_arr_2__28 (
               d_arr_2__28), .d_arr_2__27 (d_arr_2__27), .d_arr_2__26 (
               d_arr_2__26), .d_arr_2__25 (d_arr_2__25), .d_arr_2__24 (
               d_arr_2__24), .d_arr_2__23 (d_arr_2__23), .d_arr_2__22 (
               d_arr_2__22), .d_arr_2__21 (d_arr_2__21), .d_arr_2__20 (
               d_arr_2__20), .d_arr_2__19 (d_arr_2__19), .d_arr_2__18 (
               d_arr_2__18), .d_arr_2__17 (d_arr_2__17), .d_arr_2__16 (
               d_arr_2__16), .d_arr_2__15 (d_arr_2__15), .d_arr_2__14 (
               d_arr_2__14), .d_arr_2__13 (d_arr_2__13), .d_arr_2__12 (
               d_arr_2__12), .d_arr_2__11 (d_arr_2__11), .d_arr_2__10 (
               d_arr_2__10), .d_arr_2__9 (d_arr_2__9), .d_arr_2__8 (d_arr_2__8)
               , .d_arr_2__7 (d_arr_2__7), .d_arr_2__6 (d_arr_2__6), .d_arr_2__5 (
               d_arr_2__5), .d_arr_2__4 (d_arr_2__4), .d_arr_2__3 (d_arr_2__3), 
               .d_arr_2__2 (d_arr_2__2), .d_arr_2__1 (d_arr_2__1), .d_arr_2__0 (
               d_arr_2__0), .d_arr_3__31 (d_arr_3__31), .d_arr_3__30 (
               d_arr_3__30), .d_arr_3__29 (d_arr_3__29), .d_arr_3__28 (
               d_arr_3__28), .d_arr_3__27 (d_arr_3__27), .d_arr_3__26 (
               d_arr_3__26), .d_arr_3__25 (d_arr_3__25), .d_arr_3__24 (
               d_arr_3__24), .d_arr_3__23 (d_arr_3__23), .d_arr_3__22 (
               d_arr_3__22), .d_arr_3__21 (d_arr_3__21), .d_arr_3__20 (
               d_arr_3__20), .d_arr_3__19 (d_arr_3__19), .d_arr_3__18 (
               d_arr_3__18), .d_arr_3__17 (d_arr_3__17), .d_arr_3__16 (
               d_arr_3__16), .d_arr_3__15 (d_arr_3__15), .d_arr_3__14 (
               d_arr_3__14), .d_arr_3__13 (d_arr_3__13), .d_arr_3__12 (
               d_arr_3__12), .d_arr_3__11 (d_arr_3__11), .d_arr_3__10 (
               d_arr_3__10), .d_arr_3__9 (d_arr_3__9), .d_arr_3__8 (d_arr_3__8)
               , .d_arr_3__7 (d_arr_3__7), .d_arr_3__6 (d_arr_3__6), .d_arr_3__5 (
               d_arr_3__5), .d_arr_3__4 (d_arr_3__4), .d_arr_3__3 (d_arr_3__3), 
               .d_arr_3__2 (d_arr_3__2), .d_arr_3__1 (d_arr_3__1), .d_arr_3__0 (
               d_arr_3__0), .d_arr_4__31 (d_arr_4__31), .d_arr_4__30 (
               d_arr_4__30), .d_arr_4__29 (d_arr_4__29), .d_arr_4__28 (
               d_arr_4__28), .d_arr_4__27 (d_arr_4__27), .d_arr_4__26 (
               d_arr_4__26), .d_arr_4__25 (d_arr_4__25), .d_arr_4__24 (
               d_arr_4__24), .d_arr_4__23 (d_arr_4__23), .d_arr_4__22 (
               d_arr_4__22), .d_arr_4__21 (d_arr_4__21), .d_arr_4__20 (
               d_arr_4__20), .d_arr_4__19 (d_arr_4__19), .d_arr_4__18 (
               d_arr_4__18), .d_arr_4__17 (d_arr_4__17), .d_arr_4__16 (
               d_arr_4__16), .d_arr_4__15 (d_arr_4__15), .d_arr_4__14 (
               d_arr_4__14), .d_arr_4__13 (d_arr_4__13), .d_arr_4__12 (
               d_arr_4__12), .d_arr_4__11 (d_arr_4__11), .d_arr_4__10 (
               d_arr_4__10), .d_arr_4__9 (d_arr_4__9), .d_arr_4__8 (d_arr_4__8)
               , .d_arr_4__7 (d_arr_4__7), .d_arr_4__6 (d_arr_4__6), .d_arr_4__5 (
               d_arr_4__5), .d_arr_4__4 (d_arr_4__4), .d_arr_4__3 (d_arr_4__3), 
               .d_arr_4__2 (d_arr_4__2), .d_arr_4__1 (d_arr_4__1), .d_arr_4__0 (
               d_arr_4__0), .d_arr_5__31 (d_arr_5__31), .d_arr_5__30 (
               d_arr_5__30), .d_arr_5__29 (d_arr_5__29), .d_arr_5__28 (
               d_arr_5__28), .d_arr_5__27 (d_arr_5__27), .d_arr_5__26 (
               d_arr_5__26), .d_arr_5__25 (d_arr_5__25), .d_arr_5__24 (
               d_arr_5__24), .d_arr_5__23 (d_arr_5__23), .d_arr_5__22 (
               d_arr_5__22), .d_arr_5__21 (d_arr_5__21), .d_arr_5__20 (
               d_arr_5__20), .d_arr_5__19 (d_arr_5__19), .d_arr_5__18 (
               d_arr_5__18), .d_arr_5__17 (d_arr_5__17), .d_arr_5__16 (
               d_arr_5__16), .d_arr_5__15 (d_arr_5__15), .d_arr_5__14 (
               d_arr_5__14), .d_arr_5__13 (d_arr_5__13), .d_arr_5__12 (
               d_arr_5__12), .d_arr_5__11 (d_arr_5__11), .d_arr_5__10 (
               d_arr_5__10), .d_arr_5__9 (d_arr_5__9), .d_arr_5__8 (d_arr_5__8)
               , .d_arr_5__7 (d_arr_5__7), .d_arr_5__6 (d_arr_5__6), .d_arr_5__5 (
               d_arr_5__5), .d_arr_5__4 (d_arr_5__4), .d_arr_5__3 (d_arr_5__3), 
               .d_arr_5__2 (d_arr_5__2), .d_arr_5__1 (d_arr_5__1), .d_arr_5__0 (
               d_arr_5__0), .d_arr_6__31 (d_arr_6__31), .d_arr_6__30 (
               d_arr_6__30), .d_arr_6__29 (d_arr_6__29), .d_arr_6__28 (
               d_arr_6__28), .d_arr_6__27 (d_arr_6__27), .d_arr_6__26 (
               d_arr_6__26), .d_arr_6__25 (d_arr_6__25), .d_arr_6__24 (
               d_arr_6__24), .d_arr_6__23 (d_arr_6__23), .d_arr_6__22 (
               d_arr_6__22), .d_arr_6__21 (d_arr_6__21), .d_arr_6__20 (
               d_arr_6__20), .d_arr_6__19 (d_arr_6__19), .d_arr_6__18 (
               d_arr_6__18), .d_arr_6__17 (d_arr_6__17), .d_arr_6__16 (
               d_arr_6__16), .d_arr_6__15 (d_arr_6__15), .d_arr_6__14 (
               d_arr_6__14), .d_arr_6__13 (d_arr_6__13), .d_arr_6__12 (
               d_arr_6__12), .d_arr_6__11 (d_arr_6__11), .d_arr_6__10 (
               d_arr_6__10), .d_arr_6__9 (d_arr_6__9), .d_arr_6__8 (d_arr_6__8)
               , .d_arr_6__7 (d_arr_6__7), .d_arr_6__6 (d_arr_6__6), .d_arr_6__5 (
               d_arr_6__5), .d_arr_6__4 (d_arr_6__4), .d_arr_6__3 (d_arr_6__3), 
               .d_arr_6__2 (d_arr_6__2), .d_arr_6__1 (d_arr_6__1), .d_arr_6__0 (
               d_arr_6__0), .d_arr_7__31 (d_arr_7__31), .d_arr_7__30 (
               d_arr_7__30), .d_arr_7__29 (d_arr_7__29), .d_arr_7__28 (
               d_arr_7__28), .d_arr_7__27 (d_arr_7__27), .d_arr_7__26 (
               d_arr_7__26), .d_arr_7__25 (d_arr_7__25), .d_arr_7__24 (
               d_arr_7__24), .d_arr_7__23 (d_arr_7__23), .d_arr_7__22 (
               d_arr_7__22), .d_arr_7__21 (d_arr_7__21), .d_arr_7__20 (
               d_arr_7__20), .d_arr_7__19 (d_arr_7__19), .d_arr_7__18 (
               d_arr_7__18), .d_arr_7__17 (d_arr_7__17), .d_arr_7__16 (
               d_arr_7__16), .d_arr_7__15 (d_arr_7__15), .d_arr_7__14 (
               d_arr_7__14), .d_arr_7__13 (d_arr_7__13), .d_arr_7__12 (
               d_arr_7__12), .d_arr_7__11 (d_arr_7__11), .d_arr_7__10 (
               d_arr_7__10), .d_arr_7__9 (d_arr_7__9), .d_arr_7__8 (d_arr_7__8)
               , .d_arr_7__7 (d_arr_7__7), .d_arr_7__6 (d_arr_7__6), .d_arr_7__5 (
               d_arr_7__5), .d_arr_7__4 (d_arr_7__4), .d_arr_7__3 (d_arr_7__3), 
               .d_arr_7__2 (d_arr_7__2), .d_arr_7__1 (d_arr_7__1), .d_arr_7__0 (
               d_arr_7__0), .d_arr_8__31 (d_arr_8__31), .d_arr_8__30 (
               d_arr_8__30), .d_arr_8__29 (d_arr_8__29), .d_arr_8__28 (
               d_arr_8__28), .d_arr_8__27 (d_arr_8__27), .d_arr_8__26 (
               d_arr_8__26), .d_arr_8__25 (d_arr_8__25), .d_arr_8__24 (
               d_arr_8__24), .d_arr_8__23 (d_arr_8__23), .d_arr_8__22 (
               d_arr_8__22), .d_arr_8__21 (d_arr_8__21), .d_arr_8__20 (
               d_arr_8__20), .d_arr_8__19 (d_arr_8__19), .d_arr_8__18 (
               d_arr_8__18), .d_arr_8__17 (d_arr_8__17), .d_arr_8__16 (
               d_arr_8__16), .d_arr_8__15 (d_arr_8__15), .d_arr_8__14 (
               d_arr_8__14), .d_arr_8__13 (d_arr_8__13), .d_arr_8__12 (
               d_arr_8__12), .d_arr_8__11 (d_arr_8__11), .d_arr_8__10 (
               d_arr_8__10), .d_arr_8__9 (d_arr_8__9), .d_arr_8__8 (d_arr_8__8)
               , .d_arr_8__7 (d_arr_8__7), .d_arr_8__6 (d_arr_8__6), .d_arr_8__5 (
               d_arr_8__5), .d_arr_8__4 (d_arr_8__4), .d_arr_8__3 (d_arr_8__3), 
               .d_arr_8__2 (d_arr_8__2), .d_arr_8__1 (d_arr_8__1), .d_arr_8__0 (
               d_arr_8__0), .d_arr_9__31 (d_arr_9__31), .d_arr_9__30 (
               d_arr_9__30), .d_arr_9__29 (d_arr_9__29), .d_arr_9__28 (
               d_arr_9__28), .d_arr_9__27 (d_arr_9__27), .d_arr_9__26 (
               d_arr_9__26), .d_arr_9__25 (d_arr_9__25), .d_arr_9__24 (
               d_arr_9__24), .d_arr_9__23 (d_arr_9__23), .d_arr_9__22 (
               d_arr_9__22), .d_arr_9__21 (d_arr_9__21), .d_arr_9__20 (
               d_arr_9__20), .d_arr_9__19 (d_arr_9__19), .d_arr_9__18 (
               d_arr_9__18), .d_arr_9__17 (d_arr_9__17), .d_arr_9__16 (
               d_arr_9__16), .d_arr_9__15 (d_arr_9__15), .d_arr_9__14 (
               d_arr_9__14), .d_arr_9__13 (d_arr_9__13), .d_arr_9__12 (
               d_arr_9__12), .d_arr_9__11 (d_arr_9__11), .d_arr_9__10 (
               d_arr_9__10), .d_arr_9__9 (d_arr_9__9), .d_arr_9__8 (d_arr_9__8)
               , .d_arr_9__7 (d_arr_9__7), .d_arr_9__6 (d_arr_9__6), .d_arr_9__5 (
               d_arr_9__5), .d_arr_9__4 (d_arr_9__4), .d_arr_9__3 (d_arr_9__3), 
               .d_arr_9__2 (d_arr_9__2), .d_arr_9__1 (d_arr_9__1), .d_arr_9__0 (
               d_arr_9__0), .d_arr_10__31 (d_arr_10__31), .d_arr_10__30 (
               d_arr_10__30), .d_arr_10__29 (d_arr_10__29), .d_arr_10__28 (
               d_arr_10__28), .d_arr_10__27 (d_arr_10__27), .d_arr_10__26 (
               d_arr_10__26), .d_arr_10__25 (d_arr_10__25), .d_arr_10__24 (
               d_arr_10__24), .d_arr_10__23 (d_arr_10__23), .d_arr_10__22 (
               d_arr_10__22), .d_arr_10__21 (d_arr_10__21), .d_arr_10__20 (
               d_arr_10__20), .d_arr_10__19 (d_arr_10__19), .d_arr_10__18 (
               d_arr_10__18), .d_arr_10__17 (d_arr_10__17), .d_arr_10__16 (
               d_arr_10__16), .d_arr_10__15 (d_arr_10__15), .d_arr_10__14 (
               d_arr_10__14), .d_arr_10__13 (d_arr_10__13), .d_arr_10__12 (
               d_arr_10__12), .d_arr_10__11 (d_arr_10__11), .d_arr_10__10 (
               d_arr_10__10), .d_arr_10__9 (d_arr_10__9), .d_arr_10__8 (
               d_arr_10__8), .d_arr_10__7 (d_arr_10__7), .d_arr_10__6 (
               d_arr_10__6), .d_arr_10__5 (d_arr_10__5), .d_arr_10__4 (
               d_arr_10__4), .d_arr_10__3 (d_arr_10__3), .d_arr_10__2 (
               d_arr_10__2), .d_arr_10__1 (d_arr_10__1), .d_arr_10__0 (
               d_arr_10__0), .d_arr_11__31 (d_arr_11__31), .d_arr_11__30 (
               d_arr_11__30), .d_arr_11__29 (d_arr_11__29), .d_arr_11__28 (
               d_arr_11__28), .d_arr_11__27 (d_arr_11__27), .d_arr_11__26 (
               d_arr_11__26), .d_arr_11__25 (d_arr_11__25), .d_arr_11__24 (
               d_arr_11__24), .d_arr_11__23 (d_arr_11__23), .d_arr_11__22 (
               d_arr_11__22), .d_arr_11__21 (d_arr_11__21), .d_arr_11__20 (
               d_arr_11__20), .d_arr_11__19 (d_arr_11__19), .d_arr_11__18 (
               d_arr_11__18), .d_arr_11__17 (d_arr_11__17), .d_arr_11__16 (
               d_arr_11__16), .d_arr_11__15 (d_arr_11__15), .d_arr_11__14 (
               d_arr_11__14), .d_arr_11__13 (d_arr_11__13), .d_arr_11__12 (
               d_arr_11__12), .d_arr_11__11 (d_arr_11__11), .d_arr_11__10 (
               d_arr_11__10), .d_arr_11__9 (d_arr_11__9), .d_arr_11__8 (
               d_arr_11__8), .d_arr_11__7 (d_arr_11__7), .d_arr_11__6 (
               d_arr_11__6), .d_arr_11__5 (d_arr_11__5), .d_arr_11__4 (
               d_arr_11__4), .d_arr_11__3 (d_arr_11__3), .d_arr_11__2 (
               d_arr_11__2), .d_arr_11__1 (d_arr_11__1), .d_arr_11__0 (
               d_arr_11__0), .d_arr_12__31 (d_arr_12__31), .d_arr_12__30 (
               d_arr_12__30), .d_arr_12__29 (d_arr_12__29), .d_arr_12__28 (
               d_arr_12__28), .d_arr_12__27 (d_arr_12__27), .d_arr_12__26 (
               d_arr_12__26), .d_arr_12__25 (d_arr_12__25), .d_arr_12__24 (
               d_arr_12__24), .d_arr_12__23 (d_arr_12__23), .d_arr_12__22 (
               d_arr_12__22), .d_arr_12__21 (d_arr_12__21), .d_arr_12__20 (
               d_arr_12__20), .d_arr_12__19 (d_arr_12__19), .d_arr_12__18 (
               d_arr_12__18), .d_arr_12__17 (d_arr_12__17), .d_arr_12__16 (
               d_arr_12__16), .d_arr_12__15 (d_arr_12__15), .d_arr_12__14 (
               d_arr_12__14), .d_arr_12__13 (d_arr_12__13), .d_arr_12__12 (
               d_arr_12__12), .d_arr_12__11 (d_arr_12__11), .d_arr_12__10 (
               d_arr_12__10), .d_arr_12__9 (d_arr_12__9), .d_arr_12__8 (
               d_arr_12__8), .d_arr_12__7 (d_arr_12__7), .d_arr_12__6 (
               d_arr_12__6), .d_arr_12__5 (d_arr_12__5), .d_arr_12__4 (
               d_arr_12__4), .d_arr_12__3 (d_arr_12__3), .d_arr_12__2 (
               d_arr_12__2), .d_arr_12__1 (d_arr_12__1), .d_arr_12__0 (
               d_arr_12__0), .d_arr_13__31 (d_arr_13__31), .d_arr_13__30 (
               d_arr_13__30), .d_arr_13__29 (d_arr_13__29), .d_arr_13__28 (
               d_arr_13__28), .d_arr_13__27 (d_arr_13__27), .d_arr_13__26 (
               d_arr_13__26), .d_arr_13__25 (d_arr_13__25), .d_arr_13__24 (
               d_arr_13__24), .d_arr_13__23 (d_arr_13__23), .d_arr_13__22 (
               d_arr_13__22), .d_arr_13__21 (d_arr_13__21), .d_arr_13__20 (
               d_arr_13__20), .d_arr_13__19 (d_arr_13__19), .d_arr_13__18 (
               d_arr_13__18), .d_arr_13__17 (d_arr_13__17), .d_arr_13__16 (
               d_arr_13__16), .d_arr_13__15 (d_arr_13__15), .d_arr_13__14 (
               d_arr_13__14), .d_arr_13__13 (d_arr_13__13), .d_arr_13__12 (
               d_arr_13__12), .d_arr_13__11 (d_arr_13__11), .d_arr_13__10 (
               d_arr_13__10), .d_arr_13__9 (d_arr_13__9), .d_arr_13__8 (
               d_arr_13__8), .d_arr_13__7 (d_arr_13__7), .d_arr_13__6 (
               d_arr_13__6), .d_arr_13__5 (d_arr_13__5), .d_arr_13__4 (
               d_arr_13__4), .d_arr_13__3 (d_arr_13__3), .d_arr_13__2 (
               d_arr_13__2), .d_arr_13__1 (d_arr_13__1), .d_arr_13__0 (
               d_arr_13__0), .d_arr_14__31 (d_arr_14__31), .d_arr_14__30 (
               d_arr_14__30), .d_arr_14__29 (d_arr_14__29), .d_arr_14__28 (
               d_arr_14__28), .d_arr_14__27 (d_arr_14__27), .d_arr_14__26 (
               d_arr_14__26), .d_arr_14__25 (d_arr_14__25), .d_arr_14__24 (
               d_arr_14__24), .d_arr_14__23 (d_arr_14__23), .d_arr_14__22 (
               d_arr_14__22), .d_arr_14__21 (d_arr_14__21), .d_arr_14__20 (
               d_arr_14__20), .d_arr_14__19 (d_arr_14__19), .d_arr_14__18 (
               d_arr_14__18), .d_arr_14__17 (d_arr_14__17), .d_arr_14__16 (
               d_arr_14__16), .d_arr_14__15 (d_arr_14__15), .d_arr_14__14 (
               d_arr_14__14), .d_arr_14__13 (d_arr_14__13), .d_arr_14__12 (
               d_arr_14__12), .d_arr_14__11 (d_arr_14__11), .d_arr_14__10 (
               d_arr_14__10), .d_arr_14__9 (d_arr_14__9), .d_arr_14__8 (
               d_arr_14__8), .d_arr_14__7 (d_arr_14__7), .d_arr_14__6 (
               d_arr_14__6), .d_arr_14__5 (d_arr_14__5), .d_arr_14__4 (
               d_arr_14__4), .d_arr_14__3 (d_arr_14__3), .d_arr_14__2 (
               d_arr_14__2), .d_arr_14__1 (d_arr_14__1), .d_arr_14__0 (
               d_arr_14__0), .d_arr_15__31 (d_arr_15__31), .d_arr_15__30 (
               d_arr_15__30), .d_arr_15__29 (d_arr_15__29), .d_arr_15__28 (
               d_arr_15__28), .d_arr_15__27 (d_arr_15__27), .d_arr_15__26 (
               d_arr_15__26), .d_arr_15__25 (d_arr_15__25), .d_arr_15__24 (
               d_arr_15__24), .d_arr_15__23 (d_arr_15__23), .d_arr_15__22 (
               d_arr_15__22), .d_arr_15__21 (d_arr_15__21), .d_arr_15__20 (
               d_arr_15__20), .d_arr_15__19 (d_arr_15__19), .d_arr_15__18 (
               d_arr_15__18), .d_arr_15__17 (d_arr_15__17), .d_arr_15__16 (
               d_arr_15__16), .d_arr_15__15 (d_arr_15__15), .d_arr_15__14 (
               d_arr_15__14), .d_arr_15__13 (d_arr_15__13), .d_arr_15__12 (
               d_arr_15__12), .d_arr_15__11 (d_arr_15__11), .d_arr_15__10 (
               d_arr_15__10), .d_arr_15__9 (d_arr_15__9), .d_arr_15__8 (
               d_arr_15__8), .d_arr_15__7 (d_arr_15__7), .d_arr_15__6 (
               d_arr_15__6), .d_arr_15__5 (d_arr_15__5), .d_arr_15__4 (
               d_arr_15__4), .d_arr_15__3 (d_arr_15__3), .d_arr_15__2 (
               d_arr_15__2), .d_arr_15__1 (d_arr_15__1), .d_arr_15__0 (
               d_arr_15__0), .d_arr_16__31 (d_arr_16__31), .d_arr_16__30 (
               d_arr_16__30), .d_arr_16__29 (d_arr_16__29), .d_arr_16__28 (
               d_arr_16__28), .d_arr_16__27 (d_arr_16__27), .d_arr_16__26 (
               d_arr_16__26), .d_arr_16__25 (d_arr_16__25), .d_arr_16__24 (
               d_arr_16__24), .d_arr_16__23 (d_arr_16__23), .d_arr_16__22 (
               d_arr_16__22), .d_arr_16__21 (d_arr_16__21), .d_arr_16__20 (
               d_arr_16__20), .d_arr_16__19 (d_arr_16__19), .d_arr_16__18 (
               d_arr_16__18), .d_arr_16__17 (d_arr_16__17), .d_arr_16__16 (
               d_arr_16__16), .d_arr_16__15 (d_arr_16__15), .d_arr_16__14 (
               d_arr_16__14), .d_arr_16__13 (d_arr_16__13), .d_arr_16__12 (
               d_arr_16__12), .d_arr_16__11 (d_arr_16__11), .d_arr_16__10 (
               d_arr_16__10), .d_arr_16__9 (d_arr_16__9), .d_arr_16__8 (
               d_arr_16__8), .d_arr_16__7 (d_arr_16__7), .d_arr_16__6 (
               d_arr_16__6), .d_arr_16__5 (d_arr_16__5), .d_arr_16__4 (
               d_arr_16__4), .d_arr_16__3 (d_arr_16__3), .d_arr_16__2 (
               d_arr_16__2), .d_arr_16__1 (d_arr_16__1), .d_arr_16__0 (
               d_arr_16__0), .d_arr_17__31 (d_arr_17__31), .d_arr_17__30 (
               d_arr_17__30), .d_arr_17__29 (d_arr_17__29), .d_arr_17__28 (
               d_arr_17__28), .d_arr_17__27 (d_arr_17__27), .d_arr_17__26 (
               d_arr_17__26), .d_arr_17__25 (d_arr_17__25), .d_arr_17__24 (
               d_arr_17__24), .d_arr_17__23 (d_arr_17__23), .d_arr_17__22 (
               d_arr_17__22), .d_arr_17__21 (d_arr_17__21), .d_arr_17__20 (
               d_arr_17__20), .d_arr_17__19 (d_arr_17__19), .d_arr_17__18 (
               d_arr_17__18), .d_arr_17__17 (d_arr_17__17), .d_arr_17__16 (
               d_arr_17__16), .d_arr_17__15 (d_arr_17__15), .d_arr_17__14 (
               d_arr_17__14), .d_arr_17__13 (d_arr_17__13), .d_arr_17__12 (
               d_arr_17__12), .d_arr_17__11 (d_arr_17__11), .d_arr_17__10 (
               d_arr_17__10), .d_arr_17__9 (d_arr_17__9), .d_arr_17__8 (
               d_arr_17__8), .d_arr_17__7 (d_arr_17__7), .d_arr_17__6 (
               d_arr_17__6), .d_arr_17__5 (d_arr_17__5), .d_arr_17__4 (
               d_arr_17__4), .d_arr_17__3 (d_arr_17__3), .d_arr_17__2 (
               d_arr_17__2), .d_arr_17__1 (d_arr_17__1), .d_arr_17__0 (
               d_arr_17__0), .d_arr_18__31 (d_arr_18__31), .d_arr_18__30 (
               d_arr_18__30), .d_arr_18__29 (d_arr_18__29), .d_arr_18__28 (
               d_arr_18__28), .d_arr_18__27 (d_arr_18__27), .d_arr_18__26 (
               d_arr_18__26), .d_arr_18__25 (d_arr_18__25), .d_arr_18__24 (
               d_arr_18__24), .d_arr_18__23 (d_arr_18__23), .d_arr_18__22 (
               d_arr_18__22), .d_arr_18__21 (d_arr_18__21), .d_arr_18__20 (
               d_arr_18__20), .d_arr_18__19 (d_arr_18__19), .d_arr_18__18 (
               d_arr_18__18), .d_arr_18__17 (d_arr_18__17), .d_arr_18__16 (
               d_arr_18__16), .d_arr_18__15 (d_arr_18__15), .d_arr_18__14 (
               d_arr_18__14), .d_arr_18__13 (d_arr_18__13), .d_arr_18__12 (
               d_arr_18__12), .d_arr_18__11 (d_arr_18__11), .d_arr_18__10 (
               d_arr_18__10), .d_arr_18__9 (d_arr_18__9), .d_arr_18__8 (
               d_arr_18__8), .d_arr_18__7 (d_arr_18__7), .d_arr_18__6 (
               d_arr_18__6), .d_arr_18__5 (d_arr_18__5), .d_arr_18__4 (
               d_arr_18__4), .d_arr_18__3 (d_arr_18__3), .d_arr_18__2 (
               d_arr_18__2), .d_arr_18__1 (d_arr_18__1), .d_arr_18__0 (
               d_arr_18__0), .d_arr_19__31 (d_arr_19__31), .d_arr_19__30 (
               d_arr_19__30), .d_arr_19__29 (d_arr_19__29), .d_arr_19__28 (
               d_arr_19__28), .d_arr_19__27 (d_arr_19__27), .d_arr_19__26 (
               d_arr_19__26), .d_arr_19__25 (d_arr_19__25), .d_arr_19__24 (
               d_arr_19__24), .d_arr_19__23 (d_arr_19__23), .d_arr_19__22 (
               d_arr_19__22), .d_arr_19__21 (d_arr_19__21), .d_arr_19__20 (
               d_arr_19__20), .d_arr_19__19 (d_arr_19__19), .d_arr_19__18 (
               d_arr_19__18), .d_arr_19__17 (d_arr_19__17), .d_arr_19__16 (
               d_arr_19__16), .d_arr_19__15 (d_arr_19__15), .d_arr_19__14 (
               d_arr_19__14), .d_arr_19__13 (d_arr_19__13), .d_arr_19__12 (
               d_arr_19__12), .d_arr_19__11 (d_arr_19__11), .d_arr_19__10 (
               d_arr_19__10), .d_arr_19__9 (d_arr_19__9), .d_arr_19__8 (
               d_arr_19__8), .d_arr_19__7 (d_arr_19__7), .d_arr_19__6 (
               d_arr_19__6), .d_arr_19__5 (d_arr_19__5), .d_arr_19__4 (
               d_arr_19__4), .d_arr_19__3 (d_arr_19__3), .d_arr_19__2 (
               d_arr_19__2), .d_arr_19__1 (d_arr_19__1), .d_arr_19__0 (
               d_arr_19__0), .d_arr_20__31 (d_arr_20__31), .d_arr_20__30 (
               d_arr_20__30), .d_arr_20__29 (d_arr_20__29), .d_arr_20__28 (
               d_arr_20__28), .d_arr_20__27 (d_arr_20__27), .d_arr_20__26 (
               d_arr_20__26), .d_arr_20__25 (d_arr_20__25), .d_arr_20__24 (
               d_arr_20__24), .d_arr_20__23 (d_arr_20__23), .d_arr_20__22 (
               d_arr_20__22), .d_arr_20__21 (d_arr_20__21), .d_arr_20__20 (
               d_arr_20__20), .d_arr_20__19 (d_arr_20__19), .d_arr_20__18 (
               d_arr_20__18), .d_arr_20__17 (d_arr_20__17), .d_arr_20__16 (
               d_arr_20__16), .d_arr_20__15 (d_arr_20__15), .d_arr_20__14 (
               d_arr_20__14), .d_arr_20__13 (d_arr_20__13), .d_arr_20__12 (
               d_arr_20__12), .d_arr_20__11 (d_arr_20__11), .d_arr_20__10 (
               d_arr_20__10), .d_arr_20__9 (d_arr_20__9), .d_arr_20__8 (
               d_arr_20__8), .d_arr_20__7 (d_arr_20__7), .d_arr_20__6 (
               d_arr_20__6), .d_arr_20__5 (d_arr_20__5), .d_arr_20__4 (
               d_arr_20__4), .d_arr_20__3 (d_arr_20__3), .d_arr_20__2 (
               d_arr_20__2), .d_arr_20__1 (d_arr_20__1), .d_arr_20__0 (
               d_arr_20__0), .d_arr_21__31 (d_arr_21__31), .d_arr_21__30 (
               d_arr_21__30), .d_arr_21__29 (d_arr_21__29), .d_arr_21__28 (
               d_arr_21__28), .d_arr_21__27 (d_arr_21__27), .d_arr_21__26 (
               d_arr_21__26), .d_arr_21__25 (d_arr_21__25), .d_arr_21__24 (
               d_arr_21__24), .d_arr_21__23 (d_arr_21__23), .d_arr_21__22 (
               d_arr_21__22), .d_arr_21__21 (d_arr_21__21), .d_arr_21__20 (
               d_arr_21__20), .d_arr_21__19 (d_arr_21__19), .d_arr_21__18 (
               d_arr_21__18), .d_arr_21__17 (d_arr_21__17), .d_arr_21__16 (
               d_arr_21__16), .d_arr_21__15 (d_arr_21__15), .d_arr_21__14 (
               d_arr_21__14), .d_arr_21__13 (d_arr_21__13), .d_arr_21__12 (
               d_arr_21__12), .d_arr_21__11 (d_arr_21__11), .d_arr_21__10 (
               d_arr_21__10), .d_arr_21__9 (d_arr_21__9), .d_arr_21__8 (
               d_arr_21__8), .d_arr_21__7 (d_arr_21__7), .d_arr_21__6 (
               d_arr_21__6), .d_arr_21__5 (d_arr_21__5), .d_arr_21__4 (
               d_arr_21__4), .d_arr_21__3 (d_arr_21__3), .d_arr_21__2 (
               d_arr_21__2), .d_arr_21__1 (d_arr_21__1), .d_arr_21__0 (
               d_arr_21__0), .d_arr_22__31 (d_arr_22__31), .d_arr_22__30 (
               d_arr_22__30), .d_arr_22__29 (d_arr_22__29), .d_arr_22__28 (
               d_arr_22__28), .d_arr_22__27 (d_arr_22__27), .d_arr_22__26 (
               d_arr_22__26), .d_arr_22__25 (d_arr_22__25), .d_arr_22__24 (
               d_arr_22__24), .d_arr_22__23 (d_arr_22__23), .d_arr_22__22 (
               d_arr_22__22), .d_arr_22__21 (d_arr_22__21), .d_arr_22__20 (
               d_arr_22__20), .d_arr_22__19 (d_arr_22__19), .d_arr_22__18 (
               d_arr_22__18), .d_arr_22__17 (d_arr_22__17), .d_arr_22__16 (
               d_arr_22__16), .d_arr_22__15 (d_arr_22__15), .d_arr_22__14 (
               d_arr_22__14), .d_arr_22__13 (d_arr_22__13), .d_arr_22__12 (
               d_arr_22__12), .d_arr_22__11 (d_arr_22__11), .d_arr_22__10 (
               d_arr_22__10), .d_arr_22__9 (d_arr_22__9), .d_arr_22__8 (
               d_arr_22__8), .d_arr_22__7 (d_arr_22__7), .d_arr_22__6 (
               d_arr_22__6), .d_arr_22__5 (d_arr_22__5), .d_arr_22__4 (
               d_arr_22__4), .d_arr_22__3 (d_arr_22__3), .d_arr_22__2 (
               d_arr_22__2), .d_arr_22__1 (d_arr_22__1), .d_arr_22__0 (
               d_arr_22__0), .d_arr_23__31 (d_arr_23__31), .d_arr_23__30 (
               d_arr_23__30), .d_arr_23__29 (d_arr_23__29), .d_arr_23__28 (
               d_arr_23__28), .d_arr_23__27 (d_arr_23__27), .d_arr_23__26 (
               d_arr_23__26), .d_arr_23__25 (d_arr_23__25), .d_arr_23__24 (
               d_arr_23__24), .d_arr_23__23 (d_arr_23__23), .d_arr_23__22 (
               d_arr_23__22), .d_arr_23__21 (d_arr_23__21), .d_arr_23__20 (
               d_arr_23__20), .d_arr_23__19 (d_arr_23__19), .d_arr_23__18 (
               d_arr_23__18), .d_arr_23__17 (d_arr_23__17), .d_arr_23__16 (
               d_arr_23__16), .d_arr_23__15 (d_arr_23__15), .d_arr_23__14 (
               d_arr_23__14), .d_arr_23__13 (d_arr_23__13), .d_arr_23__12 (
               d_arr_23__12), .d_arr_23__11 (d_arr_23__11), .d_arr_23__10 (
               d_arr_23__10), .d_arr_23__9 (d_arr_23__9), .d_arr_23__8 (
               d_arr_23__8), .d_arr_23__7 (d_arr_23__7), .d_arr_23__6 (
               d_arr_23__6), .d_arr_23__5 (d_arr_23__5), .d_arr_23__4 (
               d_arr_23__4), .d_arr_23__3 (d_arr_23__3), .d_arr_23__2 (
               d_arr_23__2), .d_arr_23__1 (d_arr_23__1), .d_arr_23__0 (
               d_arr_23__0), .d_arr_24__31 (d_arr_24__31), .d_arr_24__30 (
               d_arr_24__30), .d_arr_24__29 (d_arr_24__29), .d_arr_24__28 (
               d_arr_24__28), .d_arr_24__27 (d_arr_24__27), .d_arr_24__26 (
               d_arr_24__26), .d_arr_24__25 (d_arr_24__25), .d_arr_24__24 (
               d_arr_24__24), .d_arr_24__23 (d_arr_24__23), .d_arr_24__22 (
               d_arr_24__22), .d_arr_24__21 (d_arr_24__21), .d_arr_24__20 (
               d_arr_24__20), .d_arr_24__19 (d_arr_24__19), .d_arr_24__18 (
               d_arr_24__18), .d_arr_24__17 (d_arr_24__17), .d_arr_24__16 (
               d_arr_24__16), .d_arr_24__15 (d_arr_24__15), .d_arr_24__14 (
               d_arr_24__14), .d_arr_24__13 (d_arr_24__13), .d_arr_24__12 (
               d_arr_24__12), .d_arr_24__11 (d_arr_24__11), .d_arr_24__10 (
               d_arr_24__10), .d_arr_24__9 (d_arr_24__9), .d_arr_24__8 (
               d_arr_24__8), .d_arr_24__7 (d_arr_24__7), .d_arr_24__6 (
               d_arr_24__6), .d_arr_24__5 (d_arr_24__5), .d_arr_24__4 (
               d_arr_24__4), .d_arr_24__3 (d_arr_24__3), .d_arr_24__2 (
               d_arr_24__2), .d_arr_24__1 (d_arr_24__1), .d_arr_24__0 (
               d_arr_24__0)) ;
    MuxLayer mux_layer_gen (.img_data_0__31 (GND0), .img_data_0__30 (GND0), .img_data_0__29 (
             GND0), .img_data_0__28 (GND0), .img_data_0__27 (GND0), .img_data_0__26 (
             GND0), .img_data_0__25 (GND0), .img_data_0__24 (GND0), .img_data_0__23 (
             GND0), .img_data_0__22 (GND0), .img_data_0__21 (GND0), .img_data_0__20 (
             GND0), .img_data_0__19 (GND0), .img_data_0__18 (GND0), .img_data_0__17 (
             GND0), .img_data_0__16 (GND0), .img_data_0__15 (GND0), .img_data_0__14 (
             GND0), .img_data_0__13 (GND0), .img_data_0__12 (GND0), .img_data_0__11 (
             GND0), .img_data_0__10 (GND0), .img_data_0__9 (GND0), .img_data_0__8 (
             GND0), .img_data_0__7 (GND0), .img_data_0__6 (GND0), .img_data_0__5 (
             GND0), .img_data_0__4 (GND0), .img_data_0__3 (GND0), .img_data_0__2 (
             GND0), .img_data_0__1 (GND0), .img_data_0__0 (GND0), .img_data_1__31 (
             img_data_1__15), .img_data_1__30 (GND0), .img_data_1__29 (GND0), .img_data_1__28 (
             GND0), .img_data_1__27 (GND0), .img_data_1__26 (GND0), .img_data_1__25 (
             GND0), .img_data_1__24 (GND0), .img_data_1__23 (GND0), .img_data_1__22 (
             GND0), .img_data_1__21 (GND0), .img_data_1__20 (GND0), .img_data_1__19 (
             GND0), .img_data_1__18 (GND0), .img_data_1__17 (GND0), .img_data_1__16 (
             GND0), .img_data_1__15 (GND0), .img_data_1__14 (nx19398), .img_data_1__13 (
             img_data_1__13), .img_data_1__12 (img_data_1__12), .img_data_1__11 (
             img_data_1__11), .img_data_1__10 (nx19402), .img_data_1__9 (
             img_data_1__9), .img_data_1__8 (img_data_1__8), .img_data_1__7 (
             img_data_1__7), .img_data_1__6 (img_data_1__6), .img_data_1__5 (
             img_data_1__5), .img_data_1__4 (img_data_1__4), .img_data_1__3 (
             img_data_1__3), .img_data_1__2 (img_data_1__2), .img_data_1__1 (
             img_data_1__1), .img_data_1__0 (img_data_1__0), .img_data_2__31 (
             img_data_2__15), .img_data_2__30 (GND0), .img_data_2__29 (GND0), .img_data_2__28 (
             GND0), .img_data_2__27 (GND0), .img_data_2__26 (GND0), .img_data_2__25 (
             GND0), .img_data_2__24 (GND0), .img_data_2__23 (GND0), .img_data_2__22 (
             GND0), .img_data_2__21 (GND0), .img_data_2__20 (GND0), .img_data_2__19 (
             GND0), .img_data_2__18 (GND0), .img_data_2__17 (GND0), .img_data_2__16 (
             GND0), .img_data_2__15 (GND0), .img_data_2__14 (nx19404), .img_data_2__13 (
             img_data_2__13), .img_data_2__12 (img_data_2__12), .img_data_2__11 (
             img_data_2__11), .img_data_2__10 (nx19408), .img_data_2__9 (
             img_data_2__9), .img_data_2__8 (img_data_2__8), .img_data_2__7 (
             img_data_2__7), .img_data_2__6 (img_data_2__6), .img_data_2__5 (
             img_data_2__5), .img_data_2__4 (img_data_2__4), .img_data_2__3 (
             img_data_2__3), .img_data_2__2 (img_data_2__2), .img_data_2__1 (
             img_data_2__1), .img_data_2__0 (img_data_2__0), .img_data_3__31 (
             img_data_3__15), .img_data_3__30 (GND0), .img_data_3__29 (GND0), .img_data_3__28 (
             GND0), .img_data_3__27 (GND0), .img_data_3__26 (GND0), .img_data_3__25 (
             GND0), .img_data_3__24 (GND0), .img_data_3__23 (GND0), .img_data_3__22 (
             GND0), .img_data_3__21 (GND0), .img_data_3__20 (GND0), .img_data_3__19 (
             GND0), .img_data_3__18 (GND0), .img_data_3__17 (GND0), .img_data_3__16 (
             GND0), .img_data_3__15 (GND0), .img_data_3__14 (img_data_3__14), .img_data_3__13 (
             img_data_3__13), .img_data_3__12 (img_data_3__12), .img_data_3__11 (
             img_data_3__11), .img_data_3__10 (img_data_3__10), .img_data_3__9 (
             img_data_3__9), .img_data_3__8 (img_data_3__8), .img_data_3__7 (
             img_data_3__7), .img_data_3__6 (img_data_3__6), .img_data_3__5 (
             img_data_3__5), .img_data_3__4 (img_data_3__4), .img_data_3__3 (
             img_data_3__3), .img_data_3__2 (img_data_3__2), .img_data_3__1 (
             img_data_3__1), .img_data_3__0 (img_data_3__0), .img_data_4__31 (
             img_data_4__15), .img_data_4__30 (GND0), .img_data_4__29 (GND0), .img_data_4__28 (
             GND0), .img_data_4__27 (GND0), .img_data_4__26 (GND0), .img_data_4__25 (
             GND0), .img_data_4__24 (GND0), .img_data_4__23 (GND0), .img_data_4__22 (
             GND0), .img_data_4__21 (GND0), .img_data_4__20 (GND0), .img_data_4__19 (
             GND0), .img_data_4__18 (GND0), .img_data_4__17 (GND0), .img_data_4__16 (
             GND0), .img_data_4__15 (GND0), .img_data_4__14 (img_data_4__14), .img_data_4__13 (
             img_data_4__13), .img_data_4__12 (img_data_4__12), .img_data_4__11 (
             img_data_4__11), .img_data_4__10 (img_data_4__10), .img_data_4__9 (
             img_data_4__9), .img_data_4__8 (img_data_4__8), .img_data_4__7 (
             img_data_4__7), .img_data_4__6 (img_data_4__6), .img_data_4__5 (
             img_data_4__5), .img_data_4__4 (img_data_4__4), .img_data_4__3 (
             img_data_4__3), .img_data_4__2 (img_data_4__2), .img_data_4__1 (
             img_data_4__1), .img_data_4__0 (img_data_4__0), .img_data_5__31 (
             GND0), .img_data_5__30 (GND0), .img_data_5__29 (GND0), .img_data_5__28 (
             GND0), .img_data_5__27 (GND0), .img_data_5__26 (GND0), .img_data_5__25 (
             GND0), .img_data_5__24 (GND0), .img_data_5__23 (GND0), .img_data_5__22 (
             GND0), .img_data_5__21 (GND0), .img_data_5__20 (GND0), .img_data_5__19 (
             GND0), .img_data_5__18 (GND0), .img_data_5__17 (GND0), .img_data_5__16 (
             GND0), .img_data_5__15 (GND0), .img_data_5__14 (GND0), .img_data_5__13 (
             GND0), .img_data_5__12 (GND0), .img_data_5__11 (GND0), .img_data_5__10 (
             GND0), .img_data_5__9 (GND0), .img_data_5__8 (GND0), .img_data_5__7 (
             GND0), .img_data_5__6 (GND0), .img_data_5__5 (GND0), .img_data_5__4 (
             GND0), .img_data_5__3 (GND0), .img_data_5__2 (GND0), .img_data_5__1 (
             GND0), .img_data_5__0 (GND0), .img_data_6__31 (img_data_6__15), .img_data_6__30 (
             GND0), .img_data_6__29 (GND0), .img_data_6__28 (GND0), .img_data_6__27 (
             GND0), .img_data_6__26 (GND0), .img_data_6__25 (GND0), .img_data_6__24 (
             GND0), .img_data_6__23 (GND0), .img_data_6__22 (GND0), .img_data_6__21 (
             GND0), .img_data_6__20 (GND0), .img_data_6__19 (GND0), .img_data_6__18 (
             GND0), .img_data_6__17 (GND0), .img_data_6__16 (GND0), .img_data_6__15 (
             GND0), .img_data_6__14 (nx19412), .img_data_6__13 (img_data_6__13)
             , .img_data_6__12 (img_data_6__12), .img_data_6__11 (img_data_6__11
             ), .img_data_6__10 (nx19416), .img_data_6__9 (img_data_6__9), .img_data_6__8 (
             img_data_6__8), .img_data_6__7 (img_data_6__7), .img_data_6__6 (
             img_data_6__6), .img_data_6__5 (img_data_6__5), .img_data_6__4 (
             img_data_6__4), .img_data_6__3 (img_data_6__3), .img_data_6__2 (
             img_data_6__2), .img_data_6__1 (img_data_6__1), .img_data_6__0 (
             img_data_6__0), .img_data_7__31 (nx16659), .img_data_7__30 (GND0), 
             .img_data_7__29 (GND0), .img_data_7__28 (GND0), .img_data_7__27 (
             GND0), .img_data_7__26 (GND0), .img_data_7__25 (GND0), .img_data_7__24 (
             GND0), .img_data_7__23 (GND0), .img_data_7__22 (GND0), .img_data_7__21 (
             GND0), .img_data_7__20 (GND0), .img_data_7__19 (GND0), .img_data_7__18 (
             GND0), .img_data_7__17 (GND0), .img_data_7__16 (GND0), .img_data_7__15 (
             GND0), .img_data_7__14 (nx19418), .img_data_7__13 (img_data_7__13)
             , .img_data_7__12 (img_data_7__12), .img_data_7__11 (img_data_7__11
             ), .img_data_7__10 (nx19422), .img_data_7__9 (img_data_7__9), .img_data_7__8 (
             img_data_7__8), .img_data_7__7 (img_data_7__7), .img_data_7__6 (
             img_data_7__6), .img_data_7__5 (img_data_7__5), .img_data_7__4 (
             img_data_7__4), .img_data_7__3 (img_data_7__3), .img_data_7__2 (
             img_data_7__2), .img_data_7__1 (img_data_7__1), .img_data_7__0 (
             img_data_7__0), .img_data_8__31 (img_data_8__15), .img_data_8__30 (
             GND0), .img_data_8__29 (GND0), .img_data_8__28 (GND0), .img_data_8__27 (
             GND0), .img_data_8__26 (GND0), .img_data_8__25 (GND0), .img_data_8__24 (
             GND0), .img_data_8__23 (GND0), .img_data_8__22 (GND0), .img_data_8__21 (
             GND0), .img_data_8__20 (GND0), .img_data_8__19 (GND0), .img_data_8__18 (
             GND0), .img_data_8__17 (GND0), .img_data_8__16 (GND0), .img_data_8__15 (
             GND0), .img_data_8__14 (img_data_8__14), .img_data_8__13 (
             img_data_8__13), .img_data_8__12 (img_data_8__12), .img_data_8__11 (
             img_data_8__11), .img_data_8__10 (img_data_8__10), .img_data_8__9 (
             img_data_8__9), .img_data_8__8 (img_data_8__8), .img_data_8__7 (
             img_data_8__7), .img_data_8__6 (img_data_8__6), .img_data_8__5 (
             img_data_8__5), .img_data_8__4 (img_data_8__4), .img_data_8__3 (
             img_data_8__3), .img_data_8__2 (img_data_8__2), .img_data_8__1 (
             img_data_8__1), .img_data_8__0 (img_data_8__0), .img_data_9__31 (
             img_data_9__15), .img_data_9__30 (GND0), .img_data_9__29 (GND0), .img_data_9__28 (
             GND0), .img_data_9__27 (GND0), .img_data_9__26 (GND0), .img_data_9__25 (
             GND0), .img_data_9__24 (GND0), .img_data_9__23 (GND0), .img_data_9__22 (
             GND0), .img_data_9__21 (GND0), .img_data_9__20 (GND0), .img_data_9__19 (
             GND0), .img_data_9__18 (GND0), .img_data_9__17 (GND0), .img_data_9__16 (
             GND0), .img_data_9__15 (GND0), .img_data_9__14 (img_data_9__14), .img_data_9__13 (
             img_data_9__13), .img_data_9__12 (img_data_9__12), .img_data_9__11 (
             img_data_9__11), .img_data_9__10 (img_data_9__10), .img_data_9__9 (
             img_data_9__9), .img_data_9__8 (img_data_9__8), .img_data_9__7 (
             img_data_9__7), .img_data_9__6 (img_data_9__6), .img_data_9__5 (
             img_data_9__5), .img_data_9__4 (img_data_9__4), .img_data_9__3 (
             img_data_9__3), .img_data_9__2 (img_data_9__2), .img_data_9__1 (
             img_data_9__1), .img_data_9__0 (img_data_9__0), .img_data_10__31 (
             GND0), .img_data_10__30 (GND0), .img_data_10__29 (GND0), .img_data_10__28 (
             GND0), .img_data_10__27 (GND0), .img_data_10__26 (GND0), .img_data_10__25 (
             GND0), .img_data_10__24 (GND0), .img_data_10__23 (GND0), .img_data_10__22 (
             GND0), .img_data_10__21 (GND0), .img_data_10__20 (GND0), .img_data_10__19 (
             GND0), .img_data_10__18 (GND0), .img_data_10__17 (GND0), .img_data_10__16 (
             GND0), .img_data_10__15 (GND0), .img_data_10__14 (GND0), .img_data_10__13 (
             GND0), .img_data_10__12 (GND0), .img_data_10__11 (GND0), .img_data_10__10 (
             GND0), .img_data_10__9 (GND0), .img_data_10__8 (GND0), .img_data_10__7 (
             GND0), .img_data_10__6 (GND0), .img_data_10__5 (GND0), .img_data_10__4 (
             GND0), .img_data_10__3 (GND0), .img_data_10__2 (GND0), .img_data_10__1 (
             GND0), .img_data_10__0 (GND0), .img_data_11__31 (nx16661), .img_data_11__30 (
             GND0), .img_data_11__29 (GND0), .img_data_11__28 (GND0), .img_data_11__27 (
             GND0), .img_data_11__26 (GND0), .img_data_11__25 (GND0), .img_data_11__24 (
             GND0), .img_data_11__23 (GND0), .img_data_11__22 (GND0), .img_data_11__21 (
             GND0), .img_data_11__20 (GND0), .img_data_11__19 (GND0), .img_data_11__18 (
             GND0), .img_data_11__17 (GND0), .img_data_11__16 (GND0), .img_data_11__15 (
             GND0), .img_data_11__14 (nx19426), .img_data_11__13 (
             img_data_11__13), .img_data_11__12 (img_data_11__12), .img_data_11__11 (
             img_data_11__11), .img_data_11__10 (nx19430), .img_data_11__9 (
             img_data_11__9), .img_data_11__8 (img_data_11__8), .img_data_11__7 (
             img_data_11__7), .img_data_11__6 (img_data_11__6), .img_data_11__5 (
             img_data_11__5), .img_data_11__4 (img_data_11__4), .img_data_11__3 (
             img_data_11__3), .img_data_11__2 (img_data_11__2), .img_data_11__1 (
             img_data_11__1), .img_data_11__0 (img_data_11__0), .img_data_12__31 (
             nx16663), .img_data_12__30 (GND0), .img_data_12__29 (GND0), .img_data_12__28 (
             GND0), .img_data_12__27 (GND0), .img_data_12__26 (GND0), .img_data_12__25 (
             GND0), .img_data_12__24 (GND0), .img_data_12__23 (GND0), .img_data_12__22 (
             GND0), .img_data_12__21 (GND0), .img_data_12__20 (GND0), .img_data_12__19 (
             GND0), .img_data_12__18 (GND0), .img_data_12__17 (GND0), .img_data_12__16 (
             GND0), .img_data_12__15 (GND0), .img_data_12__14 (nx19432), .img_data_12__13 (
             img_data_12__13), .img_data_12__12 (img_data_12__12), .img_data_12__11 (
             img_data_12__11), .img_data_12__10 (nx19436), .img_data_12__9 (
             img_data_12__9), .img_data_12__8 (img_data_12__8), .img_data_12__7 (
             img_data_12__7), .img_data_12__6 (img_data_12__6), .img_data_12__5 (
             img_data_12__5), .img_data_12__4 (img_data_12__4), .img_data_12__3 (
             img_data_12__3), .img_data_12__2 (img_data_12__2), .img_data_12__1 (
             img_data_12__1), .img_data_12__0 (img_data_12__0), .img_data_13__31 (
             img_data_13__15), .img_data_13__30 (GND0), .img_data_13__29 (GND0)
             , .img_data_13__28 (GND0), .img_data_13__27 (GND0), .img_data_13__26 (
             GND0), .img_data_13__25 (GND0), .img_data_13__24 (GND0), .img_data_13__23 (
             GND0), .img_data_13__22 (GND0), .img_data_13__21 (GND0), .img_data_13__20 (
             GND0), .img_data_13__19 (GND0), .img_data_13__18 (GND0), .img_data_13__17 (
             GND0), .img_data_13__16 (GND0), .img_data_13__15 (GND0), .img_data_13__14 (
             img_data_13__14), .img_data_13__13 (img_data_13__13), .img_data_13__12 (
             img_data_13__12), .img_data_13__11 (img_data_13__11), .img_data_13__10 (
             img_data_13__10), .img_data_13__9 (img_data_13__9), .img_data_13__8 (
             img_data_13__8), .img_data_13__7 (img_data_13__7), .img_data_13__6 (
             img_data_13__6), .img_data_13__5 (img_data_13__5), .img_data_13__4 (
             img_data_13__4), .img_data_13__3 (img_data_13__3), .img_data_13__2 (
             img_data_13__2), .img_data_13__1 (img_data_13__1), .img_data_13__0 (
             img_data_13__0), .img_data_14__31 (img_data_14__15), .img_data_14__30 (
             GND0), .img_data_14__29 (GND0), .img_data_14__28 (GND0), .img_data_14__27 (
             GND0), .img_data_14__26 (GND0), .img_data_14__25 (GND0), .img_data_14__24 (
             GND0), .img_data_14__23 (GND0), .img_data_14__22 (GND0), .img_data_14__21 (
             GND0), .img_data_14__20 (GND0), .img_data_14__19 (GND0), .img_data_14__18 (
             GND0), .img_data_14__17 (GND0), .img_data_14__16 (GND0), .img_data_14__15 (
             GND0), .img_data_14__14 (img_data_14__14), .img_data_14__13 (
             img_data_14__13), .img_data_14__12 (img_data_14__12), .img_data_14__11 (
             img_data_14__11), .img_data_14__10 (img_data_14__10), .img_data_14__9 (
             img_data_14__9), .img_data_14__8 (img_data_14__8), .img_data_14__7 (
             img_data_14__7), .img_data_14__6 (img_data_14__6), .img_data_14__5 (
             img_data_14__5), .img_data_14__4 (img_data_14__4), .img_data_14__3 (
             img_data_14__3), .img_data_14__2 (img_data_14__2), .img_data_14__1 (
             img_data_14__1), .img_data_14__0 (img_data_14__0), .img_data_15__31 (
             img_data_15__15), .img_data_15__30 (GND0), .img_data_15__29 (GND0)
             , .img_data_15__28 (GND0), .img_data_15__27 (GND0), .img_data_15__26 (
             GND0), .img_data_15__25 (GND0), .img_data_15__24 (GND0), .img_data_15__23 (
             GND0), .img_data_15__22 (GND0), .img_data_15__21 (GND0), .img_data_15__20 (
             GND0), .img_data_15__19 (GND0), .img_data_15__18 (GND0), .img_data_15__17 (
             GND0), .img_data_15__16 (GND0), .img_data_15__15 (GND0), .img_data_15__14 (
             img_data_15__14), .img_data_15__13 (img_data_15__13), .img_data_15__12 (
             img_data_15__12), .img_data_15__11 (img_data_15__11), .img_data_15__10 (
             img_data_15__10), .img_data_15__9 (img_data_15__9), .img_data_15__8 (
             img_data_15__8), .img_data_15__7 (img_data_15__7), .img_data_15__6 (
             img_data_15__6), .img_data_15__5 (img_data_15__5), .img_data_15__4 (
             img_data_15__4), .img_data_15__3 (img_data_15__3), .img_data_15__2 (
             img_data_15__2), .img_data_15__1 (img_data_15__1), .img_data_15__0 (
             img_data_15__0), .img_data_16__31 (img_data_16__15), .img_data_16__30 (
             GND0), .img_data_16__29 (GND0), .img_data_16__28 (GND0), .img_data_16__27 (
             GND0), .img_data_16__26 (GND0), .img_data_16__25 (GND0), .img_data_16__24 (
             GND0), .img_data_16__23 (GND0), .img_data_16__22 (GND0), .img_data_16__21 (
             GND0), .img_data_16__20 (GND0), .img_data_16__19 (GND0), .img_data_16__18 (
             GND0), .img_data_16__17 (GND0), .img_data_16__16 (GND0), .img_data_16__15 (
             GND0), .img_data_16__14 (img_data_16__14), .img_data_16__13 (
             img_data_16__13), .img_data_16__12 (img_data_16__12), .img_data_16__11 (
             img_data_16__11), .img_data_16__10 (img_data_16__10), .img_data_16__9 (
             img_data_16__9), .img_data_16__8 (img_data_16__8), .img_data_16__7 (
             img_data_16__7), .img_data_16__6 (img_data_16__6), .img_data_16__5 (
             img_data_16__5), .img_data_16__4 (img_data_16__4), .img_data_16__3 (
             img_data_16__3), .img_data_16__2 (img_data_16__2), .img_data_16__1 (
             img_data_16__1), .img_data_16__0 (img_data_16__0), .img_data_17__31 (
             img_data_17__15), .img_data_17__30 (GND0), .img_data_17__29 (GND0)
             , .img_data_17__28 (GND0), .img_data_17__27 (GND0), .img_data_17__26 (
             GND0), .img_data_17__25 (GND0), .img_data_17__24 (GND0), .img_data_17__23 (
             GND0), .img_data_17__22 (GND0), .img_data_17__21 (GND0), .img_data_17__20 (
             GND0), .img_data_17__19 (GND0), .img_data_17__18 (GND0), .img_data_17__17 (
             GND0), .img_data_17__16 (GND0), .img_data_17__15 (GND0), .img_data_17__14 (
             img_data_17__14), .img_data_17__13 (img_data_17__13), .img_data_17__12 (
             img_data_17__12), .img_data_17__11 (img_data_17__11), .img_data_17__10 (
             img_data_17__10), .img_data_17__9 (img_data_17__9), .img_data_17__8 (
             img_data_17__8), .img_data_17__7 (img_data_17__7), .img_data_17__6 (
             img_data_17__6), .img_data_17__5 (img_data_17__5), .img_data_17__4 (
             img_data_17__4), .img_data_17__3 (img_data_17__3), .img_data_17__2 (
             img_data_17__2), .img_data_17__1 (img_data_17__1), .img_data_17__0 (
             img_data_17__0), .img_data_18__31 (GND0), .img_data_18__30 (GND0), 
             .img_data_18__29 (GND0), .img_data_18__28 (GND0), .img_data_18__27 (
             GND0), .img_data_18__26 (GND0), .img_data_18__25 (GND0), .img_data_18__24 (
             GND0), .img_data_18__23 (GND0), .img_data_18__22 (GND0), .img_data_18__21 (
             GND0), .img_data_18__20 (GND0), .img_data_18__19 (GND0), .img_data_18__18 (
             GND0), .img_data_18__17 (GND0), .img_data_18__16 (GND0), .img_data_18__15 (
             GND0), .img_data_18__14 (GND0), .img_data_18__13 (GND0), .img_data_18__12 (
             GND0), .img_data_18__11 (GND0), .img_data_18__10 (GND0), .img_data_18__9 (
             GND0), .img_data_18__8 (GND0), .img_data_18__7 (GND0), .img_data_18__6 (
             GND0), .img_data_18__5 (GND0), .img_data_18__4 (GND0), .img_data_18__3 (
             GND0), .img_data_18__2 (GND0), .img_data_18__1 (GND0), .img_data_18__0 (
             GND0), .img_data_19__31 (GND0), .img_data_19__30 (GND0), .img_data_19__29 (
             GND0), .img_data_19__28 (GND0), .img_data_19__27 (GND0), .img_data_19__26 (
             GND0), .img_data_19__25 (GND0), .img_data_19__24 (GND0), .img_data_19__23 (
             GND0), .img_data_19__22 (GND0), .img_data_19__21 (GND0), .img_data_19__20 (
             GND0), .img_data_19__19 (GND0), .img_data_19__18 (GND0), .img_data_19__17 (
             GND0), .img_data_19__16 (GND0), .img_data_19__15 (GND0), .img_data_19__14 (
             GND0), .img_data_19__13 (GND0), .img_data_19__12 (GND0), .img_data_19__11 (
             GND0), .img_data_19__10 (GND0), .img_data_19__9 (GND0), .img_data_19__8 (
             GND0), .img_data_19__7 (GND0), .img_data_19__6 (GND0), .img_data_19__5 (
             GND0), .img_data_19__4 (GND0), .img_data_19__3 (GND0), .img_data_19__2 (
             GND0), .img_data_19__1 (GND0), .img_data_19__0 (GND0), .img_data_20__31 (
             GND0), .img_data_20__30 (GND0), .img_data_20__29 (GND0), .img_data_20__28 (
             GND0), .img_data_20__27 (GND0), .img_data_20__26 (GND0), .img_data_20__25 (
             GND0), .img_data_20__24 (GND0), .img_data_20__23 (GND0), .img_data_20__22 (
             GND0), .img_data_20__21 (GND0), .img_data_20__20 (GND0), .img_data_20__19 (
             GND0), .img_data_20__18 (GND0), .img_data_20__17 (GND0), .img_data_20__16 (
             GND0), .img_data_20__15 (GND0), .img_data_20__14 (GND0), .img_data_20__13 (
             GND0), .img_data_20__12 (GND0), .img_data_20__11 (GND0), .img_data_20__10 (
             GND0), .img_data_20__9 (GND0), .img_data_20__8 (GND0), .img_data_20__7 (
             GND0), .img_data_20__6 (GND0), .img_data_20__5 (GND0), .img_data_20__4 (
             GND0), .img_data_20__3 (GND0), .img_data_20__2 (GND0), .img_data_20__1 (
             GND0), .img_data_20__0 (GND0), .img_data_21__31 (GND0), .img_data_21__30 (
             GND0), .img_data_21__29 (GND0), .img_data_21__28 (GND0), .img_data_21__27 (
             GND0), .img_data_21__26 (GND0), .img_data_21__25 (GND0), .img_data_21__24 (
             GND0), .img_data_21__23 (GND0), .img_data_21__22 (GND0), .img_data_21__21 (
             GND0), .img_data_21__20 (GND0), .img_data_21__19 (GND0), .img_data_21__18 (
             GND0), .img_data_21__17 (GND0), .img_data_21__16 (GND0), .img_data_21__15 (
             GND0), .img_data_21__14 (GND0), .img_data_21__13 (GND0), .img_data_21__12 (
             GND0), .img_data_21__11 (GND0), .img_data_21__10 (GND0), .img_data_21__9 (
             GND0), .img_data_21__8 (GND0), .img_data_21__7 (GND0), .img_data_21__6 (
             GND0), .img_data_21__5 (GND0), .img_data_21__4 (GND0), .img_data_21__3 (
             GND0), .img_data_21__2 (GND0), .img_data_21__1 (GND0), .img_data_21__0 (
             GND0), .img_data_22__31 (GND0), .img_data_22__30 (GND0), .img_data_22__29 (
             GND0), .img_data_22__28 (GND0), .img_data_22__27 (GND0), .img_data_22__26 (
             GND0), .img_data_22__25 (GND0), .img_data_22__24 (GND0), .img_data_22__23 (
             GND0), .img_data_22__22 (GND0), .img_data_22__21 (GND0), .img_data_22__20 (
             GND0), .img_data_22__19 (GND0), .img_data_22__18 (GND0), .img_data_22__17 (
             GND0), .img_data_22__16 (GND0), .img_data_22__15 (GND0), .img_data_22__14 (
             GND0), .img_data_22__13 (GND0), .img_data_22__12 (GND0), .img_data_22__11 (
             GND0), .img_data_22__10 (GND0), .img_data_22__9 (GND0), .img_data_22__8 (
             GND0), .img_data_22__7 (GND0), .img_data_22__6 (GND0), .img_data_22__5 (
             GND0), .img_data_22__4 (GND0), .img_data_22__3 (GND0), .img_data_22__2 (
             GND0), .img_data_22__1 (GND0), .img_data_22__0 (GND0), .img_data_23__31 (
             GND0), .img_data_23__30 (GND0), .img_data_23__29 (GND0), .img_data_23__28 (
             GND0), .img_data_23__27 (GND0), .img_data_23__26 (GND0), .img_data_23__25 (
             GND0), .img_data_23__24 (GND0), .img_data_23__23 (GND0), .img_data_23__22 (
             GND0), .img_data_23__21 (GND0), .img_data_23__20 (GND0), .img_data_23__19 (
             GND0), .img_data_23__18 (GND0), .img_data_23__17 (GND0), .img_data_23__16 (
             GND0), .img_data_23__15 (GND0), .img_data_23__14 (GND0), .img_data_23__13 (
             GND0), .img_data_23__12 (GND0), .img_data_23__11 (GND0), .img_data_23__10 (
             GND0), .img_data_23__9 (GND0), .img_data_23__8 (GND0), .img_data_23__7 (
             GND0), .img_data_23__6 (GND0), .img_data_23__5 (GND0), .img_data_23__4 (
             GND0), .img_data_23__3 (GND0), .img_data_23__2 (GND0), .img_data_23__1 (
             GND0), .img_data_23__0 (GND0), .img_data_24__31 (GND0), .img_data_24__30 (
             GND0), .img_data_24__29 (GND0), .img_data_24__28 (GND0), .img_data_24__27 (
             GND0), .img_data_24__26 (GND0), .img_data_24__25 (GND0), .img_data_24__24 (
             GND0), .img_data_24__23 (GND0), .img_data_24__22 (GND0), .img_data_24__21 (
             GND0), .img_data_24__20 (GND0), .img_data_24__19 (GND0), .img_data_24__18 (
             GND0), .img_data_24__17 (GND0), .img_data_24__16 (GND0), .img_data_24__15 (
             GND0), .img_data_24__14 (GND0), .img_data_24__13 (GND0), .img_data_24__12 (
             GND0), .img_data_24__11 (GND0), .img_data_24__10 (GND0), .img_data_24__9 (
             GND0), .img_data_24__8 (GND0), .img_data_24__7 (GND0), .img_data_24__6 (
             GND0), .img_data_24__5 (GND0), .img_data_24__4 (GND0), .img_data_24__3 (
             GND0), .img_data_24__2 (GND0), .img_data_24__1 (GND0), .img_data_24__0 (
             GND0), .filter_data_0__31 (filter_data_0__15), .filter_data_0__30 (
             GND0), .filter_data_0__29 (GND0), .filter_data_0__28 (GND0), .filter_data_0__27 (
             GND0), .filter_data_0__26 (GND0), .filter_data_0__25 (GND0), .filter_data_0__24 (
             GND0), .filter_data_0__23 (GND0), .filter_data_0__22 (GND0), .filter_data_0__21 (
             GND0), .filter_data_0__20 (GND0), .filter_data_0__19 (GND0), .filter_data_0__18 (
             GND0), .filter_data_0__17 (GND0), .filter_data_0__16 (GND0), .filter_data_0__15 (
             GND0), .filter_data_0__14 (filter_data_0__14), .filter_data_0__13 (
             filter_data_0__13), .filter_data_0__12 (filter_data_0__12), .filter_data_0__11 (
             filter_data_0__11), .filter_data_0__10 (filter_data_0__10), .filter_data_0__9 (
             filter_data_0__9), .filter_data_0__8 (filter_data_0__8), .filter_data_0__7 (
             filter_data_0__7), .filter_data_0__6 (filter_data_0__6), .filter_data_0__5 (
             filter_data_0__5), .filter_data_0__4 (filter_data_0__4), .filter_data_0__3 (
             filter_data_0__3), .filter_data_0__2 (filter_data_0__2), .filter_data_0__1 (
             filter_data_0__1), .filter_data_0__0 (filter_data_0__0), .filter_data_1__31 (
             filter_data_1__15), .filter_data_1__30 (GND0), .filter_data_1__29 (
             GND0), .filter_data_1__28 (GND0), .filter_data_1__27 (GND0), .filter_data_1__26 (
             GND0), .filter_data_1__25 (GND0), .filter_data_1__24 (GND0), .filter_data_1__23 (
             GND0), .filter_data_1__22 (GND0), .filter_data_1__21 (GND0), .filter_data_1__20 (
             GND0), .filter_data_1__19 (GND0), .filter_data_1__18 (GND0), .filter_data_1__17 (
             GND0), .filter_data_1__16 (GND0), .filter_data_1__15 (GND0), .filter_data_1__14 (
             filter_data_1__14), .filter_data_1__13 (filter_data_1__13), .filter_data_1__12 (
             filter_data_1__12), .filter_data_1__11 (filter_data_1__11), .filter_data_1__10 (
             filter_data_1__10), .filter_data_1__9 (filter_data_1__9), .filter_data_1__8 (
             filter_data_1__8), .filter_data_1__7 (filter_data_1__7), .filter_data_1__6 (
             filter_data_1__6), .filter_data_1__5 (filter_data_1__5), .filter_data_1__4 (
             filter_data_1__4), .filter_data_1__3 (filter_data_1__3), .filter_data_1__2 (
             filter_data_1__2), .filter_data_1__1 (filter_data_1__1), .filter_data_1__0 (
             filter_data_1__0), .filter_data_2__31 (filter_data_2__15), .filter_data_2__30 (
             GND0), .filter_data_2__29 (GND0), .filter_data_2__28 (GND0), .filter_data_2__27 (
             GND0), .filter_data_2__26 (GND0), .filter_data_2__25 (GND0), .filter_data_2__24 (
             GND0), .filter_data_2__23 (GND0), .filter_data_2__22 (GND0), .filter_data_2__21 (
             GND0), .filter_data_2__20 (GND0), .filter_data_2__19 (GND0), .filter_data_2__18 (
             GND0), .filter_data_2__17 (GND0), .filter_data_2__16 (GND0), .filter_data_2__15 (
             GND0), .filter_data_2__14 (filter_data_2__14), .filter_data_2__13 (
             filter_data_2__13), .filter_data_2__12 (filter_data_2__12), .filter_data_2__11 (
             filter_data_2__11), .filter_data_2__10 (filter_data_2__10), .filter_data_2__9 (
             filter_data_2__9), .filter_data_2__8 (filter_data_2__8), .filter_data_2__7 (
             filter_data_2__7), .filter_data_2__6 (filter_data_2__6), .filter_data_2__5 (
             filter_data_2__5), .filter_data_2__4 (filter_data_2__4), .filter_data_2__3 (
             filter_data_2__3), .filter_data_2__2 (filter_data_2__2), .filter_data_2__1 (
             filter_data_2__1), .filter_data_2__0 (filter_data_2__0), .filter_data_3__31 (
             filter_data_3__15), .filter_data_3__30 (GND0), .filter_data_3__29 (
             GND0), .filter_data_3__28 (GND0), .filter_data_3__27 (GND0), .filter_data_3__26 (
             GND0), .filter_data_3__25 (GND0), .filter_data_3__24 (GND0), .filter_data_3__23 (
             GND0), .filter_data_3__22 (GND0), .filter_data_3__21 (GND0), .filter_data_3__20 (
             GND0), .filter_data_3__19 (GND0), .filter_data_3__18 (GND0), .filter_data_3__17 (
             GND0), .filter_data_3__16 (GND0), .filter_data_3__15 (GND0), .filter_data_3__14 (
             filter_data_3__14), .filter_data_3__13 (filter_data_3__13), .filter_data_3__12 (
             filter_data_3__12), .filter_data_3__11 (filter_data_3__11), .filter_data_3__10 (
             filter_data_3__10), .filter_data_3__9 (filter_data_3__9), .filter_data_3__8 (
             filter_data_3__8), .filter_data_3__7 (filter_data_3__7), .filter_data_3__6 (
             filter_data_3__6), .filter_data_3__5 (filter_data_3__5), .filter_data_3__4 (
             filter_data_3__4), .filter_data_3__3 (filter_data_3__3), .filter_data_3__2 (
             filter_data_3__2), .filter_data_3__1 (filter_data_3__1), .filter_data_3__0 (
             filter_data_3__0), .filter_data_4__31 (filter_data_4__15), .filter_data_4__30 (
             GND0), .filter_data_4__29 (GND0), .filter_data_4__28 (GND0), .filter_data_4__27 (
             GND0), .filter_data_4__26 (GND0), .filter_data_4__25 (GND0), .filter_data_4__24 (
             GND0), .filter_data_4__23 (GND0), .filter_data_4__22 (GND0), .filter_data_4__21 (
             GND0), .filter_data_4__20 (GND0), .filter_data_4__19 (GND0), .filter_data_4__18 (
             GND0), .filter_data_4__17 (GND0), .filter_data_4__16 (GND0), .filter_data_4__15 (
             GND0), .filter_data_4__14 (filter_data_4__14), .filter_data_4__13 (
             filter_data_4__13), .filter_data_4__12 (filter_data_4__12), .filter_data_4__11 (
             filter_data_4__11), .filter_data_4__10 (filter_data_4__10), .filter_data_4__9 (
             filter_data_4__9), .filter_data_4__8 (filter_data_4__8), .filter_data_4__7 (
             filter_data_4__7), .filter_data_4__6 (filter_data_4__6), .filter_data_4__5 (
             filter_data_4__5), .filter_data_4__4 (filter_data_4__4), .filter_data_4__3 (
             filter_data_4__3), .filter_data_4__2 (filter_data_4__2), .filter_data_4__1 (
             filter_data_4__1), .filter_data_4__0 (filter_data_4__0), .filter_data_5__31 (
             filter_data_5__15), .filter_data_5__30 (GND0), .filter_data_5__29 (
             GND0), .filter_data_5__28 (GND0), .filter_data_5__27 (GND0), .filter_data_5__26 (
             GND0), .filter_data_5__25 (GND0), .filter_data_5__24 (GND0), .filter_data_5__23 (
             GND0), .filter_data_5__22 (GND0), .filter_data_5__21 (GND0), .filter_data_5__20 (
             GND0), .filter_data_5__19 (GND0), .filter_data_5__18 (GND0), .filter_data_5__17 (
             GND0), .filter_data_5__16 (GND0), .filter_data_5__15 (GND0), .filter_data_5__14 (
             filter_data_5__14), .filter_data_5__13 (filter_data_5__13), .filter_data_5__12 (
             filter_data_5__12), .filter_data_5__11 (filter_data_5__11), .filter_data_5__10 (
             filter_data_5__10), .filter_data_5__9 (filter_data_5__9), .filter_data_5__8 (
             filter_data_5__8), .filter_data_5__7 (filter_data_5__7), .filter_data_5__6 (
             filter_data_5__6), .filter_data_5__5 (filter_data_5__5), .filter_data_5__4 (
             filter_data_5__4), .filter_data_5__3 (filter_data_5__3), .filter_data_5__2 (
             filter_data_5__2), .filter_data_5__1 (filter_data_5__1), .filter_data_5__0 (
             filter_data_5__0), .filter_data_6__31 (filter_data_6__15), .filter_data_6__30 (
             GND0), .filter_data_6__29 (GND0), .filter_data_6__28 (GND0), .filter_data_6__27 (
             GND0), .filter_data_6__26 (GND0), .filter_data_6__25 (GND0), .filter_data_6__24 (
             GND0), .filter_data_6__23 (GND0), .filter_data_6__22 (GND0), .filter_data_6__21 (
             GND0), .filter_data_6__20 (GND0), .filter_data_6__19 (GND0), .filter_data_6__18 (
             GND0), .filter_data_6__17 (GND0), .filter_data_6__16 (GND0), .filter_data_6__15 (
             GND0), .filter_data_6__14 (filter_data_6__14), .filter_data_6__13 (
             filter_data_6__13), .filter_data_6__12 (filter_data_6__12), .filter_data_6__11 (
             filter_data_6__11), .filter_data_6__10 (filter_data_6__10), .filter_data_6__9 (
             filter_data_6__9), .filter_data_6__8 (filter_data_6__8), .filter_data_6__7 (
             filter_data_6__7), .filter_data_6__6 (filter_data_6__6), .filter_data_6__5 (
             filter_data_6__5), .filter_data_6__4 (filter_data_6__4), .filter_data_6__3 (
             filter_data_6__3), .filter_data_6__2 (filter_data_6__2), .filter_data_6__1 (
             filter_data_6__1), .filter_data_6__0 (filter_data_6__0), .filter_data_7__31 (
             filter_data_7__15), .filter_data_7__30 (GND0), .filter_data_7__29 (
             GND0), .filter_data_7__28 (GND0), .filter_data_7__27 (GND0), .filter_data_7__26 (
             GND0), .filter_data_7__25 (GND0), .filter_data_7__24 (GND0), .filter_data_7__23 (
             GND0), .filter_data_7__22 (GND0), .filter_data_7__21 (GND0), .filter_data_7__20 (
             GND0), .filter_data_7__19 (GND0), .filter_data_7__18 (GND0), .filter_data_7__17 (
             GND0), .filter_data_7__16 (GND0), .filter_data_7__15 (GND0), .filter_data_7__14 (
             filter_data_7__14), .filter_data_7__13 (filter_data_7__13), .filter_data_7__12 (
             filter_data_7__12), .filter_data_7__11 (filter_data_7__11), .filter_data_7__10 (
             filter_data_7__10), .filter_data_7__9 (filter_data_7__9), .filter_data_7__8 (
             filter_data_7__8), .filter_data_7__7 (filter_data_7__7), .filter_data_7__6 (
             filter_data_7__6), .filter_data_7__5 (filter_data_7__5), .filter_data_7__4 (
             filter_data_7__4), .filter_data_7__3 (filter_data_7__3), .filter_data_7__2 (
             filter_data_7__2), .filter_data_7__1 (filter_data_7__1), .filter_data_7__0 (
             filter_data_7__0), .filter_data_8__31 (filter_data_8__15), .filter_data_8__30 (
             GND0), .filter_data_8__29 (GND0), .filter_data_8__28 (GND0), .filter_data_8__27 (
             GND0), .filter_data_8__26 (GND0), .filter_data_8__25 (GND0), .filter_data_8__24 (
             GND0), .filter_data_8__23 (GND0), .filter_data_8__22 (GND0), .filter_data_8__21 (
             GND0), .filter_data_8__20 (GND0), .filter_data_8__19 (GND0), .filter_data_8__18 (
             GND0), .filter_data_8__17 (GND0), .filter_data_8__16 (GND0), .filter_data_8__15 (
             GND0), .filter_data_8__14 (filter_data_8__14), .filter_data_8__13 (
             filter_data_8__13), .filter_data_8__12 (filter_data_8__12), .filter_data_8__11 (
             filter_data_8__11), .filter_data_8__10 (filter_data_8__10), .filter_data_8__9 (
             filter_data_8__9), .filter_data_8__8 (filter_data_8__8), .filter_data_8__7 (
             filter_data_8__7), .filter_data_8__6 (filter_data_8__6), .filter_data_8__5 (
             filter_data_8__5), .filter_data_8__4 (filter_data_8__4), .filter_data_8__3 (
             filter_data_8__3), .filter_data_8__2 (filter_data_8__2), .filter_data_8__1 (
             filter_data_8__1), .filter_data_8__0 (filter_data_8__0), .filter_data_9__31 (
             filter_data_9__15), .filter_data_9__30 (GND0), .filter_data_9__29 (
             GND0), .filter_data_9__28 (GND0), .filter_data_9__27 (GND0), .filter_data_9__26 (
             GND0), .filter_data_9__25 (GND0), .filter_data_9__24 (GND0), .filter_data_9__23 (
             GND0), .filter_data_9__22 (GND0), .filter_data_9__21 (GND0), .filter_data_9__20 (
             GND0), .filter_data_9__19 (GND0), .filter_data_9__18 (GND0), .filter_data_9__17 (
             GND0), .filter_data_9__16 (GND0), .filter_data_9__15 (GND0), .filter_data_9__14 (
             filter_data_9__14), .filter_data_9__13 (filter_data_9__13), .filter_data_9__12 (
             filter_data_9__12), .filter_data_9__11 (filter_data_9__11), .filter_data_9__10 (
             filter_data_9__10), .filter_data_9__9 (filter_data_9__9), .filter_data_9__8 (
             filter_data_9__8), .filter_data_9__7 (filter_data_9__7), .filter_data_9__6 (
             filter_data_9__6), .filter_data_9__5 (filter_data_9__5), .filter_data_9__4 (
             filter_data_9__4), .filter_data_9__3 (filter_data_9__3), .filter_data_9__2 (
             filter_data_9__2), .filter_data_9__1 (filter_data_9__1), .filter_data_9__0 (
             filter_data_9__0), .filter_data_10__31 (filter_data_10__15), .filter_data_10__30 (
             GND0), .filter_data_10__29 (GND0), .filter_data_10__28 (GND0), .filter_data_10__27 (
             GND0), .filter_data_10__26 (GND0), .filter_data_10__25 (GND0), .filter_data_10__24 (
             GND0), .filter_data_10__23 (GND0), .filter_data_10__22 (GND0), .filter_data_10__21 (
             GND0), .filter_data_10__20 (GND0), .filter_data_10__19 (GND0), .filter_data_10__18 (
             GND0), .filter_data_10__17 (GND0), .filter_data_10__16 (GND0), .filter_data_10__15 (
             GND0), .filter_data_10__14 (filter_data_10__14), .filter_data_10__13 (
             filter_data_10__13), .filter_data_10__12 (filter_data_10__12), .filter_data_10__11 (
             filter_data_10__11), .filter_data_10__10 (filter_data_10__10), .filter_data_10__9 (
             filter_data_10__9), .filter_data_10__8 (filter_data_10__8), .filter_data_10__7 (
             filter_data_10__7), .filter_data_10__6 (filter_data_10__6), .filter_data_10__5 (
             filter_data_10__5), .filter_data_10__4 (filter_data_10__4), .filter_data_10__3 (
             filter_data_10__3), .filter_data_10__2 (filter_data_10__2), .filter_data_10__1 (
             filter_data_10__1), .filter_data_10__0 (filter_data_10__0), .filter_data_11__31 (
             filter_data_11__15), .filter_data_11__30 (GND0), .filter_data_11__29 (
             GND0), .filter_data_11__28 (GND0), .filter_data_11__27 (GND0), .filter_data_11__26 (
             GND0), .filter_data_11__25 (GND0), .filter_data_11__24 (GND0), .filter_data_11__23 (
             GND0), .filter_data_11__22 (GND0), .filter_data_11__21 (GND0), .filter_data_11__20 (
             GND0), .filter_data_11__19 (GND0), .filter_data_11__18 (GND0), .filter_data_11__17 (
             GND0), .filter_data_11__16 (GND0), .filter_data_11__15 (GND0), .filter_data_11__14 (
             filter_data_11__14), .filter_data_11__13 (filter_data_11__13), .filter_data_11__12 (
             filter_data_11__12), .filter_data_11__11 (filter_data_11__11), .filter_data_11__10 (
             filter_data_11__10), .filter_data_11__9 (filter_data_11__9), .filter_data_11__8 (
             filter_data_11__8), .filter_data_11__7 (filter_data_11__7), .filter_data_11__6 (
             filter_data_11__6), .filter_data_11__5 (filter_data_11__5), .filter_data_11__4 (
             filter_data_11__4), .filter_data_11__3 (filter_data_11__3), .filter_data_11__2 (
             filter_data_11__2), .filter_data_11__1 (filter_data_11__1), .filter_data_11__0 (
             filter_data_11__0), .filter_data_12__31 (filter_data_12__15), .filter_data_12__30 (
             GND0), .filter_data_12__29 (GND0), .filter_data_12__28 (GND0), .filter_data_12__27 (
             GND0), .filter_data_12__26 (GND0), .filter_data_12__25 (GND0), .filter_data_12__24 (
             GND0), .filter_data_12__23 (GND0), .filter_data_12__22 (GND0), .filter_data_12__21 (
             GND0), .filter_data_12__20 (GND0), .filter_data_12__19 (GND0), .filter_data_12__18 (
             GND0), .filter_data_12__17 (GND0), .filter_data_12__16 (GND0), .filter_data_12__15 (
             GND0), .filter_data_12__14 (filter_data_12__14), .filter_data_12__13 (
             filter_data_12__13), .filter_data_12__12 (filter_data_12__12), .filter_data_12__11 (
             filter_data_12__11), .filter_data_12__10 (filter_data_12__10), .filter_data_12__9 (
             filter_data_12__9), .filter_data_12__8 (filter_data_12__8), .filter_data_12__7 (
             filter_data_12__7), .filter_data_12__6 (filter_data_12__6), .filter_data_12__5 (
             filter_data_12__5), .filter_data_12__4 (filter_data_12__4), .filter_data_12__3 (
             filter_data_12__3), .filter_data_12__2 (filter_data_12__2), .filter_data_12__1 (
             filter_data_12__1), .filter_data_12__0 (filter_data_12__0), .filter_data_13__31 (
             filter_data_13__15), .filter_data_13__30 (GND0), .filter_data_13__29 (
             GND0), .filter_data_13__28 (GND0), .filter_data_13__27 (GND0), .filter_data_13__26 (
             GND0), .filter_data_13__25 (GND0), .filter_data_13__24 (GND0), .filter_data_13__23 (
             GND0), .filter_data_13__22 (GND0), .filter_data_13__21 (GND0), .filter_data_13__20 (
             GND0), .filter_data_13__19 (GND0), .filter_data_13__18 (GND0), .filter_data_13__17 (
             GND0), .filter_data_13__16 (GND0), .filter_data_13__15 (GND0), .filter_data_13__14 (
             filter_data_13__14), .filter_data_13__13 (filter_data_13__13), .filter_data_13__12 (
             filter_data_13__12), .filter_data_13__11 (filter_data_13__11), .filter_data_13__10 (
             filter_data_13__10), .filter_data_13__9 (filter_data_13__9), .filter_data_13__8 (
             filter_data_13__8), .filter_data_13__7 (filter_data_13__7), .filter_data_13__6 (
             filter_data_13__6), .filter_data_13__5 (filter_data_13__5), .filter_data_13__4 (
             filter_data_13__4), .filter_data_13__3 (filter_data_13__3), .filter_data_13__2 (
             filter_data_13__2), .filter_data_13__1 (filter_data_13__1), .filter_data_13__0 (
             filter_data_13__0), .filter_data_14__31 (filter_data_14__15), .filter_data_14__30 (
             GND0), .filter_data_14__29 (GND0), .filter_data_14__28 (GND0), .filter_data_14__27 (
             GND0), .filter_data_14__26 (GND0), .filter_data_14__25 (GND0), .filter_data_14__24 (
             GND0), .filter_data_14__23 (GND0), .filter_data_14__22 (GND0), .filter_data_14__21 (
             GND0), .filter_data_14__20 (GND0), .filter_data_14__19 (GND0), .filter_data_14__18 (
             GND0), .filter_data_14__17 (GND0), .filter_data_14__16 (GND0), .filter_data_14__15 (
             GND0), .filter_data_14__14 (filter_data_14__14), .filter_data_14__13 (
             filter_data_14__13), .filter_data_14__12 (filter_data_14__12), .filter_data_14__11 (
             filter_data_14__11), .filter_data_14__10 (filter_data_14__10), .filter_data_14__9 (
             filter_data_14__9), .filter_data_14__8 (filter_data_14__8), .filter_data_14__7 (
             filter_data_14__7), .filter_data_14__6 (filter_data_14__6), .filter_data_14__5 (
             filter_data_14__5), .filter_data_14__4 (filter_data_14__4), .filter_data_14__3 (
             filter_data_14__3), .filter_data_14__2 (filter_data_14__2), .filter_data_14__1 (
             filter_data_14__1), .filter_data_14__0 (filter_data_14__0), .filter_data_15__31 (
             filter_data_15__15), .filter_data_15__30 (GND0), .filter_data_15__29 (
             GND0), .filter_data_15__28 (GND0), .filter_data_15__27 (GND0), .filter_data_15__26 (
             GND0), .filter_data_15__25 (GND0), .filter_data_15__24 (GND0), .filter_data_15__23 (
             GND0), .filter_data_15__22 (GND0), .filter_data_15__21 (GND0), .filter_data_15__20 (
             GND0), .filter_data_15__19 (GND0), .filter_data_15__18 (GND0), .filter_data_15__17 (
             GND0), .filter_data_15__16 (GND0), .filter_data_15__15 (GND0), .filter_data_15__14 (
             filter_data_15__14), .filter_data_15__13 (filter_data_15__13), .filter_data_15__12 (
             filter_data_15__12), .filter_data_15__11 (filter_data_15__11), .filter_data_15__10 (
             filter_data_15__10), .filter_data_15__9 (filter_data_15__9), .filter_data_15__8 (
             filter_data_15__8), .filter_data_15__7 (filter_data_15__7), .filter_data_15__6 (
             filter_data_15__6), .filter_data_15__5 (filter_data_15__5), .filter_data_15__4 (
             filter_data_15__4), .filter_data_15__3 (filter_data_15__3), .filter_data_15__2 (
             filter_data_15__2), .filter_data_15__1 (filter_data_15__1), .filter_data_15__0 (
             filter_data_15__0), .filter_data_16__31 (filter_data_16__15), .filter_data_16__30 (
             GND0), .filter_data_16__29 (GND0), .filter_data_16__28 (GND0), .filter_data_16__27 (
             GND0), .filter_data_16__26 (GND0), .filter_data_16__25 (GND0), .filter_data_16__24 (
             GND0), .filter_data_16__23 (GND0), .filter_data_16__22 (GND0), .filter_data_16__21 (
             GND0), .filter_data_16__20 (GND0), .filter_data_16__19 (GND0), .filter_data_16__18 (
             GND0), .filter_data_16__17 (GND0), .filter_data_16__16 (GND0), .filter_data_16__15 (
             GND0), .filter_data_16__14 (filter_data_16__14), .filter_data_16__13 (
             filter_data_16__13), .filter_data_16__12 (filter_data_16__12), .filter_data_16__11 (
             filter_data_16__11), .filter_data_16__10 (filter_data_16__10), .filter_data_16__9 (
             filter_data_16__9), .filter_data_16__8 (filter_data_16__8), .filter_data_16__7 (
             filter_data_16__7), .filter_data_16__6 (filter_data_16__6), .filter_data_16__5 (
             filter_data_16__5), .filter_data_16__4 (filter_data_16__4), .filter_data_16__3 (
             filter_data_16__3), .filter_data_16__2 (filter_data_16__2), .filter_data_16__1 (
             filter_data_16__1), .filter_data_16__0 (filter_data_16__0), .filter_data_17__31 (
             filter_data_17__15), .filter_data_17__30 (GND0), .filter_data_17__29 (
             GND0), .filter_data_17__28 (GND0), .filter_data_17__27 (GND0), .filter_data_17__26 (
             GND0), .filter_data_17__25 (GND0), .filter_data_17__24 (GND0), .filter_data_17__23 (
             GND0), .filter_data_17__22 (GND0), .filter_data_17__21 (GND0), .filter_data_17__20 (
             GND0), .filter_data_17__19 (GND0), .filter_data_17__18 (GND0), .filter_data_17__17 (
             GND0), .filter_data_17__16 (GND0), .filter_data_17__15 (GND0), .filter_data_17__14 (
             filter_data_17__14), .filter_data_17__13 (filter_data_17__13), .filter_data_17__12 (
             filter_data_17__12), .filter_data_17__11 (filter_data_17__11), .filter_data_17__10 (
             filter_data_17__10), .filter_data_17__9 (filter_data_17__9), .filter_data_17__8 (
             filter_data_17__8), .filter_data_17__7 (filter_data_17__7), .filter_data_17__6 (
             filter_data_17__6), .filter_data_17__5 (filter_data_17__5), .filter_data_17__4 (
             filter_data_17__4), .filter_data_17__3 (filter_data_17__3), .filter_data_17__2 (
             filter_data_17__2), .filter_data_17__1 (filter_data_17__1), .filter_data_17__0 (
             filter_data_17__0), .filter_data_18__31 (GND0), .filter_data_18__30 (
             GND0), .filter_data_18__29 (GND0), .filter_data_18__28 (GND0), .filter_data_18__27 (
             GND0), .filter_data_18__26 (GND0), .filter_data_18__25 (GND0), .filter_data_18__24 (
             GND0), .filter_data_18__23 (GND0), .filter_data_18__22 (GND0), .filter_data_18__21 (
             GND0), .filter_data_18__20 (GND0), .filter_data_18__19 (GND0), .filter_data_18__18 (
             GND0), .filter_data_18__17 (GND0), .filter_data_18__16 (GND0), .filter_data_18__15 (
             GND0), .filter_data_18__14 (GND0), .filter_data_18__13 (GND0), .filter_data_18__12 (
             GND0), .filter_data_18__11 (GND0), .filter_data_18__10 (GND0), .filter_data_18__9 (
             GND0), .filter_data_18__8 (GND0), .filter_data_18__7 (GND0), .filter_data_18__6 (
             GND0), .filter_data_18__5 (GND0), .filter_data_18__4 (GND0), .filter_data_18__3 (
             GND0), .filter_data_18__2 (GND0), .filter_data_18__1 (GND0), .filter_data_18__0 (
             GND0), .filter_data_19__31 (GND0), .filter_data_19__30 (GND0), .filter_data_19__29 (
             GND0), .filter_data_19__28 (GND0), .filter_data_19__27 (GND0), .filter_data_19__26 (
             GND0), .filter_data_19__25 (GND0), .filter_data_19__24 (GND0), .filter_data_19__23 (
             GND0), .filter_data_19__22 (GND0), .filter_data_19__21 (GND0), .filter_data_19__20 (
             GND0), .filter_data_19__19 (GND0), .filter_data_19__18 (GND0), .filter_data_19__17 (
             GND0), .filter_data_19__16 (GND0), .filter_data_19__15 (GND0), .filter_data_19__14 (
             GND0), .filter_data_19__13 (GND0), .filter_data_19__12 (GND0), .filter_data_19__11 (
             GND0), .filter_data_19__10 (GND0), .filter_data_19__9 (GND0), .filter_data_19__8 (
             GND0), .filter_data_19__7 (GND0), .filter_data_19__6 (GND0), .filter_data_19__5 (
             GND0), .filter_data_19__4 (GND0), .filter_data_19__3 (GND0), .filter_data_19__2 (
             GND0), .filter_data_19__1 (GND0), .filter_data_19__0 (GND0), .filter_data_20__31 (
             GND0), .filter_data_20__30 (GND0), .filter_data_20__29 (GND0), .filter_data_20__28 (
             GND0), .filter_data_20__27 (GND0), .filter_data_20__26 (GND0), .filter_data_20__25 (
             GND0), .filter_data_20__24 (GND0), .filter_data_20__23 (GND0), .filter_data_20__22 (
             GND0), .filter_data_20__21 (GND0), .filter_data_20__20 (GND0), .filter_data_20__19 (
             GND0), .filter_data_20__18 (GND0), .filter_data_20__17 (GND0), .filter_data_20__16 (
             GND0), .filter_data_20__15 (GND0), .filter_data_20__14 (GND0), .filter_data_20__13 (
             GND0), .filter_data_20__12 (GND0), .filter_data_20__11 (GND0), .filter_data_20__10 (
             GND0), .filter_data_20__9 (GND0), .filter_data_20__8 (GND0), .filter_data_20__7 (
             GND0), .filter_data_20__6 (GND0), .filter_data_20__5 (GND0), .filter_data_20__4 (
             GND0), .filter_data_20__3 (GND0), .filter_data_20__2 (GND0), .filter_data_20__1 (
             GND0), .filter_data_20__0 (GND0), .filter_data_21__31 (GND0), .filter_data_21__30 (
             GND0), .filter_data_21__29 (GND0), .filter_data_21__28 (GND0), .filter_data_21__27 (
             GND0), .filter_data_21__26 (GND0), .filter_data_21__25 (GND0), .filter_data_21__24 (
             GND0), .filter_data_21__23 (GND0), .filter_data_21__22 (GND0), .filter_data_21__21 (
             GND0), .filter_data_21__20 (GND0), .filter_data_21__19 (GND0), .filter_data_21__18 (
             GND0), .filter_data_21__17 (GND0), .filter_data_21__16 (GND0), .filter_data_21__15 (
             GND0), .filter_data_21__14 (GND0), .filter_data_21__13 (GND0), .filter_data_21__12 (
             GND0), .filter_data_21__11 (GND0), .filter_data_21__10 (GND0), .filter_data_21__9 (
             GND0), .filter_data_21__8 (GND0), .filter_data_21__7 (GND0), .filter_data_21__6 (
             GND0), .filter_data_21__5 (GND0), .filter_data_21__4 (GND0), .filter_data_21__3 (
             GND0), .filter_data_21__2 (GND0), .filter_data_21__1 (GND0), .filter_data_21__0 (
             GND0), .filter_data_22__31 (GND0), .filter_data_22__30 (GND0), .filter_data_22__29 (
             GND0), .filter_data_22__28 (GND0), .filter_data_22__27 (GND0), .filter_data_22__26 (
             GND0), .filter_data_22__25 (GND0), .filter_data_22__24 (GND0), .filter_data_22__23 (
             GND0), .filter_data_22__22 (GND0), .filter_data_22__21 (GND0), .filter_data_22__20 (
             GND0), .filter_data_22__19 (GND0), .filter_data_22__18 (GND0), .filter_data_22__17 (
             GND0), .filter_data_22__16 (GND0), .filter_data_22__15 (GND0), .filter_data_22__14 (
             GND0), .filter_data_22__13 (GND0), .filter_data_22__12 (GND0), .filter_data_22__11 (
             GND0), .filter_data_22__10 (GND0), .filter_data_22__9 (GND0), .filter_data_22__8 (
             GND0), .filter_data_22__7 (GND0), .filter_data_22__6 (GND0), .filter_data_22__5 (
             GND0), .filter_data_22__4 (GND0), .filter_data_22__3 (GND0), .filter_data_22__2 (
             GND0), .filter_data_22__1 (GND0), .filter_data_22__0 (GND0), .filter_data_23__31 (
             GND0), .filter_data_23__30 (GND0), .filter_data_23__29 (GND0), .filter_data_23__28 (
             GND0), .filter_data_23__27 (GND0), .filter_data_23__26 (GND0), .filter_data_23__25 (
             GND0), .filter_data_23__24 (GND0), .filter_data_23__23 (GND0), .filter_data_23__22 (
             GND0), .filter_data_23__21 (GND0), .filter_data_23__20 (GND0), .filter_data_23__19 (
             GND0), .filter_data_23__18 (GND0), .filter_data_23__17 (GND0), .filter_data_23__16 (
             GND0), .filter_data_23__15 (GND0), .filter_data_23__14 (GND0), .filter_data_23__13 (
             GND0), .filter_data_23__12 (GND0), .filter_data_23__11 (GND0), .filter_data_23__10 (
             GND0), .filter_data_23__9 (GND0), .filter_data_23__8 (GND0), .filter_data_23__7 (
             GND0), .filter_data_23__6 (GND0), .filter_data_23__5 (GND0), .filter_data_23__4 (
             GND0), .filter_data_23__3 (GND0), .filter_data_23__2 (GND0), .filter_data_23__1 (
             GND0), .filter_data_23__0 (GND0), .filter_data_24__31 (GND0), .filter_data_24__30 (
             GND0), .filter_data_24__29 (GND0), .filter_data_24__28 (GND0), .filter_data_24__27 (
             GND0), .filter_data_24__26 (GND0), .filter_data_24__25 (GND0), .filter_data_24__24 (
             GND0), .filter_data_24__23 (GND0), .filter_data_24__22 (GND0), .filter_data_24__21 (
             GND0), .filter_data_24__20 (GND0), .filter_data_24__19 (GND0), .filter_data_24__18 (
             GND0), .filter_data_24__17 (GND0), .filter_data_24__16 (GND0), .filter_data_24__15 (
             GND0), .filter_data_24__14 (GND0), .filter_data_24__13 (GND0), .filter_data_24__12 (
             GND0), .filter_data_24__11 (GND0), .filter_data_24__10 (GND0), .filter_data_24__9 (
             GND0), .filter_data_24__8 (GND0), .filter_data_24__7 (GND0), .filter_data_24__6 (
             GND0), .filter_data_24__5 (GND0), .filter_data_24__4 (GND0), .filter_data_24__3 (
             GND0), .filter_data_24__2 (GND0), .filter_data_24__1 (GND0), .filter_data_24__0 (
             GND0), .filter_size (nx16665), .ordered_img_data_0__31 (\$dummy [0]
             ), .ordered_img_data_0__30 (\$dummy [1]), .ordered_img_data_0__29 (
             \$dummy [2]), .ordered_img_data_0__28 (\$dummy [3]), .ordered_img_data_0__27 (
             \$dummy [4]), .ordered_img_data_0__26 (\$dummy [5]), .ordered_img_data_0__25 (
             \$dummy [6]), .ordered_img_data_0__24 (\$dummy [7]), .ordered_img_data_0__23 (
             \$dummy [8]), .ordered_img_data_0__22 (\$dummy [9]), .ordered_img_data_0__21 (
             \$dummy [10]), .ordered_img_data_0__20 (\$dummy [11]), .ordered_img_data_0__19 (
             \$dummy [12]), .ordered_img_data_0__18 (\$dummy [13]), .ordered_img_data_0__17 (
             \$dummy [14]), .ordered_img_data_0__16 (\$dummy [15]), .ordered_img_data_0__15 (
             \$dummy [16]), .ordered_img_data_0__14 (\$dummy [17]), .ordered_img_data_0__13 (
             \$dummy [18]), .ordered_img_data_0__12 (\$dummy [19]), .ordered_img_data_0__11 (
             \$dummy [20]), .ordered_img_data_0__10 (\$dummy [21]), .ordered_img_data_0__9 (
             \$dummy [22]), .ordered_img_data_0__8 (\$dummy [23]), .ordered_img_data_0__7 (
             \$dummy [24]), .ordered_img_data_0__6 (\$dummy [25]), .ordered_img_data_0__5 (
             \$dummy [26]), .ordered_img_data_0__4 (\$dummy [27]), .ordered_img_data_0__3 (
             \$dummy [28]), .ordered_img_data_0__2 (\$dummy [29]), .ordered_img_data_0__1 (
             \$dummy [30]), .ordered_img_data_0__0 (\$dummy [31]), .ordered_img_data_1__31 (
             \$dummy [32]), .ordered_img_data_1__30 (\$dummy [33]), .ordered_img_data_1__29 (
             \$dummy [34]), .ordered_img_data_1__28 (\$dummy [35]), .ordered_img_data_1__27 (
             \$dummy [36]), .ordered_img_data_1__26 (\$dummy [37]), .ordered_img_data_1__25 (
             \$dummy [38]), .ordered_img_data_1__24 (\$dummy [39]), .ordered_img_data_1__23 (
             \$dummy [40]), .ordered_img_data_1__22 (\$dummy [41]), .ordered_img_data_1__21 (
             \$dummy [42]), .ordered_img_data_1__20 (\$dummy [43]), .ordered_img_data_1__19 (
             \$dummy [44]), .ordered_img_data_1__18 (\$dummy [45]), .ordered_img_data_1__17 (
             \$dummy [46]), .ordered_img_data_1__16 (\$dummy [47]), .ordered_img_data_1__15 (
             \$dummy [48]), .ordered_img_data_1__14 (\$dummy [49]), .ordered_img_data_1__13 (
             \$dummy [50]), .ordered_img_data_1__12 (\$dummy [51]), .ordered_img_data_1__11 (
             \$dummy [52]), .ordered_img_data_1__10 (\$dummy [53]), .ordered_img_data_1__9 (
             \$dummy [54]), .ordered_img_data_1__8 (\$dummy [55]), .ordered_img_data_1__7 (
             \$dummy [56]), .ordered_img_data_1__6 (\$dummy [57]), .ordered_img_data_1__5 (
             \$dummy [58]), .ordered_img_data_1__4 (\$dummy [59]), .ordered_img_data_1__3 (
             \$dummy [60]), .ordered_img_data_1__2 (\$dummy [61]), .ordered_img_data_1__1 (
             \$dummy [62]), .ordered_img_data_1__0 (\$dummy [63]), .ordered_img_data_2__31 (
             \$dummy [64]), .ordered_img_data_2__30 (\$dummy [65]), .ordered_img_data_2__29 (
             \$dummy [66]), .ordered_img_data_2__28 (\$dummy [67]), .ordered_img_data_2__27 (
             \$dummy [68]), .ordered_img_data_2__26 (\$dummy [69]), .ordered_img_data_2__25 (
             \$dummy [70]), .ordered_img_data_2__24 (\$dummy [71]), .ordered_img_data_2__23 (
             \$dummy [72]), .ordered_img_data_2__22 (\$dummy [73]), .ordered_img_data_2__21 (
             \$dummy [74]), .ordered_img_data_2__20 (\$dummy [75]), .ordered_img_data_2__19 (
             \$dummy [76]), .ordered_img_data_2__18 (\$dummy [77]), .ordered_img_data_2__17 (
             \$dummy [78]), .ordered_img_data_2__16 (\$dummy [79]), .ordered_img_data_2__15 (
             \$dummy [80]), .ordered_img_data_2__14 (\$dummy [81]), .ordered_img_data_2__13 (
             \$dummy [82]), .ordered_img_data_2__12 (\$dummy [83]), .ordered_img_data_2__11 (
             \$dummy [84]), .ordered_img_data_2__10 (\$dummy [85]), .ordered_img_data_2__9 (
             \$dummy [86]), .ordered_img_data_2__8 (\$dummy [87]), .ordered_img_data_2__7 (
             \$dummy [88]), .ordered_img_data_2__6 (\$dummy [89]), .ordered_img_data_2__5 (
             \$dummy [90]), .ordered_img_data_2__4 (\$dummy [91]), .ordered_img_data_2__3 (
             \$dummy [92]), .ordered_img_data_2__2 (\$dummy [93]), .ordered_img_data_2__1 (
             \$dummy [94]), .ordered_img_data_2__0 (\$dummy [95]), .ordered_img_data_3__31 (
             \$dummy [96]), .ordered_img_data_3__30 (\$dummy [97]), .ordered_img_data_3__29 (
             \$dummy [98]), .ordered_img_data_3__28 (\$dummy [99]), .ordered_img_data_3__27 (
             \$dummy [100]), .ordered_img_data_3__26 (\$dummy [101]), .ordered_img_data_3__25 (
             \$dummy [102]), .ordered_img_data_3__24 (\$dummy [103]), .ordered_img_data_3__23 (
             \$dummy [104]), .ordered_img_data_3__22 (\$dummy [105]), .ordered_img_data_3__21 (
             \$dummy [106]), .ordered_img_data_3__20 (\$dummy [107]), .ordered_img_data_3__19 (
             \$dummy [108]), .ordered_img_data_3__18 (\$dummy [109]), .ordered_img_data_3__17 (
             \$dummy [110]), .ordered_img_data_3__16 (\$dummy [111]), .ordered_img_data_3__15 (
             \$dummy [112]), .ordered_img_data_3__14 (\$dummy [113]), .ordered_img_data_3__13 (
             \$dummy [114]), .ordered_img_data_3__12 (\$dummy [115]), .ordered_img_data_3__11 (
             \$dummy [116]), .ordered_img_data_3__10 (\$dummy [117]), .ordered_img_data_3__9 (
             \$dummy [118]), .ordered_img_data_3__8 (\$dummy [119]), .ordered_img_data_3__7 (
             \$dummy [120]), .ordered_img_data_3__6 (\$dummy [121]), .ordered_img_data_3__5 (
             \$dummy [122]), .ordered_img_data_3__4 (\$dummy [123]), .ordered_img_data_3__3 (
             \$dummy [124]), .ordered_img_data_3__2 (\$dummy [125]), .ordered_img_data_3__1 (
             \$dummy [126]), .ordered_img_data_3__0 (\$dummy [127]), .ordered_img_data_4__31 (
             \$dummy [128]), .ordered_img_data_4__30 (\$dummy [129]), .ordered_img_data_4__29 (
             \$dummy [130]), .ordered_img_data_4__28 (\$dummy [131]), .ordered_img_data_4__27 (
             \$dummy [132]), .ordered_img_data_4__26 (\$dummy [133]), .ordered_img_data_4__25 (
             \$dummy [134]), .ordered_img_data_4__24 (\$dummy [135]), .ordered_img_data_4__23 (
             \$dummy [136]), .ordered_img_data_4__22 (\$dummy [137]), .ordered_img_data_4__21 (
             \$dummy [138]), .ordered_img_data_4__20 (\$dummy [139]), .ordered_img_data_4__19 (
             \$dummy [140]), .ordered_img_data_4__18 (\$dummy [141]), .ordered_img_data_4__17 (
             \$dummy [142]), .ordered_img_data_4__16 (\$dummy [143]), .ordered_img_data_4__15 (
             \$dummy [144]), .ordered_img_data_4__14 (\$dummy [145]), .ordered_img_data_4__13 (
             \$dummy [146]), .ordered_img_data_4__12 (\$dummy [147]), .ordered_img_data_4__11 (
             \$dummy [148]), .ordered_img_data_4__10 (\$dummy [149]), .ordered_img_data_4__9 (
             \$dummy [150]), .ordered_img_data_4__8 (\$dummy [151]), .ordered_img_data_4__7 (
             \$dummy [152]), .ordered_img_data_4__6 (\$dummy [153]), .ordered_img_data_4__5 (
             \$dummy [154]), .ordered_img_data_4__4 (\$dummy [155]), .ordered_img_data_4__3 (
             \$dummy [156]), .ordered_img_data_4__2 (\$dummy [157]), .ordered_img_data_4__1 (
             \$dummy [158]), .ordered_img_data_4__0 (\$dummy [159]), .ordered_img_data_5__31 (
             \$dummy [160]), .ordered_img_data_5__30 (\$dummy [161]), .ordered_img_data_5__29 (
             \$dummy [162]), .ordered_img_data_5__28 (\$dummy [163]), .ordered_img_data_5__27 (
             \$dummy [164]), .ordered_img_data_5__26 (\$dummy [165]), .ordered_img_data_5__25 (
             \$dummy [166]), .ordered_img_data_5__24 (\$dummy [167]), .ordered_img_data_5__23 (
             \$dummy [168]), .ordered_img_data_5__22 (\$dummy [169]), .ordered_img_data_5__21 (
             \$dummy [170]), .ordered_img_data_5__20 (\$dummy [171]), .ordered_img_data_5__19 (
             \$dummy [172]), .ordered_img_data_5__18 (\$dummy [173]), .ordered_img_data_5__17 (
             \$dummy [174]), .ordered_img_data_5__16 (\$dummy [175]), .ordered_img_data_5__15 (
             \$dummy [176]), .ordered_img_data_5__14 (\$dummy [177]), .ordered_img_data_5__13 (
             \$dummy [178]), .ordered_img_data_5__12 (\$dummy [179]), .ordered_img_data_5__11 (
             \$dummy [180]), .ordered_img_data_5__10 (\$dummy [181]), .ordered_img_data_5__9 (
             \$dummy [182]), .ordered_img_data_5__8 (\$dummy [183]), .ordered_img_data_5__7 (
             \$dummy [184]), .ordered_img_data_5__6 (\$dummy [185]), .ordered_img_data_5__5 (
             \$dummy [186]), .ordered_img_data_5__4 (\$dummy [187]), .ordered_img_data_5__3 (
             \$dummy [188]), .ordered_img_data_5__2 (\$dummy [189]), .ordered_img_data_5__1 (
             \$dummy [190]), .ordered_img_data_5__0 (\$dummy [191]), .ordered_img_data_6__31 (
             \$dummy [192]), .ordered_img_data_6__30 (\$dummy [193]), .ordered_img_data_6__29 (
             \$dummy [194]), .ordered_img_data_6__28 (\$dummy [195]), .ordered_img_data_6__27 (
             \$dummy [196]), .ordered_img_data_6__26 (\$dummy [197]), .ordered_img_data_6__25 (
             \$dummy [198]), .ordered_img_data_6__24 (\$dummy [199]), .ordered_img_data_6__23 (
             \$dummy [200]), .ordered_img_data_6__22 (\$dummy [201]), .ordered_img_data_6__21 (
             \$dummy [202]), .ordered_img_data_6__20 (\$dummy [203]), .ordered_img_data_6__19 (
             \$dummy [204]), .ordered_img_data_6__18 (\$dummy [205]), .ordered_img_data_6__17 (
             \$dummy [206]), .ordered_img_data_6__16 (\$dummy [207]), .ordered_img_data_6__15 (
             \$dummy [208]), .ordered_img_data_6__14 (\$dummy [209]), .ordered_img_data_6__13 (
             \$dummy [210]), .ordered_img_data_6__12 (\$dummy [211]), .ordered_img_data_6__11 (
             \$dummy [212]), .ordered_img_data_6__10 (\$dummy [213]), .ordered_img_data_6__9 (
             \$dummy [214]), .ordered_img_data_6__8 (\$dummy [215]), .ordered_img_data_6__7 (
             \$dummy [216]), .ordered_img_data_6__6 (\$dummy [217]), .ordered_img_data_6__5 (
             \$dummy [218]), .ordered_img_data_6__4 (\$dummy [219]), .ordered_img_data_6__3 (
             \$dummy [220]), .ordered_img_data_6__2 (\$dummy [221]), .ordered_img_data_6__1 (
             \$dummy [222]), .ordered_img_data_6__0 (\$dummy [223]), .ordered_img_data_7__31 (
             \$dummy [224]), .ordered_img_data_7__30 (\$dummy [225]), .ordered_img_data_7__29 (
             \$dummy [226]), .ordered_img_data_7__28 (\$dummy [227]), .ordered_img_data_7__27 (
             \$dummy [228]), .ordered_img_data_7__26 (\$dummy [229]), .ordered_img_data_7__25 (
             \$dummy [230]), .ordered_img_data_7__24 (\$dummy [231]), .ordered_img_data_7__23 (
             \$dummy [232]), .ordered_img_data_7__22 (\$dummy [233]), .ordered_img_data_7__21 (
             \$dummy [234]), .ordered_img_data_7__20 (\$dummy [235]), .ordered_img_data_7__19 (
             \$dummy [236]), .ordered_img_data_7__18 (\$dummy [237]), .ordered_img_data_7__17 (
             \$dummy [238]), .ordered_img_data_7__16 (\$dummy [239]), .ordered_img_data_7__15 (
             \$dummy [240]), .ordered_img_data_7__14 (\$dummy [241]), .ordered_img_data_7__13 (
             \$dummy [242]), .ordered_img_data_7__12 (\$dummy [243]), .ordered_img_data_7__11 (
             \$dummy [244]), .ordered_img_data_7__10 (\$dummy [245]), .ordered_img_data_7__9 (
             \$dummy [246]), .ordered_img_data_7__8 (\$dummy [247]), .ordered_img_data_7__7 (
             \$dummy [248]), .ordered_img_data_7__6 (\$dummy [249]), .ordered_img_data_7__5 (
             \$dummy [250]), .ordered_img_data_7__4 (\$dummy [251]), .ordered_img_data_7__3 (
             \$dummy [252]), .ordered_img_data_7__2 (\$dummy [253]), .ordered_img_data_7__1 (
             \$dummy [254]), .ordered_img_data_7__0 (\$dummy [255]), .ordered_img_data_8__31 (
             \$dummy [256]), .ordered_img_data_8__30 (\$dummy [257]), .ordered_img_data_8__29 (
             \$dummy [258]), .ordered_img_data_8__28 (\$dummy [259]), .ordered_img_data_8__27 (
             \$dummy [260]), .ordered_img_data_8__26 (\$dummy [261]), .ordered_img_data_8__25 (
             \$dummy [262]), .ordered_img_data_8__24 (\$dummy [263]), .ordered_img_data_8__23 (
             \$dummy [264]), .ordered_img_data_8__22 (\$dummy [265]), .ordered_img_data_8__21 (
             \$dummy [266]), .ordered_img_data_8__20 (\$dummy [267]), .ordered_img_data_8__19 (
             \$dummy [268]), .ordered_img_data_8__18 (\$dummy [269]), .ordered_img_data_8__17 (
             \$dummy [270]), .ordered_img_data_8__16 (\$dummy [271]), .ordered_img_data_8__15 (
             \$dummy [272]), .ordered_img_data_8__14 (\$dummy [273]), .ordered_img_data_8__13 (
             \$dummy [274]), .ordered_img_data_8__12 (\$dummy [275]), .ordered_img_data_8__11 (
             \$dummy [276]), .ordered_img_data_8__10 (\$dummy [277]), .ordered_img_data_8__9 (
             \$dummy [278]), .ordered_img_data_8__8 (\$dummy [279]), .ordered_img_data_8__7 (
             \$dummy [280]), .ordered_img_data_8__6 (\$dummy [281]), .ordered_img_data_8__5 (
             \$dummy [282]), .ordered_img_data_8__4 (\$dummy [283]), .ordered_img_data_8__3 (
             \$dummy [284]), .ordered_img_data_8__2 (\$dummy [285]), .ordered_img_data_8__1 (
             \$dummy [286]), .ordered_img_data_8__0 (\$dummy [287]), .ordered_img_data_9__31 (
             ordered_img_data_9__31), .ordered_img_data_9__30 (\$dummy [288]), .ordered_img_data_9__29 (
             \$dummy [289]), .ordered_img_data_9__28 (\$dummy [290]), .ordered_img_data_9__27 (
             \$dummy [291]), .ordered_img_data_9__26 (\$dummy [292]), .ordered_img_data_9__25 (
             \$dummy [293]), .ordered_img_data_9__24 (\$dummy [294]), .ordered_img_data_9__23 (
             \$dummy [295]), .ordered_img_data_9__22 (\$dummy [296]), .ordered_img_data_9__21 (
             \$dummy [297]), .ordered_img_data_9__20 (\$dummy [298]), .ordered_img_data_9__19 (
             \$dummy [299]), .ordered_img_data_9__18 (\$dummy [300]), .ordered_img_data_9__17 (
             \$dummy [301]), .ordered_img_data_9__16 (\$dummy [302]), .ordered_img_data_9__15 (
             \$dummy [303]), .ordered_img_data_9__14 (ordered_img_data_9__14), .ordered_img_data_9__13 (
             ordered_img_data_9__13), .ordered_img_data_9__12 (
             ordered_img_data_9__12), .ordered_img_data_9__11 (
             ordered_img_data_9__11), .ordered_img_data_9__10 (
             ordered_img_data_9__10), .ordered_img_data_9__9 (
             ordered_img_data_9__9), .ordered_img_data_9__8 (
             ordered_img_data_9__8), .ordered_img_data_9__7 (
             ordered_img_data_9__7), .ordered_img_data_9__6 (
             ordered_img_data_9__6), .ordered_img_data_9__5 (
             ordered_img_data_9__5), .ordered_img_data_9__4 (
             ordered_img_data_9__4), .ordered_img_data_9__3 (
             ordered_img_data_9__3), .ordered_img_data_9__2 (
             ordered_img_data_9__2), .ordered_img_data_9__1 (
             ordered_img_data_9__1), .ordered_img_data_9__0 (
             ordered_img_data_9__0), .ordered_img_data_10__31 (
             ordered_img_data_10__31), .ordered_img_data_10__30 (\$dummy [304])
             , .ordered_img_data_10__29 (\$dummy [305]), .ordered_img_data_10__28 (
             \$dummy [306]), .ordered_img_data_10__27 (\$dummy [307]), .ordered_img_data_10__26 (
             \$dummy [308]), .ordered_img_data_10__25 (\$dummy [309]), .ordered_img_data_10__24 (
             \$dummy [310]), .ordered_img_data_10__23 (\$dummy [311]), .ordered_img_data_10__22 (
             \$dummy [312]), .ordered_img_data_10__21 (\$dummy [313]), .ordered_img_data_10__20 (
             \$dummy [314]), .ordered_img_data_10__19 (\$dummy [315]), .ordered_img_data_10__18 (
             \$dummy [316]), .ordered_img_data_10__17 (\$dummy [317]), .ordered_img_data_10__16 (
             \$dummy [318]), .ordered_img_data_10__15 (\$dummy [319]), .ordered_img_data_10__14 (
             ordered_img_data_10__14), .ordered_img_data_10__13 (
             ordered_img_data_10__13), .ordered_img_data_10__12 (
             ordered_img_data_10__12), .ordered_img_data_10__11 (
             ordered_img_data_10__11), .ordered_img_data_10__10 (
             ordered_img_data_10__10), .ordered_img_data_10__9 (
             ordered_img_data_10__9), .ordered_img_data_10__8 (
             ordered_img_data_10__8), .ordered_img_data_10__7 (
             ordered_img_data_10__7), .ordered_img_data_10__6 (
             ordered_img_data_10__6), .ordered_img_data_10__5 (
             ordered_img_data_10__5), .ordered_img_data_10__4 (
             ordered_img_data_10__4), .ordered_img_data_10__3 (
             ordered_img_data_10__3), .ordered_img_data_10__2 (
             ordered_img_data_10__2), .ordered_img_data_10__1 (
             ordered_img_data_10__1), .ordered_img_data_10__0 (
             ordered_img_data_10__0), .ordered_img_data_11__31 (
             ordered_img_data_11__31), .ordered_img_data_11__30 (\$dummy [320])
             , .ordered_img_data_11__29 (\$dummy [321]), .ordered_img_data_11__28 (
             \$dummy [322]), .ordered_img_data_11__27 (\$dummy [323]), .ordered_img_data_11__26 (
             \$dummy [324]), .ordered_img_data_11__25 (\$dummy [325]), .ordered_img_data_11__24 (
             \$dummy [326]), .ordered_img_data_11__23 (\$dummy [327]), .ordered_img_data_11__22 (
             \$dummy [328]), .ordered_img_data_11__21 (\$dummy [329]), .ordered_img_data_11__20 (
             \$dummy [330]), .ordered_img_data_11__19 (\$dummy [331]), .ordered_img_data_11__18 (
             \$dummy [332]), .ordered_img_data_11__17 (\$dummy [333]), .ordered_img_data_11__16 (
             \$dummy [334]), .ordered_img_data_11__15 (\$dummy [335]), .ordered_img_data_11__14 (
             ordered_img_data_11__14), .ordered_img_data_11__13 (
             ordered_img_data_11__13), .ordered_img_data_11__12 (
             ordered_img_data_11__12), .ordered_img_data_11__11 (
             ordered_img_data_11__11), .ordered_img_data_11__10 (
             ordered_img_data_11__10), .ordered_img_data_11__9 (
             ordered_img_data_11__9), .ordered_img_data_11__8 (
             ordered_img_data_11__8), .ordered_img_data_11__7 (
             ordered_img_data_11__7), .ordered_img_data_11__6 (
             ordered_img_data_11__6), .ordered_img_data_11__5 (
             ordered_img_data_11__5), .ordered_img_data_11__4 (
             ordered_img_data_11__4), .ordered_img_data_11__3 (
             ordered_img_data_11__3), .ordered_img_data_11__2 (
             ordered_img_data_11__2), .ordered_img_data_11__1 (
             ordered_img_data_11__1), .ordered_img_data_11__0 (
             ordered_img_data_11__0), .ordered_img_data_12__31 (
             ordered_img_data_12__31), .ordered_img_data_12__30 (\$dummy [336])
             , .ordered_img_data_12__29 (\$dummy [337]), .ordered_img_data_12__28 (
             \$dummy [338]), .ordered_img_data_12__27 (\$dummy [339]), .ordered_img_data_12__26 (
             \$dummy [340]), .ordered_img_data_12__25 (\$dummy [341]), .ordered_img_data_12__24 (
             \$dummy [342]), .ordered_img_data_12__23 (\$dummy [343]), .ordered_img_data_12__22 (
             \$dummy [344]), .ordered_img_data_12__21 (\$dummy [345]), .ordered_img_data_12__20 (
             \$dummy [346]), .ordered_img_data_12__19 (\$dummy [347]), .ordered_img_data_12__18 (
             \$dummy [348]), .ordered_img_data_12__17 (\$dummy [349]), .ordered_img_data_12__16 (
             \$dummy [350]), .ordered_img_data_12__15 (\$dummy [351]), .ordered_img_data_12__14 (
             ordered_img_data_12__14), .ordered_img_data_12__13 (
             ordered_img_data_12__13), .ordered_img_data_12__12 (
             ordered_img_data_12__12), .ordered_img_data_12__11 (
             ordered_img_data_12__11), .ordered_img_data_12__10 (
             ordered_img_data_12__10), .ordered_img_data_12__9 (
             ordered_img_data_12__9), .ordered_img_data_12__8 (
             ordered_img_data_12__8), .ordered_img_data_12__7 (
             ordered_img_data_12__7), .ordered_img_data_12__6 (
             ordered_img_data_12__6), .ordered_img_data_12__5 (
             ordered_img_data_12__5), .ordered_img_data_12__4 (
             ordered_img_data_12__4), .ordered_img_data_12__3 (
             ordered_img_data_12__3), .ordered_img_data_12__2 (
             ordered_img_data_12__2), .ordered_img_data_12__1 (
             ordered_img_data_12__1), .ordered_img_data_12__0 (
             ordered_img_data_12__0), .ordered_img_data_13__31 (
             ordered_img_data_13__31), .ordered_img_data_13__30 (\$dummy [352])
             , .ordered_img_data_13__29 (\$dummy [353]), .ordered_img_data_13__28 (
             \$dummy [354]), .ordered_img_data_13__27 (\$dummy [355]), .ordered_img_data_13__26 (
             \$dummy [356]), .ordered_img_data_13__25 (\$dummy [357]), .ordered_img_data_13__24 (
             \$dummy [358]), .ordered_img_data_13__23 (\$dummy [359]), .ordered_img_data_13__22 (
             \$dummy [360]), .ordered_img_data_13__21 (\$dummy [361]), .ordered_img_data_13__20 (
             \$dummy [362]), .ordered_img_data_13__19 (\$dummy [363]), .ordered_img_data_13__18 (
             \$dummy [364]), .ordered_img_data_13__17 (\$dummy [365]), .ordered_img_data_13__16 (
             \$dummy [366]), .ordered_img_data_13__15 (\$dummy [367]), .ordered_img_data_13__14 (
             ordered_img_data_13__14), .ordered_img_data_13__13 (
             ordered_img_data_13__13), .ordered_img_data_13__12 (
             ordered_img_data_13__12), .ordered_img_data_13__11 (
             ordered_img_data_13__11), .ordered_img_data_13__10 (
             ordered_img_data_13__10), .ordered_img_data_13__9 (
             ordered_img_data_13__9), .ordered_img_data_13__8 (
             ordered_img_data_13__8), .ordered_img_data_13__7 (
             ordered_img_data_13__7), .ordered_img_data_13__6 (
             ordered_img_data_13__6), .ordered_img_data_13__5 (
             ordered_img_data_13__5), .ordered_img_data_13__4 (
             ordered_img_data_13__4), .ordered_img_data_13__3 (
             ordered_img_data_13__3), .ordered_img_data_13__2 (
             ordered_img_data_13__2), .ordered_img_data_13__1 (
             ordered_img_data_13__1), .ordered_img_data_13__0 (
             ordered_img_data_13__0), .ordered_img_data_14__31 (
             ordered_img_data_14__31), .ordered_img_data_14__30 (\$dummy [368])
             , .ordered_img_data_14__29 (\$dummy [369]), .ordered_img_data_14__28 (
             \$dummy [370]), .ordered_img_data_14__27 (\$dummy [371]), .ordered_img_data_14__26 (
             \$dummy [372]), .ordered_img_data_14__25 (\$dummy [373]), .ordered_img_data_14__24 (
             \$dummy [374]), .ordered_img_data_14__23 (\$dummy [375]), .ordered_img_data_14__22 (
             \$dummy [376]), .ordered_img_data_14__21 (\$dummy [377]), .ordered_img_data_14__20 (
             \$dummy [378]), .ordered_img_data_14__19 (\$dummy [379]), .ordered_img_data_14__18 (
             \$dummy [380]), .ordered_img_data_14__17 (\$dummy [381]), .ordered_img_data_14__16 (
             \$dummy [382]), .ordered_img_data_14__15 (\$dummy [383]), .ordered_img_data_14__14 (
             ordered_img_data_14__14), .ordered_img_data_14__13 (
             ordered_img_data_14__13), .ordered_img_data_14__12 (
             ordered_img_data_14__12), .ordered_img_data_14__11 (
             ordered_img_data_14__11), .ordered_img_data_14__10 (
             ordered_img_data_14__10), .ordered_img_data_14__9 (
             ordered_img_data_14__9), .ordered_img_data_14__8 (
             ordered_img_data_14__8), .ordered_img_data_14__7 (
             ordered_img_data_14__7), .ordered_img_data_14__6 (
             ordered_img_data_14__6), .ordered_img_data_14__5 (
             ordered_img_data_14__5), .ordered_img_data_14__4 (
             ordered_img_data_14__4), .ordered_img_data_14__3 (
             ordered_img_data_14__3), .ordered_img_data_14__2 (
             ordered_img_data_14__2), .ordered_img_data_14__1 (
             ordered_img_data_14__1), .ordered_img_data_14__0 (
             ordered_img_data_14__0), .ordered_img_data_15__31 (
             ordered_img_data_15__31), .ordered_img_data_15__30 (\$dummy [384])
             , .ordered_img_data_15__29 (\$dummy [385]), .ordered_img_data_15__28 (
             \$dummy [386]), .ordered_img_data_15__27 (\$dummy [387]), .ordered_img_data_15__26 (
             \$dummy [388]), .ordered_img_data_15__25 (\$dummy [389]), .ordered_img_data_15__24 (
             \$dummy [390]), .ordered_img_data_15__23 (\$dummy [391]), .ordered_img_data_15__22 (
             \$dummy [392]), .ordered_img_data_15__21 (\$dummy [393]), .ordered_img_data_15__20 (
             \$dummy [394]), .ordered_img_data_15__19 (\$dummy [395]), .ordered_img_data_15__18 (
             \$dummy [396]), .ordered_img_data_15__17 (\$dummy [397]), .ordered_img_data_15__16 (
             \$dummy [398]), .ordered_img_data_15__15 (\$dummy [399]), .ordered_img_data_15__14 (
             ordered_img_data_15__14), .ordered_img_data_15__13 (
             ordered_img_data_15__13), .ordered_img_data_15__12 (
             ordered_img_data_15__12), .ordered_img_data_15__11 (
             ordered_img_data_15__11), .ordered_img_data_15__10 (
             ordered_img_data_15__10), .ordered_img_data_15__9 (
             ordered_img_data_15__9), .ordered_img_data_15__8 (
             ordered_img_data_15__8), .ordered_img_data_15__7 (
             ordered_img_data_15__7), .ordered_img_data_15__6 (
             ordered_img_data_15__6), .ordered_img_data_15__5 (
             ordered_img_data_15__5), .ordered_img_data_15__4 (
             ordered_img_data_15__4), .ordered_img_data_15__3 (
             ordered_img_data_15__3), .ordered_img_data_15__2 (
             ordered_img_data_15__2), .ordered_img_data_15__1 (
             ordered_img_data_15__1), .ordered_img_data_15__0 (
             ordered_img_data_15__0), .ordered_img_data_16__31 (
             ordered_img_data_16__31), .ordered_img_data_16__30 (\$dummy [400])
             , .ordered_img_data_16__29 (\$dummy [401]), .ordered_img_data_16__28 (
             \$dummy [402]), .ordered_img_data_16__27 (\$dummy [403]), .ordered_img_data_16__26 (
             \$dummy [404]), .ordered_img_data_16__25 (\$dummy [405]), .ordered_img_data_16__24 (
             \$dummy [406]), .ordered_img_data_16__23 (\$dummy [407]), .ordered_img_data_16__22 (
             \$dummy [408]), .ordered_img_data_16__21 (\$dummy [409]), .ordered_img_data_16__20 (
             \$dummy [410]), .ordered_img_data_16__19 (\$dummy [411]), .ordered_img_data_16__18 (
             \$dummy [412]), .ordered_img_data_16__17 (\$dummy [413]), .ordered_img_data_16__16 (
             \$dummy [414]), .ordered_img_data_16__15 (\$dummy [415]), .ordered_img_data_16__14 (
             ordered_img_data_16__14), .ordered_img_data_16__13 (
             ordered_img_data_16__13), .ordered_img_data_16__12 (
             ordered_img_data_16__12), .ordered_img_data_16__11 (
             ordered_img_data_16__11), .ordered_img_data_16__10 (
             ordered_img_data_16__10), .ordered_img_data_16__9 (
             ordered_img_data_16__9), .ordered_img_data_16__8 (
             ordered_img_data_16__8), .ordered_img_data_16__7 (
             ordered_img_data_16__7), .ordered_img_data_16__6 (
             ordered_img_data_16__6), .ordered_img_data_16__5 (
             ordered_img_data_16__5), .ordered_img_data_16__4 (
             ordered_img_data_16__4), .ordered_img_data_16__3 (
             ordered_img_data_16__3), .ordered_img_data_16__2 (
             ordered_img_data_16__2), .ordered_img_data_16__1 (
             ordered_img_data_16__1), .ordered_img_data_16__0 (
             ordered_img_data_16__0), .ordered_img_data_17__31 (
             ordered_img_data_17__31), .ordered_img_data_17__30 (\$dummy [416])
             , .ordered_img_data_17__29 (\$dummy [417]), .ordered_img_data_17__28 (
             \$dummy [418]), .ordered_img_data_17__27 (\$dummy [419]), .ordered_img_data_17__26 (
             \$dummy [420]), .ordered_img_data_17__25 (\$dummy [421]), .ordered_img_data_17__24 (
             \$dummy [422]), .ordered_img_data_17__23 (\$dummy [423]), .ordered_img_data_17__22 (
             \$dummy [424]), .ordered_img_data_17__21 (\$dummy [425]), .ordered_img_data_17__20 (
             \$dummy [426]), .ordered_img_data_17__19 (\$dummy [427]), .ordered_img_data_17__18 (
             \$dummy [428]), .ordered_img_data_17__17 (\$dummy [429]), .ordered_img_data_17__16 (
             \$dummy [430]), .ordered_img_data_17__15 (\$dummy [431]), .ordered_img_data_17__14 (
             ordered_img_data_17__14), .ordered_img_data_17__13 (
             ordered_img_data_17__13), .ordered_img_data_17__12 (
             ordered_img_data_17__12), .ordered_img_data_17__11 (
             ordered_img_data_17__11), .ordered_img_data_17__10 (
             ordered_img_data_17__10), .ordered_img_data_17__9 (
             ordered_img_data_17__9), .ordered_img_data_17__8 (
             ordered_img_data_17__8), .ordered_img_data_17__7 (
             ordered_img_data_17__7), .ordered_img_data_17__6 (
             ordered_img_data_17__6), .ordered_img_data_17__5 (
             ordered_img_data_17__5), .ordered_img_data_17__4 (
             ordered_img_data_17__4), .ordered_img_data_17__3 (
             ordered_img_data_17__3), .ordered_img_data_17__2 (
             ordered_img_data_17__2), .ordered_img_data_17__1 (
             ordered_img_data_17__1), .ordered_img_data_17__0 (
             ordered_img_data_17__0), .ordered_img_data_18__31 (\$dummy [432]), 
             .ordered_img_data_18__30 (\$dummy [433]), .ordered_img_data_18__29 (
             \$dummy [434]), .ordered_img_data_18__28 (\$dummy [435]), .ordered_img_data_18__27 (
             \$dummy [436]), .ordered_img_data_18__26 (\$dummy [437]), .ordered_img_data_18__25 (
             \$dummy [438]), .ordered_img_data_18__24 (\$dummy [439]), .ordered_img_data_18__23 (
             \$dummy [440]), .ordered_img_data_18__22 (\$dummy [441]), .ordered_img_data_18__21 (
             \$dummy [442]), .ordered_img_data_18__20 (\$dummy [443]), .ordered_img_data_18__19 (
             \$dummy [444]), .ordered_img_data_18__18 (\$dummy [445]), .ordered_img_data_18__17 (
             \$dummy [446]), .ordered_img_data_18__16 (\$dummy [447]), .ordered_img_data_18__15 (
             \$dummy [448]), .ordered_img_data_18__14 (\$dummy [449]), .ordered_img_data_18__13 (
             \$dummy [450]), .ordered_img_data_18__12 (\$dummy [451]), .ordered_img_data_18__11 (
             \$dummy [452]), .ordered_img_data_18__10 (\$dummy [453]), .ordered_img_data_18__9 (
             \$dummy [454]), .ordered_img_data_18__8 (\$dummy [455]), .ordered_img_data_18__7 (
             \$dummy [456]), .ordered_img_data_18__6 (\$dummy [457]), .ordered_img_data_18__5 (
             \$dummy [458]), .ordered_img_data_18__4 (\$dummy [459]), .ordered_img_data_18__3 (
             \$dummy [460]), .ordered_img_data_18__2 (\$dummy [461]), .ordered_img_data_18__1 (
             \$dummy [462]), .ordered_img_data_18__0 (\$dummy [463]), .ordered_img_data_19__31 (
             \$dummy [464]), .ordered_img_data_19__30 (\$dummy [465]), .ordered_img_data_19__29 (
             \$dummy [466]), .ordered_img_data_19__28 (\$dummy [467]), .ordered_img_data_19__27 (
             \$dummy [468]), .ordered_img_data_19__26 (\$dummy [469]), .ordered_img_data_19__25 (
             \$dummy [470]), .ordered_img_data_19__24 (\$dummy [471]), .ordered_img_data_19__23 (
             \$dummy [472]), .ordered_img_data_19__22 (\$dummy [473]), .ordered_img_data_19__21 (
             \$dummy [474]), .ordered_img_data_19__20 (\$dummy [475]), .ordered_img_data_19__19 (
             \$dummy [476]), .ordered_img_data_19__18 (\$dummy [477]), .ordered_img_data_19__17 (
             \$dummy [478]), .ordered_img_data_19__16 (\$dummy [479]), .ordered_img_data_19__15 (
             \$dummy [480]), .ordered_img_data_19__14 (\$dummy [481]), .ordered_img_data_19__13 (
             \$dummy [482]), .ordered_img_data_19__12 (\$dummy [483]), .ordered_img_data_19__11 (
             \$dummy [484]), .ordered_img_data_19__10 (\$dummy [485]), .ordered_img_data_19__9 (
             \$dummy [486]), .ordered_img_data_19__8 (\$dummy [487]), .ordered_img_data_19__7 (
             \$dummy [488]), .ordered_img_data_19__6 (\$dummy [489]), .ordered_img_data_19__5 (
             \$dummy [490]), .ordered_img_data_19__4 (\$dummy [491]), .ordered_img_data_19__3 (
             \$dummy [492]), .ordered_img_data_19__2 (\$dummy [493]), .ordered_img_data_19__1 (
             \$dummy [494]), .ordered_img_data_19__0 (\$dummy [495]), .ordered_img_data_20__31 (
             \$dummy [496]), .ordered_img_data_20__30 (\$dummy [497]), .ordered_img_data_20__29 (
             \$dummy [498]), .ordered_img_data_20__28 (\$dummy [499]), .ordered_img_data_20__27 (
             \$dummy [500]), .ordered_img_data_20__26 (\$dummy [501]), .ordered_img_data_20__25 (
             \$dummy [502]), .ordered_img_data_20__24 (\$dummy [503]), .ordered_img_data_20__23 (
             \$dummy [504]), .ordered_img_data_20__22 (\$dummy [505]), .ordered_img_data_20__21 (
             \$dummy [506]), .ordered_img_data_20__20 (\$dummy [507]), .ordered_img_data_20__19 (
             \$dummy [508]), .ordered_img_data_20__18 (\$dummy [509]), .ordered_img_data_20__17 (
             \$dummy [510]), .ordered_img_data_20__16 (\$dummy [511]), .ordered_img_data_20__15 (
             \$dummy [512]), .ordered_img_data_20__14 (\$dummy [513]), .ordered_img_data_20__13 (
             \$dummy [514]), .ordered_img_data_20__12 (\$dummy [515]), .ordered_img_data_20__11 (
             \$dummy [516]), .ordered_img_data_20__10 (\$dummy [517]), .ordered_img_data_20__9 (
             \$dummy [518]), .ordered_img_data_20__8 (\$dummy [519]), .ordered_img_data_20__7 (
             \$dummy [520]), .ordered_img_data_20__6 (\$dummy [521]), .ordered_img_data_20__5 (
             \$dummy [522]), .ordered_img_data_20__4 (\$dummy [523]), .ordered_img_data_20__3 (
             \$dummy [524]), .ordered_img_data_20__2 (\$dummy [525]), .ordered_img_data_20__1 (
             \$dummy [526]), .ordered_img_data_20__0 (\$dummy [527]), .ordered_img_data_21__31 (
             \$dummy [528]), .ordered_img_data_21__30 (\$dummy [529]), .ordered_img_data_21__29 (
             \$dummy [530]), .ordered_img_data_21__28 (\$dummy [531]), .ordered_img_data_21__27 (
             \$dummy [532]), .ordered_img_data_21__26 (\$dummy [533]), .ordered_img_data_21__25 (
             \$dummy [534]), .ordered_img_data_21__24 (\$dummy [535]), .ordered_img_data_21__23 (
             \$dummy [536]), .ordered_img_data_21__22 (\$dummy [537]), .ordered_img_data_21__21 (
             \$dummy [538]), .ordered_img_data_21__20 (\$dummy [539]), .ordered_img_data_21__19 (
             \$dummy [540]), .ordered_img_data_21__18 (\$dummy [541]), .ordered_img_data_21__17 (
             \$dummy [542]), .ordered_img_data_21__16 (\$dummy [543]), .ordered_img_data_21__15 (
             \$dummy [544]), .ordered_img_data_21__14 (\$dummy [545]), .ordered_img_data_21__13 (
             \$dummy [546]), .ordered_img_data_21__12 (\$dummy [547]), .ordered_img_data_21__11 (
             \$dummy [548]), .ordered_img_data_21__10 (\$dummy [549]), .ordered_img_data_21__9 (
             \$dummy [550]), .ordered_img_data_21__8 (\$dummy [551]), .ordered_img_data_21__7 (
             \$dummy [552]), .ordered_img_data_21__6 (\$dummy [553]), .ordered_img_data_21__5 (
             \$dummy [554]), .ordered_img_data_21__4 (\$dummy [555]), .ordered_img_data_21__3 (
             \$dummy [556]), .ordered_img_data_21__2 (\$dummy [557]), .ordered_img_data_21__1 (
             \$dummy [558]), .ordered_img_data_21__0 (\$dummy [559]), .ordered_img_data_22__31 (
             \$dummy [560]), .ordered_img_data_22__30 (\$dummy [561]), .ordered_img_data_22__29 (
             \$dummy [562]), .ordered_img_data_22__28 (\$dummy [563]), .ordered_img_data_22__27 (
             \$dummy [564]), .ordered_img_data_22__26 (\$dummy [565]), .ordered_img_data_22__25 (
             \$dummy [566]), .ordered_img_data_22__24 (\$dummy [567]), .ordered_img_data_22__23 (
             \$dummy [568]), .ordered_img_data_22__22 (\$dummy [569]), .ordered_img_data_22__21 (
             \$dummy [570]), .ordered_img_data_22__20 (\$dummy [571]), .ordered_img_data_22__19 (
             \$dummy [572]), .ordered_img_data_22__18 (\$dummy [573]), .ordered_img_data_22__17 (
             \$dummy [574]), .ordered_img_data_22__16 (\$dummy [575]), .ordered_img_data_22__15 (
             \$dummy [576]), .ordered_img_data_22__14 (\$dummy [577]), .ordered_img_data_22__13 (
             \$dummy [578]), .ordered_img_data_22__12 (\$dummy [579]), .ordered_img_data_22__11 (
             \$dummy [580]), .ordered_img_data_22__10 (\$dummy [581]), .ordered_img_data_22__9 (
             \$dummy [582]), .ordered_img_data_22__8 (\$dummy [583]), .ordered_img_data_22__7 (
             \$dummy [584]), .ordered_img_data_22__6 (\$dummy [585]), .ordered_img_data_22__5 (
             \$dummy [586]), .ordered_img_data_22__4 (\$dummy [587]), .ordered_img_data_22__3 (
             \$dummy [588]), .ordered_img_data_22__2 (\$dummy [589]), .ordered_img_data_22__1 (
             \$dummy [590]), .ordered_img_data_22__0 (\$dummy [591]), .ordered_img_data_23__31 (
             \$dummy [592]), .ordered_img_data_23__30 (\$dummy [593]), .ordered_img_data_23__29 (
             \$dummy [594]), .ordered_img_data_23__28 (\$dummy [595]), .ordered_img_data_23__27 (
             \$dummy [596]), .ordered_img_data_23__26 (\$dummy [597]), .ordered_img_data_23__25 (
             \$dummy [598]), .ordered_img_data_23__24 (\$dummy [599]), .ordered_img_data_23__23 (
             \$dummy [600]), .ordered_img_data_23__22 (\$dummy [601]), .ordered_img_data_23__21 (
             \$dummy [602]), .ordered_img_data_23__20 (\$dummy [603]), .ordered_img_data_23__19 (
             \$dummy [604]), .ordered_img_data_23__18 (\$dummy [605]), .ordered_img_data_23__17 (
             \$dummy [606]), .ordered_img_data_23__16 (\$dummy [607]), .ordered_img_data_23__15 (
             \$dummy [608]), .ordered_img_data_23__14 (\$dummy [609]), .ordered_img_data_23__13 (
             \$dummy [610]), .ordered_img_data_23__12 (\$dummy [611]), .ordered_img_data_23__11 (
             \$dummy [612]), .ordered_img_data_23__10 (\$dummy [613]), .ordered_img_data_23__9 (
             \$dummy [614]), .ordered_img_data_23__8 (\$dummy [615]), .ordered_img_data_23__7 (
             \$dummy [616]), .ordered_img_data_23__6 (\$dummy [617]), .ordered_img_data_23__5 (
             \$dummy [618]), .ordered_img_data_23__4 (\$dummy [619]), .ordered_img_data_23__3 (
             \$dummy [620]), .ordered_img_data_23__2 (\$dummy [621]), .ordered_img_data_23__1 (
             \$dummy [622]), .ordered_img_data_23__0 (\$dummy [623]), .ordered_img_data_24__31 (
             \$dummy [624]), .ordered_img_data_24__30 (\$dummy [625]), .ordered_img_data_24__29 (
             \$dummy [626]), .ordered_img_data_24__28 (\$dummy [627]), .ordered_img_data_24__27 (
             \$dummy [628]), .ordered_img_data_24__26 (\$dummy [629]), .ordered_img_data_24__25 (
             \$dummy [630]), .ordered_img_data_24__24 (\$dummy [631]), .ordered_img_data_24__23 (
             \$dummy [632]), .ordered_img_data_24__22 (\$dummy [633]), .ordered_img_data_24__21 (
             \$dummy [634]), .ordered_img_data_24__20 (\$dummy [635]), .ordered_img_data_24__19 (
             \$dummy [636]), .ordered_img_data_24__18 (\$dummy [637]), .ordered_img_data_24__17 (
             \$dummy [638]), .ordered_img_data_24__16 (\$dummy [639]), .ordered_img_data_24__15 (
             \$dummy [640]), .ordered_img_data_24__14 (\$dummy [641]), .ordered_img_data_24__13 (
             \$dummy [642]), .ordered_img_data_24__12 (\$dummy [643]), .ordered_img_data_24__11 (
             \$dummy [644]), .ordered_img_data_24__10 (\$dummy [645]), .ordered_img_data_24__9 (
             \$dummy [646]), .ordered_img_data_24__8 (\$dummy [647]), .ordered_img_data_24__7 (
             \$dummy [648]), .ordered_img_data_24__6 (\$dummy [649]), .ordered_img_data_24__5 (
             \$dummy [650]), .ordered_img_data_24__4 (\$dummy [651]), .ordered_img_data_24__3 (
             \$dummy [652]), .ordered_img_data_24__2 (\$dummy [653]), .ordered_img_data_24__1 (
             \$dummy [654]), .ordered_img_data_24__0 (\$dummy [655]), .ordered_filter_data_0__31 (
             \$dummy [656]), .ordered_filter_data_0__30 (\$dummy [657]), .ordered_filter_data_0__29 (
             \$dummy [658]), .ordered_filter_data_0__28 (\$dummy [659]), .ordered_filter_data_0__27 (
             \$dummy [660]), .ordered_filter_data_0__26 (\$dummy [661]), .ordered_filter_data_0__25 (
             \$dummy [662]), .ordered_filter_data_0__24 (\$dummy [663]), .ordered_filter_data_0__23 (
             \$dummy [664]), .ordered_filter_data_0__22 (\$dummy [665]), .ordered_filter_data_0__21 (
             \$dummy [666]), .ordered_filter_data_0__20 (\$dummy [667]), .ordered_filter_data_0__19 (
             \$dummy [668]), .ordered_filter_data_0__18 (\$dummy [669]), .ordered_filter_data_0__17 (
             \$dummy [670]), .ordered_filter_data_0__16 (\$dummy [671]), .ordered_filter_data_0__15 (
             \$dummy [672]), .ordered_filter_data_0__14 (\$dummy [673]), .ordered_filter_data_0__13 (
             \$dummy [674]), .ordered_filter_data_0__12 (\$dummy [675]), .ordered_filter_data_0__11 (
             \$dummy [676]), .ordered_filter_data_0__10 (\$dummy [677]), .ordered_filter_data_0__9 (
             \$dummy [678]), .ordered_filter_data_0__8 (\$dummy [679]), .ordered_filter_data_0__7 (
             \$dummy [680]), .ordered_filter_data_0__6 (\$dummy [681]), .ordered_filter_data_0__5 (
             \$dummy [682]), .ordered_filter_data_0__4 (\$dummy [683]), .ordered_filter_data_0__3 (
             \$dummy [684]), .ordered_filter_data_0__2 (\$dummy [685]), .ordered_filter_data_0__1 (
             \$dummy [686]), .ordered_filter_data_0__0 (\$dummy [687]), .ordered_filter_data_1__31 (
             \$dummy [688]), .ordered_filter_data_1__30 (\$dummy [689]), .ordered_filter_data_1__29 (
             \$dummy [690]), .ordered_filter_data_1__28 (\$dummy [691]), .ordered_filter_data_1__27 (
             \$dummy [692]), .ordered_filter_data_1__26 (\$dummy [693]), .ordered_filter_data_1__25 (
             \$dummy [694]), .ordered_filter_data_1__24 (\$dummy [695]), .ordered_filter_data_1__23 (
             \$dummy [696]), .ordered_filter_data_1__22 (\$dummy [697]), .ordered_filter_data_1__21 (
             \$dummy [698]), .ordered_filter_data_1__20 (\$dummy [699]), .ordered_filter_data_1__19 (
             \$dummy [700]), .ordered_filter_data_1__18 (\$dummy [701]), .ordered_filter_data_1__17 (
             \$dummy [702]), .ordered_filter_data_1__16 (\$dummy [703]), .ordered_filter_data_1__15 (
             \$dummy [704]), .ordered_filter_data_1__14 (\$dummy [705]), .ordered_filter_data_1__13 (
             \$dummy [706]), .ordered_filter_data_1__12 (\$dummy [707]), .ordered_filter_data_1__11 (
             \$dummy [708]), .ordered_filter_data_1__10 (\$dummy [709]), .ordered_filter_data_1__9 (
             \$dummy [710]), .ordered_filter_data_1__8 (\$dummy [711]), .ordered_filter_data_1__7 (
             \$dummy [712]), .ordered_filter_data_1__6 (\$dummy [713]), .ordered_filter_data_1__5 (
             \$dummy [714]), .ordered_filter_data_1__4 (\$dummy [715]), .ordered_filter_data_1__3 (
             \$dummy [716]), .ordered_filter_data_1__2 (\$dummy [717]), .ordered_filter_data_1__1 (
             \$dummy [718]), .ordered_filter_data_1__0 (\$dummy [719]), .ordered_filter_data_2__31 (
             \$dummy [720]), .ordered_filter_data_2__30 (\$dummy [721]), .ordered_filter_data_2__29 (
             \$dummy [722]), .ordered_filter_data_2__28 (\$dummy [723]), .ordered_filter_data_2__27 (
             \$dummy [724]), .ordered_filter_data_2__26 (\$dummy [725]), .ordered_filter_data_2__25 (
             \$dummy [726]), .ordered_filter_data_2__24 (\$dummy [727]), .ordered_filter_data_2__23 (
             \$dummy [728]), .ordered_filter_data_2__22 (\$dummy [729]), .ordered_filter_data_2__21 (
             \$dummy [730]), .ordered_filter_data_2__20 (\$dummy [731]), .ordered_filter_data_2__19 (
             \$dummy [732]), .ordered_filter_data_2__18 (\$dummy [733]), .ordered_filter_data_2__17 (
             \$dummy [734]), .ordered_filter_data_2__16 (\$dummy [735]), .ordered_filter_data_2__15 (
             \$dummy [736]), .ordered_filter_data_2__14 (\$dummy [737]), .ordered_filter_data_2__13 (
             \$dummy [738]), .ordered_filter_data_2__12 (\$dummy [739]), .ordered_filter_data_2__11 (
             \$dummy [740]), .ordered_filter_data_2__10 (\$dummy [741]), .ordered_filter_data_2__9 (
             \$dummy [742]), .ordered_filter_data_2__8 (\$dummy [743]), .ordered_filter_data_2__7 (
             \$dummy [744]), .ordered_filter_data_2__6 (\$dummy [745]), .ordered_filter_data_2__5 (
             \$dummy [746]), .ordered_filter_data_2__4 (\$dummy [747]), .ordered_filter_data_2__3 (
             \$dummy [748]), .ordered_filter_data_2__2 (\$dummy [749]), .ordered_filter_data_2__1 (
             \$dummy [750]), .ordered_filter_data_2__0 (\$dummy [751]), .ordered_filter_data_3__31 (
             \$dummy [752]), .ordered_filter_data_3__30 (\$dummy [753]), .ordered_filter_data_3__29 (
             \$dummy [754]), .ordered_filter_data_3__28 (\$dummy [755]), .ordered_filter_data_3__27 (
             \$dummy [756]), .ordered_filter_data_3__26 (\$dummy [757]), .ordered_filter_data_3__25 (
             \$dummy [758]), .ordered_filter_data_3__24 (\$dummy [759]), .ordered_filter_data_3__23 (
             \$dummy [760]), .ordered_filter_data_3__22 (\$dummy [761]), .ordered_filter_data_3__21 (
             \$dummy [762]), .ordered_filter_data_3__20 (\$dummy [763]), .ordered_filter_data_3__19 (
             \$dummy [764]), .ordered_filter_data_3__18 (\$dummy [765]), .ordered_filter_data_3__17 (
             \$dummy [766]), .ordered_filter_data_3__16 (\$dummy [767]), .ordered_filter_data_3__15 (
             ordered_filter_data_3__15), .ordered_filter_data_3__14 (
             ordered_filter_data_3__14), .ordered_filter_data_3__13 (
             ordered_filter_data_3__13), .ordered_filter_data_3__12 (
             ordered_filter_data_3__12), .ordered_filter_data_3__11 (
             ordered_filter_data_3__11), .ordered_filter_data_3__10 (
             ordered_filter_data_3__10), .ordered_filter_data_3__9 (
             ordered_filter_data_3__9), .ordered_filter_data_3__8 (
             ordered_filter_data_3__8), .ordered_filter_data_3__7 (
             ordered_filter_data_3__7), .ordered_filter_data_3__6 (
             ordered_filter_data_3__6), .ordered_filter_data_3__5 (
             ordered_filter_data_3__5), .ordered_filter_data_3__4 (
             ordered_filter_data_3__4), .ordered_filter_data_3__3 (
             ordered_filter_data_3__3), .ordered_filter_data_3__2 (
             ordered_filter_data_3__2), .ordered_filter_data_3__1 (
             ordered_filter_data_3__1), .ordered_filter_data_3__0 (
             ordered_filter_data_3__0), .ordered_filter_data_4__31 (
             \$dummy [768]), .ordered_filter_data_4__30 (\$dummy [769]), .ordered_filter_data_4__29 (
             \$dummy [770]), .ordered_filter_data_4__28 (\$dummy [771]), .ordered_filter_data_4__27 (
             \$dummy [772]), .ordered_filter_data_4__26 (\$dummy [773]), .ordered_filter_data_4__25 (
             \$dummy [774]), .ordered_filter_data_4__24 (\$dummy [775]), .ordered_filter_data_4__23 (
             \$dummy [776]), .ordered_filter_data_4__22 (\$dummy [777]), .ordered_filter_data_4__21 (
             \$dummy [778]), .ordered_filter_data_4__20 (\$dummy [779]), .ordered_filter_data_4__19 (
             \$dummy [780]), .ordered_filter_data_4__18 (\$dummy [781]), .ordered_filter_data_4__17 (
             \$dummy [782]), .ordered_filter_data_4__16 (\$dummy [783]), .ordered_filter_data_4__15 (
             ordered_filter_data_4__15), .ordered_filter_data_4__14 (
             ordered_filter_data_4__14), .ordered_filter_data_4__13 (
             ordered_filter_data_4__13), .ordered_filter_data_4__12 (
             ordered_filter_data_4__12), .ordered_filter_data_4__11 (
             ordered_filter_data_4__11), .ordered_filter_data_4__10 (
             ordered_filter_data_4__10), .ordered_filter_data_4__9 (
             ordered_filter_data_4__9), .ordered_filter_data_4__8 (
             ordered_filter_data_4__8), .ordered_filter_data_4__7 (
             ordered_filter_data_4__7), .ordered_filter_data_4__6 (
             ordered_filter_data_4__6), .ordered_filter_data_4__5 (
             ordered_filter_data_4__5), .ordered_filter_data_4__4 (
             ordered_filter_data_4__4), .ordered_filter_data_4__3 (
             ordered_filter_data_4__3), .ordered_filter_data_4__2 (
             ordered_filter_data_4__2), .ordered_filter_data_4__1 (
             ordered_filter_data_4__1), .ordered_filter_data_4__0 (
             ordered_filter_data_4__0), .ordered_filter_data_5__31 (
             \$dummy [784]), .ordered_filter_data_5__30 (\$dummy [785]), .ordered_filter_data_5__29 (
             \$dummy [786]), .ordered_filter_data_5__28 (\$dummy [787]), .ordered_filter_data_5__27 (
             \$dummy [788]), .ordered_filter_data_5__26 (\$dummy [789]), .ordered_filter_data_5__25 (
             \$dummy [790]), .ordered_filter_data_5__24 (\$dummy [791]), .ordered_filter_data_5__23 (
             \$dummy [792]), .ordered_filter_data_5__22 (\$dummy [793]), .ordered_filter_data_5__21 (
             \$dummy [794]), .ordered_filter_data_5__20 (\$dummy [795]), .ordered_filter_data_5__19 (
             \$dummy [796]), .ordered_filter_data_5__18 (\$dummy [797]), .ordered_filter_data_5__17 (
             \$dummy [798]), .ordered_filter_data_5__16 (\$dummy [799]), .ordered_filter_data_5__15 (
             ordered_filter_data_5__15), .ordered_filter_data_5__14 (
             ordered_filter_data_5__14), .ordered_filter_data_5__13 (
             ordered_filter_data_5__13), .ordered_filter_data_5__12 (
             ordered_filter_data_5__12), .ordered_filter_data_5__11 (
             ordered_filter_data_5__11), .ordered_filter_data_5__10 (
             ordered_filter_data_5__10), .ordered_filter_data_5__9 (
             ordered_filter_data_5__9), .ordered_filter_data_5__8 (
             ordered_filter_data_5__8), .ordered_filter_data_5__7 (
             ordered_filter_data_5__7), .ordered_filter_data_5__6 (
             ordered_filter_data_5__6), .ordered_filter_data_5__5 (
             ordered_filter_data_5__5), .ordered_filter_data_5__4 (
             ordered_filter_data_5__4), .ordered_filter_data_5__3 (
             ordered_filter_data_5__3), .ordered_filter_data_5__2 (
             ordered_filter_data_5__2), .ordered_filter_data_5__1 (
             ordered_filter_data_5__1), .ordered_filter_data_5__0 (
             ordered_filter_data_5__0), .ordered_filter_data_6__31 (
             \$dummy [800]), .ordered_filter_data_6__30 (\$dummy [801]), .ordered_filter_data_6__29 (
             \$dummy [802]), .ordered_filter_data_6__28 (\$dummy [803]), .ordered_filter_data_6__27 (
             \$dummy [804]), .ordered_filter_data_6__26 (\$dummy [805]), .ordered_filter_data_6__25 (
             \$dummy [806]), .ordered_filter_data_6__24 (\$dummy [807]), .ordered_filter_data_6__23 (
             \$dummy [808]), .ordered_filter_data_6__22 (\$dummy [809]), .ordered_filter_data_6__21 (
             \$dummy [810]), .ordered_filter_data_6__20 (\$dummy [811]), .ordered_filter_data_6__19 (
             \$dummy [812]), .ordered_filter_data_6__18 (\$dummy [813]), .ordered_filter_data_6__17 (
             \$dummy [814]), .ordered_filter_data_6__16 (\$dummy [815]), .ordered_filter_data_6__15 (
             ordered_filter_data_6__15), .ordered_filter_data_6__14 (
             ordered_filter_data_6__14), .ordered_filter_data_6__13 (
             ordered_filter_data_6__13), .ordered_filter_data_6__12 (
             ordered_filter_data_6__12), .ordered_filter_data_6__11 (
             ordered_filter_data_6__11), .ordered_filter_data_6__10 (
             ordered_filter_data_6__10), .ordered_filter_data_6__9 (
             ordered_filter_data_6__9), .ordered_filter_data_6__8 (
             ordered_filter_data_6__8), .ordered_filter_data_6__7 (
             ordered_filter_data_6__7), .ordered_filter_data_6__6 (
             ordered_filter_data_6__6), .ordered_filter_data_6__5 (
             ordered_filter_data_6__5), .ordered_filter_data_6__4 (
             ordered_filter_data_6__4), .ordered_filter_data_6__3 (
             ordered_filter_data_6__3), .ordered_filter_data_6__2 (
             ordered_filter_data_6__2), .ordered_filter_data_6__1 (
             ordered_filter_data_6__1), .ordered_filter_data_6__0 (
             ordered_filter_data_6__0), .ordered_filter_data_7__31 (
             \$dummy [816]), .ordered_filter_data_7__30 (\$dummy [817]), .ordered_filter_data_7__29 (
             \$dummy [818]), .ordered_filter_data_7__28 (\$dummy [819]), .ordered_filter_data_7__27 (
             \$dummy [820]), .ordered_filter_data_7__26 (\$dummy [821]), .ordered_filter_data_7__25 (
             \$dummy [822]), .ordered_filter_data_7__24 (\$dummy [823]), .ordered_filter_data_7__23 (
             \$dummy [824]), .ordered_filter_data_7__22 (\$dummy [825]), .ordered_filter_data_7__21 (
             \$dummy [826]), .ordered_filter_data_7__20 (\$dummy [827]), .ordered_filter_data_7__19 (
             \$dummy [828]), .ordered_filter_data_7__18 (\$dummy [829]), .ordered_filter_data_7__17 (
             \$dummy [830]), .ordered_filter_data_7__16 (\$dummy [831]), .ordered_filter_data_7__15 (
             ordered_filter_data_7__15), .ordered_filter_data_7__14 (
             ordered_filter_data_7__14), .ordered_filter_data_7__13 (
             ordered_filter_data_7__13), .ordered_filter_data_7__12 (
             ordered_filter_data_7__12), .ordered_filter_data_7__11 (
             ordered_filter_data_7__11), .ordered_filter_data_7__10 (
             ordered_filter_data_7__10), .ordered_filter_data_7__9 (
             ordered_filter_data_7__9), .ordered_filter_data_7__8 (
             ordered_filter_data_7__8), .ordered_filter_data_7__7 (
             ordered_filter_data_7__7), .ordered_filter_data_7__6 (
             ordered_filter_data_7__6), .ordered_filter_data_7__5 (
             ordered_filter_data_7__5), .ordered_filter_data_7__4 (
             ordered_filter_data_7__4), .ordered_filter_data_7__3 (
             ordered_filter_data_7__3), .ordered_filter_data_7__2 (
             ordered_filter_data_7__2), .ordered_filter_data_7__1 (
             ordered_filter_data_7__1), .ordered_filter_data_7__0 (
             ordered_filter_data_7__0), .ordered_filter_data_8__31 (
             \$dummy [832]), .ordered_filter_data_8__30 (\$dummy [833]), .ordered_filter_data_8__29 (
             \$dummy [834]), .ordered_filter_data_8__28 (\$dummy [835]), .ordered_filter_data_8__27 (
             \$dummy [836]), .ordered_filter_data_8__26 (\$dummy [837]), .ordered_filter_data_8__25 (
             \$dummy [838]), .ordered_filter_data_8__24 (\$dummy [839]), .ordered_filter_data_8__23 (
             \$dummy [840]), .ordered_filter_data_8__22 (\$dummy [841]), .ordered_filter_data_8__21 (
             \$dummy [842]), .ordered_filter_data_8__20 (\$dummy [843]), .ordered_filter_data_8__19 (
             \$dummy [844]), .ordered_filter_data_8__18 (\$dummy [845]), .ordered_filter_data_8__17 (
             \$dummy [846]), .ordered_filter_data_8__16 (\$dummy [847]), .ordered_filter_data_8__15 (
             ordered_filter_data_8__15), .ordered_filter_data_8__14 (
             ordered_filter_data_8__14), .ordered_filter_data_8__13 (
             ordered_filter_data_8__13), .ordered_filter_data_8__12 (
             ordered_filter_data_8__12), .ordered_filter_data_8__11 (
             ordered_filter_data_8__11), .ordered_filter_data_8__10 (
             ordered_filter_data_8__10), .ordered_filter_data_8__9 (
             ordered_filter_data_8__9), .ordered_filter_data_8__8 (
             ordered_filter_data_8__8), .ordered_filter_data_8__7 (
             ordered_filter_data_8__7), .ordered_filter_data_8__6 (
             ordered_filter_data_8__6), .ordered_filter_data_8__5 (
             ordered_filter_data_8__5), .ordered_filter_data_8__4 (
             ordered_filter_data_8__4), .ordered_filter_data_8__3 (
             ordered_filter_data_8__3), .ordered_filter_data_8__2 (
             ordered_filter_data_8__2), .ordered_filter_data_8__1 (
             ordered_filter_data_8__1), .ordered_filter_data_8__0 (
             ordered_filter_data_8__0), .ordered_filter_data_9__31 (
             \$dummy [848]), .ordered_filter_data_9__30 (\$dummy [849]), .ordered_filter_data_9__29 (
             \$dummy [850]), .ordered_filter_data_9__28 (\$dummy [851]), .ordered_filter_data_9__27 (
             \$dummy [852]), .ordered_filter_data_9__26 (\$dummy [853]), .ordered_filter_data_9__25 (
             \$dummy [854]), .ordered_filter_data_9__24 (\$dummy [855]), .ordered_filter_data_9__23 (
             \$dummy [856]), .ordered_filter_data_9__22 (\$dummy [857]), .ordered_filter_data_9__21 (
             \$dummy [858]), .ordered_filter_data_9__20 (\$dummy [859]), .ordered_filter_data_9__19 (
             \$dummy [860]), .ordered_filter_data_9__18 (\$dummy [861]), .ordered_filter_data_9__17 (
             \$dummy [862]), .ordered_filter_data_9__16 (\$dummy [863]), .ordered_filter_data_9__15 (
             ordered_filter_data_9__15), .ordered_filter_data_9__14 (
             ordered_filter_data_9__14), .ordered_filter_data_9__13 (
             ordered_filter_data_9__13), .ordered_filter_data_9__12 (
             ordered_filter_data_9__12), .ordered_filter_data_9__11 (
             ordered_filter_data_9__11), .ordered_filter_data_9__10 (
             ordered_filter_data_9__10), .ordered_filter_data_9__9 (
             ordered_filter_data_9__9), .ordered_filter_data_9__8 (
             ordered_filter_data_9__8), .ordered_filter_data_9__7 (
             ordered_filter_data_9__7), .ordered_filter_data_9__6 (
             ordered_filter_data_9__6), .ordered_filter_data_9__5 (
             ordered_filter_data_9__5), .ordered_filter_data_9__4 (
             ordered_filter_data_9__4), .ordered_filter_data_9__3 (
             ordered_filter_data_9__3), .ordered_filter_data_9__2 (
             ordered_filter_data_9__2), .ordered_filter_data_9__1 (
             ordered_filter_data_9__1), .ordered_filter_data_9__0 (
             ordered_filter_data_9__0), .ordered_filter_data_10__31 (
             \$dummy [864]), .ordered_filter_data_10__30 (\$dummy [865]), .ordered_filter_data_10__29 (
             \$dummy [866]), .ordered_filter_data_10__28 (\$dummy [867]), .ordered_filter_data_10__27 (
             \$dummy [868]), .ordered_filter_data_10__26 (\$dummy [869]), .ordered_filter_data_10__25 (
             \$dummy [870]), .ordered_filter_data_10__24 (\$dummy [871]), .ordered_filter_data_10__23 (
             \$dummy [872]), .ordered_filter_data_10__22 (\$dummy [873]), .ordered_filter_data_10__21 (
             \$dummy [874]), .ordered_filter_data_10__20 (\$dummy [875]), .ordered_filter_data_10__19 (
             \$dummy [876]), .ordered_filter_data_10__18 (\$dummy [877]), .ordered_filter_data_10__17 (
             \$dummy [878]), .ordered_filter_data_10__16 (\$dummy [879]), .ordered_filter_data_10__15 (
             ordered_filter_data_10__15), .ordered_filter_data_10__14 (
             ordered_filter_data_10__14), .ordered_filter_data_10__13 (
             ordered_filter_data_10__13), .ordered_filter_data_10__12 (
             ordered_filter_data_10__12), .ordered_filter_data_10__11 (
             ordered_filter_data_10__11), .ordered_filter_data_10__10 (
             ordered_filter_data_10__10), .ordered_filter_data_10__9 (
             ordered_filter_data_10__9), .ordered_filter_data_10__8 (
             ordered_filter_data_10__8), .ordered_filter_data_10__7 (
             ordered_filter_data_10__7), .ordered_filter_data_10__6 (
             ordered_filter_data_10__6), .ordered_filter_data_10__5 (
             ordered_filter_data_10__5), .ordered_filter_data_10__4 (
             ordered_filter_data_10__4), .ordered_filter_data_10__3 (
             ordered_filter_data_10__3), .ordered_filter_data_10__2 (
             ordered_filter_data_10__2), .ordered_filter_data_10__1 (
             ordered_filter_data_10__1), .ordered_filter_data_10__0 (
             ordered_filter_data_10__0), .ordered_filter_data_11__31 (
             \$dummy [880]), .ordered_filter_data_11__30 (\$dummy [881]), .ordered_filter_data_11__29 (
             \$dummy [882]), .ordered_filter_data_11__28 (\$dummy [883]), .ordered_filter_data_11__27 (
             \$dummy [884]), .ordered_filter_data_11__26 (\$dummy [885]), .ordered_filter_data_11__25 (
             \$dummy [886]), .ordered_filter_data_11__24 (\$dummy [887]), .ordered_filter_data_11__23 (
             \$dummy [888]), .ordered_filter_data_11__22 (\$dummy [889]), .ordered_filter_data_11__21 (
             \$dummy [890]), .ordered_filter_data_11__20 (\$dummy [891]), .ordered_filter_data_11__19 (
             \$dummy [892]), .ordered_filter_data_11__18 (\$dummy [893]), .ordered_filter_data_11__17 (
             \$dummy [894]), .ordered_filter_data_11__16 (\$dummy [895]), .ordered_filter_data_11__15 (
             ordered_filter_data_11__15), .ordered_filter_data_11__14 (
             ordered_filter_data_11__14), .ordered_filter_data_11__13 (
             ordered_filter_data_11__13), .ordered_filter_data_11__12 (
             ordered_filter_data_11__12), .ordered_filter_data_11__11 (
             ordered_filter_data_11__11), .ordered_filter_data_11__10 (
             ordered_filter_data_11__10), .ordered_filter_data_11__9 (
             ordered_filter_data_11__9), .ordered_filter_data_11__8 (
             ordered_filter_data_11__8), .ordered_filter_data_11__7 (
             ordered_filter_data_11__7), .ordered_filter_data_11__6 (
             ordered_filter_data_11__6), .ordered_filter_data_11__5 (
             ordered_filter_data_11__5), .ordered_filter_data_11__4 (
             ordered_filter_data_11__4), .ordered_filter_data_11__3 (
             ordered_filter_data_11__3), .ordered_filter_data_11__2 (
             ordered_filter_data_11__2), .ordered_filter_data_11__1 (
             ordered_filter_data_11__1), .ordered_filter_data_11__0 (
             ordered_filter_data_11__0), .ordered_filter_data_12__31 (
             \$dummy [896]), .ordered_filter_data_12__30 (\$dummy [897]), .ordered_filter_data_12__29 (
             \$dummy [898]), .ordered_filter_data_12__28 (\$dummy [899]), .ordered_filter_data_12__27 (
             \$dummy [900]), .ordered_filter_data_12__26 (\$dummy [901]), .ordered_filter_data_12__25 (
             \$dummy [902]), .ordered_filter_data_12__24 (\$dummy [903]), .ordered_filter_data_12__23 (
             \$dummy [904]), .ordered_filter_data_12__22 (\$dummy [905]), .ordered_filter_data_12__21 (
             \$dummy [906]), .ordered_filter_data_12__20 (\$dummy [907]), .ordered_filter_data_12__19 (
             \$dummy [908]), .ordered_filter_data_12__18 (\$dummy [909]), .ordered_filter_data_12__17 (
             \$dummy [910]), .ordered_filter_data_12__16 (\$dummy [911]), .ordered_filter_data_12__15 (
             ordered_filter_data_12__15), .ordered_filter_data_12__14 (
             ordered_filter_data_12__14), .ordered_filter_data_12__13 (
             ordered_filter_data_12__13), .ordered_filter_data_12__12 (
             ordered_filter_data_12__12), .ordered_filter_data_12__11 (
             ordered_filter_data_12__11), .ordered_filter_data_12__10 (
             ordered_filter_data_12__10), .ordered_filter_data_12__9 (
             ordered_filter_data_12__9), .ordered_filter_data_12__8 (
             ordered_filter_data_12__8), .ordered_filter_data_12__7 (
             ordered_filter_data_12__7), .ordered_filter_data_12__6 (
             ordered_filter_data_12__6), .ordered_filter_data_12__5 (
             ordered_filter_data_12__5), .ordered_filter_data_12__4 (
             ordered_filter_data_12__4), .ordered_filter_data_12__3 (
             ordered_filter_data_12__3), .ordered_filter_data_12__2 (
             ordered_filter_data_12__2), .ordered_filter_data_12__1 (
             ordered_filter_data_12__1), .ordered_filter_data_12__0 (
             ordered_filter_data_12__0), .ordered_filter_data_13__31 (
             \$dummy [912]), .ordered_filter_data_13__30 (\$dummy [913]), .ordered_filter_data_13__29 (
             \$dummy [914]), .ordered_filter_data_13__28 (\$dummy [915]), .ordered_filter_data_13__27 (
             \$dummy [916]), .ordered_filter_data_13__26 (\$dummy [917]), .ordered_filter_data_13__25 (
             \$dummy [918]), .ordered_filter_data_13__24 (\$dummy [919]), .ordered_filter_data_13__23 (
             \$dummy [920]), .ordered_filter_data_13__22 (\$dummy [921]), .ordered_filter_data_13__21 (
             \$dummy [922]), .ordered_filter_data_13__20 (\$dummy [923]), .ordered_filter_data_13__19 (
             \$dummy [924]), .ordered_filter_data_13__18 (\$dummy [925]), .ordered_filter_data_13__17 (
             \$dummy [926]), .ordered_filter_data_13__16 (\$dummy [927]), .ordered_filter_data_13__15 (
             ordered_filter_data_13__15), .ordered_filter_data_13__14 (
             ordered_filter_data_13__14), .ordered_filter_data_13__13 (
             ordered_filter_data_13__13), .ordered_filter_data_13__12 (
             ordered_filter_data_13__12), .ordered_filter_data_13__11 (
             ordered_filter_data_13__11), .ordered_filter_data_13__10 (
             ordered_filter_data_13__10), .ordered_filter_data_13__9 (
             ordered_filter_data_13__9), .ordered_filter_data_13__8 (
             ordered_filter_data_13__8), .ordered_filter_data_13__7 (
             ordered_filter_data_13__7), .ordered_filter_data_13__6 (
             ordered_filter_data_13__6), .ordered_filter_data_13__5 (
             ordered_filter_data_13__5), .ordered_filter_data_13__4 (
             ordered_filter_data_13__4), .ordered_filter_data_13__3 (
             ordered_filter_data_13__3), .ordered_filter_data_13__2 (
             ordered_filter_data_13__2), .ordered_filter_data_13__1 (
             ordered_filter_data_13__1), .ordered_filter_data_13__0 (
             ordered_filter_data_13__0), .ordered_filter_data_14__31 (
             \$dummy [928]), .ordered_filter_data_14__30 (\$dummy [929]), .ordered_filter_data_14__29 (
             \$dummy [930]), .ordered_filter_data_14__28 (\$dummy [931]), .ordered_filter_data_14__27 (
             \$dummy [932]), .ordered_filter_data_14__26 (\$dummy [933]), .ordered_filter_data_14__25 (
             \$dummy [934]), .ordered_filter_data_14__24 (\$dummy [935]), .ordered_filter_data_14__23 (
             \$dummy [936]), .ordered_filter_data_14__22 (\$dummy [937]), .ordered_filter_data_14__21 (
             \$dummy [938]), .ordered_filter_data_14__20 (\$dummy [939]), .ordered_filter_data_14__19 (
             \$dummy [940]), .ordered_filter_data_14__18 (\$dummy [941]), .ordered_filter_data_14__17 (
             \$dummy [942]), .ordered_filter_data_14__16 (\$dummy [943]), .ordered_filter_data_14__15 (
             ordered_filter_data_14__15), .ordered_filter_data_14__14 (
             ordered_filter_data_14__14), .ordered_filter_data_14__13 (
             ordered_filter_data_14__13), .ordered_filter_data_14__12 (
             ordered_filter_data_14__12), .ordered_filter_data_14__11 (
             ordered_filter_data_14__11), .ordered_filter_data_14__10 (
             ordered_filter_data_14__10), .ordered_filter_data_14__9 (
             ordered_filter_data_14__9), .ordered_filter_data_14__8 (
             ordered_filter_data_14__8), .ordered_filter_data_14__7 (
             ordered_filter_data_14__7), .ordered_filter_data_14__6 (
             ordered_filter_data_14__6), .ordered_filter_data_14__5 (
             ordered_filter_data_14__5), .ordered_filter_data_14__4 (
             ordered_filter_data_14__4), .ordered_filter_data_14__3 (
             ordered_filter_data_14__3), .ordered_filter_data_14__2 (
             ordered_filter_data_14__2), .ordered_filter_data_14__1 (
             ordered_filter_data_14__1), .ordered_filter_data_14__0 (
             ordered_filter_data_14__0), .ordered_filter_data_15__31 (
             \$dummy [944]), .ordered_filter_data_15__30 (\$dummy [945]), .ordered_filter_data_15__29 (
             \$dummy [946]), .ordered_filter_data_15__28 (\$dummy [947]), .ordered_filter_data_15__27 (
             \$dummy [948]), .ordered_filter_data_15__26 (\$dummy [949]), .ordered_filter_data_15__25 (
             \$dummy [950]), .ordered_filter_data_15__24 (\$dummy [951]), .ordered_filter_data_15__23 (
             \$dummy [952]), .ordered_filter_data_15__22 (\$dummy [953]), .ordered_filter_data_15__21 (
             \$dummy [954]), .ordered_filter_data_15__20 (\$dummy [955]), .ordered_filter_data_15__19 (
             \$dummy [956]), .ordered_filter_data_15__18 (\$dummy [957]), .ordered_filter_data_15__17 (
             \$dummy [958]), .ordered_filter_data_15__16 (\$dummy [959]), .ordered_filter_data_15__15 (
             ordered_filter_data_15__15), .ordered_filter_data_15__14 (
             ordered_filter_data_15__14), .ordered_filter_data_15__13 (
             ordered_filter_data_15__13), .ordered_filter_data_15__12 (
             ordered_filter_data_15__12), .ordered_filter_data_15__11 (
             ordered_filter_data_15__11), .ordered_filter_data_15__10 (
             ordered_filter_data_15__10), .ordered_filter_data_15__9 (
             ordered_filter_data_15__9), .ordered_filter_data_15__8 (
             ordered_filter_data_15__8), .ordered_filter_data_15__7 (
             ordered_filter_data_15__7), .ordered_filter_data_15__6 (
             ordered_filter_data_15__6), .ordered_filter_data_15__5 (
             ordered_filter_data_15__5), .ordered_filter_data_15__4 (
             ordered_filter_data_15__4), .ordered_filter_data_15__3 (
             ordered_filter_data_15__3), .ordered_filter_data_15__2 (
             ordered_filter_data_15__2), .ordered_filter_data_15__1 (
             ordered_filter_data_15__1), .ordered_filter_data_15__0 (
             ordered_filter_data_15__0), .ordered_filter_data_16__31 (
             \$dummy [960]), .ordered_filter_data_16__30 (\$dummy [961]), .ordered_filter_data_16__29 (
             \$dummy [962]), .ordered_filter_data_16__28 (\$dummy [963]), .ordered_filter_data_16__27 (
             \$dummy [964]), .ordered_filter_data_16__26 (\$dummy [965]), .ordered_filter_data_16__25 (
             \$dummy [966]), .ordered_filter_data_16__24 (\$dummy [967]), .ordered_filter_data_16__23 (
             \$dummy [968]), .ordered_filter_data_16__22 (\$dummy [969]), .ordered_filter_data_16__21 (
             \$dummy [970]), .ordered_filter_data_16__20 (\$dummy [971]), .ordered_filter_data_16__19 (
             \$dummy [972]), .ordered_filter_data_16__18 (\$dummy [973]), .ordered_filter_data_16__17 (
             \$dummy [974]), .ordered_filter_data_16__16 (\$dummy [975]), .ordered_filter_data_16__15 (
             ordered_filter_data_16__15), .ordered_filter_data_16__14 (
             ordered_filter_data_16__14), .ordered_filter_data_16__13 (
             ordered_filter_data_16__13), .ordered_filter_data_16__12 (
             ordered_filter_data_16__12), .ordered_filter_data_16__11 (
             ordered_filter_data_16__11), .ordered_filter_data_16__10 (
             ordered_filter_data_16__10), .ordered_filter_data_16__9 (
             ordered_filter_data_16__9), .ordered_filter_data_16__8 (
             ordered_filter_data_16__8), .ordered_filter_data_16__7 (
             ordered_filter_data_16__7), .ordered_filter_data_16__6 (
             ordered_filter_data_16__6), .ordered_filter_data_16__5 (
             ordered_filter_data_16__5), .ordered_filter_data_16__4 (
             ordered_filter_data_16__4), .ordered_filter_data_16__3 (
             ordered_filter_data_16__3), .ordered_filter_data_16__2 (
             ordered_filter_data_16__2), .ordered_filter_data_16__1 (
             ordered_filter_data_16__1), .ordered_filter_data_16__0 (
             ordered_filter_data_16__0), .ordered_filter_data_17__31 (
             \$dummy [976]), .ordered_filter_data_17__30 (\$dummy [977]), .ordered_filter_data_17__29 (
             \$dummy [978]), .ordered_filter_data_17__28 (\$dummy [979]), .ordered_filter_data_17__27 (
             \$dummy [980]), .ordered_filter_data_17__26 (\$dummy [981]), .ordered_filter_data_17__25 (
             \$dummy [982]), .ordered_filter_data_17__24 (\$dummy [983]), .ordered_filter_data_17__23 (
             \$dummy [984]), .ordered_filter_data_17__22 (\$dummy [985]), .ordered_filter_data_17__21 (
             \$dummy [986]), .ordered_filter_data_17__20 (\$dummy [987]), .ordered_filter_data_17__19 (
             \$dummy [988]), .ordered_filter_data_17__18 (\$dummy [989]), .ordered_filter_data_17__17 (
             \$dummy [990]), .ordered_filter_data_17__16 (\$dummy [991]), .ordered_filter_data_17__15 (
             ordered_filter_data_17__15), .ordered_filter_data_17__14 (
             ordered_filter_data_17__14), .ordered_filter_data_17__13 (
             ordered_filter_data_17__13), .ordered_filter_data_17__12 (
             ordered_filter_data_17__12), .ordered_filter_data_17__11 (
             ordered_filter_data_17__11), .ordered_filter_data_17__10 (
             ordered_filter_data_17__10), .ordered_filter_data_17__9 (
             ordered_filter_data_17__9), .ordered_filter_data_17__8 (
             ordered_filter_data_17__8), .ordered_filter_data_17__7 (
             ordered_filter_data_17__7), .ordered_filter_data_17__6 (
             ordered_filter_data_17__6), .ordered_filter_data_17__5 (
             ordered_filter_data_17__5), .ordered_filter_data_17__4 (
             ordered_filter_data_17__4), .ordered_filter_data_17__3 (
             ordered_filter_data_17__3), .ordered_filter_data_17__2 (
             ordered_filter_data_17__2), .ordered_filter_data_17__1 (
             ordered_filter_data_17__1), .ordered_filter_data_17__0 (
             ordered_filter_data_17__0), .ordered_filter_data_18__31 (
             \$dummy [992]), .ordered_filter_data_18__30 (\$dummy [993]), .ordered_filter_data_18__29 (
             \$dummy [994]), .ordered_filter_data_18__28 (\$dummy [995]), .ordered_filter_data_18__27 (
             \$dummy [996]), .ordered_filter_data_18__26 (\$dummy [997]), .ordered_filter_data_18__25 (
             \$dummy [998]), .ordered_filter_data_18__24 (\$dummy [999]), .ordered_filter_data_18__23 (
             \$dummy [1000]), .ordered_filter_data_18__22 (\$dummy [1001]), .ordered_filter_data_18__21 (
             \$dummy [1002]), .ordered_filter_data_18__20 (\$dummy [1003]), .ordered_filter_data_18__19 (
             \$dummy [1004]), .ordered_filter_data_18__18 (\$dummy [1005]), .ordered_filter_data_18__17 (
             \$dummy [1006]), .ordered_filter_data_18__16 (\$dummy [1007]), .ordered_filter_data_18__15 (
             \$dummy [1008]), .ordered_filter_data_18__14 (\$dummy [1009]), .ordered_filter_data_18__13 (
             \$dummy [1010]), .ordered_filter_data_18__12 (\$dummy [1011]), .ordered_filter_data_18__11 (
             \$dummy [1012]), .ordered_filter_data_18__10 (\$dummy [1013]), .ordered_filter_data_18__9 (
             \$dummy [1014]), .ordered_filter_data_18__8 (\$dummy [1015]), .ordered_filter_data_18__7 (
             \$dummy [1016]), .ordered_filter_data_18__6 (\$dummy [1017]), .ordered_filter_data_18__5 (
             \$dummy [1018]), .ordered_filter_data_18__4 (\$dummy [1019]), .ordered_filter_data_18__3 (
             \$dummy [1020]), .ordered_filter_data_18__2 (\$dummy [1021]), .ordered_filter_data_18__1 (
             \$dummy [1022]), .ordered_filter_data_18__0 (\$dummy [1023]), .ordered_filter_data_19__31 (
             \$dummy [1024]), .ordered_filter_data_19__30 (\$dummy [1025]), .ordered_filter_data_19__29 (
             \$dummy [1026]), .ordered_filter_data_19__28 (\$dummy [1027]), .ordered_filter_data_19__27 (
             \$dummy [1028]), .ordered_filter_data_19__26 (\$dummy [1029]), .ordered_filter_data_19__25 (
             \$dummy [1030]), .ordered_filter_data_19__24 (\$dummy [1031]), .ordered_filter_data_19__23 (
             \$dummy [1032]), .ordered_filter_data_19__22 (\$dummy [1033]), .ordered_filter_data_19__21 (
             \$dummy [1034]), .ordered_filter_data_19__20 (\$dummy [1035]), .ordered_filter_data_19__19 (
             \$dummy [1036]), .ordered_filter_data_19__18 (\$dummy [1037]), .ordered_filter_data_19__17 (
             \$dummy [1038]), .ordered_filter_data_19__16 (\$dummy [1039]), .ordered_filter_data_19__15 (
             \$dummy [1040]), .ordered_filter_data_19__14 (\$dummy [1041]), .ordered_filter_data_19__13 (
             \$dummy [1042]), .ordered_filter_data_19__12 (\$dummy [1043]), .ordered_filter_data_19__11 (
             \$dummy [1044]), .ordered_filter_data_19__10 (\$dummy [1045]), .ordered_filter_data_19__9 (
             \$dummy [1046]), .ordered_filter_data_19__8 (\$dummy [1047]), .ordered_filter_data_19__7 (
             \$dummy [1048]), .ordered_filter_data_19__6 (\$dummy [1049]), .ordered_filter_data_19__5 (
             \$dummy [1050]), .ordered_filter_data_19__4 (\$dummy [1051]), .ordered_filter_data_19__3 (
             \$dummy [1052]), .ordered_filter_data_19__2 (\$dummy [1053]), .ordered_filter_data_19__1 (
             \$dummy [1054]), .ordered_filter_data_19__0 (\$dummy [1055]), .ordered_filter_data_20__31 (
             \$dummy [1056]), .ordered_filter_data_20__30 (\$dummy [1057]), .ordered_filter_data_20__29 (
             \$dummy [1058]), .ordered_filter_data_20__28 (\$dummy [1059]), .ordered_filter_data_20__27 (
             \$dummy [1060]), .ordered_filter_data_20__26 (\$dummy [1061]), .ordered_filter_data_20__25 (
             \$dummy [1062]), .ordered_filter_data_20__24 (\$dummy [1063]), .ordered_filter_data_20__23 (
             \$dummy [1064]), .ordered_filter_data_20__22 (\$dummy [1065]), .ordered_filter_data_20__21 (
             \$dummy [1066]), .ordered_filter_data_20__20 (\$dummy [1067]), .ordered_filter_data_20__19 (
             \$dummy [1068]), .ordered_filter_data_20__18 (\$dummy [1069]), .ordered_filter_data_20__17 (
             \$dummy [1070]), .ordered_filter_data_20__16 (\$dummy [1071]), .ordered_filter_data_20__15 (
             \$dummy [1072]), .ordered_filter_data_20__14 (\$dummy [1073]), .ordered_filter_data_20__13 (
             \$dummy [1074]), .ordered_filter_data_20__12 (\$dummy [1075]), .ordered_filter_data_20__11 (
             \$dummy [1076]), .ordered_filter_data_20__10 (\$dummy [1077]), .ordered_filter_data_20__9 (
             \$dummy [1078]), .ordered_filter_data_20__8 (\$dummy [1079]), .ordered_filter_data_20__7 (
             \$dummy [1080]), .ordered_filter_data_20__6 (\$dummy [1081]), .ordered_filter_data_20__5 (
             \$dummy [1082]), .ordered_filter_data_20__4 (\$dummy [1083]), .ordered_filter_data_20__3 (
             \$dummy [1084]), .ordered_filter_data_20__2 (\$dummy [1085]), .ordered_filter_data_20__1 (
             \$dummy [1086]), .ordered_filter_data_20__0 (\$dummy [1087]), .ordered_filter_data_21__31 (
             \$dummy [1088]), .ordered_filter_data_21__30 (\$dummy [1089]), .ordered_filter_data_21__29 (
             \$dummy [1090]), .ordered_filter_data_21__28 (\$dummy [1091]), .ordered_filter_data_21__27 (
             \$dummy [1092]), .ordered_filter_data_21__26 (\$dummy [1093]), .ordered_filter_data_21__25 (
             \$dummy [1094]), .ordered_filter_data_21__24 (\$dummy [1095]), .ordered_filter_data_21__23 (
             \$dummy [1096]), .ordered_filter_data_21__22 (\$dummy [1097]), .ordered_filter_data_21__21 (
             \$dummy [1098]), .ordered_filter_data_21__20 (\$dummy [1099]), .ordered_filter_data_21__19 (
             \$dummy [1100]), .ordered_filter_data_21__18 (\$dummy [1101]), .ordered_filter_data_21__17 (
             \$dummy [1102]), .ordered_filter_data_21__16 (\$dummy [1103]), .ordered_filter_data_21__15 (
             \$dummy [1104]), .ordered_filter_data_21__14 (\$dummy [1105]), .ordered_filter_data_21__13 (
             \$dummy [1106]), .ordered_filter_data_21__12 (\$dummy [1107]), .ordered_filter_data_21__11 (
             \$dummy [1108]), .ordered_filter_data_21__10 (\$dummy [1109]), .ordered_filter_data_21__9 (
             \$dummy [1110]), .ordered_filter_data_21__8 (\$dummy [1111]), .ordered_filter_data_21__7 (
             \$dummy [1112]), .ordered_filter_data_21__6 (\$dummy [1113]), .ordered_filter_data_21__5 (
             \$dummy [1114]), .ordered_filter_data_21__4 (\$dummy [1115]), .ordered_filter_data_21__3 (
             \$dummy [1116]), .ordered_filter_data_21__2 (\$dummy [1117]), .ordered_filter_data_21__1 (
             \$dummy [1118]), .ordered_filter_data_21__0 (\$dummy [1119]), .ordered_filter_data_22__31 (
             \$dummy [1120]), .ordered_filter_data_22__30 (\$dummy [1121]), .ordered_filter_data_22__29 (
             \$dummy [1122]), .ordered_filter_data_22__28 (\$dummy [1123]), .ordered_filter_data_22__27 (
             \$dummy [1124]), .ordered_filter_data_22__26 (\$dummy [1125]), .ordered_filter_data_22__25 (
             \$dummy [1126]), .ordered_filter_data_22__24 (\$dummy [1127]), .ordered_filter_data_22__23 (
             \$dummy [1128]), .ordered_filter_data_22__22 (\$dummy [1129]), .ordered_filter_data_22__21 (
             \$dummy [1130]), .ordered_filter_data_22__20 (\$dummy [1131]), .ordered_filter_data_22__19 (
             \$dummy [1132]), .ordered_filter_data_22__18 (\$dummy [1133]), .ordered_filter_data_22__17 (
             \$dummy [1134]), .ordered_filter_data_22__16 (\$dummy [1135]), .ordered_filter_data_22__15 (
             \$dummy [1136]), .ordered_filter_data_22__14 (\$dummy [1137]), .ordered_filter_data_22__13 (
             \$dummy [1138]), .ordered_filter_data_22__12 (\$dummy [1139]), .ordered_filter_data_22__11 (
             \$dummy [1140]), .ordered_filter_data_22__10 (\$dummy [1141]), .ordered_filter_data_22__9 (
             \$dummy [1142]), .ordered_filter_data_22__8 (\$dummy [1143]), .ordered_filter_data_22__7 (
             \$dummy [1144]), .ordered_filter_data_22__6 (\$dummy [1145]), .ordered_filter_data_22__5 (
             \$dummy [1146]), .ordered_filter_data_22__4 (\$dummy [1147]), .ordered_filter_data_22__3 (
             \$dummy [1148]), .ordered_filter_data_22__2 (\$dummy [1149]), .ordered_filter_data_22__1 (
             \$dummy [1150]), .ordered_filter_data_22__0 (\$dummy [1151]), .ordered_filter_data_23__31 (
             \$dummy [1152]), .ordered_filter_data_23__30 (\$dummy [1153]), .ordered_filter_data_23__29 (
             \$dummy [1154]), .ordered_filter_data_23__28 (\$dummy [1155]), .ordered_filter_data_23__27 (
             \$dummy [1156]), .ordered_filter_data_23__26 (\$dummy [1157]), .ordered_filter_data_23__25 (
             \$dummy [1158]), .ordered_filter_data_23__24 (\$dummy [1159]), .ordered_filter_data_23__23 (
             \$dummy [1160]), .ordered_filter_data_23__22 (\$dummy [1161]), .ordered_filter_data_23__21 (
             \$dummy [1162]), .ordered_filter_data_23__20 (\$dummy [1163]), .ordered_filter_data_23__19 (
             \$dummy [1164]), .ordered_filter_data_23__18 (\$dummy [1165]), .ordered_filter_data_23__17 (
             \$dummy [1166]), .ordered_filter_data_23__16 (\$dummy [1167]), .ordered_filter_data_23__15 (
             \$dummy [1168]), .ordered_filter_data_23__14 (\$dummy [1169]), .ordered_filter_data_23__13 (
             \$dummy [1170]), .ordered_filter_data_23__12 (\$dummy [1171]), .ordered_filter_data_23__11 (
             \$dummy [1172]), .ordered_filter_data_23__10 (\$dummy [1173]), .ordered_filter_data_23__9 (
             \$dummy [1174]), .ordered_filter_data_23__8 (\$dummy [1175]), .ordered_filter_data_23__7 (
             \$dummy [1176]), .ordered_filter_data_23__6 (\$dummy [1177]), .ordered_filter_data_23__5 (
             \$dummy [1178]), .ordered_filter_data_23__4 (\$dummy [1179]), .ordered_filter_data_23__3 (
             \$dummy [1180]), .ordered_filter_data_23__2 (\$dummy [1181]), .ordered_filter_data_23__1 (
             \$dummy [1182]), .ordered_filter_data_23__0 (\$dummy [1183]), .ordered_filter_data_24__31 (
             \$dummy [1184]), .ordered_filter_data_24__30 (\$dummy [1185]), .ordered_filter_data_24__29 (
             \$dummy [1186]), .ordered_filter_data_24__28 (\$dummy [1187]), .ordered_filter_data_24__27 (
             \$dummy [1188]), .ordered_filter_data_24__26 (\$dummy [1189]), .ordered_filter_data_24__25 (
             \$dummy [1190]), .ordered_filter_data_24__24 (\$dummy [1191]), .ordered_filter_data_24__23 (
             \$dummy [1192]), .ordered_filter_data_24__22 (\$dummy [1193]), .ordered_filter_data_24__21 (
             \$dummy [1194]), .ordered_filter_data_24__20 (\$dummy [1195]), .ordered_filter_data_24__19 (
             \$dummy [1196]), .ordered_filter_data_24__18 (\$dummy [1197]), .ordered_filter_data_24__17 (
             \$dummy [1198]), .ordered_filter_data_24__16 (\$dummy [1199]), .ordered_filter_data_24__15 (
             \$dummy [1200]), .ordered_filter_data_24__14 (\$dummy [1201]), .ordered_filter_data_24__13 (
             \$dummy [1202]), .ordered_filter_data_24__12 (\$dummy [1203]), .ordered_filter_data_24__11 (
             \$dummy [1204]), .ordered_filter_data_24__10 (\$dummy [1205]), .ordered_filter_data_24__9 (
             \$dummy [1206]), .ordered_filter_data_24__8 (\$dummy [1207]), .ordered_filter_data_24__7 (
             \$dummy [1208]), .ordered_filter_data_24__6 (\$dummy [1209]), .ordered_filter_data_24__5 (
             \$dummy [1210]), .ordered_filter_data_24__4 (\$dummy [1211]), .ordered_filter_data_24__3 (
             \$dummy [1212]), .ordered_filter_data_24__2 (\$dummy [1213]), .ordered_filter_data_24__1 (
             \$dummy [1214]), .ordered_filter_data_24__0 (\$dummy [1215])) ;
    MergeLayer merge_layer1_gen (.d_arr_0__31 (d_arr_merge1_0__31), .d_arr_0__30 (
               d_arr_merge1_0__30), .d_arr_0__29 (d_arr_merge1_0__29), .d_arr_0__28 (
               d_arr_merge1_0__28), .d_arr_0__27 (d_arr_merge1_0__27), .d_arr_0__26 (
               d_arr_merge1_0__26), .d_arr_0__25 (d_arr_merge1_0__25), .d_arr_0__24 (
               d_arr_merge1_0__24), .d_arr_0__23 (d_arr_merge1_0__23), .d_arr_0__22 (
               d_arr_merge1_0__22), .d_arr_0__21 (d_arr_merge1_0__21), .d_arr_0__20 (
               d_arr_merge1_0__20), .d_arr_0__19 (d_arr_merge1_0__19), .d_arr_0__18 (
               d_arr_merge1_0__18), .d_arr_0__17 (d_arr_merge1_0__17), .d_arr_0__16 (
               d_arr_merge1_0__16), .d_arr_0__15 (d_arr_merge1_0__15), .d_arr_0__14 (
               d_arr_merge1_0__14), .d_arr_0__13 (d_arr_merge1_0__13), .d_arr_0__12 (
               d_arr_merge1_0__12), .d_arr_0__11 (d_arr_merge1_0__11), .d_arr_0__10 (
               d_arr_merge1_0__10), .d_arr_0__9 (d_arr_merge1_0__9), .d_arr_0__8 (
               d_arr_merge1_0__8), .d_arr_0__7 (d_arr_merge1_0__7), .d_arr_0__6 (
               d_arr_merge1_0__6), .d_arr_0__5 (d_arr_merge1_0__5), .d_arr_0__4 (
               d_arr_merge1_0__4), .d_arr_0__3 (d_arr_merge1_0__3), .d_arr_0__2 (
               d_arr_merge1_0__2), .d_arr_0__1 (d_arr_merge1_0__1), .d_arr_0__0 (
               d_arr_merge1_0__0), .d_arr_1__31 (d_arr_merge1_1__31), .d_arr_1__30 (
               d_arr_merge1_1__30), .d_arr_1__29 (d_arr_merge1_1__29), .d_arr_1__28 (
               d_arr_merge1_1__28), .d_arr_1__27 (d_arr_merge1_1__27), .d_arr_1__26 (
               d_arr_merge1_1__26), .d_arr_1__25 (d_arr_merge1_1__25), .d_arr_1__24 (
               d_arr_merge1_1__24), .d_arr_1__23 (d_arr_merge1_1__23), .d_arr_1__22 (
               d_arr_merge1_1__22), .d_arr_1__21 (d_arr_merge1_1__21), .d_arr_1__20 (
               d_arr_merge1_1__20), .d_arr_1__19 (d_arr_merge1_1__19), .d_arr_1__18 (
               d_arr_merge1_1__18), .d_arr_1__17 (d_arr_merge1_1__17), .d_arr_1__16 (
               d_arr_merge1_1__16), .d_arr_1__15 (d_arr_merge1_1__15), .d_arr_1__14 (
               d_arr_merge1_1__14), .d_arr_1__13 (d_arr_merge1_1__13), .d_arr_1__12 (
               d_arr_merge1_1__12), .d_arr_1__11 (d_arr_merge1_1__11), .d_arr_1__10 (
               d_arr_merge1_1__10), .d_arr_1__9 (d_arr_merge1_1__9), .d_arr_1__8 (
               d_arr_merge1_1__8), .d_arr_1__7 (d_arr_merge1_1__7), .d_arr_1__6 (
               d_arr_merge1_1__6), .d_arr_1__5 (d_arr_merge1_1__5), .d_arr_1__4 (
               d_arr_merge1_1__4), .d_arr_1__3 (d_arr_merge1_1__3), .d_arr_1__2 (
               d_arr_merge1_1__2), .d_arr_1__1 (d_arr_merge1_1__1), .d_arr_1__0 (
               d_arr_merge1_1__0), .d_arr_2__31 (\$dummy [1216]), .d_arr_2__30 (
               \$dummy [1217]), .d_arr_2__29 (\$dummy [1218]), .d_arr_2__28 (
               \$dummy [1219]), .d_arr_2__27 (\$dummy [1220]), .d_arr_2__26 (
               \$dummy [1221]), .d_arr_2__25 (\$dummy [1222]), .d_arr_2__24 (
               \$dummy [1223]), .d_arr_2__23 (\$dummy [1224]), .d_arr_2__22 (
               \$dummy [1225]), .d_arr_2__21 (\$dummy [1226]), .d_arr_2__20 (
               \$dummy [1227]), .d_arr_2__19 (\$dummy [1228]), .d_arr_2__18 (
               \$dummy [1229]), .d_arr_2__17 (\$dummy [1230]), .d_arr_2__16 (
               \$dummy [1231]), .d_arr_2__15 (\$dummy [1232]), .d_arr_2__14 (
               \$dummy [1233]), .d_arr_2__13 (\$dummy [1234]), .d_arr_2__12 (
               \$dummy [1235]), .d_arr_2__11 (\$dummy [1236]), .d_arr_2__10 (
               \$dummy [1237]), .d_arr_2__9 (\$dummy [1238]), .d_arr_2__8 (
               \$dummy [1239]), .d_arr_2__7 (\$dummy [1240]), .d_arr_2__6 (
               \$dummy [1241]), .d_arr_2__5 (\$dummy [1242]), .d_arr_2__4 (
               \$dummy [1243]), .d_arr_2__3 (\$dummy [1244]), .d_arr_2__2 (
               \$dummy [1245]), .d_arr_2__1 (\$dummy [1246]), .d_arr_2__0 (
               \$dummy [1247]), .d_arr_3__31 (\$dummy [1248]), .d_arr_3__30 (
               \$dummy [1249]), .d_arr_3__29 (\$dummy [1250]), .d_arr_3__28 (
               \$dummy [1251]), .d_arr_3__27 (\$dummy [1252]), .d_arr_3__26 (
               \$dummy [1253]), .d_arr_3__25 (\$dummy [1254]), .d_arr_3__24 (
               \$dummy [1255]), .d_arr_3__23 (\$dummy [1256]), .d_arr_3__22 (
               \$dummy [1257]), .d_arr_3__21 (\$dummy [1258]), .d_arr_3__20 (
               \$dummy [1259]), .d_arr_3__19 (\$dummy [1260]), .d_arr_3__18 (
               \$dummy [1261]), .d_arr_3__17 (\$dummy [1262]), .d_arr_3__16 (
               \$dummy [1263]), .d_arr_3__15 (\$dummy [1264]), .d_arr_3__14 (
               \$dummy [1265]), .d_arr_3__13 (\$dummy [1266]), .d_arr_3__12 (
               \$dummy [1267]), .d_arr_3__11 (\$dummy [1268]), .d_arr_3__10 (
               \$dummy [1269]), .d_arr_3__9 (\$dummy [1270]), .d_arr_3__8 (
               \$dummy [1271]), .d_arr_3__7 (\$dummy [1272]), .d_arr_3__6 (
               \$dummy [1273]), .d_arr_3__5 (\$dummy [1274]), .d_arr_3__4 (
               \$dummy [1275]), .d_arr_3__3 (\$dummy [1276]), .d_arr_3__2 (
               \$dummy [1277]), .d_arr_3__1 (\$dummy [1278]), .d_arr_3__0 (
               \$dummy [1279]), .d_arr_4__31 (\$dummy [1280]), .d_arr_4__30 (
               \$dummy [1281]), .d_arr_4__29 (\$dummy [1282]), .d_arr_4__28 (
               \$dummy [1283]), .d_arr_4__27 (\$dummy [1284]), .d_arr_4__26 (
               \$dummy [1285]), .d_arr_4__25 (\$dummy [1286]), .d_arr_4__24 (
               \$dummy [1287]), .d_arr_4__23 (\$dummy [1288]), .d_arr_4__22 (
               \$dummy [1289]), .d_arr_4__21 (\$dummy [1290]), .d_arr_4__20 (
               \$dummy [1291]), .d_arr_4__19 (\$dummy [1292]), .d_arr_4__18 (
               \$dummy [1293]), .d_arr_4__17 (\$dummy [1294]), .d_arr_4__16 (
               \$dummy [1295]), .d_arr_4__15 (\$dummy [1296]), .d_arr_4__14 (
               \$dummy [1297]), .d_arr_4__13 (\$dummy [1298]), .d_arr_4__12 (
               \$dummy [1299]), .d_arr_4__11 (\$dummy [1300]), .d_arr_4__10 (
               \$dummy [1301]), .d_arr_4__9 (\$dummy [1302]), .d_arr_4__8 (
               \$dummy [1303]), .d_arr_4__7 (\$dummy [1304]), .d_arr_4__6 (
               \$dummy [1305]), .d_arr_4__5 (\$dummy [1306]), .d_arr_4__4 (
               \$dummy [1307]), .d_arr_4__3 (\$dummy [1308]), .d_arr_4__2 (
               \$dummy [1309]), .d_arr_4__1 (\$dummy [1310]), .d_arr_4__0 (
               \$dummy [1311]), .d_arr_5__31 (\$dummy [1312]), .d_arr_5__30 (
               \$dummy [1313]), .d_arr_5__29 (\$dummy [1314]), .d_arr_5__28 (
               \$dummy [1315]), .d_arr_5__27 (\$dummy [1316]), .d_arr_5__26 (
               \$dummy [1317]), .d_arr_5__25 (\$dummy [1318]), .d_arr_5__24 (
               \$dummy [1319]), .d_arr_5__23 (\$dummy [1320]), .d_arr_5__22 (
               \$dummy [1321]), .d_arr_5__21 (\$dummy [1322]), .d_arr_5__20 (
               \$dummy [1323]), .d_arr_5__19 (\$dummy [1324]), .d_arr_5__18 (
               \$dummy [1325]), .d_arr_5__17 (\$dummy [1326]), .d_arr_5__16 (
               \$dummy [1327]), .d_arr_5__15 (\$dummy [1328]), .d_arr_5__14 (
               \$dummy [1329]), .d_arr_5__13 (\$dummy [1330]), .d_arr_5__12 (
               \$dummy [1331]), .d_arr_5__11 (\$dummy [1332]), .d_arr_5__10 (
               \$dummy [1333]), .d_arr_5__9 (\$dummy [1334]), .d_arr_5__8 (
               \$dummy [1335]), .d_arr_5__7 (\$dummy [1336]), .d_arr_5__6 (
               \$dummy [1337]), .d_arr_5__5 (\$dummy [1338]), .d_arr_5__4 (
               \$dummy [1339]), .d_arr_5__3 (\$dummy [1340]), .d_arr_5__2 (
               \$dummy [1341]), .d_arr_5__1 (\$dummy [1342]), .d_arr_5__0 (
               \$dummy [1343]), .d_arr_6__31 (\$dummy [1344]), .d_arr_6__30 (
               \$dummy [1345]), .d_arr_6__29 (\$dummy [1346]), .d_arr_6__28 (
               \$dummy [1347]), .d_arr_6__27 (\$dummy [1348]), .d_arr_6__26 (
               \$dummy [1349]), .d_arr_6__25 (\$dummy [1350]), .d_arr_6__24 (
               \$dummy [1351]), .d_arr_6__23 (\$dummy [1352]), .d_arr_6__22 (
               \$dummy [1353]), .d_arr_6__21 (\$dummy [1354]), .d_arr_6__20 (
               \$dummy [1355]), .d_arr_6__19 (\$dummy [1356]), .d_arr_6__18 (
               \$dummy [1357]), .d_arr_6__17 (\$dummy [1358]), .d_arr_6__16 (
               \$dummy [1359]), .d_arr_6__15 (\$dummy [1360]), .d_arr_6__14 (
               \$dummy [1361]), .d_arr_6__13 (\$dummy [1362]), .d_arr_6__12 (
               \$dummy [1363]), .d_arr_6__11 (\$dummy [1364]), .d_arr_6__10 (
               \$dummy [1365]), .d_arr_6__9 (\$dummy [1366]), .d_arr_6__8 (
               \$dummy [1367]), .d_arr_6__7 (\$dummy [1368]), .d_arr_6__6 (
               \$dummy [1369]), .d_arr_6__5 (\$dummy [1370]), .d_arr_6__4 (
               \$dummy [1371]), .d_arr_6__3 (\$dummy [1372]), .d_arr_6__2 (
               \$dummy [1373]), .d_arr_6__1 (\$dummy [1374]), .d_arr_6__0 (
               \$dummy [1375]), .d_arr_7__31 (\$dummy [1376]), .d_arr_7__30 (
               \$dummy [1377]), .d_arr_7__29 (\$dummy [1378]), .d_arr_7__28 (
               \$dummy [1379]), .d_arr_7__27 (\$dummy [1380]), .d_arr_7__26 (
               \$dummy [1381]), .d_arr_7__25 (\$dummy [1382]), .d_arr_7__24 (
               \$dummy [1383]), .d_arr_7__23 (\$dummy [1384]), .d_arr_7__22 (
               \$dummy [1385]), .d_arr_7__21 (\$dummy [1386]), .d_arr_7__20 (
               \$dummy [1387]), .d_arr_7__19 (\$dummy [1388]), .d_arr_7__18 (
               \$dummy [1389]), .d_arr_7__17 (\$dummy [1390]), .d_arr_7__16 (
               \$dummy [1391]), .d_arr_7__15 (\$dummy [1392]), .d_arr_7__14 (
               \$dummy [1393]), .d_arr_7__13 (\$dummy [1394]), .d_arr_7__12 (
               \$dummy [1395]), .d_arr_7__11 (\$dummy [1396]), .d_arr_7__10 (
               \$dummy [1397]), .d_arr_7__9 (\$dummy [1398]), .d_arr_7__8 (
               \$dummy [1399]), .d_arr_7__7 (\$dummy [1400]), .d_arr_7__6 (
               \$dummy [1401]), .d_arr_7__5 (\$dummy [1402]), .d_arr_7__4 (
               \$dummy [1403]), .d_arr_7__3 (\$dummy [1404]), .d_arr_7__2 (
               \$dummy [1405]), .d_arr_7__1 (\$dummy [1406]), .d_arr_7__0 (
               \$dummy [1407]), .d_arr_8__31 (\$dummy [1408]), .d_arr_8__30 (
               \$dummy [1409]), .d_arr_8__29 (\$dummy [1410]), .d_arr_8__28 (
               \$dummy [1411]), .d_arr_8__27 (\$dummy [1412]), .d_arr_8__26 (
               \$dummy [1413]), .d_arr_8__25 (\$dummy [1414]), .d_arr_8__24 (
               \$dummy [1415]), .d_arr_8__23 (\$dummy [1416]), .d_arr_8__22 (
               \$dummy [1417]), .d_arr_8__21 (\$dummy [1418]), .d_arr_8__20 (
               \$dummy [1419]), .d_arr_8__19 (\$dummy [1420]), .d_arr_8__18 (
               \$dummy [1421]), .d_arr_8__17 (\$dummy [1422]), .d_arr_8__16 (
               \$dummy [1423]), .d_arr_8__15 (\$dummy [1424]), .d_arr_8__14 (
               \$dummy [1425]), .d_arr_8__13 (\$dummy [1426]), .d_arr_8__12 (
               \$dummy [1427]), .d_arr_8__11 (\$dummy [1428]), .d_arr_8__10 (
               \$dummy [1429]), .d_arr_8__9 (\$dummy [1430]), .d_arr_8__8 (
               \$dummy [1431]), .d_arr_8__7 (\$dummy [1432]), .d_arr_8__6 (
               \$dummy [1433]), .d_arr_8__5 (\$dummy [1434]), .d_arr_8__4 (
               \$dummy [1435]), .d_arr_8__3 (\$dummy [1436]), .d_arr_8__2 (
               \$dummy [1437]), .d_arr_8__1 (\$dummy [1438]), .d_arr_8__0 (
               \$dummy [1439]), .d_arr_9__31 (\$dummy [1440]), .d_arr_9__30 (
               \$dummy [1441]), .d_arr_9__29 (\$dummy [1442]), .d_arr_9__28 (
               \$dummy [1443]), .d_arr_9__27 (\$dummy [1444]), .d_arr_9__26 (
               \$dummy [1445]), .d_arr_9__25 (\$dummy [1446]), .d_arr_9__24 (
               \$dummy [1447]), .d_arr_9__23 (\$dummy [1448]), .d_arr_9__22 (
               \$dummy [1449]), .d_arr_9__21 (\$dummy [1450]), .d_arr_9__20 (
               \$dummy [1451]), .d_arr_9__19 (\$dummy [1452]), .d_arr_9__18 (
               \$dummy [1453]), .d_arr_9__17 (\$dummy [1454]), .d_arr_9__16 (
               \$dummy [1455]), .d_arr_9__15 (\$dummy [1456]), .d_arr_9__14 (
               \$dummy [1457]), .d_arr_9__13 (\$dummy [1458]), .d_arr_9__12 (
               \$dummy [1459]), .d_arr_9__11 (\$dummy [1460]), .d_arr_9__10 (
               \$dummy [1461]), .d_arr_9__9 (\$dummy [1462]), .d_arr_9__8 (
               \$dummy [1463]), .d_arr_9__7 (\$dummy [1464]), .d_arr_9__6 (
               \$dummy [1465]), .d_arr_9__5 (\$dummy [1466]), .d_arr_9__4 (
               \$dummy [1467]), .d_arr_9__3 (\$dummy [1468]), .d_arr_9__2 (
               \$dummy [1469]), .d_arr_9__1 (\$dummy [1470]), .d_arr_9__0 (
               \$dummy [1471]), .d_arr_10__31 (\$dummy [1472]), .d_arr_10__30 (
               \$dummy [1473]), .d_arr_10__29 (\$dummy [1474]), .d_arr_10__28 (
               \$dummy [1475]), .d_arr_10__27 (\$dummy [1476]), .d_arr_10__26 (
               \$dummy [1477]), .d_arr_10__25 (\$dummy [1478]), .d_arr_10__24 (
               \$dummy [1479]), .d_arr_10__23 (\$dummy [1480]), .d_arr_10__22 (
               \$dummy [1481]), .d_arr_10__21 (\$dummy [1482]), .d_arr_10__20 (
               \$dummy [1483]), .d_arr_10__19 (\$dummy [1484]), .d_arr_10__18 (
               \$dummy [1485]), .d_arr_10__17 (\$dummy [1486]), .d_arr_10__16 (
               \$dummy [1487]), .d_arr_10__15 (\$dummy [1488]), .d_arr_10__14 (
               \$dummy [1489]), .d_arr_10__13 (\$dummy [1490]), .d_arr_10__12 (
               \$dummy [1491]), .d_arr_10__11 (\$dummy [1492]), .d_arr_10__10 (
               \$dummy [1493]), .d_arr_10__9 (\$dummy [1494]), .d_arr_10__8 (
               \$dummy [1495]), .d_arr_10__7 (\$dummy [1496]), .d_arr_10__6 (
               \$dummy [1497]), .d_arr_10__5 (\$dummy [1498]), .d_arr_10__4 (
               \$dummy [1499]), .d_arr_10__3 (\$dummy [1500]), .d_arr_10__2 (
               \$dummy [1501]), .d_arr_10__1 (\$dummy [1502]), .d_arr_10__0 (
               \$dummy [1503]), .d_arr_11__31 (\$dummy [1504]), .d_arr_11__30 (
               \$dummy [1505]), .d_arr_11__29 (\$dummy [1506]), .d_arr_11__28 (
               \$dummy [1507]), .d_arr_11__27 (\$dummy [1508]), .d_arr_11__26 (
               \$dummy [1509]), .d_arr_11__25 (\$dummy [1510]), .d_arr_11__24 (
               \$dummy [1511]), .d_arr_11__23 (\$dummy [1512]), .d_arr_11__22 (
               \$dummy [1513]), .d_arr_11__21 (\$dummy [1514]), .d_arr_11__20 (
               \$dummy [1515]), .d_arr_11__19 (\$dummy [1516]), .d_arr_11__18 (
               \$dummy [1517]), .d_arr_11__17 (\$dummy [1518]), .d_arr_11__16 (
               \$dummy [1519]), .d_arr_11__15 (\$dummy [1520]), .d_arr_11__14 (
               \$dummy [1521]), .d_arr_11__13 (\$dummy [1522]), .d_arr_11__12 (
               \$dummy [1523]), .d_arr_11__11 (\$dummy [1524]), .d_arr_11__10 (
               \$dummy [1525]), .d_arr_11__9 (\$dummy [1526]), .d_arr_11__8 (
               \$dummy [1527]), .d_arr_11__7 (\$dummy [1528]), .d_arr_11__6 (
               \$dummy [1529]), .d_arr_11__5 (\$dummy [1530]), .d_arr_11__4 (
               \$dummy [1531]), .d_arr_11__3 (\$dummy [1532]), .d_arr_11__2 (
               \$dummy [1533]), .d_arr_11__1 (\$dummy [1534]), .d_arr_11__0 (
               \$dummy [1535]), .d_arr_12__31 (\$dummy [1536]), .d_arr_12__30 (
               \$dummy [1537]), .d_arr_12__29 (\$dummy [1538]), .d_arr_12__28 (
               \$dummy [1539]), .d_arr_12__27 (\$dummy [1540]), .d_arr_12__26 (
               \$dummy [1541]), .d_arr_12__25 (\$dummy [1542]), .d_arr_12__24 (
               \$dummy [1543]), .d_arr_12__23 (\$dummy [1544]), .d_arr_12__22 (
               \$dummy [1545]), .d_arr_12__21 (\$dummy [1546]), .d_arr_12__20 (
               \$dummy [1547]), .d_arr_12__19 (\$dummy [1548]), .d_arr_12__18 (
               \$dummy [1549]), .d_arr_12__17 (\$dummy [1550]), .d_arr_12__16 (
               \$dummy [1551]), .d_arr_12__15 (\$dummy [1552]), .d_arr_12__14 (
               \$dummy [1553]), .d_arr_12__13 (\$dummy [1554]), .d_arr_12__12 (
               \$dummy [1555]), .d_arr_12__11 (\$dummy [1556]), .d_arr_12__10 (
               \$dummy [1557]), .d_arr_12__9 (\$dummy [1558]), .d_arr_12__8 (
               \$dummy [1559]), .d_arr_12__7 (\$dummy [1560]), .d_arr_12__6 (
               \$dummy [1561]), .d_arr_12__5 (\$dummy [1562]), .d_arr_12__4 (
               \$dummy [1563]), .d_arr_12__3 (\$dummy [1564]), .d_arr_12__2 (
               \$dummy [1565]), .d_arr_12__1 (\$dummy [1566]), .d_arr_12__0 (
               \$dummy [1567]), .d_arr_13__31 (\$dummy [1568]), .d_arr_13__30 (
               \$dummy [1569]), .d_arr_13__29 (\$dummy [1570]), .d_arr_13__28 (
               \$dummy [1571]), .d_arr_13__27 (\$dummy [1572]), .d_arr_13__26 (
               \$dummy [1573]), .d_arr_13__25 (\$dummy [1574]), .d_arr_13__24 (
               \$dummy [1575]), .d_arr_13__23 (\$dummy [1576]), .d_arr_13__22 (
               \$dummy [1577]), .d_arr_13__21 (\$dummy [1578]), .d_arr_13__20 (
               \$dummy [1579]), .d_arr_13__19 (\$dummy [1580]), .d_arr_13__18 (
               \$dummy [1581]), .d_arr_13__17 (\$dummy [1582]), .d_arr_13__16 (
               \$dummy [1583]), .d_arr_13__15 (\$dummy [1584]), .d_arr_13__14 (
               \$dummy [1585]), .d_arr_13__13 (\$dummy [1586]), .d_arr_13__12 (
               \$dummy [1587]), .d_arr_13__11 (\$dummy [1588]), .d_arr_13__10 (
               \$dummy [1589]), .d_arr_13__9 (\$dummy [1590]), .d_arr_13__8 (
               \$dummy [1591]), .d_arr_13__7 (\$dummy [1592]), .d_arr_13__6 (
               \$dummy [1593]), .d_arr_13__5 (\$dummy [1594]), .d_arr_13__4 (
               \$dummy [1595]), .d_arr_13__3 (\$dummy [1596]), .d_arr_13__2 (
               \$dummy [1597]), .d_arr_13__1 (\$dummy [1598]), .d_arr_13__0 (
               \$dummy [1599]), .d_arr_14__31 (\$dummy [1600]), .d_arr_14__30 (
               \$dummy [1601]), .d_arr_14__29 (\$dummy [1602]), .d_arr_14__28 (
               \$dummy [1603]), .d_arr_14__27 (\$dummy [1604]), .d_arr_14__26 (
               \$dummy [1605]), .d_arr_14__25 (\$dummy [1606]), .d_arr_14__24 (
               \$dummy [1607]), .d_arr_14__23 (\$dummy [1608]), .d_arr_14__22 (
               \$dummy [1609]), .d_arr_14__21 (\$dummy [1610]), .d_arr_14__20 (
               \$dummy [1611]), .d_arr_14__19 (\$dummy [1612]), .d_arr_14__18 (
               \$dummy [1613]), .d_arr_14__17 (\$dummy [1614]), .d_arr_14__16 (
               \$dummy [1615]), .d_arr_14__15 (\$dummy [1616]), .d_arr_14__14 (
               \$dummy [1617]), .d_arr_14__13 (\$dummy [1618]), .d_arr_14__12 (
               \$dummy [1619]), .d_arr_14__11 (\$dummy [1620]), .d_arr_14__10 (
               \$dummy [1621]), .d_arr_14__9 (\$dummy [1622]), .d_arr_14__8 (
               \$dummy [1623]), .d_arr_14__7 (\$dummy [1624]), .d_arr_14__6 (
               \$dummy [1625]), .d_arr_14__5 (\$dummy [1626]), .d_arr_14__4 (
               \$dummy [1627]), .d_arr_14__3 (\$dummy [1628]), .d_arr_14__2 (
               \$dummy [1629]), .d_arr_14__1 (\$dummy [1630]), .d_arr_14__0 (
               \$dummy [1631]), .d_arr_15__31 (\$dummy [1632]), .d_arr_15__30 (
               \$dummy [1633]), .d_arr_15__29 (\$dummy [1634]), .d_arr_15__28 (
               \$dummy [1635]), .d_arr_15__27 (\$dummy [1636]), .d_arr_15__26 (
               \$dummy [1637]), .d_arr_15__25 (\$dummy [1638]), .d_arr_15__24 (
               \$dummy [1639]), .d_arr_15__23 (\$dummy [1640]), .d_arr_15__22 (
               \$dummy [1641]), .d_arr_15__21 (\$dummy [1642]), .d_arr_15__20 (
               \$dummy [1643]), .d_arr_15__19 (\$dummy [1644]), .d_arr_15__18 (
               \$dummy [1645]), .d_arr_15__17 (\$dummy [1646]), .d_arr_15__16 (
               \$dummy [1647]), .d_arr_15__15 (\$dummy [1648]), .d_arr_15__14 (
               \$dummy [1649]), .d_arr_15__13 (\$dummy [1650]), .d_arr_15__12 (
               \$dummy [1651]), .d_arr_15__11 (\$dummy [1652]), .d_arr_15__10 (
               \$dummy [1653]), .d_arr_15__9 (\$dummy [1654]), .d_arr_15__8 (
               \$dummy [1655]), .d_arr_15__7 (\$dummy [1656]), .d_arr_15__6 (
               \$dummy [1657]), .d_arr_15__5 (\$dummy [1658]), .d_arr_15__4 (
               \$dummy [1659]), .d_arr_15__3 (\$dummy [1660]), .d_arr_15__2 (
               \$dummy [1661]), .d_arr_15__1 (\$dummy [1662]), .d_arr_15__0 (
               \$dummy [1663]), .d_arr_16__31 (\$dummy [1664]), .d_arr_16__30 (
               \$dummy [1665]), .d_arr_16__29 (\$dummy [1666]), .d_arr_16__28 (
               \$dummy [1667]), .d_arr_16__27 (\$dummy [1668]), .d_arr_16__26 (
               \$dummy [1669]), .d_arr_16__25 (\$dummy [1670]), .d_arr_16__24 (
               \$dummy [1671]), .d_arr_16__23 (\$dummy [1672]), .d_arr_16__22 (
               \$dummy [1673]), .d_arr_16__21 (\$dummy [1674]), .d_arr_16__20 (
               \$dummy [1675]), .d_arr_16__19 (\$dummy [1676]), .d_arr_16__18 (
               \$dummy [1677]), .d_arr_16__17 (\$dummy [1678]), .d_arr_16__16 (
               \$dummy [1679]), .d_arr_16__15 (\$dummy [1680]), .d_arr_16__14 (
               \$dummy [1681]), .d_arr_16__13 (\$dummy [1682]), .d_arr_16__12 (
               \$dummy [1683]), .d_arr_16__11 (\$dummy [1684]), .d_arr_16__10 (
               \$dummy [1685]), .d_arr_16__9 (\$dummy [1686]), .d_arr_16__8 (
               \$dummy [1687]), .d_arr_16__7 (\$dummy [1688]), .d_arr_16__6 (
               \$dummy [1689]), .d_arr_16__5 (\$dummy [1690]), .d_arr_16__4 (
               \$dummy [1691]), .d_arr_16__3 (\$dummy [1692]), .d_arr_16__2 (
               \$dummy [1693]), .d_arr_16__1 (\$dummy [1694]), .d_arr_16__0 (
               \$dummy [1695]), .d_arr_17__31 (\$dummy [1696]), .d_arr_17__30 (
               \$dummy [1697]), .d_arr_17__29 (\$dummy [1698]), .d_arr_17__28 (
               \$dummy [1699]), .d_arr_17__27 (\$dummy [1700]), .d_arr_17__26 (
               \$dummy [1701]), .d_arr_17__25 (\$dummy [1702]), .d_arr_17__24 (
               \$dummy [1703]), .d_arr_17__23 (\$dummy [1704]), .d_arr_17__22 (
               \$dummy [1705]), .d_arr_17__21 (\$dummy [1706]), .d_arr_17__20 (
               \$dummy [1707]), .d_arr_17__19 (\$dummy [1708]), .d_arr_17__18 (
               \$dummy [1709]), .d_arr_17__17 (\$dummy [1710]), .d_arr_17__16 (
               \$dummy [1711]), .d_arr_17__15 (\$dummy [1712]), .d_arr_17__14 (
               \$dummy [1713]), .d_arr_17__13 (\$dummy [1714]), .d_arr_17__12 (
               \$dummy [1715]), .d_arr_17__11 (\$dummy [1716]), .d_arr_17__10 (
               \$dummy [1717]), .d_arr_17__9 (\$dummy [1718]), .d_arr_17__8 (
               \$dummy [1719]), .d_arr_17__7 (\$dummy [1720]), .d_arr_17__6 (
               \$dummy [1721]), .d_arr_17__5 (\$dummy [1722]), .d_arr_17__4 (
               \$dummy [1723]), .d_arr_17__3 (\$dummy [1724]), .d_arr_17__2 (
               \$dummy [1725]), .d_arr_17__1 (\$dummy [1726]), .d_arr_17__0 (
               \$dummy [1727]), .d_arr_18__31 (\$dummy [1728]), .d_arr_18__30 (
               \$dummy [1729]), .d_arr_18__29 (\$dummy [1730]), .d_arr_18__28 (
               \$dummy [1731]), .d_arr_18__27 (\$dummy [1732]), .d_arr_18__26 (
               \$dummy [1733]), .d_arr_18__25 (\$dummy [1734]), .d_arr_18__24 (
               \$dummy [1735]), .d_arr_18__23 (\$dummy [1736]), .d_arr_18__22 (
               \$dummy [1737]), .d_arr_18__21 (\$dummy [1738]), .d_arr_18__20 (
               \$dummy [1739]), .d_arr_18__19 (\$dummy [1740]), .d_arr_18__18 (
               \$dummy [1741]), .d_arr_18__17 (\$dummy [1742]), .d_arr_18__16 (
               \$dummy [1743]), .d_arr_18__15 (\$dummy [1744]), .d_arr_18__14 (
               \$dummy [1745]), .d_arr_18__13 (\$dummy [1746]), .d_arr_18__12 (
               \$dummy [1747]), .d_arr_18__11 (\$dummy [1748]), .d_arr_18__10 (
               \$dummy [1749]), .d_arr_18__9 (\$dummy [1750]), .d_arr_18__8 (
               \$dummy [1751]), .d_arr_18__7 (\$dummy [1752]), .d_arr_18__6 (
               \$dummy [1753]), .d_arr_18__5 (\$dummy [1754]), .d_arr_18__4 (
               \$dummy [1755]), .d_arr_18__3 (\$dummy [1756]), .d_arr_18__2 (
               \$dummy [1757]), .d_arr_18__1 (\$dummy [1758]), .d_arr_18__0 (
               \$dummy [1759]), .d_arr_19__31 (\$dummy [1760]), .d_arr_19__30 (
               \$dummy [1761]), .d_arr_19__29 (\$dummy [1762]), .d_arr_19__28 (
               \$dummy [1763]), .d_arr_19__27 (\$dummy [1764]), .d_arr_19__26 (
               \$dummy [1765]), .d_arr_19__25 (\$dummy [1766]), .d_arr_19__24 (
               \$dummy [1767]), .d_arr_19__23 (\$dummy [1768]), .d_arr_19__22 (
               \$dummy [1769]), .d_arr_19__21 (\$dummy [1770]), .d_arr_19__20 (
               \$dummy [1771]), .d_arr_19__19 (\$dummy [1772]), .d_arr_19__18 (
               \$dummy [1773]), .d_arr_19__17 (\$dummy [1774]), .d_arr_19__16 (
               \$dummy [1775]), .d_arr_19__15 (\$dummy [1776]), .d_arr_19__14 (
               \$dummy [1777]), .d_arr_19__13 (\$dummy [1778]), .d_arr_19__12 (
               \$dummy [1779]), .d_arr_19__11 (\$dummy [1780]), .d_arr_19__10 (
               \$dummy [1781]), .d_arr_19__9 (\$dummy [1782]), .d_arr_19__8 (
               \$dummy [1783]), .d_arr_19__7 (\$dummy [1784]), .d_arr_19__6 (
               \$dummy [1785]), .d_arr_19__5 (\$dummy [1786]), .d_arr_19__4 (
               \$dummy [1787]), .d_arr_19__3 (\$dummy [1788]), .d_arr_19__2 (
               \$dummy [1789]), .d_arr_19__1 (\$dummy [1790]), .d_arr_19__0 (
               \$dummy [1791]), .d_arr_20__31 (\$dummy [1792]), .d_arr_20__30 (
               \$dummy [1793]), .d_arr_20__29 (\$dummy [1794]), .d_arr_20__28 (
               \$dummy [1795]), .d_arr_20__27 (\$dummy [1796]), .d_arr_20__26 (
               \$dummy [1797]), .d_arr_20__25 (\$dummy [1798]), .d_arr_20__24 (
               \$dummy [1799]), .d_arr_20__23 (\$dummy [1800]), .d_arr_20__22 (
               \$dummy [1801]), .d_arr_20__21 (\$dummy [1802]), .d_arr_20__20 (
               \$dummy [1803]), .d_arr_20__19 (\$dummy [1804]), .d_arr_20__18 (
               \$dummy [1805]), .d_arr_20__17 (\$dummy [1806]), .d_arr_20__16 (
               \$dummy [1807]), .d_arr_20__15 (\$dummy [1808]), .d_arr_20__14 (
               \$dummy [1809]), .d_arr_20__13 (\$dummy [1810]), .d_arr_20__12 (
               \$dummy [1811]), .d_arr_20__11 (\$dummy [1812]), .d_arr_20__10 (
               \$dummy [1813]), .d_arr_20__9 (\$dummy [1814]), .d_arr_20__8 (
               \$dummy [1815]), .d_arr_20__7 (\$dummy [1816]), .d_arr_20__6 (
               \$dummy [1817]), .d_arr_20__5 (\$dummy [1818]), .d_arr_20__4 (
               \$dummy [1819]), .d_arr_20__3 (\$dummy [1820]), .d_arr_20__2 (
               \$dummy [1821]), .d_arr_20__1 (\$dummy [1822]), .d_arr_20__0 (
               \$dummy [1823]), .d_arr_21__31 (\$dummy [1824]), .d_arr_21__30 (
               \$dummy [1825]), .d_arr_21__29 (\$dummy [1826]), .d_arr_21__28 (
               \$dummy [1827]), .d_arr_21__27 (\$dummy [1828]), .d_arr_21__26 (
               \$dummy [1829]), .d_arr_21__25 (\$dummy [1830]), .d_arr_21__24 (
               \$dummy [1831]), .d_arr_21__23 (\$dummy [1832]), .d_arr_21__22 (
               \$dummy [1833]), .d_arr_21__21 (\$dummy [1834]), .d_arr_21__20 (
               \$dummy [1835]), .d_arr_21__19 (\$dummy [1836]), .d_arr_21__18 (
               \$dummy [1837]), .d_arr_21__17 (\$dummy [1838]), .d_arr_21__16 (
               \$dummy [1839]), .d_arr_21__15 (\$dummy [1840]), .d_arr_21__14 (
               \$dummy [1841]), .d_arr_21__13 (\$dummy [1842]), .d_arr_21__12 (
               \$dummy [1843]), .d_arr_21__11 (\$dummy [1844]), .d_arr_21__10 (
               \$dummy [1845]), .d_arr_21__9 (\$dummy [1846]), .d_arr_21__8 (
               \$dummy [1847]), .d_arr_21__7 (\$dummy [1848]), .d_arr_21__6 (
               \$dummy [1849]), .d_arr_21__5 (\$dummy [1850]), .d_arr_21__4 (
               \$dummy [1851]), .d_arr_21__3 (\$dummy [1852]), .d_arr_21__2 (
               \$dummy [1853]), .d_arr_21__1 (\$dummy [1854]), .d_arr_21__0 (
               \$dummy [1855]), .d_arr_22__31 (\$dummy [1856]), .d_arr_22__30 (
               \$dummy [1857]), .d_arr_22__29 (\$dummy [1858]), .d_arr_22__28 (
               \$dummy [1859]), .d_arr_22__27 (\$dummy [1860]), .d_arr_22__26 (
               \$dummy [1861]), .d_arr_22__25 (\$dummy [1862]), .d_arr_22__24 (
               \$dummy [1863]), .d_arr_22__23 (\$dummy [1864]), .d_arr_22__22 (
               \$dummy [1865]), .d_arr_22__21 (\$dummy [1866]), .d_arr_22__20 (
               \$dummy [1867]), .d_arr_22__19 (\$dummy [1868]), .d_arr_22__18 (
               \$dummy [1869]), .d_arr_22__17 (\$dummy [1870]), .d_arr_22__16 (
               \$dummy [1871]), .d_arr_22__15 (\$dummy [1872]), .d_arr_22__14 (
               \$dummy [1873]), .d_arr_22__13 (\$dummy [1874]), .d_arr_22__12 (
               \$dummy [1875]), .d_arr_22__11 (\$dummy [1876]), .d_arr_22__10 (
               \$dummy [1877]), .d_arr_22__9 (\$dummy [1878]), .d_arr_22__8 (
               \$dummy [1879]), .d_arr_22__7 (\$dummy [1880]), .d_arr_22__6 (
               \$dummy [1881]), .d_arr_22__5 (\$dummy [1882]), .d_arr_22__4 (
               \$dummy [1883]), .d_arr_22__3 (\$dummy [1884]), .d_arr_22__2 (
               \$dummy [1885]), .d_arr_22__1 (\$dummy [1886]), .d_arr_22__0 (
               \$dummy [1887]), .d_arr_23__31 (\$dummy [1888]), .d_arr_23__30 (
               \$dummy [1889]), .d_arr_23__29 (\$dummy [1890]), .d_arr_23__28 (
               \$dummy [1891]), .d_arr_23__27 (\$dummy [1892]), .d_arr_23__26 (
               \$dummy [1893]), .d_arr_23__25 (\$dummy [1894]), .d_arr_23__24 (
               \$dummy [1895]), .d_arr_23__23 (\$dummy [1896]), .d_arr_23__22 (
               \$dummy [1897]), .d_arr_23__21 (\$dummy [1898]), .d_arr_23__20 (
               \$dummy [1899]), .d_arr_23__19 (\$dummy [1900]), .d_arr_23__18 (
               \$dummy [1901]), .d_arr_23__17 (\$dummy [1902]), .d_arr_23__16 (
               \$dummy [1903]), .d_arr_23__15 (\$dummy [1904]), .d_arr_23__14 (
               \$dummy [1905]), .d_arr_23__13 (\$dummy [1906]), .d_arr_23__12 (
               \$dummy [1907]), .d_arr_23__11 (\$dummy [1908]), .d_arr_23__10 (
               \$dummy [1909]), .d_arr_23__9 (\$dummy [1910]), .d_arr_23__8 (
               \$dummy [1911]), .d_arr_23__7 (\$dummy [1912]), .d_arr_23__6 (
               \$dummy [1913]), .d_arr_23__5 (\$dummy [1914]), .d_arr_23__4 (
               \$dummy [1915]), .d_arr_23__3 (\$dummy [1916]), .d_arr_23__2 (
               \$dummy [1917]), .d_arr_23__1 (\$dummy [1918]), .d_arr_23__0 (
               \$dummy [1919]), .d_arr_24__31 (\$dummy [1920]), .d_arr_24__30 (
               \$dummy [1921]), .d_arr_24__29 (\$dummy [1922]), .d_arr_24__28 (
               \$dummy [1923]), .d_arr_24__27 (\$dummy [1924]), .d_arr_24__26 (
               \$dummy [1925]), .d_arr_24__25 (\$dummy [1926]), .d_arr_24__24 (
               \$dummy [1927]), .d_arr_24__23 (\$dummy [1928]), .d_arr_24__22 (
               \$dummy [1929]), .d_arr_24__21 (\$dummy [1930]), .d_arr_24__20 (
               \$dummy [1931]), .d_arr_24__19 (\$dummy [1932]), .d_arr_24__18 (
               \$dummy [1933]), .d_arr_24__17 (\$dummy [1934]), .d_arr_24__16 (
               \$dummy [1935]), .d_arr_24__15 (\$dummy [1936]), .d_arr_24__14 (
               \$dummy [1937]), .d_arr_24__13 (\$dummy [1938]), .d_arr_24__12 (
               \$dummy [1939]), .d_arr_24__11 (\$dummy [1940]), .d_arr_24__10 (
               \$dummy [1941]), .d_arr_24__9 (\$dummy [1942]), .d_arr_24__8 (
               \$dummy [1943]), .d_arr_24__7 (\$dummy [1944]), .d_arr_24__6 (
               \$dummy [1945]), .d_arr_24__5 (\$dummy [1946]), .d_arr_24__4 (
               \$dummy [1947]), .d_arr_24__3 (\$dummy [1948]), .d_arr_24__2 (
               \$dummy [1949]), .d_arr_24__1 (\$dummy [1950]), .d_arr_24__0 (
               \$dummy [1951]), .q_arr_0__31 (nx19448), .q_arr_0__30 (nx16499), 
               .q_arr_0__29 (nx16503), .q_arr_0__28 (nx16507), .q_arr_0__27 (
               nx19388), .q_arr_0__26 (nx16515), .q_arr_0__25 (nx16519), .q_arr_0__24 (
               nx19390), .q_arr_0__23 (nx16527), .q_arr_0__22 (nx16531), .q_arr_0__21 (
               nx16535), .q_arr_0__20 (nx16539), .q_arr_0__19 (nx16543), .q_arr_0__18 (
               nx16547), .q_arr_0__17 (nx16551), .q_arr_0__16 (nx16555), .q_arr_0__15 (
               nx16559), .q_arr_0__14 (nx16563), .q_arr_0__13 (nx16567), .q_arr_0__12 (
               nx16571), .q_arr_0__11 (nx16575), .q_arr_0__10 (nx16579), .q_arr_0__9 (
               nx16583), .q_arr_0__8 (nx16587), .q_arr_0__7 (nx16591), .q_arr_0__6 (
               nx16595), .q_arr_0__5 (nx16599), .q_arr_0__4 (nx16601), .q_arr_0__3 (
               nx16603), .q_arr_0__2 (q_arr_0__2), .q_arr_0__1 (q_arr_0__1), .q_arr_0__0 (
               nx16605), .q_arr_1__31 (GND0), .q_arr_1__30 (GND0), .q_arr_1__29 (
               GND0), .q_arr_1__28 (GND0), .q_arr_1__27 (GND0), .q_arr_1__26 (
               GND0), .q_arr_1__25 (GND0), .q_arr_1__24 (GND0), .q_arr_1__23 (
               GND0), .q_arr_1__22 (GND0), .q_arr_1__21 (GND0), .q_arr_1__20 (
               GND0), .q_arr_1__19 (GND0), .q_arr_1__18 (GND0), .q_arr_1__17 (
               GND0), .q_arr_1__16 (GND0), .q_arr_1__15 (GND0), .q_arr_1__14 (
               GND0), .q_arr_1__13 (GND0), .q_arr_1__12 (GND0), .q_arr_1__11 (
               GND0), .q_arr_1__10 (GND0), .q_arr_1__9 (GND0), .q_arr_1__8 (GND0
               ), .q_arr_1__7 (GND0), .q_arr_1__6 (GND0), .q_arr_1__5 (GND0), .q_arr_1__4 (
               GND0), .q_arr_1__3 (GND0), .q_arr_1__2 (GND0), .q_arr_1__1 (GND0)
               , .q_arr_1__0 (GND0), .q_arr_2__31 (GND0), .q_arr_2__30 (GND0), .q_arr_2__29 (
               GND0), .q_arr_2__28 (GND0), .q_arr_2__27 (GND0), .q_arr_2__26 (
               GND0), .q_arr_2__25 (GND0), .q_arr_2__24 (GND0), .q_arr_2__23 (
               GND0), .q_arr_2__22 (GND0), .q_arr_2__21 (GND0), .q_arr_2__20 (
               GND0), .q_arr_2__19 (GND0), .q_arr_2__18 (GND0), .q_arr_2__17 (
               GND0), .q_arr_2__16 (GND0), .q_arr_2__15 (GND0), .q_arr_2__14 (
               GND0), .q_arr_2__13 (GND0), .q_arr_2__12 (GND0), .q_arr_2__11 (
               GND0), .q_arr_2__10 (GND0), .q_arr_2__9 (GND0), .q_arr_2__8 (GND0
               ), .q_arr_2__7 (GND0), .q_arr_2__6 (GND0), .q_arr_2__5 (GND0), .q_arr_2__4 (
               GND0), .q_arr_2__3 (GND0), .q_arr_2__2 (GND0), .q_arr_2__1 (GND0)
               , .q_arr_2__0 (GND0), .q_arr_3__31 (GND0), .q_arr_3__30 (GND0), .q_arr_3__29 (
               GND0), .q_arr_3__28 (GND0), .q_arr_3__27 (GND0), .q_arr_3__26 (
               GND0), .q_arr_3__25 (GND0), .q_arr_3__24 (GND0), .q_arr_3__23 (
               GND0), .q_arr_3__22 (GND0), .q_arr_3__21 (GND0), .q_arr_3__20 (
               GND0), .q_arr_3__19 (GND0), .q_arr_3__18 (GND0), .q_arr_3__17 (
               GND0), .q_arr_3__16 (GND0), .q_arr_3__15 (GND0), .q_arr_3__14 (
               GND0), .q_arr_3__13 (GND0), .q_arr_3__12 (GND0), .q_arr_3__11 (
               GND0), .q_arr_3__10 (GND0), .q_arr_3__9 (GND0), .q_arr_3__8 (GND0
               ), .q_arr_3__7 (GND0), .q_arr_3__6 (GND0), .q_arr_3__5 (GND0), .q_arr_3__4 (
               GND0), .q_arr_3__3 (GND0), .q_arr_3__2 (GND0), .q_arr_3__1 (GND0)
               , .q_arr_3__0 (GND0), .q_arr_4__31 (GND0), .q_arr_4__30 (GND0), .q_arr_4__29 (
               GND0), .q_arr_4__28 (GND0), .q_arr_4__27 (GND0), .q_arr_4__26 (
               GND0), .q_arr_4__25 (GND0), .q_arr_4__24 (GND0), .q_arr_4__23 (
               GND0), .q_arr_4__22 (GND0), .q_arr_4__21 (GND0), .q_arr_4__20 (
               GND0), .q_arr_4__19 (GND0), .q_arr_4__18 (GND0), .q_arr_4__17 (
               GND0), .q_arr_4__16 (GND0), .q_arr_4__15 (GND0), .q_arr_4__14 (
               GND0), .q_arr_4__13 (GND0), .q_arr_4__12 (GND0), .q_arr_4__11 (
               GND0), .q_arr_4__10 (GND0), .q_arr_4__9 (GND0), .q_arr_4__8 (GND0
               ), .q_arr_4__7 (GND0), .q_arr_4__6 (GND0), .q_arr_4__5 (GND0), .q_arr_4__4 (
               GND0), .q_arr_4__3 (GND0), .q_arr_4__2 (GND0), .q_arr_4__1 (GND0)
               , .q_arr_4__0 (GND0), .q_arr_5__31 (GND0), .q_arr_5__30 (GND0), .q_arr_5__29 (
               GND0), .q_arr_5__28 (GND0), .q_arr_5__27 (GND0), .q_arr_5__26 (
               GND0), .q_arr_5__25 (GND0), .q_arr_5__24 (GND0), .q_arr_5__23 (
               GND0), .q_arr_5__22 (GND0), .q_arr_5__21 (GND0), .q_arr_5__20 (
               GND0), .q_arr_5__19 (GND0), .q_arr_5__18 (GND0), .q_arr_5__17 (
               GND0), .q_arr_5__16 (GND0), .q_arr_5__15 (GND0), .q_arr_5__14 (
               GND0), .q_arr_5__13 (GND0), .q_arr_5__12 (GND0), .q_arr_5__11 (
               GND0), .q_arr_5__10 (GND0), .q_arr_5__9 (GND0), .q_arr_5__8 (GND0
               ), .q_arr_5__7 (GND0), .q_arr_5__6 (GND0), .q_arr_5__5 (GND0), .q_arr_5__4 (
               GND0), .q_arr_5__3 (GND0), .q_arr_5__2 (GND0), .q_arr_5__1 (GND0)
               , .q_arr_5__0 (GND0), .q_arr_6__31 (GND0), .q_arr_6__30 (GND0), .q_arr_6__29 (
               GND0), .q_arr_6__28 (GND0), .q_arr_6__27 (GND0), .q_arr_6__26 (
               GND0), .q_arr_6__25 (GND0), .q_arr_6__24 (GND0), .q_arr_6__23 (
               GND0), .q_arr_6__22 (GND0), .q_arr_6__21 (GND0), .q_arr_6__20 (
               GND0), .q_arr_6__19 (GND0), .q_arr_6__18 (GND0), .q_arr_6__17 (
               GND0), .q_arr_6__16 (GND0), .q_arr_6__15 (GND0), .q_arr_6__14 (
               GND0), .q_arr_6__13 (GND0), .q_arr_6__12 (GND0), .q_arr_6__11 (
               GND0), .q_arr_6__10 (GND0), .q_arr_6__9 (GND0), .q_arr_6__8 (GND0
               ), .q_arr_6__7 (GND0), .q_arr_6__6 (GND0), .q_arr_6__5 (GND0), .q_arr_6__4 (
               GND0), .q_arr_6__3 (GND0), .q_arr_6__2 (GND0), .q_arr_6__1 (GND0)
               , .q_arr_6__0 (GND0), .q_arr_7__31 (GND0), .q_arr_7__30 (GND0), .q_arr_7__29 (
               GND0), .q_arr_7__28 (GND0), .q_arr_7__27 (GND0), .q_arr_7__26 (
               GND0), .q_arr_7__25 (GND0), .q_arr_7__24 (GND0), .q_arr_7__23 (
               GND0), .q_arr_7__22 (GND0), .q_arr_7__21 (GND0), .q_arr_7__20 (
               GND0), .q_arr_7__19 (GND0), .q_arr_7__18 (GND0), .q_arr_7__17 (
               GND0), .q_arr_7__16 (GND0), .q_arr_7__15 (GND0), .q_arr_7__14 (
               GND0), .q_arr_7__13 (GND0), .q_arr_7__12 (GND0), .q_arr_7__11 (
               GND0), .q_arr_7__10 (GND0), .q_arr_7__9 (GND0), .q_arr_7__8 (GND0
               ), .q_arr_7__7 (GND0), .q_arr_7__6 (GND0), .q_arr_7__5 (GND0), .q_arr_7__4 (
               GND0), .q_arr_7__3 (GND0), .q_arr_7__2 (GND0), .q_arr_7__1 (GND0)
               , .q_arr_7__0 (GND0), .q_arr_8__31 (GND0), .q_arr_8__30 (GND0), .q_arr_8__29 (
               GND0), .q_arr_8__28 (GND0), .q_arr_8__27 (GND0), .q_arr_8__26 (
               GND0), .q_arr_8__25 (GND0), .q_arr_8__24 (GND0), .q_arr_8__23 (
               GND0), .q_arr_8__22 (GND0), .q_arr_8__21 (GND0), .q_arr_8__20 (
               GND0), .q_arr_8__19 (GND0), .q_arr_8__18 (GND0), .q_arr_8__17 (
               GND0), .q_arr_8__16 (GND0), .q_arr_8__15 (GND0), .q_arr_8__14 (
               GND0), .q_arr_8__13 (GND0), .q_arr_8__12 (GND0), .q_arr_8__11 (
               GND0), .q_arr_8__10 (GND0), .q_arr_8__9 (GND0), .q_arr_8__8 (GND0
               ), .q_arr_8__7 (GND0), .q_arr_8__6 (GND0), .q_arr_8__5 (GND0), .q_arr_8__4 (
               GND0), .q_arr_8__3 (GND0), .q_arr_8__2 (GND0), .q_arr_8__1 (GND0)
               , .q_arr_8__0 (GND0), .q_arr_9__31 (q_arr_9__31), .q_arr_9__30 (
               q_arr_9__30), .q_arr_9__29 (q_arr_9__29), .q_arr_9__28 (
               q_arr_9__28), .q_arr_9__27 (q_arr_9__27), .q_arr_9__26 (
               q_arr_9__26), .q_arr_9__25 (q_arr_9__25), .q_arr_9__24 (
               q_arr_9__24), .q_arr_9__23 (q_arr_9__23), .q_arr_9__22 (
               q_arr_9__22), .q_arr_9__21 (q_arr_9__21), .q_arr_9__20 (
               q_arr_9__20), .q_arr_9__19 (q_arr_9__19), .q_arr_9__18 (
               q_arr_9__18), .q_arr_9__17 (q_arr_9__17), .q_arr_9__16 (
               q_arr_9__16), .q_arr_9__15 (q_arr_9__15), .q_arr_9__14 (
               q_arr_9__14), .q_arr_9__13 (q_arr_9__13), .q_arr_9__12 (
               q_arr_9__12), .q_arr_9__11 (q_arr_9__11), .q_arr_9__10 (
               q_arr_9__10), .q_arr_9__9 (q_arr_9__9), .q_arr_9__8 (q_arr_9__8)
               , .q_arr_9__7 (q_arr_9__7), .q_arr_9__6 (q_arr_9__6), .q_arr_9__5 (
               q_arr_9__5), .q_arr_9__4 (q_arr_9__4), .q_arr_9__3 (q_arr_9__3), 
               .q_arr_9__2 (q_arr_9__2), .q_arr_9__1 (q_arr_9__1), .q_arr_9__0 (
               q_arr_9__0), .q_arr_10__31 (GND0), .q_arr_10__30 (GND0), .q_arr_10__29 (
               GND0), .q_arr_10__28 (GND0), .q_arr_10__27 (GND0), .q_arr_10__26 (
               GND0), .q_arr_10__25 (GND0), .q_arr_10__24 (GND0), .q_arr_10__23 (
               GND0), .q_arr_10__22 (GND0), .q_arr_10__21 (GND0), .q_arr_10__20 (
               GND0), .q_arr_10__19 (GND0), .q_arr_10__18 (GND0), .q_arr_10__17 (
               GND0), .q_arr_10__16 (GND0), .q_arr_10__15 (GND0), .q_arr_10__14 (
               GND0), .q_arr_10__13 (GND0), .q_arr_10__12 (GND0), .q_arr_10__11 (
               GND0), .q_arr_10__10 (GND0), .q_arr_10__9 (GND0), .q_arr_10__8 (
               GND0), .q_arr_10__7 (GND0), .q_arr_10__6 (GND0), .q_arr_10__5 (
               GND0), .q_arr_10__4 (GND0), .q_arr_10__3 (GND0), .q_arr_10__2 (
               GND0), .q_arr_10__1 (GND0), .q_arr_10__0 (GND0), .q_arr_11__31 (
               GND0), .q_arr_11__30 (GND0), .q_arr_11__29 (GND0), .q_arr_11__28 (
               GND0), .q_arr_11__27 (GND0), .q_arr_11__26 (GND0), .q_arr_11__25 (
               GND0), .q_arr_11__24 (GND0), .q_arr_11__23 (GND0), .q_arr_11__22 (
               GND0), .q_arr_11__21 (GND0), .q_arr_11__20 (GND0), .q_arr_11__19 (
               GND0), .q_arr_11__18 (GND0), .q_arr_11__17 (GND0), .q_arr_11__16 (
               GND0), .q_arr_11__15 (GND0), .q_arr_11__14 (GND0), .q_arr_11__13 (
               GND0), .q_arr_11__12 (GND0), .q_arr_11__11 (GND0), .q_arr_11__10 (
               GND0), .q_arr_11__9 (GND0), .q_arr_11__8 (GND0), .q_arr_11__7 (
               GND0), .q_arr_11__6 (GND0), .q_arr_11__5 (GND0), .q_arr_11__4 (
               GND0), .q_arr_11__3 (GND0), .q_arr_11__2 (GND0), .q_arr_11__1 (
               GND0), .q_arr_11__0 (GND0), .q_arr_12__31 (GND0), .q_arr_12__30 (
               GND0), .q_arr_12__29 (GND0), .q_arr_12__28 (GND0), .q_arr_12__27 (
               GND0), .q_arr_12__26 (GND0), .q_arr_12__25 (GND0), .q_arr_12__24 (
               GND0), .q_arr_12__23 (GND0), .q_arr_12__22 (GND0), .q_arr_12__21 (
               GND0), .q_arr_12__20 (GND0), .q_arr_12__19 (GND0), .q_arr_12__18 (
               GND0), .q_arr_12__17 (GND0), .q_arr_12__16 (GND0), .q_arr_12__15 (
               GND0), .q_arr_12__14 (GND0), .q_arr_12__13 (GND0), .q_arr_12__12 (
               GND0), .q_arr_12__11 (GND0), .q_arr_12__10 (GND0), .q_arr_12__9 (
               GND0), .q_arr_12__8 (GND0), .q_arr_12__7 (GND0), .q_arr_12__6 (
               GND0), .q_arr_12__5 (GND0), .q_arr_12__4 (GND0), .q_arr_12__3 (
               GND0), .q_arr_12__2 (GND0), .q_arr_12__1 (GND0), .q_arr_12__0 (
               GND0), .q_arr_13__31 (GND0), .q_arr_13__30 (GND0), .q_arr_13__29 (
               GND0), .q_arr_13__28 (GND0), .q_arr_13__27 (GND0), .q_arr_13__26 (
               GND0), .q_arr_13__25 (GND0), .q_arr_13__24 (GND0), .q_arr_13__23 (
               GND0), .q_arr_13__22 (GND0), .q_arr_13__21 (GND0), .q_arr_13__20 (
               GND0), .q_arr_13__19 (GND0), .q_arr_13__18 (GND0), .q_arr_13__17 (
               GND0), .q_arr_13__16 (GND0), .q_arr_13__15 (GND0), .q_arr_13__14 (
               GND0), .q_arr_13__13 (GND0), .q_arr_13__12 (GND0), .q_arr_13__11 (
               GND0), .q_arr_13__10 (GND0), .q_arr_13__9 (GND0), .q_arr_13__8 (
               GND0), .q_arr_13__7 (GND0), .q_arr_13__6 (GND0), .q_arr_13__5 (
               GND0), .q_arr_13__4 (GND0), .q_arr_13__3 (GND0), .q_arr_13__2 (
               GND0), .q_arr_13__1 (GND0), .q_arr_13__0 (GND0), .q_arr_14__31 (
               GND0), .q_arr_14__30 (GND0), .q_arr_14__29 (GND0), .q_arr_14__28 (
               GND0), .q_arr_14__27 (GND0), .q_arr_14__26 (GND0), .q_arr_14__25 (
               GND0), .q_arr_14__24 (GND0), .q_arr_14__23 (GND0), .q_arr_14__22 (
               GND0), .q_arr_14__21 (GND0), .q_arr_14__20 (GND0), .q_arr_14__19 (
               GND0), .q_arr_14__18 (GND0), .q_arr_14__17 (GND0), .q_arr_14__16 (
               GND0), .q_arr_14__15 (GND0), .q_arr_14__14 (GND0), .q_arr_14__13 (
               GND0), .q_arr_14__12 (GND0), .q_arr_14__11 (GND0), .q_arr_14__10 (
               GND0), .q_arr_14__9 (GND0), .q_arr_14__8 (GND0), .q_arr_14__7 (
               GND0), .q_arr_14__6 (GND0), .q_arr_14__5 (GND0), .q_arr_14__4 (
               GND0), .q_arr_14__3 (GND0), .q_arr_14__2 (GND0), .q_arr_14__1 (
               GND0), .q_arr_14__0 (GND0), .q_arr_15__31 (GND0), .q_arr_15__30 (
               GND0), .q_arr_15__29 (GND0), .q_arr_15__28 (GND0), .q_arr_15__27 (
               GND0), .q_arr_15__26 (GND0), .q_arr_15__25 (GND0), .q_arr_15__24 (
               GND0), .q_arr_15__23 (GND0), .q_arr_15__22 (GND0), .q_arr_15__21 (
               GND0), .q_arr_15__20 (GND0), .q_arr_15__19 (GND0), .q_arr_15__18 (
               GND0), .q_arr_15__17 (GND0), .q_arr_15__16 (GND0), .q_arr_15__15 (
               GND0), .q_arr_15__14 (GND0), .q_arr_15__13 (GND0), .q_arr_15__12 (
               GND0), .q_arr_15__11 (GND0), .q_arr_15__10 (GND0), .q_arr_15__9 (
               GND0), .q_arr_15__8 (GND0), .q_arr_15__7 (GND0), .q_arr_15__6 (
               GND0), .q_arr_15__5 (GND0), .q_arr_15__4 (GND0), .q_arr_15__3 (
               GND0), .q_arr_15__2 (GND0), .q_arr_15__1 (GND0), .q_arr_15__0 (
               GND0), .q_arr_16__31 (GND0), .q_arr_16__30 (GND0), .q_arr_16__29 (
               GND0), .q_arr_16__28 (GND0), .q_arr_16__27 (GND0), .q_arr_16__26 (
               GND0), .q_arr_16__25 (GND0), .q_arr_16__24 (GND0), .q_arr_16__23 (
               GND0), .q_arr_16__22 (GND0), .q_arr_16__21 (GND0), .q_arr_16__20 (
               GND0), .q_arr_16__19 (GND0), .q_arr_16__18 (GND0), .q_arr_16__17 (
               GND0), .q_arr_16__16 (GND0), .q_arr_16__15 (GND0), .q_arr_16__14 (
               GND0), .q_arr_16__13 (GND0), .q_arr_16__12 (GND0), .q_arr_16__11 (
               GND0), .q_arr_16__10 (GND0), .q_arr_16__9 (GND0), .q_arr_16__8 (
               GND0), .q_arr_16__7 (GND0), .q_arr_16__6 (GND0), .q_arr_16__5 (
               GND0), .q_arr_16__4 (GND0), .q_arr_16__3 (GND0), .q_arr_16__2 (
               GND0), .q_arr_16__1 (GND0), .q_arr_16__0 (GND0), .q_arr_17__31 (
               GND0), .q_arr_17__30 (GND0), .q_arr_17__29 (GND0), .q_arr_17__28 (
               GND0), .q_arr_17__27 (GND0), .q_arr_17__26 (GND0), .q_arr_17__25 (
               GND0), .q_arr_17__24 (GND0), .q_arr_17__23 (GND0), .q_arr_17__22 (
               GND0), .q_arr_17__21 (GND0), .q_arr_17__20 (GND0), .q_arr_17__19 (
               GND0), .q_arr_17__18 (GND0), .q_arr_17__17 (GND0), .q_arr_17__16 (
               GND0), .q_arr_17__15 (GND0), .q_arr_17__14 (GND0), .q_arr_17__13 (
               GND0), .q_arr_17__12 (GND0), .q_arr_17__11 (GND0), .q_arr_17__10 (
               GND0), .q_arr_17__9 (GND0), .q_arr_17__8 (GND0), .q_arr_17__7 (
               GND0), .q_arr_17__6 (GND0), .q_arr_17__5 (GND0), .q_arr_17__4 (
               GND0), .q_arr_17__3 (GND0), .q_arr_17__2 (GND0), .q_arr_17__1 (
               GND0), .q_arr_17__0 (GND0), .q_arr_18__31 (q_arr_18__31), .q_arr_18__30 (
               q_arr_18__30), .q_arr_18__29 (q_arr_18__29), .q_arr_18__28 (
               q_arr_18__28), .q_arr_18__27 (nx19488), .q_arr_18__26 (
               q_arr_18__26), .q_arr_18__25 (q_arr_18__25), .q_arr_18__24 (
               nx19492), .q_arr_18__23 (q_arr_18__23), .q_arr_18__22 (
               q_arr_18__22), .q_arr_18__21 (q_arr_18__21), .q_arr_18__20 (
               q_arr_18__20), .q_arr_18__19 (q_arr_18__19), .q_arr_18__18 (
               q_arr_18__18), .q_arr_18__17 (q_arr_18__17), .q_arr_18__16 (
               q_arr_18__16), .q_arr_18__15 (q_arr_18__15), .q_arr_18__14 (
               q_arr_18__14), .q_arr_18__13 (q_arr_18__13), .q_arr_18__12 (
               q_arr_18__12), .q_arr_18__11 (q_arr_18__11), .q_arr_18__10 (
               q_arr_18__10), .q_arr_18__9 (q_arr_18__9), .q_arr_18__8 (
               q_arr_18__8), .q_arr_18__7 (q_arr_18__7), .q_arr_18__6 (
               q_arr_18__6), .q_arr_18__5 (q_arr_18__5), .q_arr_18__4 (
               q_arr_18__4), .q_arr_18__3 (q_arr_18__3), .q_arr_18__2 (
               q_arr_18__2), .q_arr_18__1 (q_arr_18__1), .q_arr_18__0 (
               q_arr_18__0), .q_arr_19__31 (GND0), .q_arr_19__30 (GND0), .q_arr_19__29 (
               GND0), .q_arr_19__28 (GND0), .q_arr_19__27 (GND0), .q_arr_19__26 (
               GND0), .q_arr_19__25 (GND0), .q_arr_19__24 (GND0), .q_arr_19__23 (
               GND0), .q_arr_19__22 (GND0), .q_arr_19__21 (GND0), .q_arr_19__20 (
               GND0), .q_arr_19__19 (GND0), .q_arr_19__18 (GND0), .q_arr_19__17 (
               GND0), .q_arr_19__16 (GND0), .q_arr_19__15 (GND0), .q_arr_19__14 (
               GND0), .q_arr_19__13 (GND0), .q_arr_19__12 (GND0), .q_arr_19__11 (
               GND0), .q_arr_19__10 (GND0), .q_arr_19__9 (GND0), .q_arr_19__8 (
               GND0), .q_arr_19__7 (GND0), .q_arr_19__6 (GND0), .q_arr_19__5 (
               GND0), .q_arr_19__4 (GND0), .q_arr_19__3 (GND0), .q_arr_19__2 (
               GND0), .q_arr_19__1 (GND0), .q_arr_19__0 (GND0), .q_arr_20__31 (
               GND0), .q_arr_20__30 (GND0), .q_arr_20__29 (GND0), .q_arr_20__28 (
               GND0), .q_arr_20__27 (GND0), .q_arr_20__26 (GND0), .q_arr_20__25 (
               GND0), .q_arr_20__24 (GND0), .q_arr_20__23 (GND0), .q_arr_20__22 (
               GND0), .q_arr_20__21 (GND0), .q_arr_20__20 (GND0), .q_arr_20__19 (
               GND0), .q_arr_20__18 (GND0), .q_arr_20__17 (GND0), .q_arr_20__16 (
               GND0), .q_arr_20__15 (GND0), .q_arr_20__14 (GND0), .q_arr_20__13 (
               GND0), .q_arr_20__12 (GND0), .q_arr_20__11 (GND0), .q_arr_20__10 (
               GND0), .q_arr_20__9 (GND0), .q_arr_20__8 (GND0), .q_arr_20__7 (
               GND0), .q_arr_20__6 (GND0), .q_arr_20__5 (GND0), .q_arr_20__4 (
               GND0), .q_arr_20__3 (GND0), .q_arr_20__2 (GND0), .q_arr_20__1 (
               GND0), .q_arr_20__0 (GND0), .q_arr_21__31 (GND0), .q_arr_21__30 (
               GND0), .q_arr_21__29 (GND0), .q_arr_21__28 (GND0), .q_arr_21__27 (
               GND0), .q_arr_21__26 (GND0), .q_arr_21__25 (GND0), .q_arr_21__24 (
               GND0), .q_arr_21__23 (GND0), .q_arr_21__22 (GND0), .q_arr_21__21 (
               GND0), .q_arr_21__20 (GND0), .q_arr_21__19 (GND0), .q_arr_21__18 (
               GND0), .q_arr_21__17 (GND0), .q_arr_21__16 (GND0), .q_arr_21__15 (
               GND0), .q_arr_21__14 (GND0), .q_arr_21__13 (GND0), .q_arr_21__12 (
               GND0), .q_arr_21__11 (GND0), .q_arr_21__10 (GND0), .q_arr_21__9 (
               GND0), .q_arr_21__8 (GND0), .q_arr_21__7 (GND0), .q_arr_21__6 (
               GND0), .q_arr_21__5 (GND0), .q_arr_21__4 (GND0), .q_arr_21__3 (
               GND0), .q_arr_21__2 (GND0), .q_arr_21__1 (GND0), .q_arr_21__0 (
               GND0), .q_arr_22__31 (GND0), .q_arr_22__30 (GND0), .q_arr_22__29 (
               GND0), .q_arr_22__28 (GND0), .q_arr_22__27 (GND0), .q_arr_22__26 (
               GND0), .q_arr_22__25 (GND0), .q_arr_22__24 (GND0), .q_arr_22__23 (
               GND0), .q_arr_22__22 (GND0), .q_arr_22__21 (GND0), .q_arr_22__20 (
               GND0), .q_arr_22__19 (GND0), .q_arr_22__18 (GND0), .q_arr_22__17 (
               GND0), .q_arr_22__16 (GND0), .q_arr_22__15 (GND0), .q_arr_22__14 (
               GND0), .q_arr_22__13 (GND0), .q_arr_22__12 (GND0), .q_arr_22__11 (
               GND0), .q_arr_22__10 (GND0), .q_arr_22__9 (GND0), .q_arr_22__8 (
               GND0), .q_arr_22__7 (GND0), .q_arr_22__6 (GND0), .q_arr_22__5 (
               GND0), .q_arr_22__4 (GND0), .q_arr_22__3 (GND0), .q_arr_22__2 (
               GND0), .q_arr_22__1 (GND0), .q_arr_22__0 (GND0), .q_arr_23__31 (
               GND0), .q_arr_23__30 (GND0), .q_arr_23__29 (GND0), .q_arr_23__28 (
               GND0), .q_arr_23__27 (GND0), .q_arr_23__26 (GND0), .q_arr_23__25 (
               GND0), .q_arr_23__24 (GND0), .q_arr_23__23 (GND0), .q_arr_23__22 (
               GND0), .q_arr_23__21 (GND0), .q_arr_23__20 (GND0), .q_arr_23__19 (
               GND0), .q_arr_23__18 (GND0), .q_arr_23__17 (GND0), .q_arr_23__16 (
               GND0), .q_arr_23__15 (GND0), .q_arr_23__14 (GND0), .q_arr_23__13 (
               GND0), .q_arr_23__12 (GND0), .q_arr_23__11 (GND0), .q_arr_23__10 (
               GND0), .q_arr_23__9 (GND0), .q_arr_23__8 (GND0), .q_arr_23__7 (
               GND0), .q_arr_23__6 (GND0), .q_arr_23__5 (GND0), .q_arr_23__4 (
               GND0), .q_arr_23__3 (GND0), .q_arr_23__2 (GND0), .q_arr_23__1 (
               GND0), .q_arr_23__0 (GND0), .q_arr_24__31 (GND0), .q_arr_24__30 (
               GND0), .q_arr_24__29 (GND0), .q_arr_24__28 (GND0), .q_arr_24__27 (
               GND0), .q_arr_24__26 (GND0), .q_arr_24__25 (GND0), .q_arr_24__24 (
               GND0), .q_arr_24__23 (GND0), .q_arr_24__22 (GND0), .q_arr_24__21 (
               GND0), .q_arr_24__20 (GND0), .q_arr_24__19 (GND0), .q_arr_24__18 (
               GND0), .q_arr_24__17 (GND0), .q_arr_24__16 (GND0), .q_arr_24__15 (
               GND0), .q_arr_24__14 (GND0), .q_arr_24__13 (GND0), .q_arr_24__12 (
               GND0), .q_arr_24__11 (GND0), .q_arr_24__10 (GND0), .q_arr_24__9 (
               GND0), .q_arr_24__8 (GND0), .q_arr_24__7 (GND0), .q_arr_24__6 (
               GND0), .q_arr_24__5 (GND0), .q_arr_24__4 (GND0), .q_arr_24__3 (
               GND0), .q_arr_24__2 (GND0), .q_arr_24__1 (GND0), .q_arr_24__0 (
               GND0), .operation (operation), .filter_size (nx16667)) ;
    ReluLayer relu_layer_gen (.d_arr_0__31 (d_arr_relu_0__31), .d_arr_0__30 (
              d_arr_relu_0__30), .d_arr_0__29 (d_arr_relu_0__29), .d_arr_0__28 (
              d_arr_relu_0__28), .d_arr_0__27 (d_arr_relu_0__27), .d_arr_0__26 (
              d_arr_relu_0__26), .d_arr_0__25 (d_arr_relu_0__25), .d_arr_0__24 (
              d_arr_relu_0__24), .d_arr_0__23 (d_arr_relu_0__23), .d_arr_0__22 (
              d_arr_relu_0__22), .d_arr_0__21 (d_arr_relu_0__21), .d_arr_0__20 (
              d_arr_relu_0__20), .d_arr_0__19 (d_arr_relu_0__19), .d_arr_0__18 (
              d_arr_relu_0__18), .d_arr_0__17 (d_arr_relu_0__17), .d_arr_0__16 (
              d_arr_relu_0__16), .d_arr_0__15 (\$dummy [1952]), .d_arr_0__14 (
              d_arr_relu_0__14), .d_arr_0__13 (d_arr_relu_0__13), .d_arr_0__12 (
              d_arr_relu_0__12), .d_arr_0__11 (d_arr_relu_0__11), .d_arr_0__10 (
              d_arr_relu_0__10), .d_arr_0__9 (d_arr_relu_0__9), .d_arr_0__8 (
              d_arr_relu_0__8), .d_arr_0__7 (d_arr_relu_0__7), .d_arr_0__6 (
              d_arr_relu_0__6), .d_arr_0__5 (d_arr_relu_0__5), .d_arr_0__4 (
              d_arr_relu_0__4), .d_arr_0__3 (d_arr_relu_0__3), .d_arr_0__2 (
              d_arr_relu_0__2), .d_arr_0__1 (d_arr_relu_0__1), .d_arr_0__0 (
              d_arr_relu_0__0), .d_arr_1__31 (d_arr_relu_1__31), .d_arr_1__30 (
              d_arr_relu_1__30), .d_arr_1__29 (d_arr_relu_1__29), .d_arr_1__28 (
              d_arr_relu_1__28), .d_arr_1__27 (d_arr_relu_1__27), .d_arr_1__26 (
              d_arr_relu_1__26), .d_arr_1__25 (d_arr_relu_1__25), .d_arr_1__24 (
              d_arr_relu_1__24), .d_arr_1__23 (d_arr_relu_1__23), .d_arr_1__22 (
              d_arr_relu_1__22), .d_arr_1__21 (d_arr_relu_1__21), .d_arr_1__20 (
              d_arr_relu_1__20), .d_arr_1__19 (d_arr_relu_1__19), .d_arr_1__18 (
              d_arr_relu_1__18), .d_arr_1__17 (d_arr_relu_1__17), .d_arr_1__16 (
              d_arr_relu_1__16), .d_arr_1__15 (\$dummy [1953]), .d_arr_1__14 (
              d_arr_relu_1__14), .d_arr_1__13 (d_arr_relu_1__13), .d_arr_1__12 (
              d_arr_relu_1__12), .d_arr_1__11 (d_arr_relu_1__11), .d_arr_1__10 (
              d_arr_relu_1__10), .d_arr_1__9 (d_arr_relu_1__9), .d_arr_1__8 (
              d_arr_relu_1__8), .d_arr_1__7 (d_arr_relu_1__7), .d_arr_1__6 (
              d_arr_relu_1__6), .d_arr_1__5 (d_arr_relu_1__5), .d_arr_1__4 (
              d_arr_relu_1__4), .d_arr_1__3 (d_arr_relu_1__3), .d_arr_1__2 (
              d_arr_relu_1__2), .d_arr_1__1 (d_arr_relu_1__1), .d_arr_1__0 (
              d_arr_relu_1__0), .d_arr_2__31 (\$dummy [1954]), .d_arr_2__30 (
              \$dummy [1955]), .d_arr_2__29 (\$dummy [1956]), .d_arr_2__28 (
              \$dummy [1957]), .d_arr_2__27 (\$dummy [1958]), .d_arr_2__26 (
              \$dummy [1959]), .d_arr_2__25 (\$dummy [1960]), .d_arr_2__24 (
              \$dummy [1961]), .d_arr_2__23 (\$dummy [1962]), .d_arr_2__22 (
              \$dummy [1963]), .d_arr_2__21 (\$dummy [1964]), .d_arr_2__20 (
              \$dummy [1965]), .d_arr_2__19 (\$dummy [1966]), .d_arr_2__18 (
              \$dummy [1967]), .d_arr_2__17 (\$dummy [1968]), .d_arr_2__16 (
              \$dummy [1969]), .d_arr_2__15 (\$dummy [1970]), .d_arr_2__14 (
              \$dummy [1971]), .d_arr_2__13 (\$dummy [1972]), .d_arr_2__12 (
              \$dummy [1973]), .d_arr_2__11 (\$dummy [1974]), .d_arr_2__10 (
              \$dummy [1975]), .d_arr_2__9 (\$dummy [1976]), .d_arr_2__8 (
              \$dummy [1977]), .d_arr_2__7 (\$dummy [1978]), .d_arr_2__6 (
              \$dummy [1979]), .d_arr_2__5 (\$dummy [1980]), .d_arr_2__4 (
              \$dummy [1981]), .d_arr_2__3 (\$dummy [1982]), .d_arr_2__2 (
              \$dummy [1983]), .d_arr_2__1 (\$dummy [1984]), .d_arr_2__0 (
              \$dummy [1985]), .d_arr_3__31 (\$dummy [1986]), .d_arr_3__30 (
              \$dummy [1987]), .d_arr_3__29 (\$dummy [1988]), .d_arr_3__28 (
              \$dummy [1989]), .d_arr_3__27 (\$dummy [1990]), .d_arr_3__26 (
              \$dummy [1991]), .d_arr_3__25 (\$dummy [1992]), .d_arr_3__24 (
              \$dummy [1993]), .d_arr_3__23 (\$dummy [1994]), .d_arr_3__22 (
              \$dummy [1995]), .d_arr_3__21 (\$dummy [1996]), .d_arr_3__20 (
              \$dummy [1997]), .d_arr_3__19 (\$dummy [1998]), .d_arr_3__18 (
              \$dummy [1999]), .d_arr_3__17 (\$dummy [2000]), .d_arr_3__16 (
              \$dummy [2001]), .d_arr_3__15 (\$dummy [2002]), .d_arr_3__14 (
              \$dummy [2003]), .d_arr_3__13 (\$dummy [2004]), .d_arr_3__12 (
              \$dummy [2005]), .d_arr_3__11 (\$dummy [2006]), .d_arr_3__10 (
              \$dummy [2007]), .d_arr_3__9 (\$dummy [2008]), .d_arr_3__8 (
              \$dummy [2009]), .d_arr_3__7 (\$dummy [2010]), .d_arr_3__6 (
              \$dummy [2011]), .d_arr_3__5 (\$dummy [2012]), .d_arr_3__4 (
              \$dummy [2013]), .d_arr_3__3 (\$dummy [2014]), .d_arr_3__2 (
              \$dummy [2015]), .d_arr_3__1 (\$dummy [2016]), .d_arr_3__0 (
              \$dummy [2017]), .d_arr_4__31 (\$dummy [2018]), .d_arr_4__30 (
              \$dummy [2019]), .d_arr_4__29 (\$dummy [2020]), .d_arr_4__28 (
              \$dummy [2021]), .d_arr_4__27 (\$dummy [2022]), .d_arr_4__26 (
              \$dummy [2023]), .d_arr_4__25 (\$dummy [2024]), .d_arr_4__24 (
              \$dummy [2025]), .d_arr_4__23 (\$dummy [2026]), .d_arr_4__22 (
              \$dummy [2027]), .d_arr_4__21 (\$dummy [2028]), .d_arr_4__20 (
              \$dummy [2029]), .d_arr_4__19 (\$dummy [2030]), .d_arr_4__18 (
              \$dummy [2031]), .d_arr_4__17 (\$dummy [2032]), .d_arr_4__16 (
              \$dummy [2033]), .d_arr_4__15 (\$dummy [2034]), .d_arr_4__14 (
              \$dummy [2035]), .d_arr_4__13 (\$dummy [2036]), .d_arr_4__12 (
              \$dummy [2037]), .d_arr_4__11 (\$dummy [2038]), .d_arr_4__10 (
              \$dummy [2039]), .d_arr_4__9 (\$dummy [2040]), .d_arr_4__8 (
              \$dummy [2041]), .d_arr_4__7 (\$dummy [2042]), .d_arr_4__6 (
              \$dummy [2043]), .d_arr_4__5 (\$dummy [2044]), .d_arr_4__4 (
              \$dummy [2045]), .d_arr_4__3 (\$dummy [2046]), .d_arr_4__2 (
              \$dummy [2047]), .d_arr_4__1 (\$dummy [2048]), .d_arr_4__0 (
              \$dummy [2049]), .d_arr_5__31 (\$dummy [2050]), .d_arr_5__30 (
              \$dummy [2051]), .d_arr_5__29 (\$dummy [2052]), .d_arr_5__28 (
              \$dummy [2053]), .d_arr_5__27 (\$dummy [2054]), .d_arr_5__26 (
              \$dummy [2055]), .d_arr_5__25 (\$dummy [2056]), .d_arr_5__24 (
              \$dummy [2057]), .d_arr_5__23 (\$dummy [2058]), .d_arr_5__22 (
              \$dummy [2059]), .d_arr_5__21 (\$dummy [2060]), .d_arr_5__20 (
              \$dummy [2061]), .d_arr_5__19 (\$dummy [2062]), .d_arr_5__18 (
              \$dummy [2063]), .d_arr_5__17 (\$dummy [2064]), .d_arr_5__16 (
              \$dummy [2065]), .d_arr_5__15 (\$dummy [2066]), .d_arr_5__14 (
              \$dummy [2067]), .d_arr_5__13 (\$dummy [2068]), .d_arr_5__12 (
              \$dummy [2069]), .d_arr_5__11 (\$dummy [2070]), .d_arr_5__10 (
              \$dummy [2071]), .d_arr_5__9 (\$dummy [2072]), .d_arr_5__8 (
              \$dummy [2073]), .d_arr_5__7 (\$dummy [2074]), .d_arr_5__6 (
              \$dummy [2075]), .d_arr_5__5 (\$dummy [2076]), .d_arr_5__4 (
              \$dummy [2077]), .d_arr_5__3 (\$dummy [2078]), .d_arr_5__2 (
              \$dummy [2079]), .d_arr_5__1 (\$dummy [2080]), .d_arr_5__0 (
              \$dummy [2081]), .d_arr_6__31 (\$dummy [2082]), .d_arr_6__30 (
              \$dummy [2083]), .d_arr_6__29 (\$dummy [2084]), .d_arr_6__28 (
              \$dummy [2085]), .d_arr_6__27 (\$dummy [2086]), .d_arr_6__26 (
              \$dummy [2087]), .d_arr_6__25 (\$dummy [2088]), .d_arr_6__24 (
              \$dummy [2089]), .d_arr_6__23 (\$dummy [2090]), .d_arr_6__22 (
              \$dummy [2091]), .d_arr_6__21 (\$dummy [2092]), .d_arr_6__20 (
              \$dummy [2093]), .d_arr_6__19 (\$dummy [2094]), .d_arr_6__18 (
              \$dummy [2095]), .d_arr_6__17 (\$dummy [2096]), .d_arr_6__16 (
              \$dummy [2097]), .d_arr_6__15 (\$dummy [2098]), .d_arr_6__14 (
              \$dummy [2099]), .d_arr_6__13 (\$dummy [2100]), .d_arr_6__12 (
              \$dummy [2101]), .d_arr_6__11 (\$dummy [2102]), .d_arr_6__10 (
              \$dummy [2103]), .d_arr_6__9 (\$dummy [2104]), .d_arr_6__8 (
              \$dummy [2105]), .d_arr_6__7 (\$dummy [2106]), .d_arr_6__6 (
              \$dummy [2107]), .d_arr_6__5 (\$dummy [2108]), .d_arr_6__4 (
              \$dummy [2109]), .d_arr_6__3 (\$dummy [2110]), .d_arr_6__2 (
              \$dummy [2111]), .d_arr_6__1 (\$dummy [2112]), .d_arr_6__0 (
              \$dummy [2113]), .d_arr_7__31 (\$dummy [2114]), .d_arr_7__30 (
              \$dummy [2115]), .d_arr_7__29 (\$dummy [2116]), .d_arr_7__28 (
              \$dummy [2117]), .d_arr_7__27 (\$dummy [2118]), .d_arr_7__26 (
              \$dummy [2119]), .d_arr_7__25 (\$dummy [2120]), .d_arr_7__24 (
              \$dummy [2121]), .d_arr_7__23 (\$dummy [2122]), .d_arr_7__22 (
              \$dummy [2123]), .d_arr_7__21 (\$dummy [2124]), .d_arr_7__20 (
              \$dummy [2125]), .d_arr_7__19 (\$dummy [2126]), .d_arr_7__18 (
              \$dummy [2127]), .d_arr_7__17 (\$dummy [2128]), .d_arr_7__16 (
              \$dummy [2129]), .d_arr_7__15 (\$dummy [2130]), .d_arr_7__14 (
              \$dummy [2131]), .d_arr_7__13 (\$dummy [2132]), .d_arr_7__12 (
              \$dummy [2133]), .d_arr_7__11 (\$dummy [2134]), .d_arr_7__10 (
              \$dummy [2135]), .d_arr_7__9 (\$dummy [2136]), .d_arr_7__8 (
              \$dummy [2137]), .d_arr_7__7 (\$dummy [2138]), .d_arr_7__6 (
              \$dummy [2139]), .d_arr_7__5 (\$dummy [2140]), .d_arr_7__4 (
              \$dummy [2141]), .d_arr_7__3 (\$dummy [2142]), .d_arr_7__2 (
              \$dummy [2143]), .d_arr_7__1 (\$dummy [2144]), .d_arr_7__0 (
              \$dummy [2145]), .d_arr_8__31 (\$dummy [2146]), .d_arr_8__30 (
              \$dummy [2147]), .d_arr_8__29 (\$dummy [2148]), .d_arr_8__28 (
              \$dummy [2149]), .d_arr_8__27 (\$dummy [2150]), .d_arr_8__26 (
              \$dummy [2151]), .d_arr_8__25 (\$dummy [2152]), .d_arr_8__24 (
              \$dummy [2153]), .d_arr_8__23 (\$dummy [2154]), .d_arr_8__22 (
              \$dummy [2155]), .d_arr_8__21 (\$dummy [2156]), .d_arr_8__20 (
              \$dummy [2157]), .d_arr_8__19 (\$dummy [2158]), .d_arr_8__18 (
              \$dummy [2159]), .d_arr_8__17 (\$dummy [2160]), .d_arr_8__16 (
              \$dummy [2161]), .d_arr_8__15 (\$dummy [2162]), .d_arr_8__14 (
              \$dummy [2163]), .d_arr_8__13 (\$dummy [2164]), .d_arr_8__12 (
              \$dummy [2165]), .d_arr_8__11 (\$dummy [2166]), .d_arr_8__10 (
              \$dummy [2167]), .d_arr_8__9 (\$dummy [2168]), .d_arr_8__8 (
              \$dummy [2169]), .d_arr_8__7 (\$dummy [2170]), .d_arr_8__6 (
              \$dummy [2171]), .d_arr_8__5 (\$dummy [2172]), .d_arr_8__4 (
              \$dummy [2173]), .d_arr_8__3 (\$dummy [2174]), .d_arr_8__2 (
              \$dummy [2175]), .d_arr_8__1 (\$dummy [2176]), .d_arr_8__0 (
              \$dummy [2177]), .d_arr_9__31 (\$dummy [2178]), .d_arr_9__30 (
              \$dummy [2179]), .d_arr_9__29 (\$dummy [2180]), .d_arr_9__28 (
              \$dummy [2181]), .d_arr_9__27 (\$dummy [2182]), .d_arr_9__26 (
              \$dummy [2183]), .d_arr_9__25 (\$dummy [2184]), .d_arr_9__24 (
              \$dummy [2185]), .d_arr_9__23 (\$dummy [2186]), .d_arr_9__22 (
              \$dummy [2187]), .d_arr_9__21 (\$dummy [2188]), .d_arr_9__20 (
              \$dummy [2189]), .d_arr_9__19 (\$dummy [2190]), .d_arr_9__18 (
              \$dummy [2191]), .d_arr_9__17 (\$dummy [2192]), .d_arr_9__16 (
              \$dummy [2193]), .d_arr_9__15 (\$dummy [2194]), .d_arr_9__14 (
              \$dummy [2195]), .d_arr_9__13 (\$dummy [2196]), .d_arr_9__12 (
              \$dummy [2197]), .d_arr_9__11 (\$dummy [2198]), .d_arr_9__10 (
              \$dummy [2199]), .d_arr_9__9 (\$dummy [2200]), .d_arr_9__8 (
              \$dummy [2201]), .d_arr_9__7 (\$dummy [2202]), .d_arr_9__6 (
              \$dummy [2203]), .d_arr_9__5 (\$dummy [2204]), .d_arr_9__4 (
              \$dummy [2205]), .d_arr_9__3 (\$dummy [2206]), .d_arr_9__2 (
              \$dummy [2207]), .d_arr_9__1 (\$dummy [2208]), .d_arr_9__0 (
              \$dummy [2209]), .d_arr_10__31 (\$dummy [2210]), .d_arr_10__30 (
              \$dummy [2211]), .d_arr_10__29 (\$dummy [2212]), .d_arr_10__28 (
              \$dummy [2213]), .d_arr_10__27 (\$dummy [2214]), .d_arr_10__26 (
              \$dummy [2215]), .d_arr_10__25 (\$dummy [2216]), .d_arr_10__24 (
              \$dummy [2217]), .d_arr_10__23 (\$dummy [2218]), .d_arr_10__22 (
              \$dummy [2219]), .d_arr_10__21 (\$dummy [2220]), .d_arr_10__20 (
              \$dummy [2221]), .d_arr_10__19 (\$dummy [2222]), .d_arr_10__18 (
              \$dummy [2223]), .d_arr_10__17 (\$dummy [2224]), .d_arr_10__16 (
              \$dummy [2225]), .d_arr_10__15 (\$dummy [2226]), .d_arr_10__14 (
              \$dummy [2227]), .d_arr_10__13 (\$dummy [2228]), .d_arr_10__12 (
              \$dummy [2229]), .d_arr_10__11 (\$dummy [2230]), .d_arr_10__10 (
              \$dummy [2231]), .d_arr_10__9 (\$dummy [2232]), .d_arr_10__8 (
              \$dummy [2233]), .d_arr_10__7 (\$dummy [2234]), .d_arr_10__6 (
              \$dummy [2235]), .d_arr_10__5 (\$dummy [2236]), .d_arr_10__4 (
              \$dummy [2237]), .d_arr_10__3 (\$dummy [2238]), .d_arr_10__2 (
              \$dummy [2239]), .d_arr_10__1 (\$dummy [2240]), .d_arr_10__0 (
              \$dummy [2241]), .d_arr_11__31 (\$dummy [2242]), .d_arr_11__30 (
              \$dummy [2243]), .d_arr_11__29 (\$dummy [2244]), .d_arr_11__28 (
              \$dummy [2245]), .d_arr_11__27 (\$dummy [2246]), .d_arr_11__26 (
              \$dummy [2247]), .d_arr_11__25 (\$dummy [2248]), .d_arr_11__24 (
              \$dummy [2249]), .d_arr_11__23 (\$dummy [2250]), .d_arr_11__22 (
              \$dummy [2251]), .d_arr_11__21 (\$dummy [2252]), .d_arr_11__20 (
              \$dummy [2253]), .d_arr_11__19 (\$dummy [2254]), .d_arr_11__18 (
              \$dummy [2255]), .d_arr_11__17 (\$dummy [2256]), .d_arr_11__16 (
              \$dummy [2257]), .d_arr_11__15 (\$dummy [2258]), .d_arr_11__14 (
              \$dummy [2259]), .d_arr_11__13 (\$dummy [2260]), .d_arr_11__12 (
              \$dummy [2261]), .d_arr_11__11 (\$dummy [2262]), .d_arr_11__10 (
              \$dummy [2263]), .d_arr_11__9 (\$dummy [2264]), .d_arr_11__8 (
              \$dummy [2265]), .d_arr_11__7 (\$dummy [2266]), .d_arr_11__6 (
              \$dummy [2267]), .d_arr_11__5 (\$dummy [2268]), .d_arr_11__4 (
              \$dummy [2269]), .d_arr_11__3 (\$dummy [2270]), .d_arr_11__2 (
              \$dummy [2271]), .d_arr_11__1 (\$dummy [2272]), .d_arr_11__0 (
              \$dummy [2273]), .d_arr_12__31 (\$dummy [2274]), .d_arr_12__30 (
              \$dummy [2275]), .d_arr_12__29 (\$dummy [2276]), .d_arr_12__28 (
              \$dummy [2277]), .d_arr_12__27 (\$dummy [2278]), .d_arr_12__26 (
              \$dummy [2279]), .d_arr_12__25 (\$dummy [2280]), .d_arr_12__24 (
              \$dummy [2281]), .d_arr_12__23 (\$dummy [2282]), .d_arr_12__22 (
              \$dummy [2283]), .d_arr_12__21 (\$dummy [2284]), .d_arr_12__20 (
              \$dummy [2285]), .d_arr_12__19 (\$dummy [2286]), .d_arr_12__18 (
              \$dummy [2287]), .d_arr_12__17 (\$dummy [2288]), .d_arr_12__16 (
              \$dummy [2289]), .d_arr_12__15 (\$dummy [2290]), .d_arr_12__14 (
              \$dummy [2291]), .d_arr_12__13 (\$dummy [2292]), .d_arr_12__12 (
              \$dummy [2293]), .d_arr_12__11 (\$dummy [2294]), .d_arr_12__10 (
              \$dummy [2295]), .d_arr_12__9 (\$dummy [2296]), .d_arr_12__8 (
              \$dummy [2297]), .d_arr_12__7 (\$dummy [2298]), .d_arr_12__6 (
              \$dummy [2299]), .d_arr_12__5 (\$dummy [2300]), .d_arr_12__4 (
              \$dummy [2301]), .d_arr_12__3 (\$dummy [2302]), .d_arr_12__2 (
              \$dummy [2303]), .d_arr_12__1 (\$dummy [2304]), .d_arr_12__0 (
              \$dummy [2305]), .d_arr_13__31 (\$dummy [2306]), .d_arr_13__30 (
              \$dummy [2307]), .d_arr_13__29 (\$dummy [2308]), .d_arr_13__28 (
              \$dummy [2309]), .d_arr_13__27 (\$dummy [2310]), .d_arr_13__26 (
              \$dummy [2311]), .d_arr_13__25 (\$dummy [2312]), .d_arr_13__24 (
              \$dummy [2313]), .d_arr_13__23 (\$dummy [2314]), .d_arr_13__22 (
              \$dummy [2315]), .d_arr_13__21 (\$dummy [2316]), .d_arr_13__20 (
              \$dummy [2317]), .d_arr_13__19 (\$dummy [2318]), .d_arr_13__18 (
              \$dummy [2319]), .d_arr_13__17 (\$dummy [2320]), .d_arr_13__16 (
              \$dummy [2321]), .d_arr_13__15 (\$dummy [2322]), .d_arr_13__14 (
              \$dummy [2323]), .d_arr_13__13 (\$dummy [2324]), .d_arr_13__12 (
              \$dummy [2325]), .d_arr_13__11 (\$dummy [2326]), .d_arr_13__10 (
              \$dummy [2327]), .d_arr_13__9 (\$dummy [2328]), .d_arr_13__8 (
              \$dummy [2329]), .d_arr_13__7 (\$dummy [2330]), .d_arr_13__6 (
              \$dummy [2331]), .d_arr_13__5 (\$dummy [2332]), .d_arr_13__4 (
              \$dummy [2333]), .d_arr_13__3 (\$dummy [2334]), .d_arr_13__2 (
              \$dummy [2335]), .d_arr_13__1 (\$dummy [2336]), .d_arr_13__0 (
              \$dummy [2337]), .d_arr_14__31 (\$dummy [2338]), .d_arr_14__30 (
              \$dummy [2339]), .d_arr_14__29 (\$dummy [2340]), .d_arr_14__28 (
              \$dummy [2341]), .d_arr_14__27 (\$dummy [2342]), .d_arr_14__26 (
              \$dummy [2343]), .d_arr_14__25 (\$dummy [2344]), .d_arr_14__24 (
              \$dummy [2345]), .d_arr_14__23 (\$dummy [2346]), .d_arr_14__22 (
              \$dummy [2347]), .d_arr_14__21 (\$dummy [2348]), .d_arr_14__20 (
              \$dummy [2349]), .d_arr_14__19 (\$dummy [2350]), .d_arr_14__18 (
              \$dummy [2351]), .d_arr_14__17 (\$dummy [2352]), .d_arr_14__16 (
              \$dummy [2353]), .d_arr_14__15 (\$dummy [2354]), .d_arr_14__14 (
              \$dummy [2355]), .d_arr_14__13 (\$dummy [2356]), .d_arr_14__12 (
              \$dummy [2357]), .d_arr_14__11 (\$dummy [2358]), .d_arr_14__10 (
              \$dummy [2359]), .d_arr_14__9 (\$dummy [2360]), .d_arr_14__8 (
              \$dummy [2361]), .d_arr_14__7 (\$dummy [2362]), .d_arr_14__6 (
              \$dummy [2363]), .d_arr_14__5 (\$dummy [2364]), .d_arr_14__4 (
              \$dummy [2365]), .d_arr_14__3 (\$dummy [2366]), .d_arr_14__2 (
              \$dummy [2367]), .d_arr_14__1 (\$dummy [2368]), .d_arr_14__0 (
              \$dummy [2369]), .d_arr_15__31 (\$dummy [2370]), .d_arr_15__30 (
              \$dummy [2371]), .d_arr_15__29 (\$dummy [2372]), .d_arr_15__28 (
              \$dummy [2373]), .d_arr_15__27 (\$dummy [2374]), .d_arr_15__26 (
              \$dummy [2375]), .d_arr_15__25 (\$dummy [2376]), .d_arr_15__24 (
              \$dummy [2377]), .d_arr_15__23 (\$dummy [2378]), .d_arr_15__22 (
              \$dummy [2379]), .d_arr_15__21 (\$dummy [2380]), .d_arr_15__20 (
              \$dummy [2381]), .d_arr_15__19 (\$dummy [2382]), .d_arr_15__18 (
              \$dummy [2383]), .d_arr_15__17 (\$dummy [2384]), .d_arr_15__16 (
              \$dummy [2385]), .d_arr_15__15 (\$dummy [2386]), .d_arr_15__14 (
              \$dummy [2387]), .d_arr_15__13 (\$dummy [2388]), .d_arr_15__12 (
              \$dummy [2389]), .d_arr_15__11 (\$dummy [2390]), .d_arr_15__10 (
              \$dummy [2391]), .d_arr_15__9 (\$dummy [2392]), .d_arr_15__8 (
              \$dummy [2393]), .d_arr_15__7 (\$dummy [2394]), .d_arr_15__6 (
              \$dummy [2395]), .d_arr_15__5 (\$dummy [2396]), .d_arr_15__4 (
              \$dummy [2397]), .d_arr_15__3 (\$dummy [2398]), .d_arr_15__2 (
              \$dummy [2399]), .d_arr_15__1 (\$dummy [2400]), .d_arr_15__0 (
              \$dummy [2401]), .d_arr_16__31 (\$dummy [2402]), .d_arr_16__30 (
              \$dummy [2403]), .d_arr_16__29 (\$dummy [2404]), .d_arr_16__28 (
              \$dummy [2405]), .d_arr_16__27 (\$dummy [2406]), .d_arr_16__26 (
              \$dummy [2407]), .d_arr_16__25 (\$dummy [2408]), .d_arr_16__24 (
              \$dummy [2409]), .d_arr_16__23 (\$dummy [2410]), .d_arr_16__22 (
              \$dummy [2411]), .d_arr_16__21 (\$dummy [2412]), .d_arr_16__20 (
              \$dummy [2413]), .d_arr_16__19 (\$dummy [2414]), .d_arr_16__18 (
              \$dummy [2415]), .d_arr_16__17 (\$dummy [2416]), .d_arr_16__16 (
              \$dummy [2417]), .d_arr_16__15 (\$dummy [2418]), .d_arr_16__14 (
              \$dummy [2419]), .d_arr_16__13 (\$dummy [2420]), .d_arr_16__12 (
              \$dummy [2421]), .d_arr_16__11 (\$dummy [2422]), .d_arr_16__10 (
              \$dummy [2423]), .d_arr_16__9 (\$dummy [2424]), .d_arr_16__8 (
              \$dummy [2425]), .d_arr_16__7 (\$dummy [2426]), .d_arr_16__6 (
              \$dummy [2427]), .d_arr_16__5 (\$dummy [2428]), .d_arr_16__4 (
              \$dummy [2429]), .d_arr_16__3 (\$dummy [2430]), .d_arr_16__2 (
              \$dummy [2431]), .d_arr_16__1 (\$dummy [2432]), .d_arr_16__0 (
              \$dummy [2433]), .d_arr_17__31 (\$dummy [2434]), .d_arr_17__30 (
              \$dummy [2435]), .d_arr_17__29 (\$dummy [2436]), .d_arr_17__28 (
              \$dummy [2437]), .d_arr_17__27 (\$dummy [2438]), .d_arr_17__26 (
              \$dummy [2439]), .d_arr_17__25 (\$dummy [2440]), .d_arr_17__24 (
              \$dummy [2441]), .d_arr_17__23 (\$dummy [2442]), .d_arr_17__22 (
              \$dummy [2443]), .d_arr_17__21 (\$dummy [2444]), .d_arr_17__20 (
              \$dummy [2445]), .d_arr_17__19 (\$dummy [2446]), .d_arr_17__18 (
              \$dummy [2447]), .d_arr_17__17 (\$dummy [2448]), .d_arr_17__16 (
              \$dummy [2449]), .d_arr_17__15 (\$dummy [2450]), .d_arr_17__14 (
              \$dummy [2451]), .d_arr_17__13 (\$dummy [2452]), .d_arr_17__12 (
              \$dummy [2453]), .d_arr_17__11 (\$dummy [2454]), .d_arr_17__10 (
              \$dummy [2455]), .d_arr_17__9 (\$dummy [2456]), .d_arr_17__8 (
              \$dummy [2457]), .d_arr_17__7 (\$dummy [2458]), .d_arr_17__6 (
              \$dummy [2459]), .d_arr_17__5 (\$dummy [2460]), .d_arr_17__4 (
              \$dummy [2461]), .d_arr_17__3 (\$dummy [2462]), .d_arr_17__2 (
              \$dummy [2463]), .d_arr_17__1 (\$dummy [2464]), .d_arr_17__0 (
              \$dummy [2465]), .d_arr_18__31 (\$dummy [2466]), .d_arr_18__30 (
              \$dummy [2467]), .d_arr_18__29 (\$dummy [2468]), .d_arr_18__28 (
              \$dummy [2469]), .d_arr_18__27 (\$dummy [2470]), .d_arr_18__26 (
              \$dummy [2471]), .d_arr_18__25 (\$dummy [2472]), .d_arr_18__24 (
              \$dummy [2473]), .d_arr_18__23 (\$dummy [2474]), .d_arr_18__22 (
              \$dummy [2475]), .d_arr_18__21 (\$dummy [2476]), .d_arr_18__20 (
              \$dummy [2477]), .d_arr_18__19 (\$dummy [2478]), .d_arr_18__18 (
              \$dummy [2479]), .d_arr_18__17 (\$dummy [2480]), .d_arr_18__16 (
              \$dummy [2481]), .d_arr_18__15 (\$dummy [2482]), .d_arr_18__14 (
              \$dummy [2483]), .d_arr_18__13 (\$dummy [2484]), .d_arr_18__12 (
              \$dummy [2485]), .d_arr_18__11 (\$dummy [2486]), .d_arr_18__10 (
              \$dummy [2487]), .d_arr_18__9 (\$dummy [2488]), .d_arr_18__8 (
              \$dummy [2489]), .d_arr_18__7 (\$dummy [2490]), .d_arr_18__6 (
              \$dummy [2491]), .d_arr_18__5 (\$dummy [2492]), .d_arr_18__4 (
              \$dummy [2493]), .d_arr_18__3 (\$dummy [2494]), .d_arr_18__2 (
              \$dummy [2495]), .d_arr_18__1 (\$dummy [2496]), .d_arr_18__0 (
              \$dummy [2497]), .d_arr_19__31 (\$dummy [2498]), .d_arr_19__30 (
              \$dummy [2499]), .d_arr_19__29 (\$dummy [2500]), .d_arr_19__28 (
              \$dummy [2501]), .d_arr_19__27 (\$dummy [2502]), .d_arr_19__26 (
              \$dummy [2503]), .d_arr_19__25 (\$dummy [2504]), .d_arr_19__24 (
              \$dummy [2505]), .d_arr_19__23 (\$dummy [2506]), .d_arr_19__22 (
              \$dummy [2507]), .d_arr_19__21 (\$dummy [2508]), .d_arr_19__20 (
              \$dummy [2509]), .d_arr_19__19 (\$dummy [2510]), .d_arr_19__18 (
              \$dummy [2511]), .d_arr_19__17 (\$dummy [2512]), .d_arr_19__16 (
              \$dummy [2513]), .d_arr_19__15 (\$dummy [2514]), .d_arr_19__14 (
              \$dummy [2515]), .d_arr_19__13 (\$dummy [2516]), .d_arr_19__12 (
              \$dummy [2517]), .d_arr_19__11 (\$dummy [2518]), .d_arr_19__10 (
              \$dummy [2519]), .d_arr_19__9 (\$dummy [2520]), .d_arr_19__8 (
              \$dummy [2521]), .d_arr_19__7 (\$dummy [2522]), .d_arr_19__6 (
              \$dummy [2523]), .d_arr_19__5 (\$dummy [2524]), .d_arr_19__4 (
              \$dummy [2525]), .d_arr_19__3 (\$dummy [2526]), .d_arr_19__2 (
              \$dummy [2527]), .d_arr_19__1 (\$dummy [2528]), .d_arr_19__0 (
              \$dummy [2529]), .d_arr_20__31 (\$dummy [2530]), .d_arr_20__30 (
              \$dummy [2531]), .d_arr_20__29 (\$dummy [2532]), .d_arr_20__28 (
              \$dummy [2533]), .d_arr_20__27 (\$dummy [2534]), .d_arr_20__26 (
              \$dummy [2535]), .d_arr_20__25 (\$dummy [2536]), .d_arr_20__24 (
              \$dummy [2537]), .d_arr_20__23 (\$dummy [2538]), .d_arr_20__22 (
              \$dummy [2539]), .d_arr_20__21 (\$dummy [2540]), .d_arr_20__20 (
              \$dummy [2541]), .d_arr_20__19 (\$dummy [2542]), .d_arr_20__18 (
              \$dummy [2543]), .d_arr_20__17 (\$dummy [2544]), .d_arr_20__16 (
              \$dummy [2545]), .d_arr_20__15 (\$dummy [2546]), .d_arr_20__14 (
              \$dummy [2547]), .d_arr_20__13 (\$dummy [2548]), .d_arr_20__12 (
              \$dummy [2549]), .d_arr_20__11 (\$dummy [2550]), .d_arr_20__10 (
              \$dummy [2551]), .d_arr_20__9 (\$dummy [2552]), .d_arr_20__8 (
              \$dummy [2553]), .d_arr_20__7 (\$dummy [2554]), .d_arr_20__6 (
              \$dummy [2555]), .d_arr_20__5 (\$dummy [2556]), .d_arr_20__4 (
              \$dummy [2557]), .d_arr_20__3 (\$dummy [2558]), .d_arr_20__2 (
              \$dummy [2559]), .d_arr_20__1 (\$dummy [2560]), .d_arr_20__0 (
              \$dummy [2561]), .d_arr_21__31 (\$dummy [2562]), .d_arr_21__30 (
              \$dummy [2563]), .d_arr_21__29 (\$dummy [2564]), .d_arr_21__28 (
              \$dummy [2565]), .d_arr_21__27 (\$dummy [2566]), .d_arr_21__26 (
              \$dummy [2567]), .d_arr_21__25 (\$dummy [2568]), .d_arr_21__24 (
              \$dummy [2569]), .d_arr_21__23 (\$dummy [2570]), .d_arr_21__22 (
              \$dummy [2571]), .d_arr_21__21 (\$dummy [2572]), .d_arr_21__20 (
              \$dummy [2573]), .d_arr_21__19 (\$dummy [2574]), .d_arr_21__18 (
              \$dummy [2575]), .d_arr_21__17 (\$dummy [2576]), .d_arr_21__16 (
              \$dummy [2577]), .d_arr_21__15 (\$dummy [2578]), .d_arr_21__14 (
              \$dummy [2579]), .d_arr_21__13 (\$dummy [2580]), .d_arr_21__12 (
              \$dummy [2581]), .d_arr_21__11 (\$dummy [2582]), .d_arr_21__10 (
              \$dummy [2583]), .d_arr_21__9 (\$dummy [2584]), .d_arr_21__8 (
              \$dummy [2585]), .d_arr_21__7 (\$dummy [2586]), .d_arr_21__6 (
              \$dummy [2587]), .d_arr_21__5 (\$dummy [2588]), .d_arr_21__4 (
              \$dummy [2589]), .d_arr_21__3 (\$dummy [2590]), .d_arr_21__2 (
              \$dummy [2591]), .d_arr_21__1 (\$dummy [2592]), .d_arr_21__0 (
              \$dummy [2593]), .d_arr_22__31 (\$dummy [2594]), .d_arr_22__30 (
              \$dummy [2595]), .d_arr_22__29 (\$dummy [2596]), .d_arr_22__28 (
              \$dummy [2597]), .d_arr_22__27 (\$dummy [2598]), .d_arr_22__26 (
              \$dummy [2599]), .d_arr_22__25 (\$dummy [2600]), .d_arr_22__24 (
              \$dummy [2601]), .d_arr_22__23 (\$dummy [2602]), .d_arr_22__22 (
              \$dummy [2603]), .d_arr_22__21 (\$dummy [2604]), .d_arr_22__20 (
              \$dummy [2605]), .d_arr_22__19 (\$dummy [2606]), .d_arr_22__18 (
              \$dummy [2607]), .d_arr_22__17 (\$dummy [2608]), .d_arr_22__16 (
              \$dummy [2609]), .d_arr_22__15 (\$dummy [2610]), .d_arr_22__14 (
              \$dummy [2611]), .d_arr_22__13 (\$dummy [2612]), .d_arr_22__12 (
              \$dummy [2613]), .d_arr_22__11 (\$dummy [2614]), .d_arr_22__10 (
              \$dummy [2615]), .d_arr_22__9 (\$dummy [2616]), .d_arr_22__8 (
              \$dummy [2617]), .d_arr_22__7 (\$dummy [2618]), .d_arr_22__6 (
              \$dummy [2619]), .d_arr_22__5 (\$dummy [2620]), .d_arr_22__4 (
              \$dummy [2621]), .d_arr_22__3 (\$dummy [2622]), .d_arr_22__2 (
              \$dummy [2623]), .d_arr_22__1 (\$dummy [2624]), .d_arr_22__0 (
              \$dummy [2625]), .d_arr_23__31 (\$dummy [2626]), .d_arr_23__30 (
              \$dummy [2627]), .d_arr_23__29 (\$dummy [2628]), .d_arr_23__28 (
              \$dummy [2629]), .d_arr_23__27 (\$dummy [2630]), .d_arr_23__26 (
              \$dummy [2631]), .d_arr_23__25 (\$dummy [2632]), .d_arr_23__24 (
              \$dummy [2633]), .d_arr_23__23 (\$dummy [2634]), .d_arr_23__22 (
              \$dummy [2635]), .d_arr_23__21 (\$dummy [2636]), .d_arr_23__20 (
              \$dummy [2637]), .d_arr_23__19 (\$dummy [2638]), .d_arr_23__18 (
              \$dummy [2639]), .d_arr_23__17 (\$dummy [2640]), .d_arr_23__16 (
              \$dummy [2641]), .d_arr_23__15 (\$dummy [2642]), .d_arr_23__14 (
              \$dummy [2643]), .d_arr_23__13 (\$dummy [2644]), .d_arr_23__12 (
              \$dummy [2645]), .d_arr_23__11 (\$dummy [2646]), .d_arr_23__10 (
              \$dummy [2647]), .d_arr_23__9 (\$dummy [2648]), .d_arr_23__8 (
              \$dummy [2649]), .d_arr_23__7 (\$dummy [2650]), .d_arr_23__6 (
              \$dummy [2651]), .d_arr_23__5 (\$dummy [2652]), .d_arr_23__4 (
              \$dummy [2653]), .d_arr_23__3 (\$dummy [2654]), .d_arr_23__2 (
              \$dummy [2655]), .d_arr_23__1 (\$dummy [2656]), .d_arr_23__0 (
              \$dummy [2657]), .d_arr_24__31 (\$dummy [2658]), .d_arr_24__30 (
              \$dummy [2659]), .d_arr_24__29 (\$dummy [2660]), .d_arr_24__28 (
              \$dummy [2661]), .d_arr_24__27 (\$dummy [2662]), .d_arr_24__26 (
              \$dummy [2663]), .d_arr_24__25 (\$dummy [2664]), .d_arr_24__24 (
              \$dummy [2665]), .d_arr_24__23 (\$dummy [2666]), .d_arr_24__22 (
              \$dummy [2667]), .d_arr_24__21 (\$dummy [2668]), .d_arr_24__20 (
              \$dummy [2669]), .d_arr_24__19 (\$dummy [2670]), .d_arr_24__18 (
              \$dummy [2671]), .d_arr_24__17 (\$dummy [2672]), .d_arr_24__16 (
              \$dummy [2673]), .d_arr_24__15 (\$dummy [2674]), .d_arr_24__14 (
              \$dummy [2675]), .d_arr_24__13 (\$dummy [2676]), .d_arr_24__12 (
              \$dummy [2677]), .d_arr_24__11 (\$dummy [2678]), .d_arr_24__10 (
              \$dummy [2679]), .d_arr_24__9 (\$dummy [2680]), .d_arr_24__8 (
              \$dummy [2681]), .d_arr_24__7 (\$dummy [2682]), .d_arr_24__6 (
              \$dummy [2683]), .d_arr_24__5 (\$dummy [2684]), .d_arr_24__4 (
              \$dummy [2685]), .d_arr_24__3 (\$dummy [2686]), .d_arr_24__2 (
              \$dummy [2687]), .d_arr_24__1 (\$dummy [2688]), .d_arr_24__0 (
              \$dummy [2689]), .q_arr_0__31 (nx19448), .q_arr_0__30 (nx16499), .q_arr_0__29 (
              nx16503), .q_arr_0__28 (nx16507), .q_arr_0__27 (nx16511), .q_arr_0__26 (
              nx16515), .q_arr_0__25 (nx16519), .q_arr_0__24 (nx19390), .q_arr_0__23 (
              nx16527), .q_arr_0__22 (nx16531), .q_arr_0__21 (nx16535), .q_arr_0__20 (
              nx16539), .q_arr_0__19 (nx16543), .q_arr_0__18 (nx16547), .q_arr_0__17 (
              nx16551), .q_arr_0__16 (nx16555), .q_arr_0__15 (nx16559), .q_arr_0__14 (
              nx16563), .q_arr_0__13 (nx16567), .q_arr_0__12 (nx16571), .q_arr_0__11 (
              nx16575), .q_arr_0__10 (nx16579), .q_arr_0__9 (nx16583), .q_arr_0__8 (
              nx16587), .q_arr_0__7 (nx16591), .q_arr_0__6 (nx16595), .q_arr_0__5 (
              nx16599), .q_arr_0__4 (nx16601), .q_arr_0__3 (nx16603), .q_arr_0__2 (
              q_arr_0__2), .q_arr_0__1 (q_arr_0__1), .q_arr_0__0 (nx16605), .q_arr_1__31 (
              q_arr_1__31), .q_arr_1__30 (q_arr_1__30), .q_arr_1__29 (
              q_arr_1__29), .q_arr_1__28 (q_arr_1__28), .q_arr_1__27 (nx19450), 
              .q_arr_1__26 (nx19454), .q_arr_1__25 (q_arr_1__25), .q_arr_1__24 (
              nx19458), .q_arr_1__23 (q_arr_1__23), .q_arr_1__22 (q_arr_1__22), 
              .q_arr_1__21 (q_arr_1__21), .q_arr_1__20 (q_arr_1__20), .q_arr_1__19 (
              q_arr_1__19), .q_arr_1__18 (nx19462), .q_arr_1__17 (nx19466), .q_arr_1__16 (
              nx19470), .q_arr_1__15 (q_arr_1__15), .q_arr_1__14 (nx19474), .q_arr_1__13 (
              q_arr_1__13), .q_arr_1__12 (nx19476), .q_arr_1__11 (q_arr_1__11), 
              .q_arr_1__10 (nx19478), .q_arr_1__9 (q_arr_1__9), .q_arr_1__8 (
              nx19482), .q_arr_1__7 (nx19486), .q_arr_1__6 (q_arr_1__6), .q_arr_1__5 (
              q_arr_1__5), .q_arr_1__4 (q_arr_1__4), .q_arr_1__3 (q_arr_1__3), .q_arr_1__2 (
              q_arr_1__2), .q_arr_1__1 (q_arr_1__1), .q_arr_1__0 (q_arr_1__0), .q_arr_2__31 (
              GND0), .q_arr_2__30 (GND0), .q_arr_2__29 (GND0), .q_arr_2__28 (
              GND0), .q_arr_2__27 (GND0), .q_arr_2__26 (GND0), .q_arr_2__25 (
              GND0), .q_arr_2__24 (GND0), .q_arr_2__23 (GND0), .q_arr_2__22 (
              GND0), .q_arr_2__21 (GND0), .q_arr_2__20 (GND0), .q_arr_2__19 (
              GND0), .q_arr_2__18 (GND0), .q_arr_2__17 (GND0), .q_arr_2__16 (
              GND0), .q_arr_2__15 (GND0), .q_arr_2__14 (GND0), .q_arr_2__13 (
              GND0), .q_arr_2__12 (GND0), .q_arr_2__11 (GND0), .q_arr_2__10 (
              GND0), .q_arr_2__9 (GND0), .q_arr_2__8 (GND0), .q_arr_2__7 (GND0)
              , .q_arr_2__6 (GND0), .q_arr_2__5 (GND0), .q_arr_2__4 (GND0), .q_arr_2__3 (
              GND0), .q_arr_2__2 (GND0), .q_arr_2__1 (GND0), .q_arr_2__0 (GND0)
              , .q_arr_3__31 (GND0), .q_arr_3__30 (GND0), .q_arr_3__29 (GND0), .q_arr_3__28 (
              GND0), .q_arr_3__27 (GND0), .q_arr_3__26 (GND0), .q_arr_3__25 (
              GND0), .q_arr_3__24 (GND0), .q_arr_3__23 (GND0), .q_arr_3__22 (
              GND0), .q_arr_3__21 (GND0), .q_arr_3__20 (GND0), .q_arr_3__19 (
              GND0), .q_arr_3__18 (GND0), .q_arr_3__17 (GND0), .q_arr_3__16 (
              GND0), .q_arr_3__15 (GND0), .q_arr_3__14 (GND0), .q_arr_3__13 (
              GND0), .q_arr_3__12 (GND0), .q_arr_3__11 (GND0), .q_arr_3__10 (
              GND0), .q_arr_3__9 (GND0), .q_arr_3__8 (GND0), .q_arr_3__7 (GND0)
              , .q_arr_3__6 (GND0), .q_arr_3__5 (GND0), .q_arr_3__4 (GND0), .q_arr_3__3 (
              GND0), .q_arr_3__2 (GND0), .q_arr_3__1 (GND0), .q_arr_3__0 (GND0)
              , .q_arr_4__31 (GND0), .q_arr_4__30 (GND0), .q_arr_4__29 (GND0), .q_arr_4__28 (
              GND0), .q_arr_4__27 (GND0), .q_arr_4__26 (GND0), .q_arr_4__25 (
              GND0), .q_arr_4__24 (GND0), .q_arr_4__23 (GND0), .q_arr_4__22 (
              GND0), .q_arr_4__21 (GND0), .q_arr_4__20 (GND0), .q_arr_4__19 (
              GND0), .q_arr_4__18 (GND0), .q_arr_4__17 (GND0), .q_arr_4__16 (
              GND0), .q_arr_4__15 (GND0), .q_arr_4__14 (GND0), .q_arr_4__13 (
              GND0), .q_arr_4__12 (GND0), .q_arr_4__11 (GND0), .q_arr_4__10 (
              GND0), .q_arr_4__9 (GND0), .q_arr_4__8 (GND0), .q_arr_4__7 (GND0)
              , .q_arr_4__6 (GND0), .q_arr_4__5 (GND0), .q_arr_4__4 (GND0), .q_arr_4__3 (
              GND0), .q_arr_4__2 (GND0), .q_arr_4__1 (GND0), .q_arr_4__0 (GND0)
              , .q_arr_5__31 (GND0), .q_arr_5__30 (GND0), .q_arr_5__29 (GND0), .q_arr_5__28 (
              GND0), .q_arr_5__27 (GND0), .q_arr_5__26 (GND0), .q_arr_5__25 (
              GND0), .q_arr_5__24 (GND0), .q_arr_5__23 (GND0), .q_arr_5__22 (
              GND0), .q_arr_5__21 (GND0), .q_arr_5__20 (GND0), .q_arr_5__19 (
              GND0), .q_arr_5__18 (GND0), .q_arr_5__17 (GND0), .q_arr_5__16 (
              GND0), .q_arr_5__15 (GND0), .q_arr_5__14 (GND0), .q_arr_5__13 (
              GND0), .q_arr_5__12 (GND0), .q_arr_5__11 (GND0), .q_arr_5__10 (
              GND0), .q_arr_5__9 (GND0), .q_arr_5__8 (GND0), .q_arr_5__7 (GND0)
              , .q_arr_5__6 (GND0), .q_arr_5__5 (GND0), .q_arr_5__4 (GND0), .q_arr_5__3 (
              GND0), .q_arr_5__2 (GND0), .q_arr_5__1 (GND0), .q_arr_5__0 (GND0)
              , .q_arr_6__31 (GND0), .q_arr_6__30 (GND0), .q_arr_6__29 (GND0), .q_arr_6__28 (
              GND0), .q_arr_6__27 (GND0), .q_arr_6__26 (GND0), .q_arr_6__25 (
              GND0), .q_arr_6__24 (GND0), .q_arr_6__23 (GND0), .q_arr_6__22 (
              GND0), .q_arr_6__21 (GND0), .q_arr_6__20 (GND0), .q_arr_6__19 (
              GND0), .q_arr_6__18 (GND0), .q_arr_6__17 (GND0), .q_arr_6__16 (
              GND0), .q_arr_6__15 (GND0), .q_arr_6__14 (GND0), .q_arr_6__13 (
              GND0), .q_arr_6__12 (GND0), .q_arr_6__11 (GND0), .q_arr_6__10 (
              GND0), .q_arr_6__9 (GND0), .q_arr_6__8 (GND0), .q_arr_6__7 (GND0)
              , .q_arr_6__6 (GND0), .q_arr_6__5 (GND0), .q_arr_6__4 (GND0), .q_arr_6__3 (
              GND0), .q_arr_6__2 (GND0), .q_arr_6__1 (GND0), .q_arr_6__0 (GND0)
              , .q_arr_7__31 (GND0), .q_arr_7__30 (GND0), .q_arr_7__29 (GND0), .q_arr_7__28 (
              GND0), .q_arr_7__27 (GND0), .q_arr_7__26 (GND0), .q_arr_7__25 (
              GND0), .q_arr_7__24 (GND0), .q_arr_7__23 (GND0), .q_arr_7__22 (
              GND0), .q_arr_7__21 (GND0), .q_arr_7__20 (GND0), .q_arr_7__19 (
              GND0), .q_arr_7__18 (GND0), .q_arr_7__17 (GND0), .q_arr_7__16 (
              GND0), .q_arr_7__15 (GND0), .q_arr_7__14 (GND0), .q_arr_7__13 (
              GND0), .q_arr_7__12 (GND0), .q_arr_7__11 (GND0), .q_arr_7__10 (
              GND0), .q_arr_7__9 (GND0), .q_arr_7__8 (GND0), .q_arr_7__7 (GND0)
              , .q_arr_7__6 (GND0), .q_arr_7__5 (GND0), .q_arr_7__4 (GND0), .q_arr_7__3 (
              GND0), .q_arr_7__2 (GND0), .q_arr_7__1 (GND0), .q_arr_7__0 (GND0)
              , .q_arr_8__31 (GND0), .q_arr_8__30 (GND0), .q_arr_8__29 (GND0), .q_arr_8__28 (
              GND0), .q_arr_8__27 (GND0), .q_arr_8__26 (GND0), .q_arr_8__25 (
              GND0), .q_arr_8__24 (GND0), .q_arr_8__23 (GND0), .q_arr_8__22 (
              GND0), .q_arr_8__21 (GND0), .q_arr_8__20 (GND0), .q_arr_8__19 (
              GND0), .q_arr_8__18 (GND0), .q_arr_8__17 (GND0), .q_arr_8__16 (
              GND0), .q_arr_8__15 (GND0), .q_arr_8__14 (GND0), .q_arr_8__13 (
              GND0), .q_arr_8__12 (GND0), .q_arr_8__11 (GND0), .q_arr_8__10 (
              GND0), .q_arr_8__9 (GND0), .q_arr_8__8 (GND0), .q_arr_8__7 (GND0)
              , .q_arr_8__6 (GND0), .q_arr_8__5 (GND0), .q_arr_8__4 (GND0), .q_arr_8__3 (
              GND0), .q_arr_8__2 (GND0), .q_arr_8__1 (GND0), .q_arr_8__0 (GND0)
              , .q_arr_9__31 (GND0), .q_arr_9__30 (GND0), .q_arr_9__29 (GND0), .q_arr_9__28 (
              GND0), .q_arr_9__27 (GND0), .q_arr_9__26 (GND0), .q_arr_9__25 (
              GND0), .q_arr_9__24 (GND0), .q_arr_9__23 (GND0), .q_arr_9__22 (
              GND0), .q_arr_9__21 (GND0), .q_arr_9__20 (GND0), .q_arr_9__19 (
              GND0), .q_arr_9__18 (GND0), .q_arr_9__17 (GND0), .q_arr_9__16 (
              GND0), .q_arr_9__15 (GND0), .q_arr_9__14 (GND0), .q_arr_9__13 (
              GND0), .q_arr_9__12 (GND0), .q_arr_9__11 (GND0), .q_arr_9__10 (
              GND0), .q_arr_9__9 (GND0), .q_arr_9__8 (GND0), .q_arr_9__7 (GND0)
              , .q_arr_9__6 (GND0), .q_arr_9__5 (GND0), .q_arr_9__4 (GND0), .q_arr_9__3 (
              GND0), .q_arr_9__2 (GND0), .q_arr_9__1 (GND0), .q_arr_9__0 (GND0)
              , .q_arr_10__31 (GND0), .q_arr_10__30 (GND0), .q_arr_10__29 (GND0)
              , .q_arr_10__28 (GND0), .q_arr_10__27 (GND0), .q_arr_10__26 (GND0)
              , .q_arr_10__25 (GND0), .q_arr_10__24 (GND0), .q_arr_10__23 (GND0)
              , .q_arr_10__22 (GND0), .q_arr_10__21 (GND0), .q_arr_10__20 (GND0)
              , .q_arr_10__19 (GND0), .q_arr_10__18 (GND0), .q_arr_10__17 (GND0)
              , .q_arr_10__16 (GND0), .q_arr_10__15 (GND0), .q_arr_10__14 (GND0)
              , .q_arr_10__13 (GND0), .q_arr_10__12 (GND0), .q_arr_10__11 (GND0)
              , .q_arr_10__10 (GND0), .q_arr_10__9 (GND0), .q_arr_10__8 (GND0), 
              .q_arr_10__7 (GND0), .q_arr_10__6 (GND0), .q_arr_10__5 (GND0), .q_arr_10__4 (
              GND0), .q_arr_10__3 (GND0), .q_arr_10__2 (GND0), .q_arr_10__1 (
              GND0), .q_arr_10__0 (GND0), .q_arr_11__31 (GND0), .q_arr_11__30 (
              GND0), .q_arr_11__29 (GND0), .q_arr_11__28 (GND0), .q_arr_11__27 (
              GND0), .q_arr_11__26 (GND0), .q_arr_11__25 (GND0), .q_arr_11__24 (
              GND0), .q_arr_11__23 (GND0), .q_arr_11__22 (GND0), .q_arr_11__21 (
              GND0), .q_arr_11__20 (GND0), .q_arr_11__19 (GND0), .q_arr_11__18 (
              GND0), .q_arr_11__17 (GND0), .q_arr_11__16 (GND0), .q_arr_11__15 (
              GND0), .q_arr_11__14 (GND0), .q_arr_11__13 (GND0), .q_arr_11__12 (
              GND0), .q_arr_11__11 (GND0), .q_arr_11__10 (GND0), .q_arr_11__9 (
              GND0), .q_arr_11__8 (GND0), .q_arr_11__7 (GND0), .q_arr_11__6 (
              GND0), .q_arr_11__5 (GND0), .q_arr_11__4 (GND0), .q_arr_11__3 (
              GND0), .q_arr_11__2 (GND0), .q_arr_11__1 (GND0), .q_arr_11__0 (
              GND0), .q_arr_12__31 (GND0), .q_arr_12__30 (GND0), .q_arr_12__29 (
              GND0), .q_arr_12__28 (GND0), .q_arr_12__27 (GND0), .q_arr_12__26 (
              GND0), .q_arr_12__25 (GND0), .q_arr_12__24 (GND0), .q_arr_12__23 (
              GND0), .q_arr_12__22 (GND0), .q_arr_12__21 (GND0), .q_arr_12__20 (
              GND0), .q_arr_12__19 (GND0), .q_arr_12__18 (GND0), .q_arr_12__17 (
              GND0), .q_arr_12__16 (GND0), .q_arr_12__15 (GND0), .q_arr_12__14 (
              GND0), .q_arr_12__13 (GND0), .q_arr_12__12 (GND0), .q_arr_12__11 (
              GND0), .q_arr_12__10 (GND0), .q_arr_12__9 (GND0), .q_arr_12__8 (
              GND0), .q_arr_12__7 (GND0), .q_arr_12__6 (GND0), .q_arr_12__5 (
              GND0), .q_arr_12__4 (GND0), .q_arr_12__3 (GND0), .q_arr_12__2 (
              GND0), .q_arr_12__1 (GND0), .q_arr_12__0 (GND0), .q_arr_13__31 (
              GND0), .q_arr_13__30 (GND0), .q_arr_13__29 (GND0), .q_arr_13__28 (
              GND0), .q_arr_13__27 (GND0), .q_arr_13__26 (GND0), .q_arr_13__25 (
              GND0), .q_arr_13__24 (GND0), .q_arr_13__23 (GND0), .q_arr_13__22 (
              GND0), .q_arr_13__21 (GND0), .q_arr_13__20 (GND0), .q_arr_13__19 (
              GND0), .q_arr_13__18 (GND0), .q_arr_13__17 (GND0), .q_arr_13__16 (
              GND0), .q_arr_13__15 (GND0), .q_arr_13__14 (GND0), .q_arr_13__13 (
              GND0), .q_arr_13__12 (GND0), .q_arr_13__11 (GND0), .q_arr_13__10 (
              GND0), .q_arr_13__9 (GND0), .q_arr_13__8 (GND0), .q_arr_13__7 (
              GND0), .q_arr_13__6 (GND0), .q_arr_13__5 (GND0), .q_arr_13__4 (
              GND0), .q_arr_13__3 (GND0), .q_arr_13__2 (GND0), .q_arr_13__1 (
              GND0), .q_arr_13__0 (GND0), .q_arr_14__31 (GND0), .q_arr_14__30 (
              GND0), .q_arr_14__29 (GND0), .q_arr_14__28 (GND0), .q_arr_14__27 (
              GND0), .q_arr_14__26 (GND0), .q_arr_14__25 (GND0), .q_arr_14__24 (
              GND0), .q_arr_14__23 (GND0), .q_arr_14__22 (GND0), .q_arr_14__21 (
              GND0), .q_arr_14__20 (GND0), .q_arr_14__19 (GND0), .q_arr_14__18 (
              GND0), .q_arr_14__17 (GND0), .q_arr_14__16 (GND0), .q_arr_14__15 (
              GND0), .q_arr_14__14 (GND0), .q_arr_14__13 (GND0), .q_arr_14__12 (
              GND0), .q_arr_14__11 (GND0), .q_arr_14__10 (GND0), .q_arr_14__9 (
              GND0), .q_arr_14__8 (GND0), .q_arr_14__7 (GND0), .q_arr_14__6 (
              GND0), .q_arr_14__5 (GND0), .q_arr_14__4 (GND0), .q_arr_14__3 (
              GND0), .q_arr_14__2 (GND0), .q_arr_14__1 (GND0), .q_arr_14__0 (
              GND0), .q_arr_15__31 (GND0), .q_arr_15__30 (GND0), .q_arr_15__29 (
              GND0), .q_arr_15__28 (GND0), .q_arr_15__27 (GND0), .q_arr_15__26 (
              GND0), .q_arr_15__25 (GND0), .q_arr_15__24 (GND0), .q_arr_15__23 (
              GND0), .q_arr_15__22 (GND0), .q_arr_15__21 (GND0), .q_arr_15__20 (
              GND0), .q_arr_15__19 (GND0), .q_arr_15__18 (GND0), .q_arr_15__17 (
              GND0), .q_arr_15__16 (GND0), .q_arr_15__15 (GND0), .q_arr_15__14 (
              GND0), .q_arr_15__13 (GND0), .q_arr_15__12 (GND0), .q_arr_15__11 (
              GND0), .q_arr_15__10 (GND0), .q_arr_15__9 (GND0), .q_arr_15__8 (
              GND0), .q_arr_15__7 (GND0), .q_arr_15__6 (GND0), .q_arr_15__5 (
              GND0), .q_arr_15__4 (GND0), .q_arr_15__3 (GND0), .q_arr_15__2 (
              GND0), .q_arr_15__1 (GND0), .q_arr_15__0 (GND0), .q_arr_16__31 (
              GND0), .q_arr_16__30 (GND0), .q_arr_16__29 (GND0), .q_arr_16__28 (
              GND0), .q_arr_16__27 (GND0), .q_arr_16__26 (GND0), .q_arr_16__25 (
              GND0), .q_arr_16__24 (GND0), .q_arr_16__23 (GND0), .q_arr_16__22 (
              GND0), .q_arr_16__21 (GND0), .q_arr_16__20 (GND0), .q_arr_16__19 (
              GND0), .q_arr_16__18 (GND0), .q_arr_16__17 (GND0), .q_arr_16__16 (
              GND0), .q_arr_16__15 (GND0), .q_arr_16__14 (GND0), .q_arr_16__13 (
              GND0), .q_arr_16__12 (GND0), .q_arr_16__11 (GND0), .q_arr_16__10 (
              GND0), .q_arr_16__9 (GND0), .q_arr_16__8 (GND0), .q_arr_16__7 (
              GND0), .q_arr_16__6 (GND0), .q_arr_16__5 (GND0), .q_arr_16__4 (
              GND0), .q_arr_16__3 (GND0), .q_arr_16__2 (GND0), .q_arr_16__1 (
              GND0), .q_arr_16__0 (GND0), .q_arr_17__31 (GND0), .q_arr_17__30 (
              GND0), .q_arr_17__29 (GND0), .q_arr_17__28 (GND0), .q_arr_17__27 (
              GND0), .q_arr_17__26 (GND0), .q_arr_17__25 (GND0), .q_arr_17__24 (
              GND0), .q_arr_17__23 (GND0), .q_arr_17__22 (GND0), .q_arr_17__21 (
              GND0), .q_arr_17__20 (GND0), .q_arr_17__19 (GND0), .q_arr_17__18 (
              GND0), .q_arr_17__17 (GND0), .q_arr_17__16 (GND0), .q_arr_17__15 (
              GND0), .q_arr_17__14 (GND0), .q_arr_17__13 (GND0), .q_arr_17__12 (
              GND0), .q_arr_17__11 (GND0), .q_arr_17__10 (GND0), .q_arr_17__9 (
              GND0), .q_arr_17__8 (GND0), .q_arr_17__7 (GND0), .q_arr_17__6 (
              GND0), .q_arr_17__5 (GND0), .q_arr_17__4 (GND0), .q_arr_17__3 (
              GND0), .q_arr_17__2 (GND0), .q_arr_17__1 (GND0), .q_arr_17__0 (
              GND0), .q_arr_18__31 (GND0), .q_arr_18__30 (GND0), .q_arr_18__29 (
              GND0), .q_arr_18__28 (GND0), .q_arr_18__27 (GND0), .q_arr_18__26 (
              GND0), .q_arr_18__25 (GND0), .q_arr_18__24 (GND0), .q_arr_18__23 (
              GND0), .q_arr_18__22 (GND0), .q_arr_18__21 (GND0), .q_arr_18__20 (
              GND0), .q_arr_18__19 (GND0), .q_arr_18__18 (GND0), .q_arr_18__17 (
              GND0), .q_arr_18__16 (GND0), .q_arr_18__15 (GND0), .q_arr_18__14 (
              GND0), .q_arr_18__13 (GND0), .q_arr_18__12 (GND0), .q_arr_18__11 (
              GND0), .q_arr_18__10 (GND0), .q_arr_18__9 (GND0), .q_arr_18__8 (
              GND0), .q_arr_18__7 (GND0), .q_arr_18__6 (GND0), .q_arr_18__5 (
              GND0), .q_arr_18__4 (GND0), .q_arr_18__3 (GND0), .q_arr_18__2 (
              GND0), .q_arr_18__1 (GND0), .q_arr_18__0 (GND0), .q_arr_19__31 (
              GND0), .q_arr_19__30 (GND0), .q_arr_19__29 (GND0), .q_arr_19__28 (
              GND0), .q_arr_19__27 (GND0), .q_arr_19__26 (GND0), .q_arr_19__25 (
              GND0), .q_arr_19__24 (GND0), .q_arr_19__23 (GND0), .q_arr_19__22 (
              GND0), .q_arr_19__21 (GND0), .q_arr_19__20 (GND0), .q_arr_19__19 (
              GND0), .q_arr_19__18 (GND0), .q_arr_19__17 (GND0), .q_arr_19__16 (
              GND0), .q_arr_19__15 (GND0), .q_arr_19__14 (GND0), .q_arr_19__13 (
              GND0), .q_arr_19__12 (GND0), .q_arr_19__11 (GND0), .q_arr_19__10 (
              GND0), .q_arr_19__9 (GND0), .q_arr_19__8 (GND0), .q_arr_19__7 (
              GND0), .q_arr_19__6 (GND0), .q_arr_19__5 (GND0), .q_arr_19__4 (
              GND0), .q_arr_19__3 (GND0), .q_arr_19__2 (GND0), .q_arr_19__1 (
              GND0), .q_arr_19__0 (GND0), .q_arr_20__31 (GND0), .q_arr_20__30 (
              GND0), .q_arr_20__29 (GND0), .q_arr_20__28 (GND0), .q_arr_20__27 (
              GND0), .q_arr_20__26 (GND0), .q_arr_20__25 (GND0), .q_arr_20__24 (
              GND0), .q_arr_20__23 (GND0), .q_arr_20__22 (GND0), .q_arr_20__21 (
              GND0), .q_arr_20__20 (GND0), .q_arr_20__19 (GND0), .q_arr_20__18 (
              GND0), .q_arr_20__17 (GND0), .q_arr_20__16 (GND0), .q_arr_20__15 (
              GND0), .q_arr_20__14 (GND0), .q_arr_20__13 (GND0), .q_arr_20__12 (
              GND0), .q_arr_20__11 (GND0), .q_arr_20__10 (GND0), .q_arr_20__9 (
              GND0), .q_arr_20__8 (GND0), .q_arr_20__7 (GND0), .q_arr_20__6 (
              GND0), .q_arr_20__5 (GND0), .q_arr_20__4 (GND0), .q_arr_20__3 (
              GND0), .q_arr_20__2 (GND0), .q_arr_20__1 (GND0), .q_arr_20__0 (
              GND0), .q_arr_21__31 (GND0), .q_arr_21__30 (GND0), .q_arr_21__29 (
              GND0), .q_arr_21__28 (GND0), .q_arr_21__27 (GND0), .q_arr_21__26 (
              GND0), .q_arr_21__25 (GND0), .q_arr_21__24 (GND0), .q_arr_21__23 (
              GND0), .q_arr_21__22 (GND0), .q_arr_21__21 (GND0), .q_arr_21__20 (
              GND0), .q_arr_21__19 (GND0), .q_arr_21__18 (GND0), .q_arr_21__17 (
              GND0), .q_arr_21__16 (GND0), .q_arr_21__15 (GND0), .q_arr_21__14 (
              GND0), .q_arr_21__13 (GND0), .q_arr_21__12 (GND0), .q_arr_21__11 (
              GND0), .q_arr_21__10 (GND0), .q_arr_21__9 (GND0), .q_arr_21__8 (
              GND0), .q_arr_21__7 (GND0), .q_arr_21__6 (GND0), .q_arr_21__5 (
              GND0), .q_arr_21__4 (GND0), .q_arr_21__3 (GND0), .q_arr_21__2 (
              GND0), .q_arr_21__1 (GND0), .q_arr_21__0 (GND0), .q_arr_22__31 (
              GND0), .q_arr_22__30 (GND0), .q_arr_22__29 (GND0), .q_arr_22__28 (
              GND0), .q_arr_22__27 (GND0), .q_arr_22__26 (GND0), .q_arr_22__25 (
              GND0), .q_arr_22__24 (GND0), .q_arr_22__23 (GND0), .q_arr_22__22 (
              GND0), .q_arr_22__21 (GND0), .q_arr_22__20 (GND0), .q_arr_22__19 (
              GND0), .q_arr_22__18 (GND0), .q_arr_22__17 (GND0), .q_arr_22__16 (
              GND0), .q_arr_22__15 (GND0), .q_arr_22__14 (GND0), .q_arr_22__13 (
              GND0), .q_arr_22__12 (GND0), .q_arr_22__11 (GND0), .q_arr_22__10 (
              GND0), .q_arr_22__9 (GND0), .q_arr_22__8 (GND0), .q_arr_22__7 (
              GND0), .q_arr_22__6 (GND0), .q_arr_22__5 (GND0), .q_arr_22__4 (
              GND0), .q_arr_22__3 (GND0), .q_arr_22__2 (GND0), .q_arr_22__1 (
              GND0), .q_arr_22__0 (GND0), .q_arr_23__31 (GND0), .q_arr_23__30 (
              GND0), .q_arr_23__29 (GND0), .q_arr_23__28 (GND0), .q_arr_23__27 (
              GND0), .q_arr_23__26 (GND0), .q_arr_23__25 (GND0), .q_arr_23__24 (
              GND0), .q_arr_23__23 (GND0), .q_arr_23__22 (GND0), .q_arr_23__21 (
              GND0), .q_arr_23__20 (GND0), .q_arr_23__19 (GND0), .q_arr_23__18 (
              GND0), .q_arr_23__17 (GND0), .q_arr_23__16 (GND0), .q_arr_23__15 (
              GND0), .q_arr_23__14 (GND0), .q_arr_23__13 (GND0), .q_arr_23__12 (
              GND0), .q_arr_23__11 (GND0), .q_arr_23__10 (GND0), .q_arr_23__9 (
              GND0), .q_arr_23__8 (GND0), .q_arr_23__7 (GND0), .q_arr_23__6 (
              GND0), .q_arr_23__5 (GND0), .q_arr_23__4 (GND0), .q_arr_23__3 (
              GND0), .q_arr_23__2 (GND0), .q_arr_23__1 (GND0), .q_arr_23__0 (
              GND0), .q_arr_24__31 (GND0), .q_arr_24__30 (GND0), .q_arr_24__29 (
              GND0), .q_arr_24__28 (GND0), .q_arr_24__27 (GND0), .q_arr_24__26 (
              GND0), .q_arr_24__25 (GND0), .q_arr_24__24 (GND0), .q_arr_24__23 (
              GND0), .q_arr_24__22 (GND0), .q_arr_24__21 (GND0), .q_arr_24__20 (
              GND0), .q_arr_24__19 (GND0), .q_arr_24__18 (GND0), .q_arr_24__17 (
              GND0), .q_arr_24__16 (GND0), .q_arr_24__15 (GND0), .q_arr_24__14 (
              GND0), .q_arr_24__13 (GND0), .q_arr_24__12 (GND0), .q_arr_24__11 (
              GND0), .q_arr_24__10 (GND0), .q_arr_24__9 (GND0), .q_arr_24__8 (
              GND0), .q_arr_24__7 (GND0), .q_arr_24__6 (GND0), .q_arr_24__5 (
              GND0), .q_arr_24__4 (GND0), .q_arr_24__3 (GND0), .q_arr_24__2 (
              GND0), .q_arr_24__1 (GND0), .q_arr_24__0 (GND0)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_0_mul_gen_mul_gen (.M (
                            {img_data_0__15,nx19396,img_data_0__13,
                            img_data_0__12,img_data_0__11,img_data_0__10,
                            img_data_0__9,img_data_0__8,img_data_0__7,
                            img_data_0__6,img_data_0__5,img_data_0__4,
                            img_data_0__3,img_data_0__2,img_data_0__1,
                            img_data_0__0}), .R ({filter_data_0__15,
                            filter_data_0__14,filter_data_0__13,
                            filter_data_0__12,filter_data_0__11,
                            filter_data_0__10,filter_data_0__9,filter_data_0__8,
                            filter_data_0__7,filter_data_0__6,filter_data_0__5,
                            filter_data_0__4,filter_data_0__3,filter_data_0__2,
                            filter_data_0__1,filter_data_0__0}), .cnt_enable (
                            nx16627), .product ({d_arr_mul_0__31,d_arr_mul_0__30
                            ,d_arr_mul_0__29,d_arr_mul_0__28,d_arr_mul_0__27,
                            d_arr_mul_0__26,d_arr_mul_0__25,d_arr_mul_0__24,
                            d_arr_mul_0__23,d_arr_mul_0__22,d_arr_mul_0__21,
                            d_arr_mul_0__20,d_arr_mul_0__19,d_arr_mul_0__18,
                            d_arr_mul_0__17,d_arr_mul_0__16,d_arr_mul_0__15,
                            d_arr_mul_0__14,d_arr_mul_0__13,d_arr_mul_0__12,
                            d_arr_mul_0__11,d_arr_mul_0__10,d_arr_mul_0__9,
                            d_arr_mul_0__8,d_arr_mul_0__7,d_arr_mul_0__6,
                            d_arr_mul_0__5,d_arr_mul_0__4,d_arr_mul_0__3,
                            d_arr_mul_0__2,d_arr_mul_0__1,d_arr_mul_0__0}), .clk (
                            clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_1_mul_gen_mul_gen (.M (
                            {img_data_1__15,nx19400,img_data_1__13,
                            img_data_1__12,img_data_1__11,nx19402,img_data_1__9,
                            img_data_1__8,img_data_1__7,img_data_1__6,
                            img_data_1__5,img_data_1__4,img_data_1__3,
                            img_data_1__2,img_data_1__1,img_data_1__0}), .R ({
                            filter_data_1__15,filter_data_1__14,
                            filter_data_1__13,filter_data_1__12,
                            filter_data_1__11,filter_data_1__10,filter_data_1__9
                            ,filter_data_1__8,filter_data_1__7,filter_data_1__6,
                            filter_data_1__5,filter_data_1__4,filter_data_1__3,
                            filter_data_1__2,filter_data_1__1,filter_data_1__0})
                            , .cnt_enable (nx16473), .product ({d_arr_mul_1__31,
                            d_arr_mul_1__30,d_arr_mul_1__29,d_arr_mul_1__28,
                            d_arr_mul_1__27,d_arr_mul_1__26,d_arr_mul_1__25,
                            d_arr_mul_1__24,d_arr_mul_1__23,d_arr_mul_1__22,
                            d_arr_mul_1__21,d_arr_mul_1__20,d_arr_mul_1__19,
                            d_arr_mul_1__18,d_arr_mul_1__17,d_arr_mul_1__16,
                            d_arr_mul_1__15,d_arr_mul_1__14,d_arr_mul_1__13,
                            d_arr_mul_1__12,d_arr_mul_1__11,d_arr_mul_1__10,
                            d_arr_mul_1__9,d_arr_mul_1__8,d_arr_mul_1__7,
                            d_arr_mul_1__6,d_arr_mul_1__5,d_arr_mul_1__4,
                            d_arr_mul_1__3,d_arr_mul_1__2,d_arr_mul_1__1,
                            d_arr_mul_1__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_2_mul_gen_mul_gen (.M (
                            {img_data_2__15,nx19406,img_data_2__13,
                            img_data_2__12,img_data_2__11,nx19408,img_data_2__9,
                            img_data_2__8,img_data_2__7,img_data_2__6,
                            img_data_2__5,img_data_2__4,img_data_2__3,
                            img_data_2__2,img_data_2__1,img_data_2__0}), .R ({
                            filter_data_2__15,filter_data_2__14,
                            filter_data_2__13,filter_data_2__12,
                            filter_data_2__11,filter_data_2__10,filter_data_2__9
                            ,filter_data_2__8,filter_data_2__7,filter_data_2__6,
                            filter_data_2__5,filter_data_2__4,filter_data_2__3,
                            filter_data_2__2,filter_data_2__1,filter_data_2__0})
                            , .cnt_enable (nx16473), .product ({d_arr_mul_2__31,
                            d_arr_mul_2__30,d_arr_mul_2__29,d_arr_mul_2__28,
                            d_arr_mul_2__27,d_arr_mul_2__26,d_arr_mul_2__25,
                            d_arr_mul_2__24,d_arr_mul_2__23,d_arr_mul_2__22,
                            d_arr_mul_2__21,d_arr_mul_2__20,d_arr_mul_2__19,
                            d_arr_mul_2__18,d_arr_mul_2__17,d_arr_mul_2__16,
                            d_arr_mul_2__15,d_arr_mul_2__14,d_arr_mul_2__13,
                            d_arr_mul_2__12,d_arr_mul_2__11,d_arr_mul_2__10,
                            d_arr_mul_2__9,d_arr_mul_2__8,d_arr_mul_2__7,
                            d_arr_mul_2__6,d_arr_mul_2__5,d_arr_mul_2__4,
                            d_arr_mul_2__3,d_arr_mul_2__2,d_arr_mul_2__1,
                            d_arr_mul_2__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_3_mul_gen_mul_gen (.M (
                            {img_data_5__15,nx19410,img_data_5__13,
                            img_data_5__12,img_data_5__11,img_data_5__10,
                            img_data_5__9,img_data_5__8,img_data_5__7,
                            img_data_5__6,img_data_5__5,img_data_5__4,
                            img_data_5__3,img_data_5__2,img_data_5__1,
                            img_data_5__0}), .R ({ordered_filter_data_3__15,
                            ordered_filter_data_3__14,ordered_filter_data_3__13,
                            ordered_filter_data_3__12,ordered_filter_data_3__11,
                            ordered_filter_data_3__10,ordered_filter_data_3__9,
                            ordered_filter_data_3__8,ordered_filter_data_3__7,
                            ordered_filter_data_3__6,ordered_filter_data_3__5,
                            ordered_filter_data_3__4,ordered_filter_data_3__3,
                            ordered_filter_data_3__2,ordered_filter_data_3__1,
                            ordered_filter_data_3__0}), .cnt_enable (nx16629), .product (
                            {d_arr_mul_3__31,d_arr_mul_3__30,d_arr_mul_3__29,
                            d_arr_mul_3__28,d_arr_mul_3__27,d_arr_mul_3__26,
                            d_arr_mul_3__25,d_arr_mul_3__24,d_arr_mul_3__23,
                            d_arr_mul_3__22,d_arr_mul_3__21,d_arr_mul_3__20,
                            d_arr_mul_3__19,d_arr_mul_3__18,d_arr_mul_3__17,
                            d_arr_mul_3__16,d_arr_mul_3__15,d_arr_mul_3__14,
                            d_arr_mul_3__13,d_arr_mul_3__12,d_arr_mul_3__11,
                            d_arr_mul_3__10,d_arr_mul_3__9,d_arr_mul_3__8,
                            d_arr_mul_3__7,d_arr_mul_3__6,d_arr_mul_3__5,
                            d_arr_mul_3__4,d_arr_mul_3__3,d_arr_mul_3__2,
                            d_arr_mul_3__1,d_arr_mul_3__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_4_mul_gen_mul_gen (.M (
                            {img_data_6__15,nx19414,img_data_6__13,
                            img_data_6__12,img_data_6__11,nx19416,img_data_6__9,
                            img_data_6__8,img_data_6__7,img_data_6__6,
                            img_data_6__5,img_data_6__4,img_data_6__3,
                            img_data_6__2,img_data_6__1,img_data_6__0}), .R ({
                            ordered_filter_data_4__15,ordered_filter_data_4__14,
                            ordered_filter_data_4__13,ordered_filter_data_4__12,
                            ordered_filter_data_4__11,ordered_filter_data_4__10,
                            ordered_filter_data_4__9,ordered_filter_data_4__8,
                            ordered_filter_data_4__7,ordered_filter_data_4__6,
                            ordered_filter_data_4__5,ordered_filter_data_4__4,
                            ordered_filter_data_4__3,ordered_filter_data_4__2,
                            ordered_filter_data_4__1,ordered_filter_data_4__0})
                            , .cnt_enable (nx16629), .product ({d_arr_mul_4__31,
                            d_arr_mul_4__30,d_arr_mul_4__29,d_arr_mul_4__28,
                            d_arr_mul_4__27,d_arr_mul_4__26,d_arr_mul_4__25,
                            d_arr_mul_4__24,d_arr_mul_4__23,d_arr_mul_4__22,
                            d_arr_mul_4__21,d_arr_mul_4__20,d_arr_mul_4__19,
                            d_arr_mul_4__18,d_arr_mul_4__17,d_arr_mul_4__16,
                            d_arr_mul_4__15,d_arr_mul_4__14,d_arr_mul_4__13,
                            d_arr_mul_4__12,d_arr_mul_4__11,d_arr_mul_4__10,
                            d_arr_mul_4__9,d_arr_mul_4__8,d_arr_mul_4__7,
                            d_arr_mul_4__6,d_arr_mul_4__5,d_arr_mul_4__4,
                            d_arr_mul_4__3,d_arr_mul_4__2,d_arr_mul_4__1,
                            d_arr_mul_4__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_5_mul_gen_mul_gen (.M (
                            {nx16659,nx19420,img_data_7__13,img_data_7__12,
                            img_data_7__11,nx19422,img_data_7__9,img_data_7__8,
                            img_data_7__7,img_data_7__6,img_data_7__5,
                            img_data_7__4,img_data_7__3,img_data_7__2,
                            img_data_7__1,img_data_7__0}), .R ({
                            ordered_filter_data_5__15,ordered_filter_data_5__14,
                            ordered_filter_data_5__13,ordered_filter_data_5__12,
                            ordered_filter_data_5__11,ordered_filter_data_5__10,
                            ordered_filter_data_5__9,ordered_filter_data_5__8,
                            ordered_filter_data_5__7,ordered_filter_data_5__6,
                            ordered_filter_data_5__5,ordered_filter_data_5__4,
                            ordered_filter_data_5__3,ordered_filter_data_5__2,
                            ordered_filter_data_5__1,ordered_filter_data_5__0})
                            , .cnt_enable (nx16631), .product ({d_arr_mul_5__31,
                            d_arr_mul_5__30,d_arr_mul_5__29,d_arr_mul_5__28,
                            d_arr_mul_5__27,d_arr_mul_5__26,d_arr_mul_5__25,
                            d_arr_mul_5__24,d_arr_mul_5__23,d_arr_mul_5__22,
                            d_arr_mul_5__21,d_arr_mul_5__20,d_arr_mul_5__19,
                            d_arr_mul_5__18,d_arr_mul_5__17,d_arr_mul_5__16,
                            d_arr_mul_5__15,d_arr_mul_5__14,d_arr_mul_5__13,
                            d_arr_mul_5__12,d_arr_mul_5__11,d_arr_mul_5__10,
                            d_arr_mul_5__9,d_arr_mul_5__8,d_arr_mul_5__7,
                            d_arr_mul_5__6,d_arr_mul_5__5,d_arr_mul_5__4,
                            d_arr_mul_5__3,d_arr_mul_5__2,d_arr_mul_5__1,
                            d_arr_mul_5__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_6_mul_gen_mul_gen (.M (
                            {img_data_10__15,nx19424,img_data_10__13,
                            img_data_10__12,img_data_10__11,img_data_10__10,
                            img_data_10__9,img_data_10__8,img_data_10__7,
                            img_data_10__6,img_data_10__5,img_data_10__4,
                            img_data_10__3,img_data_10__2,img_data_10__1,
                            img_data_10__0}), .R ({ordered_filter_data_6__15,
                            ordered_filter_data_6__14,ordered_filter_data_6__13,
                            ordered_filter_data_6__12,ordered_filter_data_6__11,
                            ordered_filter_data_6__10,ordered_filter_data_6__9,
                            ordered_filter_data_6__8,ordered_filter_data_6__7,
                            ordered_filter_data_6__6,ordered_filter_data_6__5,
                            ordered_filter_data_6__4,ordered_filter_data_6__3,
                            ordered_filter_data_6__2,ordered_filter_data_6__1,
                            ordered_filter_data_6__0}), .cnt_enable (nx16631), .product (
                            {d_arr_mul_6__31,d_arr_mul_6__30,d_arr_mul_6__29,
                            d_arr_mul_6__28,d_arr_mul_6__27,d_arr_mul_6__26,
                            d_arr_mul_6__25,d_arr_mul_6__24,d_arr_mul_6__23,
                            d_arr_mul_6__22,d_arr_mul_6__21,d_arr_mul_6__20,
                            d_arr_mul_6__19,d_arr_mul_6__18,d_arr_mul_6__17,
                            d_arr_mul_6__16,d_arr_mul_6__15,d_arr_mul_6__14,
                            d_arr_mul_6__13,d_arr_mul_6__12,d_arr_mul_6__11,
                            d_arr_mul_6__10,d_arr_mul_6__9,d_arr_mul_6__8,
                            d_arr_mul_6__7,d_arr_mul_6__6,d_arr_mul_6__5,
                            d_arr_mul_6__4,d_arr_mul_6__3,d_arr_mul_6__2,
                            d_arr_mul_6__1,d_arr_mul_6__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_7_mul_gen_mul_gen (.M (
                            {nx16661,nx19428,img_data_11__13,img_data_11__12,
                            img_data_11__11,nx19430,img_data_11__9,
                            img_data_11__8,img_data_11__7,img_data_11__6,
                            img_data_11__5,img_data_11__4,img_data_11__3,
                            img_data_11__2,img_data_11__1,img_data_11__0}), .R (
                            {ordered_filter_data_7__15,ordered_filter_data_7__14
                            ,ordered_filter_data_7__13,ordered_filter_data_7__12
                            ,ordered_filter_data_7__11,ordered_filter_data_7__10
                            ,ordered_filter_data_7__9,ordered_filter_data_7__8,
                            ordered_filter_data_7__7,ordered_filter_data_7__6,
                            ordered_filter_data_7__5,ordered_filter_data_7__4,
                            ordered_filter_data_7__3,ordered_filter_data_7__2,
                            ordered_filter_data_7__1,ordered_filter_data_7__0})
                            , .cnt_enable (nx16633), .product ({d_arr_mul_7__31,
                            d_arr_mul_7__30,d_arr_mul_7__29,d_arr_mul_7__28,
                            d_arr_mul_7__27,d_arr_mul_7__26,d_arr_mul_7__25,
                            d_arr_mul_7__24,d_arr_mul_7__23,d_arr_mul_7__22,
                            d_arr_mul_7__21,d_arr_mul_7__20,d_arr_mul_7__19,
                            d_arr_mul_7__18,d_arr_mul_7__17,d_arr_mul_7__16,
                            d_arr_mul_7__15,d_arr_mul_7__14,d_arr_mul_7__13,
                            d_arr_mul_7__12,d_arr_mul_7__11,d_arr_mul_7__10,
                            d_arr_mul_7__9,d_arr_mul_7__8,d_arr_mul_7__7,
                            d_arr_mul_7__6,d_arr_mul_7__5,d_arr_mul_7__4,
                            d_arr_mul_7__3,d_arr_mul_7__2,d_arr_mul_7__1,
                            d_arr_mul_7__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_8_mul_gen_mul_gen (.M (
                            {nx16663,nx19434,img_data_12__13,img_data_12__12,
                            img_data_12__11,nx19436,img_data_12__9,
                            img_data_12__8,img_data_12__7,img_data_12__6,
                            img_data_12__5,img_data_12__4,img_data_12__3,
                            img_data_12__2,img_data_12__1,img_data_12__0}), .R (
                            {ordered_filter_data_8__15,ordered_filter_data_8__14
                            ,ordered_filter_data_8__13,ordered_filter_data_8__12
                            ,ordered_filter_data_8__11,ordered_filter_data_8__10
                            ,ordered_filter_data_8__9,ordered_filter_data_8__8,
                            ordered_filter_data_8__7,ordered_filter_data_8__6,
                            ordered_filter_data_8__5,ordered_filter_data_8__4,
                            ordered_filter_data_8__3,ordered_filter_data_8__2,
                            ordered_filter_data_8__1,ordered_filter_data_8__0})
                            , .cnt_enable (nx16633), .product ({d_arr_mul_8__31,
                            d_arr_mul_8__30,d_arr_mul_8__29,d_arr_mul_8__28,
                            d_arr_mul_8__27,d_arr_mul_8__26,d_arr_mul_8__25,
                            d_arr_mul_8__24,d_arr_mul_8__23,d_arr_mul_8__22,
                            d_arr_mul_8__21,d_arr_mul_8__20,d_arr_mul_8__19,
                            d_arr_mul_8__18,d_arr_mul_8__17,d_arr_mul_8__16,
                            d_arr_mul_8__15,d_arr_mul_8__14,d_arr_mul_8__13,
                            d_arr_mul_8__12,d_arr_mul_8__11,d_arr_mul_8__10,
                            d_arr_mul_8__9,d_arr_mul_8__8,d_arr_mul_8__7,
                            d_arr_mul_8__6,d_arr_mul_8__5,d_arr_mul_8__4,
                            d_arr_mul_8__3,d_arr_mul_8__2,d_arr_mul_8__1,
                            d_arr_mul_8__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_9_mul_gen_mul_gen (.M (
                            {nx16405,ordered_img_data_9__14,
                            ordered_img_data_9__13,ordered_img_data_9__12,
                            ordered_img_data_9__11,ordered_img_data_9__10,
                            ordered_img_data_9__9,ordered_img_data_9__8,
                            ordered_img_data_9__7,ordered_img_data_9__6,
                            ordered_img_data_9__5,ordered_img_data_9__4,
                            ordered_img_data_9__3,ordered_img_data_9__2,
                            ordered_img_data_9__1,ordered_img_data_9__0}), .R ({
                            ordered_filter_data_9__15,ordered_filter_data_9__14,
                            ordered_filter_data_9__13,ordered_filter_data_9__12,
                            ordered_filter_data_9__11,ordered_filter_data_9__10,
                            ordered_filter_data_9__9,ordered_filter_data_9__8,
                            ordered_filter_data_9__7,ordered_filter_data_9__6,
                            ordered_filter_data_9__5,ordered_filter_data_9__4,
                            ordered_filter_data_9__3,ordered_filter_data_9__2,
                            ordered_filter_data_9__1,ordered_filter_data_9__0})
                            , .cnt_enable (nx16475), .product ({d_arr_mul_9__31,
                            d_arr_mul_9__30,d_arr_mul_9__29,d_arr_mul_9__28,
                            d_arr_mul_9__27,d_arr_mul_9__26,d_arr_mul_9__25,
                            d_arr_mul_9__24,d_arr_mul_9__23,d_arr_mul_9__22,
                            d_arr_mul_9__21,d_arr_mul_9__20,d_arr_mul_9__19,
                            d_arr_mul_9__18,d_arr_mul_9__17,d_arr_mul_9__16,
                            d_arr_mul_9__15,d_arr_mul_9__14,d_arr_mul_9__13,
                            d_arr_mul_9__12,d_arr_mul_9__11,d_arr_mul_9__10,
                            d_arr_mul_9__9,d_arr_mul_9__8,d_arr_mul_9__7,
                            d_arr_mul_9__6,d_arr_mul_9__5,d_arr_mul_9__4,
                            d_arr_mul_9__3,d_arr_mul_9__2,d_arr_mul_9__1,
                            d_arr_mul_9__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_10_mul_gen_mul_gen (.M (
                            {nx16413,ordered_img_data_10__14,
                            ordered_img_data_10__13,ordered_img_data_10__12,
                            ordered_img_data_10__11,ordered_img_data_10__10,
                            ordered_img_data_10__9,ordered_img_data_10__8,
                            ordered_img_data_10__7,ordered_img_data_10__6,
                            ordered_img_data_10__5,ordered_img_data_10__4,
                            ordered_img_data_10__3,ordered_img_data_10__2,
                            ordered_img_data_10__1,ordered_img_data_10__0}), .R (
                            {ordered_filter_data_10__15,
                            ordered_filter_data_10__14,
                            ordered_filter_data_10__13,
                            ordered_filter_data_10__12,
                            ordered_filter_data_10__11,
                            ordered_filter_data_10__10,ordered_filter_data_10__9
                            ,ordered_filter_data_10__8,ordered_filter_data_10__7
                            ,ordered_filter_data_10__6,ordered_filter_data_10__5
                            ,ordered_filter_data_10__4,ordered_filter_data_10__3
                            ,ordered_filter_data_10__2,ordered_filter_data_10__1
                            ,ordered_filter_data_10__0}), .cnt_enable (nx16635)
                            , .product ({d_arr_mul_10__31,d_arr_mul_10__30,
                            d_arr_mul_10__29,d_arr_mul_10__28,d_arr_mul_10__27,
                            d_arr_mul_10__26,d_arr_mul_10__25,d_arr_mul_10__24,
                            d_arr_mul_10__23,d_arr_mul_10__22,d_arr_mul_10__21,
                            d_arr_mul_10__20,d_arr_mul_10__19,d_arr_mul_10__18,
                            d_arr_mul_10__17,d_arr_mul_10__16,d_arr_mul_10__15,
                            d_arr_mul_10__14,d_arr_mul_10__13,d_arr_mul_10__12,
                            d_arr_mul_10__11,d_arr_mul_10__10,d_arr_mul_10__9,
                            d_arr_mul_10__8,d_arr_mul_10__7,d_arr_mul_10__6,
                            d_arr_mul_10__5,d_arr_mul_10__4,d_arr_mul_10__3,
                            d_arr_mul_10__2,d_arr_mul_10__1,d_arr_mul_10__0}), .clk (
                            clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_11_mul_gen_mul_gen (.M (
                            {nx16421,ordered_img_data_11__14,
                            ordered_img_data_11__13,ordered_img_data_11__12,
                            ordered_img_data_11__11,ordered_img_data_11__10,
                            ordered_img_data_11__9,ordered_img_data_11__8,
                            ordered_img_data_11__7,ordered_img_data_11__6,
                            ordered_img_data_11__5,ordered_img_data_11__4,
                            ordered_img_data_11__3,ordered_img_data_11__2,
                            ordered_img_data_11__1,ordered_img_data_11__0}), .R (
                            {ordered_filter_data_11__15,
                            ordered_filter_data_11__14,
                            ordered_filter_data_11__13,
                            ordered_filter_data_11__12,
                            ordered_filter_data_11__11,
                            ordered_filter_data_11__10,ordered_filter_data_11__9
                            ,ordered_filter_data_11__8,ordered_filter_data_11__7
                            ,ordered_filter_data_11__6,ordered_filter_data_11__5
                            ,ordered_filter_data_11__4,ordered_filter_data_11__3
                            ,ordered_filter_data_11__2,ordered_filter_data_11__1
                            ,ordered_filter_data_11__0}), .cnt_enable (nx16635)
                            , .product ({d_arr_mul_11__31,d_arr_mul_11__30,
                            d_arr_mul_11__29,d_arr_mul_11__28,d_arr_mul_11__27,
                            d_arr_mul_11__26,d_arr_mul_11__25,d_arr_mul_11__24,
                            d_arr_mul_11__23,d_arr_mul_11__22,d_arr_mul_11__21,
                            d_arr_mul_11__20,d_arr_mul_11__19,d_arr_mul_11__18,
                            d_arr_mul_11__17,d_arr_mul_11__16,d_arr_mul_11__15,
                            d_arr_mul_11__14,d_arr_mul_11__13,d_arr_mul_11__12,
                            d_arr_mul_11__11,d_arr_mul_11__10,d_arr_mul_11__9,
                            d_arr_mul_11__8,d_arr_mul_11__7,d_arr_mul_11__6,
                            d_arr_mul_11__5,d_arr_mul_11__4,d_arr_mul_11__3,
                            d_arr_mul_11__2,d_arr_mul_11__1,d_arr_mul_11__0}), .clk (
                            clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_12_mul_gen_mul_gen (.M (
                            {nx16429,ordered_img_data_12__14,
                            ordered_img_data_12__13,ordered_img_data_12__12,
                            ordered_img_data_12__11,ordered_img_data_12__10,
                            ordered_img_data_12__9,ordered_img_data_12__8,
                            ordered_img_data_12__7,ordered_img_data_12__6,
                            ordered_img_data_12__5,ordered_img_data_12__4,
                            ordered_img_data_12__3,ordered_img_data_12__2,
                            ordered_img_data_12__1,ordered_img_data_12__0}), .R (
                            {ordered_filter_data_12__15,
                            ordered_filter_data_12__14,
                            ordered_filter_data_12__13,
                            ordered_filter_data_12__12,
                            ordered_filter_data_12__11,
                            ordered_filter_data_12__10,ordered_filter_data_12__9
                            ,ordered_filter_data_12__8,ordered_filter_data_12__7
                            ,ordered_filter_data_12__6,ordered_filter_data_12__5
                            ,ordered_filter_data_12__4,ordered_filter_data_12__3
                            ,ordered_filter_data_12__2,ordered_filter_data_12__1
                            ,ordered_filter_data_12__0}), .cnt_enable (nx16637)
                            , .product ({d_arr_mul_12__31,d_arr_mul_12__30,
                            d_arr_mul_12__29,d_arr_mul_12__28,d_arr_mul_12__27,
                            d_arr_mul_12__26,d_arr_mul_12__25,d_arr_mul_12__24,
                            d_arr_mul_12__23,d_arr_mul_12__22,d_arr_mul_12__21,
                            d_arr_mul_12__20,d_arr_mul_12__19,d_arr_mul_12__18,
                            d_arr_mul_12__17,d_arr_mul_12__16,d_arr_mul_12__15,
                            d_arr_mul_12__14,d_arr_mul_12__13,d_arr_mul_12__12,
                            d_arr_mul_12__11,d_arr_mul_12__10,d_arr_mul_12__9,
                            d_arr_mul_12__8,d_arr_mul_12__7,d_arr_mul_12__6,
                            d_arr_mul_12__5,d_arr_mul_12__4,d_arr_mul_12__3,
                            d_arr_mul_12__2,d_arr_mul_12__1,d_arr_mul_12__0}), .clk (
                            clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_13_mul_gen_mul_gen (.M (
                            {nx16437,ordered_img_data_13__14,
                            ordered_img_data_13__13,ordered_img_data_13__12,
                            ordered_img_data_13__11,ordered_img_data_13__10,
                            ordered_img_data_13__9,ordered_img_data_13__8,
                            ordered_img_data_13__7,ordered_img_data_13__6,
                            ordered_img_data_13__5,ordered_img_data_13__4,
                            ordered_img_data_13__3,ordered_img_data_13__2,
                            ordered_img_data_13__1,ordered_img_data_13__0}), .R (
                            {ordered_filter_data_13__15,
                            ordered_filter_data_13__14,
                            ordered_filter_data_13__13,
                            ordered_filter_data_13__12,
                            ordered_filter_data_13__11,
                            ordered_filter_data_13__10,ordered_filter_data_13__9
                            ,ordered_filter_data_13__8,ordered_filter_data_13__7
                            ,ordered_filter_data_13__6,ordered_filter_data_13__5
                            ,ordered_filter_data_13__4,ordered_filter_data_13__3
                            ,ordered_filter_data_13__2,ordered_filter_data_13__1
                            ,ordered_filter_data_13__0}), .cnt_enable (nx16637)
                            , .product ({d_arr_mul_13__31,d_arr_mul_13__30,
                            d_arr_mul_13__29,d_arr_mul_13__28,d_arr_mul_13__27,
                            d_arr_mul_13__26,d_arr_mul_13__25,d_arr_mul_13__24,
                            d_arr_mul_13__23,d_arr_mul_13__22,d_arr_mul_13__21,
                            d_arr_mul_13__20,d_arr_mul_13__19,d_arr_mul_13__18,
                            d_arr_mul_13__17,d_arr_mul_13__16,d_arr_mul_13__15,
                            d_arr_mul_13__14,d_arr_mul_13__13,d_arr_mul_13__12,
                            d_arr_mul_13__11,d_arr_mul_13__10,d_arr_mul_13__9,
                            d_arr_mul_13__8,d_arr_mul_13__7,d_arr_mul_13__6,
                            d_arr_mul_13__5,d_arr_mul_13__4,d_arr_mul_13__3,
                            d_arr_mul_13__2,d_arr_mul_13__1,d_arr_mul_13__0}), .clk (
                            clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_14_mul_gen_mul_gen (.M (
                            {nx16445,ordered_img_data_14__14,
                            ordered_img_data_14__13,ordered_img_data_14__12,
                            ordered_img_data_14__11,ordered_img_data_14__10,
                            ordered_img_data_14__9,ordered_img_data_14__8,
                            ordered_img_data_14__7,ordered_img_data_14__6,
                            ordered_img_data_14__5,ordered_img_data_14__4,
                            ordered_img_data_14__3,ordered_img_data_14__2,
                            ordered_img_data_14__1,ordered_img_data_14__0}), .R (
                            {ordered_filter_data_14__15,
                            ordered_filter_data_14__14,
                            ordered_filter_data_14__13,
                            ordered_filter_data_14__12,
                            ordered_filter_data_14__11,
                            ordered_filter_data_14__10,ordered_filter_data_14__9
                            ,ordered_filter_data_14__8,ordered_filter_data_14__7
                            ,ordered_filter_data_14__6,ordered_filter_data_14__5
                            ,ordered_filter_data_14__4,ordered_filter_data_14__3
                            ,ordered_filter_data_14__2,ordered_filter_data_14__1
                            ,ordered_filter_data_14__0}), .cnt_enable (nx16639)
                            , .product ({d_arr_mul_14__31,d_arr_mul_14__30,
                            d_arr_mul_14__29,d_arr_mul_14__28,d_arr_mul_14__27,
                            d_arr_mul_14__26,d_arr_mul_14__25,d_arr_mul_14__24,
                            d_arr_mul_14__23,d_arr_mul_14__22,d_arr_mul_14__21,
                            d_arr_mul_14__20,d_arr_mul_14__19,d_arr_mul_14__18,
                            d_arr_mul_14__17,d_arr_mul_14__16,d_arr_mul_14__15,
                            d_arr_mul_14__14,d_arr_mul_14__13,d_arr_mul_14__12,
                            d_arr_mul_14__11,d_arr_mul_14__10,d_arr_mul_14__9,
                            d_arr_mul_14__8,d_arr_mul_14__7,d_arr_mul_14__6,
                            d_arr_mul_14__5,d_arr_mul_14__4,d_arr_mul_14__3,
                            d_arr_mul_14__2,d_arr_mul_14__1,d_arr_mul_14__0}), .clk (
                            clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_15_mul_gen_mul_gen (.M (
                            {nx16453,ordered_img_data_15__14,
                            ordered_img_data_15__13,ordered_img_data_15__12,
                            ordered_img_data_15__11,ordered_img_data_15__10,
                            ordered_img_data_15__9,ordered_img_data_15__8,
                            ordered_img_data_15__7,ordered_img_data_15__6,
                            ordered_img_data_15__5,ordered_img_data_15__4,
                            ordered_img_data_15__3,ordered_img_data_15__2,
                            ordered_img_data_15__1,ordered_img_data_15__0}), .R (
                            {ordered_filter_data_15__15,
                            ordered_filter_data_15__14,
                            ordered_filter_data_15__13,
                            ordered_filter_data_15__12,
                            ordered_filter_data_15__11,
                            ordered_filter_data_15__10,ordered_filter_data_15__9
                            ,ordered_filter_data_15__8,ordered_filter_data_15__7
                            ,ordered_filter_data_15__6,ordered_filter_data_15__5
                            ,ordered_filter_data_15__4,ordered_filter_data_15__3
                            ,ordered_filter_data_15__2,ordered_filter_data_15__1
                            ,ordered_filter_data_15__0}), .cnt_enable (nx16639)
                            , .product ({d_arr_mul_15__31,d_arr_mul_15__30,
                            d_arr_mul_15__29,d_arr_mul_15__28,d_arr_mul_15__27,
                            d_arr_mul_15__26,d_arr_mul_15__25,d_arr_mul_15__24,
                            d_arr_mul_15__23,d_arr_mul_15__22,d_arr_mul_15__21,
                            d_arr_mul_15__20,d_arr_mul_15__19,d_arr_mul_15__18,
                            d_arr_mul_15__17,d_arr_mul_15__16,d_arr_mul_15__15,
                            d_arr_mul_15__14,d_arr_mul_15__13,d_arr_mul_15__12,
                            d_arr_mul_15__11,d_arr_mul_15__10,d_arr_mul_15__9,
                            d_arr_mul_15__8,d_arr_mul_15__7,d_arr_mul_15__6,
                            d_arr_mul_15__5,d_arr_mul_15__4,d_arr_mul_15__3,
                            d_arr_mul_15__2,d_arr_mul_15__1,d_arr_mul_15__0}), .clk (
                            clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_16_mul_gen_mul_gen (.M (
                            {nx16461,ordered_img_data_16__14,
                            ordered_img_data_16__13,ordered_img_data_16__12,
                            ordered_img_data_16__11,ordered_img_data_16__10,
                            ordered_img_data_16__9,ordered_img_data_16__8,
                            ordered_img_data_16__7,ordered_img_data_16__6,
                            ordered_img_data_16__5,ordered_img_data_16__4,
                            ordered_img_data_16__3,ordered_img_data_16__2,
                            ordered_img_data_16__1,ordered_img_data_16__0}), .R (
                            {ordered_filter_data_16__15,
                            ordered_filter_data_16__14,
                            ordered_filter_data_16__13,
                            ordered_filter_data_16__12,
                            ordered_filter_data_16__11,
                            ordered_filter_data_16__10,ordered_filter_data_16__9
                            ,ordered_filter_data_16__8,ordered_filter_data_16__7
                            ,ordered_filter_data_16__6,ordered_filter_data_16__5
                            ,ordered_filter_data_16__4,ordered_filter_data_16__3
                            ,ordered_filter_data_16__2,ordered_filter_data_16__1
                            ,ordered_filter_data_16__0}), .cnt_enable (nx16477)
                            , .product ({d_arr_mul_16__31,d_arr_mul_16__30,
                            d_arr_mul_16__29,d_arr_mul_16__28,d_arr_mul_16__27,
                            d_arr_mul_16__26,d_arr_mul_16__25,d_arr_mul_16__24,
                            d_arr_mul_16__23,d_arr_mul_16__22,d_arr_mul_16__21,
                            d_arr_mul_16__20,d_arr_mul_16__19,d_arr_mul_16__18,
                            d_arr_mul_16__17,d_arr_mul_16__16,d_arr_mul_16__15,
                            d_arr_mul_16__14,d_arr_mul_16__13,d_arr_mul_16__12,
                            d_arr_mul_16__11,d_arr_mul_16__10,d_arr_mul_16__9,
                            d_arr_mul_16__8,d_arr_mul_16__7,d_arr_mul_16__6,
                            d_arr_mul_16__5,d_arr_mul_16__4,d_arr_mul_16__3,
                            d_arr_mul_16__2,d_arr_mul_16__1,d_arr_mul_16__0}), .clk (
                            clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_17_mul_gen_mul_gen (.M (
                            {nx16469,ordered_img_data_17__14,
                            ordered_img_data_17__13,ordered_img_data_17__12,
                            ordered_img_data_17__11,ordered_img_data_17__10,
                            ordered_img_data_17__9,ordered_img_data_17__8,
                            ordered_img_data_17__7,ordered_img_data_17__6,
                            ordered_img_data_17__5,ordered_img_data_17__4,
                            ordered_img_data_17__3,ordered_img_data_17__2,
                            ordered_img_data_17__1,ordered_img_data_17__0}), .R (
                            {ordered_filter_data_17__15,
                            ordered_filter_data_17__14,
                            ordered_filter_data_17__13,
                            ordered_filter_data_17__12,
                            ordered_filter_data_17__11,
                            ordered_filter_data_17__10,ordered_filter_data_17__9
                            ,ordered_filter_data_17__8,ordered_filter_data_17__7
                            ,ordered_filter_data_17__6,ordered_filter_data_17__5
                            ,ordered_filter_data_17__4,ordered_filter_data_17__3
                            ,ordered_filter_data_17__2,ordered_filter_data_17__1
                            ,ordered_filter_data_17__0}), .cnt_enable (nx16641)
                            , .product ({d_arr_mul_17__31,d_arr_mul_17__30,
                            d_arr_mul_17__29,d_arr_mul_17__28,d_arr_mul_17__27,
                            d_arr_mul_17__26,d_arr_mul_17__25,d_arr_mul_17__24,
                            d_arr_mul_17__23,d_arr_mul_17__22,d_arr_mul_17__21,
                            d_arr_mul_17__20,d_arr_mul_17__19,d_arr_mul_17__18,
                            d_arr_mul_17__17,d_arr_mul_17__16,d_arr_mul_17__15,
                            d_arr_mul_17__14,d_arr_mul_17__13,d_arr_mul_17__12,
                            d_arr_mul_17__11,d_arr_mul_17__10,d_arr_mul_17__9,
                            d_arr_mul_17__8,d_arr_mul_17__7,d_arr_mul_17__6,
                            d_arr_mul_17__5,d_arr_mul_17__4,d_arr_mul_17__3,
                            d_arr_mul_17__2,d_arr_mul_17__1,d_arr_mul_17__0}), .clk (
                            clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_18_mul_gen_mul_gen (.M (
                            {img_data_18__15,nx19438,img_data_18__13,
                            img_data_18__12,img_data_18__11,img_data_18__10,
                            img_data_18__9,img_data_18__8,img_data_18__7,
                            img_data_18__6,img_data_18__5,img_data_18__4,
                            img_data_18__3,img_data_18__2,img_data_18__1,
                            img_data_18__0}), .R ({filter_data_18__15,
                            filter_data_18__14,filter_data_18__13,
                            filter_data_18__12,filter_data_18__11,
                            filter_data_18__10,filter_data_18__9,
                            filter_data_18__8,filter_data_18__7,
                            filter_data_18__6,filter_data_18__5,
                            filter_data_18__4,filter_data_18__3,
                            filter_data_18__2,filter_data_18__1,
                            filter_data_18__0}), .cnt_enable (nx16641), .product (
                            {d_arr_mul_18__31,d_arr_mul_18__30,d_arr_mul_18__29,
                            d_arr_mul_18__28,d_arr_mul_18__27,d_arr_mul_18__26,
                            d_arr_mul_18__25,d_arr_mul_18__24,d_arr_mul_18__23,
                            d_arr_mul_18__22,d_arr_mul_18__21,d_arr_mul_18__20,
                            d_arr_mul_18__19,d_arr_mul_18__18,d_arr_mul_18__17,
                            d_arr_mul_18__16,d_arr_mul_18__15,d_arr_mul_18__14,
                            d_arr_mul_18__13,d_arr_mul_18__12,d_arr_mul_18__11,
                            d_arr_mul_18__10,d_arr_mul_18__9,d_arr_mul_18__8,
                            d_arr_mul_18__7,d_arr_mul_18__6,d_arr_mul_18__5,
                            d_arr_mul_18__4,d_arr_mul_18__3,d_arr_mul_18__2,
                            d_arr_mul_18__1,d_arr_mul_18__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_19_mul_gen_mul_gen (.M (
                            {img_data_19__15,img_data_19__14,img_data_19__13,
                            img_data_19__12,img_data_19__11,img_data_19__10,
                            img_data_19__9,img_data_19__8,img_data_19__7,
                            img_data_19__6,img_data_19__5,img_data_19__4,
                            img_data_19__3,img_data_19__2,img_data_19__1,
                            img_data_19__0}), .R ({filter_data_19__15,
                            filter_data_19__14,filter_data_19__13,
                            filter_data_19__12,filter_data_19__11,
                            filter_data_19__10,filter_data_19__9,
                            filter_data_19__8,filter_data_19__7,
                            filter_data_19__6,filter_data_19__5,
                            filter_data_19__4,filter_data_19__3,
                            filter_data_19__2,filter_data_19__1,
                            filter_data_19__0}), .cnt_enable (nx16643), .product (
                            {d_arr_mul_19__31,d_arr_mul_19__30,d_arr_mul_19__29,
                            d_arr_mul_19__28,d_arr_mul_19__27,d_arr_mul_19__26,
                            d_arr_mul_19__25,d_arr_mul_19__24,d_arr_mul_19__23,
                            d_arr_mul_19__22,d_arr_mul_19__21,d_arr_mul_19__20,
                            d_arr_mul_19__19,d_arr_mul_19__18,d_arr_mul_19__17,
                            d_arr_mul_19__16,d_arr_mul_19__15,d_arr_mul_19__14,
                            d_arr_mul_19__13,d_arr_mul_19__12,d_arr_mul_19__11,
                            d_arr_mul_19__10,d_arr_mul_19__9,d_arr_mul_19__8,
                            d_arr_mul_19__7,d_arr_mul_19__6,d_arr_mul_19__5,
                            d_arr_mul_19__4,d_arr_mul_19__3,d_arr_mul_19__2,
                            d_arr_mul_19__1,d_arr_mul_19__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_20_mul_gen_mul_gen (.M (
                            {img_data_20__15,nx19440,img_data_20__13,
                            img_data_20__12,img_data_20__11,img_data_20__10,
                            img_data_20__9,img_data_20__8,img_data_20__7,
                            img_data_20__6,img_data_20__5,img_data_20__4,
                            img_data_20__3,img_data_20__2,img_data_20__1,
                            img_data_20__0}), .R ({filter_data_20__15,
                            filter_data_20__14,filter_data_20__13,
                            filter_data_20__12,filter_data_20__11,
                            filter_data_20__10,filter_data_20__9,
                            filter_data_20__8,filter_data_20__7,
                            filter_data_20__6,filter_data_20__5,
                            filter_data_20__4,filter_data_20__3,
                            filter_data_20__2,filter_data_20__1,
                            filter_data_20__0}), .cnt_enable (nx16643), .product (
                            {d_arr_mul_20__31,d_arr_mul_20__30,d_arr_mul_20__29,
                            d_arr_mul_20__28,d_arr_mul_20__27,d_arr_mul_20__26,
                            d_arr_mul_20__25,d_arr_mul_20__24,d_arr_mul_20__23,
                            d_arr_mul_20__22,d_arr_mul_20__21,d_arr_mul_20__20,
                            d_arr_mul_20__19,d_arr_mul_20__18,d_arr_mul_20__17,
                            d_arr_mul_20__16,d_arr_mul_20__15,d_arr_mul_20__14,
                            d_arr_mul_20__13,d_arr_mul_20__12,d_arr_mul_20__11,
                            d_arr_mul_20__10,d_arr_mul_20__9,d_arr_mul_20__8,
                            d_arr_mul_20__7,d_arr_mul_20__6,d_arr_mul_20__5,
                            d_arr_mul_20__4,d_arr_mul_20__3,d_arr_mul_20__2,
                            d_arr_mul_20__1,d_arr_mul_20__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_21_mul_gen_mul_gen (.M (
                            {img_data_21__15,nx19442,img_data_21__13,
                            img_data_21__12,img_data_21__11,img_data_21__10,
                            img_data_21__9,img_data_21__8,img_data_21__7,
                            img_data_21__6,img_data_21__5,img_data_21__4,
                            img_data_21__3,img_data_21__2,img_data_21__1,
                            img_data_21__0}), .R ({filter_data_21__15,
                            filter_data_21__14,filter_data_21__13,
                            filter_data_21__12,filter_data_21__11,
                            filter_data_21__10,filter_data_21__9,
                            filter_data_21__8,filter_data_21__7,
                            filter_data_21__6,filter_data_21__5,
                            filter_data_21__4,filter_data_21__3,
                            filter_data_21__2,filter_data_21__1,
                            filter_data_21__0}), .cnt_enable (nx16645), .product (
                            {d_arr_mul_21__31,d_arr_mul_21__30,d_arr_mul_21__29,
                            d_arr_mul_21__28,d_arr_mul_21__27,d_arr_mul_21__26,
                            d_arr_mul_21__25,d_arr_mul_21__24,d_arr_mul_21__23,
                            d_arr_mul_21__22,d_arr_mul_21__21,d_arr_mul_21__20,
                            d_arr_mul_21__19,d_arr_mul_21__18,d_arr_mul_21__17,
                            d_arr_mul_21__16,d_arr_mul_21__15,d_arr_mul_21__14,
                            d_arr_mul_21__13,d_arr_mul_21__12,d_arr_mul_21__11,
                            d_arr_mul_21__10,d_arr_mul_21__9,d_arr_mul_21__8,
                            d_arr_mul_21__7,d_arr_mul_21__6,d_arr_mul_21__5,
                            d_arr_mul_21__4,d_arr_mul_21__3,d_arr_mul_21__2,
                            d_arr_mul_21__1,d_arr_mul_21__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_22_mul_gen_mul_gen (.M (
                            {img_data_22__15,nx19444,img_data_22__13,
                            img_data_22__12,img_data_22__11,img_data_22__10,
                            img_data_22__9,img_data_22__8,img_data_22__7,
                            img_data_22__6,img_data_22__5,img_data_22__4,
                            img_data_22__3,img_data_22__2,img_data_22__1,
                            img_data_22__0}), .R ({filter_data_22__15,
                            filter_data_22__14,filter_data_22__13,
                            filter_data_22__12,filter_data_22__11,
                            filter_data_22__10,filter_data_22__9,
                            filter_data_22__8,filter_data_22__7,
                            filter_data_22__6,filter_data_22__5,
                            filter_data_22__4,filter_data_22__3,
                            filter_data_22__2,filter_data_22__1,
                            filter_data_22__0}), .cnt_enable (nx16645), .product (
                            {d_arr_mul_22__31,d_arr_mul_22__30,d_arr_mul_22__29,
                            d_arr_mul_22__28,d_arr_mul_22__27,d_arr_mul_22__26,
                            d_arr_mul_22__25,d_arr_mul_22__24,d_arr_mul_22__23,
                            d_arr_mul_22__22,d_arr_mul_22__21,d_arr_mul_22__20,
                            d_arr_mul_22__19,d_arr_mul_22__18,d_arr_mul_22__17,
                            d_arr_mul_22__16,d_arr_mul_22__15,d_arr_mul_22__14,
                            d_arr_mul_22__13,d_arr_mul_22__12,d_arr_mul_22__11,
                            d_arr_mul_22__10,d_arr_mul_22__9,d_arr_mul_22__8,
                            d_arr_mul_22__7,d_arr_mul_22__6,d_arr_mul_22__5,
                            d_arr_mul_22__4,d_arr_mul_22__3,d_arr_mul_22__2,
                            d_arr_mul_22__1,d_arr_mul_22__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_23_mul_gen_mul_gen (.M (
                            {img_data_23__15,nx19446,img_data_23__13,
                            img_data_23__12,img_data_23__11,img_data_23__10,
                            img_data_23__9,img_data_23__8,img_data_23__7,
                            img_data_23__6,img_data_23__5,img_data_23__4,
                            img_data_23__3,img_data_23__2,img_data_23__1,
                            img_data_23__0}), .R ({filter_data_23__15,
                            filter_data_23__14,filter_data_23__13,
                            filter_data_23__12,filter_data_23__11,
                            filter_data_23__10,filter_data_23__9,
                            filter_data_23__8,filter_data_23__7,
                            filter_data_23__6,filter_data_23__5,
                            filter_data_23__4,filter_data_23__3,
                            filter_data_23__2,filter_data_23__1,
                            filter_data_23__0}), .cnt_enable (nx16479), .product (
                            {d_arr_mul_23__31,d_arr_mul_23__30,d_arr_mul_23__29,
                            d_arr_mul_23__28,d_arr_mul_23__27,d_arr_mul_23__26,
                            d_arr_mul_23__25,d_arr_mul_23__24,d_arr_mul_23__23,
                            d_arr_mul_23__22,d_arr_mul_23__21,d_arr_mul_23__20,
                            d_arr_mul_23__19,d_arr_mul_23__18,d_arr_mul_23__17,
                            d_arr_mul_23__16,d_arr_mul_23__15,d_arr_mul_23__14,
                            d_arr_mul_23__13,d_arr_mul_23__12,d_arr_mul_23__11,
                            d_arr_mul_23__10,d_arr_mul_23__9,d_arr_mul_23__8,
                            d_arr_mul_23__7,d_arr_mul_23__6,d_arr_mul_23__5,
                            d_arr_mul_23__4,d_arr_mul_23__3,d_arr_mul_23__2,
                            d_arr_mul_23__1,d_arr_mul_23__0}), .clk (clk)) ;
    ModifiedBoothMultiplier mul_layer_gen_multipliers_gen_24_mul_gen_mul_gen (.M (
                            {img_data_24__15,img_data_24__14,img_data_24__13,
                            img_data_24__12,img_data_24__11,img_data_24__10,
                            img_data_24__9,img_data_24__8,img_data_24__7,
                            img_data_24__6,img_data_24__5,img_data_24__4,
                            img_data_24__3,img_data_24__2,img_data_24__1,
                            img_data_24__0}), .R ({filter_data_24__15,
                            filter_data_24__14,filter_data_24__13,
                            filter_data_24__12,filter_data_24__11,
                            filter_data_24__10,filter_data_24__9,
                            filter_data_24__8,filter_data_24__7,
                            filter_data_24__6,filter_data_24__5,
                            filter_data_24__4,filter_data_24__3,
                            filter_data_24__2,filter_data_24__1,
                            filter_data_24__0}), .cnt_enable (nx16481), .product (
                            {d_arr_mul_24__31,d_arr_mul_24__30,d_arr_mul_24__29,
                            d_arr_mul_24__28,d_arr_mul_24__27,d_arr_mul_24__26,
                            d_arr_mul_24__25,d_arr_mul_24__24,d_arr_mul_24__23,
                            d_arr_mul_24__22,d_arr_mul_24__21,d_arr_mul_24__20,
                            d_arr_mul_24__19,d_arr_mul_24__18,d_arr_mul_24__17,
                            d_arr_mul_24__16,d_arr_mul_24__15,d_arr_mul_24__14,
                            d_arr_mul_24__13,d_arr_mul_24__12,d_arr_mul_24__11,
                            d_arr_mul_24__10,d_arr_mul_24__9,d_arr_mul_24__8,
                            d_arr_mul_24__7,d_arr_mul_24__6,d_arr_mul_24__5,
                            d_arr_mul_24__4,d_arr_mul_24__3,d_arr_mul_24__2,
                            d_arr_mul_24__1,d_arr_mul_24__0}), .clk (clk)) ;
    NAdder_32 add_layer_gen_op9tree1_gen_loop_0_adder_gen (.a ({nx19448,nx16499,
              nx16503,nx16507,nx16511,nx16515,nx16519,nx16523,nx16527,nx16531,
              nx16535,nx16539,nx16543,nx16547,nx16551,nx16555,nx16559,nx16563,
              nx16567,nx16571,nx16575,nx16579,nx16583,nx16587,nx16591,nx16595,
              nx16599,nx16601,nx16603,q_arr_0__2,q_arr_0__1,nx16607}), .b ({
              q_arr_1__31,q_arr_1__30,q_arr_1__29,q_arr_1__28,nx19450,nx19454,
              q_arr_1__25,nx19458,q_arr_1__23,q_arr_1__22,q_arr_1__21,
              q_arr_1__20,q_arr_1__19,nx19462,nx19466,nx19470,q_arr_1__15,
              nx19474,q_arr_1__13,nx19476,q_arr_1__11,nx19478,q_arr_1__9,nx19482
              ,nx19486,q_arr_1__6,q_arr_1__5,q_arr_1__4,q_arr_1__3,q_arr_1__2,
              q_arr_1__1,q_arr_1__0}), .cin (GND0), .s ({d_arr_add_0__31,
              d_arr_add_0__30,d_arr_add_0__29,d_arr_add_0__28,d_arr_add_0__27,
              d_arr_add_0__26,d_arr_add_0__25,d_arr_add_0__24,d_arr_add_0__23,
              d_arr_add_0__22,d_arr_add_0__21,d_arr_add_0__20,d_arr_add_0__19,
              d_arr_add_0__18,d_arr_add_0__17,d_arr_add_0__16,d_arr_add_0__15,
              d_arr_add_0__14,d_arr_add_0__13,d_arr_add_0__12,d_arr_add_0__11,
              d_arr_add_0__10,d_arr_add_0__9,d_arr_add_0__8,d_arr_add_0__7,
              d_arr_add_0__6,d_arr_add_0__5,d_arr_add_0__4,d_arr_add_0__3,
              d_arr_add_0__2,d_arr_add_0__1,d_arr_add_0__0}), .cout (
              \$dummy [2690])) ;
    NAdder_32 add_layer_gen_op9tree1_gen_loop_1_adder_gen (.a ({q_arr_2__31,
              q_arr_2__30,q_arr_2__29,q_arr_2__28,q_arr_2__27,q_arr_2__26,
              q_arr_2__25,q_arr_2__24,q_arr_2__23,q_arr_2__22,q_arr_2__21,
              q_arr_2__20,q_arr_2__19,q_arr_2__18,q_arr_2__17,q_arr_2__16,
              q_arr_2__15,q_arr_2__14,q_arr_2__13,q_arr_2__12,q_arr_2__11,
              q_arr_2__10,q_arr_2__9,q_arr_2__8,q_arr_2__7,q_arr_2__6,q_arr_2__5
              ,q_arr_2__4,q_arr_2__3,q_arr_2__2,q_arr_2__1,q_arr_2__0}), .b ({
              q_arr_3__31,q_arr_3__30,q_arr_3__29,q_arr_3__28,q_arr_3__27,
              q_arr_3__26,q_arr_3__25,q_arr_3__24,q_arr_3__23,q_arr_3__22,
              q_arr_3__21,q_arr_3__20,q_arr_3__19,q_arr_3__18,q_arr_3__17,
              q_arr_3__16,q_arr_3__15,q_arr_3__14,q_arr_3__13,q_arr_3__12,
              q_arr_3__11,q_arr_3__10,q_arr_3__9,q_arr_3__8,q_arr_3__7,
              q_arr_3__6,q_arr_3__5,q_arr_3__4,q_arr_3__3,q_arr_3__2,q_arr_3__1,
              q_arr_3__0}), .cin (GND0), .s ({d_arr_add_1__31,d_arr_add_1__30,
              d_arr_add_1__29,d_arr_add_1__28,d_arr_add_1__27,d_arr_add_1__26,
              d_arr_add_1__25,d_arr_add_1__24,d_arr_add_1__23,d_arr_add_1__22,
              d_arr_add_1__21,d_arr_add_1__20,d_arr_add_1__19,d_arr_add_1__18,
              d_arr_add_1__17,d_arr_add_1__16,d_arr_add_1__15,d_arr_add_1__14,
              d_arr_add_1__13,d_arr_add_1__12,d_arr_add_1__11,d_arr_add_1__10,
              d_arr_add_1__9,d_arr_add_1__8,d_arr_add_1__7,d_arr_add_1__6,
              d_arr_add_1__5,d_arr_add_1__4,d_arr_add_1__3,d_arr_add_1__2,
              d_arr_add_1__1,d_arr_add_1__0}), .cout (\$dummy [2691])) ;
    NAdder_32 add_layer_gen_op9tree1_gen_loop_2_adder_gen (.a ({q_arr_4__31,
              q_arr_4__30,q_arr_4__29,q_arr_4__28,q_arr_4__27,q_arr_4__26,
              q_arr_4__25,q_arr_4__24,q_arr_4__23,q_arr_4__22,q_arr_4__21,
              q_arr_4__20,q_arr_4__19,q_arr_4__18,q_arr_4__17,q_arr_4__16,
              q_arr_4__15,q_arr_4__14,q_arr_4__13,q_arr_4__12,q_arr_4__11,
              q_arr_4__10,q_arr_4__9,q_arr_4__8,q_arr_4__7,q_arr_4__6,q_arr_4__5
              ,q_arr_4__4,q_arr_4__3,q_arr_4__2,q_arr_4__1,q_arr_4__0}), .b ({
              q_arr_5__31,q_arr_5__30,q_arr_5__29,q_arr_5__28,q_arr_5__27,
              q_arr_5__26,q_arr_5__25,q_arr_5__24,q_arr_5__23,q_arr_5__22,
              q_arr_5__21,q_arr_5__20,q_arr_5__19,q_arr_5__18,q_arr_5__17,
              q_arr_5__16,q_arr_5__15,q_arr_5__14,q_arr_5__13,q_arr_5__12,
              q_arr_5__11,q_arr_5__10,q_arr_5__9,q_arr_5__8,q_arr_5__7,
              q_arr_5__6,q_arr_5__5,q_arr_5__4,q_arr_5__3,q_arr_5__2,q_arr_5__1,
              q_arr_5__0}), .cin (GND0), .s ({d_arr_add_2__31,d_arr_add_2__30,
              d_arr_add_2__29,d_arr_add_2__28,d_arr_add_2__27,d_arr_add_2__26,
              d_arr_add_2__25,d_arr_add_2__24,d_arr_add_2__23,d_arr_add_2__22,
              d_arr_add_2__21,d_arr_add_2__20,d_arr_add_2__19,d_arr_add_2__18,
              d_arr_add_2__17,d_arr_add_2__16,d_arr_add_2__15,d_arr_add_2__14,
              d_arr_add_2__13,d_arr_add_2__12,d_arr_add_2__11,d_arr_add_2__10,
              d_arr_add_2__9,d_arr_add_2__8,d_arr_add_2__7,d_arr_add_2__6,
              d_arr_add_2__5,d_arr_add_2__4,d_arr_add_2__3,d_arr_add_2__2,
              d_arr_add_2__1,d_arr_add_2__0}), .cout (\$dummy [2692])) ;
    NAdder_32 add_layer_gen_op9tree1_gen_loop_3_adder_gen (.a ({q_arr_6__31,
              q_arr_6__30,q_arr_6__29,q_arr_6__28,q_arr_6__27,q_arr_6__26,
              q_arr_6__25,q_arr_6__24,q_arr_6__23,q_arr_6__22,q_arr_6__21,
              q_arr_6__20,q_arr_6__19,q_arr_6__18,q_arr_6__17,q_arr_6__16,
              q_arr_6__15,q_arr_6__14,q_arr_6__13,q_arr_6__12,q_arr_6__11,
              q_arr_6__10,q_arr_6__9,q_arr_6__8,q_arr_6__7,q_arr_6__6,q_arr_6__5
              ,q_arr_6__4,q_arr_6__3,q_arr_6__2,q_arr_6__1,q_arr_6__0}), .b ({
              q_arr_7__31,q_arr_7__30,q_arr_7__29,q_arr_7__28,q_arr_7__27,
              q_arr_7__26,q_arr_7__25,q_arr_7__24,q_arr_7__23,q_arr_7__22,
              q_arr_7__21,q_arr_7__20,q_arr_7__19,q_arr_7__18,q_arr_7__17,
              q_arr_7__16,q_arr_7__15,q_arr_7__14,q_arr_7__13,q_arr_7__12,
              q_arr_7__11,q_arr_7__10,q_arr_7__9,q_arr_7__8,q_arr_7__7,
              q_arr_7__6,q_arr_7__5,q_arr_7__4,q_arr_7__3,q_arr_7__2,q_arr_7__1,
              q_arr_7__0}), .cin (GND0), .s ({d_arr_add_3__31,d_arr_add_3__30,
              d_arr_add_3__29,d_arr_add_3__28,d_arr_add_3__27,d_arr_add_3__26,
              d_arr_add_3__25,d_arr_add_3__24,d_arr_add_3__23,d_arr_add_3__22,
              d_arr_add_3__21,d_arr_add_3__20,d_arr_add_3__19,d_arr_add_3__18,
              d_arr_add_3__17,d_arr_add_3__16,d_arr_add_3__15,d_arr_add_3__14,
              d_arr_add_3__13,d_arr_add_3__12,d_arr_add_3__11,d_arr_add_3__10,
              d_arr_add_3__9,d_arr_add_3__8,d_arr_add_3__7,d_arr_add_3__6,
              d_arr_add_3__5,d_arr_add_3__4,d_arr_add_3__3,d_arr_add_3__2,
              d_arr_add_3__1,d_arr_add_3__0}), .cout (\$dummy [2693])) ;
    NAdder_32 add_layer_gen_op9tree2_gen_loop_0_adder_gen (.a ({q_arr_9__31,
              q_arr_9__30,q_arr_9__29,q_arr_9__28,q_arr_9__27,q_arr_9__26,
              q_arr_9__25,q_arr_9__24,q_arr_9__23,q_arr_9__22,q_arr_9__21,
              q_arr_9__20,q_arr_9__19,q_arr_9__18,q_arr_9__17,q_arr_9__16,
              q_arr_9__15,q_arr_9__14,q_arr_9__13,q_arr_9__12,q_arr_9__11,
              q_arr_9__10,q_arr_9__9,q_arr_9__8,q_arr_9__7,q_arr_9__6,q_arr_9__5
              ,q_arr_9__4,q_arr_9__3,q_arr_9__2,q_arr_9__1,q_arr_9__0}), .b ({
              q_arr_10__31,q_arr_10__30,q_arr_10__29,q_arr_10__28,q_arr_10__27,
              q_arr_10__26,q_arr_10__25,q_arr_10__24,q_arr_10__23,q_arr_10__22,
              q_arr_10__21,q_arr_10__20,q_arr_10__19,q_arr_10__18,q_arr_10__17,
              q_arr_10__16,q_arr_10__15,q_arr_10__14,q_arr_10__13,q_arr_10__12,
              q_arr_10__11,q_arr_10__10,q_arr_10__9,q_arr_10__8,q_arr_10__7,
              q_arr_10__6,q_arr_10__5,q_arr_10__4,q_arr_10__3,q_arr_10__2,
              q_arr_10__1,q_arr_10__0}), .cin (GND0), .s ({d_arr_add_9__31,
              d_arr_add_9__30,d_arr_add_9__29,d_arr_add_9__28,d_arr_add_9__27,
              d_arr_add_9__26,d_arr_add_9__25,d_arr_add_9__24,d_arr_add_9__23,
              d_arr_add_9__22,d_arr_add_9__21,d_arr_add_9__20,d_arr_add_9__19,
              d_arr_add_9__18,d_arr_add_9__17,d_arr_add_9__16,d_arr_add_9__15,
              d_arr_add_9__14,d_arr_add_9__13,d_arr_add_9__12,d_arr_add_9__11,
              d_arr_add_9__10,d_arr_add_9__9,d_arr_add_9__8,d_arr_add_9__7,
              d_arr_add_9__6,d_arr_add_9__5,d_arr_add_9__4,d_arr_add_9__3,
              d_arr_add_9__2,d_arr_add_9__1,d_arr_add_9__0}), .cout (
              \$dummy [2694])) ;
    NAdder_32 add_layer_gen_op9tree2_gen_loop_1_adder_gen (.a ({q_arr_11__31,
              q_arr_11__30,q_arr_11__29,q_arr_11__28,q_arr_11__27,q_arr_11__26,
              q_arr_11__25,q_arr_11__24,q_arr_11__23,q_arr_11__22,q_arr_11__21,
              q_arr_11__20,q_arr_11__19,q_arr_11__18,q_arr_11__17,q_arr_11__16,
              q_arr_11__15,q_arr_11__14,q_arr_11__13,q_arr_11__12,q_arr_11__11,
              q_arr_11__10,q_arr_11__9,q_arr_11__8,q_arr_11__7,q_arr_11__6,
              q_arr_11__5,q_arr_11__4,q_arr_11__3,q_arr_11__2,q_arr_11__1,
              q_arr_11__0}), .b ({q_arr_12__31,q_arr_12__30,q_arr_12__29,
              q_arr_12__28,q_arr_12__27,q_arr_12__26,q_arr_12__25,q_arr_12__24,
              q_arr_12__23,q_arr_12__22,q_arr_12__21,q_arr_12__20,q_arr_12__19,
              q_arr_12__18,q_arr_12__17,q_arr_12__16,q_arr_12__15,q_arr_12__14,
              q_arr_12__13,q_arr_12__12,q_arr_12__11,q_arr_12__10,q_arr_12__9,
              q_arr_12__8,q_arr_12__7,q_arr_12__6,q_arr_12__5,q_arr_12__4,
              q_arr_12__3,q_arr_12__2,q_arr_12__1,q_arr_12__0}), .cin (GND0), .s (
              {d_arr_add_10__31,d_arr_add_10__30,d_arr_add_10__29,
              d_arr_add_10__28,d_arr_add_10__27,d_arr_add_10__26,
              d_arr_add_10__25,d_arr_add_10__24,d_arr_add_10__23,
              d_arr_add_10__22,d_arr_add_10__21,d_arr_add_10__20,
              d_arr_add_10__19,d_arr_add_10__18,d_arr_add_10__17,
              d_arr_add_10__16,d_arr_add_10__15,d_arr_add_10__14,
              d_arr_add_10__13,d_arr_add_10__12,d_arr_add_10__11,
              d_arr_add_10__10,d_arr_add_10__9,d_arr_add_10__8,d_arr_add_10__7,
              d_arr_add_10__6,d_arr_add_10__5,d_arr_add_10__4,d_arr_add_10__3,
              d_arr_add_10__2,d_arr_add_10__1,d_arr_add_10__0}), .cout (
              \$dummy [2695])) ;
    NAdder_32 add_layer_gen_op9tree2_gen_loop_2_adder_gen (.a ({q_arr_13__31,
              q_arr_13__30,q_arr_13__29,q_arr_13__28,q_arr_13__27,q_arr_13__26,
              q_arr_13__25,q_arr_13__24,q_arr_13__23,q_arr_13__22,q_arr_13__21,
              q_arr_13__20,q_arr_13__19,q_arr_13__18,q_arr_13__17,q_arr_13__16,
              q_arr_13__15,q_arr_13__14,q_arr_13__13,q_arr_13__12,q_arr_13__11,
              q_arr_13__10,q_arr_13__9,q_arr_13__8,q_arr_13__7,q_arr_13__6,
              q_arr_13__5,q_arr_13__4,q_arr_13__3,q_arr_13__2,q_arr_13__1,
              q_arr_13__0}), .b ({q_arr_14__31,q_arr_14__30,q_arr_14__29,
              q_arr_14__28,q_arr_14__27,q_arr_14__26,q_arr_14__25,q_arr_14__24,
              q_arr_14__23,q_arr_14__22,q_arr_14__21,q_arr_14__20,q_arr_14__19,
              q_arr_14__18,q_arr_14__17,q_arr_14__16,q_arr_14__15,q_arr_14__14,
              q_arr_14__13,q_arr_14__12,q_arr_14__11,q_arr_14__10,q_arr_14__9,
              q_arr_14__8,q_arr_14__7,q_arr_14__6,q_arr_14__5,q_arr_14__4,
              q_arr_14__3,q_arr_14__2,q_arr_14__1,q_arr_14__0}), .cin (GND0), .s (
              {d_arr_add_11__31,d_arr_add_11__30,d_arr_add_11__29,
              d_arr_add_11__28,d_arr_add_11__27,d_arr_add_11__26,
              d_arr_add_11__25,d_arr_add_11__24,d_arr_add_11__23,
              d_arr_add_11__22,d_arr_add_11__21,d_arr_add_11__20,
              d_arr_add_11__19,d_arr_add_11__18,d_arr_add_11__17,
              d_arr_add_11__16,d_arr_add_11__15,d_arr_add_11__14,
              d_arr_add_11__13,d_arr_add_11__12,d_arr_add_11__11,
              d_arr_add_11__10,d_arr_add_11__9,d_arr_add_11__8,d_arr_add_11__7,
              d_arr_add_11__6,d_arr_add_11__5,d_arr_add_11__4,d_arr_add_11__3,
              d_arr_add_11__2,d_arr_add_11__1,d_arr_add_11__0}), .cout (
              \$dummy [2696])) ;
    NAdder_32 add_layer_gen_op9tree2_gen_loop_3_adder_gen (.a ({q_arr_15__31,
              q_arr_15__30,q_arr_15__29,q_arr_15__28,q_arr_15__27,q_arr_15__26,
              q_arr_15__25,q_arr_15__24,q_arr_15__23,q_arr_15__22,q_arr_15__21,
              q_arr_15__20,q_arr_15__19,q_arr_15__18,q_arr_15__17,q_arr_15__16,
              q_arr_15__15,q_arr_15__14,q_arr_15__13,q_arr_15__12,q_arr_15__11,
              q_arr_15__10,q_arr_15__9,q_arr_15__8,q_arr_15__7,q_arr_15__6,
              q_arr_15__5,q_arr_15__4,q_arr_15__3,q_arr_15__2,q_arr_15__1,
              q_arr_15__0}), .b ({q_arr_16__31,q_arr_16__30,q_arr_16__29,
              q_arr_16__28,q_arr_16__27,q_arr_16__26,q_arr_16__25,q_arr_16__24,
              q_arr_16__23,q_arr_16__22,q_arr_16__21,q_arr_16__20,q_arr_16__19,
              q_arr_16__18,q_arr_16__17,q_arr_16__16,q_arr_16__15,q_arr_16__14,
              q_arr_16__13,q_arr_16__12,q_arr_16__11,q_arr_16__10,q_arr_16__9,
              q_arr_16__8,q_arr_16__7,q_arr_16__6,q_arr_16__5,q_arr_16__4,
              q_arr_16__3,q_arr_16__2,q_arr_16__1,q_arr_16__0}), .cin (GND0), .s (
              {d_arr_add_12__31,d_arr_add_12__30,d_arr_add_12__29,
              d_arr_add_12__28,d_arr_add_12__27,d_arr_add_12__26,
              d_arr_add_12__25,d_arr_add_12__24,d_arr_add_12__23,
              d_arr_add_12__22,d_arr_add_12__21,d_arr_add_12__20,
              d_arr_add_12__19,d_arr_add_12__18,d_arr_add_12__17,
              d_arr_add_12__16,d_arr_add_12__15,d_arr_add_12__14,
              d_arr_add_12__13,d_arr_add_12__12,d_arr_add_12__11,
              d_arr_add_12__10,d_arr_add_12__9,d_arr_add_12__8,d_arr_add_12__7,
              d_arr_add_12__6,d_arr_add_12__5,d_arr_add_12__4,d_arr_add_12__3,
              d_arr_add_12__2,d_arr_add_12__1,d_arr_add_12__0}), .cout (
              \$dummy [2697])) ;
    NAdder_32 add_layer_gen_op7tree1_gen_loop_0_adder_gen (.a ({q_arr_18__31,
              q_arr_18__30,q_arr_18__29,q_arr_18__28,nx19490,q_arr_18__26,
              q_arr_18__25,nx19494,q_arr_18__23,q_arr_18__22,q_arr_18__21,
              q_arr_18__20,q_arr_18__19,q_arr_18__18,q_arr_18__17,q_arr_18__16,
              q_arr_18__15,q_arr_18__14,q_arr_18__13,q_arr_18__12,q_arr_18__11,
              q_arr_18__10,q_arr_18__9,q_arr_18__8,q_arr_18__7,q_arr_18__6,
              q_arr_18__5,q_arr_18__4,q_arr_18__3,q_arr_18__2,q_arr_18__1,
              q_arr_18__0}), .b ({q_arr_19__31,q_arr_19__30,q_arr_19__29,
              q_arr_19__28,q_arr_19__27,q_arr_19__26,q_arr_19__25,q_arr_19__24,
              q_arr_19__23,q_arr_19__22,q_arr_19__21,q_arr_19__20,q_arr_19__19,
              q_arr_19__18,q_arr_19__17,q_arr_19__16,q_arr_19__15,q_arr_19__14,
              q_arr_19__13,q_arr_19__12,q_arr_19__11,q_arr_19__10,q_arr_19__9,
              q_arr_19__8,q_arr_19__7,q_arr_19__6,q_arr_19__5,q_arr_19__4,
              q_arr_19__3,q_arr_19__2,q_arr_19__1,q_arr_19__0}), .cin (GND0), .s (
              {d_arr_add_18__31,d_arr_add_18__30,d_arr_add_18__29,
              d_arr_add_18__28,d_arr_add_18__27,d_arr_add_18__26,
              d_arr_add_18__25,d_arr_add_18__24,d_arr_add_18__23,
              d_arr_add_18__22,d_arr_add_18__21,d_arr_add_18__20,
              d_arr_add_18__19,d_arr_add_18__18,d_arr_add_18__17,
              d_arr_add_18__16,d_arr_add_18__15,d_arr_add_18__14,
              d_arr_add_18__13,d_arr_add_18__12,d_arr_add_18__11,
              d_arr_add_18__10,d_arr_add_18__9,d_arr_add_18__8,d_arr_add_18__7,
              d_arr_add_18__6,d_arr_add_18__5,d_arr_add_18__4,d_arr_add_18__3,
              d_arr_add_18__2,d_arr_add_18__1,d_arr_add_18__0}), .cout (
              \$dummy [2698])) ;
    NAdder_32 add_layer_gen_op7tree1_gen_loop_1_adder_gen (.a ({q_arr_20__31,
              q_arr_20__30,q_arr_20__29,q_arr_20__28,q_arr_20__27,q_arr_20__26,
              q_arr_20__25,q_arr_20__24,q_arr_20__23,q_arr_20__22,q_arr_20__21,
              q_arr_20__20,q_arr_20__19,q_arr_20__18,q_arr_20__17,q_arr_20__16,
              q_arr_20__15,q_arr_20__14,q_arr_20__13,q_arr_20__12,q_arr_20__11,
              q_arr_20__10,q_arr_20__9,q_arr_20__8,q_arr_20__7,q_arr_20__6,
              q_arr_20__5,q_arr_20__4,q_arr_20__3,q_arr_20__2,q_arr_20__1,
              q_arr_20__0}), .b ({q_arr_21__31,q_arr_21__30,q_arr_21__29,
              q_arr_21__28,q_arr_21__27,q_arr_21__26,q_arr_21__25,q_arr_21__24,
              q_arr_21__23,q_arr_21__22,q_arr_21__21,q_arr_21__20,q_arr_21__19,
              q_arr_21__18,q_arr_21__17,q_arr_21__16,q_arr_21__15,q_arr_21__14,
              q_arr_21__13,q_arr_21__12,q_arr_21__11,q_arr_21__10,q_arr_21__9,
              q_arr_21__8,q_arr_21__7,q_arr_21__6,q_arr_21__5,q_arr_21__4,
              q_arr_21__3,q_arr_21__2,q_arr_21__1,q_arr_21__0}), .cin (GND0), .s (
              {d_arr_add_19__31,d_arr_add_19__30,d_arr_add_19__29,
              d_arr_add_19__28,d_arr_add_19__27,d_arr_add_19__26,
              d_arr_add_19__25,d_arr_add_19__24,d_arr_add_19__23,
              d_arr_add_19__22,d_arr_add_19__21,d_arr_add_19__20,
              d_arr_add_19__19,d_arr_add_19__18,d_arr_add_19__17,
              d_arr_add_19__16,d_arr_add_19__15,d_arr_add_19__14,
              d_arr_add_19__13,d_arr_add_19__12,d_arr_add_19__11,
              d_arr_add_19__10,d_arr_add_19__9,d_arr_add_19__8,d_arr_add_19__7,
              d_arr_add_19__6,d_arr_add_19__5,d_arr_add_19__4,d_arr_add_19__3,
              d_arr_add_19__2,d_arr_add_19__1,d_arr_add_19__0}), .cout (
              \$dummy [2699])) ;
    NAdder_32 add_layer_gen_op7tree1_gen_loop_2_adder_gen (.a ({q_arr_22__31,
              q_arr_22__30,q_arr_22__29,q_arr_22__28,q_arr_22__27,q_arr_22__26,
              q_arr_22__25,q_arr_22__24,q_arr_22__23,q_arr_22__22,q_arr_22__21,
              q_arr_22__20,q_arr_22__19,q_arr_22__18,q_arr_22__17,q_arr_22__16,
              q_arr_22__15,q_arr_22__14,q_arr_22__13,q_arr_22__12,q_arr_22__11,
              q_arr_22__10,q_arr_22__9,q_arr_22__8,q_arr_22__7,q_arr_22__6,
              q_arr_22__5,q_arr_22__4,q_arr_22__3,q_arr_22__2,q_arr_22__1,
              q_arr_22__0}), .b ({q_arr_23__31,q_arr_23__30,q_arr_23__29,
              q_arr_23__28,q_arr_23__27,q_arr_23__26,q_arr_23__25,q_arr_23__24,
              q_arr_23__23,q_arr_23__22,q_arr_23__21,q_arr_23__20,q_arr_23__19,
              q_arr_23__18,q_arr_23__17,q_arr_23__16,q_arr_23__15,q_arr_23__14,
              q_arr_23__13,q_arr_23__12,q_arr_23__11,q_arr_23__10,q_arr_23__9,
              q_arr_23__8,q_arr_23__7,q_arr_23__6,q_arr_23__5,q_arr_23__4,
              q_arr_23__3,q_arr_23__2,q_arr_23__1,q_arr_23__0}), .cin (GND0), .s (
              {d_arr_add_20__31,d_arr_add_20__30,d_arr_add_20__29,
              d_arr_add_20__28,d_arr_add_20__27,d_arr_add_20__26,
              d_arr_add_20__25,d_arr_add_20__24,d_arr_add_20__23,
              d_arr_add_20__22,d_arr_add_20__21,d_arr_add_20__20,
              d_arr_add_20__19,d_arr_add_20__18,d_arr_add_20__17,
              d_arr_add_20__16,d_arr_add_20__15,d_arr_add_20__14,
              d_arr_add_20__13,d_arr_add_20__12,d_arr_add_20__11,
              d_arr_add_20__10,d_arr_add_20__9,d_arr_add_20__8,d_arr_add_20__7,
              d_arr_add_20__6,d_arr_add_20__5,d_arr_add_20__4,d_arr_add_20__3,
              d_arr_add_20__2,d_arr_add_20__1,d_arr_add_20__0}), .cout (
              \$dummy [2700])) ;
    NAdder_32_unfolded2 merge_layer2_gen_adder1_gen (.a ({GND0,GND0,GND0,GND0,
                        GND0,GND0,nx19448,nx16501,nx16505,nx16509,nx16513,
                        nx16517,nx16521,nx16525,nx16529,nx16533,nx16537,nx16541,
                        nx16545,nx16549,nx16553,nx16557,nx16561,nx16565,nx16569,
                        nx16573,nx16577,nx16581,nx16585,nx16589,nx16593,nx16597}
                        ), .b ({output1_init[15],GND0,GND0,GND0,GND0,GND0,GND0,
                        GND0,GND0,GND0,GND0,GND0,GND0,GND0,GND0,GND0,GND0,
                        output1_init[14],output1_init[13],output1_init[12],
                        output1_init[11],output1_init[10],output1_init[9],
                        output1_init[8],output1_init[7],output1_init[6],
                        output1_init[5],output1_init[4],output1_init[3],
                        output1_init[2],output1_init[1],output1_init[0]}), .cin (
                        GND0), .s ({d_arr_merge2_0__31,\$dummy [2701],
                        \$dummy [2702],\$dummy [2703],\$dummy [2704],
                        d_arr_merge2_0__26,d_arr_merge2_0__25,d_arr_merge2_0__24
                        ,d_arr_merge2_0__23,d_arr_merge2_0__22,
                        d_arr_merge2_0__21,d_arr_merge2_0__20,d_arr_merge2_0__19
                        ,d_arr_merge2_0__18,d_arr_merge2_0__17,
                        d_arr_merge2_0__16,d_arr_merge2_0__15,d_arr_merge2_0__14
                        ,d_arr_merge2_0__13,d_arr_merge2_0__12,
                        d_arr_merge2_0__11,d_arr_merge2_0__10,d_arr_merge2_0__9,
                        d_arr_merge2_0__8,d_arr_merge2_0__7,d_arr_merge2_0__6,
                        d_arr_merge2_0__5,d_arr_merge2_0__4,d_arr_merge2_0__3,
                        d_arr_merge2_0__2,d_arr_merge2_0__1,d_arr_merge2_0__0})
                        , .cout (\$dummy [2705])) ;
    NAdder_32_unfolded2 merge_layer2_gen_adder2_gen (.a ({GND0,GND0,GND0,GND0,
                        GND0,GND0,q_arr_1__31,q_arr_1__30,q_arr_1__29,
                        q_arr_1__28,nx19452,nx19456,q_arr_1__25,nx19460,
                        q_arr_1__23,q_arr_1__22,q_arr_1__21,q_arr_1__20,
                        q_arr_1__19,nx19464,nx19468,nx19472,q_arr_1__15,nx19474,
                        q_arr_1__13,nx19476,q_arr_1__11,nx19480,q_arr_1__9,
                        nx19484,nx19486,q_arr_1__6}), .b ({output2_init[15],GND0
                        ,GND0,GND0,GND0,GND0,GND0,GND0,GND0,GND0,GND0,GND0,GND0,
                        GND0,GND0,GND0,GND0,output2_init[14],output2_init[13],
                        output2_init[12],output2_init[11],output2_init[10],
                        output2_init[9],output2_init[8],output2_init[7],
                        output2_init[6],output2_init[5],output2_init[4],
                        output2_init[3],output2_init[2],output2_init[1],
                        output2_init[0]}), .cin (GND0), .s ({d_arr_merge2_1__31,
                        \$dummy [2706],\$dummy [2707],\$dummy [2708],
                        \$dummy [2709],d_arr_merge2_1__26,d_arr_merge2_1__25,
                        d_arr_merge2_1__24,d_arr_merge2_1__23,d_arr_merge2_1__22
                        ,d_arr_merge2_1__21,d_arr_merge2_1__20,
                        d_arr_merge2_1__19,d_arr_merge2_1__18,d_arr_merge2_1__17
                        ,d_arr_merge2_1__16,d_arr_merge2_1__15,
                        d_arr_merge2_1__14,d_arr_merge2_1__13,d_arr_merge2_1__12
                        ,d_arr_merge2_1__11,d_arr_merge2_1__10,d_arr_merge2_1__9
                        ,d_arr_merge2_1__8,d_arr_merge2_1__7,d_arr_merge2_1__6,
                        d_arr_merge2_1__5,d_arr_merge2_1__4,d_arr_merge2_1__3,
                        d_arr_merge2_1__2,d_arr_merge2_1__1,d_arr_merge2_1__0})
                        , .cout (\$dummy [2710])) ;
    fake_gnd ix16087 (.Y (GND0)) ;
    nand02 ix201 (.Y (ready), .A0 (nx16276), .A1 (nx16625)) ;
    nand04 ix16277 (.Y (nx16276), .A0 (nx16278), .A1 (buffer_ready), .A2 (
           nx16375), .A3 (nx194)) ;
    oai21 ix16246 (.Y (nx16245), .A0 (nx16278), .A1 (nx16617), .B0 (nx16281)) ;
    nand03 ix16282 (.Y (nx16281), .A0 (counter_12), .A1 (nx16491), .A2 (nx16623)
           ) ;
    oai21 ix16236 (.Y (nx16235), .A0 (nx16285), .A1 (nx16617), .B0 (nx16289)) ;
    dffr reg_counter_12 (.Q (counter_12), .QB (nx16285), .D (nx16235), .CLK (
         nx16483), .R (nx16611)) ;
    nand03 ix16290 (.Y (nx16289), .A0 (counter_11), .A1 (nx16491), .A2 (nx16623)
           ) ;
    oai21 ix16226 (.Y (nx16225), .A0 (nx16293), .A1 (nx16617), .B0 (nx16295)) ;
    dffr reg_counter_11 (.Q (counter_11), .QB (nx16293), .D (nx16225), .CLK (
         nx16483), .R (nx16611)) ;
    nand03 ix16296 (.Y (nx16295), .A0 (counter_10), .A1 (nx16491), .A2 (nx16623)
           ) ;
    oai21 ix16216 (.Y (nx16215), .A0 (nx16299), .A1 (nx16617), .B0 (nx16301)) ;
    dffr reg_counter_10 (.Q (counter_10), .QB (nx16299), .D (nx16215), .CLK (
         nx16483), .R (nx16611)) ;
    nand03 ix16302 (.Y (nx16301), .A0 (counter_9), .A1 (nx16491), .A2 (nx16623)
           ) ;
    dffr reg_counter_9 (.Q (counter_9), .QB (\$dummy [2711]), .D (nx16205), .CLK (
         nx16487), .R (nx16615)) ;
    mux21_ni ix16206 (.Y (nx16205), .A0 (counter_9), .A1 (nx92), .S0 (nx16623)
             ) ;
    oai21 ix93 (.Y (nx92), .A0 (nx16306), .A1 (nx20), .B0 (nx16366)) ;
    dffr reg_counter_8 (.Q (\$dummy [2712]), .QB (nx16306), .D (nx16195), .CLK (
         nx16485), .R (nx16613)) ;
    oai21 ix16196 (.Y (nx16195), .A0 (nx16306), .A1 (nx16617), .B0 (nx16309)) ;
    nand03 ix16310 (.Y (nx16309), .A0 (counter_7), .A1 (nx16491), .A2 (nx16623)
           ) ;
    oai21 ix16186 (.Y (nx16185), .A0 (nx16313), .A1 (nx16617), .B0 (nx16315)) ;
    dffr reg_counter_7 (.Q (counter_7), .QB (nx16313), .D (nx16185), .CLK (
         nx16483), .R (nx16611)) ;
    nand03 ix16316 (.Y (nx16315), .A0 (counter_6), .A1 (nx16491), .A2 (nx16623)
           ) ;
    oai21 ix16176 (.Y (nx16175), .A0 (nx16319), .A1 (nx16617), .B0 (nx16321)) ;
    dffr reg_counter_6 (.Q (counter_6), .QB (nx16319), .D (nx16175), .CLK (
         nx16483), .R (nx16611)) ;
    nand03 ix16322 (.Y (nx16321), .A0 (counter_5), .A1 (nx16489), .A2 (nx16621)
           ) ;
    oai21 ix16166 (.Y (nx16165), .A0 (nx16325), .A1 (nx16619), .B0 (nx16327)) ;
    dffr reg_counter_5 (.Q (counter_5), .QB (nx16325), .D (nx16165), .CLK (
         nx16483), .R (nx16611)) ;
    nand03 ix16328 (.Y (nx16327), .A0 (counter_4), .A1 (nx16489), .A2 (nx16621)
           ) ;
    oai21 ix16156 (.Y (nx16155), .A0 (nx16331), .A1 (nx16619), .B0 (nx16333)) ;
    dffr reg_counter_4 (.Q (counter_4), .QB (nx16331), .D (nx16155), .CLK (
         nx16483), .R (nx16611)) ;
    nand03 ix16334 (.Y (nx16333), .A0 (counter_3), .A1 (nx16489), .A2 (nx16621)
           ) ;
    oai21 ix16146 (.Y (nx16145), .A0 (nx16337), .A1 (nx16619), .B0 (nx16339)) ;
    dffr reg_counter_3 (.Q (counter_3), .QB (nx16337), .D (nx16145), .CLK (
         nx16485), .R (nx16613)) ;
    nand03 ix16340 (.Y (nx16339), .A0 (counter_2), .A1 (nx16489), .A2 (nx16621)
           ) ;
    oai21 ix16136 (.Y (nx16135), .A0 (nx16343), .A1 (nx16619), .B0 (nx16345)) ;
    dffr reg_counter_2 (.Q (counter_2), .QB (nx16343), .D (nx16135), .CLK (
         nx16485), .R (nx16613)) ;
    nand03 ix16346 (.Y (nx16345), .A0 (counter_1), .A1 (nx16489), .A2 (nx16621)
           ) ;
    oai21 ix16126 (.Y (nx16125), .A0 (nx16349), .A1 (nx16619), .B0 (nx16351)) ;
    dffr reg_counter_1 (.Q (counter_1), .QB (nx16349), .D (nx16125), .CLK (
         nx16485), .R (nx16613)) ;
    nand03 ix16352 (.Y (nx16351), .A0 (nx16489), .A1 (counter_0), .A2 (nx16621)
           ) ;
    aoi21 ix16354 (.Y (nx16353), .A0 (operation), .A1 (counter_0), .B0 (nx20)) ;
    dffs_ni reg_counter_0 (.Q (counter_0), .QB (\$dummy [2713]), .D (nx16101), .CLK (
            nx16485), .S (nx16613)) ;
    nor02ii ix16102 (.Y (nx16101), .A0 (nx16619), .A1 (counter_0)) ;
    oai21 ix16116 (.Y (nx16115), .A0 (nx16361), .A1 (nx16619), .B0 (nx16363)) ;
    dffr reg_counter_14 (.Q (counter_14), .QB (nx16361), .D (nx16115), .CLK (
         nx16485), .R (nx16613)) ;
    nand03 ix16364 (.Y (nx16363), .A0 (nx16489), .A1 (counter_13), .A2 (nx16621)
           ) ;
    dffr reg_counter_13 (.Q (counter_13), .QB (nx16278), .D (nx16245), .CLK (
         nx16485), .R (nx16613)) ;
    nand02 ix16367 (.Y (nx16366), .A0 (operation), .A1 (counter_0)) ;
    oai21 ix153 (.Y (buffer_ready), .A0 (nx16481), .A1 (counter_0), .B0 (nx16625
          )) ;
    nand02 ix143 (.Y (sel_mul), .A0 (nx16371), .A1 (nx16373)) ;
    nor03_2x ix195 (.Y (nx194), .A0 (counter_14), .A1 (counter_15), .A2 (
             semi_ready)) ;
    oai21 ix16256 (.Y (nx16255), .A0 (nx16380), .A1 (nx16625), .B0 (nx16382)) ;
    dffr reg_counter_15 (.Q (counter_15), .QB (nx16380), .D (nx16255), .CLK (
         nx16487), .R (nx16615)) ;
    nand03 ix16383 (.Y (nx16382), .A0 (nx16491), .A1 (counter_14), .A2 (nx16625)
           ) ;
    dffr reg_counter_16 (.Q (semi_ready), .QB (\$dummy [2714]), .D (nx16265), .CLK (
         nx16487), .R (nx16615)) ;
    oai21 ix16266 (.Y (nx16265), .A0 (nx16386), .A1 (nx16388), .B0 (nx16390)) ;
    oai21 ix16387 (.Y (nx16386), .A0 (counter_15), .A1 (nx20), .B0 (nx16366)) ;
    inv02 ix16389 (.Y (nx16388), .A (en)) ;
    nand02 ix16391 (.Y (nx16390), .A0 (semi_ready), .A1 (nx16388)) ;
    inv01 ix159 (.Y (sel_add), .A (nx16375)) ;
    inv01 ix16398 (.Y (nx16399), .A (ordered_img_data_9__31)) ;
    inv02 ix16400 (.Y (nx16401), .A (nx16399)) ;
    inv02 ix16402 (.Y (nx16403), .A (nx16399)) ;
    inv02 ix16404 (.Y (nx16405), .A (nx16399)) ;
    inv01 ix16406 (.Y (nx16407), .A (ordered_img_data_10__31)) ;
    inv02 ix16408 (.Y (nx16409), .A (nx16407)) ;
    inv02 ix16410 (.Y (nx16411), .A (nx16407)) ;
    inv02 ix16412 (.Y (nx16413), .A (nx16407)) ;
    inv01 ix16414 (.Y (nx16415), .A (ordered_img_data_11__31)) ;
    inv02 ix16416 (.Y (nx16417), .A (nx16415)) ;
    inv02 ix16418 (.Y (nx16419), .A (nx16415)) ;
    inv02 ix16420 (.Y (nx16421), .A (nx16415)) ;
    inv01 ix16422 (.Y (nx16423), .A (ordered_img_data_12__31)) ;
    inv02 ix16424 (.Y (nx16425), .A (nx16423)) ;
    inv02 ix16426 (.Y (nx16427), .A (nx16423)) ;
    inv02 ix16428 (.Y (nx16429), .A (nx16423)) ;
    inv01 ix16430 (.Y (nx16431), .A (ordered_img_data_13__31)) ;
    inv02 ix16432 (.Y (nx16433), .A (nx16431)) ;
    inv02 ix16434 (.Y (nx16435), .A (nx16431)) ;
    inv02 ix16436 (.Y (nx16437), .A (nx16431)) ;
    inv01 ix16438 (.Y (nx16439), .A (ordered_img_data_14__31)) ;
    inv02 ix16440 (.Y (nx16441), .A (nx16439)) ;
    inv02 ix16442 (.Y (nx16443), .A (nx16439)) ;
    inv02 ix16444 (.Y (nx16445), .A (nx16439)) ;
    inv01 ix16446 (.Y (nx16447), .A (ordered_img_data_15__31)) ;
    inv02 ix16448 (.Y (nx16449), .A (nx16447)) ;
    inv02 ix16450 (.Y (nx16451), .A (nx16447)) ;
    inv02 ix16452 (.Y (nx16453), .A (nx16447)) ;
    inv01 ix16454 (.Y (nx16455), .A (ordered_img_data_16__31)) ;
    inv02 ix16456 (.Y (nx16457), .A (nx16455)) ;
    inv02 ix16458 (.Y (nx16459), .A (nx16455)) ;
    inv02 ix16460 (.Y (nx16461), .A (nx16455)) ;
    inv01 ix16462 (.Y (nx16463), .A (ordered_img_data_17__31)) ;
    inv02 ix16464 (.Y (nx16465), .A (nx16463)) ;
    inv02 ix16466 (.Y (nx16467), .A (nx16463)) ;
    inv02 ix16468 (.Y (nx16469), .A (nx16463)) ;
    inv01 ix16470 (.Y (nx16471), .A (sel_mul)) ;
    inv02 ix16472 (.Y (nx16473), .A (nx16651)) ;
    inv02 ix16474 (.Y (nx16475), .A (nx16651)) ;
    inv02 ix16476 (.Y (nx16477), .A (nx16651)) ;
    inv02 ix16478 (.Y (nx16479), .A (nx16651)) ;
    inv02 ix16480 (.Y (nx16481), .A (nx16651)) ;
    inv02 ix16482 (.Y (nx16483), .A (clk)) ;
    inv02 ix16484 (.Y (nx16485), .A (clk)) ;
    inv02 ix16486 (.Y (nx16487), .A (clk)) ;
    buf02 ix16488 (.Y (nx16489), .A (nx16353)) ;
    buf02 ix16490 (.Y (nx16491), .A (nx16353)) ;
    nor02_2x ix21 (.Y (nx20), .A0 (compute_relu), .A1 (nx16361)) ;
    and04 ix16372 (.Y (nx16371), .A0 (nx16349), .A1 (nx16343), .A2 (nx16337), .A3 (
          nx16331)) ;
    and04 ix16374 (.Y (nx16373), .A0 (nx16325), .A1 (nx16319), .A2 (nx16313), .A3 (
          nx16306)) ;
    and04 ix16376 (.Y (nx16375), .A0 (nx16497), .A1 (nx16299), .A2 (nx16293), .A3 (
          nx16285)) ;
    inv01 ix16496 (.Y (nx16497), .A (counter_9)) ;
    buf02 ix16498 (.Y (nx16499), .A (q_arr_0__30)) ;
    buf02 ix16500 (.Y (nx16501), .A (q_arr_0__30)) ;
    buf02 ix16502 (.Y (nx16503), .A (q_arr_0__29)) ;
    buf02 ix16504 (.Y (nx16505), .A (q_arr_0__29)) ;
    buf02 ix16506 (.Y (nx16507), .A (q_arr_0__28)) ;
    buf02 ix16508 (.Y (nx16509), .A (q_arr_0__28)) ;
    buf02 ix16510 (.Y (nx16511), .A (q_arr_0__27)) ;
    buf02 ix16512 (.Y (nx16513), .A (q_arr_0__27)) ;
    buf02 ix16514 (.Y (nx16515), .A (q_arr_0__26)) ;
    buf02 ix16516 (.Y (nx16517), .A (q_arr_0__26)) ;
    buf02 ix16518 (.Y (nx16519), .A (q_arr_0__25)) ;
    buf02 ix16520 (.Y (nx16521), .A (q_arr_0__25)) ;
    buf02 ix16522 (.Y (nx16523), .A (q_arr_0__24)) ;
    buf02 ix16524 (.Y (nx16525), .A (q_arr_0__24)) ;
    buf02 ix16526 (.Y (nx16527), .A (q_arr_0__23)) ;
    buf02 ix16528 (.Y (nx16529), .A (q_arr_0__23)) ;
    buf02 ix16530 (.Y (nx16531), .A (q_arr_0__22)) ;
    buf02 ix16532 (.Y (nx16533), .A (q_arr_0__22)) ;
    buf02 ix16534 (.Y (nx16535), .A (q_arr_0__21)) ;
    buf02 ix16536 (.Y (nx16537), .A (q_arr_0__21)) ;
    buf02 ix16538 (.Y (nx16539), .A (q_arr_0__20)) ;
    buf02 ix16540 (.Y (nx16541), .A (q_arr_0__20)) ;
    buf02 ix16542 (.Y (nx16543), .A (q_arr_0__19)) ;
    buf02 ix16544 (.Y (nx16545), .A (q_arr_0__19)) ;
    buf02 ix16546 (.Y (nx16547), .A (q_arr_0__18)) ;
    buf02 ix16548 (.Y (nx16549), .A (q_arr_0__18)) ;
    buf02 ix16550 (.Y (nx16551), .A (q_arr_0__17)) ;
    buf02 ix16552 (.Y (nx16553), .A (q_arr_0__17)) ;
    buf02 ix16554 (.Y (nx16555), .A (q_arr_0__16)) ;
    buf02 ix16556 (.Y (nx16557), .A (q_arr_0__16)) ;
    buf02 ix16558 (.Y (nx16559), .A (q_arr_0__15)) ;
    buf02 ix16560 (.Y (nx16561), .A (q_arr_0__15)) ;
    buf02 ix16562 (.Y (nx16563), .A (q_arr_0__14)) ;
    buf02 ix16564 (.Y (nx16565), .A (q_arr_0__14)) ;
    buf02 ix16566 (.Y (nx16567), .A (q_arr_0__13)) ;
    buf02 ix16568 (.Y (nx16569), .A (q_arr_0__13)) ;
    buf02 ix16570 (.Y (nx16571), .A (q_arr_0__12)) ;
    buf02 ix16572 (.Y (nx16573), .A (q_arr_0__12)) ;
    buf02 ix16574 (.Y (nx16575), .A (q_arr_0__11)) ;
    buf02 ix16576 (.Y (nx16577), .A (q_arr_0__11)) ;
    buf02 ix16578 (.Y (nx16579), .A (q_arr_0__10)) ;
    buf02 ix16580 (.Y (nx16581), .A (q_arr_0__10)) ;
    buf02 ix16582 (.Y (nx16583), .A (q_arr_0__9)) ;
    buf02 ix16584 (.Y (nx16585), .A (q_arr_0__9)) ;
    buf02 ix16586 (.Y (nx16587), .A (q_arr_0__8)) ;
    buf02 ix16588 (.Y (nx16589), .A (q_arr_0__8)) ;
    buf02 ix16590 (.Y (nx16591), .A (q_arr_0__7)) ;
    buf02 ix16592 (.Y (nx16593), .A (q_arr_0__7)) ;
    buf02 ix16594 (.Y (nx16595), .A (q_arr_0__6)) ;
    buf02 ix16596 (.Y (nx16597), .A (q_arr_0__6)) ;
    buf02 ix16598 (.Y (nx16599), .A (q_arr_0__5)) ;
    buf02 ix16600 (.Y (nx16601), .A (q_arr_0__4)) ;
    buf02 ix16602 (.Y (nx16603), .A (q_arr_0__3)) ;
    buf02 ix16604 (.Y (nx16605), .A (q_arr_0__0)) ;
    buf02 ix16606 (.Y (nx16607), .A (q_arr_0__0)) ;
    inv01 ix16608 (.Y (nx16609), .A (reset)) ;
    inv02 ix16610 (.Y (nx16611), .A (nx16609)) ;
    inv02 ix16612 (.Y (nx16613), .A (nx16609)) ;
    inv02 ix16614 (.Y (nx16615), .A (nx16609)) ;
    inv02 ix16616 (.Y (nx16617), .A (nx16388)) ;
    inv02 ix16618 (.Y (nx16619), .A (nx16388)) ;
    inv02 ix16620 (.Y (nx16621), .A (nx16388)) ;
    inv02 ix16622 (.Y (nx16623), .A (nx16388)) ;
    inv02 ix16624 (.Y (nx16625), .A (nx16388)) ;
    inv02 ix16626 (.Y (nx16627), .A (nx16653)) ;
    inv02 ix16628 (.Y (nx16629), .A (nx16653)) ;
    inv02 ix16630 (.Y (nx16631), .A (nx16653)) ;
    inv02 ix16632 (.Y (nx16633), .A (nx16653)) ;
    inv02 ix16634 (.Y (nx16635), .A (nx16653)) ;
    inv02 ix16636 (.Y (nx16637), .A (nx16471)) ;
    inv02 ix16638 (.Y (nx16639), .A (nx16471)) ;
    inv02 ix16640 (.Y (nx16641), .A (nx16471)) ;
    inv02 ix16642 (.Y (nx16643), .A (nx16471)) ;
    inv02 ix16644 (.Y (nx16645), .A (nx16471)) ;
    inv01 ix16650 (.Y (nx16651), .A (sel_mul)) ;
    inv01 ix16652 (.Y (nx16653), .A (sel_mul)) ;
    buf02 ix16658 (.Y (nx16659), .A (img_data_7__15)) ;
    buf02 ix16660 (.Y (nx16661), .A (img_data_11__15)) ;
    buf02 ix16662 (.Y (nx16663), .A (img_data_12__15)) ;
    buf02 ix16664 (.Y (nx16665), .A (filter_size)) ;
    buf02 ix16666 (.Y (nx16667), .A (filter_size)) ;
    buf02 ix19387 (.Y (nx19388), .A (q_arr_0__27)) ;
    buf02 ix19389 (.Y (nx19390), .A (q_arr_0__24)) ;
    buf02 ix19395 (.Y (nx19396), .A (img_data_0__14)) ;
    buf02 ix19397 (.Y (nx19398), .A (img_data_1__14)) ;
    buf02 ix19399 (.Y (nx19400), .A (img_data_1__14)) ;
    buf02 ix19401 (.Y (nx19402), .A (img_data_1__10)) ;
    buf02 ix19403 (.Y (nx19404), .A (img_data_2__14)) ;
    buf02 ix19405 (.Y (nx19406), .A (img_data_2__14)) ;
    buf02 ix19407 (.Y (nx19408), .A (img_data_2__10)) ;
    buf02 ix19409 (.Y (nx19410), .A (img_data_5__14)) ;
    buf02 ix19411 (.Y (nx19412), .A (img_data_6__14)) ;
    buf02 ix19413 (.Y (nx19414), .A (img_data_6__14)) ;
    buf02 ix19415 (.Y (nx19416), .A (img_data_6__10)) ;
    buf02 ix19417 (.Y (nx19418), .A (img_data_7__14)) ;
    buf02 ix19419 (.Y (nx19420), .A (img_data_7__14)) ;
    buf02 ix19421 (.Y (nx19422), .A (img_data_7__10)) ;
    buf02 ix19423 (.Y (nx19424), .A (img_data_10__14)) ;
    buf02 ix19425 (.Y (nx19426), .A (img_data_11__14)) ;
    buf02 ix19427 (.Y (nx19428), .A (img_data_11__14)) ;
    buf02 ix19429 (.Y (nx19430), .A (img_data_11__10)) ;
    buf02 ix19431 (.Y (nx19432), .A (img_data_12__14)) ;
    buf02 ix19433 (.Y (nx19434), .A (img_data_12__14)) ;
    buf02 ix19435 (.Y (nx19436), .A (img_data_12__10)) ;
    buf02 ix19437 (.Y (nx19438), .A (img_data_18__14)) ;
    buf02 ix19439 (.Y (nx19440), .A (img_data_20__14)) ;
    buf02 ix19441 (.Y (nx19442), .A (img_data_21__14)) ;
    buf02 ix19443 (.Y (nx19444), .A (img_data_22__14)) ;
    buf02 ix19445 (.Y (nx19446), .A (img_data_23__14)) ;
    buf02 ix19447 (.Y (nx19448), .A (q_arr_0__31)) ;
    buf02 ix19449 (.Y (nx19450), .A (q_arr_1__27)) ;
    buf02 ix19451 (.Y (nx19452), .A (q_arr_1__27)) ;
    buf02 ix19453 (.Y (nx19454), .A (q_arr_1__26)) ;
    buf02 ix19455 (.Y (nx19456), .A (q_arr_1__26)) ;
    buf02 ix19457 (.Y (nx19458), .A (q_arr_1__24)) ;
    buf02 ix19459 (.Y (nx19460), .A (q_arr_1__24)) ;
    buf02 ix19461 (.Y (nx19462), .A (q_arr_1__18)) ;
    buf02 ix19463 (.Y (nx19464), .A (q_arr_1__18)) ;
    buf02 ix19465 (.Y (nx19466), .A (q_arr_1__17)) ;
    buf02 ix19467 (.Y (nx19468), .A (q_arr_1__17)) ;
    buf02 ix19469 (.Y (nx19470), .A (q_arr_1__16)) ;
    buf02 ix19471 (.Y (nx19472), .A (q_arr_1__16)) ;
    buf02 ix19473 (.Y (nx19474), .A (q_arr_1__14)) ;
    buf02 ix19475 (.Y (nx19476), .A (q_arr_1__12)) ;
    buf02 ix19477 (.Y (nx19478), .A (q_arr_1__10)) ;
    buf02 ix19479 (.Y (nx19480), .A (q_arr_1__10)) ;
    buf02 ix19481 (.Y (nx19482), .A (q_arr_1__8)) ;
    buf02 ix19483 (.Y (nx19484), .A (q_arr_1__8)) ;
    buf02 ix19485 (.Y (nx19486), .A (q_arr_1__7)) ;
    buf02 ix19487 (.Y (nx19488), .A (q_arr_18__27)) ;
    buf02 ix19489 (.Y (nx19490), .A (q_arr_18__27)) ;
    buf02 ix19491 (.Y (nx19492), .A (q_arr_18__24)) ;
    buf02 ix19493 (.Y (nx19494), .A (q_arr_18__24)) ;
endmodule


module NAdder_32_unfolded2 ( a, b, cin, s, cout ) ;

    input [31:0]a ;
    input [31:0]b ;
    input cin ;
    output [31:0]s ;
    output cout ;

    wire nx131, nx149, nx165, nx181, nx197, nx213, nx229, nx245, nx263, nx275, 
         nx287, nx331, nx340, nx341, nx342, nx343, nx344, nx345, nx346, nx347, 
         nx348, nx349, nx350, nx351, nx352, nx353, nx354, nx355, nx356, nx357, 
         nx358, nx359, nx360, nx361, nx362, nx363, nx364, nx365, nx366, nx367, 
         nx160, nx368, nx16, nx369, nx141, nx133, nx370, nx371, nx372, nx373, 
         nx374, nx375, nx376, nx377, nx378, nx379, nx380, nx329, nx381, nx382, 
         nx383, nx384, nx385, nx386, nx387, nx311, nx388, nx389, nx144, nx390, 
         nx391, nx392, nx393, nx394, nx395, nx396, nx397, nx398, nx399, nx400, 
         nx401, nx402, nx403, nx404, nx327, nx405, nx406, nx407, nx408, nx409, 
         nx410, nx411, nx412, nx413, nx414, nx415, nx416, nx417, 
         nx329_XX0_XREP70, nx418, nx419, nx420, nx421, nx422, nx423, nx424, 
         nx425, nx128, nx426, nx427, nx249, nx255, nx112, nx237, nx428, nx429, 
         nx430, nx431, nx432, nx433, nx434, nx435, nx436, nx437, nx438, nx439, 
         nx440, nx441, nx266, nx442, nx443, nx444, nx445, nx446, nx447, nx448, 
         nx449, nx450, nx169, nx157, nx451, nx452, nx453, nx454, nx455, nx456, 
         nx457, nx458, nx459, nx460, nx461, nx462, nx233, nx463, nx464, nx465, 
         nx466, nx467, nx468, nx469, nx470, nx471, nx96, nx472, nx473, nx474, 
         nx475, nx476, nx477, nx478, nx201, nx205, nx479, nx480, nx481, nx482, 
         nx483, nx484, nx485, nx64, nx486, nx189, nx487, nx488, nx489, nx490, 
         nx491, nx492, nx493, nx494, nx495, nx185, nx496, nx173, nx497, nx498, 
         nx499, nx500, nx501, nx502, nx503, nx504, nx505, nx290, nx506, nx507, 
         nx508, nx509, nx510, nx511, nx512, nx513, nx514, nx515, nx299, nx516, 
         nx517, nx518, nx519, NOT_nx278, nx520, nx521, nx522, nx523, nx524, 
         nx525, nx526, nx527, nx528, nx529, nx530, nx531, nx32, nx532, nx533, 
         nx153, nx534, nx535, nx536, nx537, nx538, nx539, nx540, nx541, nx542, 
         nx543, nx544, nx545, nx546, nx547, nx548, nx549, nx550, nx551, nx552, 
         nx553, nx554, nx555, nx48, nx556, nx557, nx558, nx559, nx560, nx561, 
         nx562, nx563, nx564, nx565, nx566, NOT_nx302, nx567, nx568, nx569, 
         nx570, nx571, nx572, nx573, nx574, nx575, nx576, nx577, nx578, nx579, 
         nx580, nx581, nx582, nx583, nx584, nx585, nx586, nx587, nx588, nx589, 
         nx590, nx591, nx592, nx80, nx593, nx594, nx595, nx596, nx597, nx598, 
         nx137, nx599, nx600, nx601, nx602, nx603, nx604, nx605, nx606, nx607, 
         nx608, nx609, nx610, nx611, nx612, nx613, nx614, nx615, nx616, nx617, 
         nx618, nx619, nx620, nx621, nx622, nx623, nx909, nx911, nx913, nx915, 
         nx917, nx919, nx921, nx923, nx925, nx931, nx933, nx935, nx937, nx939, 
         nx941;



    assign s[30] = s[31] ;
    assign s[29] = s[31] ;
    assign s[28] = s[31] ;
    assign s[27] = s[31] ;
    fake_gnd ix73 (.Y (cout)) ;
    xor2 ix259 (.Y (s[0]), .A0 (a[0]), .A1 (b[0])) ;
    xor2 ix257 (.Y (s[1]), .A0 (nx131), .A1 (nx133)) ;
    nand02 ix132 (.Y (nx131), .A0 (b[0]), .A1 (a[0])) ;
    xor2 ix255 (.Y (s[2]), .A0 (nx925), .A1 (nx141)) ;
    xnor2 ix253 (.Y (s[3]), .A0 (nx16), .A1 (nx149)) ;
    xnor2_2x ix150 (.Y (nx149), .A0 (a[3]), .A1 (b[3])) ;
    xor2 ix251 (.Y (s[4]), .A0 (nx153), .A1 (nx157)) ;
    xnor2 ix249 (.Y (s[5]), .A0 (nx32), .A1 (nx165)) ;
    xnor2 ix166 (.Y (nx165), .A0 (a[5]), .A1 (b[5])) ;
    xor2 ix247 (.Y (s[6]), .A0 (nx169), .A1 (nx173)) ;
    xnor2 ix245 (.Y (s[7]), .A0 (nx48), .A1 (nx181)) ;
    xnor2 ix182 (.Y (nx181), .A0 (a[7]), .A1 (b[7])) ;
    xor2 ix243 (.Y (s[8]), .A0 (nx185), .A1 (nx189)) ;
    xnor2 ix241 (.Y (s[9]), .A0 (nx64), .A1 (nx197)) ;
    xnor2 ix198 (.Y (nx197), .A0 (a[9]), .A1 (b[9])) ;
    xor2 ix239 (.Y (s[10]), .A0 (nx201), .A1 (nx205)) ;
    xnor2 ix237 (.Y (s[11]), .A0 (nx80), .A1 (nx213)) ;
    xnor2 ix214 (.Y (nx213), .A0 (a[11]), .A1 (b[11])) ;
    xnor2 ix233 (.Y (s[13]), .A0 (nx96), .A1 (nx229)) ;
    xnor2 ix230 (.Y (nx229), .A0 (a[13]), .A1 (b[13])) ;
    xor2 ix231 (.Y (s[14]), .A0 (nx233), .A1 (nx237)) ;
    xnor2 ix229 (.Y (s[15]), .A0 (nx112), .A1 (nx245)) ;
    xnor2 ix246 (.Y (nx245), .A0 (a[15]), .A1 (nx935)) ;
    xor2 ix227 (.Y (s[16]), .A0 (nx249), .A1 (nx255)) ;
    xnor2 ix225 (.Y (s[17]), .A0 (nx128), .A1 (nx263)) ;
    xnor2 ix264 (.Y (nx263), .A0 (a[17]), .A1 (nx935)) ;
    xnor2 ix221 (.Y (s[19]), .A0 (nx144), .A1 (nx275)) ;
    xnor2 ix276 (.Y (nx275), .A0 (a[19]), .A1 (nx935)) ;
    xnor2 ix217 (.Y (s[21]), .A0 (nx160), .A1 (nx287)) ;
    xnor2 ix288 (.Y (nx287), .A0 (a[21]), .A1 (nx935)) ;
    inv02 ix330 (.Y (nx331), .A (b[31])) ;
    aoi21 ix624 (.Y (nx340), .A0 (nx933), .A1 (nx618), .B0 (nx311)) ;
    nor03_2x ix625 (.Y (nx341), .A0 (nx340), .A1 (nx620), .A2 (nx931)) ;
    nand02_2x ix626 (.Y (nx342), .A0 (a[23]), .A1 (nx935)) ;
    inv02 ix627 (.Y (nx343), .A (a[22])) ;
    oai21 ix628 (.Y (nx344), .A0 (a[23]), .A1 (a[22]), .B0 (nx935)) ;
    inv02 ix629 (.Y (nx345), .A (a[24])) ;
    inv02 ix630 (.Y (nx346), .A (a[25])) ;
    aoi22 ix631 (.Y (nx347), .A0 (nx620), .A1 (nx618), .B0 (nx345), .B1 (nx346)
          ) ;
    nand02_2x ix632 (.Y (nx348), .A0 (nx622), .A1 (nx931)) ;
    aoi422 ix633 (.Y (nx349), .A0 (nx618), .A1 (nx622), .A2 (nx933), .A3 (nx346)
           , .B0 (nx620), .B1 (nx345), .C0 (nx311), .C1 (nx348)) ;
    oai22 ix634 (.Y (nx350), .A0 (nx622), .A1 (nx345), .B0 (nx620), .B1 (nx933)
          ) ;
    nor02_2x ix635 (.Y (nx351), .A0 (nx935), .A1 (a[22])) ;
    inv02 ix636 (.Y (nx352), .A (a[21])) ;
    inv02 ix637 (.Y (nx353), .A (nx287)) ;
    nand02_2x ix638 (.Y (nx354), .A0 (a[20]), .A1 (nx353)) ;
    oai21 ix639 (.Y (nx355), .A0 (a[20]), .A1 (a[21]), .B0 (nx937)) ;
    aoi22 ix640 (.Y (nx356), .A0 (nx299), .A1 (nx342), .B0 (nx343), .B1 (nx618)
          ) ;
    inv02 ix641 (.Y (nx357), .A (nx343)) ;
    nor02_2x ix642 (.Y (nx358), .A0 (nx357), .A1 (nx937)) ;
    and02 ix643 (.Y (nx359), .A0 (nx516), .A1 (nx342)) ;
    nor03_2x ix644 (.Y (nx360), .A0 (nx358), .A1 (nx359), .A2 (nx344)) ;
    inv02 ix645 (.Y (nx361), .A (nx621)) ;
    inv02 ix646 (.Y (nx362), .A (nx345)) ;
    inv02 ix647 (.Y (nx363), .A (nx622)) ;
    inv02 ix648 (.Y (nx364), .A (nx933)) ;
    aoi22 ix649 (.Y (nx365), .A0 (nx361), .A1 (nx362), .B0 (nx363), .B1 (nx364)
          ) ;
    oai21 reg_s_24 (.Y (s[24]), .A0 (nx447), .A1 (nx365), .B0 (nx431)) ;
    nor02_2x ix650 (.Y (nx366), .A0 (nx937), .A1 (a[20])) ;
    inv02 ix651 (.Y (nx367), .A (a[20])) ;
    oai22 reg_nx160 (.Y (nx160), .A0 (nx366), .A1 (NOT_nx278), .B0 (nx618), .B1 (
          nx367)) ;
    nand02_2x ix652 (.Y (nx368), .A0 (b[3]), .A1 (a[3])) ;
    inv01 reg_nx16 (.Y (nx16), .A (nx451)) ;
    nor02_2x ix653 (.Y (nx369), .A0 (a[2]), .A1 (b[2])) ;
    ao21 reg_nx141 (.Y (nx141), .A0 (a[2]), .A1 (b[2]), .B0 (nx369)) ;
    ao21 reg_nx133 (.Y (nx133), .A0 (b[1]), .A1 (a[1]), .B0 (nx615)) ;
    inv02 ix654 (.Y (nx370), .A (nx341)) ;
    nand02_2x ix655 (.Y (nx371), .A0 (nx618), .A1 (nx354)) ;
    nand02_2x ix656 (.Y (nx372), .A0 (nx287), .A1 (nx352)) ;
    nand03_2x ix657 (.Y (nx373), .A0 (nx371), .A1 (nx356), .A2 (nx372)) ;
    or03 ix658 (.Y (nx374), .A0 (nx931), .A1 (nx933), .A2 (nx621)) ;
    aoi22 s_31_rename (.Y (s[31]), .A0 (nx370), .A1 (nx921), .B0 (nx374), .B1 (
          nx370)) ;
    aoi22 ix659 (.Y (nx375), .A0 (nx287), .A1 (nx352), .B0 (nx619), .B1 (nx354)
          ) ;
    inv02 ix660 (.Y (nx376), .A (a[18])) ;
    inv02 ix661 (.Y (nx377), .A (nx937)) ;
    aoi22 ix662 (.Y (nx378), .A0 (nx937), .A1 (nx376), .B0 (a[18]), .B1 (nx377)
          ) ;
    nand02_2x ix663 (.Y (nx379), .A0 (nx937), .A1 (a[19])) ;
    aoi21 ix664 (.Y (nx380), .A0 (nx355), .A1 (nx379), .B0 (nx373)) ;
    inv02 reg_nx329 (.Y (nx329), .A (nx937)) ;
    nor04_2x ix665 (.Y (nx381), .A0 (nx373), .A1 (nx275), .A2 (nx619), .A3 (
             nx376)) ;
    inv02 ix666 (.Y (nx382), .A (nx350)) ;
    inv02 ix667 (.Y (nx383), .A (nx931)) ;
    inv02 ix668 (.Y (nx384), .A (nx623)) ;
    aoi22 ix669 (.Y (nx385), .A0 (nx931), .A1 (nx623), .B0 (nx383), .B1 (nx384)
          ) ;
    or02 ix670 (.Y (nx386), .A0 (nx382), .A1 (nx385)) ;
    aoi222 ix671 (.Y (nx387), .A0 (nx931), .A1 (nx623), .B0 (nx383), .B1 (nx384)
           , .C0 (nx933), .C1 (nx939)) ;
    oai22 reg_nx311 (.Y (nx311), .A0 (nx383), .A1 (nx384), .B0 (nx931), .B1 (
          nx623)) ;
    and02 ix672 (.Y (nx388), .A0 (nx933), .A1 (nx939)) ;
    oai21 reg_s_25 (.Y (s[25]), .A0 (nx448), .A1 (nx386), .B0 (nx411)) ;
    and02 ix673 (.Y (nx389), .A0 (nx939), .A1 (a[18])) ;
    oai22 reg_nx144 (.Y (nx144), .A0 (nx378), .A1 (nx397), .B0 (nx619), .B1 (
          nx376)) ;
    inv02 ix674 (.Y (nx390), .A (nx263)) ;
    nor02_2x ix675 (.Y (nx391), .A0 (nx275), .A1 (nx378)) ;
    nor02ii ix676 (.Y (nx392), .A0 (nx329_XX0_XREP70), .A1 (a[17])) ;
    inv02 ix677 (.Y (nx393), .A (nx275)) ;
    nand02_2x ix678 (.Y (nx394), .A0 (nx389), .A1 (nx393)) ;
    nand02_2x ix679 (.Y (nx395), .A0 (nx379), .A1 (nx394)) ;
    inv01 ix680 (.Y (nx396), .A (nx375)) ;
    inv02 ix681 (.Y (nx397), .A (nx442)) ;
    nor03_2x ix682 (.Y (nx398), .A0 (nx380), .A1 (nx360), .A2 (nx381)) ;
    inv02 ix683 (.Y (nx399), .A (nx373)) ;
    inv01 ix684 (.Y (nx400), .A (nx378)) ;
    inv02 ix685 (.Y (nx401), .A (nx275)) ;
    nand03_2x ix686 (.Y (nx402), .A0 (nx399), .A1 (nx400), .A2 (nx401)) ;
    or02 ix687 (.Y (nx403), .A0 (nx621), .A1 (nx347)) ;
    and02 ix688 (.Y (nx404), .A0 (nx621), .A1 (nx349)) ;
    inv02 reg_nx327 (.Y (nx327), .A (nx621)) ;
    inv02 ix689 (.Y (nx405), .A (nx349)) ;
    oai21 reg_s_26 (.Y (s[26]), .A0 (nx921), .A1 (nx403), .B0 (nx446)) ;
    inv02 ix690 (.Y (nx406), .A (nx382)) ;
    inv02 ix691 (.Y (nx407), .A (nx311)) ;
    inv02 ix692 (.Y (nx408), .A (nx388)) ;
    aoi22 ix693 (.Y (nx409), .A0 (nx406), .A1 (nx407), .B0 (nx406), .B1 (nx408)
          ) ;
    ao21 ix694 (.Y (nx410), .A0 (nx311), .A1 (nx388), .B0 (nx387)) ;
    oai321 ix695 (.Y (nx411), .A0 (nx266), .A1 (nx409), .A2 (nx402), .B0 (nx409)
           , .B1 (nx398), .C0 (nx410)) ;
    nor02ii ix696 (.Y (nx412), .A0 (nx396), .A1 (nx391)) ;
    inv02 ix697 (.Y (nx413), .A (nx395)) ;
    nand02_2x ix698 (.Y (nx414), .A0 (nx355), .A1 (nx413)) ;
    inv02 ix699 (.Y (nx415), .A (nx396)) ;
    inv02 ix700 (.Y (nx416), .A (a[15])) ;
    inv02 ix701 (.Y (nx417), .A (a[16])) ;
    inv02 reg_nx329_XX0_XREP70 (.Y (nx329_XX0_XREP70), .A (nx939)) ;
    aoi21 ix702 (.Y (nx418), .A0 (nx416), .A1 (nx417), .B0 (nx329_XX0_XREP70)) ;
    nor02_2x ix703 (.Y (nx419), .A0 (a[14]), .A1 (b[14])) ;
    and02 ix704 (.Y (nx420), .A0 (a[14]), .A1 (b[14])) ;
    nor02_2x ix705 (.Y (nx421), .A0 (nx939), .A1 (a[16])) ;
    inv02 ix706 (.Y (nx422), .A (nx390)) ;
    inv02 ix707 (.Y (nx423), .A (nx391)) ;
    inv01 ix708 (.Y (nx424), .A (nx392)) ;
    oai21 ix709 (.Y (nx425), .A0 (nx392), .A1 (nx390), .B0 (nx391)) ;
    inv02 reg_nx128 (.Y (nx128), .A (nx527)) ;
    and02 ix710 (.Y (nx426), .A0 (a[15]), .A1 (nx939)) ;
    inv02 ix711 (.Y (nx427), .A (nx245)) ;
    oai32 reg_nx249 (.Y (nx249), .A0 (nx426), .A1 (nx462), .A2 (nx420), .B0 (
          nx427), .B1 (nx426)) ;
    oai22 reg_nx255 (.Y (nx255), .A0 (nx417), .A1 (nx329_XX0_XREP70), .B0 (nx939
          ), .B1 (a[16])) ;
    inv01 reg_nx112 (.Y (nx112), .A (nx459)) ;
    ao21 reg_nx237 (.Y (nx237), .A0 (a[14]), .A1 (b[14]), .B0 (nx419)) ;
    inv02 ix712 (.Y (nx428), .A (nx390)) ;
    inv02 ix713 (.Y (nx429), .A (nx392)) ;
    and02 ix714 (.Y (nx430), .A0 (nx365), .A1 (nx398)) ;
    oai321 ix715 (.Y (nx431), .A0 (nx527), .A1 (nx428), .A2 (nx402), .B0 (nx429)
           , .B1 (nx402), .C0 (nx430)) ;
    inv01 ix716 (.Y (nx432), .A (nx418)) ;
    aoi32 ix717 (.Y (nx433), .A0 (nx923), .A1 (nx429), .A2 (nx432), .B0 (nx429)
          , .B1 (nx428)) ;
    oai22 ix718 (.Y (nx434), .A0 (nx376), .A1 (nx377), .B0 (a[18]), .B1 (nx941)
          ) ;
    inv02 ix719 (.Y (nx435), .A (nx376)) ;
    inv02 ix720 (.Y (nx436), .A (nx377)) ;
    inv02 ix721 (.Y (nx437), .A (a[18])) ;
    inv02 ix722 (.Y (nx438), .A (nx941)) ;
    aoi22 ix723 (.Y (nx439), .A0 (nx435), .A1 (nx436), .B0 (nx437), .B1 (nx438)
          ) ;
    inv02 ix724 (.Y (nx440), .A (nx429)) ;
    inv02 ix725 (.Y (nx441), .A (nx428)) ;
    oai32 reg_nx266 (.Y (nx266), .A0 (nx482), .A1 (nx440), .A2 (nx909), .B0 (
          nx440), .B1 (nx441)) ;
    oai22 reg_s_18 (.Y (s[18]), .A0 (nx433), .A1 (nx434), .B0 (nx439), .B1 (
          nx266)) ;
    ao221 ix726 (.Y (nx442), .A0 (nx909), .A1 (nx441), .B0 (nx483), .B1 (nx441)
          , .C0 (nx440)) ;
    or02 ix727 (.Y (nx443), .A0 (nx428), .A1 (nx402)) ;
    nor02_2x ix728 (.Y (nx444), .A0 (nx545), .A1 (nx546)) ;
    and02 ix729 (.Y (nx445), .A0 (nx623), .A1 (nx405)) ;
    oai32 ix730 (.Y (nx446), .A0 (nx921), .A1 (nx445), .A2 (nx347), .B0 (nx445)
          , .B1 (nx404)) ;
    inv01 ix731 (.Y (nx447), .A (NOT_nx302)) ;
    inv01 ix732 (.Y (nx448), .A (nx921)) ;
    nand02_2x ix733 (.Y (nx449), .A0 (b[5]), .A1 (a[5])) ;
    nor02_2x ix734 (.Y (nx450), .A0 (a[4]), .A1 (b[4])) ;
    inv02 reg_nx169 (.Y (nx169), .A (nx497)) ;
    ao21 reg_nx157 (.Y (nx157), .A0 (a[4]), .A1 (b[4]), .B0 (nx450)) ;
    aoi22 ix735 (.Y (nx451), .A0 (a[2]), .A1 (b[2]), .B0 (nx609), .B1 (nx612)) ;
    inv01 ix736 (.Y (nx452), .A (nx909)) ;
    inv02 ix737 (.Y (nx453), .A (nx229)) ;
    nor03_2x ix738 (.Y (nx454), .A0 (nx419), .A1 (nx421), .A2 (nx245)) ;
    nor02_2x ix739 (.Y (nx455), .A0 (nx421), .A1 (nx245)) ;
    and02 ix740 (.Y (nx456), .A0 (b[13]), .A1 (a[13])) ;
    nor02_2x ix741 (.Y (nx457), .A0 (nx453), .A1 (nx911)) ;
    nor02_2x ix742 (.Y (nx458), .A0 (nx457), .A1 (nx419)) ;
    oai32 ix743 (.Y (nx459), .A0 (nx472), .A1 (nx911), .A2 (nx420), .B0 (nx458)
          , .B1 (nx420)) ;
    inv02 ix744 (.Y (nx460), .A (nx419)) ;
    nor02_2x ix745 (.Y (nx461), .A0 (nx229), .A1 (nx419)) ;
    ao22 ix746 (.Y (nx462), .A0 (nx460), .A1 (nx911), .B0 (nx473), .B1 (nx461)
         ) ;
    oai22 reg_nx233 (.Y (nx233), .A0 (nx911), .A1 (nx474), .B0 (nx453), .B1 (
          nx911)) ;
    or02 ix747 (.Y (nx463), .A0 (a[12]), .A1 (b[12])) ;
    or02 ix748 (.Y (nx464), .A0 (a[10]), .A1 (b[10])) ;
    and02 ix749 (.Y (nx465), .A0 (b[9]), .A1 (a[9])) ;
    nor02_2x ix750 (.Y (nx466), .A0 (a[10]), .A1 (b[10])) ;
    nor02_2x ix751 (.Y (nx467), .A0 (nx466), .A1 (nx197)) ;
    nor02_2x ix752 (.Y (nx468), .A0 (a[12]), .A1 (b[12])) ;
    aoi21 ix753 (.Y (nx469), .A0 (nx420), .A1 (nx455), .B0 (nx911)) ;
    nand02_2x ix754 (.Y (nx470), .A0 (nx420), .A1 (nx455)) ;
    oai21 ix755 (.Y (nx471), .A0 (nx453), .A1 (nx911), .B0 (nx454)) ;
    inv01 reg_nx96 (.Y (nx96), .A (nx551)) ;
    inv01 ix756 (.Y (nx472), .A (nx551)) ;
    inv01 ix757 (.Y (nx473), .A (nx551)) ;
    inv01 ix758 (.Y (nx474), .A (nx551)) ;
    nand02_2x ix759 (.Y (nx475), .A0 (b[11]), .A1 (a[11])) ;
    inv02 ix760 (.Y (nx476), .A (nx213)) ;
    aoi21 ix761 (.Y (nx477), .A0 (b[11]), .A1 (a[11]), .B0 (nx476)) ;
    inv02 ix762 (.Y (nx478), .A (nx197)) ;
    oai22 reg_nx201 (.Y (nx201), .A0 (nx465), .A1 (nx486), .B0 (nx478), .B1 (
          nx465)) ;
    ao21 reg_nx205 (.Y (nx205), .A0 (a[10]), .A1 (b[10]), .B0 (nx466)) ;
    or02 ix763 (.Y (nx479), .A0 (nx468), .A1 (nx213)) ;
    nor02_2x ix764 (.Y (nx480), .A0 (a[8]), .A1 (b[8])) ;
    and02 ix765 (.Y (nx481), .A0 (nx470), .A1 (nx471)) ;
    inv02 ix766 (.Y (nx482), .A (nx597)) ;
    inv02 ix767 (.Y (nx483), .A (nx923)) ;
    aoi22 ix768 (.Y (nx484), .A0 (a[10]), .A1 (b[10]), .B0 (nx464), .B1 (nx465)
          ) ;
    and02 ix769 (.Y (nx485), .A0 (a[8]), .A1 (b[8])) ;
    inv01 reg_nx64 (.Y (nx64), .A (nx565)) ;
    inv01 ix770 (.Y (nx486), .A (nx565)) ;
    ao21 reg_nx189 (.Y (nx189), .A0 (a[8]), .A1 (b[8]), .B0 (nx480)) ;
    inv02 ix771 (.Y (nx487), .A (b[6])) ;
    nand02_2x ix772 (.Y (nx488), .A0 (nx449), .A1 (nx487)) ;
    inv02 ix773 (.Y (nx489), .A (nx449)) ;
    nor02_2x ix774 (.Y (nx490), .A0 (b[6]), .A1 (a[6])) ;
    nor02_2x ix775 (.Y (nx491), .A0 (nx490), .A1 (nx165)) ;
    inv02 ix776 (.Y (nx492), .A (nx181)) ;
    inv02 ix777 (.Y (nx493), .A (nx468)) ;
    inv02 ix778 (.Y (nx494), .A (nx213)) ;
    nand02_2x ix779 (.Y (nx495), .A0 (b[7]), .A1 (a[7])) ;
    inv02 reg_nx185 (.Y (nx185), .A (nx595)) ;
    inv02 ix780 (.Y (nx496), .A (a[6])) ;
    oai22 reg_nx173 (.Y (nx173), .A0 (nx496), .A1 (nx487), .B0 (b[6]), .B1 (a[6]
          )) ;
    oai21 ix781 (.Y (nx497), .A0 (nx532), .A1 (nx165), .B0 (nx449)) ;
    inv02 ix782 (.Y (nx498), .A (nx619)) ;
    inv02 ix783 (.Y (nx499), .A (nx343)) ;
    inv02 ix784 (.Y (nx500), .A (nx941)) ;
    inv02 ix785 (.Y (nx501), .A (a[22])) ;
    aoi22 ix786 (.Y (nx502), .A0 (nx498), .A1 (nx499), .B0 (nx500), .B1 (nx501)
          ) ;
    nor02_2x ix787 (.Y (nx503), .A0 (nx290), .A1 (nx502)) ;
    ao21 reg_s_22 (.Y (s[22]), .A0 (nx290), .A1 (nx502), .B0 (nx503)) ;
    nand02_2x ix788 (.Y (nx504), .A0 (nx452), .A1 (nx923)) ;
    nor03_2x ix789 (.Y (nx505), .A0 (nx423), .A1 (nx422), .A2 (nx396)) ;
    aoi222 reg_nx290 (.Y (nx290), .A0 (nx414), .A1 (nx415), .B0 (nx392), .B1 (
           nx412), .C0 (nx504), .C1 (nx505)) ;
    inv02 ix790 (.Y (nx506), .A (nx619)) ;
    inv02 ix791 (.Y (nx507), .A (nx343)) ;
    nand02_2x ix792 (.Y (nx508), .A0 (nx506), .A1 (nx507)) ;
    inv02 ix793 (.Y (nx509), .A (a[23])) ;
    inv02 ix794 (.Y (nx510), .A (nx941)) ;
    aoi22 ix795 (.Y (nx511), .A0 (a[23]), .A1 (nx941), .B0 (nx509), .B1 (nx510)
          ) ;
    nand03_2x ix796 (.Y (nx512), .A0 (nx290), .A1 (nx508), .A2 (nx917)) ;
    or03 ix797 (.Y (nx513), .A0 (nx290), .A1 (nx917), .A2 (nx351)) ;
    nand03_2x ix798 (.Y (nx514), .A0 (nx917), .A1 (nx351), .A2 (nx508)) ;
    or03 ix799 (.Y (nx515), .A0 (nx917), .A1 (nx619), .A2 (nx343)) ;
    nand04_2x reg_s_23 (.Y (s[23]), .A0 (nx512), .A1 (nx513), .A2 (nx514), .A3 (
              nx515)) ;
    inv01 reg_nx299 (.Y (nx299), .A (nx511)) ;
    inv01 ix800 (.Y (nx516), .A (nx917)) ;
    inv02 ix801 (.Y (nx517), .A (nx425)) ;
    ao21 ix802 (.Y (nx518), .A0 (nx424), .A1 (nx452), .B0 (nx425)) ;
    nand02_2x ix803 (.Y (nx519), .A0 (nx413), .A1 (nx518)) ;
    aoi21 reg_NOT_nx278 (.Y (NOT_nx278), .A0 (nx547), .A1 (nx517), .B0 (nx519)
          ) ;
    inv02 ix804 (.Y (nx520), .A (nx941)) ;
    inv02 ix805 (.Y (nx521), .A (a[20])) ;
    inv02 ix806 (.Y (nx522), .A (nx619)) ;
    inv02 ix807 (.Y (nx523), .A (nx367)) ;
    aoi22 ix808 (.Y (nx524), .A0 (nx520), .A1 (nx521), .B0 (nx522), .B1 (nx523)
          ) ;
    nand02_2x ix809 (.Y (nx525), .A0 (NOT_nx278), .A1 (nx524)) ;
    oai21 reg_s_20 (.Y (s[20]), .A0 (NOT_nx278), .A1 (nx524), .B0 (nx525)) ;
    inv02 ix810 (.Y (nx526), .A (nx452)) ;
    nor02_2x ix811 (.Y (nx527), .A0 (nx526), .A1 (nx548)) ;
    nand02_2x ix812 (.Y (nx528), .A0 (nx610), .A1 (nx613)) ;
    inv02 ix813 (.Y (nx529), .A (nx608)) ;
    inv02 ix814 (.Y (nx530), .A (nx368)) ;
    nor02_2x ix815 (.Y (nx531), .A0 (nx530), .A1 (nx617)) ;
    aoi422 reg_nx32 (.Y (nx32), .A0 (nx528), .A1 (nx529), .A2 (nx368), .A3 (
           nx616), .B0 (nx450), .B1 (nx616), .C0 (nx149), .C1 (nx531)) ;
    inv02 ix816 (.Y (nx532), .A (nx32)) ;
    inv02 ix817 (.Y (nx533), .A (nx149)) ;
    oai32 reg_nx153 (.Y (nx153), .A0 (nx557), .A1 (nx530), .A2 (nx608), .B0 (
          nx533), .B1 (nx530)) ;
    inv02 ix818 (.Y (nx534), .A (nx481)) ;
    inv02 ix819 (.Y (nx535), .A (nx463)) ;
    inv02 ix820 (.Y (nx536), .A (b[11])) ;
    inv02 ix821 (.Y (nx537), .A (a[11])) ;
    inv02 ix822 (.Y (nx538), .A (a[12])) ;
    inv02 ix823 (.Y (nx539), .A (b[12])) ;
    oai321 ix824 (.Y (nx540), .A0 (nx535), .A1 (nx536), .A2 (nx537), .B0 (nx538)
           , .B1 (nx539), .C0 (nx469)) ;
    inv02 ix825 (.Y (nx541), .A (nx429)) ;
    inv02 ix826 (.Y (nx542), .A (nx402)) ;
    nand02_2x ix827 (.Y (nx543), .A0 (nx541), .A1 (nx542)) ;
    inv01 ix828 (.Y (nx544), .A (nx909)) ;
    inv02 ix829 (.Y (nx545), .A (nx398)) ;
    nor02_2x ix830 (.Y (nx546), .A0 (nx429), .A1 (nx402)) ;
    inv02 ix831 (.Y (nx547), .A (nx923)) ;
    inv02 ix832 (.Y (nx548), .A (nx923)) ;
    and03 ix833 (.Y (nx549), .A0 (nx463), .A1 (b[11]), .A2 (a[11])) ;
    and02 ix834 (.Y (nx550), .A0 (a[12]), .A1 (b[12])) ;
    nor03_2x ix835 (.Y (nx551), .A0 (nx549), .A1 (nx550), .A2 (nx554)) ;
    nand02_2x ix836 (.Y (nx552), .A0 (b[7]), .A1 (a[7])) ;
    inv02 ix837 (.Y (nx553), .A (nx480)) ;
    inv01 ix838 (.Y (nx554), .A (nx582)) ;
    inv02 ix839 (.Y (nx555), .A (nx491)) ;
    aoi22 reg_nx48 (.Y (nx48), .A0 (nx555), .A1 (nx567), .B0 (nx606), .B1 (nx567
          )) ;
    inv02 ix840 (.Y (nx556), .A (nx48)) ;
    and02 ix841 (.Y (nx557), .A0 (nx611), .A1 (nx614)) ;
    inv02 ix842 (.Y (nx558), .A (nx571)) ;
    inv02 ix843 (.Y (nx559), .A (nx484)) ;
    aoi21 ix844 (.Y (nx560), .A0 (a[12]), .A1 (b[12]), .B0 (nx468)) ;
    nand03_2x ix845 (.Y (nx561), .A0 (nx593), .A1 (nx475), .A2 (nx919)) ;
    inv02 ix846 (.Y (nx562), .A (nx475)) ;
    nor02_2x ix847 (.Y (nx563), .A0 (nx919), .A1 (nx913)) ;
    aoi22 ix848 (.Y (nx564), .A0 (nx562), .A1 (nx563), .B0 (nx913), .B1 (nx919)
          ) ;
    nand03_2x reg_s_12 (.Y (s[12]), .A0 (nx561), .A1 (nx589), .A2 (nx564)) ;
    nor02_2x ix849 (.Y (nx565), .A0 (nx594), .A1 (nx915)) ;
    and02 ix850 (.Y (nx566), .A0 (nx398), .A1 (nx544)) ;
    aoi32 reg_NOT_nx302 (.Y (NOT_nx302), .A0 (nx566), .A1 (nx923), .A2 (nx543), 
          .B0 (nx443), .B1 (nx444)) ;
    aoi22 ix851 (.Y (nx567), .A0 (a[6]), .A1 (nx488), .B0 (b[6]), .B1 (nx489)) ;
    nand02_2x ix852 (.Y (nx568), .A0 (nx553), .A1 (nx492)) ;
    oai22 ix853 (.Y (nx569), .A0 (nx480), .A1 (nx552), .B0 (nx567), .B1 (nx568)
          ) ;
    inv02 ix854 (.Y (nx570), .A (nx479)) ;
    inv02 ix855 (.Y (nx571), .A (nx467)) ;
    inv02 ix856 (.Y (nx572), .A (a[8])) ;
    inv02 ix857 (.Y (nx573), .A (b[8])) ;
    inv02 ix858 (.Y (nx574), .A (a[10])) ;
    inv02 ix859 (.Y (nx575), .A (b[10])) ;
    inv02 ix860 (.Y (nx576), .A (nx464)) ;
    inv02 ix861 (.Y (nx577), .A (nx465)) ;
    oai322 ix862 (.Y (nx578), .A0 (nx571), .A1 (nx572), .A2 (nx573), .B0 (nx574)
           , .B1 (nx575), .C0 (nx576), .C1 (nx577)) ;
    nand02_2x ix863 (.Y (nx579), .A0 (nx491), .A1 (nx467)) ;
    inv02 ix864 (.Y (nx580), .A (nx492)) ;
    nor04_2x ix865 (.Y (nx581), .A0 (nx579), .A1 (nx479), .A2 (nx580), .A3 (
             nx480)) ;
    aoi332 ix866 (.Y (nx582), .A0 (nx569), .A1 (nx467), .A2 (nx570), .B0 (nx578)
           , .B1 (nx493), .B2 (nx494), .C0 (nx607), .C1 (nx581)) ;
    nor02_2x ix867 (.Y (nx583), .A0 (nx559), .A1 (nx915)) ;
    nand03_2x ix868 (.Y (nx584), .A0 (nx583), .A1 (nx495), .A2 (nx556)) ;
    aoi21 ix869 (.Y (nx585), .A0 (nx495), .A1 (nx181), .B0 (nx480)) ;
    nor03_2x ix870 (.Y (nx586), .A0 (nx585), .A1 (nx559), .A2 (nx915)) ;
    nor02_2x ix871 (.Y (nx587), .A0 (nx558), .A1 (nx559)) ;
    nor04_2x ix872 (.Y (nx588), .A0 (nx586), .A1 (nx587), .A2 (nx919), .A3 (
             nx913)) ;
    nand02_2x ix873 (.Y (nx589), .A0 (nx584), .A1 (nx588)) ;
    inv02 ix874 (.Y (nx590), .A (nx495)) ;
    inv01 ix875 (.Y (nx591), .A (nx556)) ;
    nor04_2x ix876 (.Y (nx592), .A0 (nx559), .A1 (nx915), .A2 (nx590), .A3 (
             nx591)) ;
    nor03_2x reg_nx80 (.Y (nx80), .A0 (nx592), .A1 (nx586), .A2 (nx587)) ;
    inv02 ix877 (.Y (nx593), .A (nx80)) ;
    oai32 ix878 (.Y (nx594), .A0 (nx556), .A1 (nx480), .A2 (nx181), .B0 (nx480)
          , .B1 (nx495)) ;
    oai21 ix879 (.Y (nx595), .A0 (nx181), .A1 (nx556), .B0 (nx495)) ;
    inv01 ix880 (.Y (nx596), .A (nx582)) ;
    oai21 ix881 (.Y (nx597), .A0 (nx596), .A1 (nx540), .B0 (nx534)) ;
    or02 ix882 (.Y (nx598), .A0 (b[1]), .A1 (a[1])) ;
    aoi32 reg_nx137 (.Y (nx137), .A0 (nx598), .A1 (b[0]), .A2 (a[0]), .B0 (b[1])
          , .B1 (a[1])) ;
    nor02_2x ix883 (.Y (nx599), .A0 (a[2]), .A1 (b[2])) ;
    nor04_2x ix884 (.Y (nx600), .A0 (nx925), .A1 (nx599), .A2 (nx450), .A3 (
             nx149)) ;
    inv02 ix885 (.Y (nx601), .A (a[2])) ;
    inv02 ix886 (.Y (nx602), .A (b[2])) ;
    inv02 ix887 (.Y (nx603), .A (a[4])) ;
    inv02 ix888 (.Y (nx604), .A (b[4])) ;
    oai422 ix889 (.Y (nx605), .A0 (nx601), .A1 (nx602), .A2 (nx450), .A3 (nx149)
           , .B0 (nx368), .B1 (nx450), .C0 (nx603), .C1 (nx604)) ;
    nor02_2x ix890 (.Y (nx606), .A0 (nx600), .A1 (nx605)) ;
    inv01 ix891 (.Y (nx607), .A (nx606)) ;
    and02 ix892 (.Y (nx608), .A0 (a[2]), .A1 (b[2])) ;
    inv02 ix893 (.Y (nx609), .A (nx599)) ;
    inv02 ix894 (.Y (nx610), .A (nx599)) ;
    inv02 ix895 (.Y (nx611), .A (nx599)) ;
    inv01 ix896 (.Y (nx612), .A (nx137)) ;
    inv01 ix897 (.Y (nx613), .A (nx925)) ;
    inv01 ix898 (.Y (nx614), .A (nx925)) ;
    nor02_2x ix899 (.Y (nx615), .A0 (b[1]), .A1 (a[1])) ;
    nand02_2x ix900 (.Y (nx616), .A0 (a[4]), .A1 (b[4])) ;
    and02 ix901 (.Y (nx617), .A0 (a[4]), .A1 (b[4])) ;
    buf16 ix902 (.Y (nx618), .A (nx329)) ;
    buf16 ix903 (.Y (nx619), .A (nx329)) ;
    buf16 ix904 (.Y (nx620), .A (nx331)) ;
    buf16 ix905 (.Y (nx621), .A (nx331)) ;
    buf16 ix906 (.Y (nx622), .A (nx327)) ;
    buf16 ix907 (.Y (nx623), .A (nx327)) ;
    inv01 ix908 (.Y (nx909), .A (nx432)) ;
    buf02 ix910 (.Y (nx911), .A (nx456)) ;
    buf02 ix912 (.Y (nx913), .A (nx477)) ;
    buf02 ix914 (.Y (nx915), .A (nx485)) ;
    inv01 ix916 (.Y (nx917), .A (nx299)) ;
    buf02 ix918 (.Y (nx919), .A (nx560)) ;
    inv01 ix920 (.Y (nx921), .A (nx447)) ;
    inv02 ix922 (.Y (nx923), .A (nx482)) ;
    inv02 ix924 (.Y (nx925), .A (nx612)) ;
    inv02 ix930 (.Y (nx931), .A (nx346)) ;
    inv02 ix932 (.Y (nx933), .A (nx345)) ;
    inv02 ix934 (.Y (nx935), .A (nx331)) ;
    inv02 ix936 (.Y (nx937), .A (nx331)) ;
    inv02 ix938 (.Y (nx939), .A (nx331)) ;
    inv02 ix940 (.Y (nx941), .A (nx331)) ;
endmodule


module ModifiedBoothMultiplier ( M, R, cnt_enable, product, clk ) ;

    input [15:0]M ;
    input [15:0]R ;
    input cnt_enable ;
    output [31:0]product ;
    input clk ;

    wire aux_product_0, shifting_R_0, shifting_R_4, shifting_R_6, shifting_R_8, 
         shifting_R_10, shifting_R_12, shifting_R_14, shifting_R_16, nx30, nx40, 
         nx50, nx60, nx70, nx80, nx90, nx100, nx108, shifting_R_1, shifting_R_3, 
         shifting_R_5, shifting_R_7, shifting_R_9, shifting_R_11, shifting_R_13, 
         shifting_R_15, nx146, nx156, nx166, nx176, nx186, nx196, nx206, nx216, 
         nx228, nx254, positive_2M_1, nx258, nx268, nx270, aux_product_1, 
         negative_M_1, nx296, nx306, nx310, positive_M_1, nx338, nx350, nx354, 
         nx370, aux_product_2, positive_M_2, nx398, nx406, nx426, negative_M_2, 
         nx442, nx464, aux_product_3, positive_M_3, nx500, nx508, nx520, 
         negative_M_3, nx536, nx552, nx558, aux_product_4, positive_M_4, nx614, 
         negative_M_4, nx630, nx646, nx652, aux_product_5, positive_M_5, nx708, 
         negative_M_5, nx724, nx740, nx746, aux_product_6, positive_M_6, nx802, 
         negative_M_6, nx818, nx834, nx840, aux_product_7, positive_M_7, nx896, 
         negative_M_7, nx912, nx934, aux_product_8, positive_M_8, nx990, 
         negative_M_8, nx1006, nx1028, aux_product_9, positive_M_9, nx1084, 
         negative_M_9, nx1100, nx1122, aux_product_10, positive_M_10, nx1150, 
         nx1178, negative_M_10, nx1194, nx1216, aux_product_11, positive_M_11, 
         nx1272, negative_M_11, nx1288, nx1308, nx1310, aux_product_12, 
         positive_M_12, nx1366, negative_M_12, nx1382, nx1404, aux_product_13, 
         positive_M_13, nx1460, negative_M_13, nx1476, nx1498, aux_product_14, 
         positive_M_14, nx1526, nx1554, negative_M_14, nx1570, nx1592, 
         aux_product_15, positive_M_15, nx1616, nx1624, negative_M_15, nx1640, 
         nx1656, nx1660, nx1662, aux_product_16, positive_M_16, nx1694, 
         negative_M_16, nx1710, nx1726, nx1732, aux_product_17, positive_M_17, 
         nx1758, negative_M_17, nx1770, nx1792, aux_product_18, positive_M_18, 
         nx1818, negative_M_18, nx1830, nx1852, aux_product_19, positive_M_19, 
         nx1878, negative_M_19, nx1890, nx1906, nx1912, aux_product_20, 
         positive_M_20, nx1938, negative_M_20, nx1950, nx1966, nx1972, 
         aux_product_21, positive_M_21, nx1998, negative_M_21, nx2010, nx2026, 
         nx2032, aux_product_22, positive_M_22, nx2058, negative_M_22, nx2070, 
         nx2090, nx2092, aux_product_23, positive_M_23, nx2118, negative_M_23, 
         nx2130, aux_product_24, positive_M_24, nx2178, negative_M_24, nx2190, 
         nx2206, nx2210, aux_product_25, positive_M_25, nx2238, negative_M_25, 
         nx2250, nx2272, aux_product_26, positive_M_26, nx2298, negative_M_26, 
         nx2310, aux_product_27, positive_M_27, nx2358, negative_M_27, nx2370, 
         nx2386, nx2390, aux_product_28, positive_M_28, nx2418, negative_M_28, 
         nx2430, nx2446, aux_product_29, positive_M_29, nx2478, negative_M_29, 
         nx2490, nx2506, nx2510, aux_product_30, positive_2M_31, nx2538, 
         negative_2M_31, nx2550, nx2566, nx2570, aux_product_31, positive_M_31, 
         nx2598, negative_M_31, nx2610, nx2626, nx2630, nx3098, nx3108, nx3118, 
         nx3128, nx3138, nx3148, nx3158, nx3168, nx3178, nx3188, nx3198, nx3208, 
         nx3218, nx3228, nx3238, nx3248, nx3258, nx3268, nx3278, nx3288, nx3298, 
         nx3308, nx3318, nx3348, nx3368, nx3398, nx3421, nx3483, nx3487, nx3498, 
         nx3500, nx3508, nx3521, nx3523, nx3534, nx3540, nx3544, nx3550, nx3552, 
         nx3566, nx3568, nx3574, nx3576, nx3582, nx3591, nx3597, nx3601, nx3607, 
         nx3609, nx3615, nx3624, nx3627, nx3629, nx3635, nx3637, nx3643, nx3652, 
         nx3655, nx3657, nx3663, nx3665, nx3680, nx3683, nx3685, nx3691, nx3693, 
         nx3708, nx3711, nx3713, nx3719, nx3721, nx3736, nx3739, nx3741, nx3747, 
         nx3749, nx3764, nx3767, nx3769, nx3775, nx3777, nx3792, nx3795, nx3797, 
         nx3803, nx3805, nx3820, nx3823, nx3825, nx3831, nx3833, nx3848, nx3851, 
         nx3853, nx3859, nx3861, nx3873, nx3876, nx3879, nx3887, nx3889, nx3895, 
         nx3901, nx3904, nx3912, nx3914, nx3920, nx3924, nx3926, nx3928, nx3931, 
         nx3933, nx3943, nx3945, nx3955, nx3964, nx3966, nx3976, nx3985, nx3987, 
         nx3993, nx3997, nx4006, nx4008, nx4014, nx4018, nx4027, nx4029, nx4035, 
         nx4039, nx4048, nx4050, nx4060, nx4069, nx4081, nx4090, nx4098, nx4102, 
         nx4111, nx4113, nx4123, nx4132, nx4144, nx4153, nx4161, nx4165, nx4174, 
         nx4182, nx4186, nx4195, nx4203, nx4207, nx4216, nx4224, nx4237, nx4245, 
         nx4262, nx4268, nx4270, nx4272, nx4280, nx4284, nx4286, nx4288, nx4290, 
         nx4292, nx4294, nx4296, nx4298, nx4308, nx4310, nx4312, nx4314, nx4316, 
         nx4318, nx4320, nx4332, nx4348, nx4350, nx4352, nx4354, nx4376, nx4380, 
         nx4382, nx4384, nx4396, nx4398, nx4400, nx4402, nx4406, nx4410, nx4412, 
         nx4414, nx4416, nx4418, nx4420, nx4436, nx4438, nx4440, nx4442, nx4444, 
         nx4446, nx4448, nx4450, nx4456, nx4458, nx4460, nx4466, nx4468, nx4470, 
         nx4476, nx4480, nx4482, nx4484, nx4486, nx4488, nx4490, nx236, 
         nx4322_XX0_XREP40, nx4274, shifting_R_2, nx3454, nx3424, 
         nx4274_XX0_XREP44, nx884, nx790, nx4322, nx4478_XX0_XREP64, nx4580, 
         nx4581, nx4582, nx4583, nx4584, nx4585, nx4586, nx4587, nx4588, nx4589, 
         nx4590, nx4591, nx4592, nx4593, nx4594, nx4218, nx4595, nx4596, nx4597, 
         nx4598, nx4599, nx4600, nx4601, nx4602, nx4603, nx4604, nx4454, nx4605, 
         nx4606, nx4607, nx4608, nx4609, nx4610, nx4611, nx4612, nx4613, nx4614, 
         nx4615, nx4616, nx4617, nx4618, nx4619, nx4620, nx4304, nx4621, nx4622, 
         nx4623, nx4624, nx4625, nx4626, nx4627, nx4628, nx4629, nx4630, nx4631, 
         nx4632, nx4633, nx4634, nx4635, nx4074, nx4636, nx4637, nx4638, nx4639, 
         nx4640, nx4641, nx4642, nx4643, nx4644, nx4645, nx4646, nx4647, nx4648, 
         nx4649, nx4650, nx4651, nx4652, nx4653, nx3526, nx3492, nx4654, nx368, 
         nx4655, nx4656, nx4657, nx4658, nx4158, nx4659, nx4032, nx4660, nx4661, 
         nx4137, nx4662, nx3358, nx4663, nx4664, nx458, nx3529, nx4665, nx462, 
         nx4472, nx4462, nx4666, nx4667, nx4668, nx4669, nx4670, nx4671, nx4672, 
         nx4673, nx4674, nx4675, nx4676, nx4677, nx3990, nx3969, nx4678, nx4679, 
         nx4680, nx4681, nx4682, nx4683, nx3917, nx4684, nx4685, nx4686, nx4687, 
         nx3555, nx4688, nx4689, nx4690, nx4691, nx4692, nx4693, nx4694, nx4695, 
         nx4696, nx4697, nx4698, nx4699, nx4700, nx4701, nx4702, nx4703, nx4704, 
         nx4705, nx4706, nx4707, nx4708, nx3892, nx4709, nx3864, nx4710, nx4711, 
         nx4712, nx4713, nx4714, nx3579, nx4715, nx4716, nx556, nx4717, nx4718, 
         nx4719, nx4720, nx4721, nx4722, nx3948, nx4723, nx4724, nx4725, nx4726, 
         nx4727, nx4728, nx4729, nx4730, nx4731, nx4732, nx4733, nx4734, nx4735, 
         nx4736, nx4737, nx4738, nx4739, nx4740, nx4741, nx3808, nx3780, nx4742, 
         nx4743, nx4744, nx3612, nx4745, nx4746, nx4747, nx3752, nx4748, nx4749, 
         nx4750, nx4751, nx3724, nx3696, nx3668, nx4752, nx492, nx4753, nx4754, 
         nx4755, nx4756, nx4757, nx4758, nx4759, nx4760, nx4761, nx4762, nx4763, 
         nx4764, nx4765, nx4766, nx4767, nx4768, nx4769, nx876, nx4770, nx782, 
         nx4771, nx4772, nx696, nx688, nx4773, nx594, nx4774, nx4775, nx4776, 
         nx4777, nx4276, nx4264, nx4778, nx4779, nx928, nx3671, nx4780, nx4781, 
         nx4782, nx4783, nx4784, nx4785, nx4786, nx4787, nx3951, nx4788, nx4789, 
         nx1790, nx4790, nx4791, nx4792, nx4793, nx4794, nx4795, nx1850, nx4796, 
         nx4797, nx4798, nx4799, nx4800, nx4801, nx4802, nx4803, nx4804, nx4805, 
         nx4806, nx4807, nx4808, nx1910, nx4809, nx4810, nx4811, nx4812, nx4813, 
         nx4814, nx4815, nx4816, nx4817, nx4818, nx4819, nx4820, nx4821, nx4822, 
         nx4823, nx4824, nx4825, nx744, nx4826, nx650, nx838, nx4827, nx4828, 
         nx4829, nx4830, nx4831, nx602, nx4832, nx4833, nx4834, nx4835, nx4836, 
         nx4837, nx4838, nx1166, nx4839, nx4840, nx4841, nx1158, nx4842, nx4843, 
         nx4844, nx4845, nx4846, nx1072, nx4847, nx1064, nx4848, nx978, nx4849, 
         nx970, nx4850, nx4851, nx4852, nx4853, nx4854, nx4855, nx4856, nx4857, 
         nx4858, nx4859, nx4861, nx4862, nx1542, nx4863, nx4864, nx4865, nx4866, 
         nx4867, nx1534, nx4868, nx4869, nx1448, nx4870, nx1432, nx4871, nx4872, 
         nx1440, nx4873, nx4874, nx4875, nx1354, nx1346, nx4876, nx1260, nx1252, 
         nx4877, nx4878, nx1846, nx3972, nx4282, nx4478, nx4879, nx4880, nx4881, 
         nx4882, nx4883, nx4884, nx2270, nx4885, nx4886, nx4887, nx4888, nx4053, 
         nx4889, nx4890, nx4891, nx4892, nx4893, nx4894, nx4895, nx4896, nx4897, 
         nx4898, nx4899, nx4900, nx4901, nx4902, nx4903, nx4904, nx4905, nx4906, 
         nx4907, nx4908, nx4909, nx4910, nx4911, nx4221, nx4912, nx4913, nx4914, 
         nx4915, nx4916, nx4917, nx4918, nx4919, nx4920, nx4921, nx4922, nx4923, 
         nx4924, nx4925, nx4926, nx4927, nx1970, nx4928, nx4929, nx4930, nx2030, 
         nx4931, nx4932, nx4933, nx4934, nx4935, nx4936, nx4937, nx4938, nx4939, 
         nx4940, nx4941, nx4942, nx4943, nx4944, nx4945, nx4946, nx4947, nx4948, 
         nx3836, nx2326, nx4140, nx4949, nx4950, nx1210, nx3755, nx4951, nx4952, 
         nx4953, nx4954, nx1214, nx4955, nx4956, nx4957, nx4958, nx4959, nx4960, 
         nx4961, nx4962, nx4963, nx4964, nx4965, nx4966, nx4967, nx4968, nx4011, 
         nx4969, nx4970, nx4971, nx4155, nx4972, nx4973, nx4974, nx4975, nx1056, 
         nx4976, nx868, nx4977, nx4978, nx4979, nx4980, nx4981, nx4982, nx4983, 
         nx4984, nx4985, nx4986, nx4987, nx4988, nx3378, nx2146, nx4077, nx3408, 
         nx4989, nx4266, nx4990, nx4991, nx1398, nx3811, nx4992, nx4993, nx4994, 
         nx4995, nx1402, nx4996, nx4997, nx4998, nx4999, nx4474, nx4464, nx4278, 
         nx5000, nx1116, nx5001, nx5002, nx5003, nx5004, nx5005, nx5006, nx5007, 
         nx3699, nx5008, nx1026, nx5009, nx5010, nx5011, nx5012, nx5013, nx5014, 
         nx5015, nx1120, nx5016, nx5017, nx5018, nx5019, nx5020, nx2150, nx5021, 
         nx5022, nx5023, nx5024, nx5025, nx5026, nx5027, nx5028, nx5029, nx5030, 
         nx5031, nx5032, nx5033, nx5034, nx5035, nx5036, nx5037, nx5038, nx5039, 
         nx5040, nx5041, nx5042, nx5043, nx1022, nx5044, nx5045, nx5046, nx5047, 
         nx5048, nx5049, nx5050, nx5051, nx5052, nx5053, nx4119, nx5054, nx5055, 
         nx5056, nx5057, nx5058, nx5059, nx5060, nx5061, nx5062, nx932, nx5063, 
         nx1586, nx3867, nx5064, nx5065, nx5066, nx5067, nx1492, nx3839, nx5068, 
         nx5069, nx5070, nx5071, nx5072, nx1590, nx5073, nx5074, nx1496, nx5075, 
         nx5076, nx5077, nx5078, nx1304, nx5079, nx3640, nx5080, nx5081, nx5082, 
         nx5083, nx5084, nx5085, nx5086, nx3388, nx5087, nx5088, nx5089, nx5090, 
         nx5091, nx5092, nx5093, nx5094, nx5095, nx3783, nx5096, nx5097, nx5098, 
         nx5099, nx5100, nx5101, nx5102, nx5103, nx5104, nx5105, nx5106, nx5107, 
         nx5108, nx5109, nx5110, nx5111, nx5112, nx5113, nx5114, nx5115, nx5116, 
         nx5117, nx5118, nx5119, nx5120, nx5121, nx5122, nx3328, nx5123, nx5124, 
         nx5125, nx5126, nx5127, nx5128, nx5129, nx5130, nx5131, nx5132, nx5133, 
         nx5134, nx5135, nx5136, nx5137, nx5138, nx5139, nx5140, nx5141, nx5142, 
         nx5143, nx5144, nx5145, nx5146, nx5147, nx5148, nx5149, nx5150, nx5151, 
         nx5152, nx2450, nx1786, nx5153, nx4116, nx5154, nx5155, nx5156, nx5157, 
         nx5158, nx5159, nx5160, nx4302, nx5161, nx5162, nx5163, nx3338, nx4452, 
         nx5164, nx5165, nx5166, nx5167, nx5168, nx5169, nx5170, nx5171, nx5172, 
         nx5173, nx5174, nx5175, nx5176, nx5177, nx2330, nx5178, nx5179, nx5180, 
         nx2086, nx4056, nx5181, nx5182, nx5183, nx1730, nx5184, nx5185, nx5186, 
         nx5187, nx5188, nx5189, nx5190, nx5191, nx5192, nx5193, nx5194, nx5195, 
         nx5196, nx5197, nx5198, nx5199, nx5200, nx5201, nx5202, nx5203, nx5204, 
         nx5205, nx5206, nx5207, nx5208, nx5209, nx5210, nx5211, nx5212, nx5213, 
         nx5214, nx5215, nx5216, nx5217, nx5218, nx5219, nx5220, nx5221, nx5222, 
         nx5223, nx5224, nx5225, nx5226, nx5227, nx5228, nx5229, nx5230, nx5231, 
         nx5232, nx5233, nx5234, nx5235, nx5236, nx5237, nx5238, nx5239, nx5240, 
         nx5241, nx5905, nx5907, nx5909, nx5911, nx5913, nx5915, nx5917, nx5919, 
         nx5921, nx5923, nx5925, nx5927, nx5929, nx5931, nx5933, nx5935, nx5937, 
         nx5939, nx5941, nx5943, nx5945, nx5947, nx5949, nx5951, nx5953, nx5955, 
         nx5957, nx5959, nx5961, nx5971, nx5973, nx5975, nx5977, nx5979, nx5981, 
         nx5983, nx5985, nx5987, nx5989, nx5991, nx5993, nx5995, nx5997, nx5999, 
         nx6001, nx6003, nx6005, nx6007, nx6009;
    wire [80:0] \$dummy ;




    dff reg_product_0 (.Q (product[0]), .QB (\$dummy [0]), .D (aux_product_0), .CLK (
        clk)) ;
    oai21 ix3099 (.Y (nx3098), .A0 (nx3421), .A1 (nx4288), .B0 (nx3483)) ;
    dff reg_aux_product_0 (.Q (aux_product_0), .QB (nx3421), .D (nx3098), .CLK (
        clk)) ;
    nand04 ix255 (.Y (nx254), .A0 (nx3424), .A1 (nx4322), .A2 (nx4440), .A3 (
           nx5208)) ;
    dff reg_shifting_R_1 (.Q (shifting_R_1), .QB (\$dummy [1]), .D (nx216), .CLK (
        clk)) ;
    mux21_ni ix217 (.Y (nx216), .A0 (R[0]), .A1 (shifting_R_3), .S0 (nx4438)) ;
    dff reg_shifting_R_3 (.Q (shifting_R_3), .QB (\$dummy [2]), .D (nx206), .CLK (
        clk)) ;
    mux21_ni ix207 (.Y (nx206), .A0 (R[2]), .A1 (shifting_R_5), .S0 (nx4436)) ;
    dff reg_shifting_R_5 (.Q (shifting_R_5), .QB (\$dummy [3]), .D (nx196), .CLK (
        clk)) ;
    mux21_ni ix197 (.Y (nx196), .A0 (R[4]), .A1 (shifting_R_7), .S0 (nx4436)) ;
    dff reg_shifting_R_7 (.Q (shifting_R_7), .QB (\$dummy [4]), .D (nx186), .CLK (
        clk)) ;
    mux21_ni ix187 (.Y (nx186), .A0 (R[6]), .A1 (shifting_R_9), .S0 (nx4436)) ;
    dff reg_shifting_R_9 (.Q (shifting_R_9), .QB (\$dummy [5]), .D (nx176), .CLK (
        clk)) ;
    mux21_ni ix177 (.Y (nx176), .A0 (R[8]), .A1 (shifting_R_11), .S0 (nx4436)) ;
    dff reg_shifting_R_11 (.Q (shifting_R_11), .QB (\$dummy [6]), .D (nx166), .CLK (
        clk)) ;
    mux21_ni ix167 (.Y (nx166), .A0 (R[10]), .A1 (shifting_R_13), .S0 (nx4436)
             ) ;
    dff reg_shifting_R_13 (.Q (shifting_R_13), .QB (\$dummy [7]), .D (nx156), .CLK (
        clk)) ;
    mux21_ni ix157 (.Y (nx156), .A0 (R[12]), .A1 (shifting_R_15), .S0 (nx4436)
             ) ;
    dff reg_shifting_R_15 (.Q (shifting_R_15), .QB (\$dummy [8]), .D (nx146), .CLK (
        clk)) ;
    nor02ii ix147 (.Y (nx146), .A0 (nx4436), .A1 (R[14])) ;
    dff reg_shifting_R_0 (.Q (shifting_R_0), .QB (\$dummy [9]), .D (nx108), .CLK (
        clk)) ;
    mux21_ni ix101 (.Y (nx100), .A0 (R[1]), .A1 (shifting_R_4), .S0 (nx4440)) ;
    dff reg_shifting_R_4 (.Q (shifting_R_4), .QB (\$dummy [10]), .D (nx90), .CLK (
        clk)) ;
    mux21_ni ix91 (.Y (nx90), .A0 (R[3]), .A1 (shifting_R_6), .S0 (nx4440)) ;
    dff reg_shifting_R_6 (.Q (shifting_R_6), .QB (\$dummy [11]), .D (nx80), .CLK (
        clk)) ;
    mux21_ni ix81 (.Y (nx80), .A0 (R[5]), .A1 (shifting_R_8), .S0 (nx4438)) ;
    dff reg_shifting_R_8 (.Q (shifting_R_8), .QB (\$dummy [12]), .D (nx70), .CLK (
        clk)) ;
    mux21_ni ix71 (.Y (nx70), .A0 (R[7]), .A1 (shifting_R_10), .S0 (nx4438)) ;
    dff reg_shifting_R_10 (.Q (shifting_R_10), .QB (\$dummy [13]), .D (nx60), .CLK (
        clk)) ;
    mux21_ni ix61 (.Y (nx60), .A0 (R[9]), .A1 (shifting_R_12), .S0 (nx4438)) ;
    dff reg_shifting_R_12 (.Q (shifting_R_12), .QB (\$dummy [14]), .D (nx50), .CLK (
        clk)) ;
    mux21_ni ix51 (.Y (nx50), .A0 (R[11]), .A1 (shifting_R_14), .S0 (nx4438)) ;
    dff reg_shifting_R_14 (.Q (shifting_R_14), .QB (\$dummy [15]), .D (nx40), .CLK (
        clk)) ;
    mux21_ni ix41 (.Y (nx40), .A0 (R[13]), .A1 (shifting_R_16), .S0 (nx4438)) ;
    dff reg_shifting_R_16 (.Q (shifting_R_16), .QB (\$dummy [16]), .D (nx30), .CLK (
        clk)) ;
    nor02ii ix31 (.Y (nx30), .A0 (nx4438), .A1 (R[15])) ;
    nand04 ix3484 (.Y (nx3483), .A0 (nx270), .A1 (nx4440), .A2 (nx3492), .A3 (
           nx4288)) ;
    or02 ix271 (.Y (nx270), .A0 (nx268), .A1 (aux_product_0)) ;
    dff reg_positive_2M_1 (.Q (positive_2M_1), .QB (nx3487), .D (nx258), .CLK (
        clk)) ;
    dff reg_product_1 (.Q (product[1]), .QB (\$dummy [17]), .D (aux_product_1), 
        .CLK (clk)) ;
    oai21 ix3109 (.Y (nx3108), .A0 (nx3498), .A1 (nx4288), .B0 (nx3500)) ;
    dff reg_aux_product_1 (.Q (aux_product_1), .QB (nx3498), .D (nx3108), .CLK (
        clk)) ;
    nand03 ix3501 (.Y (nx3500), .A0 (nx4440), .A1 (nx370), .A2 (nx4288)) ;
    xnor2 ix371 (.Y (nx370), .A0 (nx3492), .A1 (nx368)) ;
    dff reg_positive_M_1 (.Q (positive_M_1), .QB (nx3508), .D (nx354), .CLK (clk
        )) ;
    nor02ii ix355 (.Y (nx354), .A0 (nx4440), .A1 (nx6003)) ;
    dff reg_negative_M_1 (.Q (negative_M_1), .QB (\$dummy [18]), .D (nx310), .CLK (
        clk)) ;
    nor02ii ix311 (.Y (nx310), .A0 (nx4440), .A1 (nx306)) ;
    aoi21 ix307 (.Y (nx306), .A0 (nx6003), .A1 (nx6007), .B0 (nx296)) ;
    nor02_2x ix297 (.Y (nx296), .A0 (nx6007), .A1 (nx6003)) ;
    dff reg_product_2 (.Q (product[2]), .QB (\$dummy [19]), .D (aux_product_2), 
        .CLK (clk)) ;
    oai21 ix3119 (.Y (nx3118), .A0 (nx3521), .A1 (nx4288), .B0 (nx3523)) ;
    dff reg_aux_product_2 (.Q (aux_product_2), .QB (nx3521), .D (nx3118), .CLK (
        clk)) ;
    nand03 ix3524 (.Y (nx3523), .A0 (nx4442), .A1 (nx464), .A2 (nx4288)) ;
    xnor2 ix465 (.Y (nx464), .A0 (nx3526), .A1 (nx462)) ;
    dff reg_negative_M_2 (.Q (negative_M_2), .QB (\$dummy [20]), .D (nx442), .CLK (
        clk)) ;
    mux21_ni ix443 (.Y (nx442), .A0 (nx406), .A1 (positive_2M_1), .S0 (nx4442)
             ) ;
    aoi21 ix407 (.Y (nx406), .A0 (nx3534), .A1 (nx5999), .B0 (nx398)) ;
    nor03_2x ix399 (.Y (nx398), .A0 (nx5999), .A1 (nx6007), .A2 (nx6003)) ;
    dff reg_positive_M_2 (.Q (positive_M_2), .QB (nx3544), .D (nx426), .CLK (clk
        )) ;
    oai21 ix427 (.Y (nx426), .A0 (nx4484), .A1 (nx3487), .B0 (nx3540)) ;
    oai21 ix3541 (.Y (nx3540), .A0 (nx350), .A1 (nx4482), .B0 (nx5999)) ;
    nor02_2x ix351 (.Y (nx350), .A0 (M[15]), .A1 (nx4442)) ;
    dff reg_product_3 (.Q (product[3]), .QB (\$dummy [21]), .D (aux_product_3), 
        .CLK (clk)) ;
    oai21 ix3129 (.Y (nx3128), .A0 (nx3550), .A1 (nx4288), .B0 (nx3552)) ;
    dff reg_aux_product_3 (.Q (aux_product_3), .QB (nx3550), .D (nx3128), .CLK (
        clk)) ;
    nand03 ix3553 (.Y (nx3552), .A0 (nx4442), .A1 (nx558), .A2 (nx4290)) ;
    xnor2 ix559 (.Y (nx558), .A0 (nx3555), .A1 (nx556)) ;
    dff reg_negative_M_3 (.Q (negative_M_3), .QB (\$dummy [22]), .D (nx536), .CLK (
        clk)) ;
    mux21_ni ix537 (.Y (nx536), .A0 (nx500), .A1 (negative_M_1), .S0 (nx4442)) ;
    xnor2 ix501 (.Y (nx500), .A0 (nx5997), .A1 (nx398)) ;
    dff reg_positive_M_3 (.Q (positive_M_3), .QB (nx3568), .D (nx520), .CLK (clk
        )) ;
    oai21 ix521 (.Y (nx520), .A0 (nx4484), .A1 (nx3508), .B0 (nx3566)) ;
    oai21 ix3567 (.Y (nx3566), .A0 (nx350), .A1 (nx4482), .B0 (nx5997)) ;
    dff reg_product_4 (.Q (product[4]), .QB (\$dummy [23]), .D (aux_product_4), 
        .CLK (clk)) ;
    oai21 ix3139 (.Y (nx3138), .A0 (nx3574), .A1 (nx4290), .B0 (nx3576)) ;
    dff reg_aux_product_4 (.Q (aux_product_4), .QB (nx3574), .D (nx3138), .CLK (
        clk)) ;
    nand03 ix3577 (.Y (nx3576), .A0 (nx4442), .A1 (nx652), .A2 (nx4290)) ;
    xnor2 ix653 (.Y (nx652), .A0 (nx3579), .A1 (nx650)) ;
    aoi221 ix3583 (.Y (nx3582), .A0 (negative_M_4), .A1 (nx4264), .B0 (
           positive_M_4), .B1 (nx4276), .C0 (nx646)) ;
    dff reg_negative_M_4 (.Q (negative_M_4), .QB (\$dummy [24]), .D (nx630), .CLK (
        clk)) ;
    mux21_ni ix631 (.Y (nx630), .A0 (nx594), .A1 (negative_M_2), .S0 (nx4442)) ;
    dff reg_positive_M_4 (.Q (positive_M_4), .QB (nx3601), .D (nx614), .CLK (clk
        )) ;
    oai322 ix615 (.Y (nx614), .A0 (nx3591), .A1 (nx5210), .A2 (nx4348), .B0 (
           nx3597), .B1 (nx4352), .C0 (nx4484), .C1 (nx3544)) ;
    nor02ii ix3592 (.Y (nx3591), .A0 (nx508), .A1 (nx594)) ;
    nor04 ix509 (.Y (nx508), .A0 (nx5997), .A1 (nx5999), .A2 (nx6007), .A3 (
          nx6003)) ;
    inv01 ix3598 (.Y (nx3597), .A (M[4])) ;
    dff reg_product_5 (.Q (product[5]), .QB (\$dummy [25]), .D (aux_product_5), 
        .CLK (clk)) ;
    oai21 ix3149 (.Y (nx3148), .A0 (nx3607), .A1 (nx4290), .B0 (nx3609)) ;
    dff reg_aux_product_5 (.Q (aux_product_5), .QB (nx3607), .D (nx3148), .CLK (
        clk)) ;
    nand03 ix3610 (.Y (nx3609), .A0 (nx4444), .A1 (nx746), .A2 (nx4290)) ;
    xnor2 ix747 (.Y (nx746), .A0 (nx3612), .A1 (nx744)) ;
    aoi221 ix3616 (.Y (nx3615), .A0 (negative_M_5), .A1 (nx4264), .B0 (
           positive_M_5), .B1 (nx4276), .C0 (nx740)) ;
    dff reg_negative_M_5 (.Q (negative_M_5), .QB (\$dummy [26]), .D (nx724), .CLK (
        clk)) ;
    mux21_ni ix725 (.Y (nx724), .A0 (nx688), .A1 (negative_M_3), .S0 (nx4444)) ;
    dff reg_positive_M_5 (.Q (positive_M_5), .QB (nx3629), .D (nx708), .CLK (clk
        )) ;
    oai322 ix709 (.Y (nx708), .A0 (nx3624), .A1 (nx696), .A2 (nx4348), .B0 (
           nx3627), .B1 (nx4352), .C0 (nx4484), .C1 (nx3568)) ;
    nor02ii ix3625 (.Y (nx3624), .A0 (nx5210), .A1 (nx4773)) ;
    inv01 ix3628 (.Y (nx3627), .A (M[5])) ;
    dff reg_product_6 (.Q (product[6]), .QB (\$dummy [27]), .D (aux_product_6), 
        .CLK (clk)) ;
    oai21 ix3159 (.Y (nx3158), .A0 (nx3635), .A1 (nx4290), .B0 (nx3637)) ;
    dff reg_aux_product_6 (.Q (aux_product_6), .QB (nx3635), .D (nx3158), .CLK (
        clk)) ;
    nand03 ix3638 (.Y (nx3637), .A0 (nx4444), .A1 (nx840), .A2 (nx4290)) ;
    xnor2 ix841 (.Y (nx840), .A0 (nx3640), .A1 (nx838)) ;
    aoi221 ix3644 (.Y (nx3643), .A0 (negative_M_6), .A1 (nx4264), .B0 (
           positive_M_6), .B1 (nx4276), .C0 (nx834)) ;
    dff reg_negative_M_6 (.Q (negative_M_6), .QB (\$dummy [28]), .D (nx818), .CLK (
        clk)) ;
    mux21_ni ix819 (.Y (nx818), .A0 (nx782), .A1 (negative_M_4), .S0 (nx4444)) ;
    dff reg_positive_M_6 (.Q (positive_M_6), .QB (nx3657), .D (nx802), .CLK (clk
        )) ;
    oai322 ix803 (.Y (nx802), .A0 (nx3652), .A1 (nx790), .A2 (nx4348), .B0 (
           nx3655), .B1 (nx4352), .C0 (nx4484), .C1 (nx3601)) ;
    nor02ii ix3653 (.Y (nx3652), .A0 (nx696), .A1 (nx4771)) ;
    inv01 ix3656 (.Y (nx3655), .A (M[6])) ;
    dff reg_product_7 (.Q (product[7]), .QB (\$dummy [29]), .D (aux_product_7), 
        .CLK (clk)) ;
    oai21 ix3169 (.Y (nx3168), .A0 (nx3663), .A1 (nx4292), .B0 (nx3665)) ;
    dff reg_aux_product_7 (.Q (aux_product_7), .QB (nx3663), .D (nx3168), .CLK (
        clk)) ;
    nand03 ix3666 (.Y (nx3665), .A0 (nx4444), .A1 (nx934), .A2 (nx4292)) ;
    xnor2 ix935 (.Y (nx934), .A0 (nx3668), .A1 (nx932)) ;
    dff reg_negative_M_7 (.Q (negative_M_7), .QB (\$dummy [30]), .D (nx912), .CLK (
        clk)) ;
    mux21_ni ix913 (.Y (nx912), .A0 (nx4580), .A1 (negative_M_5), .S0 (nx4444)
             ) ;
    dff reg_positive_M_7 (.Q (positive_M_7), .QB (nx3685), .D (nx896), .CLK (clk
        )) ;
    oai322 ix897 (.Y (nx896), .A0 (nx3680), .A1 (nx884), .A2 (nx4348), .B0 (
           nx3683), .B1 (nx4352), .C0 (nx4310), .C1 (nx3629)) ;
    nor02ii ix3681 (.Y (nx3680), .A0 (nx790), .A1 (nx4580)) ;
    inv01 ix3684 (.Y (nx3683), .A (M[7])) ;
    dff reg_product_8 (.Q (product[8]), .QB (\$dummy [31]), .D (aux_product_8), 
        .CLK (clk)) ;
    oai21 ix3179 (.Y (nx3178), .A0 (nx3691), .A1 (nx4292), .B0 (nx3693)) ;
    dff reg_aux_product_8 (.Q (aux_product_8), .QB (nx3691), .D (nx3178), .CLK (
        clk)) ;
    nand03 ix3694 (.Y (nx3693), .A0 (nx4444), .A1 (nx1028), .A2 (nx4292)) ;
    xnor2 ix1029 (.Y (nx1028), .A0 (nx5921), .A1 (nx1026)) ;
    dff reg_negative_M_8 (.Q (negative_M_8), .QB (\$dummy [32]), .D (nx1006), .CLK (
        clk)) ;
    mux21_ni ix1007 (.Y (nx1006), .A0 (nx970), .A1 (negative_M_6), .S0 (nx4446)
             ) ;
    dff reg_positive_M_8 (.Q (positive_M_8), .QB (nx3713), .D (nx990), .CLK (clk
        )) ;
    oai322 ix991 (.Y (nx990), .A0 (nx3708), .A1 (nx978), .A2 (nx4348), .B0 (
           nx3711), .B1 (nx4352), .C0 (nx4310), .C1 (nx3657)) ;
    nor02ii ix3709 (.Y (nx3708), .A0 (nx884), .A1 (nx970)) ;
    inv01 ix3712 (.Y (nx3711), .A (M[8])) ;
    dff reg_product_9 (.Q (product[9]), .QB (\$dummy [33]), .D (aux_product_9), 
        .CLK (clk)) ;
    oai21 ix3189 (.Y (nx3188), .A0 (nx3719), .A1 (nx4292), .B0 (nx3721)) ;
    dff reg_aux_product_9 (.Q (aux_product_9), .QB (nx3719), .D (nx3188), .CLK (
        clk)) ;
    nand03 ix3722 (.Y (nx3721), .A0 (nx4446), .A1 (nx1122), .A2 (nx4292)) ;
    xnor2 ix1123 (.Y (nx1122), .A0 (nx3724), .A1 (nx1120)) ;
    dff reg_negative_M_9 (.Q (negative_M_9), .QB (\$dummy [34]), .D (nx1100), .CLK (
        clk)) ;
    mux21_ni ix1101 (.Y (nx1100), .A0 (nx1064), .A1 (negative_M_7), .S0 (nx4446)
             ) ;
    dff reg_positive_M_9 (.Q (positive_M_9), .QB (nx3741), .D (nx1084), .CLK (
        clk)) ;
    oai322 ix1085 (.Y (nx1084), .A0 (nx3736), .A1 (nx1072), .A2 (nx4348), .B0 (
           nx3739), .B1 (nx4352), .C0 (nx4310), .C1 (nx3685)) ;
    nor02ii ix3737 (.Y (nx3736), .A0 (nx4849), .A1 (nx1064)) ;
    inv01 ix3740 (.Y (nx3739), .A (M[9])) ;
    dff reg_product_10 (.Q (product[10]), .QB (\$dummy [35]), .D (aux_product_10
        ), .CLK (clk)) ;
    oai21 ix3199 (.Y (nx3198), .A0 (nx3747), .A1 (nx4292), .B0 (nx3749)) ;
    dff reg_aux_product_10 (.Q (aux_product_10), .QB (nx3747), .D (nx3198), .CLK (
        clk)) ;
    nand03 ix3750 (.Y (nx3749), .A0 (nx4446), .A1 (nx1216), .A2 (nx4294)) ;
    xnor2 ix1217 (.Y (nx1216), .A0 (nx3752), .A1 (nx1214)) ;
    dff reg_negative_M_10 (.Q (negative_M_10), .QB (\$dummy [36]), .D (nx1194), 
        .CLK (clk)) ;
    mux21_ni ix1195 (.Y (nx1194), .A0 (nx1158), .A1 (negative_M_8), .S0 (nx4446)
             ) ;
    dff reg_positive_M_10 (.Q (positive_M_10), .QB (nx3769), .D (nx1178), .CLK (
        clk)) ;
    oai322 ix1179 (.Y (nx1178), .A0 (nx3764), .A1 (nx1166), .A2 (nx4348), .B0 (
           nx3767), .B1 (nx4352), .C0 (nx4310), .C1 (nx3713)) ;
    nor02ii ix3765 (.Y (nx3764), .A0 (nx4847), .A1 (nx4842)) ;
    inv01 ix3768 (.Y (nx3767), .A (M[10])) ;
    dff reg_product_11 (.Q (product[11]), .QB (\$dummy [37]), .D (aux_product_11
        ), .CLK (clk)) ;
    oai21 ix3209 (.Y (nx3208), .A0 (nx3775), .A1 (nx4294), .B0 (nx3777)) ;
    dff reg_aux_product_11 (.Q (aux_product_11), .QB (nx3775), .D (nx3208), .CLK (
        clk)) ;
    nand03 ix3778 (.Y (nx3777), .A0 (nx4446), .A1 (nx1310), .A2 (nx4294)) ;
    xnor2 ix1311 (.Y (nx1310), .A0 (nx3780), .A1 (nx5905)) ;
    dff reg_negative_M_11 (.Q (negative_M_11), .QB (\$dummy [38]), .D (nx1288), 
        .CLK (clk)) ;
    mux21_ni ix1289 (.Y (nx1288), .A0 (nx1252), .A1 (negative_M_9), .S0 (nx4446)
             ) ;
    nor02ii ix1151 (.Y (nx1150), .A0 (M[10]), .A1 (nx1056)) ;
    dff reg_positive_M_11 (.Q (positive_M_11), .QB (nx3797), .D (nx1272), .CLK (
        clk)) ;
    oai322 ix1273 (.Y (nx1272), .A0 (nx3792), .A1 (nx1260), .A2 (nx4350), .B0 (
           nx3795), .B1 (nx4354), .C0 (nx4310), .C1 (nx3741)) ;
    nor02ii ix3793 (.Y (nx3792), .A0 (nx4839), .A1 (nx1252)) ;
    inv01 ix3796 (.Y (nx3795), .A (M[11])) ;
    dff reg_product_12 (.Q (product[12]), .QB (\$dummy [39]), .D (aux_product_12
        ), .CLK (clk)) ;
    oai21 ix3219 (.Y (nx3218), .A0 (nx3803), .A1 (nx4294), .B0 (nx3805)) ;
    dff reg_aux_product_12 (.Q (aux_product_12), .QB (nx3803), .D (nx3218), .CLK (
        clk)) ;
    nand03 ix3806 (.Y (nx3805), .A0 (nx4448), .A1 (nx1404), .A2 (nx4294)) ;
    xnor2 ix1405 (.Y (nx1404), .A0 (nx3808), .A1 (nx1402)) ;
    dff reg_negative_M_12 (.Q (negative_M_12), .QB (\$dummy [40]), .D (nx1382), 
        .CLK (clk)) ;
    mux21_ni ix1383 (.Y (nx1382), .A0 (nx1346), .A1 (negative_M_10), .S0 (nx4448
             )) ;
    dff reg_positive_M_12 (.Q (positive_M_12), .QB (nx3825), .D (nx1366), .CLK (
        clk)) ;
    oai322 ix1367 (.Y (nx1366), .A0 (nx3820), .A1 (nx1354), .A2 (nx4350), .B0 (
           nx3823), .B1 (nx4354), .C0 (nx4310), .C1 (nx3769)) ;
    nor02ii ix3821 (.Y (nx3820), .A0 (nx1260), .A1 (nx1346)) ;
    inv01 ix3824 (.Y (nx3823), .A (M[12])) ;
    dff reg_product_13 (.Q (product[13]), .QB (\$dummy [41]), .D (aux_product_13
        ), .CLK (clk)) ;
    oai21 ix3229 (.Y (nx3228), .A0 (nx3831), .A1 (nx4294), .B0 (nx3833)) ;
    dff reg_aux_product_13 (.Q (aux_product_13), .QB (nx3831), .D (nx3228), .CLK (
        clk)) ;
    nand03 ix3834 (.Y (nx3833), .A0 (nx4448), .A1 (nx1498), .A2 (nx4294)) ;
    xnor2 ix1499 (.Y (nx1498), .A0 (nx3836), .A1 (nx1496)) ;
    dff reg_negative_M_13 (.Q (negative_M_13), .QB (\$dummy [42]), .D (nx1476), 
        .CLK (clk)) ;
    mux21_ni ix1477 (.Y (nx1476), .A0 (nx1440), .A1 (negative_M_11), .S0 (nx4448
             )) ;
    dff reg_positive_M_13 (.Q (positive_M_13), .QB (nx3853), .D (nx1460), .CLK (
        clk)) ;
    oai322 ix1461 (.Y (nx1460), .A0 (nx3848), .A1 (nx1448), .A2 (nx4350), .B0 (
           nx3851), .B1 (nx4354), .C0 (nx4310), .C1 (nx3797)) ;
    nor02ii ix3849 (.Y (nx3848), .A0 (nx1354), .A1 (nx4873)) ;
    inv01 ix3852 (.Y (nx3851), .A (M[13])) ;
    dff reg_product_14 (.Q (product[14]), .QB (\$dummy [43]), .D (aux_product_14
        ), .CLK (clk)) ;
    oai21 ix3239 (.Y (nx3238), .A0 (nx3859), .A1 (nx4296), .B0 (nx3861)) ;
    dff reg_aux_product_14 (.Q (aux_product_14), .QB (nx3859), .D (nx3238), .CLK (
        clk)) ;
    nand03 ix3862 (.Y (nx3861), .A0 (nx4448), .A1 (nx1592), .A2 (nx4296)) ;
    xnor2 ix1593 (.Y (nx1592), .A0 (nx3864), .A1 (nx1590)) ;
    dff reg_negative_M_14 (.Q (negative_M_14), .QB (nx3873), .D (nx1570), .CLK (
        clk)) ;
    mux21_ni ix1571 (.Y (nx1570), .A0 (nx1534), .A1 (negative_M_12), .S0 (nx4448
             )) ;
    dff reg_positive_M_14 (.Q (positive_M_14), .QB (\$dummy [44]), .D (nx1554), 
        .CLK (clk)) ;
    oai322 ix1555 (.Y (nx1554), .A0 (nx3876), .A1 (nx1542), .A2 (nx4350), .B0 (
           nx3879), .B1 (nx4354), .C0 (nx4312), .C1 (nx3825)) ;
    nor02ii ix3877 (.Y (nx3876), .A0 (nx1448), .A1 (nx4868)) ;
    inv01 ix3880 (.Y (nx3879), .A (M[14])) ;
    dff reg_product_15 (.Q (product[15]), .QB (\$dummy [45]), .D (aux_product_15
        ), .CLK (clk)) ;
    oai21 ix3249 (.Y (nx3248), .A0 (nx3887), .A1 (nx4296), .B0 (nx3889)) ;
    dff reg_aux_product_15 (.Q (aux_product_15), .QB (nx3887), .D (nx3248), .CLK (
        clk)) ;
    nand03 ix3890 (.Y (nx3889), .A0 (nx4448), .A1 (nx1662), .A2 (nx4296)) ;
    xnor2 ix1663 (.Y (nx1662), .A0 (nx3892), .A1 (nx1660)) ;
    aoi221 ix3896 (.Y (nx3895), .A0 (negative_M_15), .A1 (nx4268), .B0 (
           positive_M_15), .B1 (nx4280), .C0 (nx1656)) ;
    dff reg_negative_M_15 (.Q (negative_M_15), .QB (nx3901), .D (nx1640), .CLK (
        clk)) ;
    mux21_ni ix1641 (.Y (nx1640), .A0 (nx1616), .A1 (negative_M_13), .S0 (nx4450
             )) ;
    xnor2 ix1617 (.Y (nx1616), .A0 (M[15]), .A1 (nx1526)) ;
    nor02ii ix1527 (.Y (nx1526), .A0 (M[14]), .A1 (nx1432)) ;
    dff reg_positive_M_15 (.Q (positive_M_15), .QB (\$dummy [46]), .D (nx1624), 
        .CLK (clk)) ;
    oai22 ix1625 (.Y (nx1624), .A0 (nx3904), .A1 (nx4350), .B0 (nx4312), .B1 (
          nx3853)) ;
    xor2 ix3905 (.Y (nx3904), .A0 (nx1616), .A1 (nx1542)) ;
    dff reg_product_16 (.Q (product[16]), .QB (\$dummy [47]), .D (aux_product_16
        ), .CLK (clk)) ;
    oai21 ix3259 (.Y (nx3258), .A0 (nx3912), .A1 (nx4296), .B0 (nx3914)) ;
    dff reg_aux_product_16 (.Q (aux_product_16), .QB (nx3912), .D (nx3258), .CLK (
        clk)) ;
    nand03 ix3915 (.Y (nx3914), .A0 (nx4450), .A1 (nx1732), .A2 (nx4296)) ;
    xnor2 ix1733 (.Y (nx1732), .A0 (nx3917), .A1 (nx1730)) ;
    aoi221 ix3921 (.Y (nx3920), .A0 (negative_M_16), .A1 (nx4268), .B0 (
           positive_M_16), .B1 (nx4280), .C0 (nx1726)) ;
    dff reg_negative_M_16 (.Q (negative_M_16), .QB (nx3928), .D (nx1710), .CLK (
        clk)) ;
    oai21 ix1711 (.Y (nx1710), .A0 (nx4312), .A1 (nx3873), .B0 (nx4380)) ;
    nand02 ix3925 (.Y (nx3924), .A0 (nx3926), .A1 (nx350)) ;
    dff reg_positive_M_16 (.Q (positive_M_16), .QB (\$dummy [48]), .D (nx1694), 
        .CLK (clk)) ;
    oai21 ix3932 (.Y (nx3931), .A0 (nx3933), .A1 (nx1616), .B0 (nx4482)) ;
    dff reg_product_17 (.Q (product[17]), .QB (\$dummy [49]), .D (aux_product_17
        ), .CLK (clk)) ;
    oai21 ix3269 (.Y (nx3268), .A0 (nx3943), .A1 (nx4296), .B0 (nx3945)) ;
    dff reg_aux_product_17 (.Q (aux_product_17), .QB (nx3943), .D (nx3268), .CLK (
        clk)) ;
    nand03 ix3946 (.Y (nx3945), .A0 (nx4450), .A1 (nx1792), .A2 (nx4298)) ;
    xnor2 ix1793 (.Y (nx1792), .A0 (nx3948), .A1 (nx1790)) ;
    dff reg_negative_M_17 (.Q (negative_M_17), .QB (nx3955), .D (nx1770), .CLK (
        clk)) ;
    oai21 ix1771 (.Y (nx1770), .A0 (nx4312), .A1 (nx3901), .B0 (nx4380)) ;
    dff reg_positive_M_17 (.Q (positive_M_17), .QB (\$dummy [50]), .D (nx1758), 
        .CLK (clk)) ;
    dff reg_product_18 (.Q (product[18]), .QB (\$dummy [51]), .D (aux_product_18
        ), .CLK (clk)) ;
    oai21 ix3279 (.Y (nx3278), .A0 (nx3964), .A1 (nx4298), .B0 (nx3966)) ;
    dff reg_aux_product_18 (.Q (aux_product_18), .QB (nx3964), .D (nx3278), .CLK (
        clk)) ;
    nand03 ix3967 (.Y (nx3966), .A0 (nx4450), .A1 (nx1852), .A2 (nx4298)) ;
    xnor2 ix1853 (.Y (nx1852), .A0 (nx3969), .A1 (nx5220)) ;
    dff reg_negative_M_18 (.Q (negative_M_18), .QB (nx3976), .D (nx1830), .CLK (
        clk)) ;
    oai21 ix1831 (.Y (nx1830), .A0 (nx4312), .A1 (nx3928), .B0 (nx4380)) ;
    dff reg_positive_M_18 (.Q (positive_M_18), .QB (\$dummy [52]), .D (nx1818), 
        .CLK (clk)) ;
    dff reg_product_19 (.Q (product[19]), .QB (\$dummy [53]), .D (aux_product_19
        ), .CLK (clk)) ;
    oai21 ix3289 (.Y (nx3288), .A0 (nx3985), .A1 (nx4298), .B0 (nx3987)) ;
    dff reg_aux_product_19 (.Q (aux_product_19), .QB (nx3985), .D (nx3288), .CLK (
        clk)) ;
    nand03 ix3988 (.Y (nx3987), .A0 (nx4450), .A1 (nx1912), .A2 (nx4298)) ;
    xnor2 ix1913 (.Y (nx1912), .A0 (nx3990), .A1 (nx1910)) ;
    aoi221 ix3994 (.Y (nx3993), .A0 (negative_M_19), .A1 (nx4268), .B0 (
           positive_M_19), .B1 (nx4280), .C0 (nx1906)) ;
    dff reg_negative_M_19 (.Q (negative_M_19), .QB (nx3997), .D (nx1890), .CLK (
        clk)) ;
    oai21 ix1891 (.Y (nx1890), .A0 (nx4314), .A1 (nx3955), .B0 (nx4380)) ;
    dff reg_positive_M_19 (.Q (positive_M_19), .QB (\$dummy [54]), .D (nx1878), 
        .CLK (clk)) ;
    dff reg_product_20 (.Q (product[20]), .QB (\$dummy [55]), .D (aux_product_20
        ), .CLK (clk)) ;
    oai21 ix3299 (.Y (nx3298), .A0 (nx4006), .A1 (nx4298), .B0 (nx4008)) ;
    dff reg_aux_product_20 (.Q (aux_product_20), .QB (nx4006), .D (nx3298), .CLK (
        clk)) ;
    nand03 ix4009 (.Y (nx4008), .A0 (nx4450), .A1 (nx1972), .A2 (nx4298)) ;
    xnor2 ix1973 (.Y (nx1972), .A0 (nx4011), .A1 (nx1970)) ;
    aoi221 ix4015 (.Y (nx4014), .A0 (negative_M_20), .A1 (nx4268), .B0 (
           positive_M_20), .B1 (nx4280), .C0 (nx1966)) ;
    dff reg_negative_M_20 (.Q (negative_M_20), .QB (nx4018), .D (nx1950), .CLK (
        clk)) ;
    oai21 ix1951 (.Y (nx1950), .A0 (nx4314), .A1 (nx3976), .B0 (nx4380)) ;
    dff reg_positive_M_20 (.Q (positive_M_20), .QB (\$dummy [56]), .D (nx1938), 
        .CLK (clk)) ;
    dff reg_product_21 (.Q (product[21]), .QB (\$dummy [57]), .D (aux_product_21
        ), .CLK (clk)) ;
    oai21 ix3309 (.Y (nx3308), .A0 (nx4027), .A1 (nx5228), .B0 (nx4029)) ;
    dff reg_aux_product_21 (.Q (aux_product_21), .QB (nx4027), .D (nx3308), .CLK (
        clk)) ;
    nand03 ix4030 (.Y (nx4029), .A0 (nx4450), .A1 (nx2032), .A2 (nx5228)) ;
    xnor2 ix2033 (.Y (nx2032), .A0 (nx4032), .A1 (nx2030)) ;
    aoi221 ix4036 (.Y (nx4035), .A0 (negative_M_21), .A1 (nx4268), .B0 (
           positive_M_21), .B1 (nx4280), .C0 (nx2026)) ;
    dff reg_negative_M_21 (.Q (negative_M_21), .QB (nx4039), .D (nx2010), .CLK (
        clk)) ;
    oai21 ix2011 (.Y (nx2010), .A0 (nx4314), .A1 (nx3997), .B0 (nx4380)) ;
    dff reg_positive_M_21 (.Q (positive_M_21), .QB (\$dummy [58]), .D (nx1998), 
        .CLK (clk)) ;
    dff reg_product_22 (.Q (product[22]), .QB (\$dummy [59]), .D (aux_product_22
        ), .CLK (clk)) ;
    oai21 ix3319 (.Y (nx3318), .A0 (nx4048), .A1 (nx5228), .B0 (nx4050)) ;
    dff reg_aux_product_22 (.Q (aux_product_22), .QB (nx4048), .D (nx3318), .CLK (
        clk)) ;
    nand03 ix4051 (.Y (nx4050), .A0 (nx4452), .A1 (nx2092), .A2 (nx5228)) ;
    xnor2 ix2093 (.Y (nx2092), .A0 (nx4053), .A1 (nx5234)) ;
    dff reg_negative_M_22 (.Q (negative_M_22), .QB (nx4060), .D (nx2070), .CLK (
        clk)) ;
    oai21 ix2071 (.Y (nx2070), .A0 (nx4316), .A1 (nx4018), .B0 (nx4380)) ;
    dff reg_positive_M_22 (.Q (positive_M_22), .QB (\$dummy [60]), .D (nx2058), 
        .CLK (clk)) ;
    dff reg_product_23 (.Q (product[23]), .QB (\$dummy [61]), .D (aux_product_23
        ), .CLK (clk)) ;
    dff reg_aux_product_23 (.Q (aux_product_23), .QB (nx4069), .D (nx3328), .CLK (
        clk)) ;
    dff reg_negative_M_23 (.Q (negative_M_23), .QB (nx4081), .D (nx2130), .CLK (
        clk)) ;
    oai21 ix2131 (.Y (nx2130), .A0 (nx4316), .A1 (nx4039), .B0 (nx4382)) ;
    dff reg_positive_M_23 (.Q (positive_M_23), .QB (\$dummy [62]), .D (nx2118), 
        .CLK (clk)) ;
    dff reg_product_24 (.Q (product[24]), .QB (\$dummy [63]), .D (aux_product_24
        ), .CLK (clk)) ;
    dff reg_aux_product_24 (.Q (aux_product_24), .QB (nx4090), .D (nx3338), .CLK (
        clk)) ;
    aoi221 ix4099 (.Y (nx4098), .A0 (negative_M_24), .A1 (nx4270), .B0 (
           positive_M_24), .B1 (nx4282), .C0 (nx2206)) ;
    dff reg_negative_M_24 (.Q (negative_M_24), .QB (nx4102), .D (nx2190), .CLK (
        clk)) ;
    oai21 ix2191 (.Y (nx2190), .A0 (nx4316), .A1 (nx4060), .B0 (nx4382)) ;
    dff reg_positive_M_24 (.Q (positive_M_24), .QB (\$dummy [64]), .D (nx2178), 
        .CLK (clk)) ;
    dff reg_product_25 (.Q (product[25]), .QB (\$dummy [65]), .D (aux_product_25
        ), .CLK (clk)) ;
    oai21 ix3349 (.Y (nx3348), .A0 (nx4111), .A1 (nx5228), .B0 (nx4113)) ;
    dff reg_aux_product_25 (.Q (aux_product_25), .QB (nx4111), .D (nx3348), .CLK (
        clk)) ;
    nand03 ix4114 (.Y (nx4113), .A0 (nx4452), .A1 (nx2272), .A2 (nx5228)) ;
    xnor2 ix2273 (.Y (nx2272), .A0 (nx4116), .A1 (nx2270)) ;
    dff reg_negative_M_25 (.Q (negative_M_25), .QB (nx4123), .D (nx2250), .CLK (
        clk)) ;
    oai21 ix2251 (.Y (nx2250), .A0 (nx4316), .A1 (nx4081), .B0 (nx4382)) ;
    dff reg_positive_M_25 (.Q (positive_M_25), .QB (\$dummy [66]), .D (nx2238), 
        .CLK (clk)) ;
    dff reg_product_26 (.Q (product[26]), .QB (\$dummy [67]), .D (aux_product_26
        ), .CLK (clk)) ;
    dff reg_aux_product_26 (.Q (aux_product_26), .QB (nx4132), .D (nx3358), .CLK (
        clk)) ;
    dff reg_negative_M_26 (.Q (negative_M_26), .QB (nx4144), .D (nx2310), .CLK (
        clk)) ;
    oai21 ix2311 (.Y (nx2310), .A0 (nx4318), .A1 (nx4102), .B0 (nx4382)) ;
    dff reg_positive_M_26 (.Q (positive_M_26), .QB (\$dummy [68]), .D (nx2298), 
        .CLK (clk)) ;
    dff reg_product_27 (.Q (product[27]), .QB (\$dummy [69]), .D (aux_product_27
        ), .CLK (clk)) ;
    oai21 ix3369 (.Y (nx3368), .A0 (nx4153), .A1 (nx5228), .B0 (nx4155)) ;
    dff reg_aux_product_27 (.Q (aux_product_27), .QB (nx4153), .D (nx3368), .CLK (
        clk)) ;
    aoi221 ix4162 (.Y (nx4161), .A0 (negative_M_27), .A1 (nx4270), .B0 (
           positive_M_27), .B1 (nx4282), .C0 (nx2386)) ;
    dff reg_negative_M_27 (.Q (negative_M_27), .QB (nx4165), .D (nx2370), .CLK (
        clk)) ;
    oai21 ix2371 (.Y (nx2370), .A0 (nx4318), .A1 (nx4123), .B0 (nx4382)) ;
    dff reg_positive_M_27 (.Q (positive_M_27), .QB (\$dummy [70]), .D (nx2358), 
        .CLK (clk)) ;
    dff reg_product_28 (.Q (product[28]), .QB (\$dummy [71]), .D (aux_product_28
        ), .CLK (clk)) ;
    dff reg_aux_product_28 (.Q (aux_product_28), .QB (nx4174), .D (nx3378), .CLK (
        clk)) ;
    aoi221 ix4183 (.Y (nx4182), .A0 (negative_M_28), .A1 (nx4270), .B0 (
           positive_M_28), .B1 (nx4282), .C0 (nx2446)) ;
    dff reg_negative_M_28 (.Q (negative_M_28), .QB (nx4186), .D (nx2430), .CLK (
        clk)) ;
    oai21 ix2431 (.Y (nx2430), .A0 (nx4318), .A1 (nx4144), .B0 (nx4382)) ;
    dff reg_positive_M_28 (.Q (positive_M_28), .QB (\$dummy [72]), .D (nx2418), 
        .CLK (clk)) ;
    dff reg_product_29 (.Q (product[29]), .QB (\$dummy [73]), .D (aux_product_29
        ), .CLK (clk)) ;
    dff reg_aux_product_29 (.Q (aux_product_29), .QB (nx4195), .D (nx3388), .CLK (
        clk)) ;
    aoi221 ix4204 (.Y (nx4203), .A0 (negative_M_29), .A1 (nx4272), .B0 (
           positive_M_29), .B1 (nx4284), .C0 (nx2506)) ;
    dff reg_negative_M_29 (.Q (negative_M_29), .QB (nx4207), .D (nx2490), .CLK (
        clk)) ;
    oai21 ix2491 (.Y (nx2490), .A0 (nx4320), .A1 (nx4165), .B0 (nx4382)) ;
    dff reg_positive_M_29 (.Q (positive_M_29), .QB (\$dummy [74]), .D (nx2478), 
        .CLK (clk)) ;
    dff reg_product_30 (.Q (product[30]), .QB (\$dummy [75]), .D (aux_product_30
        ), .CLK (clk)) ;
    oai21 ix3399 (.Y (nx3398), .A0 (nx4216), .A1 (nx4304), .B0 (nx4218)) ;
    dff reg_aux_product_30 (.Q (aux_product_30), .QB (nx4216), .D (nx3398), .CLK (
        clk)) ;
    aoi221 ix4225 (.Y (nx4224), .A0 (negative_2M_31), .A1 (nx4272), .B0 (
           positive_2M_31), .B1 (nx4284), .C0 (nx2566)) ;
    dff reg_negative_2M_31 (.Q (negative_2M_31), .QB (\$dummy [76]), .D (nx2550)
        , .CLK (clk)) ;
    oai21 ix2551 (.Y (nx2550), .A0 (nx4320), .A1 (nx4186), .B0 (nx3924)) ;
    dff reg_positive_2M_31 (.Q (positive_2M_31), .QB (\$dummy [77]), .D (nx2538)
        , .CLK (clk)) ;
    dff reg_product_31 (.Q (product[31]), .QB (\$dummy [78]), .D (aux_product_31
        ), .CLK (clk)) ;
    dff reg_aux_product_31 (.Q (aux_product_31), .QB (nx4237), .D (nx3408), .CLK (
        clk)) ;
    aoi221 ix4246 (.Y (nx4245), .A0 (negative_M_31), .A1 (nx4272), .B0 (
           positive_M_31), .B1 (nx4284), .C0 (nx2626)) ;
    dff reg_negative_M_31 (.Q (negative_M_31), .QB (\$dummy [79]), .D (nx2610), 
        .CLK (clk)) ;
    oai21 ix2611 (.Y (nx2610), .A0 (nx4320), .A1 (nx4207), .B0 (nx3924)) ;
    dff reg_positive_M_31 (.Q (positive_M_31), .QB (\$dummy [80]), .D (nx2598), 
        .CLK (clk)) ;
    ao22 ix2627 (.Y (nx2626), .A0 (negative_2M_31), .A1 (nx4472), .B0 (
         positive_2M_31), .B1 (nx4462)) ;
    inv01 ix3934 (.Y (nx3933), .A (nx1542)) ;
    inv01 ix3927 (.Y (nx3926), .A (nx1526)) ;
    inv01 ix3535 (.Y (nx3534), .A (nx296)) ;
    inv02 ix4267 (.Y (nx4268), .A (nx4262)) ;
    inv02 ix4269 (.Y (nx4270), .A (nx4262)) ;
    inv02 ix4271 (.Y (nx4272), .A (nx4262)) ;
    inv02 ix4279 (.Y (nx4280), .A (nx4274)) ;
    inv02 ix4283 (.Y (nx4284), .A (nx4274)) ;
    inv01 ix4285 (.Y (nx4286), .A (nx254)) ;
    inv02 ix4287 (.Y (nx4288), .A (nx4420)) ;
    inv02 ix4289 (.Y (nx4290), .A (nx4420)) ;
    inv02 ix4291 (.Y (nx4292), .A (nx4420)) ;
    inv02 ix4293 (.Y (nx4294), .A (nx4420)) ;
    inv02 ix4295 (.Y (nx4296), .A (nx4420)) ;
    inv02 ix4297 (.Y (nx4298), .A (nx5226)) ;
    inv02 ix4307 (.Y (nx4308), .A (cnt_enable)) ;
    inv02 ix4309 (.Y (nx4310), .A (nx4454)) ;
    inv02 ix4311 (.Y (nx4312), .A (nx4454)) ;
    inv02 ix4313 (.Y (nx4314), .A (nx4454)) ;
    inv02 ix4315 (.Y (nx4316), .A (nx4454)) ;
    inv02 ix4317 (.Y (nx4318), .A (nx4456)) ;
    inv02 ix4319 (.Y (nx4320), .A (nx4456)) ;
    inv02 ix4331 (.Y (nx4332), .A (nx228)) ;
    inv04 ix4347 (.Y (nx4348), .A (nx338)) ;
    inv04 ix4349 (.Y (nx4350), .A (nx4482)) ;
    inv02 ix4351 (.Y (nx4352), .A (nx350)) ;
    inv02 ix4353 (.Y (nx4354), .A (nx350)) ;
    buf02 ix4375 (.Y (nx4376), .A (nx3895)) ;
    nand02 ix4379 (.Y (nx4380), .A0 (nx3926), .A1 (nx350)) ;
    nand02 ix4381 (.Y (nx4382), .A0 (nx3926), .A1 (nx350)) ;
    inv01 ix4383 (.Y (nx4384), .A (nx3931)) ;
    buf02 ix4395 (.Y (nx4396), .A (nx3993)) ;
    buf02 ix4397 (.Y (nx4398), .A (nx4014)) ;
    buf02 ix4399 (.Y (nx4400), .A (nx4035)) ;
    buf02 ix4401 (.Y (nx4402), .A (nx4056)) ;
    buf02 ix4405 (.Y (nx4406), .A (nx4098)) ;
    buf02 ix4409 (.Y (nx4410), .A (nx4140)) ;
    buf02 ix4411 (.Y (nx4412), .A (nx4161)) ;
    buf02 ix4413 (.Y (nx4414), .A (nx4182)) ;
    buf02 ix4415 (.Y (nx4416), .A (nx4203)) ;
    buf02 ix4417 (.Y (nx4418), .A (nx4224)) ;
    inv01 ix4419 (.Y (nx4420), .A (nx254)) ;
    and02 ix109 (.Y (nx108), .A0 (nx4456), .A1 (shifting_R_2)) ;
    and03 ix3482 (.Y (nx228), .A0 (shifting_R_0), .A1 (nx3454), .A2 (
          shifting_R_1)) ;
    nor02ii ix269 (.Y (nx268), .A0 (nx3424), .A1 (positive_2M_1)) ;
    nor02ii ix259 (.Y (nx258), .A0 (nx4456), .A1 (nx6007)) ;
    or02 ix247 (.Y (nx4262), .A0 (nx3454), .A1 (nx3424)) ;
    ao22 ix553 (.Y (nx552), .A0 (negative_M_2), .A1 (nx4472), .B0 (positive_M_2)
         , .B1 (nx4462)) ;
    nor02ii ix3596 (.Y (nx338), .A0 (nx4456), .A1 (M[15])) ;
    ao22 ix647 (.Y (nx646), .A0 (negative_M_3), .A1 (nx4472), .B0 (positive_M_3)
         , .B1 (nx4462)) ;
    ao22 ix741 (.Y (nx740), .A0 (negative_M_4), .A1 (nx4472), .B0 (positive_M_4)
         , .B1 (nx4462)) ;
    ao22 ix835 (.Y (nx834), .A0 (negative_M_5), .A1 (nx4472), .B0 (positive_M_5)
         , .B1 (nx4462)) ;
    xor2 ix1309 (.Y (nx1308), .A0 (nx3775), .A1 (nx5953)) ;
    xor2 ix1661 (.Y (nx1660), .A0 (nx3887), .A1 (nx4376)) ;
    ao22 ix1657 (.Y (nx1656), .A0 (negative_M_14), .A1 (nx4476), .B0 (
         positive_M_14), .B1 (nx4466)) ;
    ao21 ix1695 (.Y (nx1694), .A0 (nx4456), .A1 (positive_M_14), .B0 (nx4488)) ;
    ao22 ix1727 (.Y (nx1726), .A0 (negative_M_15), .A1 (nx4476), .B0 (
         positive_M_15), .B1 (nx4466)) ;
    ao21 ix1759 (.Y (nx1758), .A0 (nx4456), .A1 (positive_M_15), .B0 (nx4488)) ;
    ao21 ix1819 (.Y (nx1818), .A0 (nx4458), .A1 (positive_M_16), .B0 (nx4488)) ;
    ao21 ix1879 (.Y (nx1878), .A0 (nx4458), .A1 (positive_M_17), .B0 (nx4488)) ;
    ao22 ix1907 (.Y (nx1906), .A0 (negative_M_18), .A1 (nx4476), .B0 (
         positive_M_18), .B1 (nx4466)) ;
    ao21 ix1939 (.Y (nx1938), .A0 (nx4458), .A1 (positive_M_18), .B0 (nx4488)) ;
    ao22 ix1967 (.Y (nx1966), .A0 (negative_M_19), .A1 (nx4476), .B0 (
         positive_M_19), .B1 (nx4466)) ;
    ao21 ix1999 (.Y (nx1998), .A0 (nx4458), .A1 (positive_M_19), .B0 (nx4488)) ;
    ao22 ix2027 (.Y (nx2026), .A0 (negative_M_20), .A1 (nx4478_XX0_XREP64), .B0 (
         positive_M_20), .B1 (nx4468)) ;
    xor2 ix2091 (.Y (nx2090), .A0 (nx4048), .A1 (nx4402)) ;
    ao21 ix2059 (.Y (nx2058), .A0 (nx4458), .A1 (positive_M_20), .B0 (nx4488)) ;
    ao21 ix2119 (.Y (nx2118), .A0 (nx4458), .A1 (positive_M_21), .B0 (nx4490)) ;
    xor2_2x ix2211 (.Y (nx2210), .A0 (nx4090), .A1 (nx4406)) ;
    ao21 ix2179 (.Y (nx2178), .A0 (nx4458), .A1 (positive_M_22), .B0 (nx4490)) ;
    ao22 ix2207 (.Y (nx2206), .A0 (negative_M_23), .A1 (nx4478), .B0 (
         positive_M_23), .B1 (nx4468)) ;
    ao21 ix2239 (.Y (nx2238), .A0 (nx4460), .A1 (positive_M_23), .B0 (nx4490)) ;
    ao21 ix2299 (.Y (nx2298), .A0 (nx4460), .A1 (positive_M_24), .B0 (nx4490)) ;
    xor2 ix2391 (.Y (nx2390), .A0 (nx4153), .A1 (nx4412)) ;
    ao21 ix2359 (.Y (nx2358), .A0 (nx4460), .A1 (positive_M_25), .B0 (nx4490)) ;
    ao22 ix2387 (.Y (nx2386), .A0 (negative_M_26), .A1 (nx4478), .B0 (
         positive_M_26), .B1 (nx4468)) ;
    ao21 ix2419 (.Y (nx2418), .A0 (nx4460), .A1 (positive_M_26), .B0 (nx4490)) ;
    ao22 ix2447 (.Y (nx2446), .A0 (negative_M_27), .A1 (nx4480), .B0 (
         positive_M_27), .B1 (nx4470)) ;
    xor2 ix2511 (.Y (nx2510), .A0 (nx4195), .A1 (nx4416)) ;
    ao21 ix2479 (.Y (nx2478), .A0 (nx4460), .A1 (positive_M_27), .B0 (nx4490)) ;
    ao22 ix2507 (.Y (nx2506), .A0 (negative_M_28), .A1 (nx4480), .B0 (
         positive_M_28), .B1 (nx4470)) ;
    xor2 ix2571 (.Y (nx2570), .A0 (nx4216), .A1 (nx4418)) ;
    ao21 ix2539 (.Y (nx2538), .A0 (nx4460), .A1 (positive_M_28), .B0 (nx4384)) ;
    ao22 ix2567 (.Y (nx2566), .A0 (negative_M_29), .A1 (nx4480), .B0 (
         positive_M_29), .B1 (nx4470)) ;
    xor2 ix2631 (.Y (nx2630), .A0 (nx4237), .A1 (nx4245)) ;
    ao21 ix2599 (.Y (nx2598), .A0 (nx4460), .A1 (positive_M_29), .B0 (nx4384)) ;
    inv02 ix4435 (.Y (nx4436), .A (nx4484)) ;
    inv02 ix4437 (.Y (nx4438), .A (nx4484)) ;
    inv02 ix4439 (.Y (nx4440), .A (nx5232)) ;
    inv02 ix4441 (.Y (nx4442), .A (nx5232)) ;
    inv02 ix4443 (.Y (nx4444), .A (nx5232)) ;
    inv02 ix4445 (.Y (nx4446), .A (nx5232)) ;
    inv02 ix4447 (.Y (nx4448), .A (nx5232)) ;
    inv02 ix4449 (.Y (nx4450), .A (nx5233)) ;
    inv02 ix4455 (.Y (nx4456), .A (nx4308)) ;
    inv02 ix4457 (.Y (nx4458), .A (nx4308)) ;
    inv02 ix4459 (.Y (nx4460), .A (nx4308)) ;
    inv02 ix4465 (.Y (nx4466), .A (nx5208)) ;
    inv02 ix4467 (.Y (nx4468), .A (nx5208)) ;
    inv02 ix4469 (.Y (nx4470), .A (nx5208)) ;
    inv02 ix4475 (.Y (nx4476), .A (nx4322_XX0_XREP40)) ;
    inv02 ix4479 (.Y (nx4480), .A (nx4322)) ;
    inv02 ix4481 (.Y (nx4482), .A (nx4348)) ;
    inv02 ix4483 (.Y (nx4484), .A (cnt_enable)) ;
    inv02 ix4485 (.Y (nx4486), .A (cnt_enable)) ;
    inv01 ix4487 (.Y (nx4488), .A (nx3931)) ;
    inv01 ix4489 (.Y (nx4490), .A (nx3931)) ;
    nor03_2x ix237 (.Y (nx236), .A0 (shifting_R_0), .A1 (nx3454), .A2 (
             shifting_R_1)) ;
    inv02 ix4321_0_XREP40 (.Y (nx4322_XX0_XREP40), .A (nx236)) ;
    or02 ix251 (.Y (nx4274), .A0 (shifting_R_2), .A1 (nx3424)) ;
    dff reg_shifting_R_2 (.Q (shifting_R_2), .QB (nx3454), .D (nx100), .CLK (clk
        )) ;
    xnor2 ix3425 (.Y (nx3424), .A0 (shifting_R_1), .A1 (shifting_R_0)) ;
    or02 ix251_0_XREP44 (.Y (nx4274_XX0_XREP44), .A0 (shifting_R_2), .A1 (nx3424
         )) ;
    nor02ii ix885 (.Y (nx884), .A0 (nx4580), .A1 (nx790)) ;
    nor02ii ix791 (.Y (nx790), .A0 (nx4772), .A1 (nx696)) ;
    inv02 ix4321 (.Y (nx4322), .A (nx236)) ;
    inv02 ix4477_0_XREP64 (.Y (nx4478_XX0_XREP64), .A (nx4322)) ;
    buf04 ix5242 (.Y (nx4580), .A (nx876)) ;
    inv01 ix5243 (.Y (nx4581), .A (nx2510)) ;
    inv02 ix5244 (.Y (nx4582), .A (nx2570)) ;
    nor04_2x ix5245 (.Y (nx4583), .A0 (nx4582), .A1 (nx2630), .A2 (nx5226), .A3 (
             nx4308)) ;
    inv02 ix5246 (.Y (nx4584), .A (nx2630)) ;
    inv01 ix5247 (.Y (nx4585), .A (nx4418)) ;
    aoi22 ix5248 (.Y (nx4586), .A0 (nx2630), .A1 (nx4418), .B0 (nx4584), .B1 (
          nx4585)) ;
    nor02_2x ix5249 (.Y (nx4587), .A0 (nx5226), .A1 (nx4308)) ;
    nand03_2x ix5250 (.Y (nx4588), .A0 (nx4587), .A1 (nx2630), .A2 (nx2570)) ;
    inv02 ix5251 (.Y (nx4589), .A (nx2570)) ;
    and02 ix5252 (.Y (nx4590), .A0 (nx4416), .A1 (nx4581)) ;
    inv01 ix5253 (.Y (nx4591), .A (nx4414)) ;
    nand02_2x ix5254 (.Y (nx4592), .A0 (nx5152), .A1 (nx4591)) ;
    aoi22 ix5255 (.Y (nx4593), .A0 (nx4416), .A1 (nx4581), .B0 (nx2510), .B1 (
          nx4592)) ;
    nand02_2x ix5256 (.Y (nx4594), .A0 (nx4589), .A1 (nx4221)) ;
    nand04_2x reg_nx4218 (.Y (nx4218), .A0 (nx4594), .A1 (nx4614), .A2 (nx4454)
              , .A3 (nx4304)) ;
    inv01 ix5257 (.Y (nx4595), .A (nx5240)) ;
    nor03_2x ix5258 (.Y (nx4596), .A0 (nx4595), .A1 (nx4588), .A2 (nx4593)) ;
    nor02ii ix5259 (.Y (nx4597), .A0 (nx5240), .A1 (nx4412)) ;
    nor03_2x ix5260 (.Y (nx4598), .A0 (nx4597), .A1 (nx5152), .A2 (nx4590)) ;
    inv01 ix5261 (.Y (nx4599), .A (nx5226)) ;
    inv02 ix5262 (.Y (nx4600), .A (nx4308)) ;
    nand02_2x ix5263 (.Y (nx4601), .A0 (nx4599), .A1 (nx4600)) ;
    oai332 ix5264 (.Y (nx4602), .A0 (nx4598), .A1 (nx4588), .A2 (nx4593), .B0 (
           nx4586), .B1 (nx2570), .B2 (nx4601), .C0 (nx4304), .C1 (nx4237)) ;
    inv01 ix5265 (.Y (nx4603), .A (nx4593)) ;
    inv01 ix5266 (.Y (nx4604), .A (nx4598)) ;
    inv02 reg_nx4454 (.Y (nx4454), .A (nx4308)) ;
    nand03_2x ix5267 (.Y (nx4605), .A0 (nx2510), .A1 (nx4304), .A2 (nx4454)) ;
    inv02 ix5268 (.Y (nx4606), .A (nx2510)) ;
    nor02_2x ix5269 (.Y (nx4607), .A0 (nx5226), .A1 (nx4308)) ;
    and02 ix5270 (.Y (nx4608), .A0 (nx5240), .A1 (nx4603)) ;
    nand04_2x ix5271 (.Y (nx4609), .A0 (nx4116), .A1 (nx4608), .A2 (nx2330), .A3 (
              nx4885)) ;
    inv01 ix5272 (.Y (nx4610), .A (nx5236)) ;
    inv01 ix5273 (.Y (nx4611), .A (nx5238)) ;
    oai32 ix5274 (.Y (nx4612), .A0 (nx4886), .A1 (nx5959), .A2 (nx4610), .B0 (
          nx4611), .B1 (nx5178)) ;
    aoi321 ix5275 (.Y (nx4613), .A0 (nx4612), .A1 (nx5240), .A2 (nx4603), .B0 (
           nx4603), .B1 (nx4604), .C0 (nx4589)) ;
    nand02_2x ix5276 (.Y (nx4614), .A0 (nx4609), .A1 (nx4613)) ;
    inv01 ix5277 (.Y (nx4615), .A (nx4604)) ;
    oai321 ix5278 (.Y (nx4616), .A0 (nx5959), .A1 (nx4887), .A2 (nx5236), .B0 (
           nx5179), .B1 (nx5238), .C0 (nx5240)) ;
    inv01 ix5279 (.Y (nx4617), .A (nx4603)) ;
    inv01 ix5280 (.Y (nx4618), .A (nx2450)) ;
    inv01 ix5281 (.Y (nx4619), .A (nx4412)) ;
    inv01 ix5282 (.Y (nx4620), .A (nx4595)) ;
    inv02 reg_nx4304 (.Y (nx4304), .A (nx5227)) ;
    nand03_2x ix5283 (.Y (nx4621), .A0 (nx4618), .A1 (nx4304), .A2 (nx4452)) ;
    inv01 ix5284 (.Y (nx4622), .A (nx5236)) ;
    inv01 ix5285 (.Y (nx4623), .A (nx5238)) ;
    inv01 ix5286 (.Y (nx4624), .A (nx5234)) ;
    nor02ii ix5287 (.Y (nx4625), .A0 (nx5022), .A1 (nx5941)) ;
    inv01 ix5288 (.Y (nx4626), .A (nx2210)) ;
    aoi422 ix5289 (.Y (nx4627), .A0 (nx2210), .A1 (nx4624), .A2 (nx5023), .A3 (
           nx4402), .B0 (nx2210), .B1 (nx4625), .C0 (nx4406), .C1 (nx4626)) ;
    oai322 ix5290 (.Y (nx4628), .A0 (nx5129), .A1 (nx5143), .A2 (nx4622), .B0 (
           nx4623), .B1 (nx5139), .C0 (nx5174), .C1 (nx4627)) ;
    inv01 ix5291 (.Y (nx4629), .A (nx4402)) ;
    inv01 ix5292 (.Y (nx4630), .A (nx4077)) ;
    oai32 ix5293 (.Y (nx4631), .A0 (nx5029), .A1 (nx4629), .A2 (nx5234), .B0 (
          nx4630), .B1 (nx5024)) ;
    nor02_2x ix5294 (.Y (nx4632), .A0 (nx5959), .A1 (nx5236)) ;
    nor02_2x ix5295 (.Y (nx4633), .A0 (nx5959), .A1 (nx5052)) ;
    nor02_2x ix5296 (.Y (nx4634), .A0 (nx4629), .A1 (nx5234)) ;
    aoi22 ix5297 (.Y (nx4635), .A0 (nx5941), .A1 (nx5029), .B0 (nx5026), .B1 (
          nx4634)) ;
    ao22 reg_nx4074 (.Y (nx4074), .A0 (nx4402), .A1 (nx4624), .B0 (nx4053), .B1 (
         nx5235)) ;
    nor02_2x ix5298 (.Y (nx4636), .A0 (nx4632), .A1 (nx4633)) ;
    nor02_2x ix5299 (.Y (nx4637), .A0 (nx4619), .A1 (nx4620)) ;
    nand03_2x ix5300 (.Y (nx4638), .A0 (nx4905), .A1 (nx4907), .A2 (nx4909)) ;
    nand02_2x ix5301 (.Y (nx4639), .A0 (nx4904), .A1 (nx4638)) ;
    ao21 ix5302 (.Y (nx4640), .A0 (nx5027), .A1 (nx5235), .B0 (nx4631)) ;
    aoi22 ix5303 (.Y (nx4641), .A0 (nx2210), .A1 (nx4640), .B0 (nx4406), .B1 (
          nx4626)) ;
    and02 ix5304 (.Y (nx4642), .A0 (nx4406), .A1 (nx4626)) ;
    inv02 ix5305 (.Y (nx4643), .A (positive_M_1)) ;
    nor02_2x ix5306 (.Y (nx4644), .A0 (nx4643), .A1 (nx4274_XX0_XREP44)) ;
    inv02 ix5307 (.Y (nx4645), .A (negative_M_1)) ;
    nor02_2x ix5308 (.Y (nx4646), .A0 (nx4645), .A1 (nx4262)) ;
    nor04_2x ix5309 (.Y (nx4647), .A0 (nx4644), .A1 (nx4646), .A2 (nx4462), .A3 (
             nx4472)) ;
    inv01 ix5310 (.Y (nx4648), .A (positive_2M_1)) ;
    aoi22 ix5311 (.Y (nx4649), .A0 (nx4645), .A1 (nx4648), .B0 (nx4262), .B1 (
          nx4648)) ;
    nor02_2x ix5312 (.Y (nx4650), .A0 (nx4649), .A1 (nx4644)) ;
    inv01 ix5313 (.Y (nx4651), .A (nx3498)) ;
    and03 ix5314 (.Y (nx4652), .A0 (nx268), .A1 (aux_product_0), .A2 (nx4651)) ;
    and02 ix5315 (.Y (nx4653), .A0 (aux_product_0), .A1 (nx268)) ;
    inv02 reg_nx3526 (.Y (nx3526), .A (nx4690)) ;
    nand02_2x reg_nx3492 (.Y (nx3492), .A0 (aux_product_0), .A1 (nx268)) ;
    nor02_2x ix5316 (.Y (nx4654), .A0 (nx4711), .A1 (nx3498)) ;
    ao21 reg_nx368 (.Y (nx368), .A0 (nx3498), .A1 (nx4711), .B0 (nx4654)) ;
    and02 ix5317 (.Y (nx4655), .A0 (nx4931), .A1 (nx1970)) ;
    oai32 ix5318 (.Y (nx4656), .A0 (nx1970), .A1 (nx4922), .A2 (nx5224), .B0 (
          nx4932), .B1 (nx5230)) ;
    inv01 ix5319 (.Y (nx4657), .A (nx4641)) ;
    nand02_2x ix5320 (.Y (nx4658), .A0 (nx4639), .A1 (nx4657)) ;
    aoi322 reg_nx4158 (.Y (nx4158), .A0 (nx4683), .A1 (nx4898), .A2 (nx4655), .B0 (
           nx4656), .B1 (nx4898), .C0 (nx4658), .C1 (nx4895)) ;
    inv01 ix5321 (.Y (nx4659), .A (nx1970)) ;
    ao22 reg_nx4032 (.Y (nx4032), .A0 (nx5224), .A1 (nx4659), .B0 (nx4011), .B1 (
         nx1970)) ;
    aoi22 ix5322 (.Y (nx4660), .A0 (nx5236), .A1 (nx4880), .B0 (nx4888), .B1 (
          nx4116)) ;
    inv01 ix5323 (.Y (nx4661), .A (nx5236)) ;
    oai22 reg_nx4137 (.Y (nx4137), .A0 (nx4661), .A1 (nx5129), .B0 (nx4884), .B1 (
          nx5154)) ;
    nand03_2x ix5324 (.Y (nx4662), .A0 (nx5144), .A1 (nx5229), .A2 (nx4452)) ;
    oai422 reg_nx3358 (.Y (nx3358), .A0 (nx4660), .A1 (nx5145), .A2 (nx5227), .A3 (
           nx5233), .B0 (nx4137), .B1 (nx4662), .C0 (nx5229), .C1 (nx4132)) ;
    inv02 ix5325 (.Y (nx4663), .A (negative_M_1)) ;
    inv02 ix5326 (.Y (nx4664), .A (positive_M_1)) ;
    oai22 reg_nx458 (.Y (nx458), .A0 (nx4663), .A1 (nx4322_XX0_XREP40), .B0 (
          nx4664), .B1 (nx5208)) ;
    aoi221 reg_nx3529 (.Y (nx3529), .A0 (positive_M_2), .A1 (nx4276), .B0 (
           negative_M_2), .B1 (nx4264), .C0 (nx458)) ;
    inv02 ix5327 (.Y (nx4665), .A (nx3521)) ;
    inv01 reg_nx462 (.Y (nx462), .A (nx4692)) ;
    inv02 reg_nx4472 (.Y (nx4472), .A (nx4322_XX0_XREP40)) ;
    inv02 reg_nx4462 (.Y (nx4462), .A (nx5209)) ;
    nor02_2x ix5328 (.Y (nx4666), .A0 (nx4808), .A1 (nx4919)) ;
    and02 ix5329 (.Y (nx4667), .A0 (nx5220), .A1 (nx4790)) ;
    oai32 ix5330 (.Y (nx4668), .A0 (nx4791), .A1 (nx4786), .A2 (nx5200), .B0 (
          nx5220), .B1 (nx5931)) ;
    inv01 ix5331 (.Y (nx4669), .A (nx5222)) ;
    inv01 ix5332 (.Y (nx4670), .A (nx4655)) ;
    aoi21 ix5333 (.Y (nx4671), .A0 (nx4808), .A1 (nx4669), .B0 (nx4670)) ;
    nor02_2x ix5334 (.Y (nx4672), .A0 (nx4617), .A1 (nx4616)) ;
    oai21 ix5335 (.Y (nx4673), .A0 (nx5169), .A1 (nx4616), .B0 (nx4615)) ;
    inv01 ix5336 (.Y (nx4674), .A (nx4617)) ;
    nand03_2x ix5337 (.Y (nx4675), .A0 (nx4723), .A1 (nx5220), .A2 (nx4792)) ;
    nor02_2x ix5338 (.Y (nx4676), .A0 (nx3951), .A1 (nx4793)) ;
    aoi22 ix5339 (.Y (nx4677), .A0 (nx5931), .A1 (nx4787), .B0 (nx5221), .B1 (
          nx4676)) ;
    nand02_2x reg_nx3990 (.Y (nx3990), .A0 (nx4675), .A1 (nx4677)) ;
    ao22 reg_nx3969 (.Y (nx3969), .A0 (nx5200), .A1 (nx4804), .B0 (nx4724), .B1 (
         nx4794)) ;
    inv01 ix5340 (.Y (nx4678), .A (nx1660)) ;
    and02 ix5341 (.Y (nx4679), .A0 (nx5222), .A1 (nx4808)) ;
    nor02_2x ix5342 (.Y (nx4680), .A0 (nx4679), .A1 (nx4783)) ;
    inv01 ix5343 (.Y (nx4681), .A (nx5230)) ;
    nand02_2x ix5344 (.Y (nx4682), .A0 (nx4930), .A1 (nx4681)) ;
    inv01 ix5345 (.Y (nx4683), .A (nx4011)) ;
    ao22 reg_nx3917 (.Y (nx3917), .A0 (nx4376), .A1 (nx4678), .B0 (nx4709), .B1 (
         nx1660)) ;
    inv01 ix5346 (.Y (nx4684), .A (nx4653)) ;
    inv02 ix5347 (.Y (nx4685), .A (nx4651)) ;
    inv02 ix5348 (.Y (nx4686), .A (nx4665)) ;
    oai21 ix5349 (.Y (nx4687), .A0 (nx4653), .A1 (nx4651), .B0 (nx4665)) ;
    inv02 reg_nx3555 (.Y (nx3555), .A (nx4816)) ;
    nor02_2x ix5350 (.Y (nx4688), .A0 (nx4653), .A1 (nx4651)) ;
    nor02_2x ix5351 (.Y (nx4689), .A0 (nx4711), .A1 (nx4652)) ;
    nor02_2x ix5352 (.Y (nx4690), .A0 (nx4688), .A1 (nx4689)) ;
    inv01 ix5353 (.Y (nx4691), .A (nx3529)) ;
    oai22 ix5354 (.Y (nx4692), .A0 (nx4686), .A1 (nx5915), .B0 (nx4691), .B1 (
          nx4665)) ;
    inv01 ix5355 (.Y (nx4693), .A (nx1660)) ;
    nor03_2x ix5356 (.Y (nx4694), .A0 (nx4693), .A1 (nx5218), .A2 (nx4806)) ;
    inv01 ix5357 (.Y (nx4695), .A (nx3839)) ;
    inv01 ix5358 (.Y (nx4696), .A (nx3867)) ;
    oai32 ix5359 (.Y (nx4697), .A0 (nx5075), .A1 (nx5067), .A2 (nx4695), .B0 (
          nx4696), .B1 (nx5073)) ;
    nor02_2x ix5360 (.Y (nx4698), .A0 (nx5218), .A1 (nx5925)) ;
    inv01 ix5361 (.Y (nx4699), .A (nx3920)) ;
    oai21 ix5362 (.Y (nx4700), .A0 (nx4699), .A1 (nx5184), .B0 (nx4680)) ;
    aoi322 ix5363 (.Y (nx4701), .A0 (nx5074), .A1 (nx5951), .A2 (nx5071), .B0 (
           nx5949), .B1 (nx5067), .C0 (nx4944), .C1 (nx5072)) ;
    inv01 ix5364 (.Y (nx4702), .A (nx4678)) ;
    inv01 ix5365 (.Y (nx4703), .A (nx4376)) ;
    nor02_2x ix5366 (.Y (nx4704), .A0 (nx4376), .A1 (nx5911)) ;
    aoi33 ix5367 (.Y (nx4705), .A0 (nx5186), .A1 (nx4693), .A2 (nx4703), .B0 (
          nx5185), .B1 (nx4693), .B2 (nx4702)) ;
    aoi33 ix5368 (.Y (nx4706), .A0 (nx4693), .A1 (nx4703), .A2 (nx4699), .B0 (
          nx4702), .B1 (nx4693), .B2 (nx4699)) ;
    aoi22 ix5369 (.Y (nx4707), .A0 (nx5218), .A1 (nx4699), .B0 (nx5218), .B1 (
          nx5187)) ;
    nand03_2x ix5370 (.Y (nx4708), .A0 (nx4705), .A1 (nx4706), .A2 (nx4707)) ;
    inv01 reg_nx3892 (.Y (nx3892), .A (nx4701)) ;
    inv01 ix5371 (.Y (nx4709), .A (nx4701)) ;
    ao22 reg_nx3864 (.Y (nx3864), .A0 (nx5951), .A1 (nx5071), .B0 (nx3836), .B1 (
         nx5076)) ;
    aoi221 ix5372 (.Y (nx4710), .A0 (negative_M_3), .A1 (nx4264), .B0 (
           positive_M_3), .B1 (nx4276), .C0 (nx552)) ;
    nor02_2x ix5373 (.Y (nx4711), .A0 (nx4647), .A1 (nx4650)) ;
    inv01 ix5374 (.Y (nx4712), .A (nx4652)) ;
    aoi22 ix5375 (.Y (nx4713), .A0 (nx4686), .A1 (nx4712), .B0 (nx5915), .B1 (
          nx4712)) ;
    nor02_2x ix5376 (.Y (nx4714), .A0 (nx4711), .A1 (nx4713)) ;
    inv02 reg_nx3579 (.Y (nx3579), .A (nx4745)) ;
    inv02 ix5377 (.Y (nx4715), .A (nx3550)) ;
    nand02_2x ix5378 (.Y (nx4716), .A0 (nx4715), .A1 (nx5917)) ;
    oai21 reg_nx556 (.Y (nx556), .A0 (nx4715), .A1 (nx5917), .B0 (nx4716)) ;
    nand02_2x ix5379 (.Y (nx4717), .A0 (nx4673), .A1 (nx4674)) ;
    and02 ix5380 (.Y (nx4718), .A0 (nx4703), .A1 (nx5188)) ;
    oai22 ix5381 (.Y (nx4719), .A0 (nx4718), .A1 (nx4702), .B0 (nx4699), .B1 (
          nx5189)) ;
    nor02ii ix5382 (.Y (nx4720), .A0 (nx4704), .A1 (nx4719)) ;
    inv01 ix5383 (.Y (nx4721), .A (nx4708)) ;
    aoi22 ix5384 (.Y (nx4722), .A0 (nx4912), .A1 (nx4721), .B0 (nx4720), .B1 (
          nx4721)) ;
    inv01 reg_nx3948 (.Y (nx3948), .A (nx4722)) ;
    inv01 ix5385 (.Y (nx4723), .A (nx4722)) ;
    inv01 ix5386 (.Y (nx4724), .A (nx4722)) ;
    inv01 ix5387 (.Y (nx4725), .A (nx1308)) ;
    and02 ix5388 (.Y (nx4726), .A0 (nx5905), .A1 (nx4955)) ;
    aoi322 ix5389 (.Y (nx4727), .A0 (nx5905), .A1 (nx5935), .A2 (nx5214), .B0 (
           nx5953), .B1 (nx4725), .C0 (nx4748), .C1 (nx4726)) ;
    nand02_2x ix5390 (.Y (nx4728), .A0 (nx5072), .A1 (nx4996)) ;
    inv01 ix5391 (.Y (nx4729), .A (nx3811)) ;
    nor02_2x ix5392 (.Y (nx4730), .A0 (nx4729), .A1 (nx4997)) ;
    aoi21 ix5393 (.Y (nx4731), .A0 (nx5072), .A1 (nx4730), .B0 (nx4697)) ;
    nand02_2x ix5394 (.Y (nx4732), .A0 (nx5905), .A1 (nx4956)) ;
    inv01 ix5395 (.Y (nx4733), .A (nx3755)) ;
    inv01 ix5396 (.Y (nx4734), .A (nx3783)) ;
    aoi32 ix5397 (.Y (nx4735), .A0 (nx5905), .A1 (nx5214), .A2 (nx4733), .B0 (
          nx4725), .B1 (nx4734)) ;
    inv01 ix5398 (.Y (nx4736), .A (nx5072)) ;
    aoi21 ix5399 (.Y (nx4737), .A0 (nx4729), .A1 (nx5216), .B0 (nx4736)) ;
    inv01 ix5400 (.Y (nx4738), .A (nx4697)) ;
    and02 ix5401 (.Y (nx4739), .A0 (nx4998), .A1 (nx5905)) ;
    nor02_2x ix5402 (.Y (nx4740), .A0 (nx4733), .A1 (nx4957)) ;
    oai32 ix5403 (.Y (nx4741), .A0 (nx5905), .A1 (nx5216), .A2 (nx4734), .B0 (
          nx4729), .B1 (nx4999)) ;
    inv01 reg_nx3808 (.Y (nx3808), .A (nx4727)) ;
    ao22 reg_nx3780 (.Y (nx3780), .A0 (nx5935), .A1 (nx5214), .B0 (nx4749), .B1 (
         nx4958)) ;
    inv01 ix5404 (.Y (nx4742), .A (nx3582)) ;
    nor02_2x ix5405 (.Y (nx4743), .A0 (nx4816), .A1 (nx4814)) ;
    nor02_2x ix5406 (.Y (nx4744), .A0 (nx4743), .A1 (nx4831)) ;
    oai22 reg_nx3612 (.Y (nx3612), .A0 (nx4742), .A1 (nx650), .B0 (nx4826), .B1 (
          nx4744)) ;
    ao22 ix5407 (.Y (nx4745), .A0 (nx4816), .A1 (nx4830), .B0 (nx4814), .B1 (
         nx4830)) ;
    inv01 ix5408 (.Y (nx4746), .A (nx3643)) ;
    inv01 ix5409 (.Y (nx4747), .A (nx3671)) ;
    inv02 reg_nx3752 (.Y (nx3752), .A (nx5102)) ;
    inv01 ix5410 (.Y (nx4748), .A (nx5957)) ;
    inv01 ix5411 (.Y (nx4749), .A (nx5957)) ;
    nor02_2x ix5412 (.Y (nx4750), .A0 (nx4746), .A1 (nx4827)) ;
    aoi22 ix5413 (.Y (nx4751), .A0 (nx3671), .A1 (nx5057), .B0 (nx932), .B1 (
          nx4750)) ;
    oai422 reg_nx3724 (.Y (nx3724), .A0 (nx5945), .A1 (nx4822), .A2 (nx5058), .A3 (
           nx4825), .B0 (nx5012), .B1 (nx5009), .C0 (nx5945), .C1 (nx4751)) ;
    oai332 reg_nx3696 (.Y (nx3696), .A0 (nx5060), .A1 (nx4825), .A2 (nx4823), .B0 (
           nx5059), .B1 (nx4746), .B2 (nx4828), .C0 (nx4747), .C1 (nx932)) ;
    oai22 reg_nx3668 (.Y (nx3668), .A0 (nx4746), .A1 (nx4829), .B0 (nx4825), .B1 (
          nx4824)) ;
    or02 ix5414 (.Y (nx4752), .A0 (nx5995), .A1 (nx5997)) ;
    nor04_2x reg_nx492 (.Y (nx492), .A0 (nx5997), .A1 (nx5999), .A2 (nx6007), .A3 (
             nx6003)) ;
    inv01 ix5415 (.Y (nx4753), .A (nx4752)) ;
    nor02_2x ix5416 (.Y (nx4754), .A0 (nx5999), .A1 (nx6007)) ;
    inv01 ix5417 (.Y (nx4755), .A (M[1])) ;
    or03 ix5418 (.Y (nx4756), .A0 (nx6003), .A1 (nx5999), .A2 (nx6009)) ;
    inv02 ix5419 (.Y (nx4757), .A (nx5993)) ;
    aoi422 ix5420 (.Y (nx4758), .A0 (nx4753), .A1 (nx4754), .A2 (nx5993), .A3 (
           nx4755), .B0 (nx4756), .B1 (nx4757), .C0 (nx4752), .C1 (nx4757)) ;
    inv02 ix5421 (.Y (nx4759), .A (nx5989)) ;
    nand02_2x ix5422 (.Y (nx4760), .A0 (nx5989), .A1 (nx5991)) ;
    nand04_2x ix5423 (.Y (nx4761), .A0 (nx4978), .A1 (nx4979), .A2 (nx4759), .A3 (
              nx4980)) ;
    oai321 ix5424 (.Y (nx4762), .A0 (nx4979), .A1 (nx4759), .A2 (nx4980), .B0 (
           nx4978), .B1 (nx4760), .C0 (nx4761)) ;
    inv02 ix5425 (.Y (nx4763), .A (nx508)) ;
    inv02 ix5426 (.Y (nx4764), .A (nx5995)) ;
    inv01 ix5427 (.Y (nx4765), .A (nx492)) ;
    aoi22 ix5428 (.Y (nx4766), .A0 (nx492), .A1 (nx4764), .B0 (nx5995), .B1 (
          nx4765)) ;
    inv02 ix5429 (.Y (nx4767), .A (nx4978)) ;
    inv01 ix5430 (.Y (nx4768), .A (nx4979)) ;
    and02 ix5431 (.Y (nx4769), .A0 (nx4979), .A1 (nx4980)) ;
    oai422 reg_nx876 (.Y (nx876), .A0 (nx4767), .A1 (nx4768), .A2 (nx4759), .A3 (
           nx5991), .B0 (nx4769), .B1 (nx5989), .C0 (nx4978), .C1 (nx5989)) ;
    aoi322 ix5432 (.Y (nx4770), .A0 (nx4978), .A1 (nx5991), .A2 (nx4979), .B0 (
           nx4767), .B1 (nx4980), .C0 (nx4768), .C1 (nx4980)) ;
    inv01 reg_nx782 (.Y (nx782), .A (nx4770)) ;
    inv01 ix5433 (.Y (nx4771), .A (nx4770)) ;
    inv01 ix5434 (.Y (nx4772), .A (nx4770)) ;
    and02 reg_nx696 (.Y (nx696), .A0 (nx5210), .A1 (nx5212)) ;
    inv02 reg_nx688 (.Y (nx688), .A (nx5212)) ;
    inv02 ix5435 (.Y (nx4773), .A (nx5212)) ;
    oai22 reg_nx594 (.Y (nx594), .A0 (nx4764), .A1 (nx4765), .B0 (nx5995), .B1 (
          nx492)) ;
    inv01 ix5436 (.Y (nx4774), .A (nx4659)) ;
    nand02_2x ix5437 (.Y (nx4775), .A0 (nx5933), .A1 (nx4774)) ;
    inv01 ix5438 (.Y (nx4776), .A (nx5097)) ;
    and02 ix5439 (.Y (nx4777), .A0 (nx5224), .A1 (nx4659)) ;
    inv01 reg_nx4276 (.Y (nx4276), .A (nx4274_XX0_XREP44)) ;
    inv01 reg_nx4264 (.Y (nx4264), .A (nx4262)) ;
    inv02 ix5440 (.Y (nx4778), .A (negative_M_6)) ;
    inv02 ix5441 (.Y (nx4779), .A (positive_M_6)) ;
    oai22 reg_nx928 (.Y (nx928), .A0 (nx4778), .A1 (nx4322_XX0_XREP40), .B0 (
          nx4779), .B1 (nx5209)) ;
    aoi221 reg_nx3671 (.Y (nx3671), .A0 (positive_M_7), .A1 (nx4276), .B0 (
           negative_M_7), .B1 (nx4264), .C0 (nx928)) ;
    inv02 ix5442 (.Y (nx4780), .A (nx3663)) ;
    and02 ix5443 (.Y (nx4781), .A0 (nx3964), .A1 (nx3943)) ;
    aoi322 ix5444 (.Y (nx4782), .A0 (nx5200), .A1 (nx3943), .A2 (nx5931), .B0 (
           nx5200), .B1 (nx4781), .C0 (nx5931), .C1 (nx3964)) ;
    inv01 ix5445 (.Y (nx4783), .A (nx4782)) ;
    inv02 ix5446 (.Y (nx4784), .A (nx3964)) ;
    nor02_2x ix5447 (.Y (nx4785), .A0 (nx5931), .A1 (nx3964)) ;
    inv01 ix5448 (.Y (nx4786), .A (nx5221)) ;
    inv02 ix5449 (.Y (nx4787), .A (nx5221)) ;
    inv02 reg_nx3951 (.Y (nx3951), .A (nx5200)) ;
    inv02 ix5450 (.Y (nx4788), .A (nx3943)) ;
    and02 ix5451 (.Y (nx4789), .A0 (nx5200), .A1 (nx4788)) ;
    inv02 reg_nx1790 (.Y (nx1790), .A (nx4804)) ;
    inv01 ix5452 (.Y (nx4790), .A (nx4804)) ;
    inv01 ix5453 (.Y (nx4791), .A (nx4804)) ;
    inv02 ix5454 (.Y (nx4792), .A (nx4804)) ;
    inv02 ix5455 (.Y (nx4793), .A (nx4804)) ;
    inv02 ix5456 (.Y (nx4794), .A (nx4804)) ;
    or02 ix5457 (.Y (nx4795), .A0 (nx4784), .A1 (nx5931)) ;
    aoi21 reg_nx1850 (.Y (nx1850), .A0 (nx3964), .A1 (nx4795), .B0 (nx4785)) ;
    inv01 ix5458 (.Y (nx4796), .A (nx4782)) ;
    and02 ix5459 (.Y (nx4797), .A0 (nx5222), .A1 (nx3985)) ;
    inv01 ix5460 (.Y (nx4798), .A (nx5222)) ;
    inv02 ix5461 (.Y (nx4799), .A (nx3985)) ;
    oai21 ix5462 (.Y (nx4800), .A0 (nx4798), .A1 (nx4799), .B0 (nx4782)) ;
    oai332 ix5463 (.Y (nx4801), .A0 (nx5221), .A1 (nx4796), .A2 (nx4797), .B0 (
           nx4800), .B1 (nx4789), .B2 (nx5196), .C0 (nx5223), .C1 (nx3985)) ;
    nor02_2x ix5464 (.Y (nx4802), .A0 (nx5223), .A1 (nx3985)) ;
    inv01 ix5465 (.Y (nx4803), .A (nx4802)) ;
    nor02_2x ix5466 (.Y (nx4804), .A0 (nx4789), .A1 (nx5197)) ;
    nor02_2x ix5467 (.Y (nx4805), .A0 (nx4804), .A1 (nx4802)) ;
    aoi222 ix5468 (.Y (nx4806), .A0 (nx5223), .A1 (nx3985), .B0 (nx4803), .B1 (
           nx4796), .C0 (nx5221), .C1 (nx4805)) ;
    inv01 ix5469 (.Y (nx4807), .A (nx4806)) ;
    ao21 ix5470 (.Y (nx4808), .A0 (nx5223), .A1 (nx3985), .B0 (nx4802)) ;
    oai22 reg_nx1910 (.Y (nx1910), .A0 (nx4798), .A1 (nx3985), .B0 (nx4799), .B1 (
          nx5223)) ;
    inv01 ix5471 (.Y (nx4809), .A (nx3615)) ;
    inv02 ix5472 (.Y (nx4810), .A (nx3607)) ;
    aoi22 ix5473 (.Y (nx4811), .A0 (nx3615), .A1 (nx4810), .B0 (nx3607), .B1 (
          nx4809)) ;
    inv01 ix5474 (.Y (nx4812), .A (nx5907)) ;
    inv02 ix5475 (.Y (nx4813), .A (nx3574)) ;
    nor02_2x ix5476 (.Y (nx4814), .A0 (nx5917), .A1 (nx3550)) ;
    aoi22 ix5477 (.Y (nx4815), .A0 (nx5917), .A1 (nx3550), .B0 (nx5907), .B1 (
          nx3574)) ;
    aoi321 ix5478 (.Y (nx4816), .A0 (nx4684), .A1 (nx4685), .A2 (nx4686), .B0 (
           nx5915), .B1 (nx4687), .C0 (nx4714)) ;
    aoi222 ix5479 (.Y (nx4817), .A0 (nx4812), .A1 (nx4813), .B0 (nx4814), .B1 (
           nx4815), .C0 (nx4816), .C1 (nx4815)) ;
    inv02 ix5480 (.Y (nx4818), .A (nx3635)) ;
    inv01 ix5481 (.Y (nx4819), .A (nx5909)) ;
    aoi22 ix5482 (.Y (nx4820), .A0 (nx5909), .A1 (nx4818), .B0 (nx3635), .B1 (
          nx4819)) ;
    nor02_2x ix5483 (.Y (nx4821), .A0 (nx5061), .A1 (nx4820)) ;
    inv01 ix5484 (.Y (nx4822), .A (nx3640)) ;
    inv01 ix5485 (.Y (nx4823), .A (nx3640)) ;
    inv01 ix5486 (.Y (nx4824), .A (nx3640)) ;
    oai22 ix5487 (.Y (nx4825), .A0 (nx4818), .A1 (nx4819), .B0 (nx3635), .B1 (
          nx5909)) ;
    oai22 reg_nx744 (.Y (nx744), .A0 (nx4809), .A1 (nx3607), .B0 (nx4810), .B1 (
          nx3615)) ;
    oai22 ix5488 (.Y (nx4826), .A0 (nx4812), .A1 (nx4813), .B0 (nx5907), .B1 (
          nx3574)) ;
    oai22 reg_nx650 (.Y (nx650), .A0 (nx4813), .A1 (nx5907), .B0 (nx4812), .B1 (
          nx3574)) ;
    inv01 reg_nx838 (.Y (nx838), .A (nx4820)) ;
    inv01 ix5489 (.Y (nx4827), .A (nx4820)) ;
    inv01 ix5490 (.Y (nx4828), .A (nx4820)) ;
    inv01 ix5491 (.Y (nx4829), .A (nx4820)) ;
    nand02_2x ix5492 (.Y (nx4830), .A0 (nx5917), .A1 (nx3550)) ;
    and02 ix5493 (.Y (nx4831), .A0 (nx5917), .A1 (nx3550)) ;
    nor02_2x reg_nx602 (.Y (nx602), .A0 (nx4763), .A1 (nx4766)) ;
    inv02 ix5494 (.Y (nx4832), .A (nx5985)) ;
    inv02 ix5495 (.Y (nx4833), .A (M[10])) ;
    inv02 ix5496 (.Y (nx4834), .A (nx5981)) ;
    and04 ix5497 (.Y (nx4835), .A0 (nx5212), .A1 (nx4832), .A2 (nx4833), .A3 (
          nx4834)) ;
    and04 ix5498 (.Y (nx4836), .A0 (nx5213), .A1 (nx5985), .A2 (M[10]), .A3 (
          nx5981)) ;
    inv02 ix5499 (.Y (nx4837), .A (nx868)) ;
    aoi44 ix5500 (.Y (nx4838), .A0 (nx5211), .A1 (nx4835), .A2 (nx5939), .A3 (
          nx4762), .B0 (nx5210), .B1 (nx4836), .B2 (nx4762), .B3 (nx4837)) ;
    inv02 reg_nx1166 (.Y (nx1166), .A (nx4838)) ;
    inv02 ix5501 (.Y (nx4839), .A (nx4838)) ;
    or02 ix5502 (.Y (nx4840), .A0 (nx5985), .A1 (nx5981)) ;
    aoi422 ix5503 (.Y (nx4841), .A0 (nx5939), .A1 (nx4832), .A2 (M[10]), .A3 (
           nx4834), .B0 (nx4840), .B1 (nx4833), .C0 (nx4833), .C1 (nx4837)) ;
    inv02 reg_nx1158 (.Y (nx1158), .A (nx4841)) ;
    inv02 ix5504 (.Y (nx4842), .A (nx4841)) ;
    and02 ix5505 (.Y (nx4843), .A0 (nx5939), .A1 (nx4762)) ;
    nor02ii ix5506 (.Y (nx4844), .A0 (nx5939), .A1 (nx4762)) ;
    and02 ix5507 (.Y (nx4845), .A0 (nx5981), .A1 (nx5985)) ;
    aoi44 ix5508 (.Y (nx4846), .A0 (nx4843), .A1 (nx5211), .A2 (nx5213), .A3 (
          nx4977), .B0 (nx4844), .B1 (nx5211), .B2 (nx5213), .B3 (nx4845)) ;
    inv02 reg_nx1072 (.Y (nx1072), .A (nx4846)) ;
    inv02 ix5509 (.Y (nx4847), .A (nx4846)) ;
    oai322 reg_nx1064 (.Y (nx1064), .A0 (nx4837), .A1 (nx4834), .A2 (nx5985), .B0 (
           nx5981), .B1 (nx5939), .C0 (nx4832), .C1 (nx5981)) ;
    aoi44 ix5510 (.Y (nx4848), .A0 (nx4843), .A1 (nx5211), .A2 (nx5213), .A3 (
          nx4832), .B0 (nx4844), .B1 (nx5211), .B2 (nx5985), .B3 (nx5213)) ;
    inv02 reg_nx978 (.Y (nx978), .A (nx4848)) ;
    inv02 ix5511 (.Y (nx4849), .A (nx4848)) ;
    oai22 reg_nx970 (.Y (nx970), .A0 (nx4832), .A1 (nx4837), .B0 (nx5985), .B1 (
          nx5939)) ;
    oai21 ix5512 (.Y (nx4850), .A0 (nx5216), .A1 (nx4735), .B0 (nx4737)) ;
    nor02_2x ix5513 (.Y (nx4851), .A0 (nx5216), .A1 (nx4732)) ;
    and02 ix5514 (.Y (nx4852), .A0 (nx4738), .A1 (nx4851)) ;
    inv01 ix5515 (.Y (nx4853), .A (nx4694)) ;
    nor02_2x ix5516 (.Y (nx4854), .A0 (nx5216), .A1 (nx4735)) ;
    nor02ii ix5517 (.Y (nx4855), .A0 (nx4854), .A1 (nx4737)) ;
    nand02_2x ix5518 (.Y (nx4856), .A0 (nx5101), .A1 (nx4855)) ;
    nor02_2x ix5519 (.Y (nx4857), .A0 (M[14]), .A1 (nx5971)) ;
    inv02 ix5520 (.Y (nx4858), .A (nx5973)) ;
    inv02 ix5521 (.Y (nx4859), .A (nx5977)) ;
    and02 ix5523 (.Y (nx4861), .A0 (M[14]), .A1 (nx5971)) ;
    aoi44 ix5524 (.Y (nx4862), .A0 (nx4877), .A1 (nx4857), .A2 (nx4858), .A3 (
          nx4859), .B0 (nx5927), .B1 (nx4861), .B2 (nx5973), .B3 (nx5977)) ;
    nor02_2x reg_nx1542 (.Y (nx1542), .A0 (nx4862), .A1 (nx4838)) ;
    nor02_2x ix5525 (.Y (nx4863), .A0 (nx5973), .A1 (nx5977)) ;
    inv02 ix5526 (.Y (nx4864), .A (nx5971)) ;
    or03 ix5527 (.Y (nx4865), .A0 (nx5977), .A1 (nx5971), .A2 (nx5973)) ;
    inv02 ix5528 (.Y (nx4866), .A (M[14])) ;
    aoi422 ix5529 (.Y (nx4867), .A0 (nx4877), .A1 (nx4863), .A2 (M[14]), .A3 (
           nx4864), .B0 (nx4865), .B1 (nx4866), .C0 (nx5927), .C1 (nx4866)) ;
    inv02 reg_nx1534 (.Y (nx1534), .A (nx4867)) ;
    inv02 ix5530 (.Y (nx4868), .A (nx4867)) ;
    aoi44 ix5531 (.Y (nx4869), .A0 (nx4877), .A1 (nx4859), .A2 (nx4864), .A3 (
          nx4858), .B0 (nx5927), .B1 (nx5977), .B2 (nx5971), .B3 (nx5973)) ;
    nor02_2x reg_nx1448 (.Y (nx1448), .A0 (nx4869), .A1 (nx4838)) ;
    nor03_2x ix5532 (.Y (nx4870), .A0 (nx5977), .A1 (nx5971), .A2 (nx5973)) ;
    and02 reg_nx1432 (.Y (nx1432), .A0 (nx4877), .A1 (nx4870)) ;
    inv02 ix5533 (.Y (nx4871), .A (nx4863)) ;
    aoi422 ix5534 (.Y (nx4872), .A0 (nx4878), .A1 (nx4859), .A2 (nx5971), .A3 (
           nx4858), .B0 (nx4871), .B1 (nx4864), .C0 (nx5927), .C1 (nx4864)) ;
    inv02 reg_nx1440 (.Y (nx1440), .A (nx4872)) ;
    inv02 ix5535 (.Y (nx4873), .A (nx4872)) ;
    and02 ix5536 (.Y (nx4874), .A0 (nx5973), .A1 (nx5977)) ;
    aoi22 ix5537 (.Y (nx4875), .A0 (nx4878), .A1 (nx4863), .B0 (nx5927), .B1 (
          nx4874)) ;
    nor02_2x reg_nx1354 (.Y (nx1354), .A0 (nx4875), .A1 (nx4838)) ;
    oai322 reg_nx1346 (.Y (nx1346), .A0 (nx5927), .A1 (nx4858), .A2 (nx5979), .B0 (
           nx4878), .B1 (nx5975), .C0 (nx4859), .C1 (nx5975)) ;
    aoi22 ix5538 (.Y (nx4876), .A0 (nx4878), .A1 (nx4859), .B0 (nx5979), .B1 (
          nx5927)) ;
    nor02_2x reg_nx1260 (.Y (nx1260), .A0 (nx4876), .A1 (nx4838)) ;
    oai22 reg_nx1252 (.Y (nx1252), .A0 (nx4859), .A1 (nx5929), .B0 (nx4878), .B1 (
          nx5979)) ;
    buf04 ix5539 (.Y (nx4877), .A (nx1150)) ;
    buf04 ix5540 (.Y (nx4878), .A (nx1150)) ;
    ao22 reg_nx1846 (.Y (nx1846), .A0 (negative_M_17), .A1 (nx4476), .B0 (
         positive_M_17), .B1 (nx4466)) ;
    aoi221 reg_nx3972 (.Y (nx3972), .A0 (positive_M_18), .A1 (nx4280), .B0 (
           negative_M_18), .B1 (nx4268), .C0 (nx1846)) ;
    inv01 reg_nx4282 (.Y (nx4282), .A (nx4274)) ;
    inv01 reg_nx4478 (.Y (nx4478), .A (nx4322)) ;
    nor02_2x ix5541 (.Y (nx4879), .A0 (nx5237), .A1 (nx4111)) ;
    inv02 ix5542 (.Y (nx4880), .A (nx5129)) ;
    inv02 ix5543 (.Y (nx4881), .A (nx4111)) ;
    and02 ix5544 (.Y (nx4882), .A0 (nx5237), .A1 (nx4881)) ;
    nor02_2x ix5545 (.Y (nx4883), .A0 (nx4881), .A1 (nx5237)) ;
    nor02_2x ix5546 (.Y (nx4884), .A0 (nx4882), .A1 (nx4883)) ;
    inv02 reg_nx2270 (.Y (nx2270), .A (nx4884)) ;
    inv02 ix5547 (.Y (nx4885), .A (nx4884)) ;
    inv02 ix5548 (.Y (nx4886), .A (nx4884)) ;
    inv01 ix5549 (.Y (nx4887), .A (nx4884)) ;
    inv02 ix5550 (.Y (nx4888), .A (nx4884)) ;
    nor04_2x reg_nx4053 (.Y (nx4053), .A0 (nx5937), .A1 (nx4966), .A2 (nx5043), 
             .A3 (nx4964)) ;
    and02 ix5551 (.Y (nx4889), .A0 (nx4623), .A1 (nx5129)) ;
    oai22 ix5552 (.Y (nx4890), .A0 (nx4889), .A1 (nx5146), .B0 (nx4623), .B1 (
          nx5140)) ;
    and02 ix5553 (.Y (nx4891), .A0 (nx4636), .A1 (nx5132)) ;
    inv01 ix5554 (.Y (nx4892), .A (nx4633)) ;
    nor02_2x ix5555 (.Y (nx4893), .A0 (nx4632), .A1 (nx5124)) ;
    nand02_2x ix5556 (.Y (nx4894), .A0 (nx4623), .A1 (nx5147)) ;
    aoi44 ix5557 (.Y (nx4895), .A0 (nx4890), .A1 (nx4891), .A2 (nx4892), .A3 (
          nx4893), .B0 (nx4894), .B1 (nx5169), .B2 (nx4636), .B3 (nx5136)) ;
    inv01 ix5558 (.Y (nx4896), .A (nx4642)) ;
    inv01 ix5559 (.Y (nx4897), .A (nx4631)) ;
    and03 ix5560 (.Y (nx4898), .A0 (nx4895), .A1 (nx4896), .A2 (nx4897)) ;
    aoi21 ix5561 (.Y (nx4899), .A0 (nx5148), .A1 (nx5141), .B0 (nx4632)) ;
    nor02_2x ix5562 (.Y (nx4900), .A0 (nx5169), .A1 (nx4899)) ;
    nor02_2x ix5563 (.Y (nx4901), .A0 (nx4889), .A1 (nx4633)) ;
    nor02_2x ix5564 (.Y (nx4902), .A0 (nx5169), .A1 (nx4901)) ;
    nand02_2x ix5565 (.Y (nx4903), .A0 (nx4636), .A1 (nx5136)) ;
    or04 ix5566 (.Y (nx4904), .A0 (nx4900), .A1 (nx5171), .A2 (nx4902), .A3 (
         nx4903)) ;
    oai21 ix5567 (.Y (nx4905), .A0 (nx4889), .A1 (nx4633), .B0 (nx5175)) ;
    ao21 ix5568 (.Y (nx4906), .A0 (nx5961), .A1 (nx5142), .B0 (nx4632)) ;
    nand02_2x ix5569 (.Y (nx4907), .A0 (nx5176), .A1 (nx4906)) ;
    and02 ix5570 (.Y (nx4908), .A0 (nx4623), .A1 (nx5961)) ;
    oai21 ix5571 (.Y (nx4909), .A0 (nx4908), .A1 (nx5124), .B0 (nx5177)) ;
    nor02ii ix5572 (.Y (nx4910), .A0 (nx5155), .A1 (nx4717)) ;
    nor02ii ix5573 (.Y (nx4911), .A0 (nx4720), .A1 (nx4701)) ;
    oai22 reg_nx4221 (.Y (nx4221), .A0 (nx4910), .A1 (nx5206), .B0 (nx4911), .B1 (
          nx5205)) ;
    inv01 ix5574 (.Y (nx4912), .A (nx4701)) ;
    and02 ix5575 (.Y (nx4913), .A0 (nx5230), .A1 (nx4027)) ;
    nor02_2x ix5576 (.Y (nx4914), .A0 (nx5230), .A1 (nx4027)) ;
    inv01 ix5577 (.Y (nx4915), .A (nx5224)) ;
    inv02 ix5578 (.Y (nx4916), .A (nx4006)) ;
    nor03_2x ix5579 (.Y (nx4917), .A0 (nx4914), .A1 (nx4915), .A2 (nx4916)) ;
    nor04_2x ix5580 (.Y (nx4918), .A0 (nx4913), .A1 (nx4631), .A2 (nx4917), .A3 (
             nx4642)) ;
    inv01 ix5581 (.Y (nx4919), .A (nx4918)) ;
    inv01 ix5582 (.Y (nx4920), .A (nx4918)) ;
    aoi21 ix5583 (.Y (nx4921), .A0 (nx5230), .A1 (nx4027), .B0 (nx4914)) ;
    inv01 ix5584 (.Y (nx4922), .A (nx4921)) ;
    inv01 ix5585 (.Y (nx4923), .A (nx5933)) ;
    inv01 ix5586 (.Y (nx4924), .A (nx5933)) ;
    inv01 ix5587 (.Y (nx4925), .A (nx5933)) ;
    inv01 ix5588 (.Y (nx4926), .A (nx5933)) ;
    inv01 ix5589 (.Y (nx4927), .A (nx5933)) ;
    oai22 reg_nx1970 (.Y (nx1970), .A0 (nx4915), .A1 (nx4006), .B0 (nx4916), .B1 (
          nx5224)) ;
    inv02 ix5590 (.Y (nx4928), .A (nx4027)) ;
    inv01 ix5591 (.Y (nx4929), .A (nx5231)) ;
    aoi22 ix5592 (.Y (nx4930), .A0 (nx5231), .A1 (nx4928), .B0 (nx4027), .B1 (
          nx4929)) ;
    inv01 reg_nx2030 (.Y (nx2030), .A (nx4930)) ;
    inv01 ix5593 (.Y (nx4931), .A (nx4930)) ;
    inv01 ix5594 (.Y (nx4932), .A (nx4930)) ;
    inv01 ix5595 (.Y (nx4933), .A (nx4930)) ;
    inv01 ix5596 (.Y (nx4934), .A (nx4930)) ;
    inv01 ix5597 (.Y (nx4935), .A (nx4930)) ;
    inv02 ix5598 (.Y (nx4936), .A (nx3719)) ;
    nor02ii ix5599 (.Y (nx4937), .A0 (nx5079), .A1 (nx4821)) ;
    nand02_2x ix5600 (.Y (nx4938), .A0 (nx4809), .A1 (nx4811)) ;
    and02 ix5601 (.Y (nx4939), .A0 (nx5016), .A1 (nx5010)) ;
    aoi321 ix5602 (.Y (nx4940), .A0 (nx4937), .A1 (nx5063), .A2 (nx4938), .B0 (
           nx5192), .B1 (nx4939), .C0 (nx5005)) ;
    inv01 ix5603 (.Y (nx4941), .A (nx4739)) ;
    inv01 ix5604 (.Y (nx4942), .A (nx4740)) ;
    inv01 ix5605 (.Y (nx4943), .A (nx4741)) ;
    oai321 ix5606 (.Y (nx4944), .A0 (nx4940), .A1 (nx5214), .A2 (nx4941), .B0 (
           nx4941), .B1 (nx4942), .C0 (nx4943)) ;
    and02 ix5607 (.Y (nx4945), .A0 (nx4809), .A1 (nx4811)) ;
    ao21 ix5608 (.Y (nx4946), .A0 (nx5017), .A1 (nx5011), .B0 (nx5006)) ;
    or02 ix5609 (.Y (nx4947), .A0 (nx5007), .A1 (nx5192)) ;
    oai21 ix5610 (.Y (nx4948), .A0 (nx4740), .A1 (nx4959), .B0 (nx4739)) ;
    aoi32 reg_nx3836 (.Y (nx3836), .A0 (nx5957), .A1 (nx4943), .A2 (nx4942), .B0 (
          nx4948), .B1 (nx4943)) ;
    ao22 reg_nx2326 (.Y (nx2326), .A0 (negative_M_25), .A1 (nx4478), .B0 (
         positive_M_25), .B1 (nx4468)) ;
    aoi221 reg_nx4140 (.Y (nx4140), .A0 (positive_M_26), .A1 (nx4282), .B0 (
           negative_M_26), .B1 (nx4270), .C0 (nx2326)) ;
    inv02 ix5611 (.Y (nx4949), .A (negative_M_9)) ;
    inv02 ix5612 (.Y (nx4950), .A (positive_M_9)) ;
    oai22 reg_nx1210 (.Y (nx1210), .A0 (nx4949), .A1 (nx4322_XX0_XREP40), .B0 (
          nx4950), .B1 (nx5209)) ;
    aoi221 reg_nx3755 (.Y (nx3755), .A0 (positive_M_10), .A1 (nx4278), .B0 (
           negative_M_10), .B1 (nx4266), .C0 (nx1210)) ;
    inv02 ix5613 (.Y (nx4951), .A (nx3747)) ;
    and02 ix5614 (.Y (nx4952), .A0 (nx5935), .A1 (nx4951)) ;
    nor02_2x ix5615 (.Y (nx4953), .A0 (nx4951), .A1 (nx5935)) ;
    nor02_2x ix5616 (.Y (nx4954), .A0 (nx4952), .A1 (nx4953)) ;
    inv02 reg_nx1214 (.Y (nx1214), .A (nx5214)) ;
    inv01 ix5617 (.Y (nx4955), .A (nx5215)) ;
    inv01 ix5618 (.Y (nx4956), .A (nx5215)) ;
    inv01 ix5619 (.Y (nx4957), .A (nx5215)) ;
    inv02 ix5620 (.Y (nx4958), .A (nx5215)) ;
    inv02 ix5621 (.Y (nx4959), .A (nx5215)) ;
    nand02_2x ix5622 (.Y (nx4960), .A0 (nx4727), .A1 (nx5919)) ;
    nand02_2x ix5623 (.Y (nx4961), .A0 (nx4728), .A1 (nx5919)) ;
    inv01 ix5624 (.Y (nx4962), .A (nx4853)) ;
    inv01 ix5625 (.Y (nx4963), .A (nx5955)) ;
    aoi321 ix5626 (.Y (nx4964), .A0 (nx4960), .A1 (nx4961), .A2 (nx4962), .B0 (
           nx4682), .B1 (nx4775), .C0 (nx4963)) ;
    aoi21 ix5627 (.Y (nx4965), .A0 (nx4856), .A1 (nx4738), .B0 (nx4853)) ;
    nor04_2x ix5628 (.Y (nx4966), .A0 (nx4965), .A1 (nx4776), .A2 (nx4777), .A3 (
             nx5231)) ;
    oai22 ix5629 (.Y (nx4967), .A0 (nx4924), .A1 (nx4933), .B0 (nx5225), .B1 (
          nx4923)) ;
    nor02ii ix5630 (.Y (nx4968), .A0 (nx5098), .A1 (nx4967)) ;
    oai321 reg_nx4011 (.Y (nx4011), .A0 (nx4727), .A1 (nx4853), .A2 (nx4728), .B0 (
           nx4853), .B1 (nx5919), .C0 (nx5955)) ;
    inv01 ix5631 (.Y (nx4969), .A (nx4158)) ;
    inv02 ix5632 (.Y (nx4970), .A (nx5241)) ;
    and02 ix5633 (.Y (nx4971), .A0 (nx5229), .A1 (nx4452)) ;
    oai221 reg_nx4155 (.Y (nx4155), .A0 (nx4969), .A1 (nx5241), .B0 (nx4970), .B1 (
           nx4158), .C0 (nx4971)) ;
    nor02_2x ix5634 (.Y (nx4972), .A0 (nx5995), .A1 (nx5997)) ;
    nor02_2x ix5635 (.Y (nx4973), .A0 (nx6005), .A1 (nx5993)) ;
    nor02_2x ix5636 (.Y (nx4974), .A0 (nx5991), .A1 (nx6001)) ;
    nor04_2x ix5637 (.Y (nx4975), .A0 (nx5981), .A1 (nx6009), .A2 (nx5989), .A3 (
             nx5987)) ;
    and04 reg_nx1056 (.Y (nx1056), .A0 (nx4972), .A1 (nx4973), .A2 (nx4974), .A3 (
          nx4975)) ;
    nor02_2x ix5638 (.Y (nx4976), .A0 (nx6009), .A1 (nx5989)) ;
    and04 reg_nx868 (.Y (nx868), .A0 (nx4972), .A1 (nx4974), .A2 (nx4973), .A3 (
          nx4976)) ;
    nor02_2x ix5639 (.Y (nx4977), .A0 (nx5983), .A1 (nx5987)) ;
    nor02_2x ix5640 (.Y (nx4978), .A0 (nx6005), .A1 (nx6009)) ;
    nor04_2x ix5641 (.Y (nx4979), .A0 (nx5997), .A1 (nx6001), .A2 (nx5995), .A3 (
             nx5993)) ;
    inv02 ix5642 (.Y (nx4980), .A (nx5991)) ;
    nor03_2x ix5643 (.Y (nx4981), .A0 (nx4618), .A1 (nx5227), .A2 (nx5233)) ;
    inv01 ix5644 (.Y (nx4982), .A (nx4158)) ;
    nor02_2x ix5645 (.Y (nx4983), .A0 (nx4621), .A1 (nx4637)) ;
    aoi32 ix5646 (.Y (nx4984), .A0 (nx4158), .A1 (nx5241), .A2 (nx4981), .B0 (
          nx4982), .B1 (nx4983)) ;
    inv02 ix5647 (.Y (nx4985), .A (nx4304)) ;
    inv02 ix5648 (.Y (nx4986), .A (nx4174)) ;
    inv02 ix5649 (.Y (nx4987), .A (nx5241)) ;
    aoi322 ix5650 (.Y (nx4988), .A0 (nx4981), .A1 (nx4412), .A2 (nx4595), .B0 (
           nx4985), .B1 (nx4986), .C0 (nx4983), .C1 (nx4987)) ;
    nand02_2x reg_nx3378 (.Y (nx3378), .A0 (nx4984), .A1 (nx4988)) ;
    ao22 reg_nx2146 (.Y (nx2146), .A0 (negative_M_22), .A1 (nx4478_XX0_XREP64), 
         .B0 (positive_M_22), .B1 (nx4468)) ;
    aoi221 reg_nx4077 (.Y (nx4077), .A0 (positive_M_23), .A1 (nx4282), .B0 (
           negative_M_23), .B1 (nx4270), .C0 (nx2146)) ;
    ao221 reg_nx3408 (.Y (nx3408), .A0 (nx4158), .A1 (nx4596), .B0 (nx4583), .B1 (
          nx5045), .C0 (nx5913)) ;
    inv02 ix5651 (.Y (nx4989), .A (nx4132)) ;
    inv01 reg_nx4266 (.Y (nx4266), .A (nx4262)) ;
    inv02 ix5652 (.Y (nx4990), .A (negative_M_11)) ;
    inv02 ix5653 (.Y (nx4991), .A (positive_M_11)) ;
    oai22 reg_nx1398 (.Y (nx1398), .A0 (nx4990), .A1 (nx4322_XX0_XREP40), .B0 (
          nx4991), .B1 (nx5209)) ;
    aoi221 reg_nx3811 (.Y (nx3811), .A0 (positive_M_12), .A1 (nx4278), .B0 (
           negative_M_12), .B1 (nx4266), .C0 (nx1398)) ;
    inv02 ix5654 (.Y (nx4992), .A (nx3803)) ;
    and02 ix5655 (.Y (nx4993), .A0 (nx3811), .A1 (nx4992)) ;
    nor02_2x ix5656 (.Y (nx4994), .A0 (nx4992), .A1 (nx3811)) ;
    nor02_2x ix5657 (.Y (nx4995), .A0 (nx4993), .A1 (nx4994)) ;
    inv02 reg_nx1402 (.Y (nx1402), .A (nx5217)) ;
    inv02 ix5658 (.Y (nx4996), .A (nx5217)) ;
    inv01 ix5659 (.Y (nx4997), .A (nx5217)) ;
    inv01 ix5660 (.Y (nx4998), .A (nx5217)) ;
    inv01 ix5661 (.Y (nx4999), .A (nx5217)) ;
    inv01 reg_nx4474 (.Y (nx4474), .A (nx4322_XX0_XREP40)) ;
    inv01 reg_nx4464 (.Y (nx4464), .A (nx5209)) ;
    inv01 reg_nx4278 (.Y (nx4278), .A (nx4274_XX0_XREP44)) ;
    ao21 ix5662 (.Y (nx5000), .A0 (nx3691), .A1 (nx5947), .B0 (nx3719)) ;
    ao22 reg_nx1116 (.Y (nx1116), .A0 (negative_M_8), .A1 (nx4474), .B0 (
         positive_M_8), .B1 (nx4464)) ;
    aoi221 ix5663 (.Y (nx5001), .A0 (positive_M_9), .A1 (nx4278), .B0 (
           negative_M_9), .B1 (nx4266), .C0 (nx1116)) ;
    inv02 ix5664 (.Y (nx5002), .A (nx3691)) ;
    nor02_2x ix5665 (.Y (nx5003), .A0 (nx5002), .A1 (nx4936)) ;
    aoi22 ix5666 (.Y (nx5004), .A0 (nx5000), .A1 (nx5943), .B0 (nx5947), .B1 (
          nx5003)) ;
    inv01 ix5667 (.Y (nx5005), .A (nx5004)) ;
    inv01 ix5668 (.Y (nx5006), .A (nx5004)) ;
    inv01 ix5669 (.Y (nx5007), .A (nx5004)) ;
    inv01 reg_nx3699 (.Y (nx3699), .A (nx5044)) ;
    aoi22 ix5670 (.Y (nx5008), .A0 (nx3691), .A1 (nx3699), .B0 (nx5947), .B1 (
          nx5002)) ;
    inv01 reg_nx1026 (.Y (nx1026), .A (nx5008)) ;
    inv01 ix5671 (.Y (nx5009), .A (nx5945)) ;
    inv01 ix5672 (.Y (nx5010), .A (nx5945)) ;
    inv01 ix5673 (.Y (nx5011), .A (nx5945)) ;
    inv01 ix5674 (.Y (nx5012), .A (nx5947)) ;
    inv02 ix5675 (.Y (nx5013), .A (nx3719)) ;
    nor02_2x ix5676 (.Y (nx5014), .A0 (nx5943), .A1 (nx4936)) ;
    aoi21 ix5677 (.Y (nx5015), .A0 (nx5943), .A1 (nx5013), .B0 (nx5014)) ;
    inv01 reg_nx1120 (.Y (nx1120), .A (nx5015)) ;
    inv01 ix5678 (.Y (nx5016), .A (nx5015)) ;
    inv01 ix5679 (.Y (nx5017), .A (nx5015)) ;
    inv02 ix5680 (.Y (nx5018), .A (nx4069)) ;
    inv01 ix5681 (.Y (nx5019), .A (nx5941)) ;
    aoi22 ix5682 (.Y (nx5020), .A0 (nx5941), .A1 (nx5018), .B0 (nx4069), .B1 (
          nx5019)) ;
    inv01 reg_nx2150 (.Y (nx2150), .A (nx5028)) ;
    inv01 ix5683 (.Y (nx5021), .A (nx5028)) ;
    inv01 ix5684 (.Y (nx5022), .A (nx5028)) ;
    inv01 ix5685 (.Y (nx5023), .A (nx5028)) ;
    inv01 ix5686 (.Y (nx5024), .A (nx5029)) ;
    inv01 ix5687 (.Y (nx5025), .A (nx5029)) ;
    inv01 ix5688 (.Y (nx5026), .A (nx5029)) ;
    inv01 ix5689 (.Y (nx5027), .A (nx5029)) ;
    buf02 ix5690 (.Y (nx5028), .A (nx5020)) ;
    buf02 ix5691 (.Y (nx5029), .A (nx5020)) ;
    inv01 ix5692 (.Y (nx5030), .A (nx4655)) ;
    nor02_2x ix5693 (.Y (nx5031), .A0 (nx5225), .A1 (nx4926)) ;
    nor02_2x ix5694 (.Y (nx5032), .A0 (nx4927), .A1 (nx4934)) ;
    nand02_2x ix5695 (.Y (nx5033), .A0 (nx5225), .A1 (nx4935)) ;
    inv01 ix5696 (.Y (nx5034), .A (nx5231)) ;
    inv01 ix5697 (.Y (nx5035), .A (nx4659)) ;
    ao21 ix5698 (.Y (nx5036), .A0 (nx5033), .A1 (nx5034), .B0 (nx5035)) ;
    aoi21 ix5699 (.Y (nx5037), .A0 (nx5231), .A1 (nx4925), .B0 (nx4655)) ;
    aoi222 ix5700 (.Y (nx5038), .A0 (nx5030), .A1 (nx5031), .B0 (nx5030), .B1 (
           nx5032), .C0 (nx5036), .C1 (nx5037)) ;
    and04 ix5701 (.Y (nx5039), .A0 (nx5021), .A1 (nx5169), .A2 (nx2210), .A3 (
          nx5235)) ;
    nand02_2x ix5702 (.Y (nx5040), .A0 (nx5038), .A1 (nx5039)) ;
    nand03_2x ix5703 (.Y (nx5041), .A0 (nx4935), .A1 (nx4659), .A2 (nx5225)) ;
    oai222 ix5704 (.Y (nx5042), .A0 (nx4659), .A1 (nx4925), .B0 (nx5225), .B1 (
           nx4926), .C0 (nx4927), .C1 (nx4934)) ;
    ao32 ix5705 (.Y (nx5043), .A0 (nx5041), .A1 (nx5030), .A2 (nx5034), .B0 (
         nx5042), .B1 (nx5030)) ;
    ao22 reg_nx1022 (.Y (nx1022), .A0 (negative_M_7), .A1 (nx4474), .B0 (
         positive_M_7), .B1 (nx4464)) ;
    aoi221 ix5706 (.Y (nx5044), .A0 (positive_M_8), .A1 (nx4278), .B0 (nx4266), 
           .B1 (negative_M_8), .C0 (nx1022)) ;
    inv01 ix5707 (.Y (nx5045), .A (nx4221)) ;
    and02 ix5708 (.Y (nx5046), .A0 (positive_M_24), .A1 (nx4468)) ;
    and02 ix5709 (.Y (nx5047), .A0 (positive_M_25), .A1 (nx4282)) ;
    and02 ix5710 (.Y (nx5048), .A0 (negative_M_25), .A1 (nx4270)) ;
    inv02 ix5711 (.Y (nx5049), .A (nx4111)) ;
    ao21 ix5712 (.Y (nx5050), .A0 (negative_M_24), .A1 (nx4478), .B0 (nx5049)) ;
    nor04_2x ix5713 (.Y (nx5051), .A0 (nx5046), .A1 (nx5047), .A2 (nx5048), .A3 (
             nx5050)) ;
    inv01 ix5714 (.Y (nx5052), .A (nx5129)) ;
    and02 ix5715 (.Y (nx5053), .A0 (negative_M_24), .A1 (nx4478)) ;
    nor04_2x reg_nx4119 (.Y (nx4119), .A0 (nx5046), .A1 (nx5053), .A2 (nx5048), 
             .A3 (nx5047)) ;
    inv01 ix5716 (.Y (nx5054), .A (nx3671)) ;
    inv02 ix5717 (.Y (nx5055), .A (nx4780)) ;
    aoi22 ix5718 (.Y (nx5056), .A0 (nx4780), .A1 (nx5054), .B0 (nx3671), .B1 (
          nx5055)) ;
    inv01 ix5719 (.Y (nx5057), .A (nx5062)) ;
    inv01 ix5720 (.Y (nx5058), .A (nx5062)) ;
    inv01 ix5721 (.Y (nx5059), .A (nx5062)) ;
    inv01 ix5722 (.Y (nx5060), .A (nx5062)) ;
    inv01 ix5723 (.Y (nx5061), .A (nx932)) ;
    buf02 ix5724 (.Y (nx5062), .A (nx5056)) ;
    buf02 reg_nx932 (.Y (nx932), .A (nx5056)) ;
    nor02_2x ix5725 (.Y (nx5063), .A0 (nx5015), .A1 (nx5945)) ;
    ao22 reg_nx1586 (.Y (nx1586), .A0 (negative_M_13), .A1 (nx4476), .B0 (
         positive_M_13), .B1 (nx4466)) ;
    aoi221 reg_nx3867 (.Y (nx3867), .A0 (positive_M_14), .A1 (nx4278), .B0 (
           negative_M_14), .B1 (nx4266), .C0 (nx1586)) ;
    inv02 ix5726 (.Y (nx5064), .A (nx3859)) ;
    and02 ix5727 (.Y (nx5065), .A0 (nx5949), .A1 (nx5064)) ;
    nor02_2x ix5728 (.Y (nx5066), .A0 (nx5064), .A1 (nx5949)) ;
    nor02_2x ix5729 (.Y (nx5067), .A0 (nx5065), .A1 (nx5066)) ;
    ao22 reg_nx1492 (.Y (nx1492), .A0 (negative_M_12), .A1 (nx4474), .B0 (
         positive_M_12), .B1 (nx4464)) ;
    aoi221 reg_nx3839 (.Y (nx3839), .A0 (nx4278), .A1 (positive_M_13), .B0 (
           nx4266), .B1 (negative_M_13), .C0 (nx1492)) ;
    inv02 ix5730 (.Y (nx5068), .A (nx3831)) ;
    and02 ix5731 (.Y (nx5069), .A0 (nx5951), .A1 (nx5068)) ;
    nor02_2x ix5732 (.Y (nx5070), .A0 (nx5068), .A1 (nx5951)) ;
    nor02_2x ix5733 (.Y (nx5071), .A0 (nx5069), .A1 (nx5070)) ;
    nor02_2x ix5734 (.Y (nx5072), .A0 (nx5067), .A1 (nx5071)) ;
    inv02 reg_nx1590 (.Y (nx1590), .A (nx5067)) ;
    inv01 ix5735 (.Y (nx5073), .A (nx5067)) ;
    inv01 ix5736 (.Y (nx5074), .A (nx5067)) ;
    inv02 reg_nx1496 (.Y (nx1496), .A (nx5071)) ;
    inv01 ix5737 (.Y (nx5075), .A (nx5071)) ;
    inv02 ix5738 (.Y (nx5076), .A (nx5071)) ;
    inv02 ix5739 (.Y (nx5077), .A (nx5229)) ;
    inv02 ix5740 (.Y (nx5078), .A (nx4069)) ;
    ao22 reg_nx1304 (.Y (nx1304), .A0 (negative_M_10), .A1 (nx4474), .B0 (
         positive_M_10), .B1 (nx4464)) ;
    nor02_2x ix5741 (.Y (nx5079), .A0 (nx4811), .A1 (nx4817)) ;
    nor02_2x reg_nx3640 (.Y (nx3640), .A0 (nx5079), .A1 (nx4945)) ;
    inv01 ix5742 (.Y (nx5080), .A (nx2450)) ;
    inv02 ix5743 (.Y (nx5081), .A (nx5241)) ;
    or04 ix5744 (.Y (nx5082), .A0 (nx5117), .A1 (nx4605), .A2 (nx5080), .A3 (
         nx5081)) ;
    ao32 ix5745 (.Y (nx5083), .A0 (nx4595), .A1 (nx2450), .A2 (nx4412), .B0 (
         nx4414), .B1 (nx5152)) ;
    inv02 ix5746 (.Y (nx5084), .A (nx4605)) ;
    nand02_2x ix5747 (.Y (nx5085), .A0 (nx5083), .A1 (nx5084)) ;
    or02 ix5748 (.Y (nx5086), .A0 (nx4304), .A1 (nx4195)) ;
    nand04_2x reg_nx3388 (.Y (nx3388), .A0 (nx5082), .A1 (nx5085), .A2 (nx5114)
              , .A3 (nx5086)) ;
    inv01 ix5749 (.Y (nx5087), .A (nx5152)) ;
    inv01 ix5750 (.Y (nx5088), .A (nx4412)) ;
    inv01 ix5751 (.Y (nx5089), .A (nx4414)) ;
    inv01 ix5752 (.Y (nx5090), .A (nx4595)) ;
    nor02_2x ix5753 (.Y (nx5091), .A0 (nx4414), .A1 (nx4412)) ;
    nor02_2x ix5754 (.Y (nx5092), .A0 (nx4414), .A1 (nx5241)) ;
    aoi332 ix5755 (.Y (nx5093), .A0 (nx5081), .A1 (nx5089), .A2 (nx5088), .B0 (
           nx5090), .B1 (nx5087), .B2 (nx5081), .C0 (nx5090), .C1 (nx5092)) ;
    aoi322 ix5756 (.Y (nx5094), .A0 (nx5087), .A1 (nx5088), .A2 (nx5081), .B0 (
           nx5087), .B1 (nx5080), .C0 (nx5089), .C1 (nx5080)) ;
    nand02_2x ix5757 (.Y (nx5095), .A0 (nx5093), .A1 (nx5094)) ;
    aoi221 reg_nx3783 (.Y (nx3783), .A0 (negative_M_11), .A1 (nx4266), .B0 (
           positive_M_11), .B1 (nx4278), .C0 (nx1304)) ;
    ao221 ix5758 (.Y (nx5096), .A0 (nx4738), .A1 (nx4850), .B0 (nx5957), .B1 (
          nx4852), .C0 (nx4853)) ;
    aoi32 ix5759 (.Y (nx5097), .A0 (nx4698), .A1 (nx4376), .A2 (nx4678), .B0 (
          nx4700), .B1 (nx4807)) ;
    nand02_2x ix5760 (.Y (nx5098), .A0 (nx5096), .A1 (nx5955)) ;
    nand03_2x ix5761 (.Y (nx5099), .A0 (nx4821), .A1 (nx3640), .A2 (nx5063)) ;
    nand02_2x ix5762 (.Y (nx5100), .A0 (nx4946), .A1 (nx4947)) ;
    nand03_2x ix5763 (.Y (nx5101), .A0 (nx5099), .A1 (nx4851), .A2 (nx5100)) ;
    aoi32 ix5764 (.Y (nx5102), .A0 (nx4821), .A1 (nx3640), .A2 (nx5063), .B0 (
          nx4946), .B1 (nx4947)) ;
    inv02 ix5765 (.Y (nx5103), .A (nx5095)) ;
    inv01 ix5766 (.Y (nx5104), .A (nx4628)) ;
    or03 ix5767 (.Y (nx5105), .A0 (nx5040), .A1 (nx5937), .A2 (nx4964)) ;
    aoi22 ix5768 (.Y (nx5106), .A0 (nx4966), .A1 (nx5104), .B0 (nx5105), .B1 (
          nx5104)) ;
    nand02_2x ix5769 (.Y (nx5107), .A0 (nx5103), .A1 (nx5106)) ;
    nand02_2x ix5770 (.Y (nx5108), .A0 (nx5087), .A1 (nx5088)) ;
    inv02 ix5771 (.Y (nx5109), .A (nx5090)) ;
    inv02 ix5772 (.Y (nx5110), .A (nx5087)) ;
    inv02 ix5773 (.Y (nx5111), .A (nx5089)) ;
    aoi22 ix5774 (.Y (nx5112), .A0 (nx5108), .A1 (nx5109), .B0 (nx5110), .B1 (
          nx5111)) ;
    or03 ix5775 (.Y (nx5113), .A0 (nx5095), .A1 (nx5112), .A2 (nx5091)) ;
    nand04_2x ix5776 (.Y (nx5114), .A0 (nx5107), .A1 (nx5113), .A2 (nx4606), .A3 (
              nx4607)) ;
    inv01 ix5777 (.Y (nx5115), .A (nx4966)) ;
    nor03_2x ix5778 (.Y (nx5116), .A0 (nx5040), .A1 (nx5937), .A2 (nx4964)) ;
    oai22 ix5779 (.Y (nx5117), .A0 (nx5115), .A1 (nx4628), .B0 (nx5116), .B1 (
          nx4628)) ;
    inv02 ix5780 (.Y (nx5118), .A (nx5229)) ;
    inv02 ix5781 (.Y (nx5119), .A (nx4452)) ;
    or03 ix5782 (.Y (nx5120), .A0 (nx2150), .A1 (nx5118), .A2 (nx5119)) ;
    and02 ix5783 (.Y (nx5121), .A0 (nx5229), .A1 (nx4452)) ;
    aoi32 ix5784 (.Y (nx5122), .A0 (nx4074), .A1 (nx2150), .A2 (nx5121), .B0 (
          nx5077), .B1 (nx5078)) ;
    oai21 reg_nx3328 (.Y (nx3328), .A0 (nx4074), .A1 (nx5120), .B0 (nx5122)) ;
    inv01 ix5785 (.Y (nx5123), .A (nx5237)) ;
    nor02_2x ix5786 (.Y (nx5124), .A0 (nx5237), .A1 (nx5238)) ;
    inv02 ix5787 (.Y (nx5125), .A (nx4989)) ;
    nor02_2x ix5788 (.Y (nx5126), .A0 (nx5125), .A1 (nx5123)) ;
    and02 ix5789 (.Y (nx5127), .A0 (nx4132), .A1 (nx5237)) ;
    nor02_2x ix5790 (.Y (nx5128), .A0 (nx5126), .A1 (nx5127)) ;
    nor02_2x ix5791 (.Y (nx5129), .A0 (nx5051), .A1 (nx4879)) ;
    inv01 ix5792 (.Y (nx5130), .A (nx5239)) ;
    nor02_2x ix5793 (.Y (nx5131), .A0 (nx4132), .A1 (nx4989)) ;
    oai22 ix5794 (.Y (nx5132), .A0 (nx5128), .A1 (nx5129), .B0 (nx5130), .B1 (
          nx5131)) ;
    inv01 ix5795 (.Y (nx5133), .A (nx5123)) ;
    oai22 ix5796 (.Y (nx5134), .A0 (nx5133), .A1 (nx5127), .B0 (nx5051), .B1 (
          nx4879)) ;
    oai21 ix5797 (.Y (nx5135), .A0 (nx5239), .A1 (nx5237), .B0 (nx4132)) ;
    aoi22 ix5798 (.Y (nx5136), .A0 (nx5134), .A1 (nx5130), .B0 (nx5135), .B1 (
          nx5125)) ;
    inv02 ix5799 (.Y (nx5137), .A (nx4132)) ;
    aoi222 ix5800 (.Y (nx5138), .A0 (nx5137), .A1 (nx5125), .B0 (nx5239), .B1 (
           nx5137), .C0 (nx5130), .C1 (nx5125)) ;
    inv02 ix5801 (.Y (nx5139), .A (nx5138)) ;
    inv01 ix5802 (.Y (nx5140), .A (nx5959)) ;
    inv01 ix5803 (.Y (nx5141), .A (nx5959)) ;
    inv01 ix5804 (.Y (nx5142), .A (nx5959)) ;
    inv01 ix5805 (.Y (nx5143), .A (nx5149)) ;
    inv02 ix5806 (.Y (nx5144), .A (nx5149)) ;
    inv02 ix5807 (.Y (nx5145), .A (nx5149)) ;
    inv01 ix5808 (.Y (nx5146), .A (nx5149)) ;
    inv01 ix5809 (.Y (nx5147), .A (nx5149)) ;
    inv01 ix5810 (.Y (nx5148), .A (nx5149)) ;
    buf02 ix5811 (.Y (nx5149), .A (nx5180)) ;
    inv02 ix5812 (.Y (nx5150), .A (nx4174)) ;
    inv01 ix5813 (.Y (nx5151), .A (nx4414)) ;
    oai22 ix5814 (.Y (nx5152), .A0 (nx5150), .A1 (nx5151), .B0 (nx4174), .B1 (
          nx4414)) ;
    oai22 reg_nx2450 (.Y (nx2450), .A0 (nx5151), .A1 (nx4174), .B0 (nx5150), .B1 (
          nx4414)) ;
    ao22 reg_nx1786 (.Y (nx1786), .A0 (negative_M_16), .A1 (nx4476), .B0 (
         positive_M_16), .B1 (nx4466)) ;
    ao21 ix5815 (.Y (nx5153), .A0 (nx4708), .A1 (nx4667), .B0 (nx4668)) ;
    aoi321 reg_nx4116 (.Y (nx4116), .A0 (nx4666), .A1 (nx4911), .A2 (nx4667), .B0 (
           nx4666), .B1 (nx5153), .C0 (nx5207)) ;
    inv01 ix5816 (.Y (nx5154), .A (nx4116)) ;
    oai32 ix5817 (.Y (nx5155), .A0 (nx5207), .A1 (nx4668), .A2 (nx4667), .B0 (
          nx4666), .B1 (nx5207)) ;
    nor02_2x ix5818 (.Y (nx5156), .A0 (nx5233), .A1 (nx5227)) ;
    and04 ix5819 (.Y (nx5157), .A0 (nx5025), .A1 (nx5235), .A2 (nx2210), .A3 (
          nx5156)) ;
    inv01 ix5820 (.Y (nx5158), .A (nx4053)) ;
    inv02 ix5821 (.Y (nx5159), .A (nx2210)) ;
    and03 ix5822 (.Y (nx5160), .A0 (nx4635), .A1 (nx5159), .A2 (nx5156)) ;
    inv02 reg_nx4302 (.Y (nx4302), .A (nx5227)) ;
    and02 ix5823 (.Y (nx5161), .A0 (nx5025), .A1 (nx5235)) ;
    nand03_2x ix5824 (.Y (nx5162), .A0 (nx4635), .A1 (nx5159), .A2 (nx5156)) ;
    oai422 ix5825 (.Y (nx5163), .A0 (nx4635), .A1 (nx5159), .A2 (nx5233), .A3 (
           nx5227), .B0 (nx5229), .B1 (nx4090), .C0 (nx5161), .C1 (nx5162)) ;
    ao221 reg_nx3338 (.Y (nx3338), .A0 (nx4053), .A1 (nx5157), .B0 (nx5158), .B1 (
          nx5160), .C0 (nx5163)) ;
    inv02 reg_nx4452 (.Y (nx4452), .A (nx5233)) ;
    inv01 ix5826 (.Y (nx5164), .A (nx5125)) ;
    inv01 ix5827 (.Y (nx5165), .A (nx5130)) ;
    nand02_2x ix5828 (.Y (nx5166), .A0 (nx5125), .A1 (nx5239)) ;
    inv02 ix5829 (.Y (nx5167), .A (nx5137)) ;
    aoi22 ix5830 (.Y (nx5168), .A0 (nx5164), .A1 (nx5165), .B0 (nx5166), .B1 (
          nx5167)) ;
    nor02_2x ix5831 (.Y (nx5169), .A0 (nx5961), .A1 (nx4884)) ;
    aoi21 ix5832 (.Y (nx5170), .A0 (nx4623), .A1 (nx5961), .B0 (nx5124)) ;
    nor02_2x ix5833 (.Y (nx5171), .A0 (nx5169), .A1 (nx5170)) ;
    or02 ix5834 (.Y (nx5172), .A0 (nx5137), .A1 (nx5239)) ;
    aoi221 ix5835 (.Y (nx5173), .A0 (nx5125), .A1 (nx5172), .B0 (nx5130), .B1 (
           nx5137), .C0 (nx4884)) ;
    inv01 ix5836 (.Y (nx5174), .A (nx5173)) ;
    inv01 ix5837 (.Y (nx5175), .A (nx5173)) ;
    inv01 ix5838 (.Y (nx5176), .A (nx5173)) ;
    inv01 ix5839 (.Y (nx5177), .A (nx5173)) ;
    inv01 reg_nx2330 (.Y (nx2330), .A (nx5168)) ;
    inv01 ix5840 (.Y (nx5178), .A (nx5961)) ;
    inv01 ix5841 (.Y (nx5179), .A (nx5961)) ;
    inv01 ix5842 (.Y (nx5180), .A (nx5961)) ;
    ao22 reg_nx2086 (.Y (nx2086), .A0 (negative_M_21), .A1 (nx4478_XX0_XREP64), 
         .B0 (positive_M_21), .B1 (nx4468)) ;
    aoi221 reg_nx4056 (.Y (nx4056), .A0 (positive_M_22), .A1 (nx4282), .B0 (
           negative_M_22), .B1 (nx4270), .C0 (nx2086)) ;
    inv02 ix5843 (.Y (nx5181), .A (nx3912)) ;
    inv01 ix5844 (.Y (nx5182), .A (nx5911)) ;
    aoi22 ix5845 (.Y (nx5183), .A0 (nx5911), .A1 (nx5181), .B0 (nx3912), .B1 (
          nx5182)) ;
    inv01 reg_nx1730 (.Y (nx1730), .A (nx5218)) ;
    inv01 ix5846 (.Y (nx5184), .A (nx5219)) ;
    inv01 ix5847 (.Y (nx5185), .A (nx5219)) ;
    inv01 ix5848 (.Y (nx5186), .A (nx5219)) ;
    inv01 ix5849 (.Y (nx5187), .A (nx5219)) ;
    inv01 ix5850 (.Y (nx5188), .A (nx5219)) ;
    inv01 ix5851 (.Y (nx5189), .A (nx5219)) ;
    inv01 ix5852 (.Y (nx5190), .A (nx5062)) ;
    inv01 ix5853 (.Y (nx5191), .A (nx4820)) ;
    oai32 ix5854 (.Y (nx5192), .A0 (nx5190), .A1 (nx5191), .A2 (nx4746), .B0 (
          nx4747), .B1 (nx932)) ;
    inv02 ix5855 (.Y (nx5193), .A (nx4788)) ;
    ao22 ix5856 (.Y (nx5194), .A0 (nx4280), .A1 (positive_M_17), .B0 (nx4268), .B1 (
         negative_M_17)) ;
    aoi22 ix5857 (.Y (nx5195), .A0 (nx1786), .A1 (nx5193), .B0 (nx5194), .B1 (
          nx5193)) ;
    inv01 ix5858 (.Y (nx5196), .A (nx5195)) ;
    inv01 ix5859 (.Y (nx5197), .A (nx5195)) ;
    and02 ix5860 (.Y (nx5198), .A0 (nx4268), .A1 (negative_M_17)) ;
    and02 ix5861 (.Y (nx5199), .A0 (nx4280), .A1 (positive_M_17)) ;
    nor03_2x ix5862 (.Y (nx5200), .A0 (nx5198), .A1 (nx5199), .A2 (nx1786)) ;
    ao21 ix5863 (.Y (nx5201), .A0 (nx4673), .A1 (nx4674), .B0 (nx4672)) ;
    nor02_2x ix5864 (.Y (nx5202), .A0 (nx4671), .A1 (nx4920)) ;
    inv01 ix5865 (.Y (nx5203), .A (nx4657)) ;
    nor04_2x ix5866 (.Y (nx5204), .A0 (nx5202), .A1 (nx5203), .A2 (nx4708), .A3 (
             nx4668)) ;
    nand02_2x ix5867 (.Y (nx5205), .A0 (nx5201), .A1 (nx5204)) ;
    oai22 ix5868 (.Y (nx5206), .A0 (nx4672), .A1 (nx4673), .B0 (nx4672), .B1 (
          nx4674)) ;
    oai21 ix5869 (.Y (nx5207), .A0 (nx4671), .A1 (nx4920), .B0 (nx4657)) ;
    buf16 ix5870 (.Y (nx5208), .A (nx4332)) ;
    buf16 ix5871 (.Y (nx5209), .A (nx4332)) ;
    buf16 ix5872 (.Y (nx5210), .A (nx602)) ;
    buf16 ix5873 (.Y (nx5211), .A (nx602)) ;
    buf16 ix5874 (.Y (nx5212), .A (nx4758)) ;
    buf16 ix5875 (.Y (nx5213), .A (nx4758)) ;
    buf16 ix5876 (.Y (nx5214), .A (nx4954)) ;
    buf16 ix5877 (.Y (nx5215), .A (nx4954)) ;
    buf16 ix5878 (.Y (nx5216), .A (nx4995)) ;
    buf16 ix5879 (.Y (nx5217), .A (nx4995)) ;
    buf16 ix5880 (.Y (nx5218), .A (nx5183)) ;
    buf16 ix5881 (.Y (nx5219), .A (nx5183)) ;
    buf16 ix5882 (.Y (nx5220), .A (nx5923)) ;
    buf16 ix5883 (.Y (nx5221), .A (nx5923)) ;
    buf16 ix5884 (.Y (nx5222), .A (nx4396)) ;
    buf16 ix5885 (.Y (nx5223), .A (nx4396)) ;
    buf16 ix5886 (.Y (nx5224), .A (nx4398)) ;
    buf16 ix5887 (.Y (nx5225), .A (nx4398)) ;
    buf16 ix5888 (.Y (nx5226), .A (nx4286)) ;
    buf16 ix5889 (.Y (nx5227), .A (nx4286)) ;
    buf16 ix5890 (.Y (nx5228), .A (nx4302)) ;
    buf16 ix5891 (.Y (nx5229), .A (nx4302)) ;
    buf16 ix5892 (.Y (nx5230), .A (nx4400)) ;
    buf16 ix5893 (.Y (nx5231), .A (nx4400)) ;
    buf16 ix5894 (.Y (nx5232), .A (nx4486)) ;
    buf16 ix5895 (.Y (nx5233), .A (nx4486)) ;
    buf16 ix5896 (.Y (nx5234), .A (nx2090)) ;
    buf16 ix5897 (.Y (nx5235), .A (nx2090)) ;
    buf16 ix5898 (.Y (nx5236), .A (nx4119)) ;
    buf16 ix5899 (.Y (nx5237), .A (nx4119)) ;
    buf16 ix5900 (.Y (nx5238), .A (nx4410)) ;
    buf16 ix5901 (.Y (nx5239), .A (nx4410)) ;
    buf16 ix5902 (.Y (nx5240), .A (nx2390)) ;
    buf16 ix5903 (.Y (nx5241), .A (nx2390)) ;
    inv02 ix5904 (.Y (nx5905), .A (nx4725)) ;
    inv01 ix5906 (.Y (nx5907), .A (nx4742)) ;
    inv01 ix5908 (.Y (nx5909), .A (nx4746)) ;
    inv01 ix5910 (.Y (nx5911), .A (nx4699)) ;
    buf02 ix5912 (.Y (nx5913), .A (nx4602)) ;
    inv01 ix5914 (.Y (nx5915), .A (nx4691)) ;
    buf02 ix5916 (.Y (nx5917), .A (nx4710)) ;
    buf02 ix5918 (.Y (nx5919), .A (nx4731)) ;
    buf02 ix5920 (.Y (nx5921), .A (nx3696)) ;
    buf02 ix5922 (.Y (nx5923), .A (nx1850)) ;
    buf02 ix5924 (.Y (nx5925), .A (nx4801)) ;
    inv02 ix5926 (.Y (nx5927), .A (nx4877)) ;
    inv02 ix5928 (.Y (nx5929), .A (nx4877)) ;
    buf02 ix5930 (.Y (nx5931), .A (nx3972)) ;
    inv01 ix5932 (.Y (nx5933), .A (nx4922)) ;
    inv01 ix5934 (.Y (nx5935), .A (nx4733)) ;
    buf02 ix5936 (.Y (nx5937), .A (nx4968)) ;
    inv02 ix5938 (.Y (nx5939), .A (nx4837)) ;
    inv01 ix5940 (.Y (nx5941), .A (nx4630)) ;
    buf02 ix5942 (.Y (nx5943), .A (nx5001)) ;
    inv02 ix5944 (.Y (nx5945), .A (nx1026)) ;
    inv01 ix5946 (.Y (nx5947), .A (nx3699)) ;
    inv01 ix5948 (.Y (nx5949), .A (nx4696)) ;
    inv01 ix5950 (.Y (nx5951), .A (nx4695)) ;
    inv01 ix5952 (.Y (nx5953), .A (nx4734)) ;
    inv01 ix5954 (.Y (nx5955), .A (nx4776)) ;
    inv01 ix5956 (.Y (nx5957), .A (nx3752)) ;
    inv02 ix5958 (.Y (nx5959), .A (nx5139)) ;
    inv01 ix5960 (.Y (nx5961), .A (nx2330)) ;
    inv02 ix5970 (.Y (nx5971), .A (nx3851)) ;
    inv02 ix5972 (.Y (nx5973), .A (nx3823)) ;
    inv02 ix5974 (.Y (nx5975), .A (nx3823)) ;
    inv02 ix5976 (.Y (nx5977), .A (nx3795)) ;
    inv02 ix5978 (.Y (nx5979), .A (nx3795)) ;
    inv02 ix5980 (.Y (nx5981), .A (nx3739)) ;
    inv02 ix5982 (.Y (nx5983), .A (nx3739)) ;
    inv02 ix5984 (.Y (nx5985), .A (nx3711)) ;
    inv02 ix5986 (.Y (nx5987), .A (nx3711)) ;
    inv02 ix5988 (.Y (nx5989), .A (nx3683)) ;
    inv02 ix5990 (.Y (nx5991), .A (nx3655)) ;
    inv02 ix5992 (.Y (nx5993), .A (nx3627)) ;
    inv02 ix5994 (.Y (nx5995), .A (nx3597)) ;
    buf02 ix5996 (.Y (nx5997), .A (M[3])) ;
    buf02 ix5998 (.Y (nx5999), .A (M[2])) ;
    buf02 ix6000 (.Y (nx6001), .A (M[2])) ;
    inv02 ix6002 (.Y (nx6003), .A (nx4755)) ;
    inv02 ix6004 (.Y (nx6005), .A (nx4755)) ;
    buf02 ix6006 (.Y (nx6007), .A (M[0])) ;
    buf02 ix6008 (.Y (nx6009), .A (M[0])) ;
endmodule


module ReluLayer ( d_arr_0__31, d_arr_0__30, d_arr_0__29, d_arr_0__28, 
                   d_arr_0__27, d_arr_0__26, d_arr_0__25, d_arr_0__24, 
                   d_arr_0__23, d_arr_0__22, d_arr_0__21, d_arr_0__20, 
                   d_arr_0__19, d_arr_0__18, d_arr_0__17, d_arr_0__16, 
                   d_arr_0__15, d_arr_0__14, d_arr_0__13, d_arr_0__12, 
                   d_arr_0__11, d_arr_0__10, d_arr_0__9, d_arr_0__8, d_arr_0__7, 
                   d_arr_0__6, d_arr_0__5, d_arr_0__4, d_arr_0__3, d_arr_0__2, 
                   d_arr_0__1, d_arr_0__0, d_arr_1__31, d_arr_1__30, d_arr_1__29, 
                   d_arr_1__28, d_arr_1__27, d_arr_1__26, d_arr_1__25, 
                   d_arr_1__24, d_arr_1__23, d_arr_1__22, d_arr_1__21, 
                   d_arr_1__20, d_arr_1__19, d_arr_1__18, d_arr_1__17, 
                   d_arr_1__16, d_arr_1__15, d_arr_1__14, d_arr_1__13, 
                   d_arr_1__12, d_arr_1__11, d_arr_1__10, d_arr_1__9, d_arr_1__8, 
                   d_arr_1__7, d_arr_1__6, d_arr_1__5, d_arr_1__4, d_arr_1__3, 
                   d_arr_1__2, d_arr_1__1, d_arr_1__0, d_arr_2__31, d_arr_2__30, 
                   d_arr_2__29, d_arr_2__28, d_arr_2__27, d_arr_2__26, 
                   d_arr_2__25, d_arr_2__24, d_arr_2__23, d_arr_2__22, 
                   d_arr_2__21, d_arr_2__20, d_arr_2__19, d_arr_2__18, 
                   d_arr_2__17, d_arr_2__16, d_arr_2__15, d_arr_2__14, 
                   d_arr_2__13, d_arr_2__12, d_arr_2__11, d_arr_2__10, 
                   d_arr_2__9, d_arr_2__8, d_arr_2__7, d_arr_2__6, d_arr_2__5, 
                   d_arr_2__4, d_arr_2__3, d_arr_2__2, d_arr_2__1, d_arr_2__0, 
                   d_arr_3__31, d_arr_3__30, d_arr_3__29, d_arr_3__28, 
                   d_arr_3__27, d_arr_3__26, d_arr_3__25, d_arr_3__24, 
                   d_arr_3__23, d_arr_3__22, d_arr_3__21, d_arr_3__20, 
                   d_arr_3__19, d_arr_3__18, d_arr_3__17, d_arr_3__16, 
                   d_arr_3__15, d_arr_3__14, d_arr_3__13, d_arr_3__12, 
                   d_arr_3__11, d_arr_3__10, d_arr_3__9, d_arr_3__8, d_arr_3__7, 
                   d_arr_3__6, d_arr_3__5, d_arr_3__4, d_arr_3__3, d_arr_3__2, 
                   d_arr_3__1, d_arr_3__0, d_arr_4__31, d_arr_4__30, d_arr_4__29, 
                   d_arr_4__28, d_arr_4__27, d_arr_4__26, d_arr_4__25, 
                   d_arr_4__24, d_arr_4__23, d_arr_4__22, d_arr_4__21, 
                   d_arr_4__20, d_arr_4__19, d_arr_4__18, d_arr_4__17, 
                   d_arr_4__16, d_arr_4__15, d_arr_4__14, d_arr_4__13, 
                   d_arr_4__12, d_arr_4__11, d_arr_4__10, d_arr_4__9, d_arr_4__8, 
                   d_arr_4__7, d_arr_4__6, d_arr_4__5, d_arr_4__4, d_arr_4__3, 
                   d_arr_4__2, d_arr_4__1, d_arr_4__0, d_arr_5__31, d_arr_5__30, 
                   d_arr_5__29, d_arr_5__28, d_arr_5__27, d_arr_5__26, 
                   d_arr_5__25, d_arr_5__24, d_arr_5__23, d_arr_5__22, 
                   d_arr_5__21, d_arr_5__20, d_arr_5__19, d_arr_5__18, 
                   d_arr_5__17, d_arr_5__16, d_arr_5__15, d_arr_5__14, 
                   d_arr_5__13, d_arr_5__12, d_arr_5__11, d_arr_5__10, 
                   d_arr_5__9, d_arr_5__8, d_arr_5__7, d_arr_5__6, d_arr_5__5, 
                   d_arr_5__4, d_arr_5__3, d_arr_5__2, d_arr_5__1, d_arr_5__0, 
                   d_arr_6__31, d_arr_6__30, d_arr_6__29, d_arr_6__28, 
                   d_arr_6__27, d_arr_6__26, d_arr_6__25, d_arr_6__24, 
                   d_arr_6__23, d_arr_6__22, d_arr_6__21, d_arr_6__20, 
                   d_arr_6__19, d_arr_6__18, d_arr_6__17, d_arr_6__16, 
                   d_arr_6__15, d_arr_6__14, d_arr_6__13, d_arr_6__12, 
                   d_arr_6__11, d_arr_6__10, d_arr_6__9, d_arr_6__8, d_arr_6__7, 
                   d_arr_6__6, d_arr_6__5, d_arr_6__4, d_arr_6__3, d_arr_6__2, 
                   d_arr_6__1, d_arr_6__0, d_arr_7__31, d_arr_7__30, d_arr_7__29, 
                   d_arr_7__28, d_arr_7__27, d_arr_7__26, d_arr_7__25, 
                   d_arr_7__24, d_arr_7__23, d_arr_7__22, d_arr_7__21, 
                   d_arr_7__20, d_arr_7__19, d_arr_7__18, d_arr_7__17, 
                   d_arr_7__16, d_arr_7__15, d_arr_7__14, d_arr_7__13, 
                   d_arr_7__12, d_arr_7__11, d_arr_7__10, d_arr_7__9, d_arr_7__8, 
                   d_arr_7__7, d_arr_7__6, d_arr_7__5, d_arr_7__4, d_arr_7__3, 
                   d_arr_7__2, d_arr_7__1, d_arr_7__0, d_arr_8__31, d_arr_8__30, 
                   d_arr_8__29, d_arr_8__28, d_arr_8__27, d_arr_8__26, 
                   d_arr_8__25, d_arr_8__24, d_arr_8__23, d_arr_8__22, 
                   d_arr_8__21, d_arr_8__20, d_arr_8__19, d_arr_8__18, 
                   d_arr_8__17, d_arr_8__16, d_arr_8__15, d_arr_8__14, 
                   d_arr_8__13, d_arr_8__12, d_arr_8__11, d_arr_8__10, 
                   d_arr_8__9, d_arr_8__8, d_arr_8__7, d_arr_8__6, d_arr_8__5, 
                   d_arr_8__4, d_arr_8__3, d_arr_8__2, d_arr_8__1, d_arr_8__0, 
                   d_arr_9__31, d_arr_9__30, d_arr_9__29, d_arr_9__28, 
                   d_arr_9__27, d_arr_9__26, d_arr_9__25, d_arr_9__24, 
                   d_arr_9__23, d_arr_9__22, d_arr_9__21, d_arr_9__20, 
                   d_arr_9__19, d_arr_9__18, d_arr_9__17, d_arr_9__16, 
                   d_arr_9__15, d_arr_9__14, d_arr_9__13, d_arr_9__12, 
                   d_arr_9__11, d_arr_9__10, d_arr_9__9, d_arr_9__8, d_arr_9__7, 
                   d_arr_9__6, d_arr_9__5, d_arr_9__4, d_arr_9__3, d_arr_9__2, 
                   d_arr_9__1, d_arr_9__0, d_arr_10__31, d_arr_10__30, 
                   d_arr_10__29, d_arr_10__28, d_arr_10__27, d_arr_10__26, 
                   d_arr_10__25, d_arr_10__24, d_arr_10__23, d_arr_10__22, 
                   d_arr_10__21, d_arr_10__20, d_arr_10__19, d_arr_10__18, 
                   d_arr_10__17, d_arr_10__16, d_arr_10__15, d_arr_10__14, 
                   d_arr_10__13, d_arr_10__12, d_arr_10__11, d_arr_10__10, 
                   d_arr_10__9, d_arr_10__8, d_arr_10__7, d_arr_10__6, 
                   d_arr_10__5, d_arr_10__4, d_arr_10__3, d_arr_10__2, 
                   d_arr_10__1, d_arr_10__0, d_arr_11__31, d_arr_11__30, 
                   d_arr_11__29, d_arr_11__28, d_arr_11__27, d_arr_11__26, 
                   d_arr_11__25, d_arr_11__24, d_arr_11__23, d_arr_11__22, 
                   d_arr_11__21, d_arr_11__20, d_arr_11__19, d_arr_11__18, 
                   d_arr_11__17, d_arr_11__16, d_arr_11__15, d_arr_11__14, 
                   d_arr_11__13, d_arr_11__12, d_arr_11__11, d_arr_11__10, 
                   d_arr_11__9, d_arr_11__8, d_arr_11__7, d_arr_11__6, 
                   d_arr_11__5, d_arr_11__4, d_arr_11__3, d_arr_11__2, 
                   d_arr_11__1, d_arr_11__0, d_arr_12__31, d_arr_12__30, 
                   d_arr_12__29, d_arr_12__28, d_arr_12__27, d_arr_12__26, 
                   d_arr_12__25, d_arr_12__24, d_arr_12__23, d_arr_12__22, 
                   d_arr_12__21, d_arr_12__20, d_arr_12__19, d_arr_12__18, 
                   d_arr_12__17, d_arr_12__16, d_arr_12__15, d_arr_12__14, 
                   d_arr_12__13, d_arr_12__12, d_arr_12__11, d_arr_12__10, 
                   d_arr_12__9, d_arr_12__8, d_arr_12__7, d_arr_12__6, 
                   d_arr_12__5, d_arr_12__4, d_arr_12__3, d_arr_12__2, 
                   d_arr_12__1, d_arr_12__0, d_arr_13__31, d_arr_13__30, 
                   d_arr_13__29, d_arr_13__28, d_arr_13__27, d_arr_13__26, 
                   d_arr_13__25, d_arr_13__24, d_arr_13__23, d_arr_13__22, 
                   d_arr_13__21, d_arr_13__20, d_arr_13__19, d_arr_13__18, 
                   d_arr_13__17, d_arr_13__16, d_arr_13__15, d_arr_13__14, 
                   d_arr_13__13, d_arr_13__12, d_arr_13__11, d_arr_13__10, 
                   d_arr_13__9, d_arr_13__8, d_arr_13__7, d_arr_13__6, 
                   d_arr_13__5, d_arr_13__4, d_arr_13__3, d_arr_13__2, 
                   d_arr_13__1, d_arr_13__0, d_arr_14__31, d_arr_14__30, 
                   d_arr_14__29, d_arr_14__28, d_arr_14__27, d_arr_14__26, 
                   d_arr_14__25, d_arr_14__24, d_arr_14__23, d_arr_14__22, 
                   d_arr_14__21, d_arr_14__20, d_arr_14__19, d_arr_14__18, 
                   d_arr_14__17, d_arr_14__16, d_arr_14__15, d_arr_14__14, 
                   d_arr_14__13, d_arr_14__12, d_arr_14__11, d_arr_14__10, 
                   d_arr_14__9, d_arr_14__8, d_arr_14__7, d_arr_14__6, 
                   d_arr_14__5, d_arr_14__4, d_arr_14__3, d_arr_14__2, 
                   d_arr_14__1, d_arr_14__0, d_arr_15__31, d_arr_15__30, 
                   d_arr_15__29, d_arr_15__28, d_arr_15__27, d_arr_15__26, 
                   d_arr_15__25, d_arr_15__24, d_arr_15__23, d_arr_15__22, 
                   d_arr_15__21, d_arr_15__20, d_arr_15__19, d_arr_15__18, 
                   d_arr_15__17, d_arr_15__16, d_arr_15__15, d_arr_15__14, 
                   d_arr_15__13, d_arr_15__12, d_arr_15__11, d_arr_15__10, 
                   d_arr_15__9, d_arr_15__8, d_arr_15__7, d_arr_15__6, 
                   d_arr_15__5, d_arr_15__4, d_arr_15__3, d_arr_15__2, 
                   d_arr_15__1, d_arr_15__0, d_arr_16__31, d_arr_16__30, 
                   d_arr_16__29, d_arr_16__28, d_arr_16__27, d_arr_16__26, 
                   d_arr_16__25, d_arr_16__24, d_arr_16__23, d_arr_16__22, 
                   d_arr_16__21, d_arr_16__20, d_arr_16__19, d_arr_16__18, 
                   d_arr_16__17, d_arr_16__16, d_arr_16__15, d_arr_16__14, 
                   d_arr_16__13, d_arr_16__12, d_arr_16__11, d_arr_16__10, 
                   d_arr_16__9, d_arr_16__8, d_arr_16__7, d_arr_16__6, 
                   d_arr_16__5, d_arr_16__4, d_arr_16__3, d_arr_16__2, 
                   d_arr_16__1, d_arr_16__0, d_arr_17__31, d_arr_17__30, 
                   d_arr_17__29, d_arr_17__28, d_arr_17__27, d_arr_17__26, 
                   d_arr_17__25, d_arr_17__24, d_arr_17__23, d_arr_17__22, 
                   d_arr_17__21, d_arr_17__20, d_arr_17__19, d_arr_17__18, 
                   d_arr_17__17, d_arr_17__16, d_arr_17__15, d_arr_17__14, 
                   d_arr_17__13, d_arr_17__12, d_arr_17__11, d_arr_17__10, 
                   d_arr_17__9, d_arr_17__8, d_arr_17__7, d_arr_17__6, 
                   d_arr_17__5, d_arr_17__4, d_arr_17__3, d_arr_17__2, 
                   d_arr_17__1, d_arr_17__0, d_arr_18__31, d_arr_18__30, 
                   d_arr_18__29, d_arr_18__28, d_arr_18__27, d_arr_18__26, 
                   d_arr_18__25, d_arr_18__24, d_arr_18__23, d_arr_18__22, 
                   d_arr_18__21, d_arr_18__20, d_arr_18__19, d_arr_18__18, 
                   d_arr_18__17, d_arr_18__16, d_arr_18__15, d_arr_18__14, 
                   d_arr_18__13, d_arr_18__12, d_arr_18__11, d_arr_18__10, 
                   d_arr_18__9, d_arr_18__8, d_arr_18__7, d_arr_18__6, 
                   d_arr_18__5, d_arr_18__4, d_arr_18__3, d_arr_18__2, 
                   d_arr_18__1, d_arr_18__0, d_arr_19__31, d_arr_19__30, 
                   d_arr_19__29, d_arr_19__28, d_arr_19__27, d_arr_19__26, 
                   d_arr_19__25, d_arr_19__24, d_arr_19__23, d_arr_19__22, 
                   d_arr_19__21, d_arr_19__20, d_arr_19__19, d_arr_19__18, 
                   d_arr_19__17, d_arr_19__16, d_arr_19__15, d_arr_19__14, 
                   d_arr_19__13, d_arr_19__12, d_arr_19__11, d_arr_19__10, 
                   d_arr_19__9, d_arr_19__8, d_arr_19__7, d_arr_19__6, 
                   d_arr_19__5, d_arr_19__4, d_arr_19__3, d_arr_19__2, 
                   d_arr_19__1, d_arr_19__0, d_arr_20__31, d_arr_20__30, 
                   d_arr_20__29, d_arr_20__28, d_arr_20__27, d_arr_20__26, 
                   d_arr_20__25, d_arr_20__24, d_arr_20__23, d_arr_20__22, 
                   d_arr_20__21, d_arr_20__20, d_arr_20__19, d_arr_20__18, 
                   d_arr_20__17, d_arr_20__16, d_arr_20__15, d_arr_20__14, 
                   d_arr_20__13, d_arr_20__12, d_arr_20__11, d_arr_20__10, 
                   d_arr_20__9, d_arr_20__8, d_arr_20__7, d_arr_20__6, 
                   d_arr_20__5, d_arr_20__4, d_arr_20__3, d_arr_20__2, 
                   d_arr_20__1, d_arr_20__0, d_arr_21__31, d_arr_21__30, 
                   d_arr_21__29, d_arr_21__28, d_arr_21__27, d_arr_21__26, 
                   d_arr_21__25, d_arr_21__24, d_arr_21__23, d_arr_21__22, 
                   d_arr_21__21, d_arr_21__20, d_arr_21__19, d_arr_21__18, 
                   d_arr_21__17, d_arr_21__16, d_arr_21__15, d_arr_21__14, 
                   d_arr_21__13, d_arr_21__12, d_arr_21__11, d_arr_21__10, 
                   d_arr_21__9, d_arr_21__8, d_arr_21__7, d_arr_21__6, 
                   d_arr_21__5, d_arr_21__4, d_arr_21__3, d_arr_21__2, 
                   d_arr_21__1, d_arr_21__0, d_arr_22__31, d_arr_22__30, 
                   d_arr_22__29, d_arr_22__28, d_arr_22__27, d_arr_22__26, 
                   d_arr_22__25, d_arr_22__24, d_arr_22__23, d_arr_22__22, 
                   d_arr_22__21, d_arr_22__20, d_arr_22__19, d_arr_22__18, 
                   d_arr_22__17, d_arr_22__16, d_arr_22__15, d_arr_22__14, 
                   d_arr_22__13, d_arr_22__12, d_arr_22__11, d_arr_22__10, 
                   d_arr_22__9, d_arr_22__8, d_arr_22__7, d_arr_22__6, 
                   d_arr_22__5, d_arr_22__4, d_arr_22__3, d_arr_22__2, 
                   d_arr_22__1, d_arr_22__0, d_arr_23__31, d_arr_23__30, 
                   d_arr_23__29, d_arr_23__28, d_arr_23__27, d_arr_23__26, 
                   d_arr_23__25, d_arr_23__24, d_arr_23__23, d_arr_23__22, 
                   d_arr_23__21, d_arr_23__20, d_arr_23__19, d_arr_23__18, 
                   d_arr_23__17, d_arr_23__16, d_arr_23__15, d_arr_23__14, 
                   d_arr_23__13, d_arr_23__12, d_arr_23__11, d_arr_23__10, 
                   d_arr_23__9, d_arr_23__8, d_arr_23__7, d_arr_23__6, 
                   d_arr_23__5, d_arr_23__4, d_arr_23__3, d_arr_23__2, 
                   d_arr_23__1, d_arr_23__0, d_arr_24__31, d_arr_24__30, 
                   d_arr_24__29, d_arr_24__28, d_arr_24__27, d_arr_24__26, 
                   d_arr_24__25, d_arr_24__24, d_arr_24__23, d_arr_24__22, 
                   d_arr_24__21, d_arr_24__20, d_arr_24__19, d_arr_24__18, 
                   d_arr_24__17, d_arr_24__16, d_arr_24__15, d_arr_24__14, 
                   d_arr_24__13, d_arr_24__12, d_arr_24__11, d_arr_24__10, 
                   d_arr_24__9, d_arr_24__8, d_arr_24__7, d_arr_24__6, 
                   d_arr_24__5, d_arr_24__4, d_arr_24__3, d_arr_24__2, 
                   d_arr_24__1, d_arr_24__0, q_arr_0__31, q_arr_0__30, 
                   q_arr_0__29, q_arr_0__28, q_arr_0__27, q_arr_0__26, 
                   q_arr_0__25, q_arr_0__24, q_arr_0__23, q_arr_0__22, 
                   q_arr_0__21, q_arr_0__20, q_arr_0__19, q_arr_0__18, 
                   q_arr_0__17, q_arr_0__16, q_arr_0__15, q_arr_0__14, 
                   q_arr_0__13, q_arr_0__12, q_arr_0__11, q_arr_0__10, 
                   q_arr_0__9, q_arr_0__8, q_arr_0__7, q_arr_0__6, q_arr_0__5, 
                   q_arr_0__4, q_arr_0__3, q_arr_0__2, q_arr_0__1, q_arr_0__0, 
                   q_arr_1__31, q_arr_1__30, q_arr_1__29, q_arr_1__28, 
                   q_arr_1__27, q_arr_1__26, q_arr_1__25, q_arr_1__24, 
                   q_arr_1__23, q_arr_1__22, q_arr_1__21, q_arr_1__20, 
                   q_arr_1__19, q_arr_1__18, q_arr_1__17, q_arr_1__16, 
                   q_arr_1__15, q_arr_1__14, q_arr_1__13, q_arr_1__12, 
                   q_arr_1__11, q_arr_1__10, q_arr_1__9, q_arr_1__8, q_arr_1__7, 
                   q_arr_1__6, q_arr_1__5, q_arr_1__4, q_arr_1__3, q_arr_1__2, 
                   q_arr_1__1, q_arr_1__0, q_arr_2__31, q_arr_2__30, q_arr_2__29, 
                   q_arr_2__28, q_arr_2__27, q_arr_2__26, q_arr_2__25, 
                   q_arr_2__24, q_arr_2__23, q_arr_2__22, q_arr_2__21, 
                   q_arr_2__20, q_arr_2__19, q_arr_2__18, q_arr_2__17, 
                   q_arr_2__16, q_arr_2__15, q_arr_2__14, q_arr_2__13, 
                   q_arr_2__12, q_arr_2__11, q_arr_2__10, q_arr_2__9, q_arr_2__8, 
                   q_arr_2__7, q_arr_2__6, q_arr_2__5, q_arr_2__4, q_arr_2__3, 
                   q_arr_2__2, q_arr_2__1, q_arr_2__0, q_arr_3__31, q_arr_3__30, 
                   q_arr_3__29, q_arr_3__28, q_arr_3__27, q_arr_3__26, 
                   q_arr_3__25, q_arr_3__24, q_arr_3__23, q_arr_3__22, 
                   q_arr_3__21, q_arr_3__20, q_arr_3__19, q_arr_3__18, 
                   q_arr_3__17, q_arr_3__16, q_arr_3__15, q_arr_3__14, 
                   q_arr_3__13, q_arr_3__12, q_arr_3__11, q_arr_3__10, 
                   q_arr_3__9, q_arr_3__8, q_arr_3__7, q_arr_3__6, q_arr_3__5, 
                   q_arr_3__4, q_arr_3__3, q_arr_3__2, q_arr_3__1, q_arr_3__0, 
                   q_arr_4__31, q_arr_4__30, q_arr_4__29, q_arr_4__28, 
                   q_arr_4__27, q_arr_4__26, q_arr_4__25, q_arr_4__24, 
                   q_arr_4__23, q_arr_4__22, q_arr_4__21, q_arr_4__20, 
                   q_arr_4__19, q_arr_4__18, q_arr_4__17, q_arr_4__16, 
                   q_arr_4__15, q_arr_4__14, q_arr_4__13, q_arr_4__12, 
                   q_arr_4__11, q_arr_4__10, q_arr_4__9, q_arr_4__8, q_arr_4__7, 
                   q_arr_4__6, q_arr_4__5, q_arr_4__4, q_arr_4__3, q_arr_4__2, 
                   q_arr_4__1, q_arr_4__0, q_arr_5__31, q_arr_5__30, q_arr_5__29, 
                   q_arr_5__28, q_arr_5__27, q_arr_5__26, q_arr_5__25, 
                   q_arr_5__24, q_arr_5__23, q_arr_5__22, q_arr_5__21, 
                   q_arr_5__20, q_arr_5__19, q_arr_5__18, q_arr_5__17, 
                   q_arr_5__16, q_arr_5__15, q_arr_5__14, q_arr_5__13, 
                   q_arr_5__12, q_arr_5__11, q_arr_5__10, q_arr_5__9, q_arr_5__8, 
                   q_arr_5__7, q_arr_5__6, q_arr_5__5, q_arr_5__4, q_arr_5__3, 
                   q_arr_5__2, q_arr_5__1, q_arr_5__0, q_arr_6__31, q_arr_6__30, 
                   q_arr_6__29, q_arr_6__28, q_arr_6__27, q_arr_6__26, 
                   q_arr_6__25, q_arr_6__24, q_arr_6__23, q_arr_6__22, 
                   q_arr_6__21, q_arr_6__20, q_arr_6__19, q_arr_6__18, 
                   q_arr_6__17, q_arr_6__16, q_arr_6__15, q_arr_6__14, 
                   q_arr_6__13, q_arr_6__12, q_arr_6__11, q_arr_6__10, 
                   q_arr_6__9, q_arr_6__8, q_arr_6__7, q_arr_6__6, q_arr_6__5, 
                   q_arr_6__4, q_arr_6__3, q_arr_6__2, q_arr_6__1, q_arr_6__0, 
                   q_arr_7__31, q_arr_7__30, q_arr_7__29, q_arr_7__28, 
                   q_arr_7__27, q_arr_7__26, q_arr_7__25, q_arr_7__24, 
                   q_arr_7__23, q_arr_7__22, q_arr_7__21, q_arr_7__20, 
                   q_arr_7__19, q_arr_7__18, q_arr_7__17, q_arr_7__16, 
                   q_arr_7__15, q_arr_7__14, q_arr_7__13, q_arr_7__12, 
                   q_arr_7__11, q_arr_7__10, q_arr_7__9, q_arr_7__8, q_arr_7__7, 
                   q_arr_7__6, q_arr_7__5, q_arr_7__4, q_arr_7__3, q_arr_7__2, 
                   q_arr_7__1, q_arr_7__0, q_arr_8__31, q_arr_8__30, q_arr_8__29, 
                   q_arr_8__28, q_arr_8__27, q_arr_8__26, q_arr_8__25, 
                   q_arr_8__24, q_arr_8__23, q_arr_8__22, q_arr_8__21, 
                   q_arr_8__20, q_arr_8__19, q_arr_8__18, q_arr_8__17, 
                   q_arr_8__16, q_arr_8__15, q_arr_8__14, q_arr_8__13, 
                   q_arr_8__12, q_arr_8__11, q_arr_8__10, q_arr_8__9, q_arr_8__8, 
                   q_arr_8__7, q_arr_8__6, q_arr_8__5, q_arr_8__4, q_arr_8__3, 
                   q_arr_8__2, q_arr_8__1, q_arr_8__0, q_arr_9__31, q_arr_9__30, 
                   q_arr_9__29, q_arr_9__28, q_arr_9__27, q_arr_9__26, 
                   q_arr_9__25, q_arr_9__24, q_arr_9__23, q_arr_9__22, 
                   q_arr_9__21, q_arr_9__20, q_arr_9__19, q_arr_9__18, 
                   q_arr_9__17, q_arr_9__16, q_arr_9__15, q_arr_9__14, 
                   q_arr_9__13, q_arr_9__12, q_arr_9__11, q_arr_9__10, 
                   q_arr_9__9, q_arr_9__8, q_arr_9__7, q_arr_9__6, q_arr_9__5, 
                   q_arr_9__4, q_arr_9__3, q_arr_9__2, q_arr_9__1, q_arr_9__0, 
                   q_arr_10__31, q_arr_10__30, q_arr_10__29, q_arr_10__28, 
                   q_arr_10__27, q_arr_10__26, q_arr_10__25, q_arr_10__24, 
                   q_arr_10__23, q_arr_10__22, q_arr_10__21, q_arr_10__20, 
                   q_arr_10__19, q_arr_10__18, q_arr_10__17, q_arr_10__16, 
                   q_arr_10__15, q_arr_10__14, q_arr_10__13, q_arr_10__12, 
                   q_arr_10__11, q_arr_10__10, q_arr_10__9, q_arr_10__8, 
                   q_arr_10__7, q_arr_10__6, q_arr_10__5, q_arr_10__4, 
                   q_arr_10__3, q_arr_10__2, q_arr_10__1, q_arr_10__0, 
                   q_arr_11__31, q_arr_11__30, q_arr_11__29, q_arr_11__28, 
                   q_arr_11__27, q_arr_11__26, q_arr_11__25, q_arr_11__24, 
                   q_arr_11__23, q_arr_11__22, q_arr_11__21, q_arr_11__20, 
                   q_arr_11__19, q_arr_11__18, q_arr_11__17, q_arr_11__16, 
                   q_arr_11__15, q_arr_11__14, q_arr_11__13, q_arr_11__12, 
                   q_arr_11__11, q_arr_11__10, q_arr_11__9, q_arr_11__8, 
                   q_arr_11__7, q_arr_11__6, q_arr_11__5, q_arr_11__4, 
                   q_arr_11__3, q_arr_11__2, q_arr_11__1, q_arr_11__0, 
                   q_arr_12__31, q_arr_12__30, q_arr_12__29, q_arr_12__28, 
                   q_arr_12__27, q_arr_12__26, q_arr_12__25, q_arr_12__24, 
                   q_arr_12__23, q_arr_12__22, q_arr_12__21, q_arr_12__20, 
                   q_arr_12__19, q_arr_12__18, q_arr_12__17, q_arr_12__16, 
                   q_arr_12__15, q_arr_12__14, q_arr_12__13, q_arr_12__12, 
                   q_arr_12__11, q_arr_12__10, q_arr_12__9, q_arr_12__8, 
                   q_arr_12__7, q_arr_12__6, q_arr_12__5, q_arr_12__4, 
                   q_arr_12__3, q_arr_12__2, q_arr_12__1, q_arr_12__0, 
                   q_arr_13__31, q_arr_13__30, q_arr_13__29, q_arr_13__28, 
                   q_arr_13__27, q_arr_13__26, q_arr_13__25, q_arr_13__24, 
                   q_arr_13__23, q_arr_13__22, q_arr_13__21, q_arr_13__20, 
                   q_arr_13__19, q_arr_13__18, q_arr_13__17, q_arr_13__16, 
                   q_arr_13__15, q_arr_13__14, q_arr_13__13, q_arr_13__12, 
                   q_arr_13__11, q_arr_13__10, q_arr_13__9, q_arr_13__8, 
                   q_arr_13__7, q_arr_13__6, q_arr_13__5, q_arr_13__4, 
                   q_arr_13__3, q_arr_13__2, q_arr_13__1, q_arr_13__0, 
                   q_arr_14__31, q_arr_14__30, q_arr_14__29, q_arr_14__28, 
                   q_arr_14__27, q_arr_14__26, q_arr_14__25, q_arr_14__24, 
                   q_arr_14__23, q_arr_14__22, q_arr_14__21, q_arr_14__20, 
                   q_arr_14__19, q_arr_14__18, q_arr_14__17, q_arr_14__16, 
                   q_arr_14__15, q_arr_14__14, q_arr_14__13, q_arr_14__12, 
                   q_arr_14__11, q_arr_14__10, q_arr_14__9, q_arr_14__8, 
                   q_arr_14__7, q_arr_14__6, q_arr_14__5, q_arr_14__4, 
                   q_arr_14__3, q_arr_14__2, q_arr_14__1, q_arr_14__0, 
                   q_arr_15__31, q_arr_15__30, q_arr_15__29, q_arr_15__28, 
                   q_arr_15__27, q_arr_15__26, q_arr_15__25, q_arr_15__24, 
                   q_arr_15__23, q_arr_15__22, q_arr_15__21, q_arr_15__20, 
                   q_arr_15__19, q_arr_15__18, q_arr_15__17, q_arr_15__16, 
                   q_arr_15__15, q_arr_15__14, q_arr_15__13, q_arr_15__12, 
                   q_arr_15__11, q_arr_15__10, q_arr_15__9, q_arr_15__8, 
                   q_arr_15__7, q_arr_15__6, q_arr_15__5, q_arr_15__4, 
                   q_arr_15__3, q_arr_15__2, q_arr_15__1, q_arr_15__0, 
                   q_arr_16__31, q_arr_16__30, q_arr_16__29, q_arr_16__28, 
                   q_arr_16__27, q_arr_16__26, q_arr_16__25, q_arr_16__24, 
                   q_arr_16__23, q_arr_16__22, q_arr_16__21, q_arr_16__20, 
                   q_arr_16__19, q_arr_16__18, q_arr_16__17, q_arr_16__16, 
                   q_arr_16__15, q_arr_16__14, q_arr_16__13, q_arr_16__12, 
                   q_arr_16__11, q_arr_16__10, q_arr_16__9, q_arr_16__8, 
                   q_arr_16__7, q_arr_16__6, q_arr_16__5, q_arr_16__4, 
                   q_arr_16__3, q_arr_16__2, q_arr_16__1, q_arr_16__0, 
                   q_arr_17__31, q_arr_17__30, q_arr_17__29, q_arr_17__28, 
                   q_arr_17__27, q_arr_17__26, q_arr_17__25, q_arr_17__24, 
                   q_arr_17__23, q_arr_17__22, q_arr_17__21, q_arr_17__20, 
                   q_arr_17__19, q_arr_17__18, q_arr_17__17, q_arr_17__16, 
                   q_arr_17__15, q_arr_17__14, q_arr_17__13, q_arr_17__12, 
                   q_arr_17__11, q_arr_17__10, q_arr_17__9, q_arr_17__8, 
                   q_arr_17__7, q_arr_17__6, q_arr_17__5, q_arr_17__4, 
                   q_arr_17__3, q_arr_17__2, q_arr_17__1, q_arr_17__0, 
                   q_arr_18__31, q_arr_18__30, q_arr_18__29, q_arr_18__28, 
                   q_arr_18__27, q_arr_18__26, q_arr_18__25, q_arr_18__24, 
                   q_arr_18__23, q_arr_18__22, q_arr_18__21, q_arr_18__20, 
                   q_arr_18__19, q_arr_18__18, q_arr_18__17, q_arr_18__16, 
                   q_arr_18__15, q_arr_18__14, q_arr_18__13, q_arr_18__12, 
                   q_arr_18__11, q_arr_18__10, q_arr_18__9, q_arr_18__8, 
                   q_arr_18__7, q_arr_18__6, q_arr_18__5, q_arr_18__4, 
                   q_arr_18__3, q_arr_18__2, q_arr_18__1, q_arr_18__0, 
                   q_arr_19__31, q_arr_19__30, q_arr_19__29, q_arr_19__28, 
                   q_arr_19__27, q_arr_19__26, q_arr_19__25, q_arr_19__24, 
                   q_arr_19__23, q_arr_19__22, q_arr_19__21, q_arr_19__20, 
                   q_arr_19__19, q_arr_19__18, q_arr_19__17, q_arr_19__16, 
                   q_arr_19__15, q_arr_19__14, q_arr_19__13, q_arr_19__12, 
                   q_arr_19__11, q_arr_19__10, q_arr_19__9, q_arr_19__8, 
                   q_arr_19__7, q_arr_19__6, q_arr_19__5, q_arr_19__4, 
                   q_arr_19__3, q_arr_19__2, q_arr_19__1, q_arr_19__0, 
                   q_arr_20__31, q_arr_20__30, q_arr_20__29, q_arr_20__28, 
                   q_arr_20__27, q_arr_20__26, q_arr_20__25, q_arr_20__24, 
                   q_arr_20__23, q_arr_20__22, q_arr_20__21, q_arr_20__20, 
                   q_arr_20__19, q_arr_20__18, q_arr_20__17, q_arr_20__16, 
                   q_arr_20__15, q_arr_20__14, q_arr_20__13, q_arr_20__12, 
                   q_arr_20__11, q_arr_20__10, q_arr_20__9, q_arr_20__8, 
                   q_arr_20__7, q_arr_20__6, q_arr_20__5, q_arr_20__4, 
                   q_arr_20__3, q_arr_20__2, q_arr_20__1, q_arr_20__0, 
                   q_arr_21__31, q_arr_21__30, q_arr_21__29, q_arr_21__28, 
                   q_arr_21__27, q_arr_21__26, q_arr_21__25, q_arr_21__24, 
                   q_arr_21__23, q_arr_21__22, q_arr_21__21, q_arr_21__20, 
                   q_arr_21__19, q_arr_21__18, q_arr_21__17, q_arr_21__16, 
                   q_arr_21__15, q_arr_21__14, q_arr_21__13, q_arr_21__12, 
                   q_arr_21__11, q_arr_21__10, q_arr_21__9, q_arr_21__8, 
                   q_arr_21__7, q_arr_21__6, q_arr_21__5, q_arr_21__4, 
                   q_arr_21__3, q_arr_21__2, q_arr_21__1, q_arr_21__0, 
                   q_arr_22__31, q_arr_22__30, q_arr_22__29, q_arr_22__28, 
                   q_arr_22__27, q_arr_22__26, q_arr_22__25, q_arr_22__24, 
                   q_arr_22__23, q_arr_22__22, q_arr_22__21, q_arr_22__20, 
                   q_arr_22__19, q_arr_22__18, q_arr_22__17, q_arr_22__16, 
                   q_arr_22__15, q_arr_22__14, q_arr_22__13, q_arr_22__12, 
                   q_arr_22__11, q_arr_22__10, q_arr_22__9, q_arr_22__8, 
                   q_arr_22__7, q_arr_22__6, q_arr_22__5, q_arr_22__4, 
                   q_arr_22__3, q_arr_22__2, q_arr_22__1, q_arr_22__0, 
                   q_arr_23__31, q_arr_23__30, q_arr_23__29, q_arr_23__28, 
                   q_arr_23__27, q_arr_23__26, q_arr_23__25, q_arr_23__24, 
                   q_arr_23__23, q_arr_23__22, q_arr_23__21, q_arr_23__20, 
                   q_arr_23__19, q_arr_23__18, q_arr_23__17, q_arr_23__16, 
                   q_arr_23__15, q_arr_23__14, q_arr_23__13, q_arr_23__12, 
                   q_arr_23__11, q_arr_23__10, q_arr_23__9, q_arr_23__8, 
                   q_arr_23__7, q_arr_23__6, q_arr_23__5, q_arr_23__4, 
                   q_arr_23__3, q_arr_23__2, q_arr_23__1, q_arr_23__0, 
                   q_arr_24__31, q_arr_24__30, q_arr_24__29, q_arr_24__28, 
                   q_arr_24__27, q_arr_24__26, q_arr_24__25, q_arr_24__24, 
                   q_arr_24__23, q_arr_24__22, q_arr_24__21, q_arr_24__20, 
                   q_arr_24__19, q_arr_24__18, q_arr_24__17, q_arr_24__16, 
                   q_arr_24__15, q_arr_24__14, q_arr_24__13, q_arr_24__12, 
                   q_arr_24__11, q_arr_24__10, q_arr_24__9, q_arr_24__8, 
                   q_arr_24__7, q_arr_24__6, q_arr_24__5, q_arr_24__4, 
                   q_arr_24__3, q_arr_24__2, q_arr_24__1, q_arr_24__0 ) ;

    output d_arr_0__31 ;
    output d_arr_0__30 ;
    output d_arr_0__29 ;
    output d_arr_0__28 ;
    output d_arr_0__27 ;
    output d_arr_0__26 ;
    output d_arr_0__25 ;
    output d_arr_0__24 ;
    output d_arr_0__23 ;
    output d_arr_0__22 ;
    output d_arr_0__21 ;
    output d_arr_0__20 ;
    output d_arr_0__19 ;
    output d_arr_0__18 ;
    output d_arr_0__17 ;
    output d_arr_0__16 ;
    output d_arr_0__15 ;
    output d_arr_0__14 ;
    output d_arr_0__13 ;
    output d_arr_0__12 ;
    output d_arr_0__11 ;
    output d_arr_0__10 ;
    output d_arr_0__9 ;
    output d_arr_0__8 ;
    output d_arr_0__7 ;
    output d_arr_0__6 ;
    output d_arr_0__5 ;
    output d_arr_0__4 ;
    output d_arr_0__3 ;
    output d_arr_0__2 ;
    output d_arr_0__1 ;
    output d_arr_0__0 ;
    output d_arr_1__31 ;
    output d_arr_1__30 ;
    output d_arr_1__29 ;
    output d_arr_1__28 ;
    output d_arr_1__27 ;
    output d_arr_1__26 ;
    output d_arr_1__25 ;
    output d_arr_1__24 ;
    output d_arr_1__23 ;
    output d_arr_1__22 ;
    output d_arr_1__21 ;
    output d_arr_1__20 ;
    output d_arr_1__19 ;
    output d_arr_1__18 ;
    output d_arr_1__17 ;
    output d_arr_1__16 ;
    output d_arr_1__15 ;
    output d_arr_1__14 ;
    output d_arr_1__13 ;
    output d_arr_1__12 ;
    output d_arr_1__11 ;
    output d_arr_1__10 ;
    output d_arr_1__9 ;
    output d_arr_1__8 ;
    output d_arr_1__7 ;
    output d_arr_1__6 ;
    output d_arr_1__5 ;
    output d_arr_1__4 ;
    output d_arr_1__3 ;
    output d_arr_1__2 ;
    output d_arr_1__1 ;
    output d_arr_1__0 ;
    output d_arr_2__31 ;
    output d_arr_2__30 ;
    output d_arr_2__29 ;
    output d_arr_2__28 ;
    output d_arr_2__27 ;
    output d_arr_2__26 ;
    output d_arr_2__25 ;
    output d_arr_2__24 ;
    output d_arr_2__23 ;
    output d_arr_2__22 ;
    output d_arr_2__21 ;
    output d_arr_2__20 ;
    output d_arr_2__19 ;
    output d_arr_2__18 ;
    output d_arr_2__17 ;
    output d_arr_2__16 ;
    output d_arr_2__15 ;
    output d_arr_2__14 ;
    output d_arr_2__13 ;
    output d_arr_2__12 ;
    output d_arr_2__11 ;
    output d_arr_2__10 ;
    output d_arr_2__9 ;
    output d_arr_2__8 ;
    output d_arr_2__7 ;
    output d_arr_2__6 ;
    output d_arr_2__5 ;
    output d_arr_2__4 ;
    output d_arr_2__3 ;
    output d_arr_2__2 ;
    output d_arr_2__1 ;
    output d_arr_2__0 ;
    output d_arr_3__31 ;
    output d_arr_3__30 ;
    output d_arr_3__29 ;
    output d_arr_3__28 ;
    output d_arr_3__27 ;
    output d_arr_3__26 ;
    output d_arr_3__25 ;
    output d_arr_3__24 ;
    output d_arr_3__23 ;
    output d_arr_3__22 ;
    output d_arr_3__21 ;
    output d_arr_3__20 ;
    output d_arr_3__19 ;
    output d_arr_3__18 ;
    output d_arr_3__17 ;
    output d_arr_3__16 ;
    output d_arr_3__15 ;
    output d_arr_3__14 ;
    output d_arr_3__13 ;
    output d_arr_3__12 ;
    output d_arr_3__11 ;
    output d_arr_3__10 ;
    output d_arr_3__9 ;
    output d_arr_3__8 ;
    output d_arr_3__7 ;
    output d_arr_3__6 ;
    output d_arr_3__5 ;
    output d_arr_3__4 ;
    output d_arr_3__3 ;
    output d_arr_3__2 ;
    output d_arr_3__1 ;
    output d_arr_3__0 ;
    output d_arr_4__31 ;
    output d_arr_4__30 ;
    output d_arr_4__29 ;
    output d_arr_4__28 ;
    output d_arr_4__27 ;
    output d_arr_4__26 ;
    output d_arr_4__25 ;
    output d_arr_4__24 ;
    output d_arr_4__23 ;
    output d_arr_4__22 ;
    output d_arr_4__21 ;
    output d_arr_4__20 ;
    output d_arr_4__19 ;
    output d_arr_4__18 ;
    output d_arr_4__17 ;
    output d_arr_4__16 ;
    output d_arr_4__15 ;
    output d_arr_4__14 ;
    output d_arr_4__13 ;
    output d_arr_4__12 ;
    output d_arr_4__11 ;
    output d_arr_4__10 ;
    output d_arr_4__9 ;
    output d_arr_4__8 ;
    output d_arr_4__7 ;
    output d_arr_4__6 ;
    output d_arr_4__5 ;
    output d_arr_4__4 ;
    output d_arr_4__3 ;
    output d_arr_4__2 ;
    output d_arr_4__1 ;
    output d_arr_4__0 ;
    output d_arr_5__31 ;
    output d_arr_5__30 ;
    output d_arr_5__29 ;
    output d_arr_5__28 ;
    output d_arr_5__27 ;
    output d_arr_5__26 ;
    output d_arr_5__25 ;
    output d_arr_5__24 ;
    output d_arr_5__23 ;
    output d_arr_5__22 ;
    output d_arr_5__21 ;
    output d_arr_5__20 ;
    output d_arr_5__19 ;
    output d_arr_5__18 ;
    output d_arr_5__17 ;
    output d_arr_5__16 ;
    output d_arr_5__15 ;
    output d_arr_5__14 ;
    output d_arr_5__13 ;
    output d_arr_5__12 ;
    output d_arr_5__11 ;
    output d_arr_5__10 ;
    output d_arr_5__9 ;
    output d_arr_5__8 ;
    output d_arr_5__7 ;
    output d_arr_5__6 ;
    output d_arr_5__5 ;
    output d_arr_5__4 ;
    output d_arr_5__3 ;
    output d_arr_5__2 ;
    output d_arr_5__1 ;
    output d_arr_5__0 ;
    output d_arr_6__31 ;
    output d_arr_6__30 ;
    output d_arr_6__29 ;
    output d_arr_6__28 ;
    output d_arr_6__27 ;
    output d_arr_6__26 ;
    output d_arr_6__25 ;
    output d_arr_6__24 ;
    output d_arr_6__23 ;
    output d_arr_6__22 ;
    output d_arr_6__21 ;
    output d_arr_6__20 ;
    output d_arr_6__19 ;
    output d_arr_6__18 ;
    output d_arr_6__17 ;
    output d_arr_6__16 ;
    output d_arr_6__15 ;
    output d_arr_6__14 ;
    output d_arr_6__13 ;
    output d_arr_6__12 ;
    output d_arr_6__11 ;
    output d_arr_6__10 ;
    output d_arr_6__9 ;
    output d_arr_6__8 ;
    output d_arr_6__7 ;
    output d_arr_6__6 ;
    output d_arr_6__5 ;
    output d_arr_6__4 ;
    output d_arr_6__3 ;
    output d_arr_6__2 ;
    output d_arr_6__1 ;
    output d_arr_6__0 ;
    output d_arr_7__31 ;
    output d_arr_7__30 ;
    output d_arr_7__29 ;
    output d_arr_7__28 ;
    output d_arr_7__27 ;
    output d_arr_7__26 ;
    output d_arr_7__25 ;
    output d_arr_7__24 ;
    output d_arr_7__23 ;
    output d_arr_7__22 ;
    output d_arr_7__21 ;
    output d_arr_7__20 ;
    output d_arr_7__19 ;
    output d_arr_7__18 ;
    output d_arr_7__17 ;
    output d_arr_7__16 ;
    output d_arr_7__15 ;
    output d_arr_7__14 ;
    output d_arr_7__13 ;
    output d_arr_7__12 ;
    output d_arr_7__11 ;
    output d_arr_7__10 ;
    output d_arr_7__9 ;
    output d_arr_7__8 ;
    output d_arr_7__7 ;
    output d_arr_7__6 ;
    output d_arr_7__5 ;
    output d_arr_7__4 ;
    output d_arr_7__3 ;
    output d_arr_7__2 ;
    output d_arr_7__1 ;
    output d_arr_7__0 ;
    output d_arr_8__31 ;
    output d_arr_8__30 ;
    output d_arr_8__29 ;
    output d_arr_8__28 ;
    output d_arr_8__27 ;
    output d_arr_8__26 ;
    output d_arr_8__25 ;
    output d_arr_8__24 ;
    output d_arr_8__23 ;
    output d_arr_8__22 ;
    output d_arr_8__21 ;
    output d_arr_8__20 ;
    output d_arr_8__19 ;
    output d_arr_8__18 ;
    output d_arr_8__17 ;
    output d_arr_8__16 ;
    output d_arr_8__15 ;
    output d_arr_8__14 ;
    output d_arr_8__13 ;
    output d_arr_8__12 ;
    output d_arr_8__11 ;
    output d_arr_8__10 ;
    output d_arr_8__9 ;
    output d_arr_8__8 ;
    output d_arr_8__7 ;
    output d_arr_8__6 ;
    output d_arr_8__5 ;
    output d_arr_8__4 ;
    output d_arr_8__3 ;
    output d_arr_8__2 ;
    output d_arr_8__1 ;
    output d_arr_8__0 ;
    output d_arr_9__31 ;
    output d_arr_9__30 ;
    output d_arr_9__29 ;
    output d_arr_9__28 ;
    output d_arr_9__27 ;
    output d_arr_9__26 ;
    output d_arr_9__25 ;
    output d_arr_9__24 ;
    output d_arr_9__23 ;
    output d_arr_9__22 ;
    output d_arr_9__21 ;
    output d_arr_9__20 ;
    output d_arr_9__19 ;
    output d_arr_9__18 ;
    output d_arr_9__17 ;
    output d_arr_9__16 ;
    output d_arr_9__15 ;
    output d_arr_9__14 ;
    output d_arr_9__13 ;
    output d_arr_9__12 ;
    output d_arr_9__11 ;
    output d_arr_9__10 ;
    output d_arr_9__9 ;
    output d_arr_9__8 ;
    output d_arr_9__7 ;
    output d_arr_9__6 ;
    output d_arr_9__5 ;
    output d_arr_9__4 ;
    output d_arr_9__3 ;
    output d_arr_9__2 ;
    output d_arr_9__1 ;
    output d_arr_9__0 ;
    output d_arr_10__31 ;
    output d_arr_10__30 ;
    output d_arr_10__29 ;
    output d_arr_10__28 ;
    output d_arr_10__27 ;
    output d_arr_10__26 ;
    output d_arr_10__25 ;
    output d_arr_10__24 ;
    output d_arr_10__23 ;
    output d_arr_10__22 ;
    output d_arr_10__21 ;
    output d_arr_10__20 ;
    output d_arr_10__19 ;
    output d_arr_10__18 ;
    output d_arr_10__17 ;
    output d_arr_10__16 ;
    output d_arr_10__15 ;
    output d_arr_10__14 ;
    output d_arr_10__13 ;
    output d_arr_10__12 ;
    output d_arr_10__11 ;
    output d_arr_10__10 ;
    output d_arr_10__9 ;
    output d_arr_10__8 ;
    output d_arr_10__7 ;
    output d_arr_10__6 ;
    output d_arr_10__5 ;
    output d_arr_10__4 ;
    output d_arr_10__3 ;
    output d_arr_10__2 ;
    output d_arr_10__1 ;
    output d_arr_10__0 ;
    output d_arr_11__31 ;
    output d_arr_11__30 ;
    output d_arr_11__29 ;
    output d_arr_11__28 ;
    output d_arr_11__27 ;
    output d_arr_11__26 ;
    output d_arr_11__25 ;
    output d_arr_11__24 ;
    output d_arr_11__23 ;
    output d_arr_11__22 ;
    output d_arr_11__21 ;
    output d_arr_11__20 ;
    output d_arr_11__19 ;
    output d_arr_11__18 ;
    output d_arr_11__17 ;
    output d_arr_11__16 ;
    output d_arr_11__15 ;
    output d_arr_11__14 ;
    output d_arr_11__13 ;
    output d_arr_11__12 ;
    output d_arr_11__11 ;
    output d_arr_11__10 ;
    output d_arr_11__9 ;
    output d_arr_11__8 ;
    output d_arr_11__7 ;
    output d_arr_11__6 ;
    output d_arr_11__5 ;
    output d_arr_11__4 ;
    output d_arr_11__3 ;
    output d_arr_11__2 ;
    output d_arr_11__1 ;
    output d_arr_11__0 ;
    output d_arr_12__31 ;
    output d_arr_12__30 ;
    output d_arr_12__29 ;
    output d_arr_12__28 ;
    output d_arr_12__27 ;
    output d_arr_12__26 ;
    output d_arr_12__25 ;
    output d_arr_12__24 ;
    output d_arr_12__23 ;
    output d_arr_12__22 ;
    output d_arr_12__21 ;
    output d_arr_12__20 ;
    output d_arr_12__19 ;
    output d_arr_12__18 ;
    output d_arr_12__17 ;
    output d_arr_12__16 ;
    output d_arr_12__15 ;
    output d_arr_12__14 ;
    output d_arr_12__13 ;
    output d_arr_12__12 ;
    output d_arr_12__11 ;
    output d_arr_12__10 ;
    output d_arr_12__9 ;
    output d_arr_12__8 ;
    output d_arr_12__7 ;
    output d_arr_12__6 ;
    output d_arr_12__5 ;
    output d_arr_12__4 ;
    output d_arr_12__3 ;
    output d_arr_12__2 ;
    output d_arr_12__1 ;
    output d_arr_12__0 ;
    output d_arr_13__31 ;
    output d_arr_13__30 ;
    output d_arr_13__29 ;
    output d_arr_13__28 ;
    output d_arr_13__27 ;
    output d_arr_13__26 ;
    output d_arr_13__25 ;
    output d_arr_13__24 ;
    output d_arr_13__23 ;
    output d_arr_13__22 ;
    output d_arr_13__21 ;
    output d_arr_13__20 ;
    output d_arr_13__19 ;
    output d_arr_13__18 ;
    output d_arr_13__17 ;
    output d_arr_13__16 ;
    output d_arr_13__15 ;
    output d_arr_13__14 ;
    output d_arr_13__13 ;
    output d_arr_13__12 ;
    output d_arr_13__11 ;
    output d_arr_13__10 ;
    output d_arr_13__9 ;
    output d_arr_13__8 ;
    output d_arr_13__7 ;
    output d_arr_13__6 ;
    output d_arr_13__5 ;
    output d_arr_13__4 ;
    output d_arr_13__3 ;
    output d_arr_13__2 ;
    output d_arr_13__1 ;
    output d_arr_13__0 ;
    output d_arr_14__31 ;
    output d_arr_14__30 ;
    output d_arr_14__29 ;
    output d_arr_14__28 ;
    output d_arr_14__27 ;
    output d_arr_14__26 ;
    output d_arr_14__25 ;
    output d_arr_14__24 ;
    output d_arr_14__23 ;
    output d_arr_14__22 ;
    output d_arr_14__21 ;
    output d_arr_14__20 ;
    output d_arr_14__19 ;
    output d_arr_14__18 ;
    output d_arr_14__17 ;
    output d_arr_14__16 ;
    output d_arr_14__15 ;
    output d_arr_14__14 ;
    output d_arr_14__13 ;
    output d_arr_14__12 ;
    output d_arr_14__11 ;
    output d_arr_14__10 ;
    output d_arr_14__9 ;
    output d_arr_14__8 ;
    output d_arr_14__7 ;
    output d_arr_14__6 ;
    output d_arr_14__5 ;
    output d_arr_14__4 ;
    output d_arr_14__3 ;
    output d_arr_14__2 ;
    output d_arr_14__1 ;
    output d_arr_14__0 ;
    output d_arr_15__31 ;
    output d_arr_15__30 ;
    output d_arr_15__29 ;
    output d_arr_15__28 ;
    output d_arr_15__27 ;
    output d_arr_15__26 ;
    output d_arr_15__25 ;
    output d_arr_15__24 ;
    output d_arr_15__23 ;
    output d_arr_15__22 ;
    output d_arr_15__21 ;
    output d_arr_15__20 ;
    output d_arr_15__19 ;
    output d_arr_15__18 ;
    output d_arr_15__17 ;
    output d_arr_15__16 ;
    output d_arr_15__15 ;
    output d_arr_15__14 ;
    output d_arr_15__13 ;
    output d_arr_15__12 ;
    output d_arr_15__11 ;
    output d_arr_15__10 ;
    output d_arr_15__9 ;
    output d_arr_15__8 ;
    output d_arr_15__7 ;
    output d_arr_15__6 ;
    output d_arr_15__5 ;
    output d_arr_15__4 ;
    output d_arr_15__3 ;
    output d_arr_15__2 ;
    output d_arr_15__1 ;
    output d_arr_15__0 ;
    output d_arr_16__31 ;
    output d_arr_16__30 ;
    output d_arr_16__29 ;
    output d_arr_16__28 ;
    output d_arr_16__27 ;
    output d_arr_16__26 ;
    output d_arr_16__25 ;
    output d_arr_16__24 ;
    output d_arr_16__23 ;
    output d_arr_16__22 ;
    output d_arr_16__21 ;
    output d_arr_16__20 ;
    output d_arr_16__19 ;
    output d_arr_16__18 ;
    output d_arr_16__17 ;
    output d_arr_16__16 ;
    output d_arr_16__15 ;
    output d_arr_16__14 ;
    output d_arr_16__13 ;
    output d_arr_16__12 ;
    output d_arr_16__11 ;
    output d_arr_16__10 ;
    output d_arr_16__9 ;
    output d_arr_16__8 ;
    output d_arr_16__7 ;
    output d_arr_16__6 ;
    output d_arr_16__5 ;
    output d_arr_16__4 ;
    output d_arr_16__3 ;
    output d_arr_16__2 ;
    output d_arr_16__1 ;
    output d_arr_16__0 ;
    output d_arr_17__31 ;
    output d_arr_17__30 ;
    output d_arr_17__29 ;
    output d_arr_17__28 ;
    output d_arr_17__27 ;
    output d_arr_17__26 ;
    output d_arr_17__25 ;
    output d_arr_17__24 ;
    output d_arr_17__23 ;
    output d_arr_17__22 ;
    output d_arr_17__21 ;
    output d_arr_17__20 ;
    output d_arr_17__19 ;
    output d_arr_17__18 ;
    output d_arr_17__17 ;
    output d_arr_17__16 ;
    output d_arr_17__15 ;
    output d_arr_17__14 ;
    output d_arr_17__13 ;
    output d_arr_17__12 ;
    output d_arr_17__11 ;
    output d_arr_17__10 ;
    output d_arr_17__9 ;
    output d_arr_17__8 ;
    output d_arr_17__7 ;
    output d_arr_17__6 ;
    output d_arr_17__5 ;
    output d_arr_17__4 ;
    output d_arr_17__3 ;
    output d_arr_17__2 ;
    output d_arr_17__1 ;
    output d_arr_17__0 ;
    output d_arr_18__31 ;
    output d_arr_18__30 ;
    output d_arr_18__29 ;
    output d_arr_18__28 ;
    output d_arr_18__27 ;
    output d_arr_18__26 ;
    output d_arr_18__25 ;
    output d_arr_18__24 ;
    output d_arr_18__23 ;
    output d_arr_18__22 ;
    output d_arr_18__21 ;
    output d_arr_18__20 ;
    output d_arr_18__19 ;
    output d_arr_18__18 ;
    output d_arr_18__17 ;
    output d_arr_18__16 ;
    output d_arr_18__15 ;
    output d_arr_18__14 ;
    output d_arr_18__13 ;
    output d_arr_18__12 ;
    output d_arr_18__11 ;
    output d_arr_18__10 ;
    output d_arr_18__9 ;
    output d_arr_18__8 ;
    output d_arr_18__7 ;
    output d_arr_18__6 ;
    output d_arr_18__5 ;
    output d_arr_18__4 ;
    output d_arr_18__3 ;
    output d_arr_18__2 ;
    output d_arr_18__1 ;
    output d_arr_18__0 ;
    output d_arr_19__31 ;
    output d_arr_19__30 ;
    output d_arr_19__29 ;
    output d_arr_19__28 ;
    output d_arr_19__27 ;
    output d_arr_19__26 ;
    output d_arr_19__25 ;
    output d_arr_19__24 ;
    output d_arr_19__23 ;
    output d_arr_19__22 ;
    output d_arr_19__21 ;
    output d_arr_19__20 ;
    output d_arr_19__19 ;
    output d_arr_19__18 ;
    output d_arr_19__17 ;
    output d_arr_19__16 ;
    output d_arr_19__15 ;
    output d_arr_19__14 ;
    output d_arr_19__13 ;
    output d_arr_19__12 ;
    output d_arr_19__11 ;
    output d_arr_19__10 ;
    output d_arr_19__9 ;
    output d_arr_19__8 ;
    output d_arr_19__7 ;
    output d_arr_19__6 ;
    output d_arr_19__5 ;
    output d_arr_19__4 ;
    output d_arr_19__3 ;
    output d_arr_19__2 ;
    output d_arr_19__1 ;
    output d_arr_19__0 ;
    output d_arr_20__31 ;
    output d_arr_20__30 ;
    output d_arr_20__29 ;
    output d_arr_20__28 ;
    output d_arr_20__27 ;
    output d_arr_20__26 ;
    output d_arr_20__25 ;
    output d_arr_20__24 ;
    output d_arr_20__23 ;
    output d_arr_20__22 ;
    output d_arr_20__21 ;
    output d_arr_20__20 ;
    output d_arr_20__19 ;
    output d_arr_20__18 ;
    output d_arr_20__17 ;
    output d_arr_20__16 ;
    output d_arr_20__15 ;
    output d_arr_20__14 ;
    output d_arr_20__13 ;
    output d_arr_20__12 ;
    output d_arr_20__11 ;
    output d_arr_20__10 ;
    output d_arr_20__9 ;
    output d_arr_20__8 ;
    output d_arr_20__7 ;
    output d_arr_20__6 ;
    output d_arr_20__5 ;
    output d_arr_20__4 ;
    output d_arr_20__3 ;
    output d_arr_20__2 ;
    output d_arr_20__1 ;
    output d_arr_20__0 ;
    output d_arr_21__31 ;
    output d_arr_21__30 ;
    output d_arr_21__29 ;
    output d_arr_21__28 ;
    output d_arr_21__27 ;
    output d_arr_21__26 ;
    output d_arr_21__25 ;
    output d_arr_21__24 ;
    output d_arr_21__23 ;
    output d_arr_21__22 ;
    output d_arr_21__21 ;
    output d_arr_21__20 ;
    output d_arr_21__19 ;
    output d_arr_21__18 ;
    output d_arr_21__17 ;
    output d_arr_21__16 ;
    output d_arr_21__15 ;
    output d_arr_21__14 ;
    output d_arr_21__13 ;
    output d_arr_21__12 ;
    output d_arr_21__11 ;
    output d_arr_21__10 ;
    output d_arr_21__9 ;
    output d_arr_21__8 ;
    output d_arr_21__7 ;
    output d_arr_21__6 ;
    output d_arr_21__5 ;
    output d_arr_21__4 ;
    output d_arr_21__3 ;
    output d_arr_21__2 ;
    output d_arr_21__1 ;
    output d_arr_21__0 ;
    output d_arr_22__31 ;
    output d_arr_22__30 ;
    output d_arr_22__29 ;
    output d_arr_22__28 ;
    output d_arr_22__27 ;
    output d_arr_22__26 ;
    output d_arr_22__25 ;
    output d_arr_22__24 ;
    output d_arr_22__23 ;
    output d_arr_22__22 ;
    output d_arr_22__21 ;
    output d_arr_22__20 ;
    output d_arr_22__19 ;
    output d_arr_22__18 ;
    output d_arr_22__17 ;
    output d_arr_22__16 ;
    output d_arr_22__15 ;
    output d_arr_22__14 ;
    output d_arr_22__13 ;
    output d_arr_22__12 ;
    output d_arr_22__11 ;
    output d_arr_22__10 ;
    output d_arr_22__9 ;
    output d_arr_22__8 ;
    output d_arr_22__7 ;
    output d_arr_22__6 ;
    output d_arr_22__5 ;
    output d_arr_22__4 ;
    output d_arr_22__3 ;
    output d_arr_22__2 ;
    output d_arr_22__1 ;
    output d_arr_22__0 ;
    output d_arr_23__31 ;
    output d_arr_23__30 ;
    output d_arr_23__29 ;
    output d_arr_23__28 ;
    output d_arr_23__27 ;
    output d_arr_23__26 ;
    output d_arr_23__25 ;
    output d_arr_23__24 ;
    output d_arr_23__23 ;
    output d_arr_23__22 ;
    output d_arr_23__21 ;
    output d_arr_23__20 ;
    output d_arr_23__19 ;
    output d_arr_23__18 ;
    output d_arr_23__17 ;
    output d_arr_23__16 ;
    output d_arr_23__15 ;
    output d_arr_23__14 ;
    output d_arr_23__13 ;
    output d_arr_23__12 ;
    output d_arr_23__11 ;
    output d_arr_23__10 ;
    output d_arr_23__9 ;
    output d_arr_23__8 ;
    output d_arr_23__7 ;
    output d_arr_23__6 ;
    output d_arr_23__5 ;
    output d_arr_23__4 ;
    output d_arr_23__3 ;
    output d_arr_23__2 ;
    output d_arr_23__1 ;
    output d_arr_23__0 ;
    output d_arr_24__31 ;
    output d_arr_24__30 ;
    output d_arr_24__29 ;
    output d_arr_24__28 ;
    output d_arr_24__27 ;
    output d_arr_24__26 ;
    output d_arr_24__25 ;
    output d_arr_24__24 ;
    output d_arr_24__23 ;
    output d_arr_24__22 ;
    output d_arr_24__21 ;
    output d_arr_24__20 ;
    output d_arr_24__19 ;
    output d_arr_24__18 ;
    output d_arr_24__17 ;
    output d_arr_24__16 ;
    output d_arr_24__15 ;
    output d_arr_24__14 ;
    output d_arr_24__13 ;
    output d_arr_24__12 ;
    output d_arr_24__11 ;
    output d_arr_24__10 ;
    output d_arr_24__9 ;
    output d_arr_24__8 ;
    output d_arr_24__7 ;
    output d_arr_24__6 ;
    output d_arr_24__5 ;
    output d_arr_24__4 ;
    output d_arr_24__3 ;
    output d_arr_24__2 ;
    output d_arr_24__1 ;
    output d_arr_24__0 ;
    input q_arr_0__31 ;
    input q_arr_0__30 ;
    input q_arr_0__29 ;
    input q_arr_0__28 ;
    input q_arr_0__27 ;
    input q_arr_0__26 ;
    input q_arr_0__25 ;
    input q_arr_0__24 ;
    input q_arr_0__23 ;
    input q_arr_0__22 ;
    input q_arr_0__21 ;
    input q_arr_0__20 ;
    input q_arr_0__19 ;
    input q_arr_0__18 ;
    input q_arr_0__17 ;
    input q_arr_0__16 ;
    input q_arr_0__15 ;
    input q_arr_0__14 ;
    input q_arr_0__13 ;
    input q_arr_0__12 ;
    input q_arr_0__11 ;
    input q_arr_0__10 ;
    input q_arr_0__9 ;
    input q_arr_0__8 ;
    input q_arr_0__7 ;
    input q_arr_0__6 ;
    input q_arr_0__5 ;
    input q_arr_0__4 ;
    input q_arr_0__3 ;
    input q_arr_0__2 ;
    input q_arr_0__1 ;
    input q_arr_0__0 ;
    input q_arr_1__31 ;
    input q_arr_1__30 ;
    input q_arr_1__29 ;
    input q_arr_1__28 ;
    input q_arr_1__27 ;
    input q_arr_1__26 ;
    input q_arr_1__25 ;
    input q_arr_1__24 ;
    input q_arr_1__23 ;
    input q_arr_1__22 ;
    input q_arr_1__21 ;
    input q_arr_1__20 ;
    input q_arr_1__19 ;
    input q_arr_1__18 ;
    input q_arr_1__17 ;
    input q_arr_1__16 ;
    input q_arr_1__15 ;
    input q_arr_1__14 ;
    input q_arr_1__13 ;
    input q_arr_1__12 ;
    input q_arr_1__11 ;
    input q_arr_1__10 ;
    input q_arr_1__9 ;
    input q_arr_1__8 ;
    input q_arr_1__7 ;
    input q_arr_1__6 ;
    input q_arr_1__5 ;
    input q_arr_1__4 ;
    input q_arr_1__3 ;
    input q_arr_1__2 ;
    input q_arr_1__1 ;
    input q_arr_1__0 ;
    input q_arr_2__31 ;
    input q_arr_2__30 ;
    input q_arr_2__29 ;
    input q_arr_2__28 ;
    input q_arr_2__27 ;
    input q_arr_2__26 ;
    input q_arr_2__25 ;
    input q_arr_2__24 ;
    input q_arr_2__23 ;
    input q_arr_2__22 ;
    input q_arr_2__21 ;
    input q_arr_2__20 ;
    input q_arr_2__19 ;
    input q_arr_2__18 ;
    input q_arr_2__17 ;
    input q_arr_2__16 ;
    input q_arr_2__15 ;
    input q_arr_2__14 ;
    input q_arr_2__13 ;
    input q_arr_2__12 ;
    input q_arr_2__11 ;
    input q_arr_2__10 ;
    input q_arr_2__9 ;
    input q_arr_2__8 ;
    input q_arr_2__7 ;
    input q_arr_2__6 ;
    input q_arr_2__5 ;
    input q_arr_2__4 ;
    input q_arr_2__3 ;
    input q_arr_2__2 ;
    input q_arr_2__1 ;
    input q_arr_2__0 ;
    input q_arr_3__31 ;
    input q_arr_3__30 ;
    input q_arr_3__29 ;
    input q_arr_3__28 ;
    input q_arr_3__27 ;
    input q_arr_3__26 ;
    input q_arr_3__25 ;
    input q_arr_3__24 ;
    input q_arr_3__23 ;
    input q_arr_3__22 ;
    input q_arr_3__21 ;
    input q_arr_3__20 ;
    input q_arr_3__19 ;
    input q_arr_3__18 ;
    input q_arr_3__17 ;
    input q_arr_3__16 ;
    input q_arr_3__15 ;
    input q_arr_3__14 ;
    input q_arr_3__13 ;
    input q_arr_3__12 ;
    input q_arr_3__11 ;
    input q_arr_3__10 ;
    input q_arr_3__9 ;
    input q_arr_3__8 ;
    input q_arr_3__7 ;
    input q_arr_3__6 ;
    input q_arr_3__5 ;
    input q_arr_3__4 ;
    input q_arr_3__3 ;
    input q_arr_3__2 ;
    input q_arr_3__1 ;
    input q_arr_3__0 ;
    input q_arr_4__31 ;
    input q_arr_4__30 ;
    input q_arr_4__29 ;
    input q_arr_4__28 ;
    input q_arr_4__27 ;
    input q_arr_4__26 ;
    input q_arr_4__25 ;
    input q_arr_4__24 ;
    input q_arr_4__23 ;
    input q_arr_4__22 ;
    input q_arr_4__21 ;
    input q_arr_4__20 ;
    input q_arr_4__19 ;
    input q_arr_4__18 ;
    input q_arr_4__17 ;
    input q_arr_4__16 ;
    input q_arr_4__15 ;
    input q_arr_4__14 ;
    input q_arr_4__13 ;
    input q_arr_4__12 ;
    input q_arr_4__11 ;
    input q_arr_4__10 ;
    input q_arr_4__9 ;
    input q_arr_4__8 ;
    input q_arr_4__7 ;
    input q_arr_4__6 ;
    input q_arr_4__5 ;
    input q_arr_4__4 ;
    input q_arr_4__3 ;
    input q_arr_4__2 ;
    input q_arr_4__1 ;
    input q_arr_4__0 ;
    input q_arr_5__31 ;
    input q_arr_5__30 ;
    input q_arr_5__29 ;
    input q_arr_5__28 ;
    input q_arr_5__27 ;
    input q_arr_5__26 ;
    input q_arr_5__25 ;
    input q_arr_5__24 ;
    input q_arr_5__23 ;
    input q_arr_5__22 ;
    input q_arr_5__21 ;
    input q_arr_5__20 ;
    input q_arr_5__19 ;
    input q_arr_5__18 ;
    input q_arr_5__17 ;
    input q_arr_5__16 ;
    input q_arr_5__15 ;
    input q_arr_5__14 ;
    input q_arr_5__13 ;
    input q_arr_5__12 ;
    input q_arr_5__11 ;
    input q_arr_5__10 ;
    input q_arr_5__9 ;
    input q_arr_5__8 ;
    input q_arr_5__7 ;
    input q_arr_5__6 ;
    input q_arr_5__5 ;
    input q_arr_5__4 ;
    input q_arr_5__3 ;
    input q_arr_5__2 ;
    input q_arr_5__1 ;
    input q_arr_5__0 ;
    input q_arr_6__31 ;
    input q_arr_6__30 ;
    input q_arr_6__29 ;
    input q_arr_6__28 ;
    input q_arr_6__27 ;
    input q_arr_6__26 ;
    input q_arr_6__25 ;
    input q_arr_6__24 ;
    input q_arr_6__23 ;
    input q_arr_6__22 ;
    input q_arr_6__21 ;
    input q_arr_6__20 ;
    input q_arr_6__19 ;
    input q_arr_6__18 ;
    input q_arr_6__17 ;
    input q_arr_6__16 ;
    input q_arr_6__15 ;
    input q_arr_6__14 ;
    input q_arr_6__13 ;
    input q_arr_6__12 ;
    input q_arr_6__11 ;
    input q_arr_6__10 ;
    input q_arr_6__9 ;
    input q_arr_6__8 ;
    input q_arr_6__7 ;
    input q_arr_6__6 ;
    input q_arr_6__5 ;
    input q_arr_6__4 ;
    input q_arr_6__3 ;
    input q_arr_6__2 ;
    input q_arr_6__1 ;
    input q_arr_6__0 ;
    input q_arr_7__31 ;
    input q_arr_7__30 ;
    input q_arr_7__29 ;
    input q_arr_7__28 ;
    input q_arr_7__27 ;
    input q_arr_7__26 ;
    input q_arr_7__25 ;
    input q_arr_7__24 ;
    input q_arr_7__23 ;
    input q_arr_7__22 ;
    input q_arr_7__21 ;
    input q_arr_7__20 ;
    input q_arr_7__19 ;
    input q_arr_7__18 ;
    input q_arr_7__17 ;
    input q_arr_7__16 ;
    input q_arr_7__15 ;
    input q_arr_7__14 ;
    input q_arr_7__13 ;
    input q_arr_7__12 ;
    input q_arr_7__11 ;
    input q_arr_7__10 ;
    input q_arr_7__9 ;
    input q_arr_7__8 ;
    input q_arr_7__7 ;
    input q_arr_7__6 ;
    input q_arr_7__5 ;
    input q_arr_7__4 ;
    input q_arr_7__3 ;
    input q_arr_7__2 ;
    input q_arr_7__1 ;
    input q_arr_7__0 ;
    input q_arr_8__31 ;
    input q_arr_8__30 ;
    input q_arr_8__29 ;
    input q_arr_8__28 ;
    input q_arr_8__27 ;
    input q_arr_8__26 ;
    input q_arr_8__25 ;
    input q_arr_8__24 ;
    input q_arr_8__23 ;
    input q_arr_8__22 ;
    input q_arr_8__21 ;
    input q_arr_8__20 ;
    input q_arr_8__19 ;
    input q_arr_8__18 ;
    input q_arr_8__17 ;
    input q_arr_8__16 ;
    input q_arr_8__15 ;
    input q_arr_8__14 ;
    input q_arr_8__13 ;
    input q_arr_8__12 ;
    input q_arr_8__11 ;
    input q_arr_8__10 ;
    input q_arr_8__9 ;
    input q_arr_8__8 ;
    input q_arr_8__7 ;
    input q_arr_8__6 ;
    input q_arr_8__5 ;
    input q_arr_8__4 ;
    input q_arr_8__3 ;
    input q_arr_8__2 ;
    input q_arr_8__1 ;
    input q_arr_8__0 ;
    input q_arr_9__31 ;
    input q_arr_9__30 ;
    input q_arr_9__29 ;
    input q_arr_9__28 ;
    input q_arr_9__27 ;
    input q_arr_9__26 ;
    input q_arr_9__25 ;
    input q_arr_9__24 ;
    input q_arr_9__23 ;
    input q_arr_9__22 ;
    input q_arr_9__21 ;
    input q_arr_9__20 ;
    input q_arr_9__19 ;
    input q_arr_9__18 ;
    input q_arr_9__17 ;
    input q_arr_9__16 ;
    input q_arr_9__15 ;
    input q_arr_9__14 ;
    input q_arr_9__13 ;
    input q_arr_9__12 ;
    input q_arr_9__11 ;
    input q_arr_9__10 ;
    input q_arr_9__9 ;
    input q_arr_9__8 ;
    input q_arr_9__7 ;
    input q_arr_9__6 ;
    input q_arr_9__5 ;
    input q_arr_9__4 ;
    input q_arr_9__3 ;
    input q_arr_9__2 ;
    input q_arr_9__1 ;
    input q_arr_9__0 ;
    input q_arr_10__31 ;
    input q_arr_10__30 ;
    input q_arr_10__29 ;
    input q_arr_10__28 ;
    input q_arr_10__27 ;
    input q_arr_10__26 ;
    input q_arr_10__25 ;
    input q_arr_10__24 ;
    input q_arr_10__23 ;
    input q_arr_10__22 ;
    input q_arr_10__21 ;
    input q_arr_10__20 ;
    input q_arr_10__19 ;
    input q_arr_10__18 ;
    input q_arr_10__17 ;
    input q_arr_10__16 ;
    input q_arr_10__15 ;
    input q_arr_10__14 ;
    input q_arr_10__13 ;
    input q_arr_10__12 ;
    input q_arr_10__11 ;
    input q_arr_10__10 ;
    input q_arr_10__9 ;
    input q_arr_10__8 ;
    input q_arr_10__7 ;
    input q_arr_10__6 ;
    input q_arr_10__5 ;
    input q_arr_10__4 ;
    input q_arr_10__3 ;
    input q_arr_10__2 ;
    input q_arr_10__1 ;
    input q_arr_10__0 ;
    input q_arr_11__31 ;
    input q_arr_11__30 ;
    input q_arr_11__29 ;
    input q_arr_11__28 ;
    input q_arr_11__27 ;
    input q_arr_11__26 ;
    input q_arr_11__25 ;
    input q_arr_11__24 ;
    input q_arr_11__23 ;
    input q_arr_11__22 ;
    input q_arr_11__21 ;
    input q_arr_11__20 ;
    input q_arr_11__19 ;
    input q_arr_11__18 ;
    input q_arr_11__17 ;
    input q_arr_11__16 ;
    input q_arr_11__15 ;
    input q_arr_11__14 ;
    input q_arr_11__13 ;
    input q_arr_11__12 ;
    input q_arr_11__11 ;
    input q_arr_11__10 ;
    input q_arr_11__9 ;
    input q_arr_11__8 ;
    input q_arr_11__7 ;
    input q_arr_11__6 ;
    input q_arr_11__5 ;
    input q_arr_11__4 ;
    input q_arr_11__3 ;
    input q_arr_11__2 ;
    input q_arr_11__1 ;
    input q_arr_11__0 ;
    input q_arr_12__31 ;
    input q_arr_12__30 ;
    input q_arr_12__29 ;
    input q_arr_12__28 ;
    input q_arr_12__27 ;
    input q_arr_12__26 ;
    input q_arr_12__25 ;
    input q_arr_12__24 ;
    input q_arr_12__23 ;
    input q_arr_12__22 ;
    input q_arr_12__21 ;
    input q_arr_12__20 ;
    input q_arr_12__19 ;
    input q_arr_12__18 ;
    input q_arr_12__17 ;
    input q_arr_12__16 ;
    input q_arr_12__15 ;
    input q_arr_12__14 ;
    input q_arr_12__13 ;
    input q_arr_12__12 ;
    input q_arr_12__11 ;
    input q_arr_12__10 ;
    input q_arr_12__9 ;
    input q_arr_12__8 ;
    input q_arr_12__7 ;
    input q_arr_12__6 ;
    input q_arr_12__5 ;
    input q_arr_12__4 ;
    input q_arr_12__3 ;
    input q_arr_12__2 ;
    input q_arr_12__1 ;
    input q_arr_12__0 ;
    input q_arr_13__31 ;
    input q_arr_13__30 ;
    input q_arr_13__29 ;
    input q_arr_13__28 ;
    input q_arr_13__27 ;
    input q_arr_13__26 ;
    input q_arr_13__25 ;
    input q_arr_13__24 ;
    input q_arr_13__23 ;
    input q_arr_13__22 ;
    input q_arr_13__21 ;
    input q_arr_13__20 ;
    input q_arr_13__19 ;
    input q_arr_13__18 ;
    input q_arr_13__17 ;
    input q_arr_13__16 ;
    input q_arr_13__15 ;
    input q_arr_13__14 ;
    input q_arr_13__13 ;
    input q_arr_13__12 ;
    input q_arr_13__11 ;
    input q_arr_13__10 ;
    input q_arr_13__9 ;
    input q_arr_13__8 ;
    input q_arr_13__7 ;
    input q_arr_13__6 ;
    input q_arr_13__5 ;
    input q_arr_13__4 ;
    input q_arr_13__3 ;
    input q_arr_13__2 ;
    input q_arr_13__1 ;
    input q_arr_13__0 ;
    input q_arr_14__31 ;
    input q_arr_14__30 ;
    input q_arr_14__29 ;
    input q_arr_14__28 ;
    input q_arr_14__27 ;
    input q_arr_14__26 ;
    input q_arr_14__25 ;
    input q_arr_14__24 ;
    input q_arr_14__23 ;
    input q_arr_14__22 ;
    input q_arr_14__21 ;
    input q_arr_14__20 ;
    input q_arr_14__19 ;
    input q_arr_14__18 ;
    input q_arr_14__17 ;
    input q_arr_14__16 ;
    input q_arr_14__15 ;
    input q_arr_14__14 ;
    input q_arr_14__13 ;
    input q_arr_14__12 ;
    input q_arr_14__11 ;
    input q_arr_14__10 ;
    input q_arr_14__9 ;
    input q_arr_14__8 ;
    input q_arr_14__7 ;
    input q_arr_14__6 ;
    input q_arr_14__5 ;
    input q_arr_14__4 ;
    input q_arr_14__3 ;
    input q_arr_14__2 ;
    input q_arr_14__1 ;
    input q_arr_14__0 ;
    input q_arr_15__31 ;
    input q_arr_15__30 ;
    input q_arr_15__29 ;
    input q_arr_15__28 ;
    input q_arr_15__27 ;
    input q_arr_15__26 ;
    input q_arr_15__25 ;
    input q_arr_15__24 ;
    input q_arr_15__23 ;
    input q_arr_15__22 ;
    input q_arr_15__21 ;
    input q_arr_15__20 ;
    input q_arr_15__19 ;
    input q_arr_15__18 ;
    input q_arr_15__17 ;
    input q_arr_15__16 ;
    input q_arr_15__15 ;
    input q_arr_15__14 ;
    input q_arr_15__13 ;
    input q_arr_15__12 ;
    input q_arr_15__11 ;
    input q_arr_15__10 ;
    input q_arr_15__9 ;
    input q_arr_15__8 ;
    input q_arr_15__7 ;
    input q_arr_15__6 ;
    input q_arr_15__5 ;
    input q_arr_15__4 ;
    input q_arr_15__3 ;
    input q_arr_15__2 ;
    input q_arr_15__1 ;
    input q_arr_15__0 ;
    input q_arr_16__31 ;
    input q_arr_16__30 ;
    input q_arr_16__29 ;
    input q_arr_16__28 ;
    input q_arr_16__27 ;
    input q_arr_16__26 ;
    input q_arr_16__25 ;
    input q_arr_16__24 ;
    input q_arr_16__23 ;
    input q_arr_16__22 ;
    input q_arr_16__21 ;
    input q_arr_16__20 ;
    input q_arr_16__19 ;
    input q_arr_16__18 ;
    input q_arr_16__17 ;
    input q_arr_16__16 ;
    input q_arr_16__15 ;
    input q_arr_16__14 ;
    input q_arr_16__13 ;
    input q_arr_16__12 ;
    input q_arr_16__11 ;
    input q_arr_16__10 ;
    input q_arr_16__9 ;
    input q_arr_16__8 ;
    input q_arr_16__7 ;
    input q_arr_16__6 ;
    input q_arr_16__5 ;
    input q_arr_16__4 ;
    input q_arr_16__3 ;
    input q_arr_16__2 ;
    input q_arr_16__1 ;
    input q_arr_16__0 ;
    input q_arr_17__31 ;
    input q_arr_17__30 ;
    input q_arr_17__29 ;
    input q_arr_17__28 ;
    input q_arr_17__27 ;
    input q_arr_17__26 ;
    input q_arr_17__25 ;
    input q_arr_17__24 ;
    input q_arr_17__23 ;
    input q_arr_17__22 ;
    input q_arr_17__21 ;
    input q_arr_17__20 ;
    input q_arr_17__19 ;
    input q_arr_17__18 ;
    input q_arr_17__17 ;
    input q_arr_17__16 ;
    input q_arr_17__15 ;
    input q_arr_17__14 ;
    input q_arr_17__13 ;
    input q_arr_17__12 ;
    input q_arr_17__11 ;
    input q_arr_17__10 ;
    input q_arr_17__9 ;
    input q_arr_17__8 ;
    input q_arr_17__7 ;
    input q_arr_17__6 ;
    input q_arr_17__5 ;
    input q_arr_17__4 ;
    input q_arr_17__3 ;
    input q_arr_17__2 ;
    input q_arr_17__1 ;
    input q_arr_17__0 ;
    input q_arr_18__31 ;
    input q_arr_18__30 ;
    input q_arr_18__29 ;
    input q_arr_18__28 ;
    input q_arr_18__27 ;
    input q_arr_18__26 ;
    input q_arr_18__25 ;
    input q_arr_18__24 ;
    input q_arr_18__23 ;
    input q_arr_18__22 ;
    input q_arr_18__21 ;
    input q_arr_18__20 ;
    input q_arr_18__19 ;
    input q_arr_18__18 ;
    input q_arr_18__17 ;
    input q_arr_18__16 ;
    input q_arr_18__15 ;
    input q_arr_18__14 ;
    input q_arr_18__13 ;
    input q_arr_18__12 ;
    input q_arr_18__11 ;
    input q_arr_18__10 ;
    input q_arr_18__9 ;
    input q_arr_18__8 ;
    input q_arr_18__7 ;
    input q_arr_18__6 ;
    input q_arr_18__5 ;
    input q_arr_18__4 ;
    input q_arr_18__3 ;
    input q_arr_18__2 ;
    input q_arr_18__1 ;
    input q_arr_18__0 ;
    input q_arr_19__31 ;
    input q_arr_19__30 ;
    input q_arr_19__29 ;
    input q_arr_19__28 ;
    input q_arr_19__27 ;
    input q_arr_19__26 ;
    input q_arr_19__25 ;
    input q_arr_19__24 ;
    input q_arr_19__23 ;
    input q_arr_19__22 ;
    input q_arr_19__21 ;
    input q_arr_19__20 ;
    input q_arr_19__19 ;
    input q_arr_19__18 ;
    input q_arr_19__17 ;
    input q_arr_19__16 ;
    input q_arr_19__15 ;
    input q_arr_19__14 ;
    input q_arr_19__13 ;
    input q_arr_19__12 ;
    input q_arr_19__11 ;
    input q_arr_19__10 ;
    input q_arr_19__9 ;
    input q_arr_19__8 ;
    input q_arr_19__7 ;
    input q_arr_19__6 ;
    input q_arr_19__5 ;
    input q_arr_19__4 ;
    input q_arr_19__3 ;
    input q_arr_19__2 ;
    input q_arr_19__1 ;
    input q_arr_19__0 ;
    input q_arr_20__31 ;
    input q_arr_20__30 ;
    input q_arr_20__29 ;
    input q_arr_20__28 ;
    input q_arr_20__27 ;
    input q_arr_20__26 ;
    input q_arr_20__25 ;
    input q_arr_20__24 ;
    input q_arr_20__23 ;
    input q_arr_20__22 ;
    input q_arr_20__21 ;
    input q_arr_20__20 ;
    input q_arr_20__19 ;
    input q_arr_20__18 ;
    input q_arr_20__17 ;
    input q_arr_20__16 ;
    input q_arr_20__15 ;
    input q_arr_20__14 ;
    input q_arr_20__13 ;
    input q_arr_20__12 ;
    input q_arr_20__11 ;
    input q_arr_20__10 ;
    input q_arr_20__9 ;
    input q_arr_20__8 ;
    input q_arr_20__7 ;
    input q_arr_20__6 ;
    input q_arr_20__5 ;
    input q_arr_20__4 ;
    input q_arr_20__3 ;
    input q_arr_20__2 ;
    input q_arr_20__1 ;
    input q_arr_20__0 ;
    input q_arr_21__31 ;
    input q_arr_21__30 ;
    input q_arr_21__29 ;
    input q_arr_21__28 ;
    input q_arr_21__27 ;
    input q_arr_21__26 ;
    input q_arr_21__25 ;
    input q_arr_21__24 ;
    input q_arr_21__23 ;
    input q_arr_21__22 ;
    input q_arr_21__21 ;
    input q_arr_21__20 ;
    input q_arr_21__19 ;
    input q_arr_21__18 ;
    input q_arr_21__17 ;
    input q_arr_21__16 ;
    input q_arr_21__15 ;
    input q_arr_21__14 ;
    input q_arr_21__13 ;
    input q_arr_21__12 ;
    input q_arr_21__11 ;
    input q_arr_21__10 ;
    input q_arr_21__9 ;
    input q_arr_21__8 ;
    input q_arr_21__7 ;
    input q_arr_21__6 ;
    input q_arr_21__5 ;
    input q_arr_21__4 ;
    input q_arr_21__3 ;
    input q_arr_21__2 ;
    input q_arr_21__1 ;
    input q_arr_21__0 ;
    input q_arr_22__31 ;
    input q_arr_22__30 ;
    input q_arr_22__29 ;
    input q_arr_22__28 ;
    input q_arr_22__27 ;
    input q_arr_22__26 ;
    input q_arr_22__25 ;
    input q_arr_22__24 ;
    input q_arr_22__23 ;
    input q_arr_22__22 ;
    input q_arr_22__21 ;
    input q_arr_22__20 ;
    input q_arr_22__19 ;
    input q_arr_22__18 ;
    input q_arr_22__17 ;
    input q_arr_22__16 ;
    input q_arr_22__15 ;
    input q_arr_22__14 ;
    input q_arr_22__13 ;
    input q_arr_22__12 ;
    input q_arr_22__11 ;
    input q_arr_22__10 ;
    input q_arr_22__9 ;
    input q_arr_22__8 ;
    input q_arr_22__7 ;
    input q_arr_22__6 ;
    input q_arr_22__5 ;
    input q_arr_22__4 ;
    input q_arr_22__3 ;
    input q_arr_22__2 ;
    input q_arr_22__1 ;
    input q_arr_22__0 ;
    input q_arr_23__31 ;
    input q_arr_23__30 ;
    input q_arr_23__29 ;
    input q_arr_23__28 ;
    input q_arr_23__27 ;
    input q_arr_23__26 ;
    input q_arr_23__25 ;
    input q_arr_23__24 ;
    input q_arr_23__23 ;
    input q_arr_23__22 ;
    input q_arr_23__21 ;
    input q_arr_23__20 ;
    input q_arr_23__19 ;
    input q_arr_23__18 ;
    input q_arr_23__17 ;
    input q_arr_23__16 ;
    input q_arr_23__15 ;
    input q_arr_23__14 ;
    input q_arr_23__13 ;
    input q_arr_23__12 ;
    input q_arr_23__11 ;
    input q_arr_23__10 ;
    input q_arr_23__9 ;
    input q_arr_23__8 ;
    input q_arr_23__7 ;
    input q_arr_23__6 ;
    input q_arr_23__5 ;
    input q_arr_23__4 ;
    input q_arr_23__3 ;
    input q_arr_23__2 ;
    input q_arr_23__1 ;
    input q_arr_23__0 ;
    input q_arr_24__31 ;
    input q_arr_24__30 ;
    input q_arr_24__29 ;
    input q_arr_24__28 ;
    input q_arr_24__27 ;
    input q_arr_24__26 ;
    input q_arr_24__25 ;
    input q_arr_24__24 ;
    input q_arr_24__23 ;
    input q_arr_24__22 ;
    input q_arr_24__21 ;
    input q_arr_24__20 ;
    input q_arr_24__19 ;
    input q_arr_24__18 ;
    input q_arr_24__17 ;
    input q_arr_24__16 ;
    input q_arr_24__15 ;
    input q_arr_24__14 ;
    input q_arr_24__13 ;
    input q_arr_24__12 ;
    input q_arr_24__11 ;
    input q_arr_24__10 ;
    input q_arr_24__9 ;
    input q_arr_24__8 ;
    input q_arr_24__7 ;
    input q_arr_24__6 ;
    input q_arr_24__5 ;
    input q_arr_24__4 ;
    input q_arr_24__3 ;
    input q_arr_24__2 ;
    input q_arr_24__1 ;
    input q_arr_24__0 ;

    wire nx205, nx207, nx209, nx211, nx213, nx215, nx217, nx219, nx221, nx223, 
         nx225, nx227;



    assign d_arr_1__15 = d_arr_0__15 ;
    assign d_arr_2__31 = d_arr_0__15 ;
    assign d_arr_2__30 = d_arr_0__15 ;
    assign d_arr_2__29 = d_arr_0__15 ;
    assign d_arr_2__28 = d_arr_0__15 ;
    assign d_arr_2__27 = d_arr_0__15 ;
    assign d_arr_2__26 = d_arr_0__15 ;
    assign d_arr_2__25 = d_arr_0__15 ;
    assign d_arr_2__24 = d_arr_0__15 ;
    assign d_arr_2__23 = d_arr_0__15 ;
    assign d_arr_2__22 = d_arr_0__15 ;
    assign d_arr_2__21 = d_arr_0__15 ;
    assign d_arr_2__20 = d_arr_0__15 ;
    assign d_arr_2__19 = d_arr_0__15 ;
    assign d_arr_2__18 = d_arr_0__15 ;
    assign d_arr_2__17 = d_arr_0__15 ;
    assign d_arr_2__16 = d_arr_0__15 ;
    assign d_arr_2__15 = d_arr_0__15 ;
    assign d_arr_2__14 = d_arr_0__15 ;
    assign d_arr_2__13 = d_arr_0__15 ;
    assign d_arr_2__12 = d_arr_0__15 ;
    assign d_arr_2__11 = d_arr_0__15 ;
    assign d_arr_2__10 = d_arr_0__15 ;
    assign d_arr_2__9 = d_arr_0__15 ;
    assign d_arr_2__8 = d_arr_0__15 ;
    assign d_arr_2__7 = d_arr_0__15 ;
    assign d_arr_2__6 = d_arr_0__15 ;
    assign d_arr_2__5 = d_arr_0__15 ;
    assign d_arr_2__4 = d_arr_0__15 ;
    assign d_arr_2__3 = d_arr_0__15 ;
    assign d_arr_2__2 = d_arr_0__15 ;
    assign d_arr_2__1 = d_arr_0__15 ;
    assign d_arr_2__0 = d_arr_0__15 ;
    assign d_arr_3__31 = d_arr_0__15 ;
    assign d_arr_3__30 = d_arr_0__15 ;
    assign d_arr_3__29 = d_arr_0__15 ;
    assign d_arr_3__28 = d_arr_0__15 ;
    assign d_arr_3__27 = d_arr_0__15 ;
    assign d_arr_3__26 = d_arr_0__15 ;
    assign d_arr_3__25 = d_arr_0__15 ;
    assign d_arr_3__24 = d_arr_0__15 ;
    assign d_arr_3__23 = d_arr_0__15 ;
    assign d_arr_3__22 = d_arr_0__15 ;
    assign d_arr_3__21 = d_arr_0__15 ;
    assign d_arr_3__20 = d_arr_0__15 ;
    assign d_arr_3__19 = d_arr_0__15 ;
    assign d_arr_3__18 = d_arr_0__15 ;
    assign d_arr_3__17 = d_arr_0__15 ;
    assign d_arr_3__16 = d_arr_0__15 ;
    assign d_arr_3__15 = d_arr_0__15 ;
    assign d_arr_3__14 = d_arr_0__15 ;
    assign d_arr_3__13 = d_arr_0__15 ;
    assign d_arr_3__12 = d_arr_0__15 ;
    assign d_arr_3__11 = d_arr_0__15 ;
    assign d_arr_3__10 = d_arr_0__15 ;
    assign d_arr_3__9 = d_arr_0__15 ;
    assign d_arr_3__8 = d_arr_0__15 ;
    assign d_arr_3__7 = d_arr_0__15 ;
    assign d_arr_3__6 = d_arr_0__15 ;
    assign d_arr_3__5 = d_arr_0__15 ;
    assign d_arr_3__4 = d_arr_0__15 ;
    assign d_arr_3__3 = d_arr_0__15 ;
    assign d_arr_3__2 = d_arr_0__15 ;
    assign d_arr_3__1 = d_arr_0__15 ;
    assign d_arr_3__0 = d_arr_0__15 ;
    assign d_arr_4__31 = d_arr_0__15 ;
    assign d_arr_4__30 = d_arr_0__15 ;
    assign d_arr_4__29 = d_arr_0__15 ;
    assign d_arr_4__28 = d_arr_0__15 ;
    assign d_arr_4__27 = d_arr_0__15 ;
    assign d_arr_4__26 = d_arr_0__15 ;
    assign d_arr_4__25 = d_arr_0__15 ;
    assign d_arr_4__24 = d_arr_0__15 ;
    assign d_arr_4__23 = d_arr_0__15 ;
    assign d_arr_4__22 = d_arr_0__15 ;
    assign d_arr_4__21 = d_arr_0__15 ;
    assign d_arr_4__20 = d_arr_0__15 ;
    assign d_arr_4__19 = d_arr_0__15 ;
    assign d_arr_4__18 = d_arr_0__15 ;
    assign d_arr_4__17 = d_arr_0__15 ;
    assign d_arr_4__16 = d_arr_0__15 ;
    assign d_arr_4__15 = d_arr_0__15 ;
    assign d_arr_4__14 = d_arr_0__15 ;
    assign d_arr_4__13 = d_arr_0__15 ;
    assign d_arr_4__12 = d_arr_0__15 ;
    assign d_arr_4__11 = d_arr_0__15 ;
    assign d_arr_4__10 = d_arr_0__15 ;
    assign d_arr_4__9 = d_arr_0__15 ;
    assign d_arr_4__8 = d_arr_0__15 ;
    assign d_arr_4__7 = d_arr_0__15 ;
    assign d_arr_4__6 = d_arr_0__15 ;
    assign d_arr_4__5 = d_arr_0__15 ;
    assign d_arr_4__4 = d_arr_0__15 ;
    assign d_arr_4__3 = d_arr_0__15 ;
    assign d_arr_4__2 = d_arr_0__15 ;
    assign d_arr_4__1 = d_arr_0__15 ;
    assign d_arr_4__0 = d_arr_0__15 ;
    assign d_arr_5__31 = d_arr_0__15 ;
    assign d_arr_5__30 = d_arr_0__15 ;
    assign d_arr_5__29 = d_arr_0__15 ;
    assign d_arr_5__28 = d_arr_0__15 ;
    assign d_arr_5__27 = d_arr_0__15 ;
    assign d_arr_5__26 = d_arr_0__15 ;
    assign d_arr_5__25 = d_arr_0__15 ;
    assign d_arr_5__24 = d_arr_0__15 ;
    assign d_arr_5__23 = d_arr_0__15 ;
    assign d_arr_5__22 = d_arr_0__15 ;
    assign d_arr_5__21 = d_arr_0__15 ;
    assign d_arr_5__20 = d_arr_0__15 ;
    assign d_arr_5__19 = d_arr_0__15 ;
    assign d_arr_5__18 = d_arr_0__15 ;
    assign d_arr_5__17 = d_arr_0__15 ;
    assign d_arr_5__16 = d_arr_0__15 ;
    assign d_arr_5__15 = d_arr_0__15 ;
    assign d_arr_5__14 = d_arr_0__15 ;
    assign d_arr_5__13 = d_arr_0__15 ;
    assign d_arr_5__12 = d_arr_0__15 ;
    assign d_arr_5__11 = d_arr_0__15 ;
    assign d_arr_5__10 = d_arr_0__15 ;
    assign d_arr_5__9 = d_arr_0__15 ;
    assign d_arr_5__8 = d_arr_0__15 ;
    assign d_arr_5__7 = d_arr_0__15 ;
    assign d_arr_5__6 = d_arr_0__15 ;
    assign d_arr_5__5 = d_arr_0__15 ;
    assign d_arr_5__4 = d_arr_0__15 ;
    assign d_arr_5__3 = d_arr_0__15 ;
    assign d_arr_5__2 = d_arr_0__15 ;
    assign d_arr_5__1 = d_arr_0__15 ;
    assign d_arr_5__0 = d_arr_0__15 ;
    assign d_arr_6__31 = d_arr_0__15 ;
    assign d_arr_6__30 = d_arr_0__15 ;
    assign d_arr_6__29 = d_arr_0__15 ;
    assign d_arr_6__28 = d_arr_0__15 ;
    assign d_arr_6__27 = d_arr_0__15 ;
    assign d_arr_6__26 = d_arr_0__15 ;
    assign d_arr_6__25 = d_arr_0__15 ;
    assign d_arr_6__24 = d_arr_0__15 ;
    assign d_arr_6__23 = d_arr_0__15 ;
    assign d_arr_6__22 = d_arr_0__15 ;
    assign d_arr_6__21 = d_arr_0__15 ;
    assign d_arr_6__20 = d_arr_0__15 ;
    assign d_arr_6__19 = d_arr_0__15 ;
    assign d_arr_6__18 = d_arr_0__15 ;
    assign d_arr_6__17 = d_arr_0__15 ;
    assign d_arr_6__16 = d_arr_0__15 ;
    assign d_arr_6__15 = d_arr_0__15 ;
    assign d_arr_6__14 = d_arr_0__15 ;
    assign d_arr_6__13 = d_arr_0__15 ;
    assign d_arr_6__12 = d_arr_0__15 ;
    assign d_arr_6__11 = d_arr_0__15 ;
    assign d_arr_6__10 = d_arr_0__15 ;
    assign d_arr_6__9 = d_arr_0__15 ;
    assign d_arr_6__8 = d_arr_0__15 ;
    assign d_arr_6__7 = d_arr_0__15 ;
    assign d_arr_6__6 = d_arr_0__15 ;
    assign d_arr_6__5 = d_arr_0__15 ;
    assign d_arr_6__4 = d_arr_0__15 ;
    assign d_arr_6__3 = d_arr_0__15 ;
    assign d_arr_6__2 = d_arr_0__15 ;
    assign d_arr_6__1 = d_arr_0__15 ;
    assign d_arr_6__0 = d_arr_0__15 ;
    assign d_arr_7__31 = d_arr_0__15 ;
    assign d_arr_7__30 = d_arr_0__15 ;
    assign d_arr_7__29 = d_arr_0__15 ;
    assign d_arr_7__28 = d_arr_0__15 ;
    assign d_arr_7__27 = d_arr_0__15 ;
    assign d_arr_7__26 = d_arr_0__15 ;
    assign d_arr_7__25 = d_arr_0__15 ;
    assign d_arr_7__24 = d_arr_0__15 ;
    assign d_arr_7__23 = d_arr_0__15 ;
    assign d_arr_7__22 = d_arr_0__15 ;
    assign d_arr_7__21 = d_arr_0__15 ;
    assign d_arr_7__20 = d_arr_0__15 ;
    assign d_arr_7__19 = d_arr_0__15 ;
    assign d_arr_7__18 = d_arr_0__15 ;
    assign d_arr_7__17 = d_arr_0__15 ;
    assign d_arr_7__16 = d_arr_0__15 ;
    assign d_arr_7__15 = d_arr_0__15 ;
    assign d_arr_7__14 = d_arr_0__15 ;
    assign d_arr_7__13 = d_arr_0__15 ;
    assign d_arr_7__12 = d_arr_0__15 ;
    assign d_arr_7__11 = d_arr_0__15 ;
    assign d_arr_7__10 = d_arr_0__15 ;
    assign d_arr_7__9 = d_arr_0__15 ;
    assign d_arr_7__8 = d_arr_0__15 ;
    assign d_arr_7__7 = d_arr_0__15 ;
    assign d_arr_7__6 = d_arr_0__15 ;
    assign d_arr_7__5 = d_arr_0__15 ;
    assign d_arr_7__4 = d_arr_0__15 ;
    assign d_arr_7__3 = d_arr_0__15 ;
    assign d_arr_7__2 = d_arr_0__15 ;
    assign d_arr_7__1 = d_arr_0__15 ;
    assign d_arr_7__0 = d_arr_0__15 ;
    assign d_arr_8__31 = d_arr_0__15 ;
    assign d_arr_8__30 = d_arr_0__15 ;
    assign d_arr_8__29 = d_arr_0__15 ;
    assign d_arr_8__28 = d_arr_0__15 ;
    assign d_arr_8__27 = d_arr_0__15 ;
    assign d_arr_8__26 = d_arr_0__15 ;
    assign d_arr_8__25 = d_arr_0__15 ;
    assign d_arr_8__24 = d_arr_0__15 ;
    assign d_arr_8__23 = d_arr_0__15 ;
    assign d_arr_8__22 = d_arr_0__15 ;
    assign d_arr_8__21 = d_arr_0__15 ;
    assign d_arr_8__20 = d_arr_0__15 ;
    assign d_arr_8__19 = d_arr_0__15 ;
    assign d_arr_8__18 = d_arr_0__15 ;
    assign d_arr_8__17 = d_arr_0__15 ;
    assign d_arr_8__16 = d_arr_0__15 ;
    assign d_arr_8__15 = d_arr_0__15 ;
    assign d_arr_8__14 = d_arr_0__15 ;
    assign d_arr_8__13 = d_arr_0__15 ;
    assign d_arr_8__12 = d_arr_0__15 ;
    assign d_arr_8__11 = d_arr_0__15 ;
    assign d_arr_8__10 = d_arr_0__15 ;
    assign d_arr_8__9 = d_arr_0__15 ;
    assign d_arr_8__8 = d_arr_0__15 ;
    assign d_arr_8__7 = d_arr_0__15 ;
    assign d_arr_8__6 = d_arr_0__15 ;
    assign d_arr_8__5 = d_arr_0__15 ;
    assign d_arr_8__4 = d_arr_0__15 ;
    assign d_arr_8__3 = d_arr_0__15 ;
    assign d_arr_8__2 = d_arr_0__15 ;
    assign d_arr_8__1 = d_arr_0__15 ;
    assign d_arr_8__0 = d_arr_0__15 ;
    assign d_arr_9__31 = d_arr_0__15 ;
    assign d_arr_9__30 = d_arr_0__15 ;
    assign d_arr_9__29 = d_arr_0__15 ;
    assign d_arr_9__28 = d_arr_0__15 ;
    assign d_arr_9__27 = d_arr_0__15 ;
    assign d_arr_9__26 = d_arr_0__15 ;
    assign d_arr_9__25 = d_arr_0__15 ;
    assign d_arr_9__24 = d_arr_0__15 ;
    assign d_arr_9__23 = d_arr_0__15 ;
    assign d_arr_9__22 = d_arr_0__15 ;
    assign d_arr_9__21 = d_arr_0__15 ;
    assign d_arr_9__20 = d_arr_0__15 ;
    assign d_arr_9__19 = d_arr_0__15 ;
    assign d_arr_9__18 = d_arr_0__15 ;
    assign d_arr_9__17 = d_arr_0__15 ;
    assign d_arr_9__16 = d_arr_0__15 ;
    assign d_arr_9__15 = d_arr_0__15 ;
    assign d_arr_9__14 = d_arr_0__15 ;
    assign d_arr_9__13 = d_arr_0__15 ;
    assign d_arr_9__12 = d_arr_0__15 ;
    assign d_arr_9__11 = d_arr_0__15 ;
    assign d_arr_9__10 = d_arr_0__15 ;
    assign d_arr_9__9 = d_arr_0__15 ;
    assign d_arr_9__8 = d_arr_0__15 ;
    assign d_arr_9__7 = d_arr_0__15 ;
    assign d_arr_9__6 = d_arr_0__15 ;
    assign d_arr_9__5 = d_arr_0__15 ;
    assign d_arr_9__4 = d_arr_0__15 ;
    assign d_arr_9__3 = d_arr_0__15 ;
    assign d_arr_9__2 = d_arr_0__15 ;
    assign d_arr_9__1 = d_arr_0__15 ;
    assign d_arr_9__0 = d_arr_0__15 ;
    assign d_arr_10__31 = d_arr_0__15 ;
    assign d_arr_10__30 = d_arr_0__15 ;
    assign d_arr_10__29 = d_arr_0__15 ;
    assign d_arr_10__28 = d_arr_0__15 ;
    assign d_arr_10__27 = d_arr_0__15 ;
    assign d_arr_10__26 = d_arr_0__15 ;
    assign d_arr_10__25 = d_arr_0__15 ;
    assign d_arr_10__24 = d_arr_0__15 ;
    assign d_arr_10__23 = d_arr_0__15 ;
    assign d_arr_10__22 = d_arr_0__15 ;
    assign d_arr_10__21 = d_arr_0__15 ;
    assign d_arr_10__20 = d_arr_0__15 ;
    assign d_arr_10__19 = d_arr_0__15 ;
    assign d_arr_10__18 = d_arr_0__15 ;
    assign d_arr_10__17 = d_arr_0__15 ;
    assign d_arr_10__16 = d_arr_0__15 ;
    assign d_arr_10__15 = d_arr_0__15 ;
    assign d_arr_10__14 = d_arr_0__15 ;
    assign d_arr_10__13 = d_arr_0__15 ;
    assign d_arr_10__12 = d_arr_0__15 ;
    assign d_arr_10__11 = d_arr_0__15 ;
    assign d_arr_10__10 = d_arr_0__15 ;
    assign d_arr_10__9 = d_arr_0__15 ;
    assign d_arr_10__8 = d_arr_0__15 ;
    assign d_arr_10__7 = d_arr_0__15 ;
    assign d_arr_10__6 = d_arr_0__15 ;
    assign d_arr_10__5 = d_arr_0__15 ;
    assign d_arr_10__4 = d_arr_0__15 ;
    assign d_arr_10__3 = d_arr_0__15 ;
    assign d_arr_10__2 = d_arr_0__15 ;
    assign d_arr_10__1 = d_arr_0__15 ;
    assign d_arr_10__0 = d_arr_0__15 ;
    assign d_arr_11__31 = d_arr_0__15 ;
    assign d_arr_11__30 = d_arr_0__15 ;
    assign d_arr_11__29 = d_arr_0__15 ;
    assign d_arr_11__28 = d_arr_0__15 ;
    assign d_arr_11__27 = d_arr_0__15 ;
    assign d_arr_11__26 = d_arr_0__15 ;
    assign d_arr_11__25 = d_arr_0__15 ;
    assign d_arr_11__24 = d_arr_0__15 ;
    assign d_arr_11__23 = d_arr_0__15 ;
    assign d_arr_11__22 = d_arr_0__15 ;
    assign d_arr_11__21 = d_arr_0__15 ;
    assign d_arr_11__20 = d_arr_0__15 ;
    assign d_arr_11__19 = d_arr_0__15 ;
    assign d_arr_11__18 = d_arr_0__15 ;
    assign d_arr_11__17 = d_arr_0__15 ;
    assign d_arr_11__16 = d_arr_0__15 ;
    assign d_arr_11__15 = d_arr_0__15 ;
    assign d_arr_11__14 = d_arr_0__15 ;
    assign d_arr_11__13 = d_arr_0__15 ;
    assign d_arr_11__12 = d_arr_0__15 ;
    assign d_arr_11__11 = d_arr_0__15 ;
    assign d_arr_11__10 = d_arr_0__15 ;
    assign d_arr_11__9 = d_arr_0__15 ;
    assign d_arr_11__8 = d_arr_0__15 ;
    assign d_arr_11__7 = d_arr_0__15 ;
    assign d_arr_11__6 = d_arr_0__15 ;
    assign d_arr_11__5 = d_arr_0__15 ;
    assign d_arr_11__4 = d_arr_0__15 ;
    assign d_arr_11__3 = d_arr_0__15 ;
    assign d_arr_11__2 = d_arr_0__15 ;
    assign d_arr_11__1 = d_arr_0__15 ;
    assign d_arr_11__0 = d_arr_0__15 ;
    assign d_arr_12__31 = d_arr_0__15 ;
    assign d_arr_12__30 = d_arr_0__15 ;
    assign d_arr_12__29 = d_arr_0__15 ;
    assign d_arr_12__28 = d_arr_0__15 ;
    assign d_arr_12__27 = d_arr_0__15 ;
    assign d_arr_12__26 = d_arr_0__15 ;
    assign d_arr_12__25 = d_arr_0__15 ;
    assign d_arr_12__24 = d_arr_0__15 ;
    assign d_arr_12__23 = d_arr_0__15 ;
    assign d_arr_12__22 = d_arr_0__15 ;
    assign d_arr_12__21 = d_arr_0__15 ;
    assign d_arr_12__20 = d_arr_0__15 ;
    assign d_arr_12__19 = d_arr_0__15 ;
    assign d_arr_12__18 = d_arr_0__15 ;
    assign d_arr_12__17 = d_arr_0__15 ;
    assign d_arr_12__16 = d_arr_0__15 ;
    assign d_arr_12__15 = d_arr_0__15 ;
    assign d_arr_12__14 = d_arr_0__15 ;
    assign d_arr_12__13 = d_arr_0__15 ;
    assign d_arr_12__12 = d_arr_0__15 ;
    assign d_arr_12__11 = d_arr_0__15 ;
    assign d_arr_12__10 = d_arr_0__15 ;
    assign d_arr_12__9 = d_arr_0__15 ;
    assign d_arr_12__8 = d_arr_0__15 ;
    assign d_arr_12__7 = d_arr_0__15 ;
    assign d_arr_12__6 = d_arr_0__15 ;
    assign d_arr_12__5 = d_arr_0__15 ;
    assign d_arr_12__4 = d_arr_0__15 ;
    assign d_arr_12__3 = d_arr_0__15 ;
    assign d_arr_12__2 = d_arr_0__15 ;
    assign d_arr_12__1 = d_arr_0__15 ;
    assign d_arr_12__0 = d_arr_0__15 ;
    assign d_arr_13__31 = d_arr_0__15 ;
    assign d_arr_13__30 = d_arr_0__15 ;
    assign d_arr_13__29 = d_arr_0__15 ;
    assign d_arr_13__28 = d_arr_0__15 ;
    assign d_arr_13__27 = d_arr_0__15 ;
    assign d_arr_13__26 = d_arr_0__15 ;
    assign d_arr_13__25 = d_arr_0__15 ;
    assign d_arr_13__24 = d_arr_0__15 ;
    assign d_arr_13__23 = d_arr_0__15 ;
    assign d_arr_13__22 = d_arr_0__15 ;
    assign d_arr_13__21 = d_arr_0__15 ;
    assign d_arr_13__20 = d_arr_0__15 ;
    assign d_arr_13__19 = d_arr_0__15 ;
    assign d_arr_13__18 = d_arr_0__15 ;
    assign d_arr_13__17 = d_arr_0__15 ;
    assign d_arr_13__16 = d_arr_0__15 ;
    assign d_arr_13__15 = d_arr_0__15 ;
    assign d_arr_13__14 = d_arr_0__15 ;
    assign d_arr_13__13 = d_arr_0__15 ;
    assign d_arr_13__12 = d_arr_0__15 ;
    assign d_arr_13__11 = d_arr_0__15 ;
    assign d_arr_13__10 = d_arr_0__15 ;
    assign d_arr_13__9 = d_arr_0__15 ;
    assign d_arr_13__8 = d_arr_0__15 ;
    assign d_arr_13__7 = d_arr_0__15 ;
    assign d_arr_13__6 = d_arr_0__15 ;
    assign d_arr_13__5 = d_arr_0__15 ;
    assign d_arr_13__4 = d_arr_0__15 ;
    assign d_arr_13__3 = d_arr_0__15 ;
    assign d_arr_13__2 = d_arr_0__15 ;
    assign d_arr_13__1 = d_arr_0__15 ;
    assign d_arr_13__0 = d_arr_0__15 ;
    assign d_arr_14__31 = d_arr_0__15 ;
    assign d_arr_14__30 = d_arr_0__15 ;
    assign d_arr_14__29 = d_arr_0__15 ;
    assign d_arr_14__28 = d_arr_0__15 ;
    assign d_arr_14__27 = d_arr_0__15 ;
    assign d_arr_14__26 = d_arr_0__15 ;
    assign d_arr_14__25 = d_arr_0__15 ;
    assign d_arr_14__24 = d_arr_0__15 ;
    assign d_arr_14__23 = d_arr_0__15 ;
    assign d_arr_14__22 = d_arr_0__15 ;
    assign d_arr_14__21 = d_arr_0__15 ;
    assign d_arr_14__20 = d_arr_0__15 ;
    assign d_arr_14__19 = d_arr_0__15 ;
    assign d_arr_14__18 = d_arr_0__15 ;
    assign d_arr_14__17 = d_arr_0__15 ;
    assign d_arr_14__16 = d_arr_0__15 ;
    assign d_arr_14__15 = d_arr_0__15 ;
    assign d_arr_14__14 = d_arr_0__15 ;
    assign d_arr_14__13 = d_arr_0__15 ;
    assign d_arr_14__12 = d_arr_0__15 ;
    assign d_arr_14__11 = d_arr_0__15 ;
    assign d_arr_14__10 = d_arr_0__15 ;
    assign d_arr_14__9 = d_arr_0__15 ;
    assign d_arr_14__8 = d_arr_0__15 ;
    assign d_arr_14__7 = d_arr_0__15 ;
    assign d_arr_14__6 = d_arr_0__15 ;
    assign d_arr_14__5 = d_arr_0__15 ;
    assign d_arr_14__4 = d_arr_0__15 ;
    assign d_arr_14__3 = d_arr_0__15 ;
    assign d_arr_14__2 = d_arr_0__15 ;
    assign d_arr_14__1 = d_arr_0__15 ;
    assign d_arr_14__0 = d_arr_0__15 ;
    assign d_arr_15__31 = d_arr_0__15 ;
    assign d_arr_15__30 = d_arr_0__15 ;
    assign d_arr_15__29 = d_arr_0__15 ;
    assign d_arr_15__28 = d_arr_0__15 ;
    assign d_arr_15__27 = d_arr_0__15 ;
    assign d_arr_15__26 = d_arr_0__15 ;
    assign d_arr_15__25 = d_arr_0__15 ;
    assign d_arr_15__24 = d_arr_0__15 ;
    assign d_arr_15__23 = d_arr_0__15 ;
    assign d_arr_15__22 = d_arr_0__15 ;
    assign d_arr_15__21 = d_arr_0__15 ;
    assign d_arr_15__20 = d_arr_0__15 ;
    assign d_arr_15__19 = d_arr_0__15 ;
    assign d_arr_15__18 = d_arr_0__15 ;
    assign d_arr_15__17 = d_arr_0__15 ;
    assign d_arr_15__16 = d_arr_0__15 ;
    assign d_arr_15__15 = d_arr_0__15 ;
    assign d_arr_15__14 = d_arr_0__15 ;
    assign d_arr_15__13 = d_arr_0__15 ;
    assign d_arr_15__12 = d_arr_0__15 ;
    assign d_arr_15__11 = d_arr_0__15 ;
    assign d_arr_15__10 = d_arr_0__15 ;
    assign d_arr_15__9 = d_arr_0__15 ;
    assign d_arr_15__8 = d_arr_0__15 ;
    assign d_arr_15__7 = d_arr_0__15 ;
    assign d_arr_15__6 = d_arr_0__15 ;
    assign d_arr_15__5 = d_arr_0__15 ;
    assign d_arr_15__4 = d_arr_0__15 ;
    assign d_arr_15__3 = d_arr_0__15 ;
    assign d_arr_15__2 = d_arr_0__15 ;
    assign d_arr_15__1 = d_arr_0__15 ;
    assign d_arr_15__0 = d_arr_0__15 ;
    assign d_arr_16__31 = d_arr_0__15 ;
    assign d_arr_16__30 = d_arr_0__15 ;
    assign d_arr_16__29 = d_arr_0__15 ;
    assign d_arr_16__28 = d_arr_0__15 ;
    assign d_arr_16__27 = d_arr_0__15 ;
    assign d_arr_16__26 = d_arr_0__15 ;
    assign d_arr_16__25 = d_arr_0__15 ;
    assign d_arr_16__24 = d_arr_0__15 ;
    assign d_arr_16__23 = d_arr_0__15 ;
    assign d_arr_16__22 = d_arr_0__15 ;
    assign d_arr_16__21 = d_arr_0__15 ;
    assign d_arr_16__20 = d_arr_0__15 ;
    assign d_arr_16__19 = d_arr_0__15 ;
    assign d_arr_16__18 = d_arr_0__15 ;
    assign d_arr_16__17 = d_arr_0__15 ;
    assign d_arr_16__16 = d_arr_0__15 ;
    assign d_arr_16__15 = d_arr_0__15 ;
    assign d_arr_16__14 = d_arr_0__15 ;
    assign d_arr_16__13 = d_arr_0__15 ;
    assign d_arr_16__12 = d_arr_0__15 ;
    assign d_arr_16__11 = d_arr_0__15 ;
    assign d_arr_16__10 = d_arr_0__15 ;
    assign d_arr_16__9 = d_arr_0__15 ;
    assign d_arr_16__8 = d_arr_0__15 ;
    assign d_arr_16__7 = d_arr_0__15 ;
    assign d_arr_16__6 = d_arr_0__15 ;
    assign d_arr_16__5 = d_arr_0__15 ;
    assign d_arr_16__4 = d_arr_0__15 ;
    assign d_arr_16__3 = d_arr_0__15 ;
    assign d_arr_16__2 = d_arr_0__15 ;
    assign d_arr_16__1 = d_arr_0__15 ;
    assign d_arr_16__0 = d_arr_0__15 ;
    assign d_arr_17__31 = d_arr_0__15 ;
    assign d_arr_17__30 = d_arr_0__15 ;
    assign d_arr_17__29 = d_arr_0__15 ;
    assign d_arr_17__28 = d_arr_0__15 ;
    assign d_arr_17__27 = d_arr_0__15 ;
    assign d_arr_17__26 = d_arr_0__15 ;
    assign d_arr_17__25 = d_arr_0__15 ;
    assign d_arr_17__24 = d_arr_0__15 ;
    assign d_arr_17__23 = d_arr_0__15 ;
    assign d_arr_17__22 = d_arr_0__15 ;
    assign d_arr_17__21 = d_arr_0__15 ;
    assign d_arr_17__20 = d_arr_0__15 ;
    assign d_arr_17__19 = d_arr_0__15 ;
    assign d_arr_17__18 = d_arr_0__15 ;
    assign d_arr_17__17 = d_arr_0__15 ;
    assign d_arr_17__16 = d_arr_0__15 ;
    assign d_arr_17__15 = d_arr_0__15 ;
    assign d_arr_17__14 = d_arr_0__15 ;
    assign d_arr_17__13 = d_arr_0__15 ;
    assign d_arr_17__12 = d_arr_0__15 ;
    assign d_arr_17__11 = d_arr_0__15 ;
    assign d_arr_17__10 = d_arr_0__15 ;
    assign d_arr_17__9 = d_arr_0__15 ;
    assign d_arr_17__8 = d_arr_0__15 ;
    assign d_arr_17__7 = d_arr_0__15 ;
    assign d_arr_17__6 = d_arr_0__15 ;
    assign d_arr_17__5 = d_arr_0__15 ;
    assign d_arr_17__4 = d_arr_0__15 ;
    assign d_arr_17__3 = d_arr_0__15 ;
    assign d_arr_17__2 = d_arr_0__15 ;
    assign d_arr_17__1 = d_arr_0__15 ;
    assign d_arr_17__0 = d_arr_0__15 ;
    assign d_arr_18__31 = d_arr_0__15 ;
    assign d_arr_18__30 = d_arr_0__15 ;
    assign d_arr_18__29 = d_arr_0__15 ;
    assign d_arr_18__28 = d_arr_0__15 ;
    assign d_arr_18__27 = d_arr_0__15 ;
    assign d_arr_18__26 = d_arr_0__15 ;
    assign d_arr_18__25 = d_arr_0__15 ;
    assign d_arr_18__24 = d_arr_0__15 ;
    assign d_arr_18__23 = d_arr_0__15 ;
    assign d_arr_18__22 = d_arr_0__15 ;
    assign d_arr_18__21 = d_arr_0__15 ;
    assign d_arr_18__20 = d_arr_0__15 ;
    assign d_arr_18__19 = d_arr_0__15 ;
    assign d_arr_18__18 = d_arr_0__15 ;
    assign d_arr_18__17 = d_arr_0__15 ;
    assign d_arr_18__16 = d_arr_0__15 ;
    assign d_arr_18__15 = d_arr_0__15 ;
    assign d_arr_18__14 = d_arr_0__15 ;
    assign d_arr_18__13 = d_arr_0__15 ;
    assign d_arr_18__12 = d_arr_0__15 ;
    assign d_arr_18__11 = d_arr_0__15 ;
    assign d_arr_18__10 = d_arr_0__15 ;
    assign d_arr_18__9 = d_arr_0__15 ;
    assign d_arr_18__8 = d_arr_0__15 ;
    assign d_arr_18__7 = d_arr_0__15 ;
    assign d_arr_18__6 = d_arr_0__15 ;
    assign d_arr_18__5 = d_arr_0__15 ;
    assign d_arr_18__4 = d_arr_0__15 ;
    assign d_arr_18__3 = d_arr_0__15 ;
    assign d_arr_18__2 = d_arr_0__15 ;
    assign d_arr_18__1 = d_arr_0__15 ;
    assign d_arr_18__0 = d_arr_0__15 ;
    assign d_arr_19__31 = d_arr_0__15 ;
    assign d_arr_19__30 = d_arr_0__15 ;
    assign d_arr_19__29 = d_arr_0__15 ;
    assign d_arr_19__28 = d_arr_0__15 ;
    assign d_arr_19__27 = d_arr_0__15 ;
    assign d_arr_19__26 = d_arr_0__15 ;
    assign d_arr_19__25 = d_arr_0__15 ;
    assign d_arr_19__24 = d_arr_0__15 ;
    assign d_arr_19__23 = d_arr_0__15 ;
    assign d_arr_19__22 = d_arr_0__15 ;
    assign d_arr_19__21 = d_arr_0__15 ;
    assign d_arr_19__20 = d_arr_0__15 ;
    assign d_arr_19__19 = d_arr_0__15 ;
    assign d_arr_19__18 = d_arr_0__15 ;
    assign d_arr_19__17 = d_arr_0__15 ;
    assign d_arr_19__16 = d_arr_0__15 ;
    assign d_arr_19__15 = d_arr_0__15 ;
    assign d_arr_19__14 = d_arr_0__15 ;
    assign d_arr_19__13 = d_arr_0__15 ;
    assign d_arr_19__12 = d_arr_0__15 ;
    assign d_arr_19__11 = d_arr_0__15 ;
    assign d_arr_19__10 = d_arr_0__15 ;
    assign d_arr_19__9 = d_arr_0__15 ;
    assign d_arr_19__8 = d_arr_0__15 ;
    assign d_arr_19__7 = d_arr_0__15 ;
    assign d_arr_19__6 = d_arr_0__15 ;
    assign d_arr_19__5 = d_arr_0__15 ;
    assign d_arr_19__4 = d_arr_0__15 ;
    assign d_arr_19__3 = d_arr_0__15 ;
    assign d_arr_19__2 = d_arr_0__15 ;
    assign d_arr_19__1 = d_arr_0__15 ;
    assign d_arr_19__0 = d_arr_0__15 ;
    assign d_arr_20__31 = d_arr_0__15 ;
    assign d_arr_20__30 = d_arr_0__15 ;
    assign d_arr_20__29 = d_arr_0__15 ;
    assign d_arr_20__28 = d_arr_0__15 ;
    assign d_arr_20__27 = d_arr_0__15 ;
    assign d_arr_20__26 = d_arr_0__15 ;
    assign d_arr_20__25 = d_arr_0__15 ;
    assign d_arr_20__24 = d_arr_0__15 ;
    assign d_arr_20__23 = d_arr_0__15 ;
    assign d_arr_20__22 = d_arr_0__15 ;
    assign d_arr_20__21 = d_arr_0__15 ;
    assign d_arr_20__20 = d_arr_0__15 ;
    assign d_arr_20__19 = d_arr_0__15 ;
    assign d_arr_20__18 = d_arr_0__15 ;
    assign d_arr_20__17 = d_arr_0__15 ;
    assign d_arr_20__16 = d_arr_0__15 ;
    assign d_arr_20__15 = d_arr_0__15 ;
    assign d_arr_20__14 = d_arr_0__15 ;
    assign d_arr_20__13 = d_arr_0__15 ;
    assign d_arr_20__12 = d_arr_0__15 ;
    assign d_arr_20__11 = d_arr_0__15 ;
    assign d_arr_20__10 = d_arr_0__15 ;
    assign d_arr_20__9 = d_arr_0__15 ;
    assign d_arr_20__8 = d_arr_0__15 ;
    assign d_arr_20__7 = d_arr_0__15 ;
    assign d_arr_20__6 = d_arr_0__15 ;
    assign d_arr_20__5 = d_arr_0__15 ;
    assign d_arr_20__4 = d_arr_0__15 ;
    assign d_arr_20__3 = d_arr_0__15 ;
    assign d_arr_20__2 = d_arr_0__15 ;
    assign d_arr_20__1 = d_arr_0__15 ;
    assign d_arr_20__0 = d_arr_0__15 ;
    assign d_arr_21__31 = d_arr_0__15 ;
    assign d_arr_21__30 = d_arr_0__15 ;
    assign d_arr_21__29 = d_arr_0__15 ;
    assign d_arr_21__28 = d_arr_0__15 ;
    assign d_arr_21__27 = d_arr_0__15 ;
    assign d_arr_21__26 = d_arr_0__15 ;
    assign d_arr_21__25 = d_arr_0__15 ;
    assign d_arr_21__24 = d_arr_0__15 ;
    assign d_arr_21__23 = d_arr_0__15 ;
    assign d_arr_21__22 = d_arr_0__15 ;
    assign d_arr_21__21 = d_arr_0__15 ;
    assign d_arr_21__20 = d_arr_0__15 ;
    assign d_arr_21__19 = d_arr_0__15 ;
    assign d_arr_21__18 = d_arr_0__15 ;
    assign d_arr_21__17 = d_arr_0__15 ;
    assign d_arr_21__16 = d_arr_0__15 ;
    assign d_arr_21__15 = d_arr_0__15 ;
    assign d_arr_21__14 = d_arr_0__15 ;
    assign d_arr_21__13 = d_arr_0__15 ;
    assign d_arr_21__12 = d_arr_0__15 ;
    assign d_arr_21__11 = d_arr_0__15 ;
    assign d_arr_21__10 = d_arr_0__15 ;
    assign d_arr_21__9 = d_arr_0__15 ;
    assign d_arr_21__8 = d_arr_0__15 ;
    assign d_arr_21__7 = d_arr_0__15 ;
    assign d_arr_21__6 = d_arr_0__15 ;
    assign d_arr_21__5 = d_arr_0__15 ;
    assign d_arr_21__4 = d_arr_0__15 ;
    assign d_arr_21__3 = d_arr_0__15 ;
    assign d_arr_21__2 = d_arr_0__15 ;
    assign d_arr_21__1 = d_arr_0__15 ;
    assign d_arr_21__0 = d_arr_0__15 ;
    assign d_arr_22__31 = d_arr_0__15 ;
    assign d_arr_22__30 = d_arr_0__15 ;
    assign d_arr_22__29 = d_arr_0__15 ;
    assign d_arr_22__28 = d_arr_0__15 ;
    assign d_arr_22__27 = d_arr_0__15 ;
    assign d_arr_22__26 = d_arr_0__15 ;
    assign d_arr_22__25 = d_arr_0__15 ;
    assign d_arr_22__24 = d_arr_0__15 ;
    assign d_arr_22__23 = d_arr_0__15 ;
    assign d_arr_22__22 = d_arr_0__15 ;
    assign d_arr_22__21 = d_arr_0__15 ;
    assign d_arr_22__20 = d_arr_0__15 ;
    assign d_arr_22__19 = d_arr_0__15 ;
    assign d_arr_22__18 = d_arr_0__15 ;
    assign d_arr_22__17 = d_arr_0__15 ;
    assign d_arr_22__16 = d_arr_0__15 ;
    assign d_arr_22__15 = d_arr_0__15 ;
    assign d_arr_22__14 = d_arr_0__15 ;
    assign d_arr_22__13 = d_arr_0__15 ;
    assign d_arr_22__12 = d_arr_0__15 ;
    assign d_arr_22__11 = d_arr_0__15 ;
    assign d_arr_22__10 = d_arr_0__15 ;
    assign d_arr_22__9 = d_arr_0__15 ;
    assign d_arr_22__8 = d_arr_0__15 ;
    assign d_arr_22__7 = d_arr_0__15 ;
    assign d_arr_22__6 = d_arr_0__15 ;
    assign d_arr_22__5 = d_arr_0__15 ;
    assign d_arr_22__4 = d_arr_0__15 ;
    assign d_arr_22__3 = d_arr_0__15 ;
    assign d_arr_22__2 = d_arr_0__15 ;
    assign d_arr_22__1 = d_arr_0__15 ;
    assign d_arr_22__0 = d_arr_0__15 ;
    assign d_arr_23__31 = d_arr_0__15 ;
    assign d_arr_23__30 = d_arr_0__15 ;
    assign d_arr_23__29 = d_arr_0__15 ;
    assign d_arr_23__28 = d_arr_0__15 ;
    assign d_arr_23__27 = d_arr_0__15 ;
    assign d_arr_23__26 = d_arr_0__15 ;
    assign d_arr_23__25 = d_arr_0__15 ;
    assign d_arr_23__24 = d_arr_0__15 ;
    assign d_arr_23__23 = d_arr_0__15 ;
    assign d_arr_23__22 = d_arr_0__15 ;
    assign d_arr_23__21 = d_arr_0__15 ;
    assign d_arr_23__20 = d_arr_0__15 ;
    assign d_arr_23__19 = d_arr_0__15 ;
    assign d_arr_23__18 = d_arr_0__15 ;
    assign d_arr_23__17 = d_arr_0__15 ;
    assign d_arr_23__16 = d_arr_0__15 ;
    assign d_arr_23__15 = d_arr_0__15 ;
    assign d_arr_23__14 = d_arr_0__15 ;
    assign d_arr_23__13 = d_arr_0__15 ;
    assign d_arr_23__12 = d_arr_0__15 ;
    assign d_arr_23__11 = d_arr_0__15 ;
    assign d_arr_23__10 = d_arr_0__15 ;
    assign d_arr_23__9 = d_arr_0__15 ;
    assign d_arr_23__8 = d_arr_0__15 ;
    assign d_arr_23__7 = d_arr_0__15 ;
    assign d_arr_23__6 = d_arr_0__15 ;
    assign d_arr_23__5 = d_arr_0__15 ;
    assign d_arr_23__4 = d_arr_0__15 ;
    assign d_arr_23__3 = d_arr_0__15 ;
    assign d_arr_23__2 = d_arr_0__15 ;
    assign d_arr_23__1 = d_arr_0__15 ;
    assign d_arr_23__0 = d_arr_0__15 ;
    assign d_arr_24__31 = d_arr_0__15 ;
    assign d_arr_24__30 = d_arr_0__15 ;
    assign d_arr_24__29 = d_arr_0__15 ;
    assign d_arr_24__28 = d_arr_0__15 ;
    assign d_arr_24__27 = d_arr_0__15 ;
    assign d_arr_24__26 = d_arr_0__15 ;
    assign d_arr_24__25 = d_arr_0__15 ;
    assign d_arr_24__24 = d_arr_0__15 ;
    assign d_arr_24__23 = d_arr_0__15 ;
    assign d_arr_24__22 = d_arr_0__15 ;
    assign d_arr_24__21 = d_arr_0__15 ;
    assign d_arr_24__20 = d_arr_0__15 ;
    assign d_arr_24__19 = d_arr_0__15 ;
    assign d_arr_24__18 = d_arr_0__15 ;
    assign d_arr_24__17 = d_arr_0__15 ;
    assign d_arr_24__16 = d_arr_0__15 ;
    assign d_arr_24__15 = d_arr_0__15 ;
    assign d_arr_24__14 = d_arr_0__15 ;
    assign d_arr_24__13 = d_arr_0__15 ;
    assign d_arr_24__12 = d_arr_0__15 ;
    assign d_arr_24__11 = d_arr_0__15 ;
    assign d_arr_24__10 = d_arr_0__15 ;
    assign d_arr_24__9 = d_arr_0__15 ;
    assign d_arr_24__8 = d_arr_0__15 ;
    assign d_arr_24__7 = d_arr_0__15 ;
    assign d_arr_24__6 = d_arr_0__15 ;
    assign d_arr_24__5 = d_arr_0__15 ;
    assign d_arr_24__4 = d_arr_0__15 ;
    assign d_arr_24__3 = d_arr_0__15 ;
    assign d_arr_24__2 = d_arr_0__15 ;
    assign d_arr_24__1 = d_arr_0__15 ;
    assign d_arr_24__0 = d_arr_0__15 ;
    fake_gnd ix42 (.Y (d_arr_0__15)) ;
    nor02ii ix3 (.Y (d_arr_1__0), .A0 (nx219), .A1 (q_arr_1__0)) ;
    nor02ii ix7 (.Y (d_arr_1__1), .A0 (nx219), .A1 (q_arr_1__1)) ;
    nor02ii ix11 (.Y (d_arr_1__2), .A0 (nx219), .A1 (q_arr_1__2)) ;
    nor02ii ix15 (.Y (d_arr_1__3), .A0 (nx219), .A1 (q_arr_1__3)) ;
    nor02ii ix19 (.Y (d_arr_1__4), .A0 (nx219), .A1 (q_arr_1__4)) ;
    nor02ii ix23 (.Y (d_arr_1__5), .A0 (nx219), .A1 (q_arr_1__5)) ;
    nor02ii ix27 (.Y (d_arr_1__6), .A0 (nx219), .A1 (q_arr_1__6)) ;
    nor02ii ix31 (.Y (d_arr_1__7), .A0 (nx221), .A1 (q_arr_1__7)) ;
    nor02ii ix35 (.Y (d_arr_1__8), .A0 (nx221), .A1 (q_arr_1__8)) ;
    nor02ii ix39 (.Y (d_arr_1__9), .A0 (nx221), .A1 (q_arr_1__9)) ;
    nor02ii ix43 (.Y (d_arr_1__10), .A0 (nx221), .A1 (q_arr_1__10)) ;
    nor02ii ix47 (.Y (d_arr_1__11), .A0 (nx221), .A1 (q_arr_1__11)) ;
    nor02ii ix51 (.Y (d_arr_1__12), .A0 (nx221), .A1 (q_arr_1__12)) ;
    nor02ii ix55 (.Y (d_arr_1__13), .A0 (nx221), .A1 (q_arr_1__13)) ;
    nor02ii ix59 (.Y (d_arr_1__14), .A0 (nx223), .A1 (q_arr_1__14)) ;
    nor02ii ix63 (.Y (d_arr_1__16), .A0 (nx223), .A1 (q_arr_1__16)) ;
    nor02ii ix67 (.Y (d_arr_1__17), .A0 (nx223), .A1 (q_arr_1__17)) ;
    nor02ii ix71 (.Y (d_arr_1__18), .A0 (nx223), .A1 (q_arr_1__18)) ;
    nor02ii ix75 (.Y (d_arr_1__19), .A0 (nx223), .A1 (q_arr_1__19)) ;
    nor02ii ix79 (.Y (d_arr_1__20), .A0 (nx223), .A1 (q_arr_1__20)) ;
    nor02ii ix83 (.Y (d_arr_1__21), .A0 (nx223), .A1 (q_arr_1__21)) ;
    nor02ii ix87 (.Y (d_arr_1__22), .A0 (nx225), .A1 (q_arr_1__22)) ;
    nor02ii ix91 (.Y (d_arr_1__23), .A0 (nx225), .A1 (q_arr_1__23)) ;
    nor02ii ix95 (.Y (d_arr_1__24), .A0 (nx225), .A1 (q_arr_1__24)) ;
    nor02ii ix99 (.Y (d_arr_1__25), .A0 (nx225), .A1 (q_arr_1__25)) ;
    nor02ii ix103 (.Y (d_arr_1__26), .A0 (nx225), .A1 (q_arr_1__26)) ;
    nor02ii ix107 (.Y (d_arr_1__27), .A0 (nx225), .A1 (q_arr_1__27)) ;
    nor02ii ix111 (.Y (d_arr_1__28), .A0 (nx225), .A1 (q_arr_1__28)) ;
    nor02ii ix115 (.Y (d_arr_1__29), .A0 (nx227), .A1 (q_arr_1__29)) ;
    nor02ii ix119 (.Y (d_arr_1__30), .A0 (nx227), .A1 (q_arr_1__30)) ;
    nor02ii ix123 (.Y (d_arr_1__31), .A0 (nx227), .A1 (q_arr_1__31)) ;
    nor02ii ix127 (.Y (d_arr_0__0), .A0 (nx207), .A1 (q_arr_0__0)) ;
    nor02ii ix131 (.Y (d_arr_0__1), .A0 (nx207), .A1 (q_arr_0__1)) ;
    nor02ii ix135 (.Y (d_arr_0__2), .A0 (nx207), .A1 (q_arr_0__2)) ;
    nor02ii ix139 (.Y (d_arr_0__3), .A0 (nx207), .A1 (q_arr_0__3)) ;
    nor02ii ix143 (.Y (d_arr_0__4), .A0 (nx207), .A1 (q_arr_0__4)) ;
    nor02ii ix147 (.Y (d_arr_0__5), .A0 (nx207), .A1 (q_arr_0__5)) ;
    nor02ii ix151 (.Y (d_arr_0__6), .A0 (nx207), .A1 (q_arr_0__6)) ;
    nor02ii ix155 (.Y (d_arr_0__7), .A0 (nx209), .A1 (q_arr_0__7)) ;
    nor02ii ix159 (.Y (d_arr_0__8), .A0 (nx209), .A1 (q_arr_0__8)) ;
    nor02ii ix163 (.Y (d_arr_0__9), .A0 (nx209), .A1 (q_arr_0__9)) ;
    nor02ii ix167 (.Y (d_arr_0__10), .A0 (nx209), .A1 (q_arr_0__10)) ;
    nor02ii ix171 (.Y (d_arr_0__11), .A0 (nx209), .A1 (q_arr_0__11)) ;
    nor02ii ix175 (.Y (d_arr_0__12), .A0 (nx209), .A1 (q_arr_0__12)) ;
    nor02ii ix179 (.Y (d_arr_0__13), .A0 (nx209), .A1 (q_arr_0__13)) ;
    nor02ii ix183 (.Y (d_arr_0__14), .A0 (nx211), .A1 (q_arr_0__14)) ;
    nor02ii ix187 (.Y (d_arr_0__16), .A0 (nx211), .A1 (q_arr_0__16)) ;
    nor02ii ix191 (.Y (d_arr_0__17), .A0 (nx211), .A1 (q_arr_0__17)) ;
    nor02ii ix195 (.Y (d_arr_0__18), .A0 (nx211), .A1 (q_arr_0__18)) ;
    nor02ii ix199 (.Y (d_arr_0__19), .A0 (nx211), .A1 (q_arr_0__19)) ;
    nor02ii ix203 (.Y (d_arr_0__20), .A0 (nx211), .A1 (q_arr_0__20)) ;
    nor02ii ix207 (.Y (d_arr_0__21), .A0 (nx211), .A1 (q_arr_0__21)) ;
    nor02ii ix211 (.Y (d_arr_0__22), .A0 (nx213), .A1 (q_arr_0__22)) ;
    nor02ii ix215 (.Y (d_arr_0__23), .A0 (nx213), .A1 (q_arr_0__23)) ;
    nor02ii ix219 (.Y (d_arr_0__24), .A0 (nx213), .A1 (q_arr_0__24)) ;
    nor02ii ix223 (.Y (d_arr_0__25), .A0 (nx213), .A1 (q_arr_0__25)) ;
    nor02ii ix227 (.Y (d_arr_0__26), .A0 (nx213), .A1 (q_arr_0__26)) ;
    nor02ii ix231 (.Y (d_arr_0__27), .A0 (nx213), .A1 (q_arr_0__27)) ;
    nor02ii ix235 (.Y (d_arr_0__28), .A0 (nx213), .A1 (q_arr_0__28)) ;
    nor02ii ix239 (.Y (d_arr_0__29), .A0 (nx215), .A1 (q_arr_0__29)) ;
    nor02ii ix243 (.Y (d_arr_0__30), .A0 (nx215), .A1 (q_arr_0__30)) ;
    nor02ii ix247 (.Y (d_arr_0__31), .A0 (nx215), .A1 (q_arr_0__31)) ;
    inv01 ix204 (.Y (nx205), .A (q_arr_0__15)) ;
    inv01 ix206 (.Y (nx207), .A (nx205)) ;
    inv01 ix208 (.Y (nx209), .A (nx205)) ;
    inv01 ix210 (.Y (nx211), .A (nx205)) ;
    inv01 ix212 (.Y (nx213), .A (nx205)) ;
    inv01 ix214 (.Y (nx215), .A (nx205)) ;
    inv01 ix216 (.Y (nx217), .A (q_arr_1__15)) ;
    inv01 ix218 (.Y (nx219), .A (nx217)) ;
    inv01 ix220 (.Y (nx221), .A (nx217)) ;
    inv01 ix222 (.Y (nx223), .A (nx217)) ;
    inv01 ix224 (.Y (nx225), .A (nx217)) ;
    inv01 ix226 (.Y (nx227), .A (nx217)) ;
endmodule


module MergeLayer ( d_arr_0__31, d_arr_0__30, d_arr_0__29, d_arr_0__28, 
                    d_arr_0__27, d_arr_0__26, d_arr_0__25, d_arr_0__24, 
                    d_arr_0__23, d_arr_0__22, d_arr_0__21, d_arr_0__20, 
                    d_arr_0__19, d_arr_0__18, d_arr_0__17, d_arr_0__16, 
                    d_arr_0__15, d_arr_0__14, d_arr_0__13, d_arr_0__12, 
                    d_arr_0__11, d_arr_0__10, d_arr_0__9, d_arr_0__8, d_arr_0__7, 
                    d_arr_0__6, d_arr_0__5, d_arr_0__4, d_arr_0__3, d_arr_0__2, 
                    d_arr_0__1, d_arr_0__0, d_arr_1__31, d_arr_1__30, 
                    d_arr_1__29, d_arr_1__28, d_arr_1__27, d_arr_1__26, 
                    d_arr_1__25, d_arr_1__24, d_arr_1__23, d_arr_1__22, 
                    d_arr_1__21, d_arr_1__20, d_arr_1__19, d_arr_1__18, 
                    d_arr_1__17, d_arr_1__16, d_arr_1__15, d_arr_1__14, 
                    d_arr_1__13, d_arr_1__12, d_arr_1__11, d_arr_1__10, 
                    d_arr_1__9, d_arr_1__8, d_arr_1__7, d_arr_1__6, d_arr_1__5, 
                    d_arr_1__4, d_arr_1__3, d_arr_1__2, d_arr_1__1, d_arr_1__0, 
                    d_arr_2__31, d_arr_2__30, d_arr_2__29, d_arr_2__28, 
                    d_arr_2__27, d_arr_2__26, d_arr_2__25, d_arr_2__24, 
                    d_arr_2__23, d_arr_2__22, d_arr_2__21, d_arr_2__20, 
                    d_arr_2__19, d_arr_2__18, d_arr_2__17, d_arr_2__16, 
                    d_arr_2__15, d_arr_2__14, d_arr_2__13, d_arr_2__12, 
                    d_arr_2__11, d_arr_2__10, d_arr_2__9, d_arr_2__8, d_arr_2__7, 
                    d_arr_2__6, d_arr_2__5, d_arr_2__4, d_arr_2__3, d_arr_2__2, 
                    d_arr_2__1, d_arr_2__0, d_arr_3__31, d_arr_3__30, 
                    d_arr_3__29, d_arr_3__28, d_arr_3__27, d_arr_3__26, 
                    d_arr_3__25, d_arr_3__24, d_arr_3__23, d_arr_3__22, 
                    d_arr_3__21, d_arr_3__20, d_arr_3__19, d_arr_3__18, 
                    d_arr_3__17, d_arr_3__16, d_arr_3__15, d_arr_3__14, 
                    d_arr_3__13, d_arr_3__12, d_arr_3__11, d_arr_3__10, 
                    d_arr_3__9, d_arr_3__8, d_arr_3__7, d_arr_3__6, d_arr_3__5, 
                    d_arr_3__4, d_arr_3__3, d_arr_3__2, d_arr_3__1, d_arr_3__0, 
                    d_arr_4__31, d_arr_4__30, d_arr_4__29, d_arr_4__28, 
                    d_arr_4__27, d_arr_4__26, d_arr_4__25, d_arr_4__24, 
                    d_arr_4__23, d_arr_4__22, d_arr_4__21, d_arr_4__20, 
                    d_arr_4__19, d_arr_4__18, d_arr_4__17, d_arr_4__16, 
                    d_arr_4__15, d_arr_4__14, d_arr_4__13, d_arr_4__12, 
                    d_arr_4__11, d_arr_4__10, d_arr_4__9, d_arr_4__8, d_arr_4__7, 
                    d_arr_4__6, d_arr_4__5, d_arr_4__4, d_arr_4__3, d_arr_4__2, 
                    d_arr_4__1, d_arr_4__0, d_arr_5__31, d_arr_5__30, 
                    d_arr_5__29, d_arr_5__28, d_arr_5__27, d_arr_5__26, 
                    d_arr_5__25, d_arr_5__24, d_arr_5__23, d_arr_5__22, 
                    d_arr_5__21, d_arr_5__20, d_arr_5__19, d_arr_5__18, 
                    d_arr_5__17, d_arr_5__16, d_arr_5__15, d_arr_5__14, 
                    d_arr_5__13, d_arr_5__12, d_arr_5__11, d_arr_5__10, 
                    d_arr_5__9, d_arr_5__8, d_arr_5__7, d_arr_5__6, d_arr_5__5, 
                    d_arr_5__4, d_arr_5__3, d_arr_5__2, d_arr_5__1, d_arr_5__0, 
                    d_arr_6__31, d_arr_6__30, d_arr_6__29, d_arr_6__28, 
                    d_arr_6__27, d_arr_6__26, d_arr_6__25, d_arr_6__24, 
                    d_arr_6__23, d_arr_6__22, d_arr_6__21, d_arr_6__20, 
                    d_arr_6__19, d_arr_6__18, d_arr_6__17, d_arr_6__16, 
                    d_arr_6__15, d_arr_6__14, d_arr_6__13, d_arr_6__12, 
                    d_arr_6__11, d_arr_6__10, d_arr_6__9, d_arr_6__8, d_arr_6__7, 
                    d_arr_6__6, d_arr_6__5, d_arr_6__4, d_arr_6__3, d_arr_6__2, 
                    d_arr_6__1, d_arr_6__0, d_arr_7__31, d_arr_7__30, 
                    d_arr_7__29, d_arr_7__28, d_arr_7__27, d_arr_7__26, 
                    d_arr_7__25, d_arr_7__24, d_arr_7__23, d_arr_7__22, 
                    d_arr_7__21, d_arr_7__20, d_arr_7__19, d_arr_7__18, 
                    d_arr_7__17, d_arr_7__16, d_arr_7__15, d_arr_7__14, 
                    d_arr_7__13, d_arr_7__12, d_arr_7__11, d_arr_7__10, 
                    d_arr_7__9, d_arr_7__8, d_arr_7__7, d_arr_7__6, d_arr_7__5, 
                    d_arr_7__4, d_arr_7__3, d_arr_7__2, d_arr_7__1, d_arr_7__0, 
                    d_arr_8__31, d_arr_8__30, d_arr_8__29, d_arr_8__28, 
                    d_arr_8__27, d_arr_8__26, d_arr_8__25, d_arr_8__24, 
                    d_arr_8__23, d_arr_8__22, d_arr_8__21, d_arr_8__20, 
                    d_arr_8__19, d_arr_8__18, d_arr_8__17, d_arr_8__16, 
                    d_arr_8__15, d_arr_8__14, d_arr_8__13, d_arr_8__12, 
                    d_arr_8__11, d_arr_8__10, d_arr_8__9, d_arr_8__8, d_arr_8__7, 
                    d_arr_8__6, d_arr_8__5, d_arr_8__4, d_arr_8__3, d_arr_8__2, 
                    d_arr_8__1, d_arr_8__0, d_arr_9__31, d_arr_9__30, 
                    d_arr_9__29, d_arr_9__28, d_arr_9__27, d_arr_9__26, 
                    d_arr_9__25, d_arr_9__24, d_arr_9__23, d_arr_9__22, 
                    d_arr_9__21, d_arr_9__20, d_arr_9__19, d_arr_9__18, 
                    d_arr_9__17, d_arr_9__16, d_arr_9__15, d_arr_9__14, 
                    d_arr_9__13, d_arr_9__12, d_arr_9__11, d_arr_9__10, 
                    d_arr_9__9, d_arr_9__8, d_arr_9__7, d_arr_9__6, d_arr_9__5, 
                    d_arr_9__4, d_arr_9__3, d_arr_9__2, d_arr_9__1, d_arr_9__0, 
                    d_arr_10__31, d_arr_10__30, d_arr_10__29, d_arr_10__28, 
                    d_arr_10__27, d_arr_10__26, d_arr_10__25, d_arr_10__24, 
                    d_arr_10__23, d_arr_10__22, d_arr_10__21, d_arr_10__20, 
                    d_arr_10__19, d_arr_10__18, d_arr_10__17, d_arr_10__16, 
                    d_arr_10__15, d_arr_10__14, d_arr_10__13, d_arr_10__12, 
                    d_arr_10__11, d_arr_10__10, d_arr_10__9, d_arr_10__8, 
                    d_arr_10__7, d_arr_10__6, d_arr_10__5, d_arr_10__4, 
                    d_arr_10__3, d_arr_10__2, d_arr_10__1, d_arr_10__0, 
                    d_arr_11__31, d_arr_11__30, d_arr_11__29, d_arr_11__28, 
                    d_arr_11__27, d_arr_11__26, d_arr_11__25, d_arr_11__24, 
                    d_arr_11__23, d_arr_11__22, d_arr_11__21, d_arr_11__20, 
                    d_arr_11__19, d_arr_11__18, d_arr_11__17, d_arr_11__16, 
                    d_arr_11__15, d_arr_11__14, d_arr_11__13, d_arr_11__12, 
                    d_arr_11__11, d_arr_11__10, d_arr_11__9, d_arr_11__8, 
                    d_arr_11__7, d_arr_11__6, d_arr_11__5, d_arr_11__4, 
                    d_arr_11__3, d_arr_11__2, d_arr_11__1, d_arr_11__0, 
                    d_arr_12__31, d_arr_12__30, d_arr_12__29, d_arr_12__28, 
                    d_arr_12__27, d_arr_12__26, d_arr_12__25, d_arr_12__24, 
                    d_arr_12__23, d_arr_12__22, d_arr_12__21, d_arr_12__20, 
                    d_arr_12__19, d_arr_12__18, d_arr_12__17, d_arr_12__16, 
                    d_arr_12__15, d_arr_12__14, d_arr_12__13, d_arr_12__12, 
                    d_arr_12__11, d_arr_12__10, d_arr_12__9, d_arr_12__8, 
                    d_arr_12__7, d_arr_12__6, d_arr_12__5, d_arr_12__4, 
                    d_arr_12__3, d_arr_12__2, d_arr_12__1, d_arr_12__0, 
                    d_arr_13__31, d_arr_13__30, d_arr_13__29, d_arr_13__28, 
                    d_arr_13__27, d_arr_13__26, d_arr_13__25, d_arr_13__24, 
                    d_arr_13__23, d_arr_13__22, d_arr_13__21, d_arr_13__20, 
                    d_arr_13__19, d_arr_13__18, d_arr_13__17, d_arr_13__16, 
                    d_arr_13__15, d_arr_13__14, d_arr_13__13, d_arr_13__12, 
                    d_arr_13__11, d_arr_13__10, d_arr_13__9, d_arr_13__8, 
                    d_arr_13__7, d_arr_13__6, d_arr_13__5, d_arr_13__4, 
                    d_arr_13__3, d_arr_13__2, d_arr_13__1, d_arr_13__0, 
                    d_arr_14__31, d_arr_14__30, d_arr_14__29, d_arr_14__28, 
                    d_arr_14__27, d_arr_14__26, d_arr_14__25, d_arr_14__24, 
                    d_arr_14__23, d_arr_14__22, d_arr_14__21, d_arr_14__20, 
                    d_arr_14__19, d_arr_14__18, d_arr_14__17, d_arr_14__16, 
                    d_arr_14__15, d_arr_14__14, d_arr_14__13, d_arr_14__12, 
                    d_arr_14__11, d_arr_14__10, d_arr_14__9, d_arr_14__8, 
                    d_arr_14__7, d_arr_14__6, d_arr_14__5, d_arr_14__4, 
                    d_arr_14__3, d_arr_14__2, d_arr_14__1, d_arr_14__0, 
                    d_arr_15__31, d_arr_15__30, d_arr_15__29, d_arr_15__28, 
                    d_arr_15__27, d_arr_15__26, d_arr_15__25, d_arr_15__24, 
                    d_arr_15__23, d_arr_15__22, d_arr_15__21, d_arr_15__20, 
                    d_arr_15__19, d_arr_15__18, d_arr_15__17, d_arr_15__16, 
                    d_arr_15__15, d_arr_15__14, d_arr_15__13, d_arr_15__12, 
                    d_arr_15__11, d_arr_15__10, d_arr_15__9, d_arr_15__8, 
                    d_arr_15__7, d_arr_15__6, d_arr_15__5, d_arr_15__4, 
                    d_arr_15__3, d_arr_15__2, d_arr_15__1, d_arr_15__0, 
                    d_arr_16__31, d_arr_16__30, d_arr_16__29, d_arr_16__28, 
                    d_arr_16__27, d_arr_16__26, d_arr_16__25, d_arr_16__24, 
                    d_arr_16__23, d_arr_16__22, d_arr_16__21, d_arr_16__20, 
                    d_arr_16__19, d_arr_16__18, d_arr_16__17, d_arr_16__16, 
                    d_arr_16__15, d_arr_16__14, d_arr_16__13, d_arr_16__12, 
                    d_arr_16__11, d_arr_16__10, d_arr_16__9, d_arr_16__8, 
                    d_arr_16__7, d_arr_16__6, d_arr_16__5, d_arr_16__4, 
                    d_arr_16__3, d_arr_16__2, d_arr_16__1, d_arr_16__0, 
                    d_arr_17__31, d_arr_17__30, d_arr_17__29, d_arr_17__28, 
                    d_arr_17__27, d_arr_17__26, d_arr_17__25, d_arr_17__24, 
                    d_arr_17__23, d_arr_17__22, d_arr_17__21, d_arr_17__20, 
                    d_arr_17__19, d_arr_17__18, d_arr_17__17, d_arr_17__16, 
                    d_arr_17__15, d_arr_17__14, d_arr_17__13, d_arr_17__12, 
                    d_arr_17__11, d_arr_17__10, d_arr_17__9, d_arr_17__8, 
                    d_arr_17__7, d_arr_17__6, d_arr_17__5, d_arr_17__4, 
                    d_arr_17__3, d_arr_17__2, d_arr_17__1, d_arr_17__0, 
                    d_arr_18__31, d_arr_18__30, d_arr_18__29, d_arr_18__28, 
                    d_arr_18__27, d_arr_18__26, d_arr_18__25, d_arr_18__24, 
                    d_arr_18__23, d_arr_18__22, d_arr_18__21, d_arr_18__20, 
                    d_arr_18__19, d_arr_18__18, d_arr_18__17, d_arr_18__16, 
                    d_arr_18__15, d_arr_18__14, d_arr_18__13, d_arr_18__12, 
                    d_arr_18__11, d_arr_18__10, d_arr_18__9, d_arr_18__8, 
                    d_arr_18__7, d_arr_18__6, d_arr_18__5, d_arr_18__4, 
                    d_arr_18__3, d_arr_18__2, d_arr_18__1, d_arr_18__0, 
                    d_arr_19__31, d_arr_19__30, d_arr_19__29, d_arr_19__28, 
                    d_arr_19__27, d_arr_19__26, d_arr_19__25, d_arr_19__24, 
                    d_arr_19__23, d_arr_19__22, d_arr_19__21, d_arr_19__20, 
                    d_arr_19__19, d_arr_19__18, d_arr_19__17, d_arr_19__16, 
                    d_arr_19__15, d_arr_19__14, d_arr_19__13, d_arr_19__12, 
                    d_arr_19__11, d_arr_19__10, d_arr_19__9, d_arr_19__8, 
                    d_arr_19__7, d_arr_19__6, d_arr_19__5, d_arr_19__4, 
                    d_arr_19__3, d_arr_19__2, d_arr_19__1, d_arr_19__0, 
                    d_arr_20__31, d_arr_20__30, d_arr_20__29, d_arr_20__28, 
                    d_arr_20__27, d_arr_20__26, d_arr_20__25, d_arr_20__24, 
                    d_arr_20__23, d_arr_20__22, d_arr_20__21, d_arr_20__20, 
                    d_arr_20__19, d_arr_20__18, d_arr_20__17, d_arr_20__16, 
                    d_arr_20__15, d_arr_20__14, d_arr_20__13, d_arr_20__12, 
                    d_arr_20__11, d_arr_20__10, d_arr_20__9, d_arr_20__8, 
                    d_arr_20__7, d_arr_20__6, d_arr_20__5, d_arr_20__4, 
                    d_arr_20__3, d_arr_20__2, d_arr_20__1, d_arr_20__0, 
                    d_arr_21__31, d_arr_21__30, d_arr_21__29, d_arr_21__28, 
                    d_arr_21__27, d_arr_21__26, d_arr_21__25, d_arr_21__24, 
                    d_arr_21__23, d_arr_21__22, d_arr_21__21, d_arr_21__20, 
                    d_arr_21__19, d_arr_21__18, d_arr_21__17, d_arr_21__16, 
                    d_arr_21__15, d_arr_21__14, d_arr_21__13, d_arr_21__12, 
                    d_arr_21__11, d_arr_21__10, d_arr_21__9, d_arr_21__8, 
                    d_arr_21__7, d_arr_21__6, d_arr_21__5, d_arr_21__4, 
                    d_arr_21__3, d_arr_21__2, d_arr_21__1, d_arr_21__0, 
                    d_arr_22__31, d_arr_22__30, d_arr_22__29, d_arr_22__28, 
                    d_arr_22__27, d_arr_22__26, d_arr_22__25, d_arr_22__24, 
                    d_arr_22__23, d_arr_22__22, d_arr_22__21, d_arr_22__20, 
                    d_arr_22__19, d_arr_22__18, d_arr_22__17, d_arr_22__16, 
                    d_arr_22__15, d_arr_22__14, d_arr_22__13, d_arr_22__12, 
                    d_arr_22__11, d_arr_22__10, d_arr_22__9, d_arr_22__8, 
                    d_arr_22__7, d_arr_22__6, d_arr_22__5, d_arr_22__4, 
                    d_arr_22__3, d_arr_22__2, d_arr_22__1, d_arr_22__0, 
                    d_arr_23__31, d_arr_23__30, d_arr_23__29, d_arr_23__28, 
                    d_arr_23__27, d_arr_23__26, d_arr_23__25, d_arr_23__24, 
                    d_arr_23__23, d_arr_23__22, d_arr_23__21, d_arr_23__20, 
                    d_arr_23__19, d_arr_23__18, d_arr_23__17, d_arr_23__16, 
                    d_arr_23__15, d_arr_23__14, d_arr_23__13, d_arr_23__12, 
                    d_arr_23__11, d_arr_23__10, d_arr_23__9, d_arr_23__8, 
                    d_arr_23__7, d_arr_23__6, d_arr_23__5, d_arr_23__4, 
                    d_arr_23__3, d_arr_23__2, d_arr_23__1, d_arr_23__0, 
                    d_arr_24__31, d_arr_24__30, d_arr_24__29, d_arr_24__28, 
                    d_arr_24__27, d_arr_24__26, d_arr_24__25, d_arr_24__24, 
                    d_arr_24__23, d_arr_24__22, d_arr_24__21, d_arr_24__20, 
                    d_arr_24__19, d_arr_24__18, d_arr_24__17, d_arr_24__16, 
                    d_arr_24__15, d_arr_24__14, d_arr_24__13, d_arr_24__12, 
                    d_arr_24__11, d_arr_24__10, d_arr_24__9, d_arr_24__8, 
                    d_arr_24__7, d_arr_24__6, d_arr_24__5, d_arr_24__4, 
                    d_arr_24__3, d_arr_24__2, d_arr_24__1, d_arr_24__0, 
                    q_arr_0__31, q_arr_0__30, q_arr_0__29, q_arr_0__28, 
                    q_arr_0__27, q_arr_0__26, q_arr_0__25, q_arr_0__24, 
                    q_arr_0__23, q_arr_0__22, q_arr_0__21, q_arr_0__20, 
                    q_arr_0__19, q_arr_0__18, q_arr_0__17, q_arr_0__16, 
                    q_arr_0__15, q_arr_0__14, q_arr_0__13, q_arr_0__12, 
                    q_arr_0__11, q_arr_0__10, q_arr_0__9, q_arr_0__8, q_arr_0__7, 
                    q_arr_0__6, q_arr_0__5, q_arr_0__4, q_arr_0__3, q_arr_0__2, 
                    q_arr_0__1, q_arr_0__0, q_arr_1__31, q_arr_1__30, 
                    q_arr_1__29, q_arr_1__28, q_arr_1__27, q_arr_1__26, 
                    q_arr_1__25, q_arr_1__24, q_arr_1__23, q_arr_1__22, 
                    q_arr_1__21, q_arr_1__20, q_arr_1__19, q_arr_1__18, 
                    q_arr_1__17, q_arr_1__16, q_arr_1__15, q_arr_1__14, 
                    q_arr_1__13, q_arr_1__12, q_arr_1__11, q_arr_1__10, 
                    q_arr_1__9, q_arr_1__8, q_arr_1__7, q_arr_1__6, q_arr_1__5, 
                    q_arr_1__4, q_arr_1__3, q_arr_1__2, q_arr_1__1, q_arr_1__0, 
                    q_arr_2__31, q_arr_2__30, q_arr_2__29, q_arr_2__28, 
                    q_arr_2__27, q_arr_2__26, q_arr_2__25, q_arr_2__24, 
                    q_arr_2__23, q_arr_2__22, q_arr_2__21, q_arr_2__20, 
                    q_arr_2__19, q_arr_2__18, q_arr_2__17, q_arr_2__16, 
                    q_arr_2__15, q_arr_2__14, q_arr_2__13, q_arr_2__12, 
                    q_arr_2__11, q_arr_2__10, q_arr_2__9, q_arr_2__8, q_arr_2__7, 
                    q_arr_2__6, q_arr_2__5, q_arr_2__4, q_arr_2__3, q_arr_2__2, 
                    q_arr_2__1, q_arr_2__0, q_arr_3__31, q_arr_3__30, 
                    q_arr_3__29, q_arr_3__28, q_arr_3__27, q_arr_3__26, 
                    q_arr_3__25, q_arr_3__24, q_arr_3__23, q_arr_3__22, 
                    q_arr_3__21, q_arr_3__20, q_arr_3__19, q_arr_3__18, 
                    q_arr_3__17, q_arr_3__16, q_arr_3__15, q_arr_3__14, 
                    q_arr_3__13, q_arr_3__12, q_arr_3__11, q_arr_3__10, 
                    q_arr_3__9, q_arr_3__8, q_arr_3__7, q_arr_3__6, q_arr_3__5, 
                    q_arr_3__4, q_arr_3__3, q_arr_3__2, q_arr_3__1, q_arr_3__0, 
                    q_arr_4__31, q_arr_4__30, q_arr_4__29, q_arr_4__28, 
                    q_arr_4__27, q_arr_4__26, q_arr_4__25, q_arr_4__24, 
                    q_arr_4__23, q_arr_4__22, q_arr_4__21, q_arr_4__20, 
                    q_arr_4__19, q_arr_4__18, q_arr_4__17, q_arr_4__16, 
                    q_arr_4__15, q_arr_4__14, q_arr_4__13, q_arr_4__12, 
                    q_arr_4__11, q_arr_4__10, q_arr_4__9, q_arr_4__8, q_arr_4__7, 
                    q_arr_4__6, q_arr_4__5, q_arr_4__4, q_arr_4__3, q_arr_4__2, 
                    q_arr_4__1, q_arr_4__0, q_arr_5__31, q_arr_5__30, 
                    q_arr_5__29, q_arr_5__28, q_arr_5__27, q_arr_5__26, 
                    q_arr_5__25, q_arr_5__24, q_arr_5__23, q_arr_5__22, 
                    q_arr_5__21, q_arr_5__20, q_arr_5__19, q_arr_5__18, 
                    q_arr_5__17, q_arr_5__16, q_arr_5__15, q_arr_5__14, 
                    q_arr_5__13, q_arr_5__12, q_arr_5__11, q_arr_5__10, 
                    q_arr_5__9, q_arr_5__8, q_arr_5__7, q_arr_5__6, q_arr_5__5, 
                    q_arr_5__4, q_arr_5__3, q_arr_5__2, q_arr_5__1, q_arr_5__0, 
                    q_arr_6__31, q_arr_6__30, q_arr_6__29, q_arr_6__28, 
                    q_arr_6__27, q_arr_6__26, q_arr_6__25, q_arr_6__24, 
                    q_arr_6__23, q_arr_6__22, q_arr_6__21, q_arr_6__20, 
                    q_arr_6__19, q_arr_6__18, q_arr_6__17, q_arr_6__16, 
                    q_arr_6__15, q_arr_6__14, q_arr_6__13, q_arr_6__12, 
                    q_arr_6__11, q_arr_6__10, q_arr_6__9, q_arr_6__8, q_arr_6__7, 
                    q_arr_6__6, q_arr_6__5, q_arr_6__4, q_arr_6__3, q_arr_6__2, 
                    q_arr_6__1, q_arr_6__0, q_arr_7__31, q_arr_7__30, 
                    q_arr_7__29, q_arr_7__28, q_arr_7__27, q_arr_7__26, 
                    q_arr_7__25, q_arr_7__24, q_arr_7__23, q_arr_7__22, 
                    q_arr_7__21, q_arr_7__20, q_arr_7__19, q_arr_7__18, 
                    q_arr_7__17, q_arr_7__16, q_arr_7__15, q_arr_7__14, 
                    q_arr_7__13, q_arr_7__12, q_arr_7__11, q_arr_7__10, 
                    q_arr_7__9, q_arr_7__8, q_arr_7__7, q_arr_7__6, q_arr_7__5, 
                    q_arr_7__4, q_arr_7__3, q_arr_7__2, q_arr_7__1, q_arr_7__0, 
                    q_arr_8__31, q_arr_8__30, q_arr_8__29, q_arr_8__28, 
                    q_arr_8__27, q_arr_8__26, q_arr_8__25, q_arr_8__24, 
                    q_arr_8__23, q_arr_8__22, q_arr_8__21, q_arr_8__20, 
                    q_arr_8__19, q_arr_8__18, q_arr_8__17, q_arr_8__16, 
                    q_arr_8__15, q_arr_8__14, q_arr_8__13, q_arr_8__12, 
                    q_arr_8__11, q_arr_8__10, q_arr_8__9, q_arr_8__8, q_arr_8__7, 
                    q_arr_8__6, q_arr_8__5, q_arr_8__4, q_arr_8__3, q_arr_8__2, 
                    q_arr_8__1, q_arr_8__0, q_arr_9__31, q_arr_9__30, 
                    q_arr_9__29, q_arr_9__28, q_arr_9__27, q_arr_9__26, 
                    q_arr_9__25, q_arr_9__24, q_arr_9__23, q_arr_9__22, 
                    q_arr_9__21, q_arr_9__20, q_arr_9__19, q_arr_9__18, 
                    q_arr_9__17, q_arr_9__16, q_arr_9__15, q_arr_9__14, 
                    q_arr_9__13, q_arr_9__12, q_arr_9__11, q_arr_9__10, 
                    q_arr_9__9, q_arr_9__8, q_arr_9__7, q_arr_9__6, q_arr_9__5, 
                    q_arr_9__4, q_arr_9__3, q_arr_9__2, q_arr_9__1, q_arr_9__0, 
                    q_arr_10__31, q_arr_10__30, q_arr_10__29, q_arr_10__28, 
                    q_arr_10__27, q_arr_10__26, q_arr_10__25, q_arr_10__24, 
                    q_arr_10__23, q_arr_10__22, q_arr_10__21, q_arr_10__20, 
                    q_arr_10__19, q_arr_10__18, q_arr_10__17, q_arr_10__16, 
                    q_arr_10__15, q_arr_10__14, q_arr_10__13, q_arr_10__12, 
                    q_arr_10__11, q_arr_10__10, q_arr_10__9, q_arr_10__8, 
                    q_arr_10__7, q_arr_10__6, q_arr_10__5, q_arr_10__4, 
                    q_arr_10__3, q_arr_10__2, q_arr_10__1, q_arr_10__0, 
                    q_arr_11__31, q_arr_11__30, q_arr_11__29, q_arr_11__28, 
                    q_arr_11__27, q_arr_11__26, q_arr_11__25, q_arr_11__24, 
                    q_arr_11__23, q_arr_11__22, q_arr_11__21, q_arr_11__20, 
                    q_arr_11__19, q_arr_11__18, q_arr_11__17, q_arr_11__16, 
                    q_arr_11__15, q_arr_11__14, q_arr_11__13, q_arr_11__12, 
                    q_arr_11__11, q_arr_11__10, q_arr_11__9, q_arr_11__8, 
                    q_arr_11__7, q_arr_11__6, q_arr_11__5, q_arr_11__4, 
                    q_arr_11__3, q_arr_11__2, q_arr_11__1, q_arr_11__0, 
                    q_arr_12__31, q_arr_12__30, q_arr_12__29, q_arr_12__28, 
                    q_arr_12__27, q_arr_12__26, q_arr_12__25, q_arr_12__24, 
                    q_arr_12__23, q_arr_12__22, q_arr_12__21, q_arr_12__20, 
                    q_arr_12__19, q_arr_12__18, q_arr_12__17, q_arr_12__16, 
                    q_arr_12__15, q_arr_12__14, q_arr_12__13, q_arr_12__12, 
                    q_arr_12__11, q_arr_12__10, q_arr_12__9, q_arr_12__8, 
                    q_arr_12__7, q_arr_12__6, q_arr_12__5, q_arr_12__4, 
                    q_arr_12__3, q_arr_12__2, q_arr_12__1, q_arr_12__0, 
                    q_arr_13__31, q_arr_13__30, q_arr_13__29, q_arr_13__28, 
                    q_arr_13__27, q_arr_13__26, q_arr_13__25, q_arr_13__24, 
                    q_arr_13__23, q_arr_13__22, q_arr_13__21, q_arr_13__20, 
                    q_arr_13__19, q_arr_13__18, q_arr_13__17, q_arr_13__16, 
                    q_arr_13__15, q_arr_13__14, q_arr_13__13, q_arr_13__12, 
                    q_arr_13__11, q_arr_13__10, q_arr_13__9, q_arr_13__8, 
                    q_arr_13__7, q_arr_13__6, q_arr_13__5, q_arr_13__4, 
                    q_arr_13__3, q_arr_13__2, q_arr_13__1, q_arr_13__0, 
                    q_arr_14__31, q_arr_14__30, q_arr_14__29, q_arr_14__28, 
                    q_arr_14__27, q_arr_14__26, q_arr_14__25, q_arr_14__24, 
                    q_arr_14__23, q_arr_14__22, q_arr_14__21, q_arr_14__20, 
                    q_arr_14__19, q_arr_14__18, q_arr_14__17, q_arr_14__16, 
                    q_arr_14__15, q_arr_14__14, q_arr_14__13, q_arr_14__12, 
                    q_arr_14__11, q_arr_14__10, q_arr_14__9, q_arr_14__8, 
                    q_arr_14__7, q_arr_14__6, q_arr_14__5, q_arr_14__4, 
                    q_arr_14__3, q_arr_14__2, q_arr_14__1, q_arr_14__0, 
                    q_arr_15__31, q_arr_15__30, q_arr_15__29, q_arr_15__28, 
                    q_arr_15__27, q_arr_15__26, q_arr_15__25, q_arr_15__24, 
                    q_arr_15__23, q_arr_15__22, q_arr_15__21, q_arr_15__20, 
                    q_arr_15__19, q_arr_15__18, q_arr_15__17, q_arr_15__16, 
                    q_arr_15__15, q_arr_15__14, q_arr_15__13, q_arr_15__12, 
                    q_arr_15__11, q_arr_15__10, q_arr_15__9, q_arr_15__8, 
                    q_arr_15__7, q_arr_15__6, q_arr_15__5, q_arr_15__4, 
                    q_arr_15__3, q_arr_15__2, q_arr_15__1, q_arr_15__0, 
                    q_arr_16__31, q_arr_16__30, q_arr_16__29, q_arr_16__28, 
                    q_arr_16__27, q_arr_16__26, q_arr_16__25, q_arr_16__24, 
                    q_arr_16__23, q_arr_16__22, q_arr_16__21, q_arr_16__20, 
                    q_arr_16__19, q_arr_16__18, q_arr_16__17, q_arr_16__16, 
                    q_arr_16__15, q_arr_16__14, q_arr_16__13, q_arr_16__12, 
                    q_arr_16__11, q_arr_16__10, q_arr_16__9, q_arr_16__8, 
                    q_arr_16__7, q_arr_16__6, q_arr_16__5, q_arr_16__4, 
                    q_arr_16__3, q_arr_16__2, q_arr_16__1, q_arr_16__0, 
                    q_arr_17__31, q_arr_17__30, q_arr_17__29, q_arr_17__28, 
                    q_arr_17__27, q_arr_17__26, q_arr_17__25, q_arr_17__24, 
                    q_arr_17__23, q_arr_17__22, q_arr_17__21, q_arr_17__20, 
                    q_arr_17__19, q_arr_17__18, q_arr_17__17, q_arr_17__16, 
                    q_arr_17__15, q_arr_17__14, q_arr_17__13, q_arr_17__12, 
                    q_arr_17__11, q_arr_17__10, q_arr_17__9, q_arr_17__8, 
                    q_arr_17__7, q_arr_17__6, q_arr_17__5, q_arr_17__4, 
                    q_arr_17__3, q_arr_17__2, q_arr_17__1, q_arr_17__0, 
                    q_arr_18__31, q_arr_18__30, q_arr_18__29, q_arr_18__28, 
                    q_arr_18__27, q_arr_18__26, q_arr_18__25, q_arr_18__24, 
                    q_arr_18__23, q_arr_18__22, q_arr_18__21, q_arr_18__20, 
                    q_arr_18__19, q_arr_18__18, q_arr_18__17, q_arr_18__16, 
                    q_arr_18__15, q_arr_18__14, q_arr_18__13, q_arr_18__12, 
                    q_arr_18__11, q_arr_18__10, q_arr_18__9, q_arr_18__8, 
                    q_arr_18__7, q_arr_18__6, q_arr_18__5, q_arr_18__4, 
                    q_arr_18__3, q_arr_18__2, q_arr_18__1, q_arr_18__0, 
                    q_arr_19__31, q_arr_19__30, q_arr_19__29, q_arr_19__28, 
                    q_arr_19__27, q_arr_19__26, q_arr_19__25, q_arr_19__24, 
                    q_arr_19__23, q_arr_19__22, q_arr_19__21, q_arr_19__20, 
                    q_arr_19__19, q_arr_19__18, q_arr_19__17, q_arr_19__16, 
                    q_arr_19__15, q_arr_19__14, q_arr_19__13, q_arr_19__12, 
                    q_arr_19__11, q_arr_19__10, q_arr_19__9, q_arr_19__8, 
                    q_arr_19__7, q_arr_19__6, q_arr_19__5, q_arr_19__4, 
                    q_arr_19__3, q_arr_19__2, q_arr_19__1, q_arr_19__0, 
                    q_arr_20__31, q_arr_20__30, q_arr_20__29, q_arr_20__28, 
                    q_arr_20__27, q_arr_20__26, q_arr_20__25, q_arr_20__24, 
                    q_arr_20__23, q_arr_20__22, q_arr_20__21, q_arr_20__20, 
                    q_arr_20__19, q_arr_20__18, q_arr_20__17, q_arr_20__16, 
                    q_arr_20__15, q_arr_20__14, q_arr_20__13, q_arr_20__12, 
                    q_arr_20__11, q_arr_20__10, q_arr_20__9, q_arr_20__8, 
                    q_arr_20__7, q_arr_20__6, q_arr_20__5, q_arr_20__4, 
                    q_arr_20__3, q_arr_20__2, q_arr_20__1, q_arr_20__0, 
                    q_arr_21__31, q_arr_21__30, q_arr_21__29, q_arr_21__28, 
                    q_arr_21__27, q_arr_21__26, q_arr_21__25, q_arr_21__24, 
                    q_arr_21__23, q_arr_21__22, q_arr_21__21, q_arr_21__20, 
                    q_arr_21__19, q_arr_21__18, q_arr_21__17, q_arr_21__16, 
                    q_arr_21__15, q_arr_21__14, q_arr_21__13, q_arr_21__12, 
                    q_arr_21__11, q_arr_21__10, q_arr_21__9, q_arr_21__8, 
                    q_arr_21__7, q_arr_21__6, q_arr_21__5, q_arr_21__4, 
                    q_arr_21__3, q_arr_21__2, q_arr_21__1, q_arr_21__0, 
                    q_arr_22__31, q_arr_22__30, q_arr_22__29, q_arr_22__28, 
                    q_arr_22__27, q_arr_22__26, q_arr_22__25, q_arr_22__24, 
                    q_arr_22__23, q_arr_22__22, q_arr_22__21, q_arr_22__20, 
                    q_arr_22__19, q_arr_22__18, q_arr_22__17, q_arr_22__16, 
                    q_arr_22__15, q_arr_22__14, q_arr_22__13, q_arr_22__12, 
                    q_arr_22__11, q_arr_22__10, q_arr_22__9, q_arr_22__8, 
                    q_arr_22__7, q_arr_22__6, q_arr_22__5, q_arr_22__4, 
                    q_arr_22__3, q_arr_22__2, q_arr_22__1, q_arr_22__0, 
                    q_arr_23__31, q_arr_23__30, q_arr_23__29, q_arr_23__28, 
                    q_arr_23__27, q_arr_23__26, q_arr_23__25, q_arr_23__24, 
                    q_arr_23__23, q_arr_23__22, q_arr_23__21, q_arr_23__20, 
                    q_arr_23__19, q_arr_23__18, q_arr_23__17, q_arr_23__16, 
                    q_arr_23__15, q_arr_23__14, q_arr_23__13, q_arr_23__12, 
                    q_arr_23__11, q_arr_23__10, q_arr_23__9, q_arr_23__8, 
                    q_arr_23__7, q_arr_23__6, q_arr_23__5, q_arr_23__4, 
                    q_arr_23__3, q_arr_23__2, q_arr_23__1, q_arr_23__0, 
                    q_arr_24__31, q_arr_24__30, q_arr_24__29, q_arr_24__28, 
                    q_arr_24__27, q_arr_24__26, q_arr_24__25, q_arr_24__24, 
                    q_arr_24__23, q_arr_24__22, q_arr_24__21, q_arr_24__20, 
                    q_arr_24__19, q_arr_24__18, q_arr_24__17, q_arr_24__16, 
                    q_arr_24__15, q_arr_24__14, q_arr_24__13, q_arr_24__12, 
                    q_arr_24__11, q_arr_24__10, q_arr_24__9, q_arr_24__8, 
                    q_arr_24__7, q_arr_24__6, q_arr_24__5, q_arr_24__4, 
                    q_arr_24__3, q_arr_24__2, q_arr_24__1, q_arr_24__0, 
                    operation, filter_size ) ;

    output d_arr_0__31 ;
    output d_arr_0__30 ;
    output d_arr_0__29 ;
    output d_arr_0__28 ;
    output d_arr_0__27 ;
    output d_arr_0__26 ;
    output d_arr_0__25 ;
    output d_arr_0__24 ;
    output d_arr_0__23 ;
    output d_arr_0__22 ;
    output d_arr_0__21 ;
    output d_arr_0__20 ;
    output d_arr_0__19 ;
    output d_arr_0__18 ;
    output d_arr_0__17 ;
    output d_arr_0__16 ;
    output d_arr_0__15 ;
    output d_arr_0__14 ;
    output d_arr_0__13 ;
    output d_arr_0__12 ;
    output d_arr_0__11 ;
    output d_arr_0__10 ;
    output d_arr_0__9 ;
    output d_arr_0__8 ;
    output d_arr_0__7 ;
    output d_arr_0__6 ;
    output d_arr_0__5 ;
    output d_arr_0__4 ;
    output d_arr_0__3 ;
    output d_arr_0__2 ;
    output d_arr_0__1 ;
    output d_arr_0__0 ;
    output d_arr_1__31 ;
    output d_arr_1__30 ;
    output d_arr_1__29 ;
    output d_arr_1__28 ;
    output d_arr_1__27 ;
    output d_arr_1__26 ;
    output d_arr_1__25 ;
    output d_arr_1__24 ;
    output d_arr_1__23 ;
    output d_arr_1__22 ;
    output d_arr_1__21 ;
    output d_arr_1__20 ;
    output d_arr_1__19 ;
    output d_arr_1__18 ;
    output d_arr_1__17 ;
    output d_arr_1__16 ;
    output d_arr_1__15 ;
    output d_arr_1__14 ;
    output d_arr_1__13 ;
    output d_arr_1__12 ;
    output d_arr_1__11 ;
    output d_arr_1__10 ;
    output d_arr_1__9 ;
    output d_arr_1__8 ;
    output d_arr_1__7 ;
    output d_arr_1__6 ;
    output d_arr_1__5 ;
    output d_arr_1__4 ;
    output d_arr_1__3 ;
    output d_arr_1__2 ;
    output d_arr_1__1 ;
    output d_arr_1__0 ;
    output d_arr_2__31 ;
    output d_arr_2__30 ;
    output d_arr_2__29 ;
    output d_arr_2__28 ;
    output d_arr_2__27 ;
    output d_arr_2__26 ;
    output d_arr_2__25 ;
    output d_arr_2__24 ;
    output d_arr_2__23 ;
    output d_arr_2__22 ;
    output d_arr_2__21 ;
    output d_arr_2__20 ;
    output d_arr_2__19 ;
    output d_arr_2__18 ;
    output d_arr_2__17 ;
    output d_arr_2__16 ;
    output d_arr_2__15 ;
    output d_arr_2__14 ;
    output d_arr_2__13 ;
    output d_arr_2__12 ;
    output d_arr_2__11 ;
    output d_arr_2__10 ;
    output d_arr_2__9 ;
    output d_arr_2__8 ;
    output d_arr_2__7 ;
    output d_arr_2__6 ;
    output d_arr_2__5 ;
    output d_arr_2__4 ;
    output d_arr_2__3 ;
    output d_arr_2__2 ;
    output d_arr_2__1 ;
    output d_arr_2__0 ;
    output d_arr_3__31 ;
    output d_arr_3__30 ;
    output d_arr_3__29 ;
    output d_arr_3__28 ;
    output d_arr_3__27 ;
    output d_arr_3__26 ;
    output d_arr_3__25 ;
    output d_arr_3__24 ;
    output d_arr_3__23 ;
    output d_arr_3__22 ;
    output d_arr_3__21 ;
    output d_arr_3__20 ;
    output d_arr_3__19 ;
    output d_arr_3__18 ;
    output d_arr_3__17 ;
    output d_arr_3__16 ;
    output d_arr_3__15 ;
    output d_arr_3__14 ;
    output d_arr_3__13 ;
    output d_arr_3__12 ;
    output d_arr_3__11 ;
    output d_arr_3__10 ;
    output d_arr_3__9 ;
    output d_arr_3__8 ;
    output d_arr_3__7 ;
    output d_arr_3__6 ;
    output d_arr_3__5 ;
    output d_arr_3__4 ;
    output d_arr_3__3 ;
    output d_arr_3__2 ;
    output d_arr_3__1 ;
    output d_arr_3__0 ;
    output d_arr_4__31 ;
    output d_arr_4__30 ;
    output d_arr_4__29 ;
    output d_arr_4__28 ;
    output d_arr_4__27 ;
    output d_arr_4__26 ;
    output d_arr_4__25 ;
    output d_arr_4__24 ;
    output d_arr_4__23 ;
    output d_arr_4__22 ;
    output d_arr_4__21 ;
    output d_arr_4__20 ;
    output d_arr_4__19 ;
    output d_arr_4__18 ;
    output d_arr_4__17 ;
    output d_arr_4__16 ;
    output d_arr_4__15 ;
    output d_arr_4__14 ;
    output d_arr_4__13 ;
    output d_arr_4__12 ;
    output d_arr_4__11 ;
    output d_arr_4__10 ;
    output d_arr_4__9 ;
    output d_arr_4__8 ;
    output d_arr_4__7 ;
    output d_arr_4__6 ;
    output d_arr_4__5 ;
    output d_arr_4__4 ;
    output d_arr_4__3 ;
    output d_arr_4__2 ;
    output d_arr_4__1 ;
    output d_arr_4__0 ;
    output d_arr_5__31 ;
    output d_arr_5__30 ;
    output d_arr_5__29 ;
    output d_arr_5__28 ;
    output d_arr_5__27 ;
    output d_arr_5__26 ;
    output d_arr_5__25 ;
    output d_arr_5__24 ;
    output d_arr_5__23 ;
    output d_arr_5__22 ;
    output d_arr_5__21 ;
    output d_arr_5__20 ;
    output d_arr_5__19 ;
    output d_arr_5__18 ;
    output d_arr_5__17 ;
    output d_arr_5__16 ;
    output d_arr_5__15 ;
    output d_arr_5__14 ;
    output d_arr_5__13 ;
    output d_arr_5__12 ;
    output d_arr_5__11 ;
    output d_arr_5__10 ;
    output d_arr_5__9 ;
    output d_arr_5__8 ;
    output d_arr_5__7 ;
    output d_arr_5__6 ;
    output d_arr_5__5 ;
    output d_arr_5__4 ;
    output d_arr_5__3 ;
    output d_arr_5__2 ;
    output d_arr_5__1 ;
    output d_arr_5__0 ;
    output d_arr_6__31 ;
    output d_arr_6__30 ;
    output d_arr_6__29 ;
    output d_arr_6__28 ;
    output d_arr_6__27 ;
    output d_arr_6__26 ;
    output d_arr_6__25 ;
    output d_arr_6__24 ;
    output d_arr_6__23 ;
    output d_arr_6__22 ;
    output d_arr_6__21 ;
    output d_arr_6__20 ;
    output d_arr_6__19 ;
    output d_arr_6__18 ;
    output d_arr_6__17 ;
    output d_arr_6__16 ;
    output d_arr_6__15 ;
    output d_arr_6__14 ;
    output d_arr_6__13 ;
    output d_arr_6__12 ;
    output d_arr_6__11 ;
    output d_arr_6__10 ;
    output d_arr_6__9 ;
    output d_arr_6__8 ;
    output d_arr_6__7 ;
    output d_arr_6__6 ;
    output d_arr_6__5 ;
    output d_arr_6__4 ;
    output d_arr_6__3 ;
    output d_arr_6__2 ;
    output d_arr_6__1 ;
    output d_arr_6__0 ;
    output d_arr_7__31 ;
    output d_arr_7__30 ;
    output d_arr_7__29 ;
    output d_arr_7__28 ;
    output d_arr_7__27 ;
    output d_arr_7__26 ;
    output d_arr_7__25 ;
    output d_arr_7__24 ;
    output d_arr_7__23 ;
    output d_arr_7__22 ;
    output d_arr_7__21 ;
    output d_arr_7__20 ;
    output d_arr_7__19 ;
    output d_arr_7__18 ;
    output d_arr_7__17 ;
    output d_arr_7__16 ;
    output d_arr_7__15 ;
    output d_arr_7__14 ;
    output d_arr_7__13 ;
    output d_arr_7__12 ;
    output d_arr_7__11 ;
    output d_arr_7__10 ;
    output d_arr_7__9 ;
    output d_arr_7__8 ;
    output d_arr_7__7 ;
    output d_arr_7__6 ;
    output d_arr_7__5 ;
    output d_arr_7__4 ;
    output d_arr_7__3 ;
    output d_arr_7__2 ;
    output d_arr_7__1 ;
    output d_arr_7__0 ;
    output d_arr_8__31 ;
    output d_arr_8__30 ;
    output d_arr_8__29 ;
    output d_arr_8__28 ;
    output d_arr_8__27 ;
    output d_arr_8__26 ;
    output d_arr_8__25 ;
    output d_arr_8__24 ;
    output d_arr_8__23 ;
    output d_arr_8__22 ;
    output d_arr_8__21 ;
    output d_arr_8__20 ;
    output d_arr_8__19 ;
    output d_arr_8__18 ;
    output d_arr_8__17 ;
    output d_arr_8__16 ;
    output d_arr_8__15 ;
    output d_arr_8__14 ;
    output d_arr_8__13 ;
    output d_arr_8__12 ;
    output d_arr_8__11 ;
    output d_arr_8__10 ;
    output d_arr_8__9 ;
    output d_arr_8__8 ;
    output d_arr_8__7 ;
    output d_arr_8__6 ;
    output d_arr_8__5 ;
    output d_arr_8__4 ;
    output d_arr_8__3 ;
    output d_arr_8__2 ;
    output d_arr_8__1 ;
    output d_arr_8__0 ;
    output d_arr_9__31 ;
    output d_arr_9__30 ;
    output d_arr_9__29 ;
    output d_arr_9__28 ;
    output d_arr_9__27 ;
    output d_arr_9__26 ;
    output d_arr_9__25 ;
    output d_arr_9__24 ;
    output d_arr_9__23 ;
    output d_arr_9__22 ;
    output d_arr_9__21 ;
    output d_arr_9__20 ;
    output d_arr_9__19 ;
    output d_arr_9__18 ;
    output d_arr_9__17 ;
    output d_arr_9__16 ;
    output d_arr_9__15 ;
    output d_arr_9__14 ;
    output d_arr_9__13 ;
    output d_arr_9__12 ;
    output d_arr_9__11 ;
    output d_arr_9__10 ;
    output d_arr_9__9 ;
    output d_arr_9__8 ;
    output d_arr_9__7 ;
    output d_arr_9__6 ;
    output d_arr_9__5 ;
    output d_arr_9__4 ;
    output d_arr_9__3 ;
    output d_arr_9__2 ;
    output d_arr_9__1 ;
    output d_arr_9__0 ;
    output d_arr_10__31 ;
    output d_arr_10__30 ;
    output d_arr_10__29 ;
    output d_arr_10__28 ;
    output d_arr_10__27 ;
    output d_arr_10__26 ;
    output d_arr_10__25 ;
    output d_arr_10__24 ;
    output d_arr_10__23 ;
    output d_arr_10__22 ;
    output d_arr_10__21 ;
    output d_arr_10__20 ;
    output d_arr_10__19 ;
    output d_arr_10__18 ;
    output d_arr_10__17 ;
    output d_arr_10__16 ;
    output d_arr_10__15 ;
    output d_arr_10__14 ;
    output d_arr_10__13 ;
    output d_arr_10__12 ;
    output d_arr_10__11 ;
    output d_arr_10__10 ;
    output d_arr_10__9 ;
    output d_arr_10__8 ;
    output d_arr_10__7 ;
    output d_arr_10__6 ;
    output d_arr_10__5 ;
    output d_arr_10__4 ;
    output d_arr_10__3 ;
    output d_arr_10__2 ;
    output d_arr_10__1 ;
    output d_arr_10__0 ;
    output d_arr_11__31 ;
    output d_arr_11__30 ;
    output d_arr_11__29 ;
    output d_arr_11__28 ;
    output d_arr_11__27 ;
    output d_arr_11__26 ;
    output d_arr_11__25 ;
    output d_arr_11__24 ;
    output d_arr_11__23 ;
    output d_arr_11__22 ;
    output d_arr_11__21 ;
    output d_arr_11__20 ;
    output d_arr_11__19 ;
    output d_arr_11__18 ;
    output d_arr_11__17 ;
    output d_arr_11__16 ;
    output d_arr_11__15 ;
    output d_arr_11__14 ;
    output d_arr_11__13 ;
    output d_arr_11__12 ;
    output d_arr_11__11 ;
    output d_arr_11__10 ;
    output d_arr_11__9 ;
    output d_arr_11__8 ;
    output d_arr_11__7 ;
    output d_arr_11__6 ;
    output d_arr_11__5 ;
    output d_arr_11__4 ;
    output d_arr_11__3 ;
    output d_arr_11__2 ;
    output d_arr_11__1 ;
    output d_arr_11__0 ;
    output d_arr_12__31 ;
    output d_arr_12__30 ;
    output d_arr_12__29 ;
    output d_arr_12__28 ;
    output d_arr_12__27 ;
    output d_arr_12__26 ;
    output d_arr_12__25 ;
    output d_arr_12__24 ;
    output d_arr_12__23 ;
    output d_arr_12__22 ;
    output d_arr_12__21 ;
    output d_arr_12__20 ;
    output d_arr_12__19 ;
    output d_arr_12__18 ;
    output d_arr_12__17 ;
    output d_arr_12__16 ;
    output d_arr_12__15 ;
    output d_arr_12__14 ;
    output d_arr_12__13 ;
    output d_arr_12__12 ;
    output d_arr_12__11 ;
    output d_arr_12__10 ;
    output d_arr_12__9 ;
    output d_arr_12__8 ;
    output d_arr_12__7 ;
    output d_arr_12__6 ;
    output d_arr_12__5 ;
    output d_arr_12__4 ;
    output d_arr_12__3 ;
    output d_arr_12__2 ;
    output d_arr_12__1 ;
    output d_arr_12__0 ;
    output d_arr_13__31 ;
    output d_arr_13__30 ;
    output d_arr_13__29 ;
    output d_arr_13__28 ;
    output d_arr_13__27 ;
    output d_arr_13__26 ;
    output d_arr_13__25 ;
    output d_arr_13__24 ;
    output d_arr_13__23 ;
    output d_arr_13__22 ;
    output d_arr_13__21 ;
    output d_arr_13__20 ;
    output d_arr_13__19 ;
    output d_arr_13__18 ;
    output d_arr_13__17 ;
    output d_arr_13__16 ;
    output d_arr_13__15 ;
    output d_arr_13__14 ;
    output d_arr_13__13 ;
    output d_arr_13__12 ;
    output d_arr_13__11 ;
    output d_arr_13__10 ;
    output d_arr_13__9 ;
    output d_arr_13__8 ;
    output d_arr_13__7 ;
    output d_arr_13__6 ;
    output d_arr_13__5 ;
    output d_arr_13__4 ;
    output d_arr_13__3 ;
    output d_arr_13__2 ;
    output d_arr_13__1 ;
    output d_arr_13__0 ;
    output d_arr_14__31 ;
    output d_arr_14__30 ;
    output d_arr_14__29 ;
    output d_arr_14__28 ;
    output d_arr_14__27 ;
    output d_arr_14__26 ;
    output d_arr_14__25 ;
    output d_arr_14__24 ;
    output d_arr_14__23 ;
    output d_arr_14__22 ;
    output d_arr_14__21 ;
    output d_arr_14__20 ;
    output d_arr_14__19 ;
    output d_arr_14__18 ;
    output d_arr_14__17 ;
    output d_arr_14__16 ;
    output d_arr_14__15 ;
    output d_arr_14__14 ;
    output d_arr_14__13 ;
    output d_arr_14__12 ;
    output d_arr_14__11 ;
    output d_arr_14__10 ;
    output d_arr_14__9 ;
    output d_arr_14__8 ;
    output d_arr_14__7 ;
    output d_arr_14__6 ;
    output d_arr_14__5 ;
    output d_arr_14__4 ;
    output d_arr_14__3 ;
    output d_arr_14__2 ;
    output d_arr_14__1 ;
    output d_arr_14__0 ;
    output d_arr_15__31 ;
    output d_arr_15__30 ;
    output d_arr_15__29 ;
    output d_arr_15__28 ;
    output d_arr_15__27 ;
    output d_arr_15__26 ;
    output d_arr_15__25 ;
    output d_arr_15__24 ;
    output d_arr_15__23 ;
    output d_arr_15__22 ;
    output d_arr_15__21 ;
    output d_arr_15__20 ;
    output d_arr_15__19 ;
    output d_arr_15__18 ;
    output d_arr_15__17 ;
    output d_arr_15__16 ;
    output d_arr_15__15 ;
    output d_arr_15__14 ;
    output d_arr_15__13 ;
    output d_arr_15__12 ;
    output d_arr_15__11 ;
    output d_arr_15__10 ;
    output d_arr_15__9 ;
    output d_arr_15__8 ;
    output d_arr_15__7 ;
    output d_arr_15__6 ;
    output d_arr_15__5 ;
    output d_arr_15__4 ;
    output d_arr_15__3 ;
    output d_arr_15__2 ;
    output d_arr_15__1 ;
    output d_arr_15__0 ;
    output d_arr_16__31 ;
    output d_arr_16__30 ;
    output d_arr_16__29 ;
    output d_arr_16__28 ;
    output d_arr_16__27 ;
    output d_arr_16__26 ;
    output d_arr_16__25 ;
    output d_arr_16__24 ;
    output d_arr_16__23 ;
    output d_arr_16__22 ;
    output d_arr_16__21 ;
    output d_arr_16__20 ;
    output d_arr_16__19 ;
    output d_arr_16__18 ;
    output d_arr_16__17 ;
    output d_arr_16__16 ;
    output d_arr_16__15 ;
    output d_arr_16__14 ;
    output d_arr_16__13 ;
    output d_arr_16__12 ;
    output d_arr_16__11 ;
    output d_arr_16__10 ;
    output d_arr_16__9 ;
    output d_arr_16__8 ;
    output d_arr_16__7 ;
    output d_arr_16__6 ;
    output d_arr_16__5 ;
    output d_arr_16__4 ;
    output d_arr_16__3 ;
    output d_arr_16__2 ;
    output d_arr_16__1 ;
    output d_arr_16__0 ;
    output d_arr_17__31 ;
    output d_arr_17__30 ;
    output d_arr_17__29 ;
    output d_arr_17__28 ;
    output d_arr_17__27 ;
    output d_arr_17__26 ;
    output d_arr_17__25 ;
    output d_arr_17__24 ;
    output d_arr_17__23 ;
    output d_arr_17__22 ;
    output d_arr_17__21 ;
    output d_arr_17__20 ;
    output d_arr_17__19 ;
    output d_arr_17__18 ;
    output d_arr_17__17 ;
    output d_arr_17__16 ;
    output d_arr_17__15 ;
    output d_arr_17__14 ;
    output d_arr_17__13 ;
    output d_arr_17__12 ;
    output d_arr_17__11 ;
    output d_arr_17__10 ;
    output d_arr_17__9 ;
    output d_arr_17__8 ;
    output d_arr_17__7 ;
    output d_arr_17__6 ;
    output d_arr_17__5 ;
    output d_arr_17__4 ;
    output d_arr_17__3 ;
    output d_arr_17__2 ;
    output d_arr_17__1 ;
    output d_arr_17__0 ;
    output d_arr_18__31 ;
    output d_arr_18__30 ;
    output d_arr_18__29 ;
    output d_arr_18__28 ;
    output d_arr_18__27 ;
    output d_arr_18__26 ;
    output d_arr_18__25 ;
    output d_arr_18__24 ;
    output d_arr_18__23 ;
    output d_arr_18__22 ;
    output d_arr_18__21 ;
    output d_arr_18__20 ;
    output d_arr_18__19 ;
    output d_arr_18__18 ;
    output d_arr_18__17 ;
    output d_arr_18__16 ;
    output d_arr_18__15 ;
    output d_arr_18__14 ;
    output d_arr_18__13 ;
    output d_arr_18__12 ;
    output d_arr_18__11 ;
    output d_arr_18__10 ;
    output d_arr_18__9 ;
    output d_arr_18__8 ;
    output d_arr_18__7 ;
    output d_arr_18__6 ;
    output d_arr_18__5 ;
    output d_arr_18__4 ;
    output d_arr_18__3 ;
    output d_arr_18__2 ;
    output d_arr_18__1 ;
    output d_arr_18__0 ;
    output d_arr_19__31 ;
    output d_arr_19__30 ;
    output d_arr_19__29 ;
    output d_arr_19__28 ;
    output d_arr_19__27 ;
    output d_arr_19__26 ;
    output d_arr_19__25 ;
    output d_arr_19__24 ;
    output d_arr_19__23 ;
    output d_arr_19__22 ;
    output d_arr_19__21 ;
    output d_arr_19__20 ;
    output d_arr_19__19 ;
    output d_arr_19__18 ;
    output d_arr_19__17 ;
    output d_arr_19__16 ;
    output d_arr_19__15 ;
    output d_arr_19__14 ;
    output d_arr_19__13 ;
    output d_arr_19__12 ;
    output d_arr_19__11 ;
    output d_arr_19__10 ;
    output d_arr_19__9 ;
    output d_arr_19__8 ;
    output d_arr_19__7 ;
    output d_arr_19__6 ;
    output d_arr_19__5 ;
    output d_arr_19__4 ;
    output d_arr_19__3 ;
    output d_arr_19__2 ;
    output d_arr_19__1 ;
    output d_arr_19__0 ;
    output d_arr_20__31 ;
    output d_arr_20__30 ;
    output d_arr_20__29 ;
    output d_arr_20__28 ;
    output d_arr_20__27 ;
    output d_arr_20__26 ;
    output d_arr_20__25 ;
    output d_arr_20__24 ;
    output d_arr_20__23 ;
    output d_arr_20__22 ;
    output d_arr_20__21 ;
    output d_arr_20__20 ;
    output d_arr_20__19 ;
    output d_arr_20__18 ;
    output d_arr_20__17 ;
    output d_arr_20__16 ;
    output d_arr_20__15 ;
    output d_arr_20__14 ;
    output d_arr_20__13 ;
    output d_arr_20__12 ;
    output d_arr_20__11 ;
    output d_arr_20__10 ;
    output d_arr_20__9 ;
    output d_arr_20__8 ;
    output d_arr_20__7 ;
    output d_arr_20__6 ;
    output d_arr_20__5 ;
    output d_arr_20__4 ;
    output d_arr_20__3 ;
    output d_arr_20__2 ;
    output d_arr_20__1 ;
    output d_arr_20__0 ;
    output d_arr_21__31 ;
    output d_arr_21__30 ;
    output d_arr_21__29 ;
    output d_arr_21__28 ;
    output d_arr_21__27 ;
    output d_arr_21__26 ;
    output d_arr_21__25 ;
    output d_arr_21__24 ;
    output d_arr_21__23 ;
    output d_arr_21__22 ;
    output d_arr_21__21 ;
    output d_arr_21__20 ;
    output d_arr_21__19 ;
    output d_arr_21__18 ;
    output d_arr_21__17 ;
    output d_arr_21__16 ;
    output d_arr_21__15 ;
    output d_arr_21__14 ;
    output d_arr_21__13 ;
    output d_arr_21__12 ;
    output d_arr_21__11 ;
    output d_arr_21__10 ;
    output d_arr_21__9 ;
    output d_arr_21__8 ;
    output d_arr_21__7 ;
    output d_arr_21__6 ;
    output d_arr_21__5 ;
    output d_arr_21__4 ;
    output d_arr_21__3 ;
    output d_arr_21__2 ;
    output d_arr_21__1 ;
    output d_arr_21__0 ;
    output d_arr_22__31 ;
    output d_arr_22__30 ;
    output d_arr_22__29 ;
    output d_arr_22__28 ;
    output d_arr_22__27 ;
    output d_arr_22__26 ;
    output d_arr_22__25 ;
    output d_arr_22__24 ;
    output d_arr_22__23 ;
    output d_arr_22__22 ;
    output d_arr_22__21 ;
    output d_arr_22__20 ;
    output d_arr_22__19 ;
    output d_arr_22__18 ;
    output d_arr_22__17 ;
    output d_arr_22__16 ;
    output d_arr_22__15 ;
    output d_arr_22__14 ;
    output d_arr_22__13 ;
    output d_arr_22__12 ;
    output d_arr_22__11 ;
    output d_arr_22__10 ;
    output d_arr_22__9 ;
    output d_arr_22__8 ;
    output d_arr_22__7 ;
    output d_arr_22__6 ;
    output d_arr_22__5 ;
    output d_arr_22__4 ;
    output d_arr_22__3 ;
    output d_arr_22__2 ;
    output d_arr_22__1 ;
    output d_arr_22__0 ;
    output d_arr_23__31 ;
    output d_arr_23__30 ;
    output d_arr_23__29 ;
    output d_arr_23__28 ;
    output d_arr_23__27 ;
    output d_arr_23__26 ;
    output d_arr_23__25 ;
    output d_arr_23__24 ;
    output d_arr_23__23 ;
    output d_arr_23__22 ;
    output d_arr_23__21 ;
    output d_arr_23__20 ;
    output d_arr_23__19 ;
    output d_arr_23__18 ;
    output d_arr_23__17 ;
    output d_arr_23__16 ;
    output d_arr_23__15 ;
    output d_arr_23__14 ;
    output d_arr_23__13 ;
    output d_arr_23__12 ;
    output d_arr_23__11 ;
    output d_arr_23__10 ;
    output d_arr_23__9 ;
    output d_arr_23__8 ;
    output d_arr_23__7 ;
    output d_arr_23__6 ;
    output d_arr_23__5 ;
    output d_arr_23__4 ;
    output d_arr_23__3 ;
    output d_arr_23__2 ;
    output d_arr_23__1 ;
    output d_arr_23__0 ;
    output d_arr_24__31 ;
    output d_arr_24__30 ;
    output d_arr_24__29 ;
    output d_arr_24__28 ;
    output d_arr_24__27 ;
    output d_arr_24__26 ;
    output d_arr_24__25 ;
    output d_arr_24__24 ;
    output d_arr_24__23 ;
    output d_arr_24__22 ;
    output d_arr_24__21 ;
    output d_arr_24__20 ;
    output d_arr_24__19 ;
    output d_arr_24__18 ;
    output d_arr_24__17 ;
    output d_arr_24__16 ;
    output d_arr_24__15 ;
    output d_arr_24__14 ;
    output d_arr_24__13 ;
    output d_arr_24__12 ;
    output d_arr_24__11 ;
    output d_arr_24__10 ;
    output d_arr_24__9 ;
    output d_arr_24__8 ;
    output d_arr_24__7 ;
    output d_arr_24__6 ;
    output d_arr_24__5 ;
    output d_arr_24__4 ;
    output d_arr_24__3 ;
    output d_arr_24__2 ;
    output d_arr_24__1 ;
    output d_arr_24__0 ;
    input q_arr_0__31 ;
    input q_arr_0__30 ;
    input q_arr_0__29 ;
    input q_arr_0__28 ;
    input q_arr_0__27 ;
    input q_arr_0__26 ;
    input q_arr_0__25 ;
    input q_arr_0__24 ;
    input q_arr_0__23 ;
    input q_arr_0__22 ;
    input q_arr_0__21 ;
    input q_arr_0__20 ;
    input q_arr_0__19 ;
    input q_arr_0__18 ;
    input q_arr_0__17 ;
    input q_arr_0__16 ;
    input q_arr_0__15 ;
    input q_arr_0__14 ;
    input q_arr_0__13 ;
    input q_arr_0__12 ;
    input q_arr_0__11 ;
    input q_arr_0__10 ;
    input q_arr_0__9 ;
    input q_arr_0__8 ;
    input q_arr_0__7 ;
    input q_arr_0__6 ;
    input q_arr_0__5 ;
    input q_arr_0__4 ;
    input q_arr_0__3 ;
    input q_arr_0__2 ;
    input q_arr_0__1 ;
    input q_arr_0__0 ;
    input q_arr_1__31 ;
    input q_arr_1__30 ;
    input q_arr_1__29 ;
    input q_arr_1__28 ;
    input q_arr_1__27 ;
    input q_arr_1__26 ;
    input q_arr_1__25 ;
    input q_arr_1__24 ;
    input q_arr_1__23 ;
    input q_arr_1__22 ;
    input q_arr_1__21 ;
    input q_arr_1__20 ;
    input q_arr_1__19 ;
    input q_arr_1__18 ;
    input q_arr_1__17 ;
    input q_arr_1__16 ;
    input q_arr_1__15 ;
    input q_arr_1__14 ;
    input q_arr_1__13 ;
    input q_arr_1__12 ;
    input q_arr_1__11 ;
    input q_arr_1__10 ;
    input q_arr_1__9 ;
    input q_arr_1__8 ;
    input q_arr_1__7 ;
    input q_arr_1__6 ;
    input q_arr_1__5 ;
    input q_arr_1__4 ;
    input q_arr_1__3 ;
    input q_arr_1__2 ;
    input q_arr_1__1 ;
    input q_arr_1__0 ;
    input q_arr_2__31 ;
    input q_arr_2__30 ;
    input q_arr_2__29 ;
    input q_arr_2__28 ;
    input q_arr_2__27 ;
    input q_arr_2__26 ;
    input q_arr_2__25 ;
    input q_arr_2__24 ;
    input q_arr_2__23 ;
    input q_arr_2__22 ;
    input q_arr_2__21 ;
    input q_arr_2__20 ;
    input q_arr_2__19 ;
    input q_arr_2__18 ;
    input q_arr_2__17 ;
    input q_arr_2__16 ;
    input q_arr_2__15 ;
    input q_arr_2__14 ;
    input q_arr_2__13 ;
    input q_arr_2__12 ;
    input q_arr_2__11 ;
    input q_arr_2__10 ;
    input q_arr_2__9 ;
    input q_arr_2__8 ;
    input q_arr_2__7 ;
    input q_arr_2__6 ;
    input q_arr_2__5 ;
    input q_arr_2__4 ;
    input q_arr_2__3 ;
    input q_arr_2__2 ;
    input q_arr_2__1 ;
    input q_arr_2__0 ;
    input q_arr_3__31 ;
    input q_arr_3__30 ;
    input q_arr_3__29 ;
    input q_arr_3__28 ;
    input q_arr_3__27 ;
    input q_arr_3__26 ;
    input q_arr_3__25 ;
    input q_arr_3__24 ;
    input q_arr_3__23 ;
    input q_arr_3__22 ;
    input q_arr_3__21 ;
    input q_arr_3__20 ;
    input q_arr_3__19 ;
    input q_arr_3__18 ;
    input q_arr_3__17 ;
    input q_arr_3__16 ;
    input q_arr_3__15 ;
    input q_arr_3__14 ;
    input q_arr_3__13 ;
    input q_arr_3__12 ;
    input q_arr_3__11 ;
    input q_arr_3__10 ;
    input q_arr_3__9 ;
    input q_arr_3__8 ;
    input q_arr_3__7 ;
    input q_arr_3__6 ;
    input q_arr_3__5 ;
    input q_arr_3__4 ;
    input q_arr_3__3 ;
    input q_arr_3__2 ;
    input q_arr_3__1 ;
    input q_arr_3__0 ;
    input q_arr_4__31 ;
    input q_arr_4__30 ;
    input q_arr_4__29 ;
    input q_arr_4__28 ;
    input q_arr_4__27 ;
    input q_arr_4__26 ;
    input q_arr_4__25 ;
    input q_arr_4__24 ;
    input q_arr_4__23 ;
    input q_arr_4__22 ;
    input q_arr_4__21 ;
    input q_arr_4__20 ;
    input q_arr_4__19 ;
    input q_arr_4__18 ;
    input q_arr_4__17 ;
    input q_arr_4__16 ;
    input q_arr_4__15 ;
    input q_arr_4__14 ;
    input q_arr_4__13 ;
    input q_arr_4__12 ;
    input q_arr_4__11 ;
    input q_arr_4__10 ;
    input q_arr_4__9 ;
    input q_arr_4__8 ;
    input q_arr_4__7 ;
    input q_arr_4__6 ;
    input q_arr_4__5 ;
    input q_arr_4__4 ;
    input q_arr_4__3 ;
    input q_arr_4__2 ;
    input q_arr_4__1 ;
    input q_arr_4__0 ;
    input q_arr_5__31 ;
    input q_arr_5__30 ;
    input q_arr_5__29 ;
    input q_arr_5__28 ;
    input q_arr_5__27 ;
    input q_arr_5__26 ;
    input q_arr_5__25 ;
    input q_arr_5__24 ;
    input q_arr_5__23 ;
    input q_arr_5__22 ;
    input q_arr_5__21 ;
    input q_arr_5__20 ;
    input q_arr_5__19 ;
    input q_arr_5__18 ;
    input q_arr_5__17 ;
    input q_arr_5__16 ;
    input q_arr_5__15 ;
    input q_arr_5__14 ;
    input q_arr_5__13 ;
    input q_arr_5__12 ;
    input q_arr_5__11 ;
    input q_arr_5__10 ;
    input q_arr_5__9 ;
    input q_arr_5__8 ;
    input q_arr_5__7 ;
    input q_arr_5__6 ;
    input q_arr_5__5 ;
    input q_arr_5__4 ;
    input q_arr_5__3 ;
    input q_arr_5__2 ;
    input q_arr_5__1 ;
    input q_arr_5__0 ;
    input q_arr_6__31 ;
    input q_arr_6__30 ;
    input q_arr_6__29 ;
    input q_arr_6__28 ;
    input q_arr_6__27 ;
    input q_arr_6__26 ;
    input q_arr_6__25 ;
    input q_arr_6__24 ;
    input q_arr_6__23 ;
    input q_arr_6__22 ;
    input q_arr_6__21 ;
    input q_arr_6__20 ;
    input q_arr_6__19 ;
    input q_arr_6__18 ;
    input q_arr_6__17 ;
    input q_arr_6__16 ;
    input q_arr_6__15 ;
    input q_arr_6__14 ;
    input q_arr_6__13 ;
    input q_arr_6__12 ;
    input q_arr_6__11 ;
    input q_arr_6__10 ;
    input q_arr_6__9 ;
    input q_arr_6__8 ;
    input q_arr_6__7 ;
    input q_arr_6__6 ;
    input q_arr_6__5 ;
    input q_arr_6__4 ;
    input q_arr_6__3 ;
    input q_arr_6__2 ;
    input q_arr_6__1 ;
    input q_arr_6__0 ;
    input q_arr_7__31 ;
    input q_arr_7__30 ;
    input q_arr_7__29 ;
    input q_arr_7__28 ;
    input q_arr_7__27 ;
    input q_arr_7__26 ;
    input q_arr_7__25 ;
    input q_arr_7__24 ;
    input q_arr_7__23 ;
    input q_arr_7__22 ;
    input q_arr_7__21 ;
    input q_arr_7__20 ;
    input q_arr_7__19 ;
    input q_arr_7__18 ;
    input q_arr_7__17 ;
    input q_arr_7__16 ;
    input q_arr_7__15 ;
    input q_arr_7__14 ;
    input q_arr_7__13 ;
    input q_arr_7__12 ;
    input q_arr_7__11 ;
    input q_arr_7__10 ;
    input q_arr_7__9 ;
    input q_arr_7__8 ;
    input q_arr_7__7 ;
    input q_arr_7__6 ;
    input q_arr_7__5 ;
    input q_arr_7__4 ;
    input q_arr_7__3 ;
    input q_arr_7__2 ;
    input q_arr_7__1 ;
    input q_arr_7__0 ;
    input q_arr_8__31 ;
    input q_arr_8__30 ;
    input q_arr_8__29 ;
    input q_arr_8__28 ;
    input q_arr_8__27 ;
    input q_arr_8__26 ;
    input q_arr_8__25 ;
    input q_arr_8__24 ;
    input q_arr_8__23 ;
    input q_arr_8__22 ;
    input q_arr_8__21 ;
    input q_arr_8__20 ;
    input q_arr_8__19 ;
    input q_arr_8__18 ;
    input q_arr_8__17 ;
    input q_arr_8__16 ;
    input q_arr_8__15 ;
    input q_arr_8__14 ;
    input q_arr_8__13 ;
    input q_arr_8__12 ;
    input q_arr_8__11 ;
    input q_arr_8__10 ;
    input q_arr_8__9 ;
    input q_arr_8__8 ;
    input q_arr_8__7 ;
    input q_arr_8__6 ;
    input q_arr_8__5 ;
    input q_arr_8__4 ;
    input q_arr_8__3 ;
    input q_arr_8__2 ;
    input q_arr_8__1 ;
    input q_arr_8__0 ;
    input q_arr_9__31 ;
    input q_arr_9__30 ;
    input q_arr_9__29 ;
    input q_arr_9__28 ;
    input q_arr_9__27 ;
    input q_arr_9__26 ;
    input q_arr_9__25 ;
    input q_arr_9__24 ;
    input q_arr_9__23 ;
    input q_arr_9__22 ;
    input q_arr_9__21 ;
    input q_arr_9__20 ;
    input q_arr_9__19 ;
    input q_arr_9__18 ;
    input q_arr_9__17 ;
    input q_arr_9__16 ;
    input q_arr_9__15 ;
    input q_arr_9__14 ;
    input q_arr_9__13 ;
    input q_arr_9__12 ;
    input q_arr_9__11 ;
    input q_arr_9__10 ;
    input q_arr_9__9 ;
    input q_arr_9__8 ;
    input q_arr_9__7 ;
    input q_arr_9__6 ;
    input q_arr_9__5 ;
    input q_arr_9__4 ;
    input q_arr_9__3 ;
    input q_arr_9__2 ;
    input q_arr_9__1 ;
    input q_arr_9__0 ;
    input q_arr_10__31 ;
    input q_arr_10__30 ;
    input q_arr_10__29 ;
    input q_arr_10__28 ;
    input q_arr_10__27 ;
    input q_arr_10__26 ;
    input q_arr_10__25 ;
    input q_arr_10__24 ;
    input q_arr_10__23 ;
    input q_arr_10__22 ;
    input q_arr_10__21 ;
    input q_arr_10__20 ;
    input q_arr_10__19 ;
    input q_arr_10__18 ;
    input q_arr_10__17 ;
    input q_arr_10__16 ;
    input q_arr_10__15 ;
    input q_arr_10__14 ;
    input q_arr_10__13 ;
    input q_arr_10__12 ;
    input q_arr_10__11 ;
    input q_arr_10__10 ;
    input q_arr_10__9 ;
    input q_arr_10__8 ;
    input q_arr_10__7 ;
    input q_arr_10__6 ;
    input q_arr_10__5 ;
    input q_arr_10__4 ;
    input q_arr_10__3 ;
    input q_arr_10__2 ;
    input q_arr_10__1 ;
    input q_arr_10__0 ;
    input q_arr_11__31 ;
    input q_arr_11__30 ;
    input q_arr_11__29 ;
    input q_arr_11__28 ;
    input q_arr_11__27 ;
    input q_arr_11__26 ;
    input q_arr_11__25 ;
    input q_arr_11__24 ;
    input q_arr_11__23 ;
    input q_arr_11__22 ;
    input q_arr_11__21 ;
    input q_arr_11__20 ;
    input q_arr_11__19 ;
    input q_arr_11__18 ;
    input q_arr_11__17 ;
    input q_arr_11__16 ;
    input q_arr_11__15 ;
    input q_arr_11__14 ;
    input q_arr_11__13 ;
    input q_arr_11__12 ;
    input q_arr_11__11 ;
    input q_arr_11__10 ;
    input q_arr_11__9 ;
    input q_arr_11__8 ;
    input q_arr_11__7 ;
    input q_arr_11__6 ;
    input q_arr_11__5 ;
    input q_arr_11__4 ;
    input q_arr_11__3 ;
    input q_arr_11__2 ;
    input q_arr_11__1 ;
    input q_arr_11__0 ;
    input q_arr_12__31 ;
    input q_arr_12__30 ;
    input q_arr_12__29 ;
    input q_arr_12__28 ;
    input q_arr_12__27 ;
    input q_arr_12__26 ;
    input q_arr_12__25 ;
    input q_arr_12__24 ;
    input q_arr_12__23 ;
    input q_arr_12__22 ;
    input q_arr_12__21 ;
    input q_arr_12__20 ;
    input q_arr_12__19 ;
    input q_arr_12__18 ;
    input q_arr_12__17 ;
    input q_arr_12__16 ;
    input q_arr_12__15 ;
    input q_arr_12__14 ;
    input q_arr_12__13 ;
    input q_arr_12__12 ;
    input q_arr_12__11 ;
    input q_arr_12__10 ;
    input q_arr_12__9 ;
    input q_arr_12__8 ;
    input q_arr_12__7 ;
    input q_arr_12__6 ;
    input q_arr_12__5 ;
    input q_arr_12__4 ;
    input q_arr_12__3 ;
    input q_arr_12__2 ;
    input q_arr_12__1 ;
    input q_arr_12__0 ;
    input q_arr_13__31 ;
    input q_arr_13__30 ;
    input q_arr_13__29 ;
    input q_arr_13__28 ;
    input q_arr_13__27 ;
    input q_arr_13__26 ;
    input q_arr_13__25 ;
    input q_arr_13__24 ;
    input q_arr_13__23 ;
    input q_arr_13__22 ;
    input q_arr_13__21 ;
    input q_arr_13__20 ;
    input q_arr_13__19 ;
    input q_arr_13__18 ;
    input q_arr_13__17 ;
    input q_arr_13__16 ;
    input q_arr_13__15 ;
    input q_arr_13__14 ;
    input q_arr_13__13 ;
    input q_arr_13__12 ;
    input q_arr_13__11 ;
    input q_arr_13__10 ;
    input q_arr_13__9 ;
    input q_arr_13__8 ;
    input q_arr_13__7 ;
    input q_arr_13__6 ;
    input q_arr_13__5 ;
    input q_arr_13__4 ;
    input q_arr_13__3 ;
    input q_arr_13__2 ;
    input q_arr_13__1 ;
    input q_arr_13__0 ;
    input q_arr_14__31 ;
    input q_arr_14__30 ;
    input q_arr_14__29 ;
    input q_arr_14__28 ;
    input q_arr_14__27 ;
    input q_arr_14__26 ;
    input q_arr_14__25 ;
    input q_arr_14__24 ;
    input q_arr_14__23 ;
    input q_arr_14__22 ;
    input q_arr_14__21 ;
    input q_arr_14__20 ;
    input q_arr_14__19 ;
    input q_arr_14__18 ;
    input q_arr_14__17 ;
    input q_arr_14__16 ;
    input q_arr_14__15 ;
    input q_arr_14__14 ;
    input q_arr_14__13 ;
    input q_arr_14__12 ;
    input q_arr_14__11 ;
    input q_arr_14__10 ;
    input q_arr_14__9 ;
    input q_arr_14__8 ;
    input q_arr_14__7 ;
    input q_arr_14__6 ;
    input q_arr_14__5 ;
    input q_arr_14__4 ;
    input q_arr_14__3 ;
    input q_arr_14__2 ;
    input q_arr_14__1 ;
    input q_arr_14__0 ;
    input q_arr_15__31 ;
    input q_arr_15__30 ;
    input q_arr_15__29 ;
    input q_arr_15__28 ;
    input q_arr_15__27 ;
    input q_arr_15__26 ;
    input q_arr_15__25 ;
    input q_arr_15__24 ;
    input q_arr_15__23 ;
    input q_arr_15__22 ;
    input q_arr_15__21 ;
    input q_arr_15__20 ;
    input q_arr_15__19 ;
    input q_arr_15__18 ;
    input q_arr_15__17 ;
    input q_arr_15__16 ;
    input q_arr_15__15 ;
    input q_arr_15__14 ;
    input q_arr_15__13 ;
    input q_arr_15__12 ;
    input q_arr_15__11 ;
    input q_arr_15__10 ;
    input q_arr_15__9 ;
    input q_arr_15__8 ;
    input q_arr_15__7 ;
    input q_arr_15__6 ;
    input q_arr_15__5 ;
    input q_arr_15__4 ;
    input q_arr_15__3 ;
    input q_arr_15__2 ;
    input q_arr_15__1 ;
    input q_arr_15__0 ;
    input q_arr_16__31 ;
    input q_arr_16__30 ;
    input q_arr_16__29 ;
    input q_arr_16__28 ;
    input q_arr_16__27 ;
    input q_arr_16__26 ;
    input q_arr_16__25 ;
    input q_arr_16__24 ;
    input q_arr_16__23 ;
    input q_arr_16__22 ;
    input q_arr_16__21 ;
    input q_arr_16__20 ;
    input q_arr_16__19 ;
    input q_arr_16__18 ;
    input q_arr_16__17 ;
    input q_arr_16__16 ;
    input q_arr_16__15 ;
    input q_arr_16__14 ;
    input q_arr_16__13 ;
    input q_arr_16__12 ;
    input q_arr_16__11 ;
    input q_arr_16__10 ;
    input q_arr_16__9 ;
    input q_arr_16__8 ;
    input q_arr_16__7 ;
    input q_arr_16__6 ;
    input q_arr_16__5 ;
    input q_arr_16__4 ;
    input q_arr_16__3 ;
    input q_arr_16__2 ;
    input q_arr_16__1 ;
    input q_arr_16__0 ;
    input q_arr_17__31 ;
    input q_arr_17__30 ;
    input q_arr_17__29 ;
    input q_arr_17__28 ;
    input q_arr_17__27 ;
    input q_arr_17__26 ;
    input q_arr_17__25 ;
    input q_arr_17__24 ;
    input q_arr_17__23 ;
    input q_arr_17__22 ;
    input q_arr_17__21 ;
    input q_arr_17__20 ;
    input q_arr_17__19 ;
    input q_arr_17__18 ;
    input q_arr_17__17 ;
    input q_arr_17__16 ;
    input q_arr_17__15 ;
    input q_arr_17__14 ;
    input q_arr_17__13 ;
    input q_arr_17__12 ;
    input q_arr_17__11 ;
    input q_arr_17__10 ;
    input q_arr_17__9 ;
    input q_arr_17__8 ;
    input q_arr_17__7 ;
    input q_arr_17__6 ;
    input q_arr_17__5 ;
    input q_arr_17__4 ;
    input q_arr_17__3 ;
    input q_arr_17__2 ;
    input q_arr_17__1 ;
    input q_arr_17__0 ;
    input q_arr_18__31 ;
    input q_arr_18__30 ;
    input q_arr_18__29 ;
    input q_arr_18__28 ;
    input q_arr_18__27 ;
    input q_arr_18__26 ;
    input q_arr_18__25 ;
    input q_arr_18__24 ;
    input q_arr_18__23 ;
    input q_arr_18__22 ;
    input q_arr_18__21 ;
    input q_arr_18__20 ;
    input q_arr_18__19 ;
    input q_arr_18__18 ;
    input q_arr_18__17 ;
    input q_arr_18__16 ;
    input q_arr_18__15 ;
    input q_arr_18__14 ;
    input q_arr_18__13 ;
    input q_arr_18__12 ;
    input q_arr_18__11 ;
    input q_arr_18__10 ;
    input q_arr_18__9 ;
    input q_arr_18__8 ;
    input q_arr_18__7 ;
    input q_arr_18__6 ;
    input q_arr_18__5 ;
    input q_arr_18__4 ;
    input q_arr_18__3 ;
    input q_arr_18__2 ;
    input q_arr_18__1 ;
    input q_arr_18__0 ;
    input q_arr_19__31 ;
    input q_arr_19__30 ;
    input q_arr_19__29 ;
    input q_arr_19__28 ;
    input q_arr_19__27 ;
    input q_arr_19__26 ;
    input q_arr_19__25 ;
    input q_arr_19__24 ;
    input q_arr_19__23 ;
    input q_arr_19__22 ;
    input q_arr_19__21 ;
    input q_arr_19__20 ;
    input q_arr_19__19 ;
    input q_arr_19__18 ;
    input q_arr_19__17 ;
    input q_arr_19__16 ;
    input q_arr_19__15 ;
    input q_arr_19__14 ;
    input q_arr_19__13 ;
    input q_arr_19__12 ;
    input q_arr_19__11 ;
    input q_arr_19__10 ;
    input q_arr_19__9 ;
    input q_arr_19__8 ;
    input q_arr_19__7 ;
    input q_arr_19__6 ;
    input q_arr_19__5 ;
    input q_arr_19__4 ;
    input q_arr_19__3 ;
    input q_arr_19__2 ;
    input q_arr_19__1 ;
    input q_arr_19__0 ;
    input q_arr_20__31 ;
    input q_arr_20__30 ;
    input q_arr_20__29 ;
    input q_arr_20__28 ;
    input q_arr_20__27 ;
    input q_arr_20__26 ;
    input q_arr_20__25 ;
    input q_arr_20__24 ;
    input q_arr_20__23 ;
    input q_arr_20__22 ;
    input q_arr_20__21 ;
    input q_arr_20__20 ;
    input q_arr_20__19 ;
    input q_arr_20__18 ;
    input q_arr_20__17 ;
    input q_arr_20__16 ;
    input q_arr_20__15 ;
    input q_arr_20__14 ;
    input q_arr_20__13 ;
    input q_arr_20__12 ;
    input q_arr_20__11 ;
    input q_arr_20__10 ;
    input q_arr_20__9 ;
    input q_arr_20__8 ;
    input q_arr_20__7 ;
    input q_arr_20__6 ;
    input q_arr_20__5 ;
    input q_arr_20__4 ;
    input q_arr_20__3 ;
    input q_arr_20__2 ;
    input q_arr_20__1 ;
    input q_arr_20__0 ;
    input q_arr_21__31 ;
    input q_arr_21__30 ;
    input q_arr_21__29 ;
    input q_arr_21__28 ;
    input q_arr_21__27 ;
    input q_arr_21__26 ;
    input q_arr_21__25 ;
    input q_arr_21__24 ;
    input q_arr_21__23 ;
    input q_arr_21__22 ;
    input q_arr_21__21 ;
    input q_arr_21__20 ;
    input q_arr_21__19 ;
    input q_arr_21__18 ;
    input q_arr_21__17 ;
    input q_arr_21__16 ;
    input q_arr_21__15 ;
    input q_arr_21__14 ;
    input q_arr_21__13 ;
    input q_arr_21__12 ;
    input q_arr_21__11 ;
    input q_arr_21__10 ;
    input q_arr_21__9 ;
    input q_arr_21__8 ;
    input q_arr_21__7 ;
    input q_arr_21__6 ;
    input q_arr_21__5 ;
    input q_arr_21__4 ;
    input q_arr_21__3 ;
    input q_arr_21__2 ;
    input q_arr_21__1 ;
    input q_arr_21__0 ;
    input q_arr_22__31 ;
    input q_arr_22__30 ;
    input q_arr_22__29 ;
    input q_arr_22__28 ;
    input q_arr_22__27 ;
    input q_arr_22__26 ;
    input q_arr_22__25 ;
    input q_arr_22__24 ;
    input q_arr_22__23 ;
    input q_arr_22__22 ;
    input q_arr_22__21 ;
    input q_arr_22__20 ;
    input q_arr_22__19 ;
    input q_arr_22__18 ;
    input q_arr_22__17 ;
    input q_arr_22__16 ;
    input q_arr_22__15 ;
    input q_arr_22__14 ;
    input q_arr_22__13 ;
    input q_arr_22__12 ;
    input q_arr_22__11 ;
    input q_arr_22__10 ;
    input q_arr_22__9 ;
    input q_arr_22__8 ;
    input q_arr_22__7 ;
    input q_arr_22__6 ;
    input q_arr_22__5 ;
    input q_arr_22__4 ;
    input q_arr_22__3 ;
    input q_arr_22__2 ;
    input q_arr_22__1 ;
    input q_arr_22__0 ;
    input q_arr_23__31 ;
    input q_arr_23__30 ;
    input q_arr_23__29 ;
    input q_arr_23__28 ;
    input q_arr_23__27 ;
    input q_arr_23__26 ;
    input q_arr_23__25 ;
    input q_arr_23__24 ;
    input q_arr_23__23 ;
    input q_arr_23__22 ;
    input q_arr_23__21 ;
    input q_arr_23__20 ;
    input q_arr_23__19 ;
    input q_arr_23__18 ;
    input q_arr_23__17 ;
    input q_arr_23__16 ;
    input q_arr_23__15 ;
    input q_arr_23__14 ;
    input q_arr_23__13 ;
    input q_arr_23__12 ;
    input q_arr_23__11 ;
    input q_arr_23__10 ;
    input q_arr_23__9 ;
    input q_arr_23__8 ;
    input q_arr_23__7 ;
    input q_arr_23__6 ;
    input q_arr_23__5 ;
    input q_arr_23__4 ;
    input q_arr_23__3 ;
    input q_arr_23__2 ;
    input q_arr_23__1 ;
    input q_arr_23__0 ;
    input q_arr_24__31 ;
    input q_arr_24__30 ;
    input q_arr_24__29 ;
    input q_arr_24__28 ;
    input q_arr_24__27 ;
    input q_arr_24__26 ;
    input q_arr_24__25 ;
    input q_arr_24__24 ;
    input q_arr_24__23 ;
    input q_arr_24__22 ;
    input q_arr_24__21 ;
    input q_arr_24__20 ;
    input q_arr_24__19 ;
    input q_arr_24__18 ;
    input q_arr_24__17 ;
    input q_arr_24__16 ;
    input q_arr_24__15 ;
    input q_arr_24__14 ;
    input q_arr_24__13 ;
    input q_arr_24__12 ;
    input q_arr_24__11 ;
    input q_arr_24__10 ;
    input q_arr_24__9 ;
    input q_arr_24__8 ;
    input q_arr_24__7 ;
    input q_arr_24__6 ;
    input q_arr_24__5 ;
    input q_arr_24__4 ;
    input q_arr_24__3 ;
    input q_arr_24__2 ;
    input q_arr_24__1 ;
    input q_arr_24__0 ;
    input operation ;
    input filter_size ;

    wire s1_31, s1_30, s1_29, s1_28, s1_27, s1_26, s1_25, s1_24, s1_23, s1_22, 
         s1_21, s1_20, s1_19, s1_18, s1_17, s1_16, s1_15, s1_14, s1_13, s1_12, 
         s1_11, s1_10, s1_9, s1_8, s1_7, s1_6, s1_5, s1_4, s1_3, s1_2, s1_1, 
         s1_0, s2_31, s2_30, s2_29, s2_28, s2_27, s2_26, s2_25, s2_24, s2_23, 
         s2_22, s2_21, s2_20, s2_19, s2_18, s2_17, s2_16, s2_15, s2_14, s2_13, 
         s2_12, s2_11, s2_10, s2_9, s2_8, s2_7, s2_6, s2_5, s2_4, s2_3, s2_2, 
         s2_1, s2_0, nx6, nx10, nx350, nx153, nx165, nx169, nx173, nx177, nx181, 
         nx185, nx189, nx193, nx197, nx201, nx205, nx209, nx213, nx217, nx221, 
         nx225, nx229, nx233, nx237, nx241, nx245, nx249, nx253, nx257, nx261, 
         nx265, nx277, nx279, nx285, nx287, nx291, nx293, nx297, nx299, nx303, 
         nx305, nx309, nx311, nx315, nx317, nx321, nx323, nx327, nx329, nx333, 
         nx335, nx339, nx341, nx345, nx347, nx351, nx353, nx357, nx359, nx363, 
         nx365, nx369, nx371, nx375, nx377, nx381, nx383, nx387, nx389, nx393, 
         nx395, nx399, nx401, nx405, nx407, nx411, nx413, nx417, nx419, nx423, 
         nx425, nx429, nx431, nx435, nx437, nx441, nx445, nx458, nx460, nx462, 
         nx464, nx466, nx469, nx471, nx473, nx475, nx477, nx479, nx481, nx483, 
         nx485, nx487, nx489, nx491, nx493, nx495, nx497, nx499, nx501, nx503, 
         nx505, nx507, nx509, nx511, nx513, nx515, nx517, nx519, nx521, nx523, 
         nx525, nx527, nx529, nx531, nx533, nx540, nx542, nx550, nx553, nx555;
    wire [1:0] \$dummy ;




    assign d_arr_2__30 = d_arr_2__31 ;
    assign d_arr_2__29 = d_arr_2__31 ;
    assign d_arr_2__28 = d_arr_2__31 ;
    assign d_arr_2__27 = d_arr_2__31 ;
    assign d_arr_2__26 = d_arr_2__31 ;
    assign d_arr_2__25 = d_arr_2__31 ;
    assign d_arr_2__24 = d_arr_2__31 ;
    assign d_arr_2__23 = d_arr_2__31 ;
    assign d_arr_2__22 = d_arr_2__31 ;
    assign d_arr_2__21 = d_arr_2__31 ;
    assign d_arr_2__20 = d_arr_2__31 ;
    assign d_arr_2__19 = d_arr_2__31 ;
    assign d_arr_2__18 = d_arr_2__31 ;
    assign d_arr_2__17 = d_arr_2__31 ;
    assign d_arr_2__16 = d_arr_2__31 ;
    assign d_arr_2__15 = d_arr_2__31 ;
    assign d_arr_2__14 = d_arr_2__31 ;
    assign d_arr_2__13 = d_arr_2__31 ;
    assign d_arr_2__12 = d_arr_2__31 ;
    assign d_arr_2__11 = d_arr_2__31 ;
    assign d_arr_2__10 = d_arr_2__31 ;
    assign d_arr_2__9 = d_arr_2__31 ;
    assign d_arr_2__8 = d_arr_2__31 ;
    assign d_arr_2__7 = d_arr_2__31 ;
    assign d_arr_2__6 = d_arr_2__31 ;
    assign d_arr_2__5 = d_arr_2__31 ;
    assign d_arr_2__4 = d_arr_2__31 ;
    assign d_arr_2__3 = d_arr_2__31 ;
    assign d_arr_2__2 = d_arr_2__31 ;
    assign d_arr_2__1 = d_arr_2__31 ;
    assign d_arr_2__0 = d_arr_2__31 ;
    assign d_arr_3__31 = d_arr_2__31 ;
    assign d_arr_3__30 = d_arr_2__31 ;
    assign d_arr_3__29 = d_arr_2__31 ;
    assign d_arr_3__28 = d_arr_2__31 ;
    assign d_arr_3__27 = d_arr_2__31 ;
    assign d_arr_3__26 = d_arr_2__31 ;
    assign d_arr_3__25 = d_arr_2__31 ;
    assign d_arr_3__24 = d_arr_2__31 ;
    assign d_arr_3__23 = d_arr_2__31 ;
    assign d_arr_3__22 = d_arr_2__31 ;
    assign d_arr_3__21 = d_arr_2__31 ;
    assign d_arr_3__20 = d_arr_2__31 ;
    assign d_arr_3__19 = d_arr_2__31 ;
    assign d_arr_3__18 = d_arr_2__31 ;
    assign d_arr_3__17 = d_arr_2__31 ;
    assign d_arr_3__16 = d_arr_2__31 ;
    assign d_arr_3__15 = d_arr_2__31 ;
    assign d_arr_3__14 = d_arr_2__31 ;
    assign d_arr_3__13 = d_arr_2__31 ;
    assign d_arr_3__12 = d_arr_2__31 ;
    assign d_arr_3__11 = d_arr_2__31 ;
    assign d_arr_3__10 = d_arr_2__31 ;
    assign d_arr_3__9 = d_arr_2__31 ;
    assign d_arr_3__8 = d_arr_2__31 ;
    assign d_arr_3__7 = d_arr_2__31 ;
    assign d_arr_3__6 = d_arr_2__31 ;
    assign d_arr_3__5 = d_arr_2__31 ;
    assign d_arr_3__4 = d_arr_2__31 ;
    assign d_arr_3__3 = d_arr_2__31 ;
    assign d_arr_3__2 = d_arr_2__31 ;
    assign d_arr_3__1 = d_arr_2__31 ;
    assign d_arr_3__0 = d_arr_2__31 ;
    assign d_arr_4__31 = d_arr_2__31 ;
    assign d_arr_4__30 = d_arr_2__31 ;
    assign d_arr_4__29 = d_arr_2__31 ;
    assign d_arr_4__28 = d_arr_2__31 ;
    assign d_arr_4__27 = d_arr_2__31 ;
    assign d_arr_4__26 = d_arr_2__31 ;
    assign d_arr_4__25 = d_arr_2__31 ;
    assign d_arr_4__24 = d_arr_2__31 ;
    assign d_arr_4__23 = d_arr_2__31 ;
    assign d_arr_4__22 = d_arr_2__31 ;
    assign d_arr_4__21 = d_arr_2__31 ;
    assign d_arr_4__20 = d_arr_2__31 ;
    assign d_arr_4__19 = d_arr_2__31 ;
    assign d_arr_4__18 = d_arr_2__31 ;
    assign d_arr_4__17 = d_arr_2__31 ;
    assign d_arr_4__16 = d_arr_2__31 ;
    assign d_arr_4__15 = d_arr_2__31 ;
    assign d_arr_4__14 = d_arr_2__31 ;
    assign d_arr_4__13 = d_arr_2__31 ;
    assign d_arr_4__12 = d_arr_2__31 ;
    assign d_arr_4__11 = d_arr_2__31 ;
    assign d_arr_4__10 = d_arr_2__31 ;
    assign d_arr_4__9 = d_arr_2__31 ;
    assign d_arr_4__8 = d_arr_2__31 ;
    assign d_arr_4__7 = d_arr_2__31 ;
    assign d_arr_4__6 = d_arr_2__31 ;
    assign d_arr_4__5 = d_arr_2__31 ;
    assign d_arr_4__4 = d_arr_2__31 ;
    assign d_arr_4__3 = d_arr_2__31 ;
    assign d_arr_4__2 = d_arr_2__31 ;
    assign d_arr_4__1 = d_arr_2__31 ;
    assign d_arr_4__0 = d_arr_2__31 ;
    assign d_arr_5__31 = d_arr_2__31 ;
    assign d_arr_5__30 = d_arr_2__31 ;
    assign d_arr_5__29 = d_arr_2__31 ;
    assign d_arr_5__28 = d_arr_2__31 ;
    assign d_arr_5__27 = d_arr_2__31 ;
    assign d_arr_5__26 = d_arr_2__31 ;
    assign d_arr_5__25 = d_arr_2__31 ;
    assign d_arr_5__24 = d_arr_2__31 ;
    assign d_arr_5__23 = d_arr_2__31 ;
    assign d_arr_5__22 = d_arr_2__31 ;
    assign d_arr_5__21 = d_arr_2__31 ;
    assign d_arr_5__20 = d_arr_2__31 ;
    assign d_arr_5__19 = d_arr_2__31 ;
    assign d_arr_5__18 = d_arr_2__31 ;
    assign d_arr_5__17 = d_arr_2__31 ;
    assign d_arr_5__16 = d_arr_2__31 ;
    assign d_arr_5__15 = d_arr_2__31 ;
    assign d_arr_5__14 = d_arr_2__31 ;
    assign d_arr_5__13 = d_arr_2__31 ;
    assign d_arr_5__12 = d_arr_2__31 ;
    assign d_arr_5__11 = d_arr_2__31 ;
    assign d_arr_5__10 = d_arr_2__31 ;
    assign d_arr_5__9 = d_arr_2__31 ;
    assign d_arr_5__8 = d_arr_2__31 ;
    assign d_arr_5__7 = d_arr_2__31 ;
    assign d_arr_5__6 = d_arr_2__31 ;
    assign d_arr_5__5 = d_arr_2__31 ;
    assign d_arr_5__4 = d_arr_2__31 ;
    assign d_arr_5__3 = d_arr_2__31 ;
    assign d_arr_5__2 = d_arr_2__31 ;
    assign d_arr_5__1 = d_arr_2__31 ;
    assign d_arr_5__0 = d_arr_2__31 ;
    assign d_arr_6__31 = d_arr_2__31 ;
    assign d_arr_6__30 = d_arr_2__31 ;
    assign d_arr_6__29 = d_arr_2__31 ;
    assign d_arr_6__28 = d_arr_2__31 ;
    assign d_arr_6__27 = d_arr_2__31 ;
    assign d_arr_6__26 = d_arr_2__31 ;
    assign d_arr_6__25 = d_arr_2__31 ;
    assign d_arr_6__24 = d_arr_2__31 ;
    assign d_arr_6__23 = d_arr_2__31 ;
    assign d_arr_6__22 = d_arr_2__31 ;
    assign d_arr_6__21 = d_arr_2__31 ;
    assign d_arr_6__20 = d_arr_2__31 ;
    assign d_arr_6__19 = d_arr_2__31 ;
    assign d_arr_6__18 = d_arr_2__31 ;
    assign d_arr_6__17 = d_arr_2__31 ;
    assign d_arr_6__16 = d_arr_2__31 ;
    assign d_arr_6__15 = d_arr_2__31 ;
    assign d_arr_6__14 = d_arr_2__31 ;
    assign d_arr_6__13 = d_arr_2__31 ;
    assign d_arr_6__12 = d_arr_2__31 ;
    assign d_arr_6__11 = d_arr_2__31 ;
    assign d_arr_6__10 = d_arr_2__31 ;
    assign d_arr_6__9 = d_arr_2__31 ;
    assign d_arr_6__8 = d_arr_2__31 ;
    assign d_arr_6__7 = d_arr_2__31 ;
    assign d_arr_6__6 = d_arr_2__31 ;
    assign d_arr_6__5 = d_arr_2__31 ;
    assign d_arr_6__4 = d_arr_2__31 ;
    assign d_arr_6__3 = d_arr_2__31 ;
    assign d_arr_6__2 = d_arr_2__31 ;
    assign d_arr_6__1 = d_arr_2__31 ;
    assign d_arr_6__0 = d_arr_2__31 ;
    assign d_arr_7__31 = d_arr_2__31 ;
    assign d_arr_7__30 = d_arr_2__31 ;
    assign d_arr_7__29 = d_arr_2__31 ;
    assign d_arr_7__28 = d_arr_2__31 ;
    assign d_arr_7__27 = d_arr_2__31 ;
    assign d_arr_7__26 = d_arr_2__31 ;
    assign d_arr_7__25 = d_arr_2__31 ;
    assign d_arr_7__24 = d_arr_2__31 ;
    assign d_arr_7__23 = d_arr_2__31 ;
    assign d_arr_7__22 = d_arr_2__31 ;
    assign d_arr_7__21 = d_arr_2__31 ;
    assign d_arr_7__20 = d_arr_2__31 ;
    assign d_arr_7__19 = d_arr_2__31 ;
    assign d_arr_7__18 = d_arr_2__31 ;
    assign d_arr_7__17 = d_arr_2__31 ;
    assign d_arr_7__16 = d_arr_2__31 ;
    assign d_arr_7__15 = d_arr_2__31 ;
    assign d_arr_7__14 = d_arr_2__31 ;
    assign d_arr_7__13 = d_arr_2__31 ;
    assign d_arr_7__12 = d_arr_2__31 ;
    assign d_arr_7__11 = d_arr_2__31 ;
    assign d_arr_7__10 = d_arr_2__31 ;
    assign d_arr_7__9 = d_arr_2__31 ;
    assign d_arr_7__8 = d_arr_2__31 ;
    assign d_arr_7__7 = d_arr_2__31 ;
    assign d_arr_7__6 = d_arr_2__31 ;
    assign d_arr_7__5 = d_arr_2__31 ;
    assign d_arr_7__4 = d_arr_2__31 ;
    assign d_arr_7__3 = d_arr_2__31 ;
    assign d_arr_7__2 = d_arr_2__31 ;
    assign d_arr_7__1 = d_arr_2__31 ;
    assign d_arr_7__0 = d_arr_2__31 ;
    assign d_arr_8__31 = d_arr_2__31 ;
    assign d_arr_8__30 = d_arr_2__31 ;
    assign d_arr_8__29 = d_arr_2__31 ;
    assign d_arr_8__28 = d_arr_2__31 ;
    assign d_arr_8__27 = d_arr_2__31 ;
    assign d_arr_8__26 = d_arr_2__31 ;
    assign d_arr_8__25 = d_arr_2__31 ;
    assign d_arr_8__24 = d_arr_2__31 ;
    assign d_arr_8__23 = d_arr_2__31 ;
    assign d_arr_8__22 = d_arr_2__31 ;
    assign d_arr_8__21 = d_arr_2__31 ;
    assign d_arr_8__20 = d_arr_2__31 ;
    assign d_arr_8__19 = d_arr_2__31 ;
    assign d_arr_8__18 = d_arr_2__31 ;
    assign d_arr_8__17 = d_arr_2__31 ;
    assign d_arr_8__16 = d_arr_2__31 ;
    assign d_arr_8__15 = d_arr_2__31 ;
    assign d_arr_8__14 = d_arr_2__31 ;
    assign d_arr_8__13 = d_arr_2__31 ;
    assign d_arr_8__12 = d_arr_2__31 ;
    assign d_arr_8__11 = d_arr_2__31 ;
    assign d_arr_8__10 = d_arr_2__31 ;
    assign d_arr_8__9 = d_arr_2__31 ;
    assign d_arr_8__8 = d_arr_2__31 ;
    assign d_arr_8__7 = d_arr_2__31 ;
    assign d_arr_8__6 = d_arr_2__31 ;
    assign d_arr_8__5 = d_arr_2__31 ;
    assign d_arr_8__4 = d_arr_2__31 ;
    assign d_arr_8__3 = d_arr_2__31 ;
    assign d_arr_8__2 = d_arr_2__31 ;
    assign d_arr_8__1 = d_arr_2__31 ;
    assign d_arr_8__0 = d_arr_2__31 ;
    assign d_arr_9__31 = d_arr_2__31 ;
    assign d_arr_9__30 = d_arr_2__31 ;
    assign d_arr_9__29 = d_arr_2__31 ;
    assign d_arr_9__28 = d_arr_2__31 ;
    assign d_arr_9__27 = d_arr_2__31 ;
    assign d_arr_9__26 = d_arr_2__31 ;
    assign d_arr_9__25 = d_arr_2__31 ;
    assign d_arr_9__24 = d_arr_2__31 ;
    assign d_arr_9__23 = d_arr_2__31 ;
    assign d_arr_9__22 = d_arr_2__31 ;
    assign d_arr_9__21 = d_arr_2__31 ;
    assign d_arr_9__20 = d_arr_2__31 ;
    assign d_arr_9__19 = d_arr_2__31 ;
    assign d_arr_9__18 = d_arr_2__31 ;
    assign d_arr_9__17 = d_arr_2__31 ;
    assign d_arr_9__16 = d_arr_2__31 ;
    assign d_arr_9__15 = d_arr_2__31 ;
    assign d_arr_9__14 = d_arr_2__31 ;
    assign d_arr_9__13 = d_arr_2__31 ;
    assign d_arr_9__12 = d_arr_2__31 ;
    assign d_arr_9__11 = d_arr_2__31 ;
    assign d_arr_9__10 = d_arr_2__31 ;
    assign d_arr_9__9 = d_arr_2__31 ;
    assign d_arr_9__8 = d_arr_2__31 ;
    assign d_arr_9__7 = d_arr_2__31 ;
    assign d_arr_9__6 = d_arr_2__31 ;
    assign d_arr_9__5 = d_arr_2__31 ;
    assign d_arr_9__4 = d_arr_2__31 ;
    assign d_arr_9__3 = d_arr_2__31 ;
    assign d_arr_9__2 = d_arr_2__31 ;
    assign d_arr_9__1 = d_arr_2__31 ;
    assign d_arr_9__0 = d_arr_2__31 ;
    assign d_arr_10__31 = d_arr_2__31 ;
    assign d_arr_10__30 = d_arr_2__31 ;
    assign d_arr_10__29 = d_arr_2__31 ;
    assign d_arr_10__28 = d_arr_2__31 ;
    assign d_arr_10__27 = d_arr_2__31 ;
    assign d_arr_10__26 = d_arr_2__31 ;
    assign d_arr_10__25 = d_arr_2__31 ;
    assign d_arr_10__24 = d_arr_2__31 ;
    assign d_arr_10__23 = d_arr_2__31 ;
    assign d_arr_10__22 = d_arr_2__31 ;
    assign d_arr_10__21 = d_arr_2__31 ;
    assign d_arr_10__20 = d_arr_2__31 ;
    assign d_arr_10__19 = d_arr_2__31 ;
    assign d_arr_10__18 = d_arr_2__31 ;
    assign d_arr_10__17 = d_arr_2__31 ;
    assign d_arr_10__16 = d_arr_2__31 ;
    assign d_arr_10__15 = d_arr_2__31 ;
    assign d_arr_10__14 = d_arr_2__31 ;
    assign d_arr_10__13 = d_arr_2__31 ;
    assign d_arr_10__12 = d_arr_2__31 ;
    assign d_arr_10__11 = d_arr_2__31 ;
    assign d_arr_10__10 = d_arr_2__31 ;
    assign d_arr_10__9 = d_arr_2__31 ;
    assign d_arr_10__8 = d_arr_2__31 ;
    assign d_arr_10__7 = d_arr_2__31 ;
    assign d_arr_10__6 = d_arr_2__31 ;
    assign d_arr_10__5 = d_arr_2__31 ;
    assign d_arr_10__4 = d_arr_2__31 ;
    assign d_arr_10__3 = d_arr_2__31 ;
    assign d_arr_10__2 = d_arr_2__31 ;
    assign d_arr_10__1 = d_arr_2__31 ;
    assign d_arr_10__0 = d_arr_2__31 ;
    assign d_arr_11__31 = d_arr_2__31 ;
    assign d_arr_11__30 = d_arr_2__31 ;
    assign d_arr_11__29 = d_arr_2__31 ;
    assign d_arr_11__28 = d_arr_2__31 ;
    assign d_arr_11__27 = d_arr_2__31 ;
    assign d_arr_11__26 = d_arr_2__31 ;
    assign d_arr_11__25 = d_arr_2__31 ;
    assign d_arr_11__24 = d_arr_2__31 ;
    assign d_arr_11__23 = d_arr_2__31 ;
    assign d_arr_11__22 = d_arr_2__31 ;
    assign d_arr_11__21 = d_arr_2__31 ;
    assign d_arr_11__20 = d_arr_2__31 ;
    assign d_arr_11__19 = d_arr_2__31 ;
    assign d_arr_11__18 = d_arr_2__31 ;
    assign d_arr_11__17 = d_arr_2__31 ;
    assign d_arr_11__16 = d_arr_2__31 ;
    assign d_arr_11__15 = d_arr_2__31 ;
    assign d_arr_11__14 = d_arr_2__31 ;
    assign d_arr_11__13 = d_arr_2__31 ;
    assign d_arr_11__12 = d_arr_2__31 ;
    assign d_arr_11__11 = d_arr_2__31 ;
    assign d_arr_11__10 = d_arr_2__31 ;
    assign d_arr_11__9 = d_arr_2__31 ;
    assign d_arr_11__8 = d_arr_2__31 ;
    assign d_arr_11__7 = d_arr_2__31 ;
    assign d_arr_11__6 = d_arr_2__31 ;
    assign d_arr_11__5 = d_arr_2__31 ;
    assign d_arr_11__4 = d_arr_2__31 ;
    assign d_arr_11__3 = d_arr_2__31 ;
    assign d_arr_11__2 = d_arr_2__31 ;
    assign d_arr_11__1 = d_arr_2__31 ;
    assign d_arr_11__0 = d_arr_2__31 ;
    assign d_arr_12__31 = d_arr_2__31 ;
    assign d_arr_12__30 = d_arr_2__31 ;
    assign d_arr_12__29 = d_arr_2__31 ;
    assign d_arr_12__28 = d_arr_2__31 ;
    assign d_arr_12__27 = d_arr_2__31 ;
    assign d_arr_12__26 = d_arr_2__31 ;
    assign d_arr_12__25 = d_arr_2__31 ;
    assign d_arr_12__24 = d_arr_2__31 ;
    assign d_arr_12__23 = d_arr_2__31 ;
    assign d_arr_12__22 = d_arr_2__31 ;
    assign d_arr_12__21 = d_arr_2__31 ;
    assign d_arr_12__20 = d_arr_2__31 ;
    assign d_arr_12__19 = d_arr_2__31 ;
    assign d_arr_12__18 = d_arr_2__31 ;
    assign d_arr_12__17 = d_arr_2__31 ;
    assign d_arr_12__16 = d_arr_2__31 ;
    assign d_arr_12__15 = d_arr_2__31 ;
    assign d_arr_12__14 = d_arr_2__31 ;
    assign d_arr_12__13 = d_arr_2__31 ;
    assign d_arr_12__12 = d_arr_2__31 ;
    assign d_arr_12__11 = d_arr_2__31 ;
    assign d_arr_12__10 = d_arr_2__31 ;
    assign d_arr_12__9 = d_arr_2__31 ;
    assign d_arr_12__8 = d_arr_2__31 ;
    assign d_arr_12__7 = d_arr_2__31 ;
    assign d_arr_12__6 = d_arr_2__31 ;
    assign d_arr_12__5 = d_arr_2__31 ;
    assign d_arr_12__4 = d_arr_2__31 ;
    assign d_arr_12__3 = d_arr_2__31 ;
    assign d_arr_12__2 = d_arr_2__31 ;
    assign d_arr_12__1 = d_arr_2__31 ;
    assign d_arr_12__0 = d_arr_2__31 ;
    assign d_arr_13__31 = d_arr_2__31 ;
    assign d_arr_13__30 = d_arr_2__31 ;
    assign d_arr_13__29 = d_arr_2__31 ;
    assign d_arr_13__28 = d_arr_2__31 ;
    assign d_arr_13__27 = d_arr_2__31 ;
    assign d_arr_13__26 = d_arr_2__31 ;
    assign d_arr_13__25 = d_arr_2__31 ;
    assign d_arr_13__24 = d_arr_2__31 ;
    assign d_arr_13__23 = d_arr_2__31 ;
    assign d_arr_13__22 = d_arr_2__31 ;
    assign d_arr_13__21 = d_arr_2__31 ;
    assign d_arr_13__20 = d_arr_2__31 ;
    assign d_arr_13__19 = d_arr_2__31 ;
    assign d_arr_13__18 = d_arr_2__31 ;
    assign d_arr_13__17 = d_arr_2__31 ;
    assign d_arr_13__16 = d_arr_2__31 ;
    assign d_arr_13__15 = d_arr_2__31 ;
    assign d_arr_13__14 = d_arr_2__31 ;
    assign d_arr_13__13 = d_arr_2__31 ;
    assign d_arr_13__12 = d_arr_2__31 ;
    assign d_arr_13__11 = d_arr_2__31 ;
    assign d_arr_13__10 = d_arr_2__31 ;
    assign d_arr_13__9 = d_arr_2__31 ;
    assign d_arr_13__8 = d_arr_2__31 ;
    assign d_arr_13__7 = d_arr_2__31 ;
    assign d_arr_13__6 = d_arr_2__31 ;
    assign d_arr_13__5 = d_arr_2__31 ;
    assign d_arr_13__4 = d_arr_2__31 ;
    assign d_arr_13__3 = d_arr_2__31 ;
    assign d_arr_13__2 = d_arr_2__31 ;
    assign d_arr_13__1 = d_arr_2__31 ;
    assign d_arr_13__0 = d_arr_2__31 ;
    assign d_arr_14__31 = d_arr_2__31 ;
    assign d_arr_14__30 = d_arr_2__31 ;
    assign d_arr_14__29 = d_arr_2__31 ;
    assign d_arr_14__28 = d_arr_2__31 ;
    assign d_arr_14__27 = d_arr_2__31 ;
    assign d_arr_14__26 = d_arr_2__31 ;
    assign d_arr_14__25 = d_arr_2__31 ;
    assign d_arr_14__24 = d_arr_2__31 ;
    assign d_arr_14__23 = d_arr_2__31 ;
    assign d_arr_14__22 = d_arr_2__31 ;
    assign d_arr_14__21 = d_arr_2__31 ;
    assign d_arr_14__20 = d_arr_2__31 ;
    assign d_arr_14__19 = d_arr_2__31 ;
    assign d_arr_14__18 = d_arr_2__31 ;
    assign d_arr_14__17 = d_arr_2__31 ;
    assign d_arr_14__16 = d_arr_2__31 ;
    assign d_arr_14__15 = d_arr_2__31 ;
    assign d_arr_14__14 = d_arr_2__31 ;
    assign d_arr_14__13 = d_arr_2__31 ;
    assign d_arr_14__12 = d_arr_2__31 ;
    assign d_arr_14__11 = d_arr_2__31 ;
    assign d_arr_14__10 = d_arr_2__31 ;
    assign d_arr_14__9 = d_arr_2__31 ;
    assign d_arr_14__8 = d_arr_2__31 ;
    assign d_arr_14__7 = d_arr_2__31 ;
    assign d_arr_14__6 = d_arr_2__31 ;
    assign d_arr_14__5 = d_arr_2__31 ;
    assign d_arr_14__4 = d_arr_2__31 ;
    assign d_arr_14__3 = d_arr_2__31 ;
    assign d_arr_14__2 = d_arr_2__31 ;
    assign d_arr_14__1 = d_arr_2__31 ;
    assign d_arr_14__0 = d_arr_2__31 ;
    assign d_arr_15__31 = d_arr_2__31 ;
    assign d_arr_15__30 = d_arr_2__31 ;
    assign d_arr_15__29 = d_arr_2__31 ;
    assign d_arr_15__28 = d_arr_2__31 ;
    assign d_arr_15__27 = d_arr_2__31 ;
    assign d_arr_15__26 = d_arr_2__31 ;
    assign d_arr_15__25 = d_arr_2__31 ;
    assign d_arr_15__24 = d_arr_2__31 ;
    assign d_arr_15__23 = d_arr_2__31 ;
    assign d_arr_15__22 = d_arr_2__31 ;
    assign d_arr_15__21 = d_arr_2__31 ;
    assign d_arr_15__20 = d_arr_2__31 ;
    assign d_arr_15__19 = d_arr_2__31 ;
    assign d_arr_15__18 = d_arr_2__31 ;
    assign d_arr_15__17 = d_arr_2__31 ;
    assign d_arr_15__16 = d_arr_2__31 ;
    assign d_arr_15__15 = d_arr_2__31 ;
    assign d_arr_15__14 = d_arr_2__31 ;
    assign d_arr_15__13 = d_arr_2__31 ;
    assign d_arr_15__12 = d_arr_2__31 ;
    assign d_arr_15__11 = d_arr_2__31 ;
    assign d_arr_15__10 = d_arr_2__31 ;
    assign d_arr_15__9 = d_arr_2__31 ;
    assign d_arr_15__8 = d_arr_2__31 ;
    assign d_arr_15__7 = d_arr_2__31 ;
    assign d_arr_15__6 = d_arr_2__31 ;
    assign d_arr_15__5 = d_arr_2__31 ;
    assign d_arr_15__4 = d_arr_2__31 ;
    assign d_arr_15__3 = d_arr_2__31 ;
    assign d_arr_15__2 = d_arr_2__31 ;
    assign d_arr_15__1 = d_arr_2__31 ;
    assign d_arr_15__0 = d_arr_2__31 ;
    assign d_arr_16__31 = d_arr_2__31 ;
    assign d_arr_16__30 = d_arr_2__31 ;
    assign d_arr_16__29 = d_arr_2__31 ;
    assign d_arr_16__28 = d_arr_2__31 ;
    assign d_arr_16__27 = d_arr_2__31 ;
    assign d_arr_16__26 = d_arr_2__31 ;
    assign d_arr_16__25 = d_arr_2__31 ;
    assign d_arr_16__24 = d_arr_2__31 ;
    assign d_arr_16__23 = d_arr_2__31 ;
    assign d_arr_16__22 = d_arr_2__31 ;
    assign d_arr_16__21 = d_arr_2__31 ;
    assign d_arr_16__20 = d_arr_2__31 ;
    assign d_arr_16__19 = d_arr_2__31 ;
    assign d_arr_16__18 = d_arr_2__31 ;
    assign d_arr_16__17 = d_arr_2__31 ;
    assign d_arr_16__16 = d_arr_2__31 ;
    assign d_arr_16__15 = d_arr_2__31 ;
    assign d_arr_16__14 = d_arr_2__31 ;
    assign d_arr_16__13 = d_arr_2__31 ;
    assign d_arr_16__12 = d_arr_2__31 ;
    assign d_arr_16__11 = d_arr_2__31 ;
    assign d_arr_16__10 = d_arr_2__31 ;
    assign d_arr_16__9 = d_arr_2__31 ;
    assign d_arr_16__8 = d_arr_2__31 ;
    assign d_arr_16__7 = d_arr_2__31 ;
    assign d_arr_16__6 = d_arr_2__31 ;
    assign d_arr_16__5 = d_arr_2__31 ;
    assign d_arr_16__4 = d_arr_2__31 ;
    assign d_arr_16__3 = d_arr_2__31 ;
    assign d_arr_16__2 = d_arr_2__31 ;
    assign d_arr_16__1 = d_arr_2__31 ;
    assign d_arr_16__0 = d_arr_2__31 ;
    assign d_arr_17__31 = d_arr_2__31 ;
    assign d_arr_17__30 = d_arr_2__31 ;
    assign d_arr_17__29 = d_arr_2__31 ;
    assign d_arr_17__28 = d_arr_2__31 ;
    assign d_arr_17__27 = d_arr_2__31 ;
    assign d_arr_17__26 = d_arr_2__31 ;
    assign d_arr_17__25 = d_arr_2__31 ;
    assign d_arr_17__24 = d_arr_2__31 ;
    assign d_arr_17__23 = d_arr_2__31 ;
    assign d_arr_17__22 = d_arr_2__31 ;
    assign d_arr_17__21 = d_arr_2__31 ;
    assign d_arr_17__20 = d_arr_2__31 ;
    assign d_arr_17__19 = d_arr_2__31 ;
    assign d_arr_17__18 = d_arr_2__31 ;
    assign d_arr_17__17 = d_arr_2__31 ;
    assign d_arr_17__16 = d_arr_2__31 ;
    assign d_arr_17__15 = d_arr_2__31 ;
    assign d_arr_17__14 = d_arr_2__31 ;
    assign d_arr_17__13 = d_arr_2__31 ;
    assign d_arr_17__12 = d_arr_2__31 ;
    assign d_arr_17__11 = d_arr_2__31 ;
    assign d_arr_17__10 = d_arr_2__31 ;
    assign d_arr_17__9 = d_arr_2__31 ;
    assign d_arr_17__8 = d_arr_2__31 ;
    assign d_arr_17__7 = d_arr_2__31 ;
    assign d_arr_17__6 = d_arr_2__31 ;
    assign d_arr_17__5 = d_arr_2__31 ;
    assign d_arr_17__4 = d_arr_2__31 ;
    assign d_arr_17__3 = d_arr_2__31 ;
    assign d_arr_17__2 = d_arr_2__31 ;
    assign d_arr_17__1 = d_arr_2__31 ;
    assign d_arr_17__0 = d_arr_2__31 ;
    assign d_arr_18__31 = d_arr_2__31 ;
    assign d_arr_18__30 = d_arr_2__31 ;
    assign d_arr_18__29 = d_arr_2__31 ;
    assign d_arr_18__28 = d_arr_2__31 ;
    assign d_arr_18__27 = d_arr_2__31 ;
    assign d_arr_18__26 = d_arr_2__31 ;
    assign d_arr_18__25 = d_arr_2__31 ;
    assign d_arr_18__24 = d_arr_2__31 ;
    assign d_arr_18__23 = d_arr_2__31 ;
    assign d_arr_18__22 = d_arr_2__31 ;
    assign d_arr_18__21 = d_arr_2__31 ;
    assign d_arr_18__20 = d_arr_2__31 ;
    assign d_arr_18__19 = d_arr_2__31 ;
    assign d_arr_18__18 = d_arr_2__31 ;
    assign d_arr_18__17 = d_arr_2__31 ;
    assign d_arr_18__16 = d_arr_2__31 ;
    assign d_arr_18__15 = d_arr_2__31 ;
    assign d_arr_18__14 = d_arr_2__31 ;
    assign d_arr_18__13 = d_arr_2__31 ;
    assign d_arr_18__12 = d_arr_2__31 ;
    assign d_arr_18__11 = d_arr_2__31 ;
    assign d_arr_18__10 = d_arr_2__31 ;
    assign d_arr_18__9 = d_arr_2__31 ;
    assign d_arr_18__8 = d_arr_2__31 ;
    assign d_arr_18__7 = d_arr_2__31 ;
    assign d_arr_18__6 = d_arr_2__31 ;
    assign d_arr_18__5 = d_arr_2__31 ;
    assign d_arr_18__4 = d_arr_2__31 ;
    assign d_arr_18__3 = d_arr_2__31 ;
    assign d_arr_18__2 = d_arr_2__31 ;
    assign d_arr_18__1 = d_arr_2__31 ;
    assign d_arr_18__0 = d_arr_2__31 ;
    assign d_arr_19__31 = d_arr_2__31 ;
    assign d_arr_19__30 = d_arr_2__31 ;
    assign d_arr_19__29 = d_arr_2__31 ;
    assign d_arr_19__28 = d_arr_2__31 ;
    assign d_arr_19__27 = d_arr_2__31 ;
    assign d_arr_19__26 = d_arr_2__31 ;
    assign d_arr_19__25 = d_arr_2__31 ;
    assign d_arr_19__24 = d_arr_2__31 ;
    assign d_arr_19__23 = d_arr_2__31 ;
    assign d_arr_19__22 = d_arr_2__31 ;
    assign d_arr_19__21 = d_arr_2__31 ;
    assign d_arr_19__20 = d_arr_2__31 ;
    assign d_arr_19__19 = d_arr_2__31 ;
    assign d_arr_19__18 = d_arr_2__31 ;
    assign d_arr_19__17 = d_arr_2__31 ;
    assign d_arr_19__16 = d_arr_2__31 ;
    assign d_arr_19__15 = d_arr_2__31 ;
    assign d_arr_19__14 = d_arr_2__31 ;
    assign d_arr_19__13 = d_arr_2__31 ;
    assign d_arr_19__12 = d_arr_2__31 ;
    assign d_arr_19__11 = d_arr_2__31 ;
    assign d_arr_19__10 = d_arr_2__31 ;
    assign d_arr_19__9 = d_arr_2__31 ;
    assign d_arr_19__8 = d_arr_2__31 ;
    assign d_arr_19__7 = d_arr_2__31 ;
    assign d_arr_19__6 = d_arr_2__31 ;
    assign d_arr_19__5 = d_arr_2__31 ;
    assign d_arr_19__4 = d_arr_2__31 ;
    assign d_arr_19__3 = d_arr_2__31 ;
    assign d_arr_19__2 = d_arr_2__31 ;
    assign d_arr_19__1 = d_arr_2__31 ;
    assign d_arr_19__0 = d_arr_2__31 ;
    assign d_arr_20__31 = d_arr_2__31 ;
    assign d_arr_20__30 = d_arr_2__31 ;
    assign d_arr_20__29 = d_arr_2__31 ;
    assign d_arr_20__28 = d_arr_2__31 ;
    assign d_arr_20__27 = d_arr_2__31 ;
    assign d_arr_20__26 = d_arr_2__31 ;
    assign d_arr_20__25 = d_arr_2__31 ;
    assign d_arr_20__24 = d_arr_2__31 ;
    assign d_arr_20__23 = d_arr_2__31 ;
    assign d_arr_20__22 = d_arr_2__31 ;
    assign d_arr_20__21 = d_arr_2__31 ;
    assign d_arr_20__20 = d_arr_2__31 ;
    assign d_arr_20__19 = d_arr_2__31 ;
    assign d_arr_20__18 = d_arr_2__31 ;
    assign d_arr_20__17 = d_arr_2__31 ;
    assign d_arr_20__16 = d_arr_2__31 ;
    assign d_arr_20__15 = d_arr_2__31 ;
    assign d_arr_20__14 = d_arr_2__31 ;
    assign d_arr_20__13 = d_arr_2__31 ;
    assign d_arr_20__12 = d_arr_2__31 ;
    assign d_arr_20__11 = d_arr_2__31 ;
    assign d_arr_20__10 = d_arr_2__31 ;
    assign d_arr_20__9 = d_arr_2__31 ;
    assign d_arr_20__8 = d_arr_2__31 ;
    assign d_arr_20__7 = d_arr_2__31 ;
    assign d_arr_20__6 = d_arr_2__31 ;
    assign d_arr_20__5 = d_arr_2__31 ;
    assign d_arr_20__4 = d_arr_2__31 ;
    assign d_arr_20__3 = d_arr_2__31 ;
    assign d_arr_20__2 = d_arr_2__31 ;
    assign d_arr_20__1 = d_arr_2__31 ;
    assign d_arr_20__0 = d_arr_2__31 ;
    assign d_arr_21__31 = d_arr_2__31 ;
    assign d_arr_21__30 = d_arr_2__31 ;
    assign d_arr_21__29 = d_arr_2__31 ;
    assign d_arr_21__28 = d_arr_2__31 ;
    assign d_arr_21__27 = d_arr_2__31 ;
    assign d_arr_21__26 = d_arr_2__31 ;
    assign d_arr_21__25 = d_arr_2__31 ;
    assign d_arr_21__24 = d_arr_2__31 ;
    assign d_arr_21__23 = d_arr_2__31 ;
    assign d_arr_21__22 = d_arr_2__31 ;
    assign d_arr_21__21 = d_arr_2__31 ;
    assign d_arr_21__20 = d_arr_2__31 ;
    assign d_arr_21__19 = d_arr_2__31 ;
    assign d_arr_21__18 = d_arr_2__31 ;
    assign d_arr_21__17 = d_arr_2__31 ;
    assign d_arr_21__16 = d_arr_2__31 ;
    assign d_arr_21__15 = d_arr_2__31 ;
    assign d_arr_21__14 = d_arr_2__31 ;
    assign d_arr_21__13 = d_arr_2__31 ;
    assign d_arr_21__12 = d_arr_2__31 ;
    assign d_arr_21__11 = d_arr_2__31 ;
    assign d_arr_21__10 = d_arr_2__31 ;
    assign d_arr_21__9 = d_arr_2__31 ;
    assign d_arr_21__8 = d_arr_2__31 ;
    assign d_arr_21__7 = d_arr_2__31 ;
    assign d_arr_21__6 = d_arr_2__31 ;
    assign d_arr_21__5 = d_arr_2__31 ;
    assign d_arr_21__4 = d_arr_2__31 ;
    assign d_arr_21__3 = d_arr_2__31 ;
    assign d_arr_21__2 = d_arr_2__31 ;
    assign d_arr_21__1 = d_arr_2__31 ;
    assign d_arr_21__0 = d_arr_2__31 ;
    assign d_arr_22__31 = d_arr_2__31 ;
    assign d_arr_22__30 = d_arr_2__31 ;
    assign d_arr_22__29 = d_arr_2__31 ;
    assign d_arr_22__28 = d_arr_2__31 ;
    assign d_arr_22__27 = d_arr_2__31 ;
    assign d_arr_22__26 = d_arr_2__31 ;
    assign d_arr_22__25 = d_arr_2__31 ;
    assign d_arr_22__24 = d_arr_2__31 ;
    assign d_arr_22__23 = d_arr_2__31 ;
    assign d_arr_22__22 = d_arr_2__31 ;
    assign d_arr_22__21 = d_arr_2__31 ;
    assign d_arr_22__20 = d_arr_2__31 ;
    assign d_arr_22__19 = d_arr_2__31 ;
    assign d_arr_22__18 = d_arr_2__31 ;
    assign d_arr_22__17 = d_arr_2__31 ;
    assign d_arr_22__16 = d_arr_2__31 ;
    assign d_arr_22__15 = d_arr_2__31 ;
    assign d_arr_22__14 = d_arr_2__31 ;
    assign d_arr_22__13 = d_arr_2__31 ;
    assign d_arr_22__12 = d_arr_2__31 ;
    assign d_arr_22__11 = d_arr_2__31 ;
    assign d_arr_22__10 = d_arr_2__31 ;
    assign d_arr_22__9 = d_arr_2__31 ;
    assign d_arr_22__8 = d_arr_2__31 ;
    assign d_arr_22__7 = d_arr_2__31 ;
    assign d_arr_22__6 = d_arr_2__31 ;
    assign d_arr_22__5 = d_arr_2__31 ;
    assign d_arr_22__4 = d_arr_2__31 ;
    assign d_arr_22__3 = d_arr_2__31 ;
    assign d_arr_22__2 = d_arr_2__31 ;
    assign d_arr_22__1 = d_arr_2__31 ;
    assign d_arr_22__0 = d_arr_2__31 ;
    assign d_arr_23__31 = d_arr_2__31 ;
    assign d_arr_23__30 = d_arr_2__31 ;
    assign d_arr_23__29 = d_arr_2__31 ;
    assign d_arr_23__28 = d_arr_2__31 ;
    assign d_arr_23__27 = d_arr_2__31 ;
    assign d_arr_23__26 = d_arr_2__31 ;
    assign d_arr_23__25 = d_arr_2__31 ;
    assign d_arr_23__24 = d_arr_2__31 ;
    assign d_arr_23__23 = d_arr_2__31 ;
    assign d_arr_23__22 = d_arr_2__31 ;
    assign d_arr_23__21 = d_arr_2__31 ;
    assign d_arr_23__20 = d_arr_2__31 ;
    assign d_arr_23__19 = d_arr_2__31 ;
    assign d_arr_23__18 = d_arr_2__31 ;
    assign d_arr_23__17 = d_arr_2__31 ;
    assign d_arr_23__16 = d_arr_2__31 ;
    assign d_arr_23__15 = d_arr_2__31 ;
    assign d_arr_23__14 = d_arr_2__31 ;
    assign d_arr_23__13 = d_arr_2__31 ;
    assign d_arr_23__12 = d_arr_2__31 ;
    assign d_arr_23__11 = d_arr_2__31 ;
    assign d_arr_23__10 = d_arr_2__31 ;
    assign d_arr_23__9 = d_arr_2__31 ;
    assign d_arr_23__8 = d_arr_2__31 ;
    assign d_arr_23__7 = d_arr_2__31 ;
    assign d_arr_23__6 = d_arr_2__31 ;
    assign d_arr_23__5 = d_arr_2__31 ;
    assign d_arr_23__4 = d_arr_2__31 ;
    assign d_arr_23__3 = d_arr_2__31 ;
    assign d_arr_23__2 = d_arr_2__31 ;
    assign d_arr_23__1 = d_arr_2__31 ;
    assign d_arr_23__0 = d_arr_2__31 ;
    assign d_arr_24__31 = d_arr_2__31 ;
    assign d_arr_24__30 = d_arr_2__31 ;
    assign d_arr_24__29 = d_arr_2__31 ;
    assign d_arr_24__28 = d_arr_2__31 ;
    assign d_arr_24__27 = d_arr_2__31 ;
    assign d_arr_24__26 = d_arr_2__31 ;
    assign d_arr_24__25 = d_arr_2__31 ;
    assign d_arr_24__24 = d_arr_2__31 ;
    assign d_arr_24__23 = d_arr_2__31 ;
    assign d_arr_24__22 = d_arr_2__31 ;
    assign d_arr_24__21 = d_arr_2__31 ;
    assign d_arr_24__20 = d_arr_2__31 ;
    assign d_arr_24__19 = d_arr_2__31 ;
    assign d_arr_24__18 = d_arr_2__31 ;
    assign d_arr_24__17 = d_arr_2__31 ;
    assign d_arr_24__16 = d_arr_2__31 ;
    assign d_arr_24__15 = d_arr_2__31 ;
    assign d_arr_24__14 = d_arr_2__31 ;
    assign d_arr_24__13 = d_arr_2__31 ;
    assign d_arr_24__12 = d_arr_2__31 ;
    assign d_arr_24__11 = d_arr_2__31 ;
    assign d_arr_24__10 = d_arr_2__31 ;
    assign d_arr_24__9 = d_arr_2__31 ;
    assign d_arr_24__8 = d_arr_2__31 ;
    assign d_arr_24__7 = d_arr_2__31 ;
    assign d_arr_24__6 = d_arr_2__31 ;
    assign d_arr_24__5 = d_arr_2__31 ;
    assign d_arr_24__4 = d_arr_2__31 ;
    assign d_arr_24__3 = d_arr_2__31 ;
    assign d_arr_24__2 = d_arr_2__31 ;
    assign d_arr_24__1 = d_arr_2__31 ;
    assign d_arr_24__0 = d_arr_2__31 ;
    NAdder_32 adder1_gen (.a ({q_arr_9__31,q_arr_9__30,q_arr_9__29,q_arr_9__28,
              nx550,q_arr_9__26,q_arr_9__25,nx555,q_arr_9__23,q_arr_9__22,
              q_arr_9__21,q_arr_9__20,q_arr_9__19,q_arr_9__18,q_arr_9__17,
              q_arr_9__16,q_arr_9__15,q_arr_9__14,q_arr_9__13,q_arr_9__12,
              q_arr_9__11,q_arr_9__10,q_arr_9__9,q_arr_9__8,q_arr_9__7,
              q_arr_9__6,q_arr_9__5,q_arr_9__4,q_arr_9__3,q_arr_9__2,q_arr_9__1,
              q_arr_9__0}), .b ({q_arr_18__31,q_arr_18__30,q_arr_18__29,
              q_arr_18__28,q_arr_18__27,q_arr_18__26,q_arr_18__25,q_arr_18__24,
              q_arr_18__23,q_arr_18__22,q_arr_18__21,q_arr_18__20,q_arr_18__19,
              q_arr_18__18,q_arr_18__17,q_arr_18__16,q_arr_18__15,q_arr_18__14,
              q_arr_18__13,q_arr_18__12,q_arr_18__11,q_arr_18__10,q_arr_18__9,
              q_arr_18__8,q_arr_18__7,q_arr_18__6,q_arr_18__5,q_arr_18__4,
              q_arr_18__3,q_arr_18__2,q_arr_18__1,q_arr_18__0}), .cin (
              d_arr_2__31), .s ({s1_31,s1_30,s1_29,s1_28,s1_27,s1_26,s1_25,s1_24
              ,s1_23,s1_22,s1_21,s1_20,s1_19,s1_18,s1_17,s1_16,s1_15,s1_14,s1_13
              ,s1_12,s1_11,s1_10,s1_9,s1_8,s1_7,s1_6,s1_5,s1_4,s1_3,s1_2,s1_1,
              s1_0}), .cout (\$dummy [0])) ;
    NAdder_32 adder2_gen (.a ({q_arr_0__31,q_arr_0__30,q_arr_0__29,q_arr_0__28,
              q_arr_0__27,q_arr_0__26,q_arr_0__25,q_arr_0__24,q_arr_0__23,
              q_arr_0__22,q_arr_0__21,q_arr_0__20,q_arr_0__19,q_arr_0__18,
              q_arr_0__17,q_arr_0__16,q_arr_0__15,q_arr_0__14,q_arr_0__13,
              q_arr_0__12,q_arr_0__11,q_arr_0__10,q_arr_0__9,q_arr_0__8,
              q_arr_0__7,q_arr_0__6,q_arr_0__5,q_arr_0__4,q_arr_0__3,q_arr_0__2,
              q_arr_0__1,q_arr_0__0}), .b ({s1_31,s1_30,s1_29,s1_28,s1_27,s1_26,
              s1_25,s1_24,s1_23,s1_22,s1_21,s1_20,s1_19,s1_18,s1_17,s1_16,s1_15,
              s1_14,s1_13,s1_12,s1_11,s1_10,s1_9,s1_8,s1_7,s1_6,s1_5,s1_4,s1_3,
              s1_2,s1_1,s1_0}), .cin (d_arr_2__31), .s ({s2_31,s2_30,s2_29,s2_28
              ,s2_27,s2_26,s2_25,s2_24,s2_23,s2_22,s2_21,s2_20,s2_19,s2_18,s2_17
              ,s2_16,s2_15,s2_14,s2_13,s2_12,s2_11,s2_10,s2_9,s2_8,s2_7,s2_6,
              s2_5,s2_4,s2_3,s2_2,s2_1,s2_0}), .cout (\$dummy [1])) ;
    fake_gnd ix41 (.Y (d_arr_2__31)) ;
    inv01 ix17 (.Y (d_arr_1__0), .A (nx153)) ;
    aoi222 ix154 (.Y (nx153), .A0 (q_arr_9__0), .A1 (nx521), .B0 (q_arr_9__5), .B1 (
           nx460), .C0 (q_arr_9__3), .C1 (nx479)) ;
    inv01 ix29 (.Y (d_arr_1__1), .A (nx165)) ;
    aoi222 ix166 (.Y (nx165), .A0 (q_arr_9__1), .A1 (nx521), .B0 (q_arr_9__6), .B1 (
           nx460), .C0 (q_arr_9__4), .C1 (nx479)) ;
    inv01 ix43 (.Y (d_arr_1__2), .A (nx169)) ;
    aoi222 ix170 (.Y (nx169), .A0 (q_arr_9__2), .A1 (nx521), .B0 (q_arr_9__7), .B1 (
           nx460), .C0 (q_arr_9__5), .C1 (nx479)) ;
    inv01 ix53 (.Y (d_arr_1__3), .A (nx173)) ;
    aoi222 ix174 (.Y (nx173), .A0 (q_arr_9__3), .A1 (nx521), .B0 (q_arr_9__8), .B1 (
           nx460), .C0 (q_arr_9__6), .C1 (nx479)) ;
    inv01 ix65 (.Y (d_arr_1__4), .A (nx177)) ;
    aoi222 ix178 (.Y (nx177), .A0 (q_arr_9__4), .A1 (nx521), .B0 (q_arr_9__9), .B1 (
           nx460), .C0 (q_arr_9__7), .C1 (nx479)) ;
    inv01 ix77 (.Y (d_arr_1__5), .A (nx181)) ;
    aoi222 ix182 (.Y (nx181), .A0 (q_arr_9__5), .A1 (nx523), .B0 (q_arr_9__10), 
           .B1 (nx460), .C0 (q_arr_9__8), .C1 (nx479)) ;
    inv01 ix89 (.Y (d_arr_1__6), .A (nx185)) ;
    aoi222 ix186 (.Y (nx185), .A0 (q_arr_9__6), .A1 (nx523), .B0 (q_arr_9__11), 
           .B1 (nx460), .C0 (q_arr_9__9), .C1 (nx479)) ;
    inv01 ix101 (.Y (d_arr_1__7), .A (nx189)) ;
    aoi222 ix190 (.Y (nx189), .A0 (q_arr_9__7), .A1 (nx523), .B0 (q_arr_9__12), 
           .B1 (nx462), .C0 (q_arr_9__10), .C1 (nx481)) ;
    inv01 ix113 (.Y (d_arr_1__8), .A (nx193)) ;
    aoi222 ix194 (.Y (nx193), .A0 (q_arr_9__8), .A1 (nx523), .B0 (q_arr_9__13), 
           .B1 (nx462), .C0 (q_arr_9__11), .C1 (nx481)) ;
    inv01 ix125 (.Y (d_arr_1__9), .A (nx197)) ;
    aoi222 ix198 (.Y (nx197), .A0 (q_arr_9__9), .A1 (nx523), .B0 (q_arr_9__14), 
           .B1 (nx462), .C0 (q_arr_9__12), .C1 (nx481)) ;
    inv01 ix137 (.Y (d_arr_1__10), .A (nx201)) ;
    aoi222 ix202 (.Y (nx201), .A0 (q_arr_9__10), .A1 (nx523), .B0 (q_arr_9__15)
           , .B1 (nx462), .C0 (q_arr_9__13), .C1 (nx481)) ;
    inv01 ix149 (.Y (d_arr_1__11), .A (nx205)) ;
    aoi222 ix206 (.Y (nx205), .A0 (q_arr_9__11), .A1 (nx523), .B0 (q_arr_9__16)
           , .B1 (nx462), .C0 (q_arr_9__14), .C1 (nx481)) ;
    inv01 ix161 (.Y (d_arr_1__12), .A (nx209)) ;
    aoi222 ix210 (.Y (nx209), .A0 (q_arr_9__12), .A1 (nx525), .B0 (q_arr_9__17)
           , .B1 (nx462), .C0 (q_arr_9__15), .C1 (nx481)) ;
    inv01 ix173 (.Y (d_arr_1__13), .A (nx213)) ;
    aoi222 ix214 (.Y (nx213), .A0 (q_arr_9__13), .A1 (nx525), .B0 (q_arr_9__18)
           , .B1 (nx462), .C0 (q_arr_9__16), .C1 (nx481)) ;
    inv01 ix185 (.Y (d_arr_1__14), .A (nx217)) ;
    aoi222 ix218 (.Y (nx217), .A0 (q_arr_9__14), .A1 (nx525), .B0 (q_arr_9__19)
           , .B1 (nx464), .C0 (q_arr_9__17), .C1 (nx483)) ;
    inv01 ix197 (.Y (d_arr_1__15), .A (nx221)) ;
    aoi222 ix222 (.Y (nx221), .A0 (q_arr_9__15), .A1 (nx525), .B0 (q_arr_9__20)
           , .B1 (nx464), .C0 (q_arr_9__18), .C1 (nx483)) ;
    inv01 ix209 (.Y (d_arr_1__16), .A (nx225)) ;
    aoi222 ix226 (.Y (nx225), .A0 (q_arr_9__16), .A1 (nx525), .B0 (q_arr_9__21)
           , .B1 (nx464), .C0 (q_arr_9__19), .C1 (nx483)) ;
    inv01 ix221 (.Y (d_arr_1__17), .A (nx229)) ;
    aoi222 ix230 (.Y (nx229), .A0 (q_arr_9__17), .A1 (nx525), .B0 (q_arr_9__22)
           , .B1 (nx464), .C0 (q_arr_9__20), .C1 (nx483)) ;
    inv01 ix233 (.Y (d_arr_1__18), .A (nx233)) ;
    aoi222 ix234 (.Y (nx233), .A0 (q_arr_9__18), .A1 (nx525), .B0 (q_arr_9__23)
           , .B1 (nx464), .C0 (q_arr_9__21), .C1 (nx483)) ;
    inv01 ix245 (.Y (d_arr_1__19), .A (nx237)) ;
    aoi222 ix238 (.Y (nx237), .A0 (q_arr_9__19), .A1 (nx527), .B0 (nx555), .B1 (
           nx464), .C0 (q_arr_9__22), .C1 (nx483)) ;
    inv01 ix257 (.Y (d_arr_1__20), .A (nx241)) ;
    aoi222 ix242 (.Y (nx241), .A0 (q_arr_9__20), .A1 (nx527), .B0 (q_arr_9__25)
           , .B1 (nx464), .C0 (q_arr_9__23), .C1 (nx483)) ;
    inv01 ix269 (.Y (d_arr_1__21), .A (nx245)) ;
    aoi222 ix246 (.Y (nx245), .A0 (q_arr_9__21), .A1 (nx527), .B0 (q_arr_9__26)
           , .B1 (nx466), .C0 (nx555), .C1 (nx485)) ;
    inv01 ix281 (.Y (d_arr_1__22), .A (nx249)) ;
    aoi222 ix250 (.Y (nx249), .A0 (q_arr_9__22), .A1 (nx527), .B0 (nx550), .B1 (
           nx466), .C0 (q_arr_9__25), .C1 (nx485)) ;
    inv01 ix293 (.Y (d_arr_1__23), .A (nx253)) ;
    aoi222 ix254 (.Y (nx253), .A0 (q_arr_9__23), .A1 (nx527), .B0 (q_arr_9__28)
           , .B1 (nx466), .C0 (q_arr_9__26), .C1 (nx485)) ;
    inv01 ix305 (.Y (d_arr_1__24), .A (nx257)) ;
    aoi222 ix258 (.Y (nx257), .A0 (nx555), .A1 (nx527), .B0 (q_arr_9__29), .B1 (
           nx466), .C0 (nx550), .C1 (nx485)) ;
    inv01 ix317 (.Y (d_arr_1__25), .A (nx261)) ;
    aoi222 ix262 (.Y (nx261), .A0 (q_arr_9__25), .A1 (nx527), .B0 (q_arr_9__30)
           , .B1 (nx466), .C0 (q_arr_9__28), .C1 (nx485)) ;
    inv01 ix329 (.Y (d_arr_1__26), .A (nx265)) ;
    aoi222 ix266 (.Y (nx265), .A0 (q_arr_9__26), .A1 (nx529), .B0 (q_arr_9__31)
           , .B1 (nx466), .C0 (q_arr_9__29), .C1 (nx485)) ;
    ao22 ix337 (.Y (d_arr_1__27), .A0 (nx553), .A1 (nx529), .B0 (q_arr_9__30), .B1 (
         nx485)) ;
    ao22 ix345 (.Y (d_arr_1__28), .A0 (q_arr_9__28), .A1 (nx529), .B0 (
         q_arr_9__31), .B1 (nx487)) ;
    nor02ii ix757 (.Y (d_arr_1__29), .A0 (nx540), .A1 (q_arr_9__29)) ;
    nor02ii ix761 (.Y (d_arr_1__30), .A0 (nx540), .A1 (q_arr_9__30)) ;
    nor02ii ix765 (.Y (d_arr_1__31), .A0 (nx540), .A1 (q_arr_9__31)) ;
    nand02 ix369 (.Y (d_arr_0__0), .A0 (nx277), .A1 (nx279)) ;
    aoi22 ix278 (.Y (nx277), .A0 (s2_5), .A1 (nx466), .B0 (q_arr_0__3), .B1 (
          nx487)) ;
    aoi22 ix280 (.Y (nx279), .A0 (s2_0), .A1 (nx499), .B0 (q_arr_0__0), .B1 (
          nx511)) ;
    nor02_2x ix351 (.Y (nx350), .A0 (filter_size), .A1 (nx540)) ;
    nand02 ix383 (.Y (d_arr_0__1), .A0 (nx285), .A1 (nx287)) ;
    aoi22 ix286 (.Y (nx285), .A0 (s2_6), .A1 (nx469), .B0 (q_arr_0__4), .B1 (
          nx487)) ;
    aoi22 ix288 (.Y (nx287), .A0 (s2_1), .A1 (nx499), .B0 (q_arr_0__1), .B1 (
          nx511)) ;
    nand02 ix397 (.Y (d_arr_0__2), .A0 (nx291), .A1 (nx293)) ;
    aoi22 ix292 (.Y (nx291), .A0 (s2_7), .A1 (nx469), .B0 (q_arr_0__5), .B1 (
          nx487)) ;
    aoi22 ix294 (.Y (nx293), .A0 (s2_2), .A1 (nx499), .B0 (q_arr_0__2), .B1 (
          nx511)) ;
    nand02 ix411 (.Y (d_arr_0__3), .A0 (nx297), .A1 (nx299)) ;
    aoi22 ix298 (.Y (nx297), .A0 (s2_8), .A1 (nx469), .B0 (q_arr_0__6), .B1 (
          nx487)) ;
    aoi22 ix300 (.Y (nx299), .A0 (s2_3), .A1 (nx499), .B0 (q_arr_0__3), .B1 (
          nx511)) ;
    nand02 ix425 (.Y (d_arr_0__4), .A0 (nx303), .A1 (nx305)) ;
    aoi22 ix304 (.Y (nx303), .A0 (s2_9), .A1 (nx469), .B0 (q_arr_0__7), .B1 (
          nx487)) ;
    aoi22 ix306 (.Y (nx305), .A0 (s2_4), .A1 (nx499), .B0 (q_arr_0__4), .B1 (
          nx511)) ;
    nand02 ix439 (.Y (d_arr_0__5), .A0 (nx309), .A1 (nx311)) ;
    aoi22 ix310 (.Y (nx309), .A0 (s2_10), .A1 (nx469), .B0 (q_arr_0__8), .B1 (
          nx487)) ;
    aoi22 ix312 (.Y (nx311), .A0 (s2_5), .A1 (nx499), .B0 (q_arr_0__5), .B1 (
          nx511)) ;
    nand02 ix453 (.Y (d_arr_0__6), .A0 (nx315), .A1 (nx317)) ;
    aoi22 ix316 (.Y (nx315), .A0 (s2_11), .A1 (nx469), .B0 (q_arr_0__9), .B1 (
          nx489)) ;
    aoi22 ix318 (.Y (nx317), .A0 (s2_6), .A1 (nx499), .B0 (q_arr_0__6), .B1 (
          nx511)) ;
    nand02 ix467 (.Y (d_arr_0__7), .A0 (nx321), .A1 (nx323)) ;
    aoi22 ix322 (.Y (nx321), .A0 (s2_12), .A1 (nx469), .B0 (q_arr_0__10), .B1 (
          nx489)) ;
    aoi22 ix324 (.Y (nx323), .A0 (s2_7), .A1 (nx501), .B0 (q_arr_0__7), .B1 (
          nx513)) ;
    nand02 ix481 (.Y (d_arr_0__8), .A0 (nx327), .A1 (nx329)) ;
    aoi22 ix328 (.Y (nx327), .A0 (s2_13), .A1 (nx471), .B0 (q_arr_0__11), .B1 (
          nx489)) ;
    aoi22 ix330 (.Y (nx329), .A0 (s2_8), .A1 (nx501), .B0 (q_arr_0__8), .B1 (
          nx513)) ;
    nand02 ix495 (.Y (d_arr_0__9), .A0 (nx333), .A1 (nx335)) ;
    aoi22 ix334 (.Y (nx333), .A0 (s2_14), .A1 (nx471), .B0 (q_arr_0__12), .B1 (
          nx489)) ;
    aoi22 ix336 (.Y (nx335), .A0 (s2_9), .A1 (nx501), .B0 (q_arr_0__9), .B1 (
          nx513)) ;
    nand02 ix509 (.Y (d_arr_0__10), .A0 (nx339), .A1 (nx341)) ;
    aoi22 ix340 (.Y (nx339), .A0 (s2_15), .A1 (nx471), .B0 (q_arr_0__13), .B1 (
          nx489)) ;
    aoi22 ix342 (.Y (nx341), .A0 (s2_10), .A1 (nx501), .B0 (q_arr_0__10), .B1 (
          nx513)) ;
    nand02 ix523 (.Y (d_arr_0__11), .A0 (nx345), .A1 (nx347)) ;
    aoi22 ix346 (.Y (nx345), .A0 (s2_16), .A1 (nx471), .B0 (q_arr_0__14), .B1 (
          nx489)) ;
    aoi22 ix348 (.Y (nx347), .A0 (s2_11), .A1 (nx501), .B0 (q_arr_0__11), .B1 (
          nx513)) ;
    nand02 ix537 (.Y (d_arr_0__12), .A0 (nx351), .A1 (nx353)) ;
    aoi22 ix352 (.Y (nx351), .A0 (s2_17), .A1 (nx471), .B0 (q_arr_0__15), .B1 (
          nx489)) ;
    aoi22 ix354 (.Y (nx353), .A0 (s2_12), .A1 (nx501), .B0 (q_arr_0__12), .B1 (
          nx513)) ;
    nand02 ix551 (.Y (d_arr_0__13), .A0 (nx357), .A1 (nx359)) ;
    aoi22 ix358 (.Y (nx357), .A0 (s2_18), .A1 (nx471), .B0 (q_arr_0__16), .B1 (
          nx491)) ;
    aoi22 ix360 (.Y (nx359), .A0 (s2_13), .A1 (nx501), .B0 (q_arr_0__13), .B1 (
          nx513)) ;
    nand02 ix565 (.Y (d_arr_0__14), .A0 (nx363), .A1 (nx365)) ;
    aoi22 ix364 (.Y (nx363), .A0 (s2_19), .A1 (nx471), .B0 (q_arr_0__17), .B1 (
          nx491)) ;
    aoi22 ix366 (.Y (nx365), .A0 (s2_14), .A1 (nx503), .B0 (q_arr_0__14), .B1 (
          nx515)) ;
    nand02 ix579 (.Y (d_arr_0__15), .A0 (nx369), .A1 (nx371)) ;
    aoi22 ix370 (.Y (nx369), .A0 (s2_20), .A1 (nx473), .B0 (q_arr_0__18), .B1 (
          nx491)) ;
    aoi22 ix372 (.Y (nx371), .A0 (s2_15), .A1 (nx503), .B0 (q_arr_0__15), .B1 (
          nx515)) ;
    nand02 ix593 (.Y (d_arr_0__16), .A0 (nx375), .A1 (nx377)) ;
    aoi22 ix376 (.Y (nx375), .A0 (s2_21), .A1 (nx473), .B0 (q_arr_0__19), .B1 (
          nx491)) ;
    aoi22 ix378 (.Y (nx377), .A0 (s2_16), .A1 (nx503), .B0 (q_arr_0__16), .B1 (
          nx515)) ;
    nand02 ix607 (.Y (d_arr_0__17), .A0 (nx381), .A1 (nx383)) ;
    aoi22 ix382 (.Y (nx381), .A0 (s2_22), .A1 (nx473), .B0 (q_arr_0__20), .B1 (
          nx491)) ;
    aoi22 ix384 (.Y (nx383), .A0 (s2_17), .A1 (nx503), .B0 (q_arr_0__17), .B1 (
          nx515)) ;
    nand02 ix621 (.Y (d_arr_0__18), .A0 (nx387), .A1 (nx389)) ;
    aoi22 ix388 (.Y (nx387), .A0 (s2_23), .A1 (nx473), .B0 (q_arr_0__21), .B1 (
          nx491)) ;
    aoi22 ix390 (.Y (nx389), .A0 (s2_18), .A1 (nx503), .B0 (q_arr_0__18), .B1 (
          nx515)) ;
    nand02 ix635 (.Y (d_arr_0__19), .A0 (nx393), .A1 (nx395)) ;
    aoi22 ix394 (.Y (nx393), .A0 (s2_24), .A1 (nx473), .B0 (q_arr_0__22), .B1 (
          nx491)) ;
    aoi22 ix396 (.Y (nx395), .A0 (s2_19), .A1 (nx503), .B0 (q_arr_0__19), .B1 (
          nx515)) ;
    nand02 ix649 (.Y (d_arr_0__20), .A0 (nx399), .A1 (nx401)) ;
    aoi22 ix400 (.Y (nx399), .A0 (s2_25), .A1 (nx473), .B0 (q_arr_0__23), .B1 (
          nx493)) ;
    aoi22 ix402 (.Y (nx401), .A0 (s2_20), .A1 (nx503), .B0 (q_arr_0__20), .B1 (
          nx515)) ;
    nand02 ix663 (.Y (d_arr_0__21), .A0 (nx405), .A1 (nx407)) ;
    aoi22 ix406 (.Y (nx405), .A0 (s2_26), .A1 (nx473), .B0 (q_arr_0__24), .B1 (
          nx493)) ;
    aoi22 ix408 (.Y (nx407), .A0 (s2_21), .A1 (nx505), .B0 (q_arr_0__21), .B1 (
          nx517)) ;
    nand02 ix677 (.Y (d_arr_0__22), .A0 (nx411), .A1 (nx413)) ;
    aoi22 ix412 (.Y (nx411), .A0 (s2_27), .A1 (nx475), .B0 (q_arr_0__25), .B1 (
          nx493)) ;
    aoi22 ix414 (.Y (nx413), .A0 (s2_22), .A1 (nx505), .B0 (q_arr_0__22), .B1 (
          nx517)) ;
    nand02 ix691 (.Y (d_arr_0__23), .A0 (nx417), .A1 (nx419)) ;
    aoi22 ix418 (.Y (nx417), .A0 (s2_28), .A1 (nx475), .B0 (q_arr_0__26), .B1 (
          nx493)) ;
    aoi22 ix420 (.Y (nx419), .A0 (s2_23), .A1 (nx505), .B0 (q_arr_0__23), .B1 (
          nx517)) ;
    nand02 ix705 (.Y (d_arr_0__24), .A0 (nx423), .A1 (nx425)) ;
    aoi22 ix424 (.Y (nx423), .A0 (s2_29), .A1 (nx475), .B0 (q_arr_0__27), .B1 (
          nx493)) ;
    aoi22 ix426 (.Y (nx425), .A0 (s2_24), .A1 (nx505), .B0 (q_arr_0__24), .B1 (
          nx517)) ;
    nand02 ix719 (.Y (d_arr_0__25), .A0 (nx429), .A1 (nx431)) ;
    aoi22 ix430 (.Y (nx429), .A0 (s2_30), .A1 (nx475), .B0 (q_arr_0__28), .B1 (
          nx493)) ;
    aoi22 ix432 (.Y (nx431), .A0 (s2_25), .A1 (nx505), .B0 (q_arr_0__25), .B1 (
          nx517)) ;
    nand02 ix733 (.Y (d_arr_0__26), .A0 (nx435), .A1 (nx437)) ;
    aoi22 ix436 (.Y (nx435), .A0 (s2_31), .A1 (nx475), .B0 (q_arr_0__29), .B1 (
          nx493)) ;
    aoi22 ix438 (.Y (nx437), .A0 (s2_26), .A1 (nx505), .B0 (q_arr_0__26), .B1 (
          nx517)) ;
    inv01 ix743 (.Y (d_arr_0__27), .A (nx441)) ;
    aoi222 ix442 (.Y (nx441), .A0 (s2_27), .A1 (nx505), .B0 (q_arr_0__27), .B1 (
           nx517), .C0 (q_arr_0__30), .C1 (nx495)) ;
    inv01 ix753 (.Y (d_arr_0__28), .A (nx445)) ;
    aoi222 ix446 (.Y (nx445), .A0 (s2_28), .A1 (nx507), .B0 (q_arr_0__28), .B1 (
           nx519), .C0 (q_arr_0__31), .C1 (nx495)) ;
    ao32 ix771 (.Y (d_arr_0__29), .A0 (q_arr_0__29), .A1 (filter_size), .A2 (
         nx529), .B0 (s2_29), .B1 (nx507)) ;
    ao32 ix777 (.Y (d_arr_0__30), .A0 (q_arr_0__30), .A1 (filter_size), .A2 (
         nx529), .B0 (s2_30), .B1 (nx507)) ;
    ao32 ix783 (.Y (d_arr_0__31), .A0 (q_arr_0__31), .A1 (filter_size), .A2 (
         nx529), .B0 (s2_31), .B1 (nx507)) ;
    inv01 ix457 (.Y (nx458), .A (nx6)) ;
    inv02 ix459 (.Y (nx460), .A (nx531)) ;
    inv02 ix461 (.Y (nx462), .A (nx531)) ;
    inv02 ix463 (.Y (nx464), .A (nx531)) ;
    inv02 ix465 (.Y (nx466), .A (nx531)) ;
    inv02 ix468 (.Y (nx469), .A (nx531)) ;
    inv02 ix470 (.Y (nx471), .A (nx458)) ;
    inv02 ix472 (.Y (nx473), .A (nx458)) ;
    inv02 ix474 (.Y (nx475), .A (nx458)) ;
    inv01 ix476 (.Y (nx477), .A (nx10)) ;
    inv02 ix478 (.Y (nx479), .A (nx533)) ;
    inv02 ix480 (.Y (nx481), .A (nx533)) ;
    inv02 ix482 (.Y (nx483), .A (nx533)) ;
    inv02 ix484 (.Y (nx485), .A (nx533)) ;
    inv02 ix486 (.Y (nx487), .A (nx533)) ;
    inv02 ix488 (.Y (nx489), .A (nx477)) ;
    inv02 ix490 (.Y (nx491), .A (nx477)) ;
    inv02 ix492 (.Y (nx493), .A (nx477)) ;
    inv02 ix494 (.Y (nx495), .A (nx477)) ;
    inv01 ix496 (.Y (nx497), .A (nx350)) ;
    inv02 ix498 (.Y (nx499), .A (nx497)) ;
    inv02 ix500 (.Y (nx501), .A (nx497)) ;
    inv02 ix502 (.Y (nx503), .A (nx497)) ;
    inv02 ix504 (.Y (nx505), .A (nx497)) ;
    inv02 ix506 (.Y (nx507), .A (nx497)) ;
    inv02 ix510 (.Y (nx511), .A (nx509)) ;
    inv02 ix512 (.Y (nx513), .A (nx509)) ;
    inv02 ix514 (.Y (nx515), .A (nx509)) ;
    inv02 ix516 (.Y (nx517), .A (nx509)) ;
    inv02 ix518 (.Y (nx519), .A (nx509)) ;
    inv02 ix520 (.Y (nx521), .A (operation)) ;
    inv02 ix522 (.Y (nx523), .A (nx540)) ;
    inv02 ix524 (.Y (nx525), .A (nx540)) ;
    inv02 ix526 (.Y (nx527), .A (nx540)) ;
    inv02 ix528 (.Y (nx529), .A (nx542)) ;
    inv01 ix530 (.Y (nx531), .A (nx6)) ;
    inv01 ix532 (.Y (nx533), .A (nx10)) ;
    nor02ii ix7 (.Y (nx6), .A0 (filter_size), .A1 (nx542)) ;
    and02 ix11 (.Y (nx10), .A0 (filter_size), .A1 (nx542)) ;
    nand02 ix357 (.Y (nx509), .A0 (filter_size), .A1 (nx521)) ;
    inv02 ix539 (.Y (nx540), .A (nx521)) ;
    inv02 ix541 (.Y (nx542), .A (nx521)) ;
    buf02 ix549 (.Y (nx550), .A (q_arr_9__27)) ;
    buf02 ix552 (.Y (nx553), .A (q_arr_9__27)) ;
    buf02 ix554 (.Y (nx555), .A (q_arr_9__24)) ;
endmodule


module NAdder_32 ( a, b, cin, s, cout ) ;

    input [31:0]a ;
    input [31:0]b ;
    input cin ;
    output [31:0]s ;
    output cout ;

    wire nx2, nx16, nx18, nx32, nx34, nx48, nx50, nx64, nx66, nx80, nx82, nx96, 
         nx98, nx112, nx114, nx128, nx130, nx144, nx146, nx160, nx162, nx176, 
         nx178, nx210, nx224, nx226, nx240, nx153, nx155, nx159, nx163, nx169, 
         nx171, nx175, nx179, nx185, nx187, nx191, nx195, nx201, nx203, nx207, 
         nx211, nx217, nx219, nx223, nx227, nx233, nx235, nx239, nx243, nx249, 
         nx251, nx255, nx259, nx265, nx267, nx271, nx275, nx281, nx283, nx287, 
         nx291, nx297, nx299, nx303, nx307, nx313, nx315, nx318, nx321, nx325, 
         nx327, nx339, nx345, nx349, nx354, nx357, nx361, nx363, nx366, nx369, 
         nx373, nx375, nx385, nx386, nx387, nx388, nx208, nx389, nx390, nx391, 
         nx392, nx393, nx394, nx395, nx351, nx342, nx192, nx330, nx396, nx333;



    fake_gnd ix73 (.Y (cout)) ;
    xor2 ix311 (.Y (s[0]), .A0 (b[0]), .A1 (a[0])) ;
    xor2 ix305 (.Y (s[1]), .A0 (nx153), .A1 (nx155)) ;
    nand02 ix154 (.Y (nx153), .A0 (b[0]), .A1 (a[0])) ;
    xnor2 ix156 (.Y (nx155), .A0 (a[1]), .A1 (b[1])) ;
    xor2 ix303 (.Y (s[2]), .A0 (nx159), .A1 (nx163)) ;
    aoi32 ix160 (.Y (nx159), .A0 (b[0]), .A1 (a[0]), .A2 (nx2), .B0 (b[1]), .B1 (
          a[1])) ;
    xnor2 ix164 (.Y (nx163), .A0 (a[2]), .A1 (b[2])) ;
    xnor2 ix301 (.Y (s[3]), .A0 (nx16), .A1 (nx171)) ;
    oai21 ix17 (.Y (nx16), .A0 (nx159), .A1 (nx163), .B0 (nx169)) ;
    nand02 ix170 (.Y (nx169), .A0 (b[2]), .A1 (a[2])) ;
    xnor2 ix172 (.Y (nx171), .A0 (a[3]), .A1 (b[3])) ;
    xor2 ix299 (.Y (s[4]), .A0 (nx175), .A1 (nx179)) ;
    aoi22 ix176 (.Y (nx175), .A0 (b[3]), .A1 (a[3]), .B0 (nx16), .B1 (nx18)) ;
    xnor2 ix180 (.Y (nx179), .A0 (a[4]), .A1 (b[4])) ;
    xnor2 ix297 (.Y (s[5]), .A0 (nx32), .A1 (nx187)) ;
    oai21 ix33 (.Y (nx32), .A0 (nx175), .A1 (nx179), .B0 (nx185)) ;
    nand02 ix186 (.Y (nx185), .A0 (b[4]), .A1 (a[4])) ;
    xnor2 ix188 (.Y (nx187), .A0 (a[5]), .A1 (b[5])) ;
    xor2 ix295 (.Y (s[6]), .A0 (nx191), .A1 (nx195)) ;
    aoi22 ix192 (.Y (nx191), .A0 (b[5]), .A1 (a[5]), .B0 (nx32), .B1 (nx34)) ;
    xnor2 ix196 (.Y (nx195), .A0 (a[6]), .A1 (b[6])) ;
    xnor2 ix293 (.Y (s[7]), .A0 (nx48), .A1 (nx203)) ;
    oai21 ix49 (.Y (nx48), .A0 (nx191), .A1 (nx195), .B0 (nx201)) ;
    nand02 ix202 (.Y (nx201), .A0 (b[6]), .A1 (a[6])) ;
    xnor2 ix204 (.Y (nx203), .A0 (a[7]), .A1 (b[7])) ;
    xor2 ix291 (.Y (s[8]), .A0 (nx207), .A1 (nx211)) ;
    aoi22 ix208 (.Y (nx207), .A0 (b[7]), .A1 (a[7]), .B0 (nx48), .B1 (nx50)) ;
    xnor2 ix212 (.Y (nx211), .A0 (a[8]), .A1 (b[8])) ;
    xnor2 ix289 (.Y (s[9]), .A0 (nx64), .A1 (nx219)) ;
    oai21 ix65 (.Y (nx64), .A0 (nx207), .A1 (nx211), .B0 (nx217)) ;
    nand02 ix218 (.Y (nx217), .A0 (b[8]), .A1 (a[8])) ;
    xnor2 ix220 (.Y (nx219), .A0 (a[9]), .A1 (b[9])) ;
    xor2 ix287 (.Y (s[10]), .A0 (nx223), .A1 (nx227)) ;
    aoi22 ix224 (.Y (nx223), .A0 (b[9]), .A1 (a[9]), .B0 (nx64), .B1 (nx66)) ;
    xnor2 ix228 (.Y (nx227), .A0 (a[10]), .A1 (b[10])) ;
    xnor2 ix285 (.Y (s[11]), .A0 (nx80), .A1 (nx235)) ;
    oai21 ix81 (.Y (nx80), .A0 (nx223), .A1 (nx227), .B0 (nx233)) ;
    nand02 ix234 (.Y (nx233), .A0 (b[10]), .A1 (a[10])) ;
    xnor2 ix236 (.Y (nx235), .A0 (a[11]), .A1 (b[11])) ;
    xor2 ix283 (.Y (s[12]), .A0 (nx239), .A1 (nx243)) ;
    aoi22 ix240 (.Y (nx239), .A0 (b[11]), .A1 (a[11]), .B0 (nx80), .B1 (nx82)) ;
    xnor2 ix244 (.Y (nx243), .A0 (a[12]), .A1 (b[12])) ;
    xnor2 ix281 (.Y (s[13]), .A0 (nx96), .A1 (nx251)) ;
    oai21 ix97 (.Y (nx96), .A0 (nx239), .A1 (nx243), .B0 (nx249)) ;
    nand02 ix250 (.Y (nx249), .A0 (b[12]), .A1 (a[12])) ;
    xnor2 ix252 (.Y (nx251), .A0 (a[13]), .A1 (b[13])) ;
    xor2 ix279 (.Y (s[14]), .A0 (nx255), .A1 (nx259)) ;
    aoi22 ix256 (.Y (nx255), .A0 (b[13]), .A1 (a[13]), .B0 (nx96), .B1 (nx98)) ;
    xnor2 ix260 (.Y (nx259), .A0 (a[14]), .A1 (b[14])) ;
    xnor2 ix277 (.Y (s[15]), .A0 (nx112), .A1 (nx267)) ;
    oai21 ix113 (.Y (nx112), .A0 (nx255), .A1 (nx259), .B0 (nx265)) ;
    nand02 ix266 (.Y (nx265), .A0 (b[14]), .A1 (a[14])) ;
    xnor2 ix268 (.Y (nx267), .A0 (a[15]), .A1 (b[15])) ;
    xor2 ix275 (.Y (s[16]), .A0 (nx271), .A1 (nx275)) ;
    aoi22 ix272 (.Y (nx271), .A0 (b[15]), .A1 (a[15]), .B0 (nx112), .B1 (nx114)
          ) ;
    xnor2 ix276 (.Y (nx275), .A0 (a[16]), .A1 (b[16])) ;
    xnor2 ix273 (.Y (s[17]), .A0 (nx128), .A1 (nx283)) ;
    oai21 ix129 (.Y (nx128), .A0 (nx271), .A1 (nx275), .B0 (nx281)) ;
    nand02 ix282 (.Y (nx281), .A0 (b[16]), .A1 (a[16])) ;
    xnor2 ix284 (.Y (nx283), .A0 (a[17]), .A1 (b[17])) ;
    xor2 ix271 (.Y (s[18]), .A0 (nx287), .A1 (nx291)) ;
    aoi22 ix288 (.Y (nx287), .A0 (b[17]), .A1 (a[17]), .B0 (nx128), .B1 (nx130)
          ) ;
    xnor2 ix292 (.Y (nx291), .A0 (a[18]), .A1 (b[18])) ;
    xnor2 ix269 (.Y (s[19]), .A0 (nx144), .A1 (nx299)) ;
    oai21 ix145 (.Y (nx144), .A0 (nx287), .A1 (nx291), .B0 (nx297)) ;
    nand02 ix298 (.Y (nx297), .A0 (b[18]), .A1 (a[18])) ;
    xnor2 ix300 (.Y (nx299), .A0 (a[19]), .A1 (b[19])) ;
    xor2 ix267 (.Y (s[20]), .A0 (nx303), .A1 (nx307)) ;
    aoi22 ix304 (.Y (nx303), .A0 (b[19]), .A1 (a[19]), .B0 (nx144), .B1 (nx146)
          ) ;
    xnor2 ix308 (.Y (nx307), .A0 (a[20]), .A1 (b[20])) ;
    xnor2 ix265 (.Y (s[21]), .A0 (nx160), .A1 (nx315)) ;
    oai21 ix161 (.Y (nx160), .A0 (nx303), .A1 (nx307), .B0 (nx313)) ;
    nand02 ix314 (.Y (nx313), .A0 (b[20]), .A1 (a[20])) ;
    xnor2 ix316 (.Y (nx315), .A0 (a[21]), .A1 (b[21])) ;
    xor2 ix263 (.Y (s[22]), .A0 (nx318), .A1 (nx321)) ;
    aoi22 ix319 (.Y (nx318), .A0 (b[21]), .A1 (a[21]), .B0 (nx160), .B1 (nx162)
          ) ;
    xnor2 ix322 (.Y (nx321), .A0 (a[22]), .A1 (b[22])) ;
    xnor2 ix261 (.Y (s[23]), .A0 (nx176), .A1 (nx327)) ;
    oai21 ix177 (.Y (nx176), .A0 (nx318), .A1 (nx321), .B0 (nx325)) ;
    nand02 ix326 (.Y (nx325), .A0 (b[22]), .A1 (a[22])) ;
    xnor2 ix328 (.Y (nx327), .A0 (a[23]), .A1 (b[23])) ;
    xor2 ix259 (.Y (s[24]), .A0 (nx330), .A1 (nx333)) ;
    xnor2 ix257 (.Y (s[25]), .A0 (nx192), .A1 (nx339)) ;
    xnor2 ix340 (.Y (nx339), .A0 (a[25]), .A1 (b[25])) ;
    xor2 ix255 (.Y (s[26]), .A0 (nx342), .A1 (nx345)) ;
    xnor2 ix346 (.Y (nx345), .A0 (a[26]), .A1 (b[26])) ;
    nand02 ix350 (.Y (nx349), .A0 (b[26]), .A1 (a[26])) ;
    xor2 ix251 (.Y (s[28]), .A0 (nx354), .A1 (nx357)) ;
    aoi22 ix355 (.Y (nx354), .A0 (b[27]), .A1 (a[27]), .B0 (nx395), .B1 (nx210)
          ) ;
    xnor2 ix358 (.Y (nx357), .A0 (a[28]), .A1 (b[28])) ;
    xnor2 ix249 (.Y (s[29]), .A0 (nx224), .A1 (nx363)) ;
    oai21 ix225 (.Y (nx224), .A0 (nx354), .A1 (nx357), .B0 (nx361)) ;
    nand02 ix362 (.Y (nx361), .A0 (b[28]), .A1 (a[28])) ;
    xnor2 ix364 (.Y (nx363), .A0 (a[29]), .A1 (b[29])) ;
    xor2 ix247 (.Y (s[30]), .A0 (nx366), .A1 (nx369)) ;
    aoi22 ix367 (.Y (nx366), .A0 (b[29]), .A1 (a[29]), .B0 (nx224), .B1 (nx226)
          ) ;
    xnor2 ix370 (.Y (nx369), .A0 (a[30]), .A1 (b[30])) ;
    xnor2 ix245 (.Y (s[31]), .A0 (nx240), .A1 (nx375)) ;
    oai21 ix241 (.Y (nx240), .A0 (nx366), .A1 (nx369), .B0 (nx373)) ;
    nand02 ix374 (.Y (nx373), .A0 (b[30]), .A1 (a[30])) ;
    xnor2 ix376 (.Y (nx375), .A0 (a[31]), .A1 (b[31])) ;
    inv01 ix227 (.Y (nx226), .A (nx363)) ;
    inv01 ix211 (.Y (nx210), .A (nx351)) ;
    inv01 ix179 (.Y (nx178), .A (nx327)) ;
    inv01 ix163 (.Y (nx162), .A (nx315)) ;
    inv01 ix147 (.Y (nx146), .A (nx299)) ;
    inv01 ix131 (.Y (nx130), .A (nx283)) ;
    inv01 ix115 (.Y (nx114), .A (nx267)) ;
    inv01 ix99 (.Y (nx98), .A (nx251)) ;
    inv01 ix83 (.Y (nx82), .A (nx235)) ;
    inv01 ix67 (.Y (nx66), .A (nx219)) ;
    inv01 ix51 (.Y (nx50), .A (nx203)) ;
    inv01 ix35 (.Y (nx34), .A (nx187)) ;
    inv01 ix19 (.Y (nx18), .A (nx171)) ;
    inv01 ix3 (.Y (nx2), .A (nx155)) ;
    or02 ix397 (.Y (nx385), .A0 (a[24]), .A1 (b[24])) ;
    and02 ix398 (.Y (nx386), .A0 (b[23]), .A1 (a[23])) ;
    aoi322 ix399 (.Y (nx387), .A0 (nx176), .A1 (nx178), .A2 (nx385), .B0 (nx385)
           , .B1 (nx386), .C0 (a[24]), .C1 (b[24])) ;
    nand02_2x ix400 (.Y (nx388), .A0 (b[25]), .A1 (a[25])) ;
    oai321 reg_nx208 (.Y (nx208), .A0 (nx387), .A1 (nx345), .A2 (nx339), .B0 (
           nx345), .B1 (nx388), .C0 (nx349)) ;
    inv02 ix401 (.Y (nx389), .A (nx208)) ;
    inv02 ix402 (.Y (nx390), .A (a[27])) ;
    inv02 ix403 (.Y (nx391), .A (b[27])) ;
    aoi22 ix404 (.Y (nx392), .A0 (a[27]), .A1 (b[27]), .B0 (nx390), .B1 (nx391)
          ) ;
    oai22 ix405 (.Y (nx393), .A0 (nx391), .A1 (a[27]), .B0 (nx390), .B1 (b[27])
          ) ;
    nand02_2x ix406 (.Y (nx394), .A0 (nx393), .A1 (nx389)) ;
    oai21 reg_s_27 (.Y (s[27]), .A0 (nx389), .A1 (nx392), .B0 (nx394)) ;
    inv02 ix407 (.Y (nx395), .A (nx389)) ;
    oai22 reg_nx351 (.Y (nx351), .A0 (nx390), .A1 (nx391), .B0 (a[27]), .B1 (
          b[27])) ;
    ao22 reg_nx342 (.Y (nx342), .A0 (nx388), .A1 (nx387), .B0 (nx339), .B1 (
         nx388)) ;
    inv01 reg_nx192 (.Y (nx192), .A (nx387)) ;
    oai22 reg_nx330 (.Y (nx330), .A0 (nx386), .A1 (nx176), .B0 (nx386), .B1 (
          nx178)) ;
    nor02_2x ix408 (.Y (nx396), .A0 (a[24]), .A1 (b[24])) ;
    ao21 reg_nx333 (.Y (nx333), .A0 (a[24]), .A1 (b[24]), .B0 (nx396)) ;
endmodule


module MuxLayer ( img_data_0__31, img_data_0__30, img_data_0__29, img_data_0__28, 
                  img_data_0__27, img_data_0__26, img_data_0__25, img_data_0__24, 
                  img_data_0__23, img_data_0__22, img_data_0__21, img_data_0__20, 
                  img_data_0__19, img_data_0__18, img_data_0__17, img_data_0__16, 
                  img_data_0__15, img_data_0__14, img_data_0__13, img_data_0__12, 
                  img_data_0__11, img_data_0__10, img_data_0__9, img_data_0__8, 
                  img_data_0__7, img_data_0__6, img_data_0__5, img_data_0__4, 
                  img_data_0__3, img_data_0__2, img_data_0__1, img_data_0__0, 
                  img_data_1__31, img_data_1__30, img_data_1__29, img_data_1__28, 
                  img_data_1__27, img_data_1__26, img_data_1__25, img_data_1__24, 
                  img_data_1__23, img_data_1__22, img_data_1__21, img_data_1__20, 
                  img_data_1__19, img_data_1__18, img_data_1__17, img_data_1__16, 
                  img_data_1__15, img_data_1__14, img_data_1__13, img_data_1__12, 
                  img_data_1__11, img_data_1__10, img_data_1__9, img_data_1__8, 
                  img_data_1__7, img_data_1__6, img_data_1__5, img_data_1__4, 
                  img_data_1__3, img_data_1__2, img_data_1__1, img_data_1__0, 
                  img_data_2__31, img_data_2__30, img_data_2__29, img_data_2__28, 
                  img_data_2__27, img_data_2__26, img_data_2__25, img_data_2__24, 
                  img_data_2__23, img_data_2__22, img_data_2__21, img_data_2__20, 
                  img_data_2__19, img_data_2__18, img_data_2__17, img_data_2__16, 
                  img_data_2__15, img_data_2__14, img_data_2__13, img_data_2__12, 
                  img_data_2__11, img_data_2__10, img_data_2__9, img_data_2__8, 
                  img_data_2__7, img_data_2__6, img_data_2__5, img_data_2__4, 
                  img_data_2__3, img_data_2__2, img_data_2__1, img_data_2__0, 
                  img_data_3__31, img_data_3__30, img_data_3__29, img_data_3__28, 
                  img_data_3__27, img_data_3__26, img_data_3__25, img_data_3__24, 
                  img_data_3__23, img_data_3__22, img_data_3__21, img_data_3__20, 
                  img_data_3__19, img_data_3__18, img_data_3__17, img_data_3__16, 
                  img_data_3__15, img_data_3__14, img_data_3__13, img_data_3__12, 
                  img_data_3__11, img_data_3__10, img_data_3__9, img_data_3__8, 
                  img_data_3__7, img_data_3__6, img_data_3__5, img_data_3__4, 
                  img_data_3__3, img_data_3__2, img_data_3__1, img_data_3__0, 
                  img_data_4__31, img_data_4__30, img_data_4__29, img_data_4__28, 
                  img_data_4__27, img_data_4__26, img_data_4__25, img_data_4__24, 
                  img_data_4__23, img_data_4__22, img_data_4__21, img_data_4__20, 
                  img_data_4__19, img_data_4__18, img_data_4__17, img_data_4__16, 
                  img_data_4__15, img_data_4__14, img_data_4__13, img_data_4__12, 
                  img_data_4__11, img_data_4__10, img_data_4__9, img_data_4__8, 
                  img_data_4__7, img_data_4__6, img_data_4__5, img_data_4__4, 
                  img_data_4__3, img_data_4__2, img_data_4__1, img_data_4__0, 
                  img_data_5__31, img_data_5__30, img_data_5__29, img_data_5__28, 
                  img_data_5__27, img_data_5__26, img_data_5__25, img_data_5__24, 
                  img_data_5__23, img_data_5__22, img_data_5__21, img_data_5__20, 
                  img_data_5__19, img_data_5__18, img_data_5__17, img_data_5__16, 
                  img_data_5__15, img_data_5__14, img_data_5__13, img_data_5__12, 
                  img_data_5__11, img_data_5__10, img_data_5__9, img_data_5__8, 
                  img_data_5__7, img_data_5__6, img_data_5__5, img_data_5__4, 
                  img_data_5__3, img_data_5__2, img_data_5__1, img_data_5__0, 
                  img_data_6__31, img_data_6__30, img_data_6__29, img_data_6__28, 
                  img_data_6__27, img_data_6__26, img_data_6__25, img_data_6__24, 
                  img_data_6__23, img_data_6__22, img_data_6__21, img_data_6__20, 
                  img_data_6__19, img_data_6__18, img_data_6__17, img_data_6__16, 
                  img_data_6__15, img_data_6__14, img_data_6__13, img_data_6__12, 
                  img_data_6__11, img_data_6__10, img_data_6__9, img_data_6__8, 
                  img_data_6__7, img_data_6__6, img_data_6__5, img_data_6__4, 
                  img_data_6__3, img_data_6__2, img_data_6__1, img_data_6__0, 
                  img_data_7__31, img_data_7__30, img_data_7__29, img_data_7__28, 
                  img_data_7__27, img_data_7__26, img_data_7__25, img_data_7__24, 
                  img_data_7__23, img_data_7__22, img_data_7__21, img_data_7__20, 
                  img_data_7__19, img_data_7__18, img_data_7__17, img_data_7__16, 
                  img_data_7__15, img_data_7__14, img_data_7__13, img_data_7__12, 
                  img_data_7__11, img_data_7__10, img_data_7__9, img_data_7__8, 
                  img_data_7__7, img_data_7__6, img_data_7__5, img_data_7__4, 
                  img_data_7__3, img_data_7__2, img_data_7__1, img_data_7__0, 
                  img_data_8__31, img_data_8__30, img_data_8__29, img_data_8__28, 
                  img_data_8__27, img_data_8__26, img_data_8__25, img_data_8__24, 
                  img_data_8__23, img_data_8__22, img_data_8__21, img_data_8__20, 
                  img_data_8__19, img_data_8__18, img_data_8__17, img_data_8__16, 
                  img_data_8__15, img_data_8__14, img_data_8__13, img_data_8__12, 
                  img_data_8__11, img_data_8__10, img_data_8__9, img_data_8__8, 
                  img_data_8__7, img_data_8__6, img_data_8__5, img_data_8__4, 
                  img_data_8__3, img_data_8__2, img_data_8__1, img_data_8__0, 
                  img_data_9__31, img_data_9__30, img_data_9__29, img_data_9__28, 
                  img_data_9__27, img_data_9__26, img_data_9__25, img_data_9__24, 
                  img_data_9__23, img_data_9__22, img_data_9__21, img_data_9__20, 
                  img_data_9__19, img_data_9__18, img_data_9__17, img_data_9__16, 
                  img_data_9__15, img_data_9__14, img_data_9__13, img_data_9__12, 
                  img_data_9__11, img_data_9__10, img_data_9__9, img_data_9__8, 
                  img_data_9__7, img_data_9__6, img_data_9__5, img_data_9__4, 
                  img_data_9__3, img_data_9__2, img_data_9__1, img_data_9__0, 
                  img_data_10__31, img_data_10__30, img_data_10__29, 
                  img_data_10__28, img_data_10__27, img_data_10__26, 
                  img_data_10__25, img_data_10__24, img_data_10__23, 
                  img_data_10__22, img_data_10__21, img_data_10__20, 
                  img_data_10__19, img_data_10__18, img_data_10__17, 
                  img_data_10__16, img_data_10__15, img_data_10__14, 
                  img_data_10__13, img_data_10__12, img_data_10__11, 
                  img_data_10__10, img_data_10__9, img_data_10__8, 
                  img_data_10__7, img_data_10__6, img_data_10__5, img_data_10__4, 
                  img_data_10__3, img_data_10__2, img_data_10__1, img_data_10__0, 
                  img_data_11__31, img_data_11__30, img_data_11__29, 
                  img_data_11__28, img_data_11__27, img_data_11__26, 
                  img_data_11__25, img_data_11__24, img_data_11__23, 
                  img_data_11__22, img_data_11__21, img_data_11__20, 
                  img_data_11__19, img_data_11__18, img_data_11__17, 
                  img_data_11__16, img_data_11__15, img_data_11__14, 
                  img_data_11__13, img_data_11__12, img_data_11__11, 
                  img_data_11__10, img_data_11__9, img_data_11__8, 
                  img_data_11__7, img_data_11__6, img_data_11__5, img_data_11__4, 
                  img_data_11__3, img_data_11__2, img_data_11__1, img_data_11__0, 
                  img_data_12__31, img_data_12__30, img_data_12__29, 
                  img_data_12__28, img_data_12__27, img_data_12__26, 
                  img_data_12__25, img_data_12__24, img_data_12__23, 
                  img_data_12__22, img_data_12__21, img_data_12__20, 
                  img_data_12__19, img_data_12__18, img_data_12__17, 
                  img_data_12__16, img_data_12__15, img_data_12__14, 
                  img_data_12__13, img_data_12__12, img_data_12__11, 
                  img_data_12__10, img_data_12__9, img_data_12__8, 
                  img_data_12__7, img_data_12__6, img_data_12__5, img_data_12__4, 
                  img_data_12__3, img_data_12__2, img_data_12__1, img_data_12__0, 
                  img_data_13__31, img_data_13__30, img_data_13__29, 
                  img_data_13__28, img_data_13__27, img_data_13__26, 
                  img_data_13__25, img_data_13__24, img_data_13__23, 
                  img_data_13__22, img_data_13__21, img_data_13__20, 
                  img_data_13__19, img_data_13__18, img_data_13__17, 
                  img_data_13__16, img_data_13__15, img_data_13__14, 
                  img_data_13__13, img_data_13__12, img_data_13__11, 
                  img_data_13__10, img_data_13__9, img_data_13__8, 
                  img_data_13__7, img_data_13__6, img_data_13__5, img_data_13__4, 
                  img_data_13__3, img_data_13__2, img_data_13__1, img_data_13__0, 
                  img_data_14__31, img_data_14__30, img_data_14__29, 
                  img_data_14__28, img_data_14__27, img_data_14__26, 
                  img_data_14__25, img_data_14__24, img_data_14__23, 
                  img_data_14__22, img_data_14__21, img_data_14__20, 
                  img_data_14__19, img_data_14__18, img_data_14__17, 
                  img_data_14__16, img_data_14__15, img_data_14__14, 
                  img_data_14__13, img_data_14__12, img_data_14__11, 
                  img_data_14__10, img_data_14__9, img_data_14__8, 
                  img_data_14__7, img_data_14__6, img_data_14__5, img_data_14__4, 
                  img_data_14__3, img_data_14__2, img_data_14__1, img_data_14__0, 
                  img_data_15__31, img_data_15__30, img_data_15__29, 
                  img_data_15__28, img_data_15__27, img_data_15__26, 
                  img_data_15__25, img_data_15__24, img_data_15__23, 
                  img_data_15__22, img_data_15__21, img_data_15__20, 
                  img_data_15__19, img_data_15__18, img_data_15__17, 
                  img_data_15__16, img_data_15__15, img_data_15__14, 
                  img_data_15__13, img_data_15__12, img_data_15__11, 
                  img_data_15__10, img_data_15__9, img_data_15__8, 
                  img_data_15__7, img_data_15__6, img_data_15__5, img_data_15__4, 
                  img_data_15__3, img_data_15__2, img_data_15__1, img_data_15__0, 
                  img_data_16__31, img_data_16__30, img_data_16__29, 
                  img_data_16__28, img_data_16__27, img_data_16__26, 
                  img_data_16__25, img_data_16__24, img_data_16__23, 
                  img_data_16__22, img_data_16__21, img_data_16__20, 
                  img_data_16__19, img_data_16__18, img_data_16__17, 
                  img_data_16__16, img_data_16__15, img_data_16__14, 
                  img_data_16__13, img_data_16__12, img_data_16__11, 
                  img_data_16__10, img_data_16__9, img_data_16__8, 
                  img_data_16__7, img_data_16__6, img_data_16__5, img_data_16__4, 
                  img_data_16__3, img_data_16__2, img_data_16__1, img_data_16__0, 
                  img_data_17__31, img_data_17__30, img_data_17__29, 
                  img_data_17__28, img_data_17__27, img_data_17__26, 
                  img_data_17__25, img_data_17__24, img_data_17__23, 
                  img_data_17__22, img_data_17__21, img_data_17__20, 
                  img_data_17__19, img_data_17__18, img_data_17__17, 
                  img_data_17__16, img_data_17__15, img_data_17__14, 
                  img_data_17__13, img_data_17__12, img_data_17__11, 
                  img_data_17__10, img_data_17__9, img_data_17__8, 
                  img_data_17__7, img_data_17__6, img_data_17__5, img_data_17__4, 
                  img_data_17__3, img_data_17__2, img_data_17__1, img_data_17__0, 
                  img_data_18__31, img_data_18__30, img_data_18__29, 
                  img_data_18__28, img_data_18__27, img_data_18__26, 
                  img_data_18__25, img_data_18__24, img_data_18__23, 
                  img_data_18__22, img_data_18__21, img_data_18__20, 
                  img_data_18__19, img_data_18__18, img_data_18__17, 
                  img_data_18__16, img_data_18__15, img_data_18__14, 
                  img_data_18__13, img_data_18__12, img_data_18__11, 
                  img_data_18__10, img_data_18__9, img_data_18__8, 
                  img_data_18__7, img_data_18__6, img_data_18__5, img_data_18__4, 
                  img_data_18__3, img_data_18__2, img_data_18__1, img_data_18__0, 
                  img_data_19__31, img_data_19__30, img_data_19__29, 
                  img_data_19__28, img_data_19__27, img_data_19__26, 
                  img_data_19__25, img_data_19__24, img_data_19__23, 
                  img_data_19__22, img_data_19__21, img_data_19__20, 
                  img_data_19__19, img_data_19__18, img_data_19__17, 
                  img_data_19__16, img_data_19__15, img_data_19__14, 
                  img_data_19__13, img_data_19__12, img_data_19__11, 
                  img_data_19__10, img_data_19__9, img_data_19__8, 
                  img_data_19__7, img_data_19__6, img_data_19__5, img_data_19__4, 
                  img_data_19__3, img_data_19__2, img_data_19__1, img_data_19__0, 
                  img_data_20__31, img_data_20__30, img_data_20__29, 
                  img_data_20__28, img_data_20__27, img_data_20__26, 
                  img_data_20__25, img_data_20__24, img_data_20__23, 
                  img_data_20__22, img_data_20__21, img_data_20__20, 
                  img_data_20__19, img_data_20__18, img_data_20__17, 
                  img_data_20__16, img_data_20__15, img_data_20__14, 
                  img_data_20__13, img_data_20__12, img_data_20__11, 
                  img_data_20__10, img_data_20__9, img_data_20__8, 
                  img_data_20__7, img_data_20__6, img_data_20__5, img_data_20__4, 
                  img_data_20__3, img_data_20__2, img_data_20__1, img_data_20__0, 
                  img_data_21__31, img_data_21__30, img_data_21__29, 
                  img_data_21__28, img_data_21__27, img_data_21__26, 
                  img_data_21__25, img_data_21__24, img_data_21__23, 
                  img_data_21__22, img_data_21__21, img_data_21__20, 
                  img_data_21__19, img_data_21__18, img_data_21__17, 
                  img_data_21__16, img_data_21__15, img_data_21__14, 
                  img_data_21__13, img_data_21__12, img_data_21__11, 
                  img_data_21__10, img_data_21__9, img_data_21__8, 
                  img_data_21__7, img_data_21__6, img_data_21__5, img_data_21__4, 
                  img_data_21__3, img_data_21__2, img_data_21__1, img_data_21__0, 
                  img_data_22__31, img_data_22__30, img_data_22__29, 
                  img_data_22__28, img_data_22__27, img_data_22__26, 
                  img_data_22__25, img_data_22__24, img_data_22__23, 
                  img_data_22__22, img_data_22__21, img_data_22__20, 
                  img_data_22__19, img_data_22__18, img_data_22__17, 
                  img_data_22__16, img_data_22__15, img_data_22__14, 
                  img_data_22__13, img_data_22__12, img_data_22__11, 
                  img_data_22__10, img_data_22__9, img_data_22__8, 
                  img_data_22__7, img_data_22__6, img_data_22__5, img_data_22__4, 
                  img_data_22__3, img_data_22__2, img_data_22__1, img_data_22__0, 
                  img_data_23__31, img_data_23__30, img_data_23__29, 
                  img_data_23__28, img_data_23__27, img_data_23__26, 
                  img_data_23__25, img_data_23__24, img_data_23__23, 
                  img_data_23__22, img_data_23__21, img_data_23__20, 
                  img_data_23__19, img_data_23__18, img_data_23__17, 
                  img_data_23__16, img_data_23__15, img_data_23__14, 
                  img_data_23__13, img_data_23__12, img_data_23__11, 
                  img_data_23__10, img_data_23__9, img_data_23__8, 
                  img_data_23__7, img_data_23__6, img_data_23__5, img_data_23__4, 
                  img_data_23__3, img_data_23__2, img_data_23__1, img_data_23__0, 
                  img_data_24__31, img_data_24__30, img_data_24__29, 
                  img_data_24__28, img_data_24__27, img_data_24__26, 
                  img_data_24__25, img_data_24__24, img_data_24__23, 
                  img_data_24__22, img_data_24__21, img_data_24__20, 
                  img_data_24__19, img_data_24__18, img_data_24__17, 
                  img_data_24__16, img_data_24__15, img_data_24__14, 
                  img_data_24__13, img_data_24__12, img_data_24__11, 
                  img_data_24__10, img_data_24__9, img_data_24__8, 
                  img_data_24__7, img_data_24__6, img_data_24__5, img_data_24__4, 
                  img_data_24__3, img_data_24__2, img_data_24__1, img_data_24__0, 
                  filter_data_0__31, filter_data_0__30, filter_data_0__29, 
                  filter_data_0__28, filter_data_0__27, filter_data_0__26, 
                  filter_data_0__25, filter_data_0__24, filter_data_0__23, 
                  filter_data_0__22, filter_data_0__21, filter_data_0__20, 
                  filter_data_0__19, filter_data_0__18, filter_data_0__17, 
                  filter_data_0__16, filter_data_0__15, filter_data_0__14, 
                  filter_data_0__13, filter_data_0__12, filter_data_0__11, 
                  filter_data_0__10, filter_data_0__9, filter_data_0__8, 
                  filter_data_0__7, filter_data_0__6, filter_data_0__5, 
                  filter_data_0__4, filter_data_0__3, filter_data_0__2, 
                  filter_data_0__1, filter_data_0__0, filter_data_1__31, 
                  filter_data_1__30, filter_data_1__29, filter_data_1__28, 
                  filter_data_1__27, filter_data_1__26, filter_data_1__25, 
                  filter_data_1__24, filter_data_1__23, filter_data_1__22, 
                  filter_data_1__21, filter_data_1__20, filter_data_1__19, 
                  filter_data_1__18, filter_data_1__17, filter_data_1__16, 
                  filter_data_1__15, filter_data_1__14, filter_data_1__13, 
                  filter_data_1__12, filter_data_1__11, filter_data_1__10, 
                  filter_data_1__9, filter_data_1__8, filter_data_1__7, 
                  filter_data_1__6, filter_data_1__5, filter_data_1__4, 
                  filter_data_1__3, filter_data_1__2, filter_data_1__1, 
                  filter_data_1__0, filter_data_2__31, filter_data_2__30, 
                  filter_data_2__29, filter_data_2__28, filter_data_2__27, 
                  filter_data_2__26, filter_data_2__25, filter_data_2__24, 
                  filter_data_2__23, filter_data_2__22, filter_data_2__21, 
                  filter_data_2__20, filter_data_2__19, filter_data_2__18, 
                  filter_data_2__17, filter_data_2__16, filter_data_2__15, 
                  filter_data_2__14, filter_data_2__13, filter_data_2__12, 
                  filter_data_2__11, filter_data_2__10, filter_data_2__9, 
                  filter_data_2__8, filter_data_2__7, filter_data_2__6, 
                  filter_data_2__5, filter_data_2__4, filter_data_2__3, 
                  filter_data_2__2, filter_data_2__1, filter_data_2__0, 
                  filter_data_3__31, filter_data_3__30, filter_data_3__29, 
                  filter_data_3__28, filter_data_3__27, filter_data_3__26, 
                  filter_data_3__25, filter_data_3__24, filter_data_3__23, 
                  filter_data_3__22, filter_data_3__21, filter_data_3__20, 
                  filter_data_3__19, filter_data_3__18, filter_data_3__17, 
                  filter_data_3__16, filter_data_3__15, filter_data_3__14, 
                  filter_data_3__13, filter_data_3__12, filter_data_3__11, 
                  filter_data_3__10, filter_data_3__9, filter_data_3__8, 
                  filter_data_3__7, filter_data_3__6, filter_data_3__5, 
                  filter_data_3__4, filter_data_3__3, filter_data_3__2, 
                  filter_data_3__1, filter_data_3__0, filter_data_4__31, 
                  filter_data_4__30, filter_data_4__29, filter_data_4__28, 
                  filter_data_4__27, filter_data_4__26, filter_data_4__25, 
                  filter_data_4__24, filter_data_4__23, filter_data_4__22, 
                  filter_data_4__21, filter_data_4__20, filter_data_4__19, 
                  filter_data_4__18, filter_data_4__17, filter_data_4__16, 
                  filter_data_4__15, filter_data_4__14, filter_data_4__13, 
                  filter_data_4__12, filter_data_4__11, filter_data_4__10, 
                  filter_data_4__9, filter_data_4__8, filter_data_4__7, 
                  filter_data_4__6, filter_data_4__5, filter_data_4__4, 
                  filter_data_4__3, filter_data_4__2, filter_data_4__1, 
                  filter_data_4__0, filter_data_5__31, filter_data_5__30, 
                  filter_data_5__29, filter_data_5__28, filter_data_5__27, 
                  filter_data_5__26, filter_data_5__25, filter_data_5__24, 
                  filter_data_5__23, filter_data_5__22, filter_data_5__21, 
                  filter_data_5__20, filter_data_5__19, filter_data_5__18, 
                  filter_data_5__17, filter_data_5__16, filter_data_5__15, 
                  filter_data_5__14, filter_data_5__13, filter_data_5__12, 
                  filter_data_5__11, filter_data_5__10, filter_data_5__9, 
                  filter_data_5__8, filter_data_5__7, filter_data_5__6, 
                  filter_data_5__5, filter_data_5__4, filter_data_5__3, 
                  filter_data_5__2, filter_data_5__1, filter_data_5__0, 
                  filter_data_6__31, filter_data_6__30, filter_data_6__29, 
                  filter_data_6__28, filter_data_6__27, filter_data_6__26, 
                  filter_data_6__25, filter_data_6__24, filter_data_6__23, 
                  filter_data_6__22, filter_data_6__21, filter_data_6__20, 
                  filter_data_6__19, filter_data_6__18, filter_data_6__17, 
                  filter_data_6__16, filter_data_6__15, filter_data_6__14, 
                  filter_data_6__13, filter_data_6__12, filter_data_6__11, 
                  filter_data_6__10, filter_data_6__9, filter_data_6__8, 
                  filter_data_6__7, filter_data_6__6, filter_data_6__5, 
                  filter_data_6__4, filter_data_6__3, filter_data_6__2, 
                  filter_data_6__1, filter_data_6__0, filter_data_7__31, 
                  filter_data_7__30, filter_data_7__29, filter_data_7__28, 
                  filter_data_7__27, filter_data_7__26, filter_data_7__25, 
                  filter_data_7__24, filter_data_7__23, filter_data_7__22, 
                  filter_data_7__21, filter_data_7__20, filter_data_7__19, 
                  filter_data_7__18, filter_data_7__17, filter_data_7__16, 
                  filter_data_7__15, filter_data_7__14, filter_data_7__13, 
                  filter_data_7__12, filter_data_7__11, filter_data_7__10, 
                  filter_data_7__9, filter_data_7__8, filter_data_7__7, 
                  filter_data_7__6, filter_data_7__5, filter_data_7__4, 
                  filter_data_7__3, filter_data_7__2, filter_data_7__1, 
                  filter_data_7__0, filter_data_8__31, filter_data_8__30, 
                  filter_data_8__29, filter_data_8__28, filter_data_8__27, 
                  filter_data_8__26, filter_data_8__25, filter_data_8__24, 
                  filter_data_8__23, filter_data_8__22, filter_data_8__21, 
                  filter_data_8__20, filter_data_8__19, filter_data_8__18, 
                  filter_data_8__17, filter_data_8__16, filter_data_8__15, 
                  filter_data_8__14, filter_data_8__13, filter_data_8__12, 
                  filter_data_8__11, filter_data_8__10, filter_data_8__9, 
                  filter_data_8__8, filter_data_8__7, filter_data_8__6, 
                  filter_data_8__5, filter_data_8__4, filter_data_8__3, 
                  filter_data_8__2, filter_data_8__1, filter_data_8__0, 
                  filter_data_9__31, filter_data_9__30, filter_data_9__29, 
                  filter_data_9__28, filter_data_9__27, filter_data_9__26, 
                  filter_data_9__25, filter_data_9__24, filter_data_9__23, 
                  filter_data_9__22, filter_data_9__21, filter_data_9__20, 
                  filter_data_9__19, filter_data_9__18, filter_data_9__17, 
                  filter_data_9__16, filter_data_9__15, filter_data_9__14, 
                  filter_data_9__13, filter_data_9__12, filter_data_9__11, 
                  filter_data_9__10, filter_data_9__9, filter_data_9__8, 
                  filter_data_9__7, filter_data_9__6, filter_data_9__5, 
                  filter_data_9__4, filter_data_9__3, filter_data_9__2, 
                  filter_data_9__1, filter_data_9__0, filter_data_10__31, 
                  filter_data_10__30, filter_data_10__29, filter_data_10__28, 
                  filter_data_10__27, filter_data_10__26, filter_data_10__25, 
                  filter_data_10__24, filter_data_10__23, filter_data_10__22, 
                  filter_data_10__21, filter_data_10__20, filter_data_10__19, 
                  filter_data_10__18, filter_data_10__17, filter_data_10__16, 
                  filter_data_10__15, filter_data_10__14, filter_data_10__13, 
                  filter_data_10__12, filter_data_10__11, filter_data_10__10, 
                  filter_data_10__9, filter_data_10__8, filter_data_10__7, 
                  filter_data_10__6, filter_data_10__5, filter_data_10__4, 
                  filter_data_10__3, filter_data_10__2, filter_data_10__1, 
                  filter_data_10__0, filter_data_11__31, filter_data_11__30, 
                  filter_data_11__29, filter_data_11__28, filter_data_11__27, 
                  filter_data_11__26, filter_data_11__25, filter_data_11__24, 
                  filter_data_11__23, filter_data_11__22, filter_data_11__21, 
                  filter_data_11__20, filter_data_11__19, filter_data_11__18, 
                  filter_data_11__17, filter_data_11__16, filter_data_11__15, 
                  filter_data_11__14, filter_data_11__13, filter_data_11__12, 
                  filter_data_11__11, filter_data_11__10, filter_data_11__9, 
                  filter_data_11__8, filter_data_11__7, filter_data_11__6, 
                  filter_data_11__5, filter_data_11__4, filter_data_11__3, 
                  filter_data_11__2, filter_data_11__1, filter_data_11__0, 
                  filter_data_12__31, filter_data_12__30, filter_data_12__29, 
                  filter_data_12__28, filter_data_12__27, filter_data_12__26, 
                  filter_data_12__25, filter_data_12__24, filter_data_12__23, 
                  filter_data_12__22, filter_data_12__21, filter_data_12__20, 
                  filter_data_12__19, filter_data_12__18, filter_data_12__17, 
                  filter_data_12__16, filter_data_12__15, filter_data_12__14, 
                  filter_data_12__13, filter_data_12__12, filter_data_12__11, 
                  filter_data_12__10, filter_data_12__9, filter_data_12__8, 
                  filter_data_12__7, filter_data_12__6, filter_data_12__5, 
                  filter_data_12__4, filter_data_12__3, filter_data_12__2, 
                  filter_data_12__1, filter_data_12__0, filter_data_13__31, 
                  filter_data_13__30, filter_data_13__29, filter_data_13__28, 
                  filter_data_13__27, filter_data_13__26, filter_data_13__25, 
                  filter_data_13__24, filter_data_13__23, filter_data_13__22, 
                  filter_data_13__21, filter_data_13__20, filter_data_13__19, 
                  filter_data_13__18, filter_data_13__17, filter_data_13__16, 
                  filter_data_13__15, filter_data_13__14, filter_data_13__13, 
                  filter_data_13__12, filter_data_13__11, filter_data_13__10, 
                  filter_data_13__9, filter_data_13__8, filter_data_13__7, 
                  filter_data_13__6, filter_data_13__5, filter_data_13__4, 
                  filter_data_13__3, filter_data_13__2, filter_data_13__1, 
                  filter_data_13__0, filter_data_14__31, filter_data_14__30, 
                  filter_data_14__29, filter_data_14__28, filter_data_14__27, 
                  filter_data_14__26, filter_data_14__25, filter_data_14__24, 
                  filter_data_14__23, filter_data_14__22, filter_data_14__21, 
                  filter_data_14__20, filter_data_14__19, filter_data_14__18, 
                  filter_data_14__17, filter_data_14__16, filter_data_14__15, 
                  filter_data_14__14, filter_data_14__13, filter_data_14__12, 
                  filter_data_14__11, filter_data_14__10, filter_data_14__9, 
                  filter_data_14__8, filter_data_14__7, filter_data_14__6, 
                  filter_data_14__5, filter_data_14__4, filter_data_14__3, 
                  filter_data_14__2, filter_data_14__1, filter_data_14__0, 
                  filter_data_15__31, filter_data_15__30, filter_data_15__29, 
                  filter_data_15__28, filter_data_15__27, filter_data_15__26, 
                  filter_data_15__25, filter_data_15__24, filter_data_15__23, 
                  filter_data_15__22, filter_data_15__21, filter_data_15__20, 
                  filter_data_15__19, filter_data_15__18, filter_data_15__17, 
                  filter_data_15__16, filter_data_15__15, filter_data_15__14, 
                  filter_data_15__13, filter_data_15__12, filter_data_15__11, 
                  filter_data_15__10, filter_data_15__9, filter_data_15__8, 
                  filter_data_15__7, filter_data_15__6, filter_data_15__5, 
                  filter_data_15__4, filter_data_15__3, filter_data_15__2, 
                  filter_data_15__1, filter_data_15__0, filter_data_16__31, 
                  filter_data_16__30, filter_data_16__29, filter_data_16__28, 
                  filter_data_16__27, filter_data_16__26, filter_data_16__25, 
                  filter_data_16__24, filter_data_16__23, filter_data_16__22, 
                  filter_data_16__21, filter_data_16__20, filter_data_16__19, 
                  filter_data_16__18, filter_data_16__17, filter_data_16__16, 
                  filter_data_16__15, filter_data_16__14, filter_data_16__13, 
                  filter_data_16__12, filter_data_16__11, filter_data_16__10, 
                  filter_data_16__9, filter_data_16__8, filter_data_16__7, 
                  filter_data_16__6, filter_data_16__5, filter_data_16__4, 
                  filter_data_16__3, filter_data_16__2, filter_data_16__1, 
                  filter_data_16__0, filter_data_17__31, filter_data_17__30, 
                  filter_data_17__29, filter_data_17__28, filter_data_17__27, 
                  filter_data_17__26, filter_data_17__25, filter_data_17__24, 
                  filter_data_17__23, filter_data_17__22, filter_data_17__21, 
                  filter_data_17__20, filter_data_17__19, filter_data_17__18, 
                  filter_data_17__17, filter_data_17__16, filter_data_17__15, 
                  filter_data_17__14, filter_data_17__13, filter_data_17__12, 
                  filter_data_17__11, filter_data_17__10, filter_data_17__9, 
                  filter_data_17__8, filter_data_17__7, filter_data_17__6, 
                  filter_data_17__5, filter_data_17__4, filter_data_17__3, 
                  filter_data_17__2, filter_data_17__1, filter_data_17__0, 
                  filter_data_18__31, filter_data_18__30, filter_data_18__29, 
                  filter_data_18__28, filter_data_18__27, filter_data_18__26, 
                  filter_data_18__25, filter_data_18__24, filter_data_18__23, 
                  filter_data_18__22, filter_data_18__21, filter_data_18__20, 
                  filter_data_18__19, filter_data_18__18, filter_data_18__17, 
                  filter_data_18__16, filter_data_18__15, filter_data_18__14, 
                  filter_data_18__13, filter_data_18__12, filter_data_18__11, 
                  filter_data_18__10, filter_data_18__9, filter_data_18__8, 
                  filter_data_18__7, filter_data_18__6, filter_data_18__5, 
                  filter_data_18__4, filter_data_18__3, filter_data_18__2, 
                  filter_data_18__1, filter_data_18__0, filter_data_19__31, 
                  filter_data_19__30, filter_data_19__29, filter_data_19__28, 
                  filter_data_19__27, filter_data_19__26, filter_data_19__25, 
                  filter_data_19__24, filter_data_19__23, filter_data_19__22, 
                  filter_data_19__21, filter_data_19__20, filter_data_19__19, 
                  filter_data_19__18, filter_data_19__17, filter_data_19__16, 
                  filter_data_19__15, filter_data_19__14, filter_data_19__13, 
                  filter_data_19__12, filter_data_19__11, filter_data_19__10, 
                  filter_data_19__9, filter_data_19__8, filter_data_19__7, 
                  filter_data_19__6, filter_data_19__5, filter_data_19__4, 
                  filter_data_19__3, filter_data_19__2, filter_data_19__1, 
                  filter_data_19__0, filter_data_20__31, filter_data_20__30, 
                  filter_data_20__29, filter_data_20__28, filter_data_20__27, 
                  filter_data_20__26, filter_data_20__25, filter_data_20__24, 
                  filter_data_20__23, filter_data_20__22, filter_data_20__21, 
                  filter_data_20__20, filter_data_20__19, filter_data_20__18, 
                  filter_data_20__17, filter_data_20__16, filter_data_20__15, 
                  filter_data_20__14, filter_data_20__13, filter_data_20__12, 
                  filter_data_20__11, filter_data_20__10, filter_data_20__9, 
                  filter_data_20__8, filter_data_20__7, filter_data_20__6, 
                  filter_data_20__5, filter_data_20__4, filter_data_20__3, 
                  filter_data_20__2, filter_data_20__1, filter_data_20__0, 
                  filter_data_21__31, filter_data_21__30, filter_data_21__29, 
                  filter_data_21__28, filter_data_21__27, filter_data_21__26, 
                  filter_data_21__25, filter_data_21__24, filter_data_21__23, 
                  filter_data_21__22, filter_data_21__21, filter_data_21__20, 
                  filter_data_21__19, filter_data_21__18, filter_data_21__17, 
                  filter_data_21__16, filter_data_21__15, filter_data_21__14, 
                  filter_data_21__13, filter_data_21__12, filter_data_21__11, 
                  filter_data_21__10, filter_data_21__9, filter_data_21__8, 
                  filter_data_21__7, filter_data_21__6, filter_data_21__5, 
                  filter_data_21__4, filter_data_21__3, filter_data_21__2, 
                  filter_data_21__1, filter_data_21__0, filter_data_22__31, 
                  filter_data_22__30, filter_data_22__29, filter_data_22__28, 
                  filter_data_22__27, filter_data_22__26, filter_data_22__25, 
                  filter_data_22__24, filter_data_22__23, filter_data_22__22, 
                  filter_data_22__21, filter_data_22__20, filter_data_22__19, 
                  filter_data_22__18, filter_data_22__17, filter_data_22__16, 
                  filter_data_22__15, filter_data_22__14, filter_data_22__13, 
                  filter_data_22__12, filter_data_22__11, filter_data_22__10, 
                  filter_data_22__9, filter_data_22__8, filter_data_22__7, 
                  filter_data_22__6, filter_data_22__5, filter_data_22__4, 
                  filter_data_22__3, filter_data_22__2, filter_data_22__1, 
                  filter_data_22__0, filter_data_23__31, filter_data_23__30, 
                  filter_data_23__29, filter_data_23__28, filter_data_23__27, 
                  filter_data_23__26, filter_data_23__25, filter_data_23__24, 
                  filter_data_23__23, filter_data_23__22, filter_data_23__21, 
                  filter_data_23__20, filter_data_23__19, filter_data_23__18, 
                  filter_data_23__17, filter_data_23__16, filter_data_23__15, 
                  filter_data_23__14, filter_data_23__13, filter_data_23__12, 
                  filter_data_23__11, filter_data_23__10, filter_data_23__9, 
                  filter_data_23__8, filter_data_23__7, filter_data_23__6, 
                  filter_data_23__5, filter_data_23__4, filter_data_23__3, 
                  filter_data_23__2, filter_data_23__1, filter_data_23__0, 
                  filter_data_24__31, filter_data_24__30, filter_data_24__29, 
                  filter_data_24__28, filter_data_24__27, filter_data_24__26, 
                  filter_data_24__25, filter_data_24__24, filter_data_24__23, 
                  filter_data_24__22, filter_data_24__21, filter_data_24__20, 
                  filter_data_24__19, filter_data_24__18, filter_data_24__17, 
                  filter_data_24__16, filter_data_24__15, filter_data_24__14, 
                  filter_data_24__13, filter_data_24__12, filter_data_24__11, 
                  filter_data_24__10, filter_data_24__9, filter_data_24__8, 
                  filter_data_24__7, filter_data_24__6, filter_data_24__5, 
                  filter_data_24__4, filter_data_24__3, filter_data_24__2, 
                  filter_data_24__1, filter_data_24__0, filter_size, 
                  ordered_img_data_0__31, ordered_img_data_0__30, 
                  ordered_img_data_0__29, ordered_img_data_0__28, 
                  ordered_img_data_0__27, ordered_img_data_0__26, 
                  ordered_img_data_0__25, ordered_img_data_0__24, 
                  ordered_img_data_0__23, ordered_img_data_0__22, 
                  ordered_img_data_0__21, ordered_img_data_0__20, 
                  ordered_img_data_0__19, ordered_img_data_0__18, 
                  ordered_img_data_0__17, ordered_img_data_0__16, 
                  ordered_img_data_0__15, ordered_img_data_0__14, 
                  ordered_img_data_0__13, ordered_img_data_0__12, 
                  ordered_img_data_0__11, ordered_img_data_0__10, 
                  ordered_img_data_0__9, ordered_img_data_0__8, 
                  ordered_img_data_0__7, ordered_img_data_0__6, 
                  ordered_img_data_0__5, ordered_img_data_0__4, 
                  ordered_img_data_0__3, ordered_img_data_0__2, 
                  ordered_img_data_0__1, ordered_img_data_0__0, 
                  ordered_img_data_1__31, ordered_img_data_1__30, 
                  ordered_img_data_1__29, ordered_img_data_1__28, 
                  ordered_img_data_1__27, ordered_img_data_1__26, 
                  ordered_img_data_1__25, ordered_img_data_1__24, 
                  ordered_img_data_1__23, ordered_img_data_1__22, 
                  ordered_img_data_1__21, ordered_img_data_1__20, 
                  ordered_img_data_1__19, ordered_img_data_1__18, 
                  ordered_img_data_1__17, ordered_img_data_1__16, 
                  ordered_img_data_1__15, ordered_img_data_1__14, 
                  ordered_img_data_1__13, ordered_img_data_1__12, 
                  ordered_img_data_1__11, ordered_img_data_1__10, 
                  ordered_img_data_1__9, ordered_img_data_1__8, 
                  ordered_img_data_1__7, ordered_img_data_1__6, 
                  ordered_img_data_1__5, ordered_img_data_1__4, 
                  ordered_img_data_1__3, ordered_img_data_1__2, 
                  ordered_img_data_1__1, ordered_img_data_1__0, 
                  ordered_img_data_2__31, ordered_img_data_2__30, 
                  ordered_img_data_2__29, ordered_img_data_2__28, 
                  ordered_img_data_2__27, ordered_img_data_2__26, 
                  ordered_img_data_2__25, ordered_img_data_2__24, 
                  ordered_img_data_2__23, ordered_img_data_2__22, 
                  ordered_img_data_2__21, ordered_img_data_2__20, 
                  ordered_img_data_2__19, ordered_img_data_2__18, 
                  ordered_img_data_2__17, ordered_img_data_2__16, 
                  ordered_img_data_2__15, ordered_img_data_2__14, 
                  ordered_img_data_2__13, ordered_img_data_2__12, 
                  ordered_img_data_2__11, ordered_img_data_2__10, 
                  ordered_img_data_2__9, ordered_img_data_2__8, 
                  ordered_img_data_2__7, ordered_img_data_2__6, 
                  ordered_img_data_2__5, ordered_img_data_2__4, 
                  ordered_img_data_2__3, ordered_img_data_2__2, 
                  ordered_img_data_2__1, ordered_img_data_2__0, 
                  ordered_img_data_3__31, ordered_img_data_3__30, 
                  ordered_img_data_3__29, ordered_img_data_3__28, 
                  ordered_img_data_3__27, ordered_img_data_3__26, 
                  ordered_img_data_3__25, ordered_img_data_3__24, 
                  ordered_img_data_3__23, ordered_img_data_3__22, 
                  ordered_img_data_3__21, ordered_img_data_3__20, 
                  ordered_img_data_3__19, ordered_img_data_3__18, 
                  ordered_img_data_3__17, ordered_img_data_3__16, 
                  ordered_img_data_3__15, ordered_img_data_3__14, 
                  ordered_img_data_3__13, ordered_img_data_3__12, 
                  ordered_img_data_3__11, ordered_img_data_3__10, 
                  ordered_img_data_3__9, ordered_img_data_3__8, 
                  ordered_img_data_3__7, ordered_img_data_3__6, 
                  ordered_img_data_3__5, ordered_img_data_3__4, 
                  ordered_img_data_3__3, ordered_img_data_3__2, 
                  ordered_img_data_3__1, ordered_img_data_3__0, 
                  ordered_img_data_4__31, ordered_img_data_4__30, 
                  ordered_img_data_4__29, ordered_img_data_4__28, 
                  ordered_img_data_4__27, ordered_img_data_4__26, 
                  ordered_img_data_4__25, ordered_img_data_4__24, 
                  ordered_img_data_4__23, ordered_img_data_4__22, 
                  ordered_img_data_4__21, ordered_img_data_4__20, 
                  ordered_img_data_4__19, ordered_img_data_4__18, 
                  ordered_img_data_4__17, ordered_img_data_4__16, 
                  ordered_img_data_4__15, ordered_img_data_4__14, 
                  ordered_img_data_4__13, ordered_img_data_4__12, 
                  ordered_img_data_4__11, ordered_img_data_4__10, 
                  ordered_img_data_4__9, ordered_img_data_4__8, 
                  ordered_img_data_4__7, ordered_img_data_4__6, 
                  ordered_img_data_4__5, ordered_img_data_4__4, 
                  ordered_img_data_4__3, ordered_img_data_4__2, 
                  ordered_img_data_4__1, ordered_img_data_4__0, 
                  ordered_img_data_5__31, ordered_img_data_5__30, 
                  ordered_img_data_5__29, ordered_img_data_5__28, 
                  ordered_img_data_5__27, ordered_img_data_5__26, 
                  ordered_img_data_5__25, ordered_img_data_5__24, 
                  ordered_img_data_5__23, ordered_img_data_5__22, 
                  ordered_img_data_5__21, ordered_img_data_5__20, 
                  ordered_img_data_5__19, ordered_img_data_5__18, 
                  ordered_img_data_5__17, ordered_img_data_5__16, 
                  ordered_img_data_5__15, ordered_img_data_5__14, 
                  ordered_img_data_5__13, ordered_img_data_5__12, 
                  ordered_img_data_5__11, ordered_img_data_5__10, 
                  ordered_img_data_5__9, ordered_img_data_5__8, 
                  ordered_img_data_5__7, ordered_img_data_5__6, 
                  ordered_img_data_5__5, ordered_img_data_5__4, 
                  ordered_img_data_5__3, ordered_img_data_5__2, 
                  ordered_img_data_5__1, ordered_img_data_5__0, 
                  ordered_img_data_6__31, ordered_img_data_6__30, 
                  ordered_img_data_6__29, ordered_img_data_6__28, 
                  ordered_img_data_6__27, ordered_img_data_6__26, 
                  ordered_img_data_6__25, ordered_img_data_6__24, 
                  ordered_img_data_6__23, ordered_img_data_6__22, 
                  ordered_img_data_6__21, ordered_img_data_6__20, 
                  ordered_img_data_6__19, ordered_img_data_6__18, 
                  ordered_img_data_6__17, ordered_img_data_6__16, 
                  ordered_img_data_6__15, ordered_img_data_6__14, 
                  ordered_img_data_6__13, ordered_img_data_6__12, 
                  ordered_img_data_6__11, ordered_img_data_6__10, 
                  ordered_img_data_6__9, ordered_img_data_6__8, 
                  ordered_img_data_6__7, ordered_img_data_6__6, 
                  ordered_img_data_6__5, ordered_img_data_6__4, 
                  ordered_img_data_6__3, ordered_img_data_6__2, 
                  ordered_img_data_6__1, ordered_img_data_6__0, 
                  ordered_img_data_7__31, ordered_img_data_7__30, 
                  ordered_img_data_7__29, ordered_img_data_7__28, 
                  ordered_img_data_7__27, ordered_img_data_7__26, 
                  ordered_img_data_7__25, ordered_img_data_7__24, 
                  ordered_img_data_7__23, ordered_img_data_7__22, 
                  ordered_img_data_7__21, ordered_img_data_7__20, 
                  ordered_img_data_7__19, ordered_img_data_7__18, 
                  ordered_img_data_7__17, ordered_img_data_7__16, 
                  ordered_img_data_7__15, ordered_img_data_7__14, 
                  ordered_img_data_7__13, ordered_img_data_7__12, 
                  ordered_img_data_7__11, ordered_img_data_7__10, 
                  ordered_img_data_7__9, ordered_img_data_7__8, 
                  ordered_img_data_7__7, ordered_img_data_7__6, 
                  ordered_img_data_7__5, ordered_img_data_7__4, 
                  ordered_img_data_7__3, ordered_img_data_7__2, 
                  ordered_img_data_7__1, ordered_img_data_7__0, 
                  ordered_img_data_8__31, ordered_img_data_8__30, 
                  ordered_img_data_8__29, ordered_img_data_8__28, 
                  ordered_img_data_8__27, ordered_img_data_8__26, 
                  ordered_img_data_8__25, ordered_img_data_8__24, 
                  ordered_img_data_8__23, ordered_img_data_8__22, 
                  ordered_img_data_8__21, ordered_img_data_8__20, 
                  ordered_img_data_8__19, ordered_img_data_8__18, 
                  ordered_img_data_8__17, ordered_img_data_8__16, 
                  ordered_img_data_8__15, ordered_img_data_8__14, 
                  ordered_img_data_8__13, ordered_img_data_8__12, 
                  ordered_img_data_8__11, ordered_img_data_8__10, 
                  ordered_img_data_8__9, ordered_img_data_8__8, 
                  ordered_img_data_8__7, ordered_img_data_8__6, 
                  ordered_img_data_8__5, ordered_img_data_8__4, 
                  ordered_img_data_8__3, ordered_img_data_8__2, 
                  ordered_img_data_8__1, ordered_img_data_8__0, 
                  ordered_img_data_9__31, ordered_img_data_9__30, 
                  ordered_img_data_9__29, ordered_img_data_9__28, 
                  ordered_img_data_9__27, ordered_img_data_9__26, 
                  ordered_img_data_9__25, ordered_img_data_9__24, 
                  ordered_img_data_9__23, ordered_img_data_9__22, 
                  ordered_img_data_9__21, ordered_img_data_9__20, 
                  ordered_img_data_9__19, ordered_img_data_9__18, 
                  ordered_img_data_9__17, ordered_img_data_9__16, 
                  ordered_img_data_9__15, ordered_img_data_9__14, 
                  ordered_img_data_9__13, ordered_img_data_9__12, 
                  ordered_img_data_9__11, ordered_img_data_9__10, 
                  ordered_img_data_9__9, ordered_img_data_9__8, 
                  ordered_img_data_9__7, ordered_img_data_9__6, 
                  ordered_img_data_9__5, ordered_img_data_9__4, 
                  ordered_img_data_9__3, ordered_img_data_9__2, 
                  ordered_img_data_9__1, ordered_img_data_9__0, 
                  ordered_img_data_10__31, ordered_img_data_10__30, 
                  ordered_img_data_10__29, ordered_img_data_10__28, 
                  ordered_img_data_10__27, ordered_img_data_10__26, 
                  ordered_img_data_10__25, ordered_img_data_10__24, 
                  ordered_img_data_10__23, ordered_img_data_10__22, 
                  ordered_img_data_10__21, ordered_img_data_10__20, 
                  ordered_img_data_10__19, ordered_img_data_10__18, 
                  ordered_img_data_10__17, ordered_img_data_10__16, 
                  ordered_img_data_10__15, ordered_img_data_10__14, 
                  ordered_img_data_10__13, ordered_img_data_10__12, 
                  ordered_img_data_10__11, ordered_img_data_10__10, 
                  ordered_img_data_10__9, ordered_img_data_10__8, 
                  ordered_img_data_10__7, ordered_img_data_10__6, 
                  ordered_img_data_10__5, ordered_img_data_10__4, 
                  ordered_img_data_10__3, ordered_img_data_10__2, 
                  ordered_img_data_10__1, ordered_img_data_10__0, 
                  ordered_img_data_11__31, ordered_img_data_11__30, 
                  ordered_img_data_11__29, ordered_img_data_11__28, 
                  ordered_img_data_11__27, ordered_img_data_11__26, 
                  ordered_img_data_11__25, ordered_img_data_11__24, 
                  ordered_img_data_11__23, ordered_img_data_11__22, 
                  ordered_img_data_11__21, ordered_img_data_11__20, 
                  ordered_img_data_11__19, ordered_img_data_11__18, 
                  ordered_img_data_11__17, ordered_img_data_11__16, 
                  ordered_img_data_11__15, ordered_img_data_11__14, 
                  ordered_img_data_11__13, ordered_img_data_11__12, 
                  ordered_img_data_11__11, ordered_img_data_11__10, 
                  ordered_img_data_11__9, ordered_img_data_11__8, 
                  ordered_img_data_11__7, ordered_img_data_11__6, 
                  ordered_img_data_11__5, ordered_img_data_11__4, 
                  ordered_img_data_11__3, ordered_img_data_11__2, 
                  ordered_img_data_11__1, ordered_img_data_11__0, 
                  ordered_img_data_12__31, ordered_img_data_12__30, 
                  ordered_img_data_12__29, ordered_img_data_12__28, 
                  ordered_img_data_12__27, ordered_img_data_12__26, 
                  ordered_img_data_12__25, ordered_img_data_12__24, 
                  ordered_img_data_12__23, ordered_img_data_12__22, 
                  ordered_img_data_12__21, ordered_img_data_12__20, 
                  ordered_img_data_12__19, ordered_img_data_12__18, 
                  ordered_img_data_12__17, ordered_img_data_12__16, 
                  ordered_img_data_12__15, ordered_img_data_12__14, 
                  ordered_img_data_12__13, ordered_img_data_12__12, 
                  ordered_img_data_12__11, ordered_img_data_12__10, 
                  ordered_img_data_12__9, ordered_img_data_12__8, 
                  ordered_img_data_12__7, ordered_img_data_12__6, 
                  ordered_img_data_12__5, ordered_img_data_12__4, 
                  ordered_img_data_12__3, ordered_img_data_12__2, 
                  ordered_img_data_12__1, ordered_img_data_12__0, 
                  ordered_img_data_13__31, ordered_img_data_13__30, 
                  ordered_img_data_13__29, ordered_img_data_13__28, 
                  ordered_img_data_13__27, ordered_img_data_13__26, 
                  ordered_img_data_13__25, ordered_img_data_13__24, 
                  ordered_img_data_13__23, ordered_img_data_13__22, 
                  ordered_img_data_13__21, ordered_img_data_13__20, 
                  ordered_img_data_13__19, ordered_img_data_13__18, 
                  ordered_img_data_13__17, ordered_img_data_13__16, 
                  ordered_img_data_13__15, ordered_img_data_13__14, 
                  ordered_img_data_13__13, ordered_img_data_13__12, 
                  ordered_img_data_13__11, ordered_img_data_13__10, 
                  ordered_img_data_13__9, ordered_img_data_13__8, 
                  ordered_img_data_13__7, ordered_img_data_13__6, 
                  ordered_img_data_13__5, ordered_img_data_13__4, 
                  ordered_img_data_13__3, ordered_img_data_13__2, 
                  ordered_img_data_13__1, ordered_img_data_13__0, 
                  ordered_img_data_14__31, ordered_img_data_14__30, 
                  ordered_img_data_14__29, ordered_img_data_14__28, 
                  ordered_img_data_14__27, ordered_img_data_14__26, 
                  ordered_img_data_14__25, ordered_img_data_14__24, 
                  ordered_img_data_14__23, ordered_img_data_14__22, 
                  ordered_img_data_14__21, ordered_img_data_14__20, 
                  ordered_img_data_14__19, ordered_img_data_14__18, 
                  ordered_img_data_14__17, ordered_img_data_14__16, 
                  ordered_img_data_14__15, ordered_img_data_14__14, 
                  ordered_img_data_14__13, ordered_img_data_14__12, 
                  ordered_img_data_14__11, ordered_img_data_14__10, 
                  ordered_img_data_14__9, ordered_img_data_14__8, 
                  ordered_img_data_14__7, ordered_img_data_14__6, 
                  ordered_img_data_14__5, ordered_img_data_14__4, 
                  ordered_img_data_14__3, ordered_img_data_14__2, 
                  ordered_img_data_14__1, ordered_img_data_14__0, 
                  ordered_img_data_15__31, ordered_img_data_15__30, 
                  ordered_img_data_15__29, ordered_img_data_15__28, 
                  ordered_img_data_15__27, ordered_img_data_15__26, 
                  ordered_img_data_15__25, ordered_img_data_15__24, 
                  ordered_img_data_15__23, ordered_img_data_15__22, 
                  ordered_img_data_15__21, ordered_img_data_15__20, 
                  ordered_img_data_15__19, ordered_img_data_15__18, 
                  ordered_img_data_15__17, ordered_img_data_15__16, 
                  ordered_img_data_15__15, ordered_img_data_15__14, 
                  ordered_img_data_15__13, ordered_img_data_15__12, 
                  ordered_img_data_15__11, ordered_img_data_15__10, 
                  ordered_img_data_15__9, ordered_img_data_15__8, 
                  ordered_img_data_15__7, ordered_img_data_15__6, 
                  ordered_img_data_15__5, ordered_img_data_15__4, 
                  ordered_img_data_15__3, ordered_img_data_15__2, 
                  ordered_img_data_15__1, ordered_img_data_15__0, 
                  ordered_img_data_16__31, ordered_img_data_16__30, 
                  ordered_img_data_16__29, ordered_img_data_16__28, 
                  ordered_img_data_16__27, ordered_img_data_16__26, 
                  ordered_img_data_16__25, ordered_img_data_16__24, 
                  ordered_img_data_16__23, ordered_img_data_16__22, 
                  ordered_img_data_16__21, ordered_img_data_16__20, 
                  ordered_img_data_16__19, ordered_img_data_16__18, 
                  ordered_img_data_16__17, ordered_img_data_16__16, 
                  ordered_img_data_16__15, ordered_img_data_16__14, 
                  ordered_img_data_16__13, ordered_img_data_16__12, 
                  ordered_img_data_16__11, ordered_img_data_16__10, 
                  ordered_img_data_16__9, ordered_img_data_16__8, 
                  ordered_img_data_16__7, ordered_img_data_16__6, 
                  ordered_img_data_16__5, ordered_img_data_16__4, 
                  ordered_img_data_16__3, ordered_img_data_16__2, 
                  ordered_img_data_16__1, ordered_img_data_16__0, 
                  ordered_img_data_17__31, ordered_img_data_17__30, 
                  ordered_img_data_17__29, ordered_img_data_17__28, 
                  ordered_img_data_17__27, ordered_img_data_17__26, 
                  ordered_img_data_17__25, ordered_img_data_17__24, 
                  ordered_img_data_17__23, ordered_img_data_17__22, 
                  ordered_img_data_17__21, ordered_img_data_17__20, 
                  ordered_img_data_17__19, ordered_img_data_17__18, 
                  ordered_img_data_17__17, ordered_img_data_17__16, 
                  ordered_img_data_17__15, ordered_img_data_17__14, 
                  ordered_img_data_17__13, ordered_img_data_17__12, 
                  ordered_img_data_17__11, ordered_img_data_17__10, 
                  ordered_img_data_17__9, ordered_img_data_17__8, 
                  ordered_img_data_17__7, ordered_img_data_17__6, 
                  ordered_img_data_17__5, ordered_img_data_17__4, 
                  ordered_img_data_17__3, ordered_img_data_17__2, 
                  ordered_img_data_17__1, ordered_img_data_17__0, 
                  ordered_img_data_18__31, ordered_img_data_18__30, 
                  ordered_img_data_18__29, ordered_img_data_18__28, 
                  ordered_img_data_18__27, ordered_img_data_18__26, 
                  ordered_img_data_18__25, ordered_img_data_18__24, 
                  ordered_img_data_18__23, ordered_img_data_18__22, 
                  ordered_img_data_18__21, ordered_img_data_18__20, 
                  ordered_img_data_18__19, ordered_img_data_18__18, 
                  ordered_img_data_18__17, ordered_img_data_18__16, 
                  ordered_img_data_18__15, ordered_img_data_18__14, 
                  ordered_img_data_18__13, ordered_img_data_18__12, 
                  ordered_img_data_18__11, ordered_img_data_18__10, 
                  ordered_img_data_18__9, ordered_img_data_18__8, 
                  ordered_img_data_18__7, ordered_img_data_18__6, 
                  ordered_img_data_18__5, ordered_img_data_18__4, 
                  ordered_img_data_18__3, ordered_img_data_18__2, 
                  ordered_img_data_18__1, ordered_img_data_18__0, 
                  ordered_img_data_19__31, ordered_img_data_19__30, 
                  ordered_img_data_19__29, ordered_img_data_19__28, 
                  ordered_img_data_19__27, ordered_img_data_19__26, 
                  ordered_img_data_19__25, ordered_img_data_19__24, 
                  ordered_img_data_19__23, ordered_img_data_19__22, 
                  ordered_img_data_19__21, ordered_img_data_19__20, 
                  ordered_img_data_19__19, ordered_img_data_19__18, 
                  ordered_img_data_19__17, ordered_img_data_19__16, 
                  ordered_img_data_19__15, ordered_img_data_19__14, 
                  ordered_img_data_19__13, ordered_img_data_19__12, 
                  ordered_img_data_19__11, ordered_img_data_19__10, 
                  ordered_img_data_19__9, ordered_img_data_19__8, 
                  ordered_img_data_19__7, ordered_img_data_19__6, 
                  ordered_img_data_19__5, ordered_img_data_19__4, 
                  ordered_img_data_19__3, ordered_img_data_19__2, 
                  ordered_img_data_19__1, ordered_img_data_19__0, 
                  ordered_img_data_20__31, ordered_img_data_20__30, 
                  ordered_img_data_20__29, ordered_img_data_20__28, 
                  ordered_img_data_20__27, ordered_img_data_20__26, 
                  ordered_img_data_20__25, ordered_img_data_20__24, 
                  ordered_img_data_20__23, ordered_img_data_20__22, 
                  ordered_img_data_20__21, ordered_img_data_20__20, 
                  ordered_img_data_20__19, ordered_img_data_20__18, 
                  ordered_img_data_20__17, ordered_img_data_20__16, 
                  ordered_img_data_20__15, ordered_img_data_20__14, 
                  ordered_img_data_20__13, ordered_img_data_20__12, 
                  ordered_img_data_20__11, ordered_img_data_20__10, 
                  ordered_img_data_20__9, ordered_img_data_20__8, 
                  ordered_img_data_20__7, ordered_img_data_20__6, 
                  ordered_img_data_20__5, ordered_img_data_20__4, 
                  ordered_img_data_20__3, ordered_img_data_20__2, 
                  ordered_img_data_20__1, ordered_img_data_20__0, 
                  ordered_img_data_21__31, ordered_img_data_21__30, 
                  ordered_img_data_21__29, ordered_img_data_21__28, 
                  ordered_img_data_21__27, ordered_img_data_21__26, 
                  ordered_img_data_21__25, ordered_img_data_21__24, 
                  ordered_img_data_21__23, ordered_img_data_21__22, 
                  ordered_img_data_21__21, ordered_img_data_21__20, 
                  ordered_img_data_21__19, ordered_img_data_21__18, 
                  ordered_img_data_21__17, ordered_img_data_21__16, 
                  ordered_img_data_21__15, ordered_img_data_21__14, 
                  ordered_img_data_21__13, ordered_img_data_21__12, 
                  ordered_img_data_21__11, ordered_img_data_21__10, 
                  ordered_img_data_21__9, ordered_img_data_21__8, 
                  ordered_img_data_21__7, ordered_img_data_21__6, 
                  ordered_img_data_21__5, ordered_img_data_21__4, 
                  ordered_img_data_21__3, ordered_img_data_21__2, 
                  ordered_img_data_21__1, ordered_img_data_21__0, 
                  ordered_img_data_22__31, ordered_img_data_22__30, 
                  ordered_img_data_22__29, ordered_img_data_22__28, 
                  ordered_img_data_22__27, ordered_img_data_22__26, 
                  ordered_img_data_22__25, ordered_img_data_22__24, 
                  ordered_img_data_22__23, ordered_img_data_22__22, 
                  ordered_img_data_22__21, ordered_img_data_22__20, 
                  ordered_img_data_22__19, ordered_img_data_22__18, 
                  ordered_img_data_22__17, ordered_img_data_22__16, 
                  ordered_img_data_22__15, ordered_img_data_22__14, 
                  ordered_img_data_22__13, ordered_img_data_22__12, 
                  ordered_img_data_22__11, ordered_img_data_22__10, 
                  ordered_img_data_22__9, ordered_img_data_22__8, 
                  ordered_img_data_22__7, ordered_img_data_22__6, 
                  ordered_img_data_22__5, ordered_img_data_22__4, 
                  ordered_img_data_22__3, ordered_img_data_22__2, 
                  ordered_img_data_22__1, ordered_img_data_22__0, 
                  ordered_img_data_23__31, ordered_img_data_23__30, 
                  ordered_img_data_23__29, ordered_img_data_23__28, 
                  ordered_img_data_23__27, ordered_img_data_23__26, 
                  ordered_img_data_23__25, ordered_img_data_23__24, 
                  ordered_img_data_23__23, ordered_img_data_23__22, 
                  ordered_img_data_23__21, ordered_img_data_23__20, 
                  ordered_img_data_23__19, ordered_img_data_23__18, 
                  ordered_img_data_23__17, ordered_img_data_23__16, 
                  ordered_img_data_23__15, ordered_img_data_23__14, 
                  ordered_img_data_23__13, ordered_img_data_23__12, 
                  ordered_img_data_23__11, ordered_img_data_23__10, 
                  ordered_img_data_23__9, ordered_img_data_23__8, 
                  ordered_img_data_23__7, ordered_img_data_23__6, 
                  ordered_img_data_23__5, ordered_img_data_23__4, 
                  ordered_img_data_23__3, ordered_img_data_23__2, 
                  ordered_img_data_23__1, ordered_img_data_23__0, 
                  ordered_img_data_24__31, ordered_img_data_24__30, 
                  ordered_img_data_24__29, ordered_img_data_24__28, 
                  ordered_img_data_24__27, ordered_img_data_24__26, 
                  ordered_img_data_24__25, ordered_img_data_24__24, 
                  ordered_img_data_24__23, ordered_img_data_24__22, 
                  ordered_img_data_24__21, ordered_img_data_24__20, 
                  ordered_img_data_24__19, ordered_img_data_24__18, 
                  ordered_img_data_24__17, ordered_img_data_24__16, 
                  ordered_img_data_24__15, ordered_img_data_24__14, 
                  ordered_img_data_24__13, ordered_img_data_24__12, 
                  ordered_img_data_24__11, ordered_img_data_24__10, 
                  ordered_img_data_24__9, ordered_img_data_24__8, 
                  ordered_img_data_24__7, ordered_img_data_24__6, 
                  ordered_img_data_24__5, ordered_img_data_24__4, 
                  ordered_img_data_24__3, ordered_img_data_24__2, 
                  ordered_img_data_24__1, ordered_img_data_24__0, 
                  ordered_filter_data_0__31, ordered_filter_data_0__30, 
                  ordered_filter_data_0__29, ordered_filter_data_0__28, 
                  ordered_filter_data_0__27, ordered_filter_data_0__26, 
                  ordered_filter_data_0__25, ordered_filter_data_0__24, 
                  ordered_filter_data_0__23, ordered_filter_data_0__22, 
                  ordered_filter_data_0__21, ordered_filter_data_0__20, 
                  ordered_filter_data_0__19, ordered_filter_data_0__18, 
                  ordered_filter_data_0__17, ordered_filter_data_0__16, 
                  ordered_filter_data_0__15, ordered_filter_data_0__14, 
                  ordered_filter_data_0__13, ordered_filter_data_0__12, 
                  ordered_filter_data_0__11, ordered_filter_data_0__10, 
                  ordered_filter_data_0__9, ordered_filter_data_0__8, 
                  ordered_filter_data_0__7, ordered_filter_data_0__6, 
                  ordered_filter_data_0__5, ordered_filter_data_0__4, 
                  ordered_filter_data_0__3, ordered_filter_data_0__2, 
                  ordered_filter_data_0__1, ordered_filter_data_0__0, 
                  ordered_filter_data_1__31, ordered_filter_data_1__30, 
                  ordered_filter_data_1__29, ordered_filter_data_1__28, 
                  ordered_filter_data_1__27, ordered_filter_data_1__26, 
                  ordered_filter_data_1__25, ordered_filter_data_1__24, 
                  ordered_filter_data_1__23, ordered_filter_data_1__22, 
                  ordered_filter_data_1__21, ordered_filter_data_1__20, 
                  ordered_filter_data_1__19, ordered_filter_data_1__18, 
                  ordered_filter_data_1__17, ordered_filter_data_1__16, 
                  ordered_filter_data_1__15, ordered_filter_data_1__14, 
                  ordered_filter_data_1__13, ordered_filter_data_1__12, 
                  ordered_filter_data_1__11, ordered_filter_data_1__10, 
                  ordered_filter_data_1__9, ordered_filter_data_1__8, 
                  ordered_filter_data_1__7, ordered_filter_data_1__6, 
                  ordered_filter_data_1__5, ordered_filter_data_1__4, 
                  ordered_filter_data_1__3, ordered_filter_data_1__2, 
                  ordered_filter_data_1__1, ordered_filter_data_1__0, 
                  ordered_filter_data_2__31, ordered_filter_data_2__30, 
                  ordered_filter_data_2__29, ordered_filter_data_2__28, 
                  ordered_filter_data_2__27, ordered_filter_data_2__26, 
                  ordered_filter_data_2__25, ordered_filter_data_2__24, 
                  ordered_filter_data_2__23, ordered_filter_data_2__22, 
                  ordered_filter_data_2__21, ordered_filter_data_2__20, 
                  ordered_filter_data_2__19, ordered_filter_data_2__18, 
                  ordered_filter_data_2__17, ordered_filter_data_2__16, 
                  ordered_filter_data_2__15, ordered_filter_data_2__14, 
                  ordered_filter_data_2__13, ordered_filter_data_2__12, 
                  ordered_filter_data_2__11, ordered_filter_data_2__10, 
                  ordered_filter_data_2__9, ordered_filter_data_2__8, 
                  ordered_filter_data_2__7, ordered_filter_data_2__6, 
                  ordered_filter_data_2__5, ordered_filter_data_2__4, 
                  ordered_filter_data_2__3, ordered_filter_data_2__2, 
                  ordered_filter_data_2__1, ordered_filter_data_2__0, 
                  ordered_filter_data_3__31, ordered_filter_data_3__30, 
                  ordered_filter_data_3__29, ordered_filter_data_3__28, 
                  ordered_filter_data_3__27, ordered_filter_data_3__26, 
                  ordered_filter_data_3__25, ordered_filter_data_3__24, 
                  ordered_filter_data_3__23, ordered_filter_data_3__22, 
                  ordered_filter_data_3__21, ordered_filter_data_3__20, 
                  ordered_filter_data_3__19, ordered_filter_data_3__18, 
                  ordered_filter_data_3__17, ordered_filter_data_3__16, 
                  ordered_filter_data_3__15, ordered_filter_data_3__14, 
                  ordered_filter_data_3__13, ordered_filter_data_3__12, 
                  ordered_filter_data_3__11, ordered_filter_data_3__10, 
                  ordered_filter_data_3__9, ordered_filter_data_3__8, 
                  ordered_filter_data_3__7, ordered_filter_data_3__6, 
                  ordered_filter_data_3__5, ordered_filter_data_3__4, 
                  ordered_filter_data_3__3, ordered_filter_data_3__2, 
                  ordered_filter_data_3__1, ordered_filter_data_3__0, 
                  ordered_filter_data_4__31, ordered_filter_data_4__30, 
                  ordered_filter_data_4__29, ordered_filter_data_4__28, 
                  ordered_filter_data_4__27, ordered_filter_data_4__26, 
                  ordered_filter_data_4__25, ordered_filter_data_4__24, 
                  ordered_filter_data_4__23, ordered_filter_data_4__22, 
                  ordered_filter_data_4__21, ordered_filter_data_4__20, 
                  ordered_filter_data_4__19, ordered_filter_data_4__18, 
                  ordered_filter_data_4__17, ordered_filter_data_4__16, 
                  ordered_filter_data_4__15, ordered_filter_data_4__14, 
                  ordered_filter_data_4__13, ordered_filter_data_4__12, 
                  ordered_filter_data_4__11, ordered_filter_data_4__10, 
                  ordered_filter_data_4__9, ordered_filter_data_4__8, 
                  ordered_filter_data_4__7, ordered_filter_data_4__6, 
                  ordered_filter_data_4__5, ordered_filter_data_4__4, 
                  ordered_filter_data_4__3, ordered_filter_data_4__2, 
                  ordered_filter_data_4__1, ordered_filter_data_4__0, 
                  ordered_filter_data_5__31, ordered_filter_data_5__30, 
                  ordered_filter_data_5__29, ordered_filter_data_5__28, 
                  ordered_filter_data_5__27, ordered_filter_data_5__26, 
                  ordered_filter_data_5__25, ordered_filter_data_5__24, 
                  ordered_filter_data_5__23, ordered_filter_data_5__22, 
                  ordered_filter_data_5__21, ordered_filter_data_5__20, 
                  ordered_filter_data_5__19, ordered_filter_data_5__18, 
                  ordered_filter_data_5__17, ordered_filter_data_5__16, 
                  ordered_filter_data_5__15, ordered_filter_data_5__14, 
                  ordered_filter_data_5__13, ordered_filter_data_5__12, 
                  ordered_filter_data_5__11, ordered_filter_data_5__10, 
                  ordered_filter_data_5__9, ordered_filter_data_5__8, 
                  ordered_filter_data_5__7, ordered_filter_data_5__6, 
                  ordered_filter_data_5__5, ordered_filter_data_5__4, 
                  ordered_filter_data_5__3, ordered_filter_data_5__2, 
                  ordered_filter_data_5__1, ordered_filter_data_5__0, 
                  ordered_filter_data_6__31, ordered_filter_data_6__30, 
                  ordered_filter_data_6__29, ordered_filter_data_6__28, 
                  ordered_filter_data_6__27, ordered_filter_data_6__26, 
                  ordered_filter_data_6__25, ordered_filter_data_6__24, 
                  ordered_filter_data_6__23, ordered_filter_data_6__22, 
                  ordered_filter_data_6__21, ordered_filter_data_6__20, 
                  ordered_filter_data_6__19, ordered_filter_data_6__18, 
                  ordered_filter_data_6__17, ordered_filter_data_6__16, 
                  ordered_filter_data_6__15, ordered_filter_data_6__14, 
                  ordered_filter_data_6__13, ordered_filter_data_6__12, 
                  ordered_filter_data_6__11, ordered_filter_data_6__10, 
                  ordered_filter_data_6__9, ordered_filter_data_6__8, 
                  ordered_filter_data_6__7, ordered_filter_data_6__6, 
                  ordered_filter_data_6__5, ordered_filter_data_6__4, 
                  ordered_filter_data_6__3, ordered_filter_data_6__2, 
                  ordered_filter_data_6__1, ordered_filter_data_6__0, 
                  ordered_filter_data_7__31, ordered_filter_data_7__30, 
                  ordered_filter_data_7__29, ordered_filter_data_7__28, 
                  ordered_filter_data_7__27, ordered_filter_data_7__26, 
                  ordered_filter_data_7__25, ordered_filter_data_7__24, 
                  ordered_filter_data_7__23, ordered_filter_data_7__22, 
                  ordered_filter_data_7__21, ordered_filter_data_7__20, 
                  ordered_filter_data_7__19, ordered_filter_data_7__18, 
                  ordered_filter_data_7__17, ordered_filter_data_7__16, 
                  ordered_filter_data_7__15, ordered_filter_data_7__14, 
                  ordered_filter_data_7__13, ordered_filter_data_7__12, 
                  ordered_filter_data_7__11, ordered_filter_data_7__10, 
                  ordered_filter_data_7__9, ordered_filter_data_7__8, 
                  ordered_filter_data_7__7, ordered_filter_data_7__6, 
                  ordered_filter_data_7__5, ordered_filter_data_7__4, 
                  ordered_filter_data_7__3, ordered_filter_data_7__2, 
                  ordered_filter_data_7__1, ordered_filter_data_7__0, 
                  ordered_filter_data_8__31, ordered_filter_data_8__30, 
                  ordered_filter_data_8__29, ordered_filter_data_8__28, 
                  ordered_filter_data_8__27, ordered_filter_data_8__26, 
                  ordered_filter_data_8__25, ordered_filter_data_8__24, 
                  ordered_filter_data_8__23, ordered_filter_data_8__22, 
                  ordered_filter_data_8__21, ordered_filter_data_8__20, 
                  ordered_filter_data_8__19, ordered_filter_data_8__18, 
                  ordered_filter_data_8__17, ordered_filter_data_8__16, 
                  ordered_filter_data_8__15, ordered_filter_data_8__14, 
                  ordered_filter_data_8__13, ordered_filter_data_8__12, 
                  ordered_filter_data_8__11, ordered_filter_data_8__10, 
                  ordered_filter_data_8__9, ordered_filter_data_8__8, 
                  ordered_filter_data_8__7, ordered_filter_data_8__6, 
                  ordered_filter_data_8__5, ordered_filter_data_8__4, 
                  ordered_filter_data_8__3, ordered_filter_data_8__2, 
                  ordered_filter_data_8__1, ordered_filter_data_8__0, 
                  ordered_filter_data_9__31, ordered_filter_data_9__30, 
                  ordered_filter_data_9__29, ordered_filter_data_9__28, 
                  ordered_filter_data_9__27, ordered_filter_data_9__26, 
                  ordered_filter_data_9__25, ordered_filter_data_9__24, 
                  ordered_filter_data_9__23, ordered_filter_data_9__22, 
                  ordered_filter_data_9__21, ordered_filter_data_9__20, 
                  ordered_filter_data_9__19, ordered_filter_data_9__18, 
                  ordered_filter_data_9__17, ordered_filter_data_9__16, 
                  ordered_filter_data_9__15, ordered_filter_data_9__14, 
                  ordered_filter_data_9__13, ordered_filter_data_9__12, 
                  ordered_filter_data_9__11, ordered_filter_data_9__10, 
                  ordered_filter_data_9__9, ordered_filter_data_9__8, 
                  ordered_filter_data_9__7, ordered_filter_data_9__6, 
                  ordered_filter_data_9__5, ordered_filter_data_9__4, 
                  ordered_filter_data_9__3, ordered_filter_data_9__2, 
                  ordered_filter_data_9__1, ordered_filter_data_9__0, 
                  ordered_filter_data_10__31, ordered_filter_data_10__30, 
                  ordered_filter_data_10__29, ordered_filter_data_10__28, 
                  ordered_filter_data_10__27, ordered_filter_data_10__26, 
                  ordered_filter_data_10__25, ordered_filter_data_10__24, 
                  ordered_filter_data_10__23, ordered_filter_data_10__22, 
                  ordered_filter_data_10__21, ordered_filter_data_10__20, 
                  ordered_filter_data_10__19, ordered_filter_data_10__18, 
                  ordered_filter_data_10__17, ordered_filter_data_10__16, 
                  ordered_filter_data_10__15, ordered_filter_data_10__14, 
                  ordered_filter_data_10__13, ordered_filter_data_10__12, 
                  ordered_filter_data_10__11, ordered_filter_data_10__10, 
                  ordered_filter_data_10__9, ordered_filter_data_10__8, 
                  ordered_filter_data_10__7, ordered_filter_data_10__6, 
                  ordered_filter_data_10__5, ordered_filter_data_10__4, 
                  ordered_filter_data_10__3, ordered_filter_data_10__2, 
                  ordered_filter_data_10__1, ordered_filter_data_10__0, 
                  ordered_filter_data_11__31, ordered_filter_data_11__30, 
                  ordered_filter_data_11__29, ordered_filter_data_11__28, 
                  ordered_filter_data_11__27, ordered_filter_data_11__26, 
                  ordered_filter_data_11__25, ordered_filter_data_11__24, 
                  ordered_filter_data_11__23, ordered_filter_data_11__22, 
                  ordered_filter_data_11__21, ordered_filter_data_11__20, 
                  ordered_filter_data_11__19, ordered_filter_data_11__18, 
                  ordered_filter_data_11__17, ordered_filter_data_11__16, 
                  ordered_filter_data_11__15, ordered_filter_data_11__14, 
                  ordered_filter_data_11__13, ordered_filter_data_11__12, 
                  ordered_filter_data_11__11, ordered_filter_data_11__10, 
                  ordered_filter_data_11__9, ordered_filter_data_11__8, 
                  ordered_filter_data_11__7, ordered_filter_data_11__6, 
                  ordered_filter_data_11__5, ordered_filter_data_11__4, 
                  ordered_filter_data_11__3, ordered_filter_data_11__2, 
                  ordered_filter_data_11__1, ordered_filter_data_11__0, 
                  ordered_filter_data_12__31, ordered_filter_data_12__30, 
                  ordered_filter_data_12__29, ordered_filter_data_12__28, 
                  ordered_filter_data_12__27, ordered_filter_data_12__26, 
                  ordered_filter_data_12__25, ordered_filter_data_12__24, 
                  ordered_filter_data_12__23, ordered_filter_data_12__22, 
                  ordered_filter_data_12__21, ordered_filter_data_12__20, 
                  ordered_filter_data_12__19, ordered_filter_data_12__18, 
                  ordered_filter_data_12__17, ordered_filter_data_12__16, 
                  ordered_filter_data_12__15, ordered_filter_data_12__14, 
                  ordered_filter_data_12__13, ordered_filter_data_12__12, 
                  ordered_filter_data_12__11, ordered_filter_data_12__10, 
                  ordered_filter_data_12__9, ordered_filter_data_12__8, 
                  ordered_filter_data_12__7, ordered_filter_data_12__6, 
                  ordered_filter_data_12__5, ordered_filter_data_12__4, 
                  ordered_filter_data_12__3, ordered_filter_data_12__2, 
                  ordered_filter_data_12__1, ordered_filter_data_12__0, 
                  ordered_filter_data_13__31, ordered_filter_data_13__30, 
                  ordered_filter_data_13__29, ordered_filter_data_13__28, 
                  ordered_filter_data_13__27, ordered_filter_data_13__26, 
                  ordered_filter_data_13__25, ordered_filter_data_13__24, 
                  ordered_filter_data_13__23, ordered_filter_data_13__22, 
                  ordered_filter_data_13__21, ordered_filter_data_13__20, 
                  ordered_filter_data_13__19, ordered_filter_data_13__18, 
                  ordered_filter_data_13__17, ordered_filter_data_13__16, 
                  ordered_filter_data_13__15, ordered_filter_data_13__14, 
                  ordered_filter_data_13__13, ordered_filter_data_13__12, 
                  ordered_filter_data_13__11, ordered_filter_data_13__10, 
                  ordered_filter_data_13__9, ordered_filter_data_13__8, 
                  ordered_filter_data_13__7, ordered_filter_data_13__6, 
                  ordered_filter_data_13__5, ordered_filter_data_13__4, 
                  ordered_filter_data_13__3, ordered_filter_data_13__2, 
                  ordered_filter_data_13__1, ordered_filter_data_13__0, 
                  ordered_filter_data_14__31, ordered_filter_data_14__30, 
                  ordered_filter_data_14__29, ordered_filter_data_14__28, 
                  ordered_filter_data_14__27, ordered_filter_data_14__26, 
                  ordered_filter_data_14__25, ordered_filter_data_14__24, 
                  ordered_filter_data_14__23, ordered_filter_data_14__22, 
                  ordered_filter_data_14__21, ordered_filter_data_14__20, 
                  ordered_filter_data_14__19, ordered_filter_data_14__18, 
                  ordered_filter_data_14__17, ordered_filter_data_14__16, 
                  ordered_filter_data_14__15, ordered_filter_data_14__14, 
                  ordered_filter_data_14__13, ordered_filter_data_14__12, 
                  ordered_filter_data_14__11, ordered_filter_data_14__10, 
                  ordered_filter_data_14__9, ordered_filter_data_14__8, 
                  ordered_filter_data_14__7, ordered_filter_data_14__6, 
                  ordered_filter_data_14__5, ordered_filter_data_14__4, 
                  ordered_filter_data_14__3, ordered_filter_data_14__2, 
                  ordered_filter_data_14__1, ordered_filter_data_14__0, 
                  ordered_filter_data_15__31, ordered_filter_data_15__30, 
                  ordered_filter_data_15__29, ordered_filter_data_15__28, 
                  ordered_filter_data_15__27, ordered_filter_data_15__26, 
                  ordered_filter_data_15__25, ordered_filter_data_15__24, 
                  ordered_filter_data_15__23, ordered_filter_data_15__22, 
                  ordered_filter_data_15__21, ordered_filter_data_15__20, 
                  ordered_filter_data_15__19, ordered_filter_data_15__18, 
                  ordered_filter_data_15__17, ordered_filter_data_15__16, 
                  ordered_filter_data_15__15, ordered_filter_data_15__14, 
                  ordered_filter_data_15__13, ordered_filter_data_15__12, 
                  ordered_filter_data_15__11, ordered_filter_data_15__10, 
                  ordered_filter_data_15__9, ordered_filter_data_15__8, 
                  ordered_filter_data_15__7, ordered_filter_data_15__6, 
                  ordered_filter_data_15__5, ordered_filter_data_15__4, 
                  ordered_filter_data_15__3, ordered_filter_data_15__2, 
                  ordered_filter_data_15__1, ordered_filter_data_15__0, 
                  ordered_filter_data_16__31, ordered_filter_data_16__30, 
                  ordered_filter_data_16__29, ordered_filter_data_16__28, 
                  ordered_filter_data_16__27, ordered_filter_data_16__26, 
                  ordered_filter_data_16__25, ordered_filter_data_16__24, 
                  ordered_filter_data_16__23, ordered_filter_data_16__22, 
                  ordered_filter_data_16__21, ordered_filter_data_16__20, 
                  ordered_filter_data_16__19, ordered_filter_data_16__18, 
                  ordered_filter_data_16__17, ordered_filter_data_16__16, 
                  ordered_filter_data_16__15, ordered_filter_data_16__14, 
                  ordered_filter_data_16__13, ordered_filter_data_16__12, 
                  ordered_filter_data_16__11, ordered_filter_data_16__10, 
                  ordered_filter_data_16__9, ordered_filter_data_16__8, 
                  ordered_filter_data_16__7, ordered_filter_data_16__6, 
                  ordered_filter_data_16__5, ordered_filter_data_16__4, 
                  ordered_filter_data_16__3, ordered_filter_data_16__2, 
                  ordered_filter_data_16__1, ordered_filter_data_16__0, 
                  ordered_filter_data_17__31, ordered_filter_data_17__30, 
                  ordered_filter_data_17__29, ordered_filter_data_17__28, 
                  ordered_filter_data_17__27, ordered_filter_data_17__26, 
                  ordered_filter_data_17__25, ordered_filter_data_17__24, 
                  ordered_filter_data_17__23, ordered_filter_data_17__22, 
                  ordered_filter_data_17__21, ordered_filter_data_17__20, 
                  ordered_filter_data_17__19, ordered_filter_data_17__18, 
                  ordered_filter_data_17__17, ordered_filter_data_17__16, 
                  ordered_filter_data_17__15, ordered_filter_data_17__14, 
                  ordered_filter_data_17__13, ordered_filter_data_17__12, 
                  ordered_filter_data_17__11, ordered_filter_data_17__10, 
                  ordered_filter_data_17__9, ordered_filter_data_17__8, 
                  ordered_filter_data_17__7, ordered_filter_data_17__6, 
                  ordered_filter_data_17__5, ordered_filter_data_17__4, 
                  ordered_filter_data_17__3, ordered_filter_data_17__2, 
                  ordered_filter_data_17__1, ordered_filter_data_17__0, 
                  ordered_filter_data_18__31, ordered_filter_data_18__30, 
                  ordered_filter_data_18__29, ordered_filter_data_18__28, 
                  ordered_filter_data_18__27, ordered_filter_data_18__26, 
                  ordered_filter_data_18__25, ordered_filter_data_18__24, 
                  ordered_filter_data_18__23, ordered_filter_data_18__22, 
                  ordered_filter_data_18__21, ordered_filter_data_18__20, 
                  ordered_filter_data_18__19, ordered_filter_data_18__18, 
                  ordered_filter_data_18__17, ordered_filter_data_18__16, 
                  ordered_filter_data_18__15, ordered_filter_data_18__14, 
                  ordered_filter_data_18__13, ordered_filter_data_18__12, 
                  ordered_filter_data_18__11, ordered_filter_data_18__10, 
                  ordered_filter_data_18__9, ordered_filter_data_18__8, 
                  ordered_filter_data_18__7, ordered_filter_data_18__6, 
                  ordered_filter_data_18__5, ordered_filter_data_18__4, 
                  ordered_filter_data_18__3, ordered_filter_data_18__2, 
                  ordered_filter_data_18__1, ordered_filter_data_18__0, 
                  ordered_filter_data_19__31, ordered_filter_data_19__30, 
                  ordered_filter_data_19__29, ordered_filter_data_19__28, 
                  ordered_filter_data_19__27, ordered_filter_data_19__26, 
                  ordered_filter_data_19__25, ordered_filter_data_19__24, 
                  ordered_filter_data_19__23, ordered_filter_data_19__22, 
                  ordered_filter_data_19__21, ordered_filter_data_19__20, 
                  ordered_filter_data_19__19, ordered_filter_data_19__18, 
                  ordered_filter_data_19__17, ordered_filter_data_19__16, 
                  ordered_filter_data_19__15, ordered_filter_data_19__14, 
                  ordered_filter_data_19__13, ordered_filter_data_19__12, 
                  ordered_filter_data_19__11, ordered_filter_data_19__10, 
                  ordered_filter_data_19__9, ordered_filter_data_19__8, 
                  ordered_filter_data_19__7, ordered_filter_data_19__6, 
                  ordered_filter_data_19__5, ordered_filter_data_19__4, 
                  ordered_filter_data_19__3, ordered_filter_data_19__2, 
                  ordered_filter_data_19__1, ordered_filter_data_19__0, 
                  ordered_filter_data_20__31, ordered_filter_data_20__30, 
                  ordered_filter_data_20__29, ordered_filter_data_20__28, 
                  ordered_filter_data_20__27, ordered_filter_data_20__26, 
                  ordered_filter_data_20__25, ordered_filter_data_20__24, 
                  ordered_filter_data_20__23, ordered_filter_data_20__22, 
                  ordered_filter_data_20__21, ordered_filter_data_20__20, 
                  ordered_filter_data_20__19, ordered_filter_data_20__18, 
                  ordered_filter_data_20__17, ordered_filter_data_20__16, 
                  ordered_filter_data_20__15, ordered_filter_data_20__14, 
                  ordered_filter_data_20__13, ordered_filter_data_20__12, 
                  ordered_filter_data_20__11, ordered_filter_data_20__10, 
                  ordered_filter_data_20__9, ordered_filter_data_20__8, 
                  ordered_filter_data_20__7, ordered_filter_data_20__6, 
                  ordered_filter_data_20__5, ordered_filter_data_20__4, 
                  ordered_filter_data_20__3, ordered_filter_data_20__2, 
                  ordered_filter_data_20__1, ordered_filter_data_20__0, 
                  ordered_filter_data_21__31, ordered_filter_data_21__30, 
                  ordered_filter_data_21__29, ordered_filter_data_21__28, 
                  ordered_filter_data_21__27, ordered_filter_data_21__26, 
                  ordered_filter_data_21__25, ordered_filter_data_21__24, 
                  ordered_filter_data_21__23, ordered_filter_data_21__22, 
                  ordered_filter_data_21__21, ordered_filter_data_21__20, 
                  ordered_filter_data_21__19, ordered_filter_data_21__18, 
                  ordered_filter_data_21__17, ordered_filter_data_21__16, 
                  ordered_filter_data_21__15, ordered_filter_data_21__14, 
                  ordered_filter_data_21__13, ordered_filter_data_21__12, 
                  ordered_filter_data_21__11, ordered_filter_data_21__10, 
                  ordered_filter_data_21__9, ordered_filter_data_21__8, 
                  ordered_filter_data_21__7, ordered_filter_data_21__6, 
                  ordered_filter_data_21__5, ordered_filter_data_21__4, 
                  ordered_filter_data_21__3, ordered_filter_data_21__2, 
                  ordered_filter_data_21__1, ordered_filter_data_21__0, 
                  ordered_filter_data_22__31, ordered_filter_data_22__30, 
                  ordered_filter_data_22__29, ordered_filter_data_22__28, 
                  ordered_filter_data_22__27, ordered_filter_data_22__26, 
                  ordered_filter_data_22__25, ordered_filter_data_22__24, 
                  ordered_filter_data_22__23, ordered_filter_data_22__22, 
                  ordered_filter_data_22__21, ordered_filter_data_22__20, 
                  ordered_filter_data_22__19, ordered_filter_data_22__18, 
                  ordered_filter_data_22__17, ordered_filter_data_22__16, 
                  ordered_filter_data_22__15, ordered_filter_data_22__14, 
                  ordered_filter_data_22__13, ordered_filter_data_22__12, 
                  ordered_filter_data_22__11, ordered_filter_data_22__10, 
                  ordered_filter_data_22__9, ordered_filter_data_22__8, 
                  ordered_filter_data_22__7, ordered_filter_data_22__6, 
                  ordered_filter_data_22__5, ordered_filter_data_22__4, 
                  ordered_filter_data_22__3, ordered_filter_data_22__2, 
                  ordered_filter_data_22__1, ordered_filter_data_22__0, 
                  ordered_filter_data_23__31, ordered_filter_data_23__30, 
                  ordered_filter_data_23__29, ordered_filter_data_23__28, 
                  ordered_filter_data_23__27, ordered_filter_data_23__26, 
                  ordered_filter_data_23__25, ordered_filter_data_23__24, 
                  ordered_filter_data_23__23, ordered_filter_data_23__22, 
                  ordered_filter_data_23__21, ordered_filter_data_23__20, 
                  ordered_filter_data_23__19, ordered_filter_data_23__18, 
                  ordered_filter_data_23__17, ordered_filter_data_23__16, 
                  ordered_filter_data_23__15, ordered_filter_data_23__14, 
                  ordered_filter_data_23__13, ordered_filter_data_23__12, 
                  ordered_filter_data_23__11, ordered_filter_data_23__10, 
                  ordered_filter_data_23__9, ordered_filter_data_23__8, 
                  ordered_filter_data_23__7, ordered_filter_data_23__6, 
                  ordered_filter_data_23__5, ordered_filter_data_23__4, 
                  ordered_filter_data_23__3, ordered_filter_data_23__2, 
                  ordered_filter_data_23__1, ordered_filter_data_23__0, 
                  ordered_filter_data_24__31, ordered_filter_data_24__30, 
                  ordered_filter_data_24__29, ordered_filter_data_24__28, 
                  ordered_filter_data_24__27, ordered_filter_data_24__26, 
                  ordered_filter_data_24__25, ordered_filter_data_24__24, 
                  ordered_filter_data_24__23, ordered_filter_data_24__22, 
                  ordered_filter_data_24__21, ordered_filter_data_24__20, 
                  ordered_filter_data_24__19, ordered_filter_data_24__18, 
                  ordered_filter_data_24__17, ordered_filter_data_24__16, 
                  ordered_filter_data_24__15, ordered_filter_data_24__14, 
                  ordered_filter_data_24__13, ordered_filter_data_24__12, 
                  ordered_filter_data_24__11, ordered_filter_data_24__10, 
                  ordered_filter_data_24__9, ordered_filter_data_24__8, 
                  ordered_filter_data_24__7, ordered_filter_data_24__6, 
                  ordered_filter_data_24__5, ordered_filter_data_24__4, 
                  ordered_filter_data_24__3, ordered_filter_data_24__2, 
                  ordered_filter_data_24__1, ordered_filter_data_24__0 ) ;

    input img_data_0__31 ;
    input img_data_0__30 ;
    input img_data_0__29 ;
    input img_data_0__28 ;
    input img_data_0__27 ;
    input img_data_0__26 ;
    input img_data_0__25 ;
    input img_data_0__24 ;
    input img_data_0__23 ;
    input img_data_0__22 ;
    input img_data_0__21 ;
    input img_data_0__20 ;
    input img_data_0__19 ;
    input img_data_0__18 ;
    input img_data_0__17 ;
    input img_data_0__16 ;
    input img_data_0__15 ;
    input img_data_0__14 ;
    input img_data_0__13 ;
    input img_data_0__12 ;
    input img_data_0__11 ;
    input img_data_0__10 ;
    input img_data_0__9 ;
    input img_data_0__8 ;
    input img_data_0__7 ;
    input img_data_0__6 ;
    input img_data_0__5 ;
    input img_data_0__4 ;
    input img_data_0__3 ;
    input img_data_0__2 ;
    input img_data_0__1 ;
    input img_data_0__0 ;
    input img_data_1__31 ;
    input img_data_1__30 ;
    input img_data_1__29 ;
    input img_data_1__28 ;
    input img_data_1__27 ;
    input img_data_1__26 ;
    input img_data_1__25 ;
    input img_data_1__24 ;
    input img_data_1__23 ;
    input img_data_1__22 ;
    input img_data_1__21 ;
    input img_data_1__20 ;
    input img_data_1__19 ;
    input img_data_1__18 ;
    input img_data_1__17 ;
    input img_data_1__16 ;
    input img_data_1__15 ;
    input img_data_1__14 ;
    input img_data_1__13 ;
    input img_data_1__12 ;
    input img_data_1__11 ;
    input img_data_1__10 ;
    input img_data_1__9 ;
    input img_data_1__8 ;
    input img_data_1__7 ;
    input img_data_1__6 ;
    input img_data_1__5 ;
    input img_data_1__4 ;
    input img_data_1__3 ;
    input img_data_1__2 ;
    input img_data_1__1 ;
    input img_data_1__0 ;
    input img_data_2__31 ;
    input img_data_2__30 ;
    input img_data_2__29 ;
    input img_data_2__28 ;
    input img_data_2__27 ;
    input img_data_2__26 ;
    input img_data_2__25 ;
    input img_data_2__24 ;
    input img_data_2__23 ;
    input img_data_2__22 ;
    input img_data_2__21 ;
    input img_data_2__20 ;
    input img_data_2__19 ;
    input img_data_2__18 ;
    input img_data_2__17 ;
    input img_data_2__16 ;
    input img_data_2__15 ;
    input img_data_2__14 ;
    input img_data_2__13 ;
    input img_data_2__12 ;
    input img_data_2__11 ;
    input img_data_2__10 ;
    input img_data_2__9 ;
    input img_data_2__8 ;
    input img_data_2__7 ;
    input img_data_2__6 ;
    input img_data_2__5 ;
    input img_data_2__4 ;
    input img_data_2__3 ;
    input img_data_2__2 ;
    input img_data_2__1 ;
    input img_data_2__0 ;
    input img_data_3__31 ;
    input img_data_3__30 ;
    input img_data_3__29 ;
    input img_data_3__28 ;
    input img_data_3__27 ;
    input img_data_3__26 ;
    input img_data_3__25 ;
    input img_data_3__24 ;
    input img_data_3__23 ;
    input img_data_3__22 ;
    input img_data_3__21 ;
    input img_data_3__20 ;
    input img_data_3__19 ;
    input img_data_3__18 ;
    input img_data_3__17 ;
    input img_data_3__16 ;
    input img_data_3__15 ;
    input img_data_3__14 ;
    input img_data_3__13 ;
    input img_data_3__12 ;
    input img_data_3__11 ;
    input img_data_3__10 ;
    input img_data_3__9 ;
    input img_data_3__8 ;
    input img_data_3__7 ;
    input img_data_3__6 ;
    input img_data_3__5 ;
    input img_data_3__4 ;
    input img_data_3__3 ;
    input img_data_3__2 ;
    input img_data_3__1 ;
    input img_data_3__0 ;
    input img_data_4__31 ;
    input img_data_4__30 ;
    input img_data_4__29 ;
    input img_data_4__28 ;
    input img_data_4__27 ;
    input img_data_4__26 ;
    input img_data_4__25 ;
    input img_data_4__24 ;
    input img_data_4__23 ;
    input img_data_4__22 ;
    input img_data_4__21 ;
    input img_data_4__20 ;
    input img_data_4__19 ;
    input img_data_4__18 ;
    input img_data_4__17 ;
    input img_data_4__16 ;
    input img_data_4__15 ;
    input img_data_4__14 ;
    input img_data_4__13 ;
    input img_data_4__12 ;
    input img_data_4__11 ;
    input img_data_4__10 ;
    input img_data_4__9 ;
    input img_data_4__8 ;
    input img_data_4__7 ;
    input img_data_4__6 ;
    input img_data_4__5 ;
    input img_data_4__4 ;
    input img_data_4__3 ;
    input img_data_4__2 ;
    input img_data_4__1 ;
    input img_data_4__0 ;
    input img_data_5__31 ;
    input img_data_5__30 ;
    input img_data_5__29 ;
    input img_data_5__28 ;
    input img_data_5__27 ;
    input img_data_5__26 ;
    input img_data_5__25 ;
    input img_data_5__24 ;
    input img_data_5__23 ;
    input img_data_5__22 ;
    input img_data_5__21 ;
    input img_data_5__20 ;
    input img_data_5__19 ;
    input img_data_5__18 ;
    input img_data_5__17 ;
    input img_data_5__16 ;
    input img_data_5__15 ;
    input img_data_5__14 ;
    input img_data_5__13 ;
    input img_data_5__12 ;
    input img_data_5__11 ;
    input img_data_5__10 ;
    input img_data_5__9 ;
    input img_data_5__8 ;
    input img_data_5__7 ;
    input img_data_5__6 ;
    input img_data_5__5 ;
    input img_data_5__4 ;
    input img_data_5__3 ;
    input img_data_5__2 ;
    input img_data_5__1 ;
    input img_data_5__0 ;
    input img_data_6__31 ;
    input img_data_6__30 ;
    input img_data_6__29 ;
    input img_data_6__28 ;
    input img_data_6__27 ;
    input img_data_6__26 ;
    input img_data_6__25 ;
    input img_data_6__24 ;
    input img_data_6__23 ;
    input img_data_6__22 ;
    input img_data_6__21 ;
    input img_data_6__20 ;
    input img_data_6__19 ;
    input img_data_6__18 ;
    input img_data_6__17 ;
    input img_data_6__16 ;
    input img_data_6__15 ;
    input img_data_6__14 ;
    input img_data_6__13 ;
    input img_data_6__12 ;
    input img_data_6__11 ;
    input img_data_6__10 ;
    input img_data_6__9 ;
    input img_data_6__8 ;
    input img_data_6__7 ;
    input img_data_6__6 ;
    input img_data_6__5 ;
    input img_data_6__4 ;
    input img_data_6__3 ;
    input img_data_6__2 ;
    input img_data_6__1 ;
    input img_data_6__0 ;
    input img_data_7__31 ;
    input img_data_7__30 ;
    input img_data_7__29 ;
    input img_data_7__28 ;
    input img_data_7__27 ;
    input img_data_7__26 ;
    input img_data_7__25 ;
    input img_data_7__24 ;
    input img_data_7__23 ;
    input img_data_7__22 ;
    input img_data_7__21 ;
    input img_data_7__20 ;
    input img_data_7__19 ;
    input img_data_7__18 ;
    input img_data_7__17 ;
    input img_data_7__16 ;
    input img_data_7__15 ;
    input img_data_7__14 ;
    input img_data_7__13 ;
    input img_data_7__12 ;
    input img_data_7__11 ;
    input img_data_7__10 ;
    input img_data_7__9 ;
    input img_data_7__8 ;
    input img_data_7__7 ;
    input img_data_7__6 ;
    input img_data_7__5 ;
    input img_data_7__4 ;
    input img_data_7__3 ;
    input img_data_7__2 ;
    input img_data_7__1 ;
    input img_data_7__0 ;
    input img_data_8__31 ;
    input img_data_8__30 ;
    input img_data_8__29 ;
    input img_data_8__28 ;
    input img_data_8__27 ;
    input img_data_8__26 ;
    input img_data_8__25 ;
    input img_data_8__24 ;
    input img_data_8__23 ;
    input img_data_8__22 ;
    input img_data_8__21 ;
    input img_data_8__20 ;
    input img_data_8__19 ;
    input img_data_8__18 ;
    input img_data_8__17 ;
    input img_data_8__16 ;
    input img_data_8__15 ;
    input img_data_8__14 ;
    input img_data_8__13 ;
    input img_data_8__12 ;
    input img_data_8__11 ;
    input img_data_8__10 ;
    input img_data_8__9 ;
    input img_data_8__8 ;
    input img_data_8__7 ;
    input img_data_8__6 ;
    input img_data_8__5 ;
    input img_data_8__4 ;
    input img_data_8__3 ;
    input img_data_8__2 ;
    input img_data_8__1 ;
    input img_data_8__0 ;
    input img_data_9__31 ;
    input img_data_9__30 ;
    input img_data_9__29 ;
    input img_data_9__28 ;
    input img_data_9__27 ;
    input img_data_9__26 ;
    input img_data_9__25 ;
    input img_data_9__24 ;
    input img_data_9__23 ;
    input img_data_9__22 ;
    input img_data_9__21 ;
    input img_data_9__20 ;
    input img_data_9__19 ;
    input img_data_9__18 ;
    input img_data_9__17 ;
    input img_data_9__16 ;
    input img_data_9__15 ;
    input img_data_9__14 ;
    input img_data_9__13 ;
    input img_data_9__12 ;
    input img_data_9__11 ;
    input img_data_9__10 ;
    input img_data_9__9 ;
    input img_data_9__8 ;
    input img_data_9__7 ;
    input img_data_9__6 ;
    input img_data_9__5 ;
    input img_data_9__4 ;
    input img_data_9__3 ;
    input img_data_9__2 ;
    input img_data_9__1 ;
    input img_data_9__0 ;
    input img_data_10__31 ;
    input img_data_10__30 ;
    input img_data_10__29 ;
    input img_data_10__28 ;
    input img_data_10__27 ;
    input img_data_10__26 ;
    input img_data_10__25 ;
    input img_data_10__24 ;
    input img_data_10__23 ;
    input img_data_10__22 ;
    input img_data_10__21 ;
    input img_data_10__20 ;
    input img_data_10__19 ;
    input img_data_10__18 ;
    input img_data_10__17 ;
    input img_data_10__16 ;
    input img_data_10__15 ;
    input img_data_10__14 ;
    input img_data_10__13 ;
    input img_data_10__12 ;
    input img_data_10__11 ;
    input img_data_10__10 ;
    input img_data_10__9 ;
    input img_data_10__8 ;
    input img_data_10__7 ;
    input img_data_10__6 ;
    input img_data_10__5 ;
    input img_data_10__4 ;
    input img_data_10__3 ;
    input img_data_10__2 ;
    input img_data_10__1 ;
    input img_data_10__0 ;
    input img_data_11__31 ;
    input img_data_11__30 ;
    input img_data_11__29 ;
    input img_data_11__28 ;
    input img_data_11__27 ;
    input img_data_11__26 ;
    input img_data_11__25 ;
    input img_data_11__24 ;
    input img_data_11__23 ;
    input img_data_11__22 ;
    input img_data_11__21 ;
    input img_data_11__20 ;
    input img_data_11__19 ;
    input img_data_11__18 ;
    input img_data_11__17 ;
    input img_data_11__16 ;
    input img_data_11__15 ;
    input img_data_11__14 ;
    input img_data_11__13 ;
    input img_data_11__12 ;
    input img_data_11__11 ;
    input img_data_11__10 ;
    input img_data_11__9 ;
    input img_data_11__8 ;
    input img_data_11__7 ;
    input img_data_11__6 ;
    input img_data_11__5 ;
    input img_data_11__4 ;
    input img_data_11__3 ;
    input img_data_11__2 ;
    input img_data_11__1 ;
    input img_data_11__0 ;
    input img_data_12__31 ;
    input img_data_12__30 ;
    input img_data_12__29 ;
    input img_data_12__28 ;
    input img_data_12__27 ;
    input img_data_12__26 ;
    input img_data_12__25 ;
    input img_data_12__24 ;
    input img_data_12__23 ;
    input img_data_12__22 ;
    input img_data_12__21 ;
    input img_data_12__20 ;
    input img_data_12__19 ;
    input img_data_12__18 ;
    input img_data_12__17 ;
    input img_data_12__16 ;
    input img_data_12__15 ;
    input img_data_12__14 ;
    input img_data_12__13 ;
    input img_data_12__12 ;
    input img_data_12__11 ;
    input img_data_12__10 ;
    input img_data_12__9 ;
    input img_data_12__8 ;
    input img_data_12__7 ;
    input img_data_12__6 ;
    input img_data_12__5 ;
    input img_data_12__4 ;
    input img_data_12__3 ;
    input img_data_12__2 ;
    input img_data_12__1 ;
    input img_data_12__0 ;
    input img_data_13__31 ;
    input img_data_13__30 ;
    input img_data_13__29 ;
    input img_data_13__28 ;
    input img_data_13__27 ;
    input img_data_13__26 ;
    input img_data_13__25 ;
    input img_data_13__24 ;
    input img_data_13__23 ;
    input img_data_13__22 ;
    input img_data_13__21 ;
    input img_data_13__20 ;
    input img_data_13__19 ;
    input img_data_13__18 ;
    input img_data_13__17 ;
    input img_data_13__16 ;
    input img_data_13__15 ;
    input img_data_13__14 ;
    input img_data_13__13 ;
    input img_data_13__12 ;
    input img_data_13__11 ;
    input img_data_13__10 ;
    input img_data_13__9 ;
    input img_data_13__8 ;
    input img_data_13__7 ;
    input img_data_13__6 ;
    input img_data_13__5 ;
    input img_data_13__4 ;
    input img_data_13__3 ;
    input img_data_13__2 ;
    input img_data_13__1 ;
    input img_data_13__0 ;
    input img_data_14__31 ;
    input img_data_14__30 ;
    input img_data_14__29 ;
    input img_data_14__28 ;
    input img_data_14__27 ;
    input img_data_14__26 ;
    input img_data_14__25 ;
    input img_data_14__24 ;
    input img_data_14__23 ;
    input img_data_14__22 ;
    input img_data_14__21 ;
    input img_data_14__20 ;
    input img_data_14__19 ;
    input img_data_14__18 ;
    input img_data_14__17 ;
    input img_data_14__16 ;
    input img_data_14__15 ;
    input img_data_14__14 ;
    input img_data_14__13 ;
    input img_data_14__12 ;
    input img_data_14__11 ;
    input img_data_14__10 ;
    input img_data_14__9 ;
    input img_data_14__8 ;
    input img_data_14__7 ;
    input img_data_14__6 ;
    input img_data_14__5 ;
    input img_data_14__4 ;
    input img_data_14__3 ;
    input img_data_14__2 ;
    input img_data_14__1 ;
    input img_data_14__0 ;
    input img_data_15__31 ;
    input img_data_15__30 ;
    input img_data_15__29 ;
    input img_data_15__28 ;
    input img_data_15__27 ;
    input img_data_15__26 ;
    input img_data_15__25 ;
    input img_data_15__24 ;
    input img_data_15__23 ;
    input img_data_15__22 ;
    input img_data_15__21 ;
    input img_data_15__20 ;
    input img_data_15__19 ;
    input img_data_15__18 ;
    input img_data_15__17 ;
    input img_data_15__16 ;
    input img_data_15__15 ;
    input img_data_15__14 ;
    input img_data_15__13 ;
    input img_data_15__12 ;
    input img_data_15__11 ;
    input img_data_15__10 ;
    input img_data_15__9 ;
    input img_data_15__8 ;
    input img_data_15__7 ;
    input img_data_15__6 ;
    input img_data_15__5 ;
    input img_data_15__4 ;
    input img_data_15__3 ;
    input img_data_15__2 ;
    input img_data_15__1 ;
    input img_data_15__0 ;
    input img_data_16__31 ;
    input img_data_16__30 ;
    input img_data_16__29 ;
    input img_data_16__28 ;
    input img_data_16__27 ;
    input img_data_16__26 ;
    input img_data_16__25 ;
    input img_data_16__24 ;
    input img_data_16__23 ;
    input img_data_16__22 ;
    input img_data_16__21 ;
    input img_data_16__20 ;
    input img_data_16__19 ;
    input img_data_16__18 ;
    input img_data_16__17 ;
    input img_data_16__16 ;
    input img_data_16__15 ;
    input img_data_16__14 ;
    input img_data_16__13 ;
    input img_data_16__12 ;
    input img_data_16__11 ;
    input img_data_16__10 ;
    input img_data_16__9 ;
    input img_data_16__8 ;
    input img_data_16__7 ;
    input img_data_16__6 ;
    input img_data_16__5 ;
    input img_data_16__4 ;
    input img_data_16__3 ;
    input img_data_16__2 ;
    input img_data_16__1 ;
    input img_data_16__0 ;
    input img_data_17__31 ;
    input img_data_17__30 ;
    input img_data_17__29 ;
    input img_data_17__28 ;
    input img_data_17__27 ;
    input img_data_17__26 ;
    input img_data_17__25 ;
    input img_data_17__24 ;
    input img_data_17__23 ;
    input img_data_17__22 ;
    input img_data_17__21 ;
    input img_data_17__20 ;
    input img_data_17__19 ;
    input img_data_17__18 ;
    input img_data_17__17 ;
    input img_data_17__16 ;
    input img_data_17__15 ;
    input img_data_17__14 ;
    input img_data_17__13 ;
    input img_data_17__12 ;
    input img_data_17__11 ;
    input img_data_17__10 ;
    input img_data_17__9 ;
    input img_data_17__8 ;
    input img_data_17__7 ;
    input img_data_17__6 ;
    input img_data_17__5 ;
    input img_data_17__4 ;
    input img_data_17__3 ;
    input img_data_17__2 ;
    input img_data_17__1 ;
    input img_data_17__0 ;
    input img_data_18__31 ;
    input img_data_18__30 ;
    input img_data_18__29 ;
    input img_data_18__28 ;
    input img_data_18__27 ;
    input img_data_18__26 ;
    input img_data_18__25 ;
    input img_data_18__24 ;
    input img_data_18__23 ;
    input img_data_18__22 ;
    input img_data_18__21 ;
    input img_data_18__20 ;
    input img_data_18__19 ;
    input img_data_18__18 ;
    input img_data_18__17 ;
    input img_data_18__16 ;
    input img_data_18__15 ;
    input img_data_18__14 ;
    input img_data_18__13 ;
    input img_data_18__12 ;
    input img_data_18__11 ;
    input img_data_18__10 ;
    input img_data_18__9 ;
    input img_data_18__8 ;
    input img_data_18__7 ;
    input img_data_18__6 ;
    input img_data_18__5 ;
    input img_data_18__4 ;
    input img_data_18__3 ;
    input img_data_18__2 ;
    input img_data_18__1 ;
    input img_data_18__0 ;
    input img_data_19__31 ;
    input img_data_19__30 ;
    input img_data_19__29 ;
    input img_data_19__28 ;
    input img_data_19__27 ;
    input img_data_19__26 ;
    input img_data_19__25 ;
    input img_data_19__24 ;
    input img_data_19__23 ;
    input img_data_19__22 ;
    input img_data_19__21 ;
    input img_data_19__20 ;
    input img_data_19__19 ;
    input img_data_19__18 ;
    input img_data_19__17 ;
    input img_data_19__16 ;
    input img_data_19__15 ;
    input img_data_19__14 ;
    input img_data_19__13 ;
    input img_data_19__12 ;
    input img_data_19__11 ;
    input img_data_19__10 ;
    input img_data_19__9 ;
    input img_data_19__8 ;
    input img_data_19__7 ;
    input img_data_19__6 ;
    input img_data_19__5 ;
    input img_data_19__4 ;
    input img_data_19__3 ;
    input img_data_19__2 ;
    input img_data_19__1 ;
    input img_data_19__0 ;
    input img_data_20__31 ;
    input img_data_20__30 ;
    input img_data_20__29 ;
    input img_data_20__28 ;
    input img_data_20__27 ;
    input img_data_20__26 ;
    input img_data_20__25 ;
    input img_data_20__24 ;
    input img_data_20__23 ;
    input img_data_20__22 ;
    input img_data_20__21 ;
    input img_data_20__20 ;
    input img_data_20__19 ;
    input img_data_20__18 ;
    input img_data_20__17 ;
    input img_data_20__16 ;
    input img_data_20__15 ;
    input img_data_20__14 ;
    input img_data_20__13 ;
    input img_data_20__12 ;
    input img_data_20__11 ;
    input img_data_20__10 ;
    input img_data_20__9 ;
    input img_data_20__8 ;
    input img_data_20__7 ;
    input img_data_20__6 ;
    input img_data_20__5 ;
    input img_data_20__4 ;
    input img_data_20__3 ;
    input img_data_20__2 ;
    input img_data_20__1 ;
    input img_data_20__0 ;
    input img_data_21__31 ;
    input img_data_21__30 ;
    input img_data_21__29 ;
    input img_data_21__28 ;
    input img_data_21__27 ;
    input img_data_21__26 ;
    input img_data_21__25 ;
    input img_data_21__24 ;
    input img_data_21__23 ;
    input img_data_21__22 ;
    input img_data_21__21 ;
    input img_data_21__20 ;
    input img_data_21__19 ;
    input img_data_21__18 ;
    input img_data_21__17 ;
    input img_data_21__16 ;
    input img_data_21__15 ;
    input img_data_21__14 ;
    input img_data_21__13 ;
    input img_data_21__12 ;
    input img_data_21__11 ;
    input img_data_21__10 ;
    input img_data_21__9 ;
    input img_data_21__8 ;
    input img_data_21__7 ;
    input img_data_21__6 ;
    input img_data_21__5 ;
    input img_data_21__4 ;
    input img_data_21__3 ;
    input img_data_21__2 ;
    input img_data_21__1 ;
    input img_data_21__0 ;
    input img_data_22__31 ;
    input img_data_22__30 ;
    input img_data_22__29 ;
    input img_data_22__28 ;
    input img_data_22__27 ;
    input img_data_22__26 ;
    input img_data_22__25 ;
    input img_data_22__24 ;
    input img_data_22__23 ;
    input img_data_22__22 ;
    input img_data_22__21 ;
    input img_data_22__20 ;
    input img_data_22__19 ;
    input img_data_22__18 ;
    input img_data_22__17 ;
    input img_data_22__16 ;
    input img_data_22__15 ;
    input img_data_22__14 ;
    input img_data_22__13 ;
    input img_data_22__12 ;
    input img_data_22__11 ;
    input img_data_22__10 ;
    input img_data_22__9 ;
    input img_data_22__8 ;
    input img_data_22__7 ;
    input img_data_22__6 ;
    input img_data_22__5 ;
    input img_data_22__4 ;
    input img_data_22__3 ;
    input img_data_22__2 ;
    input img_data_22__1 ;
    input img_data_22__0 ;
    input img_data_23__31 ;
    input img_data_23__30 ;
    input img_data_23__29 ;
    input img_data_23__28 ;
    input img_data_23__27 ;
    input img_data_23__26 ;
    input img_data_23__25 ;
    input img_data_23__24 ;
    input img_data_23__23 ;
    input img_data_23__22 ;
    input img_data_23__21 ;
    input img_data_23__20 ;
    input img_data_23__19 ;
    input img_data_23__18 ;
    input img_data_23__17 ;
    input img_data_23__16 ;
    input img_data_23__15 ;
    input img_data_23__14 ;
    input img_data_23__13 ;
    input img_data_23__12 ;
    input img_data_23__11 ;
    input img_data_23__10 ;
    input img_data_23__9 ;
    input img_data_23__8 ;
    input img_data_23__7 ;
    input img_data_23__6 ;
    input img_data_23__5 ;
    input img_data_23__4 ;
    input img_data_23__3 ;
    input img_data_23__2 ;
    input img_data_23__1 ;
    input img_data_23__0 ;
    input img_data_24__31 ;
    input img_data_24__30 ;
    input img_data_24__29 ;
    input img_data_24__28 ;
    input img_data_24__27 ;
    input img_data_24__26 ;
    input img_data_24__25 ;
    input img_data_24__24 ;
    input img_data_24__23 ;
    input img_data_24__22 ;
    input img_data_24__21 ;
    input img_data_24__20 ;
    input img_data_24__19 ;
    input img_data_24__18 ;
    input img_data_24__17 ;
    input img_data_24__16 ;
    input img_data_24__15 ;
    input img_data_24__14 ;
    input img_data_24__13 ;
    input img_data_24__12 ;
    input img_data_24__11 ;
    input img_data_24__10 ;
    input img_data_24__9 ;
    input img_data_24__8 ;
    input img_data_24__7 ;
    input img_data_24__6 ;
    input img_data_24__5 ;
    input img_data_24__4 ;
    input img_data_24__3 ;
    input img_data_24__2 ;
    input img_data_24__1 ;
    input img_data_24__0 ;
    input filter_data_0__31 ;
    input filter_data_0__30 ;
    input filter_data_0__29 ;
    input filter_data_0__28 ;
    input filter_data_0__27 ;
    input filter_data_0__26 ;
    input filter_data_0__25 ;
    input filter_data_0__24 ;
    input filter_data_0__23 ;
    input filter_data_0__22 ;
    input filter_data_0__21 ;
    input filter_data_0__20 ;
    input filter_data_0__19 ;
    input filter_data_0__18 ;
    input filter_data_0__17 ;
    input filter_data_0__16 ;
    input filter_data_0__15 ;
    input filter_data_0__14 ;
    input filter_data_0__13 ;
    input filter_data_0__12 ;
    input filter_data_0__11 ;
    input filter_data_0__10 ;
    input filter_data_0__9 ;
    input filter_data_0__8 ;
    input filter_data_0__7 ;
    input filter_data_0__6 ;
    input filter_data_0__5 ;
    input filter_data_0__4 ;
    input filter_data_0__3 ;
    input filter_data_0__2 ;
    input filter_data_0__1 ;
    input filter_data_0__0 ;
    input filter_data_1__31 ;
    input filter_data_1__30 ;
    input filter_data_1__29 ;
    input filter_data_1__28 ;
    input filter_data_1__27 ;
    input filter_data_1__26 ;
    input filter_data_1__25 ;
    input filter_data_1__24 ;
    input filter_data_1__23 ;
    input filter_data_1__22 ;
    input filter_data_1__21 ;
    input filter_data_1__20 ;
    input filter_data_1__19 ;
    input filter_data_1__18 ;
    input filter_data_1__17 ;
    input filter_data_1__16 ;
    input filter_data_1__15 ;
    input filter_data_1__14 ;
    input filter_data_1__13 ;
    input filter_data_1__12 ;
    input filter_data_1__11 ;
    input filter_data_1__10 ;
    input filter_data_1__9 ;
    input filter_data_1__8 ;
    input filter_data_1__7 ;
    input filter_data_1__6 ;
    input filter_data_1__5 ;
    input filter_data_1__4 ;
    input filter_data_1__3 ;
    input filter_data_1__2 ;
    input filter_data_1__1 ;
    input filter_data_1__0 ;
    input filter_data_2__31 ;
    input filter_data_2__30 ;
    input filter_data_2__29 ;
    input filter_data_2__28 ;
    input filter_data_2__27 ;
    input filter_data_2__26 ;
    input filter_data_2__25 ;
    input filter_data_2__24 ;
    input filter_data_2__23 ;
    input filter_data_2__22 ;
    input filter_data_2__21 ;
    input filter_data_2__20 ;
    input filter_data_2__19 ;
    input filter_data_2__18 ;
    input filter_data_2__17 ;
    input filter_data_2__16 ;
    input filter_data_2__15 ;
    input filter_data_2__14 ;
    input filter_data_2__13 ;
    input filter_data_2__12 ;
    input filter_data_2__11 ;
    input filter_data_2__10 ;
    input filter_data_2__9 ;
    input filter_data_2__8 ;
    input filter_data_2__7 ;
    input filter_data_2__6 ;
    input filter_data_2__5 ;
    input filter_data_2__4 ;
    input filter_data_2__3 ;
    input filter_data_2__2 ;
    input filter_data_2__1 ;
    input filter_data_2__0 ;
    input filter_data_3__31 ;
    input filter_data_3__30 ;
    input filter_data_3__29 ;
    input filter_data_3__28 ;
    input filter_data_3__27 ;
    input filter_data_3__26 ;
    input filter_data_3__25 ;
    input filter_data_3__24 ;
    input filter_data_3__23 ;
    input filter_data_3__22 ;
    input filter_data_3__21 ;
    input filter_data_3__20 ;
    input filter_data_3__19 ;
    input filter_data_3__18 ;
    input filter_data_3__17 ;
    input filter_data_3__16 ;
    input filter_data_3__15 ;
    input filter_data_3__14 ;
    input filter_data_3__13 ;
    input filter_data_3__12 ;
    input filter_data_3__11 ;
    input filter_data_3__10 ;
    input filter_data_3__9 ;
    input filter_data_3__8 ;
    input filter_data_3__7 ;
    input filter_data_3__6 ;
    input filter_data_3__5 ;
    input filter_data_3__4 ;
    input filter_data_3__3 ;
    input filter_data_3__2 ;
    input filter_data_3__1 ;
    input filter_data_3__0 ;
    input filter_data_4__31 ;
    input filter_data_4__30 ;
    input filter_data_4__29 ;
    input filter_data_4__28 ;
    input filter_data_4__27 ;
    input filter_data_4__26 ;
    input filter_data_4__25 ;
    input filter_data_4__24 ;
    input filter_data_4__23 ;
    input filter_data_4__22 ;
    input filter_data_4__21 ;
    input filter_data_4__20 ;
    input filter_data_4__19 ;
    input filter_data_4__18 ;
    input filter_data_4__17 ;
    input filter_data_4__16 ;
    input filter_data_4__15 ;
    input filter_data_4__14 ;
    input filter_data_4__13 ;
    input filter_data_4__12 ;
    input filter_data_4__11 ;
    input filter_data_4__10 ;
    input filter_data_4__9 ;
    input filter_data_4__8 ;
    input filter_data_4__7 ;
    input filter_data_4__6 ;
    input filter_data_4__5 ;
    input filter_data_4__4 ;
    input filter_data_4__3 ;
    input filter_data_4__2 ;
    input filter_data_4__1 ;
    input filter_data_4__0 ;
    input filter_data_5__31 ;
    input filter_data_5__30 ;
    input filter_data_5__29 ;
    input filter_data_5__28 ;
    input filter_data_5__27 ;
    input filter_data_5__26 ;
    input filter_data_5__25 ;
    input filter_data_5__24 ;
    input filter_data_5__23 ;
    input filter_data_5__22 ;
    input filter_data_5__21 ;
    input filter_data_5__20 ;
    input filter_data_5__19 ;
    input filter_data_5__18 ;
    input filter_data_5__17 ;
    input filter_data_5__16 ;
    input filter_data_5__15 ;
    input filter_data_5__14 ;
    input filter_data_5__13 ;
    input filter_data_5__12 ;
    input filter_data_5__11 ;
    input filter_data_5__10 ;
    input filter_data_5__9 ;
    input filter_data_5__8 ;
    input filter_data_5__7 ;
    input filter_data_5__6 ;
    input filter_data_5__5 ;
    input filter_data_5__4 ;
    input filter_data_5__3 ;
    input filter_data_5__2 ;
    input filter_data_5__1 ;
    input filter_data_5__0 ;
    input filter_data_6__31 ;
    input filter_data_6__30 ;
    input filter_data_6__29 ;
    input filter_data_6__28 ;
    input filter_data_6__27 ;
    input filter_data_6__26 ;
    input filter_data_6__25 ;
    input filter_data_6__24 ;
    input filter_data_6__23 ;
    input filter_data_6__22 ;
    input filter_data_6__21 ;
    input filter_data_6__20 ;
    input filter_data_6__19 ;
    input filter_data_6__18 ;
    input filter_data_6__17 ;
    input filter_data_6__16 ;
    input filter_data_6__15 ;
    input filter_data_6__14 ;
    input filter_data_6__13 ;
    input filter_data_6__12 ;
    input filter_data_6__11 ;
    input filter_data_6__10 ;
    input filter_data_6__9 ;
    input filter_data_6__8 ;
    input filter_data_6__7 ;
    input filter_data_6__6 ;
    input filter_data_6__5 ;
    input filter_data_6__4 ;
    input filter_data_6__3 ;
    input filter_data_6__2 ;
    input filter_data_6__1 ;
    input filter_data_6__0 ;
    input filter_data_7__31 ;
    input filter_data_7__30 ;
    input filter_data_7__29 ;
    input filter_data_7__28 ;
    input filter_data_7__27 ;
    input filter_data_7__26 ;
    input filter_data_7__25 ;
    input filter_data_7__24 ;
    input filter_data_7__23 ;
    input filter_data_7__22 ;
    input filter_data_7__21 ;
    input filter_data_7__20 ;
    input filter_data_7__19 ;
    input filter_data_7__18 ;
    input filter_data_7__17 ;
    input filter_data_7__16 ;
    input filter_data_7__15 ;
    input filter_data_7__14 ;
    input filter_data_7__13 ;
    input filter_data_7__12 ;
    input filter_data_7__11 ;
    input filter_data_7__10 ;
    input filter_data_7__9 ;
    input filter_data_7__8 ;
    input filter_data_7__7 ;
    input filter_data_7__6 ;
    input filter_data_7__5 ;
    input filter_data_7__4 ;
    input filter_data_7__3 ;
    input filter_data_7__2 ;
    input filter_data_7__1 ;
    input filter_data_7__0 ;
    input filter_data_8__31 ;
    input filter_data_8__30 ;
    input filter_data_8__29 ;
    input filter_data_8__28 ;
    input filter_data_8__27 ;
    input filter_data_8__26 ;
    input filter_data_8__25 ;
    input filter_data_8__24 ;
    input filter_data_8__23 ;
    input filter_data_8__22 ;
    input filter_data_8__21 ;
    input filter_data_8__20 ;
    input filter_data_8__19 ;
    input filter_data_8__18 ;
    input filter_data_8__17 ;
    input filter_data_8__16 ;
    input filter_data_8__15 ;
    input filter_data_8__14 ;
    input filter_data_8__13 ;
    input filter_data_8__12 ;
    input filter_data_8__11 ;
    input filter_data_8__10 ;
    input filter_data_8__9 ;
    input filter_data_8__8 ;
    input filter_data_8__7 ;
    input filter_data_8__6 ;
    input filter_data_8__5 ;
    input filter_data_8__4 ;
    input filter_data_8__3 ;
    input filter_data_8__2 ;
    input filter_data_8__1 ;
    input filter_data_8__0 ;
    input filter_data_9__31 ;
    input filter_data_9__30 ;
    input filter_data_9__29 ;
    input filter_data_9__28 ;
    input filter_data_9__27 ;
    input filter_data_9__26 ;
    input filter_data_9__25 ;
    input filter_data_9__24 ;
    input filter_data_9__23 ;
    input filter_data_9__22 ;
    input filter_data_9__21 ;
    input filter_data_9__20 ;
    input filter_data_9__19 ;
    input filter_data_9__18 ;
    input filter_data_9__17 ;
    input filter_data_9__16 ;
    input filter_data_9__15 ;
    input filter_data_9__14 ;
    input filter_data_9__13 ;
    input filter_data_9__12 ;
    input filter_data_9__11 ;
    input filter_data_9__10 ;
    input filter_data_9__9 ;
    input filter_data_9__8 ;
    input filter_data_9__7 ;
    input filter_data_9__6 ;
    input filter_data_9__5 ;
    input filter_data_9__4 ;
    input filter_data_9__3 ;
    input filter_data_9__2 ;
    input filter_data_9__1 ;
    input filter_data_9__0 ;
    input filter_data_10__31 ;
    input filter_data_10__30 ;
    input filter_data_10__29 ;
    input filter_data_10__28 ;
    input filter_data_10__27 ;
    input filter_data_10__26 ;
    input filter_data_10__25 ;
    input filter_data_10__24 ;
    input filter_data_10__23 ;
    input filter_data_10__22 ;
    input filter_data_10__21 ;
    input filter_data_10__20 ;
    input filter_data_10__19 ;
    input filter_data_10__18 ;
    input filter_data_10__17 ;
    input filter_data_10__16 ;
    input filter_data_10__15 ;
    input filter_data_10__14 ;
    input filter_data_10__13 ;
    input filter_data_10__12 ;
    input filter_data_10__11 ;
    input filter_data_10__10 ;
    input filter_data_10__9 ;
    input filter_data_10__8 ;
    input filter_data_10__7 ;
    input filter_data_10__6 ;
    input filter_data_10__5 ;
    input filter_data_10__4 ;
    input filter_data_10__3 ;
    input filter_data_10__2 ;
    input filter_data_10__1 ;
    input filter_data_10__0 ;
    input filter_data_11__31 ;
    input filter_data_11__30 ;
    input filter_data_11__29 ;
    input filter_data_11__28 ;
    input filter_data_11__27 ;
    input filter_data_11__26 ;
    input filter_data_11__25 ;
    input filter_data_11__24 ;
    input filter_data_11__23 ;
    input filter_data_11__22 ;
    input filter_data_11__21 ;
    input filter_data_11__20 ;
    input filter_data_11__19 ;
    input filter_data_11__18 ;
    input filter_data_11__17 ;
    input filter_data_11__16 ;
    input filter_data_11__15 ;
    input filter_data_11__14 ;
    input filter_data_11__13 ;
    input filter_data_11__12 ;
    input filter_data_11__11 ;
    input filter_data_11__10 ;
    input filter_data_11__9 ;
    input filter_data_11__8 ;
    input filter_data_11__7 ;
    input filter_data_11__6 ;
    input filter_data_11__5 ;
    input filter_data_11__4 ;
    input filter_data_11__3 ;
    input filter_data_11__2 ;
    input filter_data_11__1 ;
    input filter_data_11__0 ;
    input filter_data_12__31 ;
    input filter_data_12__30 ;
    input filter_data_12__29 ;
    input filter_data_12__28 ;
    input filter_data_12__27 ;
    input filter_data_12__26 ;
    input filter_data_12__25 ;
    input filter_data_12__24 ;
    input filter_data_12__23 ;
    input filter_data_12__22 ;
    input filter_data_12__21 ;
    input filter_data_12__20 ;
    input filter_data_12__19 ;
    input filter_data_12__18 ;
    input filter_data_12__17 ;
    input filter_data_12__16 ;
    input filter_data_12__15 ;
    input filter_data_12__14 ;
    input filter_data_12__13 ;
    input filter_data_12__12 ;
    input filter_data_12__11 ;
    input filter_data_12__10 ;
    input filter_data_12__9 ;
    input filter_data_12__8 ;
    input filter_data_12__7 ;
    input filter_data_12__6 ;
    input filter_data_12__5 ;
    input filter_data_12__4 ;
    input filter_data_12__3 ;
    input filter_data_12__2 ;
    input filter_data_12__1 ;
    input filter_data_12__0 ;
    input filter_data_13__31 ;
    input filter_data_13__30 ;
    input filter_data_13__29 ;
    input filter_data_13__28 ;
    input filter_data_13__27 ;
    input filter_data_13__26 ;
    input filter_data_13__25 ;
    input filter_data_13__24 ;
    input filter_data_13__23 ;
    input filter_data_13__22 ;
    input filter_data_13__21 ;
    input filter_data_13__20 ;
    input filter_data_13__19 ;
    input filter_data_13__18 ;
    input filter_data_13__17 ;
    input filter_data_13__16 ;
    input filter_data_13__15 ;
    input filter_data_13__14 ;
    input filter_data_13__13 ;
    input filter_data_13__12 ;
    input filter_data_13__11 ;
    input filter_data_13__10 ;
    input filter_data_13__9 ;
    input filter_data_13__8 ;
    input filter_data_13__7 ;
    input filter_data_13__6 ;
    input filter_data_13__5 ;
    input filter_data_13__4 ;
    input filter_data_13__3 ;
    input filter_data_13__2 ;
    input filter_data_13__1 ;
    input filter_data_13__0 ;
    input filter_data_14__31 ;
    input filter_data_14__30 ;
    input filter_data_14__29 ;
    input filter_data_14__28 ;
    input filter_data_14__27 ;
    input filter_data_14__26 ;
    input filter_data_14__25 ;
    input filter_data_14__24 ;
    input filter_data_14__23 ;
    input filter_data_14__22 ;
    input filter_data_14__21 ;
    input filter_data_14__20 ;
    input filter_data_14__19 ;
    input filter_data_14__18 ;
    input filter_data_14__17 ;
    input filter_data_14__16 ;
    input filter_data_14__15 ;
    input filter_data_14__14 ;
    input filter_data_14__13 ;
    input filter_data_14__12 ;
    input filter_data_14__11 ;
    input filter_data_14__10 ;
    input filter_data_14__9 ;
    input filter_data_14__8 ;
    input filter_data_14__7 ;
    input filter_data_14__6 ;
    input filter_data_14__5 ;
    input filter_data_14__4 ;
    input filter_data_14__3 ;
    input filter_data_14__2 ;
    input filter_data_14__1 ;
    input filter_data_14__0 ;
    input filter_data_15__31 ;
    input filter_data_15__30 ;
    input filter_data_15__29 ;
    input filter_data_15__28 ;
    input filter_data_15__27 ;
    input filter_data_15__26 ;
    input filter_data_15__25 ;
    input filter_data_15__24 ;
    input filter_data_15__23 ;
    input filter_data_15__22 ;
    input filter_data_15__21 ;
    input filter_data_15__20 ;
    input filter_data_15__19 ;
    input filter_data_15__18 ;
    input filter_data_15__17 ;
    input filter_data_15__16 ;
    input filter_data_15__15 ;
    input filter_data_15__14 ;
    input filter_data_15__13 ;
    input filter_data_15__12 ;
    input filter_data_15__11 ;
    input filter_data_15__10 ;
    input filter_data_15__9 ;
    input filter_data_15__8 ;
    input filter_data_15__7 ;
    input filter_data_15__6 ;
    input filter_data_15__5 ;
    input filter_data_15__4 ;
    input filter_data_15__3 ;
    input filter_data_15__2 ;
    input filter_data_15__1 ;
    input filter_data_15__0 ;
    input filter_data_16__31 ;
    input filter_data_16__30 ;
    input filter_data_16__29 ;
    input filter_data_16__28 ;
    input filter_data_16__27 ;
    input filter_data_16__26 ;
    input filter_data_16__25 ;
    input filter_data_16__24 ;
    input filter_data_16__23 ;
    input filter_data_16__22 ;
    input filter_data_16__21 ;
    input filter_data_16__20 ;
    input filter_data_16__19 ;
    input filter_data_16__18 ;
    input filter_data_16__17 ;
    input filter_data_16__16 ;
    input filter_data_16__15 ;
    input filter_data_16__14 ;
    input filter_data_16__13 ;
    input filter_data_16__12 ;
    input filter_data_16__11 ;
    input filter_data_16__10 ;
    input filter_data_16__9 ;
    input filter_data_16__8 ;
    input filter_data_16__7 ;
    input filter_data_16__6 ;
    input filter_data_16__5 ;
    input filter_data_16__4 ;
    input filter_data_16__3 ;
    input filter_data_16__2 ;
    input filter_data_16__1 ;
    input filter_data_16__0 ;
    input filter_data_17__31 ;
    input filter_data_17__30 ;
    input filter_data_17__29 ;
    input filter_data_17__28 ;
    input filter_data_17__27 ;
    input filter_data_17__26 ;
    input filter_data_17__25 ;
    input filter_data_17__24 ;
    input filter_data_17__23 ;
    input filter_data_17__22 ;
    input filter_data_17__21 ;
    input filter_data_17__20 ;
    input filter_data_17__19 ;
    input filter_data_17__18 ;
    input filter_data_17__17 ;
    input filter_data_17__16 ;
    input filter_data_17__15 ;
    input filter_data_17__14 ;
    input filter_data_17__13 ;
    input filter_data_17__12 ;
    input filter_data_17__11 ;
    input filter_data_17__10 ;
    input filter_data_17__9 ;
    input filter_data_17__8 ;
    input filter_data_17__7 ;
    input filter_data_17__6 ;
    input filter_data_17__5 ;
    input filter_data_17__4 ;
    input filter_data_17__3 ;
    input filter_data_17__2 ;
    input filter_data_17__1 ;
    input filter_data_17__0 ;
    input filter_data_18__31 ;
    input filter_data_18__30 ;
    input filter_data_18__29 ;
    input filter_data_18__28 ;
    input filter_data_18__27 ;
    input filter_data_18__26 ;
    input filter_data_18__25 ;
    input filter_data_18__24 ;
    input filter_data_18__23 ;
    input filter_data_18__22 ;
    input filter_data_18__21 ;
    input filter_data_18__20 ;
    input filter_data_18__19 ;
    input filter_data_18__18 ;
    input filter_data_18__17 ;
    input filter_data_18__16 ;
    input filter_data_18__15 ;
    input filter_data_18__14 ;
    input filter_data_18__13 ;
    input filter_data_18__12 ;
    input filter_data_18__11 ;
    input filter_data_18__10 ;
    input filter_data_18__9 ;
    input filter_data_18__8 ;
    input filter_data_18__7 ;
    input filter_data_18__6 ;
    input filter_data_18__5 ;
    input filter_data_18__4 ;
    input filter_data_18__3 ;
    input filter_data_18__2 ;
    input filter_data_18__1 ;
    input filter_data_18__0 ;
    input filter_data_19__31 ;
    input filter_data_19__30 ;
    input filter_data_19__29 ;
    input filter_data_19__28 ;
    input filter_data_19__27 ;
    input filter_data_19__26 ;
    input filter_data_19__25 ;
    input filter_data_19__24 ;
    input filter_data_19__23 ;
    input filter_data_19__22 ;
    input filter_data_19__21 ;
    input filter_data_19__20 ;
    input filter_data_19__19 ;
    input filter_data_19__18 ;
    input filter_data_19__17 ;
    input filter_data_19__16 ;
    input filter_data_19__15 ;
    input filter_data_19__14 ;
    input filter_data_19__13 ;
    input filter_data_19__12 ;
    input filter_data_19__11 ;
    input filter_data_19__10 ;
    input filter_data_19__9 ;
    input filter_data_19__8 ;
    input filter_data_19__7 ;
    input filter_data_19__6 ;
    input filter_data_19__5 ;
    input filter_data_19__4 ;
    input filter_data_19__3 ;
    input filter_data_19__2 ;
    input filter_data_19__1 ;
    input filter_data_19__0 ;
    input filter_data_20__31 ;
    input filter_data_20__30 ;
    input filter_data_20__29 ;
    input filter_data_20__28 ;
    input filter_data_20__27 ;
    input filter_data_20__26 ;
    input filter_data_20__25 ;
    input filter_data_20__24 ;
    input filter_data_20__23 ;
    input filter_data_20__22 ;
    input filter_data_20__21 ;
    input filter_data_20__20 ;
    input filter_data_20__19 ;
    input filter_data_20__18 ;
    input filter_data_20__17 ;
    input filter_data_20__16 ;
    input filter_data_20__15 ;
    input filter_data_20__14 ;
    input filter_data_20__13 ;
    input filter_data_20__12 ;
    input filter_data_20__11 ;
    input filter_data_20__10 ;
    input filter_data_20__9 ;
    input filter_data_20__8 ;
    input filter_data_20__7 ;
    input filter_data_20__6 ;
    input filter_data_20__5 ;
    input filter_data_20__4 ;
    input filter_data_20__3 ;
    input filter_data_20__2 ;
    input filter_data_20__1 ;
    input filter_data_20__0 ;
    input filter_data_21__31 ;
    input filter_data_21__30 ;
    input filter_data_21__29 ;
    input filter_data_21__28 ;
    input filter_data_21__27 ;
    input filter_data_21__26 ;
    input filter_data_21__25 ;
    input filter_data_21__24 ;
    input filter_data_21__23 ;
    input filter_data_21__22 ;
    input filter_data_21__21 ;
    input filter_data_21__20 ;
    input filter_data_21__19 ;
    input filter_data_21__18 ;
    input filter_data_21__17 ;
    input filter_data_21__16 ;
    input filter_data_21__15 ;
    input filter_data_21__14 ;
    input filter_data_21__13 ;
    input filter_data_21__12 ;
    input filter_data_21__11 ;
    input filter_data_21__10 ;
    input filter_data_21__9 ;
    input filter_data_21__8 ;
    input filter_data_21__7 ;
    input filter_data_21__6 ;
    input filter_data_21__5 ;
    input filter_data_21__4 ;
    input filter_data_21__3 ;
    input filter_data_21__2 ;
    input filter_data_21__1 ;
    input filter_data_21__0 ;
    input filter_data_22__31 ;
    input filter_data_22__30 ;
    input filter_data_22__29 ;
    input filter_data_22__28 ;
    input filter_data_22__27 ;
    input filter_data_22__26 ;
    input filter_data_22__25 ;
    input filter_data_22__24 ;
    input filter_data_22__23 ;
    input filter_data_22__22 ;
    input filter_data_22__21 ;
    input filter_data_22__20 ;
    input filter_data_22__19 ;
    input filter_data_22__18 ;
    input filter_data_22__17 ;
    input filter_data_22__16 ;
    input filter_data_22__15 ;
    input filter_data_22__14 ;
    input filter_data_22__13 ;
    input filter_data_22__12 ;
    input filter_data_22__11 ;
    input filter_data_22__10 ;
    input filter_data_22__9 ;
    input filter_data_22__8 ;
    input filter_data_22__7 ;
    input filter_data_22__6 ;
    input filter_data_22__5 ;
    input filter_data_22__4 ;
    input filter_data_22__3 ;
    input filter_data_22__2 ;
    input filter_data_22__1 ;
    input filter_data_22__0 ;
    input filter_data_23__31 ;
    input filter_data_23__30 ;
    input filter_data_23__29 ;
    input filter_data_23__28 ;
    input filter_data_23__27 ;
    input filter_data_23__26 ;
    input filter_data_23__25 ;
    input filter_data_23__24 ;
    input filter_data_23__23 ;
    input filter_data_23__22 ;
    input filter_data_23__21 ;
    input filter_data_23__20 ;
    input filter_data_23__19 ;
    input filter_data_23__18 ;
    input filter_data_23__17 ;
    input filter_data_23__16 ;
    input filter_data_23__15 ;
    input filter_data_23__14 ;
    input filter_data_23__13 ;
    input filter_data_23__12 ;
    input filter_data_23__11 ;
    input filter_data_23__10 ;
    input filter_data_23__9 ;
    input filter_data_23__8 ;
    input filter_data_23__7 ;
    input filter_data_23__6 ;
    input filter_data_23__5 ;
    input filter_data_23__4 ;
    input filter_data_23__3 ;
    input filter_data_23__2 ;
    input filter_data_23__1 ;
    input filter_data_23__0 ;
    input filter_data_24__31 ;
    input filter_data_24__30 ;
    input filter_data_24__29 ;
    input filter_data_24__28 ;
    input filter_data_24__27 ;
    input filter_data_24__26 ;
    input filter_data_24__25 ;
    input filter_data_24__24 ;
    input filter_data_24__23 ;
    input filter_data_24__22 ;
    input filter_data_24__21 ;
    input filter_data_24__20 ;
    input filter_data_24__19 ;
    input filter_data_24__18 ;
    input filter_data_24__17 ;
    input filter_data_24__16 ;
    input filter_data_24__15 ;
    input filter_data_24__14 ;
    input filter_data_24__13 ;
    input filter_data_24__12 ;
    input filter_data_24__11 ;
    input filter_data_24__10 ;
    input filter_data_24__9 ;
    input filter_data_24__8 ;
    input filter_data_24__7 ;
    input filter_data_24__6 ;
    input filter_data_24__5 ;
    input filter_data_24__4 ;
    input filter_data_24__3 ;
    input filter_data_24__2 ;
    input filter_data_24__1 ;
    input filter_data_24__0 ;
    input filter_size ;
    output ordered_img_data_0__31 ;
    output ordered_img_data_0__30 ;
    output ordered_img_data_0__29 ;
    output ordered_img_data_0__28 ;
    output ordered_img_data_0__27 ;
    output ordered_img_data_0__26 ;
    output ordered_img_data_0__25 ;
    output ordered_img_data_0__24 ;
    output ordered_img_data_0__23 ;
    output ordered_img_data_0__22 ;
    output ordered_img_data_0__21 ;
    output ordered_img_data_0__20 ;
    output ordered_img_data_0__19 ;
    output ordered_img_data_0__18 ;
    output ordered_img_data_0__17 ;
    output ordered_img_data_0__16 ;
    output ordered_img_data_0__15 ;
    output ordered_img_data_0__14 ;
    output ordered_img_data_0__13 ;
    output ordered_img_data_0__12 ;
    output ordered_img_data_0__11 ;
    output ordered_img_data_0__10 ;
    output ordered_img_data_0__9 ;
    output ordered_img_data_0__8 ;
    output ordered_img_data_0__7 ;
    output ordered_img_data_0__6 ;
    output ordered_img_data_0__5 ;
    output ordered_img_data_0__4 ;
    output ordered_img_data_0__3 ;
    output ordered_img_data_0__2 ;
    output ordered_img_data_0__1 ;
    output ordered_img_data_0__0 ;
    output ordered_img_data_1__31 ;
    output ordered_img_data_1__30 ;
    output ordered_img_data_1__29 ;
    output ordered_img_data_1__28 ;
    output ordered_img_data_1__27 ;
    output ordered_img_data_1__26 ;
    output ordered_img_data_1__25 ;
    output ordered_img_data_1__24 ;
    output ordered_img_data_1__23 ;
    output ordered_img_data_1__22 ;
    output ordered_img_data_1__21 ;
    output ordered_img_data_1__20 ;
    output ordered_img_data_1__19 ;
    output ordered_img_data_1__18 ;
    output ordered_img_data_1__17 ;
    output ordered_img_data_1__16 ;
    output ordered_img_data_1__15 ;
    output ordered_img_data_1__14 ;
    output ordered_img_data_1__13 ;
    output ordered_img_data_1__12 ;
    output ordered_img_data_1__11 ;
    output ordered_img_data_1__10 ;
    output ordered_img_data_1__9 ;
    output ordered_img_data_1__8 ;
    output ordered_img_data_1__7 ;
    output ordered_img_data_1__6 ;
    output ordered_img_data_1__5 ;
    output ordered_img_data_1__4 ;
    output ordered_img_data_1__3 ;
    output ordered_img_data_1__2 ;
    output ordered_img_data_1__1 ;
    output ordered_img_data_1__0 ;
    output ordered_img_data_2__31 ;
    output ordered_img_data_2__30 ;
    output ordered_img_data_2__29 ;
    output ordered_img_data_2__28 ;
    output ordered_img_data_2__27 ;
    output ordered_img_data_2__26 ;
    output ordered_img_data_2__25 ;
    output ordered_img_data_2__24 ;
    output ordered_img_data_2__23 ;
    output ordered_img_data_2__22 ;
    output ordered_img_data_2__21 ;
    output ordered_img_data_2__20 ;
    output ordered_img_data_2__19 ;
    output ordered_img_data_2__18 ;
    output ordered_img_data_2__17 ;
    output ordered_img_data_2__16 ;
    output ordered_img_data_2__15 ;
    output ordered_img_data_2__14 ;
    output ordered_img_data_2__13 ;
    output ordered_img_data_2__12 ;
    output ordered_img_data_2__11 ;
    output ordered_img_data_2__10 ;
    output ordered_img_data_2__9 ;
    output ordered_img_data_2__8 ;
    output ordered_img_data_2__7 ;
    output ordered_img_data_2__6 ;
    output ordered_img_data_2__5 ;
    output ordered_img_data_2__4 ;
    output ordered_img_data_2__3 ;
    output ordered_img_data_2__2 ;
    output ordered_img_data_2__1 ;
    output ordered_img_data_2__0 ;
    output ordered_img_data_3__31 ;
    output ordered_img_data_3__30 ;
    output ordered_img_data_3__29 ;
    output ordered_img_data_3__28 ;
    output ordered_img_data_3__27 ;
    output ordered_img_data_3__26 ;
    output ordered_img_data_3__25 ;
    output ordered_img_data_3__24 ;
    output ordered_img_data_3__23 ;
    output ordered_img_data_3__22 ;
    output ordered_img_data_3__21 ;
    output ordered_img_data_3__20 ;
    output ordered_img_data_3__19 ;
    output ordered_img_data_3__18 ;
    output ordered_img_data_3__17 ;
    output ordered_img_data_3__16 ;
    output ordered_img_data_3__15 ;
    output ordered_img_data_3__14 ;
    output ordered_img_data_3__13 ;
    output ordered_img_data_3__12 ;
    output ordered_img_data_3__11 ;
    output ordered_img_data_3__10 ;
    output ordered_img_data_3__9 ;
    output ordered_img_data_3__8 ;
    output ordered_img_data_3__7 ;
    output ordered_img_data_3__6 ;
    output ordered_img_data_3__5 ;
    output ordered_img_data_3__4 ;
    output ordered_img_data_3__3 ;
    output ordered_img_data_3__2 ;
    output ordered_img_data_3__1 ;
    output ordered_img_data_3__0 ;
    output ordered_img_data_4__31 ;
    output ordered_img_data_4__30 ;
    output ordered_img_data_4__29 ;
    output ordered_img_data_4__28 ;
    output ordered_img_data_4__27 ;
    output ordered_img_data_4__26 ;
    output ordered_img_data_4__25 ;
    output ordered_img_data_4__24 ;
    output ordered_img_data_4__23 ;
    output ordered_img_data_4__22 ;
    output ordered_img_data_4__21 ;
    output ordered_img_data_4__20 ;
    output ordered_img_data_4__19 ;
    output ordered_img_data_4__18 ;
    output ordered_img_data_4__17 ;
    output ordered_img_data_4__16 ;
    output ordered_img_data_4__15 ;
    output ordered_img_data_4__14 ;
    output ordered_img_data_4__13 ;
    output ordered_img_data_4__12 ;
    output ordered_img_data_4__11 ;
    output ordered_img_data_4__10 ;
    output ordered_img_data_4__9 ;
    output ordered_img_data_4__8 ;
    output ordered_img_data_4__7 ;
    output ordered_img_data_4__6 ;
    output ordered_img_data_4__5 ;
    output ordered_img_data_4__4 ;
    output ordered_img_data_4__3 ;
    output ordered_img_data_4__2 ;
    output ordered_img_data_4__1 ;
    output ordered_img_data_4__0 ;
    output ordered_img_data_5__31 ;
    output ordered_img_data_5__30 ;
    output ordered_img_data_5__29 ;
    output ordered_img_data_5__28 ;
    output ordered_img_data_5__27 ;
    output ordered_img_data_5__26 ;
    output ordered_img_data_5__25 ;
    output ordered_img_data_5__24 ;
    output ordered_img_data_5__23 ;
    output ordered_img_data_5__22 ;
    output ordered_img_data_5__21 ;
    output ordered_img_data_5__20 ;
    output ordered_img_data_5__19 ;
    output ordered_img_data_5__18 ;
    output ordered_img_data_5__17 ;
    output ordered_img_data_5__16 ;
    output ordered_img_data_5__15 ;
    output ordered_img_data_5__14 ;
    output ordered_img_data_5__13 ;
    output ordered_img_data_5__12 ;
    output ordered_img_data_5__11 ;
    output ordered_img_data_5__10 ;
    output ordered_img_data_5__9 ;
    output ordered_img_data_5__8 ;
    output ordered_img_data_5__7 ;
    output ordered_img_data_5__6 ;
    output ordered_img_data_5__5 ;
    output ordered_img_data_5__4 ;
    output ordered_img_data_5__3 ;
    output ordered_img_data_5__2 ;
    output ordered_img_data_5__1 ;
    output ordered_img_data_5__0 ;
    output ordered_img_data_6__31 ;
    output ordered_img_data_6__30 ;
    output ordered_img_data_6__29 ;
    output ordered_img_data_6__28 ;
    output ordered_img_data_6__27 ;
    output ordered_img_data_6__26 ;
    output ordered_img_data_6__25 ;
    output ordered_img_data_6__24 ;
    output ordered_img_data_6__23 ;
    output ordered_img_data_6__22 ;
    output ordered_img_data_6__21 ;
    output ordered_img_data_6__20 ;
    output ordered_img_data_6__19 ;
    output ordered_img_data_6__18 ;
    output ordered_img_data_6__17 ;
    output ordered_img_data_6__16 ;
    output ordered_img_data_6__15 ;
    output ordered_img_data_6__14 ;
    output ordered_img_data_6__13 ;
    output ordered_img_data_6__12 ;
    output ordered_img_data_6__11 ;
    output ordered_img_data_6__10 ;
    output ordered_img_data_6__9 ;
    output ordered_img_data_6__8 ;
    output ordered_img_data_6__7 ;
    output ordered_img_data_6__6 ;
    output ordered_img_data_6__5 ;
    output ordered_img_data_6__4 ;
    output ordered_img_data_6__3 ;
    output ordered_img_data_6__2 ;
    output ordered_img_data_6__1 ;
    output ordered_img_data_6__0 ;
    output ordered_img_data_7__31 ;
    output ordered_img_data_7__30 ;
    output ordered_img_data_7__29 ;
    output ordered_img_data_7__28 ;
    output ordered_img_data_7__27 ;
    output ordered_img_data_7__26 ;
    output ordered_img_data_7__25 ;
    output ordered_img_data_7__24 ;
    output ordered_img_data_7__23 ;
    output ordered_img_data_7__22 ;
    output ordered_img_data_7__21 ;
    output ordered_img_data_7__20 ;
    output ordered_img_data_7__19 ;
    output ordered_img_data_7__18 ;
    output ordered_img_data_7__17 ;
    output ordered_img_data_7__16 ;
    output ordered_img_data_7__15 ;
    output ordered_img_data_7__14 ;
    output ordered_img_data_7__13 ;
    output ordered_img_data_7__12 ;
    output ordered_img_data_7__11 ;
    output ordered_img_data_7__10 ;
    output ordered_img_data_7__9 ;
    output ordered_img_data_7__8 ;
    output ordered_img_data_7__7 ;
    output ordered_img_data_7__6 ;
    output ordered_img_data_7__5 ;
    output ordered_img_data_7__4 ;
    output ordered_img_data_7__3 ;
    output ordered_img_data_7__2 ;
    output ordered_img_data_7__1 ;
    output ordered_img_data_7__0 ;
    output ordered_img_data_8__31 ;
    output ordered_img_data_8__30 ;
    output ordered_img_data_8__29 ;
    output ordered_img_data_8__28 ;
    output ordered_img_data_8__27 ;
    output ordered_img_data_8__26 ;
    output ordered_img_data_8__25 ;
    output ordered_img_data_8__24 ;
    output ordered_img_data_8__23 ;
    output ordered_img_data_8__22 ;
    output ordered_img_data_8__21 ;
    output ordered_img_data_8__20 ;
    output ordered_img_data_8__19 ;
    output ordered_img_data_8__18 ;
    output ordered_img_data_8__17 ;
    output ordered_img_data_8__16 ;
    output ordered_img_data_8__15 ;
    output ordered_img_data_8__14 ;
    output ordered_img_data_8__13 ;
    output ordered_img_data_8__12 ;
    output ordered_img_data_8__11 ;
    output ordered_img_data_8__10 ;
    output ordered_img_data_8__9 ;
    output ordered_img_data_8__8 ;
    output ordered_img_data_8__7 ;
    output ordered_img_data_8__6 ;
    output ordered_img_data_8__5 ;
    output ordered_img_data_8__4 ;
    output ordered_img_data_8__3 ;
    output ordered_img_data_8__2 ;
    output ordered_img_data_8__1 ;
    output ordered_img_data_8__0 ;
    output ordered_img_data_9__31 ;
    output ordered_img_data_9__30 ;
    output ordered_img_data_9__29 ;
    output ordered_img_data_9__28 ;
    output ordered_img_data_9__27 ;
    output ordered_img_data_9__26 ;
    output ordered_img_data_9__25 ;
    output ordered_img_data_9__24 ;
    output ordered_img_data_9__23 ;
    output ordered_img_data_9__22 ;
    output ordered_img_data_9__21 ;
    output ordered_img_data_9__20 ;
    output ordered_img_data_9__19 ;
    output ordered_img_data_9__18 ;
    output ordered_img_data_9__17 ;
    output ordered_img_data_9__16 ;
    output ordered_img_data_9__15 ;
    output ordered_img_data_9__14 ;
    output ordered_img_data_9__13 ;
    output ordered_img_data_9__12 ;
    output ordered_img_data_9__11 ;
    output ordered_img_data_9__10 ;
    output ordered_img_data_9__9 ;
    output ordered_img_data_9__8 ;
    output ordered_img_data_9__7 ;
    output ordered_img_data_9__6 ;
    output ordered_img_data_9__5 ;
    output ordered_img_data_9__4 ;
    output ordered_img_data_9__3 ;
    output ordered_img_data_9__2 ;
    output ordered_img_data_9__1 ;
    output ordered_img_data_9__0 ;
    output ordered_img_data_10__31 ;
    output ordered_img_data_10__30 ;
    output ordered_img_data_10__29 ;
    output ordered_img_data_10__28 ;
    output ordered_img_data_10__27 ;
    output ordered_img_data_10__26 ;
    output ordered_img_data_10__25 ;
    output ordered_img_data_10__24 ;
    output ordered_img_data_10__23 ;
    output ordered_img_data_10__22 ;
    output ordered_img_data_10__21 ;
    output ordered_img_data_10__20 ;
    output ordered_img_data_10__19 ;
    output ordered_img_data_10__18 ;
    output ordered_img_data_10__17 ;
    output ordered_img_data_10__16 ;
    output ordered_img_data_10__15 ;
    output ordered_img_data_10__14 ;
    output ordered_img_data_10__13 ;
    output ordered_img_data_10__12 ;
    output ordered_img_data_10__11 ;
    output ordered_img_data_10__10 ;
    output ordered_img_data_10__9 ;
    output ordered_img_data_10__8 ;
    output ordered_img_data_10__7 ;
    output ordered_img_data_10__6 ;
    output ordered_img_data_10__5 ;
    output ordered_img_data_10__4 ;
    output ordered_img_data_10__3 ;
    output ordered_img_data_10__2 ;
    output ordered_img_data_10__1 ;
    output ordered_img_data_10__0 ;
    output ordered_img_data_11__31 ;
    output ordered_img_data_11__30 ;
    output ordered_img_data_11__29 ;
    output ordered_img_data_11__28 ;
    output ordered_img_data_11__27 ;
    output ordered_img_data_11__26 ;
    output ordered_img_data_11__25 ;
    output ordered_img_data_11__24 ;
    output ordered_img_data_11__23 ;
    output ordered_img_data_11__22 ;
    output ordered_img_data_11__21 ;
    output ordered_img_data_11__20 ;
    output ordered_img_data_11__19 ;
    output ordered_img_data_11__18 ;
    output ordered_img_data_11__17 ;
    output ordered_img_data_11__16 ;
    output ordered_img_data_11__15 ;
    output ordered_img_data_11__14 ;
    output ordered_img_data_11__13 ;
    output ordered_img_data_11__12 ;
    output ordered_img_data_11__11 ;
    output ordered_img_data_11__10 ;
    output ordered_img_data_11__9 ;
    output ordered_img_data_11__8 ;
    output ordered_img_data_11__7 ;
    output ordered_img_data_11__6 ;
    output ordered_img_data_11__5 ;
    output ordered_img_data_11__4 ;
    output ordered_img_data_11__3 ;
    output ordered_img_data_11__2 ;
    output ordered_img_data_11__1 ;
    output ordered_img_data_11__0 ;
    output ordered_img_data_12__31 ;
    output ordered_img_data_12__30 ;
    output ordered_img_data_12__29 ;
    output ordered_img_data_12__28 ;
    output ordered_img_data_12__27 ;
    output ordered_img_data_12__26 ;
    output ordered_img_data_12__25 ;
    output ordered_img_data_12__24 ;
    output ordered_img_data_12__23 ;
    output ordered_img_data_12__22 ;
    output ordered_img_data_12__21 ;
    output ordered_img_data_12__20 ;
    output ordered_img_data_12__19 ;
    output ordered_img_data_12__18 ;
    output ordered_img_data_12__17 ;
    output ordered_img_data_12__16 ;
    output ordered_img_data_12__15 ;
    output ordered_img_data_12__14 ;
    output ordered_img_data_12__13 ;
    output ordered_img_data_12__12 ;
    output ordered_img_data_12__11 ;
    output ordered_img_data_12__10 ;
    output ordered_img_data_12__9 ;
    output ordered_img_data_12__8 ;
    output ordered_img_data_12__7 ;
    output ordered_img_data_12__6 ;
    output ordered_img_data_12__5 ;
    output ordered_img_data_12__4 ;
    output ordered_img_data_12__3 ;
    output ordered_img_data_12__2 ;
    output ordered_img_data_12__1 ;
    output ordered_img_data_12__0 ;
    output ordered_img_data_13__31 ;
    output ordered_img_data_13__30 ;
    output ordered_img_data_13__29 ;
    output ordered_img_data_13__28 ;
    output ordered_img_data_13__27 ;
    output ordered_img_data_13__26 ;
    output ordered_img_data_13__25 ;
    output ordered_img_data_13__24 ;
    output ordered_img_data_13__23 ;
    output ordered_img_data_13__22 ;
    output ordered_img_data_13__21 ;
    output ordered_img_data_13__20 ;
    output ordered_img_data_13__19 ;
    output ordered_img_data_13__18 ;
    output ordered_img_data_13__17 ;
    output ordered_img_data_13__16 ;
    output ordered_img_data_13__15 ;
    output ordered_img_data_13__14 ;
    output ordered_img_data_13__13 ;
    output ordered_img_data_13__12 ;
    output ordered_img_data_13__11 ;
    output ordered_img_data_13__10 ;
    output ordered_img_data_13__9 ;
    output ordered_img_data_13__8 ;
    output ordered_img_data_13__7 ;
    output ordered_img_data_13__6 ;
    output ordered_img_data_13__5 ;
    output ordered_img_data_13__4 ;
    output ordered_img_data_13__3 ;
    output ordered_img_data_13__2 ;
    output ordered_img_data_13__1 ;
    output ordered_img_data_13__0 ;
    output ordered_img_data_14__31 ;
    output ordered_img_data_14__30 ;
    output ordered_img_data_14__29 ;
    output ordered_img_data_14__28 ;
    output ordered_img_data_14__27 ;
    output ordered_img_data_14__26 ;
    output ordered_img_data_14__25 ;
    output ordered_img_data_14__24 ;
    output ordered_img_data_14__23 ;
    output ordered_img_data_14__22 ;
    output ordered_img_data_14__21 ;
    output ordered_img_data_14__20 ;
    output ordered_img_data_14__19 ;
    output ordered_img_data_14__18 ;
    output ordered_img_data_14__17 ;
    output ordered_img_data_14__16 ;
    output ordered_img_data_14__15 ;
    output ordered_img_data_14__14 ;
    output ordered_img_data_14__13 ;
    output ordered_img_data_14__12 ;
    output ordered_img_data_14__11 ;
    output ordered_img_data_14__10 ;
    output ordered_img_data_14__9 ;
    output ordered_img_data_14__8 ;
    output ordered_img_data_14__7 ;
    output ordered_img_data_14__6 ;
    output ordered_img_data_14__5 ;
    output ordered_img_data_14__4 ;
    output ordered_img_data_14__3 ;
    output ordered_img_data_14__2 ;
    output ordered_img_data_14__1 ;
    output ordered_img_data_14__0 ;
    output ordered_img_data_15__31 ;
    output ordered_img_data_15__30 ;
    output ordered_img_data_15__29 ;
    output ordered_img_data_15__28 ;
    output ordered_img_data_15__27 ;
    output ordered_img_data_15__26 ;
    output ordered_img_data_15__25 ;
    output ordered_img_data_15__24 ;
    output ordered_img_data_15__23 ;
    output ordered_img_data_15__22 ;
    output ordered_img_data_15__21 ;
    output ordered_img_data_15__20 ;
    output ordered_img_data_15__19 ;
    output ordered_img_data_15__18 ;
    output ordered_img_data_15__17 ;
    output ordered_img_data_15__16 ;
    output ordered_img_data_15__15 ;
    output ordered_img_data_15__14 ;
    output ordered_img_data_15__13 ;
    output ordered_img_data_15__12 ;
    output ordered_img_data_15__11 ;
    output ordered_img_data_15__10 ;
    output ordered_img_data_15__9 ;
    output ordered_img_data_15__8 ;
    output ordered_img_data_15__7 ;
    output ordered_img_data_15__6 ;
    output ordered_img_data_15__5 ;
    output ordered_img_data_15__4 ;
    output ordered_img_data_15__3 ;
    output ordered_img_data_15__2 ;
    output ordered_img_data_15__1 ;
    output ordered_img_data_15__0 ;
    output ordered_img_data_16__31 ;
    output ordered_img_data_16__30 ;
    output ordered_img_data_16__29 ;
    output ordered_img_data_16__28 ;
    output ordered_img_data_16__27 ;
    output ordered_img_data_16__26 ;
    output ordered_img_data_16__25 ;
    output ordered_img_data_16__24 ;
    output ordered_img_data_16__23 ;
    output ordered_img_data_16__22 ;
    output ordered_img_data_16__21 ;
    output ordered_img_data_16__20 ;
    output ordered_img_data_16__19 ;
    output ordered_img_data_16__18 ;
    output ordered_img_data_16__17 ;
    output ordered_img_data_16__16 ;
    output ordered_img_data_16__15 ;
    output ordered_img_data_16__14 ;
    output ordered_img_data_16__13 ;
    output ordered_img_data_16__12 ;
    output ordered_img_data_16__11 ;
    output ordered_img_data_16__10 ;
    output ordered_img_data_16__9 ;
    output ordered_img_data_16__8 ;
    output ordered_img_data_16__7 ;
    output ordered_img_data_16__6 ;
    output ordered_img_data_16__5 ;
    output ordered_img_data_16__4 ;
    output ordered_img_data_16__3 ;
    output ordered_img_data_16__2 ;
    output ordered_img_data_16__1 ;
    output ordered_img_data_16__0 ;
    output ordered_img_data_17__31 ;
    output ordered_img_data_17__30 ;
    output ordered_img_data_17__29 ;
    output ordered_img_data_17__28 ;
    output ordered_img_data_17__27 ;
    output ordered_img_data_17__26 ;
    output ordered_img_data_17__25 ;
    output ordered_img_data_17__24 ;
    output ordered_img_data_17__23 ;
    output ordered_img_data_17__22 ;
    output ordered_img_data_17__21 ;
    output ordered_img_data_17__20 ;
    output ordered_img_data_17__19 ;
    output ordered_img_data_17__18 ;
    output ordered_img_data_17__17 ;
    output ordered_img_data_17__16 ;
    output ordered_img_data_17__15 ;
    output ordered_img_data_17__14 ;
    output ordered_img_data_17__13 ;
    output ordered_img_data_17__12 ;
    output ordered_img_data_17__11 ;
    output ordered_img_data_17__10 ;
    output ordered_img_data_17__9 ;
    output ordered_img_data_17__8 ;
    output ordered_img_data_17__7 ;
    output ordered_img_data_17__6 ;
    output ordered_img_data_17__5 ;
    output ordered_img_data_17__4 ;
    output ordered_img_data_17__3 ;
    output ordered_img_data_17__2 ;
    output ordered_img_data_17__1 ;
    output ordered_img_data_17__0 ;
    output ordered_img_data_18__31 ;
    output ordered_img_data_18__30 ;
    output ordered_img_data_18__29 ;
    output ordered_img_data_18__28 ;
    output ordered_img_data_18__27 ;
    output ordered_img_data_18__26 ;
    output ordered_img_data_18__25 ;
    output ordered_img_data_18__24 ;
    output ordered_img_data_18__23 ;
    output ordered_img_data_18__22 ;
    output ordered_img_data_18__21 ;
    output ordered_img_data_18__20 ;
    output ordered_img_data_18__19 ;
    output ordered_img_data_18__18 ;
    output ordered_img_data_18__17 ;
    output ordered_img_data_18__16 ;
    output ordered_img_data_18__15 ;
    output ordered_img_data_18__14 ;
    output ordered_img_data_18__13 ;
    output ordered_img_data_18__12 ;
    output ordered_img_data_18__11 ;
    output ordered_img_data_18__10 ;
    output ordered_img_data_18__9 ;
    output ordered_img_data_18__8 ;
    output ordered_img_data_18__7 ;
    output ordered_img_data_18__6 ;
    output ordered_img_data_18__5 ;
    output ordered_img_data_18__4 ;
    output ordered_img_data_18__3 ;
    output ordered_img_data_18__2 ;
    output ordered_img_data_18__1 ;
    output ordered_img_data_18__0 ;
    output ordered_img_data_19__31 ;
    output ordered_img_data_19__30 ;
    output ordered_img_data_19__29 ;
    output ordered_img_data_19__28 ;
    output ordered_img_data_19__27 ;
    output ordered_img_data_19__26 ;
    output ordered_img_data_19__25 ;
    output ordered_img_data_19__24 ;
    output ordered_img_data_19__23 ;
    output ordered_img_data_19__22 ;
    output ordered_img_data_19__21 ;
    output ordered_img_data_19__20 ;
    output ordered_img_data_19__19 ;
    output ordered_img_data_19__18 ;
    output ordered_img_data_19__17 ;
    output ordered_img_data_19__16 ;
    output ordered_img_data_19__15 ;
    output ordered_img_data_19__14 ;
    output ordered_img_data_19__13 ;
    output ordered_img_data_19__12 ;
    output ordered_img_data_19__11 ;
    output ordered_img_data_19__10 ;
    output ordered_img_data_19__9 ;
    output ordered_img_data_19__8 ;
    output ordered_img_data_19__7 ;
    output ordered_img_data_19__6 ;
    output ordered_img_data_19__5 ;
    output ordered_img_data_19__4 ;
    output ordered_img_data_19__3 ;
    output ordered_img_data_19__2 ;
    output ordered_img_data_19__1 ;
    output ordered_img_data_19__0 ;
    output ordered_img_data_20__31 ;
    output ordered_img_data_20__30 ;
    output ordered_img_data_20__29 ;
    output ordered_img_data_20__28 ;
    output ordered_img_data_20__27 ;
    output ordered_img_data_20__26 ;
    output ordered_img_data_20__25 ;
    output ordered_img_data_20__24 ;
    output ordered_img_data_20__23 ;
    output ordered_img_data_20__22 ;
    output ordered_img_data_20__21 ;
    output ordered_img_data_20__20 ;
    output ordered_img_data_20__19 ;
    output ordered_img_data_20__18 ;
    output ordered_img_data_20__17 ;
    output ordered_img_data_20__16 ;
    output ordered_img_data_20__15 ;
    output ordered_img_data_20__14 ;
    output ordered_img_data_20__13 ;
    output ordered_img_data_20__12 ;
    output ordered_img_data_20__11 ;
    output ordered_img_data_20__10 ;
    output ordered_img_data_20__9 ;
    output ordered_img_data_20__8 ;
    output ordered_img_data_20__7 ;
    output ordered_img_data_20__6 ;
    output ordered_img_data_20__5 ;
    output ordered_img_data_20__4 ;
    output ordered_img_data_20__3 ;
    output ordered_img_data_20__2 ;
    output ordered_img_data_20__1 ;
    output ordered_img_data_20__0 ;
    output ordered_img_data_21__31 ;
    output ordered_img_data_21__30 ;
    output ordered_img_data_21__29 ;
    output ordered_img_data_21__28 ;
    output ordered_img_data_21__27 ;
    output ordered_img_data_21__26 ;
    output ordered_img_data_21__25 ;
    output ordered_img_data_21__24 ;
    output ordered_img_data_21__23 ;
    output ordered_img_data_21__22 ;
    output ordered_img_data_21__21 ;
    output ordered_img_data_21__20 ;
    output ordered_img_data_21__19 ;
    output ordered_img_data_21__18 ;
    output ordered_img_data_21__17 ;
    output ordered_img_data_21__16 ;
    output ordered_img_data_21__15 ;
    output ordered_img_data_21__14 ;
    output ordered_img_data_21__13 ;
    output ordered_img_data_21__12 ;
    output ordered_img_data_21__11 ;
    output ordered_img_data_21__10 ;
    output ordered_img_data_21__9 ;
    output ordered_img_data_21__8 ;
    output ordered_img_data_21__7 ;
    output ordered_img_data_21__6 ;
    output ordered_img_data_21__5 ;
    output ordered_img_data_21__4 ;
    output ordered_img_data_21__3 ;
    output ordered_img_data_21__2 ;
    output ordered_img_data_21__1 ;
    output ordered_img_data_21__0 ;
    output ordered_img_data_22__31 ;
    output ordered_img_data_22__30 ;
    output ordered_img_data_22__29 ;
    output ordered_img_data_22__28 ;
    output ordered_img_data_22__27 ;
    output ordered_img_data_22__26 ;
    output ordered_img_data_22__25 ;
    output ordered_img_data_22__24 ;
    output ordered_img_data_22__23 ;
    output ordered_img_data_22__22 ;
    output ordered_img_data_22__21 ;
    output ordered_img_data_22__20 ;
    output ordered_img_data_22__19 ;
    output ordered_img_data_22__18 ;
    output ordered_img_data_22__17 ;
    output ordered_img_data_22__16 ;
    output ordered_img_data_22__15 ;
    output ordered_img_data_22__14 ;
    output ordered_img_data_22__13 ;
    output ordered_img_data_22__12 ;
    output ordered_img_data_22__11 ;
    output ordered_img_data_22__10 ;
    output ordered_img_data_22__9 ;
    output ordered_img_data_22__8 ;
    output ordered_img_data_22__7 ;
    output ordered_img_data_22__6 ;
    output ordered_img_data_22__5 ;
    output ordered_img_data_22__4 ;
    output ordered_img_data_22__3 ;
    output ordered_img_data_22__2 ;
    output ordered_img_data_22__1 ;
    output ordered_img_data_22__0 ;
    output ordered_img_data_23__31 ;
    output ordered_img_data_23__30 ;
    output ordered_img_data_23__29 ;
    output ordered_img_data_23__28 ;
    output ordered_img_data_23__27 ;
    output ordered_img_data_23__26 ;
    output ordered_img_data_23__25 ;
    output ordered_img_data_23__24 ;
    output ordered_img_data_23__23 ;
    output ordered_img_data_23__22 ;
    output ordered_img_data_23__21 ;
    output ordered_img_data_23__20 ;
    output ordered_img_data_23__19 ;
    output ordered_img_data_23__18 ;
    output ordered_img_data_23__17 ;
    output ordered_img_data_23__16 ;
    output ordered_img_data_23__15 ;
    output ordered_img_data_23__14 ;
    output ordered_img_data_23__13 ;
    output ordered_img_data_23__12 ;
    output ordered_img_data_23__11 ;
    output ordered_img_data_23__10 ;
    output ordered_img_data_23__9 ;
    output ordered_img_data_23__8 ;
    output ordered_img_data_23__7 ;
    output ordered_img_data_23__6 ;
    output ordered_img_data_23__5 ;
    output ordered_img_data_23__4 ;
    output ordered_img_data_23__3 ;
    output ordered_img_data_23__2 ;
    output ordered_img_data_23__1 ;
    output ordered_img_data_23__0 ;
    output ordered_img_data_24__31 ;
    output ordered_img_data_24__30 ;
    output ordered_img_data_24__29 ;
    output ordered_img_data_24__28 ;
    output ordered_img_data_24__27 ;
    output ordered_img_data_24__26 ;
    output ordered_img_data_24__25 ;
    output ordered_img_data_24__24 ;
    output ordered_img_data_24__23 ;
    output ordered_img_data_24__22 ;
    output ordered_img_data_24__21 ;
    output ordered_img_data_24__20 ;
    output ordered_img_data_24__19 ;
    output ordered_img_data_24__18 ;
    output ordered_img_data_24__17 ;
    output ordered_img_data_24__16 ;
    output ordered_img_data_24__15 ;
    output ordered_img_data_24__14 ;
    output ordered_img_data_24__13 ;
    output ordered_img_data_24__12 ;
    output ordered_img_data_24__11 ;
    output ordered_img_data_24__10 ;
    output ordered_img_data_24__9 ;
    output ordered_img_data_24__8 ;
    output ordered_img_data_24__7 ;
    output ordered_img_data_24__6 ;
    output ordered_img_data_24__5 ;
    output ordered_img_data_24__4 ;
    output ordered_img_data_24__3 ;
    output ordered_img_data_24__2 ;
    output ordered_img_data_24__1 ;
    output ordered_img_data_24__0 ;
    output ordered_filter_data_0__31 ;
    output ordered_filter_data_0__30 ;
    output ordered_filter_data_0__29 ;
    output ordered_filter_data_0__28 ;
    output ordered_filter_data_0__27 ;
    output ordered_filter_data_0__26 ;
    output ordered_filter_data_0__25 ;
    output ordered_filter_data_0__24 ;
    output ordered_filter_data_0__23 ;
    output ordered_filter_data_0__22 ;
    output ordered_filter_data_0__21 ;
    output ordered_filter_data_0__20 ;
    output ordered_filter_data_0__19 ;
    output ordered_filter_data_0__18 ;
    output ordered_filter_data_0__17 ;
    output ordered_filter_data_0__16 ;
    output ordered_filter_data_0__15 ;
    output ordered_filter_data_0__14 ;
    output ordered_filter_data_0__13 ;
    output ordered_filter_data_0__12 ;
    output ordered_filter_data_0__11 ;
    output ordered_filter_data_0__10 ;
    output ordered_filter_data_0__9 ;
    output ordered_filter_data_0__8 ;
    output ordered_filter_data_0__7 ;
    output ordered_filter_data_0__6 ;
    output ordered_filter_data_0__5 ;
    output ordered_filter_data_0__4 ;
    output ordered_filter_data_0__3 ;
    output ordered_filter_data_0__2 ;
    output ordered_filter_data_0__1 ;
    output ordered_filter_data_0__0 ;
    output ordered_filter_data_1__31 ;
    output ordered_filter_data_1__30 ;
    output ordered_filter_data_1__29 ;
    output ordered_filter_data_1__28 ;
    output ordered_filter_data_1__27 ;
    output ordered_filter_data_1__26 ;
    output ordered_filter_data_1__25 ;
    output ordered_filter_data_1__24 ;
    output ordered_filter_data_1__23 ;
    output ordered_filter_data_1__22 ;
    output ordered_filter_data_1__21 ;
    output ordered_filter_data_1__20 ;
    output ordered_filter_data_1__19 ;
    output ordered_filter_data_1__18 ;
    output ordered_filter_data_1__17 ;
    output ordered_filter_data_1__16 ;
    output ordered_filter_data_1__15 ;
    output ordered_filter_data_1__14 ;
    output ordered_filter_data_1__13 ;
    output ordered_filter_data_1__12 ;
    output ordered_filter_data_1__11 ;
    output ordered_filter_data_1__10 ;
    output ordered_filter_data_1__9 ;
    output ordered_filter_data_1__8 ;
    output ordered_filter_data_1__7 ;
    output ordered_filter_data_1__6 ;
    output ordered_filter_data_1__5 ;
    output ordered_filter_data_1__4 ;
    output ordered_filter_data_1__3 ;
    output ordered_filter_data_1__2 ;
    output ordered_filter_data_1__1 ;
    output ordered_filter_data_1__0 ;
    output ordered_filter_data_2__31 ;
    output ordered_filter_data_2__30 ;
    output ordered_filter_data_2__29 ;
    output ordered_filter_data_2__28 ;
    output ordered_filter_data_2__27 ;
    output ordered_filter_data_2__26 ;
    output ordered_filter_data_2__25 ;
    output ordered_filter_data_2__24 ;
    output ordered_filter_data_2__23 ;
    output ordered_filter_data_2__22 ;
    output ordered_filter_data_2__21 ;
    output ordered_filter_data_2__20 ;
    output ordered_filter_data_2__19 ;
    output ordered_filter_data_2__18 ;
    output ordered_filter_data_2__17 ;
    output ordered_filter_data_2__16 ;
    output ordered_filter_data_2__15 ;
    output ordered_filter_data_2__14 ;
    output ordered_filter_data_2__13 ;
    output ordered_filter_data_2__12 ;
    output ordered_filter_data_2__11 ;
    output ordered_filter_data_2__10 ;
    output ordered_filter_data_2__9 ;
    output ordered_filter_data_2__8 ;
    output ordered_filter_data_2__7 ;
    output ordered_filter_data_2__6 ;
    output ordered_filter_data_2__5 ;
    output ordered_filter_data_2__4 ;
    output ordered_filter_data_2__3 ;
    output ordered_filter_data_2__2 ;
    output ordered_filter_data_2__1 ;
    output ordered_filter_data_2__0 ;
    output ordered_filter_data_3__31 ;
    output ordered_filter_data_3__30 ;
    output ordered_filter_data_3__29 ;
    output ordered_filter_data_3__28 ;
    output ordered_filter_data_3__27 ;
    output ordered_filter_data_3__26 ;
    output ordered_filter_data_3__25 ;
    output ordered_filter_data_3__24 ;
    output ordered_filter_data_3__23 ;
    output ordered_filter_data_3__22 ;
    output ordered_filter_data_3__21 ;
    output ordered_filter_data_3__20 ;
    output ordered_filter_data_3__19 ;
    output ordered_filter_data_3__18 ;
    output ordered_filter_data_3__17 ;
    output ordered_filter_data_3__16 ;
    output ordered_filter_data_3__15 ;
    output ordered_filter_data_3__14 ;
    output ordered_filter_data_3__13 ;
    output ordered_filter_data_3__12 ;
    output ordered_filter_data_3__11 ;
    output ordered_filter_data_3__10 ;
    output ordered_filter_data_3__9 ;
    output ordered_filter_data_3__8 ;
    output ordered_filter_data_3__7 ;
    output ordered_filter_data_3__6 ;
    output ordered_filter_data_3__5 ;
    output ordered_filter_data_3__4 ;
    output ordered_filter_data_3__3 ;
    output ordered_filter_data_3__2 ;
    output ordered_filter_data_3__1 ;
    output ordered_filter_data_3__0 ;
    output ordered_filter_data_4__31 ;
    output ordered_filter_data_4__30 ;
    output ordered_filter_data_4__29 ;
    output ordered_filter_data_4__28 ;
    output ordered_filter_data_4__27 ;
    output ordered_filter_data_4__26 ;
    output ordered_filter_data_4__25 ;
    output ordered_filter_data_4__24 ;
    output ordered_filter_data_4__23 ;
    output ordered_filter_data_4__22 ;
    output ordered_filter_data_4__21 ;
    output ordered_filter_data_4__20 ;
    output ordered_filter_data_4__19 ;
    output ordered_filter_data_4__18 ;
    output ordered_filter_data_4__17 ;
    output ordered_filter_data_4__16 ;
    output ordered_filter_data_4__15 ;
    output ordered_filter_data_4__14 ;
    output ordered_filter_data_4__13 ;
    output ordered_filter_data_4__12 ;
    output ordered_filter_data_4__11 ;
    output ordered_filter_data_4__10 ;
    output ordered_filter_data_4__9 ;
    output ordered_filter_data_4__8 ;
    output ordered_filter_data_4__7 ;
    output ordered_filter_data_4__6 ;
    output ordered_filter_data_4__5 ;
    output ordered_filter_data_4__4 ;
    output ordered_filter_data_4__3 ;
    output ordered_filter_data_4__2 ;
    output ordered_filter_data_4__1 ;
    output ordered_filter_data_4__0 ;
    output ordered_filter_data_5__31 ;
    output ordered_filter_data_5__30 ;
    output ordered_filter_data_5__29 ;
    output ordered_filter_data_5__28 ;
    output ordered_filter_data_5__27 ;
    output ordered_filter_data_5__26 ;
    output ordered_filter_data_5__25 ;
    output ordered_filter_data_5__24 ;
    output ordered_filter_data_5__23 ;
    output ordered_filter_data_5__22 ;
    output ordered_filter_data_5__21 ;
    output ordered_filter_data_5__20 ;
    output ordered_filter_data_5__19 ;
    output ordered_filter_data_5__18 ;
    output ordered_filter_data_5__17 ;
    output ordered_filter_data_5__16 ;
    output ordered_filter_data_5__15 ;
    output ordered_filter_data_5__14 ;
    output ordered_filter_data_5__13 ;
    output ordered_filter_data_5__12 ;
    output ordered_filter_data_5__11 ;
    output ordered_filter_data_5__10 ;
    output ordered_filter_data_5__9 ;
    output ordered_filter_data_5__8 ;
    output ordered_filter_data_5__7 ;
    output ordered_filter_data_5__6 ;
    output ordered_filter_data_5__5 ;
    output ordered_filter_data_5__4 ;
    output ordered_filter_data_5__3 ;
    output ordered_filter_data_5__2 ;
    output ordered_filter_data_5__1 ;
    output ordered_filter_data_5__0 ;
    output ordered_filter_data_6__31 ;
    output ordered_filter_data_6__30 ;
    output ordered_filter_data_6__29 ;
    output ordered_filter_data_6__28 ;
    output ordered_filter_data_6__27 ;
    output ordered_filter_data_6__26 ;
    output ordered_filter_data_6__25 ;
    output ordered_filter_data_6__24 ;
    output ordered_filter_data_6__23 ;
    output ordered_filter_data_6__22 ;
    output ordered_filter_data_6__21 ;
    output ordered_filter_data_6__20 ;
    output ordered_filter_data_6__19 ;
    output ordered_filter_data_6__18 ;
    output ordered_filter_data_6__17 ;
    output ordered_filter_data_6__16 ;
    output ordered_filter_data_6__15 ;
    output ordered_filter_data_6__14 ;
    output ordered_filter_data_6__13 ;
    output ordered_filter_data_6__12 ;
    output ordered_filter_data_6__11 ;
    output ordered_filter_data_6__10 ;
    output ordered_filter_data_6__9 ;
    output ordered_filter_data_6__8 ;
    output ordered_filter_data_6__7 ;
    output ordered_filter_data_6__6 ;
    output ordered_filter_data_6__5 ;
    output ordered_filter_data_6__4 ;
    output ordered_filter_data_6__3 ;
    output ordered_filter_data_6__2 ;
    output ordered_filter_data_6__1 ;
    output ordered_filter_data_6__0 ;
    output ordered_filter_data_7__31 ;
    output ordered_filter_data_7__30 ;
    output ordered_filter_data_7__29 ;
    output ordered_filter_data_7__28 ;
    output ordered_filter_data_7__27 ;
    output ordered_filter_data_7__26 ;
    output ordered_filter_data_7__25 ;
    output ordered_filter_data_7__24 ;
    output ordered_filter_data_7__23 ;
    output ordered_filter_data_7__22 ;
    output ordered_filter_data_7__21 ;
    output ordered_filter_data_7__20 ;
    output ordered_filter_data_7__19 ;
    output ordered_filter_data_7__18 ;
    output ordered_filter_data_7__17 ;
    output ordered_filter_data_7__16 ;
    output ordered_filter_data_7__15 ;
    output ordered_filter_data_7__14 ;
    output ordered_filter_data_7__13 ;
    output ordered_filter_data_7__12 ;
    output ordered_filter_data_7__11 ;
    output ordered_filter_data_7__10 ;
    output ordered_filter_data_7__9 ;
    output ordered_filter_data_7__8 ;
    output ordered_filter_data_7__7 ;
    output ordered_filter_data_7__6 ;
    output ordered_filter_data_7__5 ;
    output ordered_filter_data_7__4 ;
    output ordered_filter_data_7__3 ;
    output ordered_filter_data_7__2 ;
    output ordered_filter_data_7__1 ;
    output ordered_filter_data_7__0 ;
    output ordered_filter_data_8__31 ;
    output ordered_filter_data_8__30 ;
    output ordered_filter_data_8__29 ;
    output ordered_filter_data_8__28 ;
    output ordered_filter_data_8__27 ;
    output ordered_filter_data_8__26 ;
    output ordered_filter_data_8__25 ;
    output ordered_filter_data_8__24 ;
    output ordered_filter_data_8__23 ;
    output ordered_filter_data_8__22 ;
    output ordered_filter_data_8__21 ;
    output ordered_filter_data_8__20 ;
    output ordered_filter_data_8__19 ;
    output ordered_filter_data_8__18 ;
    output ordered_filter_data_8__17 ;
    output ordered_filter_data_8__16 ;
    output ordered_filter_data_8__15 ;
    output ordered_filter_data_8__14 ;
    output ordered_filter_data_8__13 ;
    output ordered_filter_data_8__12 ;
    output ordered_filter_data_8__11 ;
    output ordered_filter_data_8__10 ;
    output ordered_filter_data_8__9 ;
    output ordered_filter_data_8__8 ;
    output ordered_filter_data_8__7 ;
    output ordered_filter_data_8__6 ;
    output ordered_filter_data_8__5 ;
    output ordered_filter_data_8__4 ;
    output ordered_filter_data_8__3 ;
    output ordered_filter_data_8__2 ;
    output ordered_filter_data_8__1 ;
    output ordered_filter_data_8__0 ;
    output ordered_filter_data_9__31 ;
    output ordered_filter_data_9__30 ;
    output ordered_filter_data_9__29 ;
    output ordered_filter_data_9__28 ;
    output ordered_filter_data_9__27 ;
    output ordered_filter_data_9__26 ;
    output ordered_filter_data_9__25 ;
    output ordered_filter_data_9__24 ;
    output ordered_filter_data_9__23 ;
    output ordered_filter_data_9__22 ;
    output ordered_filter_data_9__21 ;
    output ordered_filter_data_9__20 ;
    output ordered_filter_data_9__19 ;
    output ordered_filter_data_9__18 ;
    output ordered_filter_data_9__17 ;
    output ordered_filter_data_9__16 ;
    output ordered_filter_data_9__15 ;
    output ordered_filter_data_9__14 ;
    output ordered_filter_data_9__13 ;
    output ordered_filter_data_9__12 ;
    output ordered_filter_data_9__11 ;
    output ordered_filter_data_9__10 ;
    output ordered_filter_data_9__9 ;
    output ordered_filter_data_9__8 ;
    output ordered_filter_data_9__7 ;
    output ordered_filter_data_9__6 ;
    output ordered_filter_data_9__5 ;
    output ordered_filter_data_9__4 ;
    output ordered_filter_data_9__3 ;
    output ordered_filter_data_9__2 ;
    output ordered_filter_data_9__1 ;
    output ordered_filter_data_9__0 ;
    output ordered_filter_data_10__31 ;
    output ordered_filter_data_10__30 ;
    output ordered_filter_data_10__29 ;
    output ordered_filter_data_10__28 ;
    output ordered_filter_data_10__27 ;
    output ordered_filter_data_10__26 ;
    output ordered_filter_data_10__25 ;
    output ordered_filter_data_10__24 ;
    output ordered_filter_data_10__23 ;
    output ordered_filter_data_10__22 ;
    output ordered_filter_data_10__21 ;
    output ordered_filter_data_10__20 ;
    output ordered_filter_data_10__19 ;
    output ordered_filter_data_10__18 ;
    output ordered_filter_data_10__17 ;
    output ordered_filter_data_10__16 ;
    output ordered_filter_data_10__15 ;
    output ordered_filter_data_10__14 ;
    output ordered_filter_data_10__13 ;
    output ordered_filter_data_10__12 ;
    output ordered_filter_data_10__11 ;
    output ordered_filter_data_10__10 ;
    output ordered_filter_data_10__9 ;
    output ordered_filter_data_10__8 ;
    output ordered_filter_data_10__7 ;
    output ordered_filter_data_10__6 ;
    output ordered_filter_data_10__5 ;
    output ordered_filter_data_10__4 ;
    output ordered_filter_data_10__3 ;
    output ordered_filter_data_10__2 ;
    output ordered_filter_data_10__1 ;
    output ordered_filter_data_10__0 ;
    output ordered_filter_data_11__31 ;
    output ordered_filter_data_11__30 ;
    output ordered_filter_data_11__29 ;
    output ordered_filter_data_11__28 ;
    output ordered_filter_data_11__27 ;
    output ordered_filter_data_11__26 ;
    output ordered_filter_data_11__25 ;
    output ordered_filter_data_11__24 ;
    output ordered_filter_data_11__23 ;
    output ordered_filter_data_11__22 ;
    output ordered_filter_data_11__21 ;
    output ordered_filter_data_11__20 ;
    output ordered_filter_data_11__19 ;
    output ordered_filter_data_11__18 ;
    output ordered_filter_data_11__17 ;
    output ordered_filter_data_11__16 ;
    output ordered_filter_data_11__15 ;
    output ordered_filter_data_11__14 ;
    output ordered_filter_data_11__13 ;
    output ordered_filter_data_11__12 ;
    output ordered_filter_data_11__11 ;
    output ordered_filter_data_11__10 ;
    output ordered_filter_data_11__9 ;
    output ordered_filter_data_11__8 ;
    output ordered_filter_data_11__7 ;
    output ordered_filter_data_11__6 ;
    output ordered_filter_data_11__5 ;
    output ordered_filter_data_11__4 ;
    output ordered_filter_data_11__3 ;
    output ordered_filter_data_11__2 ;
    output ordered_filter_data_11__1 ;
    output ordered_filter_data_11__0 ;
    output ordered_filter_data_12__31 ;
    output ordered_filter_data_12__30 ;
    output ordered_filter_data_12__29 ;
    output ordered_filter_data_12__28 ;
    output ordered_filter_data_12__27 ;
    output ordered_filter_data_12__26 ;
    output ordered_filter_data_12__25 ;
    output ordered_filter_data_12__24 ;
    output ordered_filter_data_12__23 ;
    output ordered_filter_data_12__22 ;
    output ordered_filter_data_12__21 ;
    output ordered_filter_data_12__20 ;
    output ordered_filter_data_12__19 ;
    output ordered_filter_data_12__18 ;
    output ordered_filter_data_12__17 ;
    output ordered_filter_data_12__16 ;
    output ordered_filter_data_12__15 ;
    output ordered_filter_data_12__14 ;
    output ordered_filter_data_12__13 ;
    output ordered_filter_data_12__12 ;
    output ordered_filter_data_12__11 ;
    output ordered_filter_data_12__10 ;
    output ordered_filter_data_12__9 ;
    output ordered_filter_data_12__8 ;
    output ordered_filter_data_12__7 ;
    output ordered_filter_data_12__6 ;
    output ordered_filter_data_12__5 ;
    output ordered_filter_data_12__4 ;
    output ordered_filter_data_12__3 ;
    output ordered_filter_data_12__2 ;
    output ordered_filter_data_12__1 ;
    output ordered_filter_data_12__0 ;
    output ordered_filter_data_13__31 ;
    output ordered_filter_data_13__30 ;
    output ordered_filter_data_13__29 ;
    output ordered_filter_data_13__28 ;
    output ordered_filter_data_13__27 ;
    output ordered_filter_data_13__26 ;
    output ordered_filter_data_13__25 ;
    output ordered_filter_data_13__24 ;
    output ordered_filter_data_13__23 ;
    output ordered_filter_data_13__22 ;
    output ordered_filter_data_13__21 ;
    output ordered_filter_data_13__20 ;
    output ordered_filter_data_13__19 ;
    output ordered_filter_data_13__18 ;
    output ordered_filter_data_13__17 ;
    output ordered_filter_data_13__16 ;
    output ordered_filter_data_13__15 ;
    output ordered_filter_data_13__14 ;
    output ordered_filter_data_13__13 ;
    output ordered_filter_data_13__12 ;
    output ordered_filter_data_13__11 ;
    output ordered_filter_data_13__10 ;
    output ordered_filter_data_13__9 ;
    output ordered_filter_data_13__8 ;
    output ordered_filter_data_13__7 ;
    output ordered_filter_data_13__6 ;
    output ordered_filter_data_13__5 ;
    output ordered_filter_data_13__4 ;
    output ordered_filter_data_13__3 ;
    output ordered_filter_data_13__2 ;
    output ordered_filter_data_13__1 ;
    output ordered_filter_data_13__0 ;
    output ordered_filter_data_14__31 ;
    output ordered_filter_data_14__30 ;
    output ordered_filter_data_14__29 ;
    output ordered_filter_data_14__28 ;
    output ordered_filter_data_14__27 ;
    output ordered_filter_data_14__26 ;
    output ordered_filter_data_14__25 ;
    output ordered_filter_data_14__24 ;
    output ordered_filter_data_14__23 ;
    output ordered_filter_data_14__22 ;
    output ordered_filter_data_14__21 ;
    output ordered_filter_data_14__20 ;
    output ordered_filter_data_14__19 ;
    output ordered_filter_data_14__18 ;
    output ordered_filter_data_14__17 ;
    output ordered_filter_data_14__16 ;
    output ordered_filter_data_14__15 ;
    output ordered_filter_data_14__14 ;
    output ordered_filter_data_14__13 ;
    output ordered_filter_data_14__12 ;
    output ordered_filter_data_14__11 ;
    output ordered_filter_data_14__10 ;
    output ordered_filter_data_14__9 ;
    output ordered_filter_data_14__8 ;
    output ordered_filter_data_14__7 ;
    output ordered_filter_data_14__6 ;
    output ordered_filter_data_14__5 ;
    output ordered_filter_data_14__4 ;
    output ordered_filter_data_14__3 ;
    output ordered_filter_data_14__2 ;
    output ordered_filter_data_14__1 ;
    output ordered_filter_data_14__0 ;
    output ordered_filter_data_15__31 ;
    output ordered_filter_data_15__30 ;
    output ordered_filter_data_15__29 ;
    output ordered_filter_data_15__28 ;
    output ordered_filter_data_15__27 ;
    output ordered_filter_data_15__26 ;
    output ordered_filter_data_15__25 ;
    output ordered_filter_data_15__24 ;
    output ordered_filter_data_15__23 ;
    output ordered_filter_data_15__22 ;
    output ordered_filter_data_15__21 ;
    output ordered_filter_data_15__20 ;
    output ordered_filter_data_15__19 ;
    output ordered_filter_data_15__18 ;
    output ordered_filter_data_15__17 ;
    output ordered_filter_data_15__16 ;
    output ordered_filter_data_15__15 ;
    output ordered_filter_data_15__14 ;
    output ordered_filter_data_15__13 ;
    output ordered_filter_data_15__12 ;
    output ordered_filter_data_15__11 ;
    output ordered_filter_data_15__10 ;
    output ordered_filter_data_15__9 ;
    output ordered_filter_data_15__8 ;
    output ordered_filter_data_15__7 ;
    output ordered_filter_data_15__6 ;
    output ordered_filter_data_15__5 ;
    output ordered_filter_data_15__4 ;
    output ordered_filter_data_15__3 ;
    output ordered_filter_data_15__2 ;
    output ordered_filter_data_15__1 ;
    output ordered_filter_data_15__0 ;
    output ordered_filter_data_16__31 ;
    output ordered_filter_data_16__30 ;
    output ordered_filter_data_16__29 ;
    output ordered_filter_data_16__28 ;
    output ordered_filter_data_16__27 ;
    output ordered_filter_data_16__26 ;
    output ordered_filter_data_16__25 ;
    output ordered_filter_data_16__24 ;
    output ordered_filter_data_16__23 ;
    output ordered_filter_data_16__22 ;
    output ordered_filter_data_16__21 ;
    output ordered_filter_data_16__20 ;
    output ordered_filter_data_16__19 ;
    output ordered_filter_data_16__18 ;
    output ordered_filter_data_16__17 ;
    output ordered_filter_data_16__16 ;
    output ordered_filter_data_16__15 ;
    output ordered_filter_data_16__14 ;
    output ordered_filter_data_16__13 ;
    output ordered_filter_data_16__12 ;
    output ordered_filter_data_16__11 ;
    output ordered_filter_data_16__10 ;
    output ordered_filter_data_16__9 ;
    output ordered_filter_data_16__8 ;
    output ordered_filter_data_16__7 ;
    output ordered_filter_data_16__6 ;
    output ordered_filter_data_16__5 ;
    output ordered_filter_data_16__4 ;
    output ordered_filter_data_16__3 ;
    output ordered_filter_data_16__2 ;
    output ordered_filter_data_16__1 ;
    output ordered_filter_data_16__0 ;
    output ordered_filter_data_17__31 ;
    output ordered_filter_data_17__30 ;
    output ordered_filter_data_17__29 ;
    output ordered_filter_data_17__28 ;
    output ordered_filter_data_17__27 ;
    output ordered_filter_data_17__26 ;
    output ordered_filter_data_17__25 ;
    output ordered_filter_data_17__24 ;
    output ordered_filter_data_17__23 ;
    output ordered_filter_data_17__22 ;
    output ordered_filter_data_17__21 ;
    output ordered_filter_data_17__20 ;
    output ordered_filter_data_17__19 ;
    output ordered_filter_data_17__18 ;
    output ordered_filter_data_17__17 ;
    output ordered_filter_data_17__16 ;
    output ordered_filter_data_17__15 ;
    output ordered_filter_data_17__14 ;
    output ordered_filter_data_17__13 ;
    output ordered_filter_data_17__12 ;
    output ordered_filter_data_17__11 ;
    output ordered_filter_data_17__10 ;
    output ordered_filter_data_17__9 ;
    output ordered_filter_data_17__8 ;
    output ordered_filter_data_17__7 ;
    output ordered_filter_data_17__6 ;
    output ordered_filter_data_17__5 ;
    output ordered_filter_data_17__4 ;
    output ordered_filter_data_17__3 ;
    output ordered_filter_data_17__2 ;
    output ordered_filter_data_17__1 ;
    output ordered_filter_data_17__0 ;
    output ordered_filter_data_18__31 ;
    output ordered_filter_data_18__30 ;
    output ordered_filter_data_18__29 ;
    output ordered_filter_data_18__28 ;
    output ordered_filter_data_18__27 ;
    output ordered_filter_data_18__26 ;
    output ordered_filter_data_18__25 ;
    output ordered_filter_data_18__24 ;
    output ordered_filter_data_18__23 ;
    output ordered_filter_data_18__22 ;
    output ordered_filter_data_18__21 ;
    output ordered_filter_data_18__20 ;
    output ordered_filter_data_18__19 ;
    output ordered_filter_data_18__18 ;
    output ordered_filter_data_18__17 ;
    output ordered_filter_data_18__16 ;
    output ordered_filter_data_18__15 ;
    output ordered_filter_data_18__14 ;
    output ordered_filter_data_18__13 ;
    output ordered_filter_data_18__12 ;
    output ordered_filter_data_18__11 ;
    output ordered_filter_data_18__10 ;
    output ordered_filter_data_18__9 ;
    output ordered_filter_data_18__8 ;
    output ordered_filter_data_18__7 ;
    output ordered_filter_data_18__6 ;
    output ordered_filter_data_18__5 ;
    output ordered_filter_data_18__4 ;
    output ordered_filter_data_18__3 ;
    output ordered_filter_data_18__2 ;
    output ordered_filter_data_18__1 ;
    output ordered_filter_data_18__0 ;
    output ordered_filter_data_19__31 ;
    output ordered_filter_data_19__30 ;
    output ordered_filter_data_19__29 ;
    output ordered_filter_data_19__28 ;
    output ordered_filter_data_19__27 ;
    output ordered_filter_data_19__26 ;
    output ordered_filter_data_19__25 ;
    output ordered_filter_data_19__24 ;
    output ordered_filter_data_19__23 ;
    output ordered_filter_data_19__22 ;
    output ordered_filter_data_19__21 ;
    output ordered_filter_data_19__20 ;
    output ordered_filter_data_19__19 ;
    output ordered_filter_data_19__18 ;
    output ordered_filter_data_19__17 ;
    output ordered_filter_data_19__16 ;
    output ordered_filter_data_19__15 ;
    output ordered_filter_data_19__14 ;
    output ordered_filter_data_19__13 ;
    output ordered_filter_data_19__12 ;
    output ordered_filter_data_19__11 ;
    output ordered_filter_data_19__10 ;
    output ordered_filter_data_19__9 ;
    output ordered_filter_data_19__8 ;
    output ordered_filter_data_19__7 ;
    output ordered_filter_data_19__6 ;
    output ordered_filter_data_19__5 ;
    output ordered_filter_data_19__4 ;
    output ordered_filter_data_19__3 ;
    output ordered_filter_data_19__2 ;
    output ordered_filter_data_19__1 ;
    output ordered_filter_data_19__0 ;
    output ordered_filter_data_20__31 ;
    output ordered_filter_data_20__30 ;
    output ordered_filter_data_20__29 ;
    output ordered_filter_data_20__28 ;
    output ordered_filter_data_20__27 ;
    output ordered_filter_data_20__26 ;
    output ordered_filter_data_20__25 ;
    output ordered_filter_data_20__24 ;
    output ordered_filter_data_20__23 ;
    output ordered_filter_data_20__22 ;
    output ordered_filter_data_20__21 ;
    output ordered_filter_data_20__20 ;
    output ordered_filter_data_20__19 ;
    output ordered_filter_data_20__18 ;
    output ordered_filter_data_20__17 ;
    output ordered_filter_data_20__16 ;
    output ordered_filter_data_20__15 ;
    output ordered_filter_data_20__14 ;
    output ordered_filter_data_20__13 ;
    output ordered_filter_data_20__12 ;
    output ordered_filter_data_20__11 ;
    output ordered_filter_data_20__10 ;
    output ordered_filter_data_20__9 ;
    output ordered_filter_data_20__8 ;
    output ordered_filter_data_20__7 ;
    output ordered_filter_data_20__6 ;
    output ordered_filter_data_20__5 ;
    output ordered_filter_data_20__4 ;
    output ordered_filter_data_20__3 ;
    output ordered_filter_data_20__2 ;
    output ordered_filter_data_20__1 ;
    output ordered_filter_data_20__0 ;
    output ordered_filter_data_21__31 ;
    output ordered_filter_data_21__30 ;
    output ordered_filter_data_21__29 ;
    output ordered_filter_data_21__28 ;
    output ordered_filter_data_21__27 ;
    output ordered_filter_data_21__26 ;
    output ordered_filter_data_21__25 ;
    output ordered_filter_data_21__24 ;
    output ordered_filter_data_21__23 ;
    output ordered_filter_data_21__22 ;
    output ordered_filter_data_21__21 ;
    output ordered_filter_data_21__20 ;
    output ordered_filter_data_21__19 ;
    output ordered_filter_data_21__18 ;
    output ordered_filter_data_21__17 ;
    output ordered_filter_data_21__16 ;
    output ordered_filter_data_21__15 ;
    output ordered_filter_data_21__14 ;
    output ordered_filter_data_21__13 ;
    output ordered_filter_data_21__12 ;
    output ordered_filter_data_21__11 ;
    output ordered_filter_data_21__10 ;
    output ordered_filter_data_21__9 ;
    output ordered_filter_data_21__8 ;
    output ordered_filter_data_21__7 ;
    output ordered_filter_data_21__6 ;
    output ordered_filter_data_21__5 ;
    output ordered_filter_data_21__4 ;
    output ordered_filter_data_21__3 ;
    output ordered_filter_data_21__2 ;
    output ordered_filter_data_21__1 ;
    output ordered_filter_data_21__0 ;
    output ordered_filter_data_22__31 ;
    output ordered_filter_data_22__30 ;
    output ordered_filter_data_22__29 ;
    output ordered_filter_data_22__28 ;
    output ordered_filter_data_22__27 ;
    output ordered_filter_data_22__26 ;
    output ordered_filter_data_22__25 ;
    output ordered_filter_data_22__24 ;
    output ordered_filter_data_22__23 ;
    output ordered_filter_data_22__22 ;
    output ordered_filter_data_22__21 ;
    output ordered_filter_data_22__20 ;
    output ordered_filter_data_22__19 ;
    output ordered_filter_data_22__18 ;
    output ordered_filter_data_22__17 ;
    output ordered_filter_data_22__16 ;
    output ordered_filter_data_22__15 ;
    output ordered_filter_data_22__14 ;
    output ordered_filter_data_22__13 ;
    output ordered_filter_data_22__12 ;
    output ordered_filter_data_22__11 ;
    output ordered_filter_data_22__10 ;
    output ordered_filter_data_22__9 ;
    output ordered_filter_data_22__8 ;
    output ordered_filter_data_22__7 ;
    output ordered_filter_data_22__6 ;
    output ordered_filter_data_22__5 ;
    output ordered_filter_data_22__4 ;
    output ordered_filter_data_22__3 ;
    output ordered_filter_data_22__2 ;
    output ordered_filter_data_22__1 ;
    output ordered_filter_data_22__0 ;
    output ordered_filter_data_23__31 ;
    output ordered_filter_data_23__30 ;
    output ordered_filter_data_23__29 ;
    output ordered_filter_data_23__28 ;
    output ordered_filter_data_23__27 ;
    output ordered_filter_data_23__26 ;
    output ordered_filter_data_23__25 ;
    output ordered_filter_data_23__24 ;
    output ordered_filter_data_23__23 ;
    output ordered_filter_data_23__22 ;
    output ordered_filter_data_23__21 ;
    output ordered_filter_data_23__20 ;
    output ordered_filter_data_23__19 ;
    output ordered_filter_data_23__18 ;
    output ordered_filter_data_23__17 ;
    output ordered_filter_data_23__16 ;
    output ordered_filter_data_23__15 ;
    output ordered_filter_data_23__14 ;
    output ordered_filter_data_23__13 ;
    output ordered_filter_data_23__12 ;
    output ordered_filter_data_23__11 ;
    output ordered_filter_data_23__10 ;
    output ordered_filter_data_23__9 ;
    output ordered_filter_data_23__8 ;
    output ordered_filter_data_23__7 ;
    output ordered_filter_data_23__6 ;
    output ordered_filter_data_23__5 ;
    output ordered_filter_data_23__4 ;
    output ordered_filter_data_23__3 ;
    output ordered_filter_data_23__2 ;
    output ordered_filter_data_23__1 ;
    output ordered_filter_data_23__0 ;
    output ordered_filter_data_24__31 ;
    output ordered_filter_data_24__30 ;
    output ordered_filter_data_24__29 ;
    output ordered_filter_data_24__28 ;
    output ordered_filter_data_24__27 ;
    output ordered_filter_data_24__26 ;
    output ordered_filter_data_24__25 ;
    output ordered_filter_data_24__24 ;
    output ordered_filter_data_24__23 ;
    output ordered_filter_data_24__22 ;
    output ordered_filter_data_24__21 ;
    output ordered_filter_data_24__20 ;
    output ordered_filter_data_24__19 ;
    output ordered_filter_data_24__18 ;
    output ordered_filter_data_24__17 ;
    output ordered_filter_data_24__16 ;
    output ordered_filter_data_24__15 ;
    output ordered_filter_data_24__14 ;
    output ordered_filter_data_24__13 ;
    output ordered_filter_data_24__12 ;
    output ordered_filter_data_24__11 ;
    output ordered_filter_data_24__10 ;
    output ordered_filter_data_24__9 ;
    output ordered_filter_data_24__8 ;
    output ordered_filter_data_24__7 ;
    output ordered_filter_data_24__6 ;
    output ordered_filter_data_24__5 ;
    output ordered_filter_data_24__4 ;
    output ordered_filter_data_24__3 ;
    output ordered_filter_data_24__2 ;
    output ordered_filter_data_24__1 ;
    output ordered_filter_data_24__0 ;

    wire nx1206, nx1209, nx1211, nx1213, nx1215, nx1217, nx1219, nx1221, nx1223, 
         nx1225, nx1227, nx1229, nx1231, nx1233, nx1235, nx1237, nx1239, nx1241, 
         nx1243, nx1245, nx1247, nx1249, nx1251, nx1253, nx1255, nx1257, nx1259, 
         nx1261, nx1263, nx1265, nx1267, nx1269, nx1271, nx1273, nx1287, nx1301, 
         nx1315, nx1319, nx1321, nx1323, nx1317, nx1317_XX0_XREP32, nx1325, 
         nx1331, nx1345, nx1346, nx1354, nx1356, nx1358, nx1361, nx1363, nx1365, 
         nx1367, nx1369, nx1371, nx1373, nx1375, nx1377, nx1379, nx1381, nx1383, 
         nx1385, nx1387, nx1389, nx1391;



    assign ordered_img_data_0__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_0__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_1__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_2__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_3__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_4__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_5__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_6__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_7__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_8__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_9__30 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__29 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__28 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__27 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__26 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__25 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__24 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__23 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__22 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__21 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__20 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__19 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__18 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__17 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__16 = ordered_img_data_9__31 ;
    assign ordered_img_data_9__15 = ordered_img_data_9__31 ;
    assign ordered_img_data_10__30 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__29 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__28 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__27 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__26 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__25 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__24 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__23 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__22 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__21 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__20 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__19 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__18 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__17 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__16 = ordered_img_data_10__31 ;
    assign ordered_img_data_10__15 = ordered_img_data_10__31 ;
    assign ordered_img_data_11__30 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__29 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__28 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__27 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__26 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__25 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__24 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__23 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__22 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__21 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__20 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__19 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__18 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__17 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__16 = ordered_img_data_11__31 ;
    assign ordered_img_data_11__15 = ordered_img_data_11__31 ;
    assign ordered_img_data_12__30 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__29 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__28 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__27 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__26 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__25 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__24 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__23 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__22 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__21 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__20 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__19 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__18 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__17 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__16 = ordered_img_data_12__31 ;
    assign ordered_img_data_12__15 = ordered_img_data_12__31 ;
    assign ordered_img_data_13__30 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__29 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__28 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__27 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__26 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__25 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__24 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__23 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__22 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__21 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__20 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__19 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__18 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__17 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__16 = ordered_img_data_13__31 ;
    assign ordered_img_data_13__15 = ordered_img_data_13__31 ;
    assign ordered_img_data_14__30 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__29 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__28 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__27 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__26 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__25 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__24 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__23 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__22 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__21 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__20 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__19 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__18 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__17 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__16 = ordered_img_data_14__31 ;
    assign ordered_img_data_14__15 = ordered_img_data_14__31 ;
    assign ordered_img_data_15__30 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__29 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__28 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__27 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__26 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__25 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__24 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__23 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__22 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__21 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__20 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__19 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__18 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__17 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__16 = ordered_img_data_15__31 ;
    assign ordered_img_data_15__15 = ordered_img_data_15__31 ;
    assign ordered_img_data_16__30 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__29 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__28 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__27 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__26 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__25 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__24 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__23 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__22 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__21 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__20 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__19 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__18 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__17 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__16 = ordered_img_data_16__31 ;
    assign ordered_img_data_16__15 = ordered_img_data_16__31 ;
    assign ordered_img_data_17__30 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__29 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__28 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__27 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__26 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__25 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__24 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__23 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__22 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__21 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__20 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__19 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__18 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__17 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__16 = ordered_img_data_17__31 ;
    assign ordered_img_data_17__15 = ordered_img_data_17__31 ;
    assign ordered_img_data_18__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_18__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_19__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_20__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_21__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_22__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_23__0 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__31 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__30 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__29 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__28 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__27 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__26 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__25 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__24 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__23 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__22 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__21 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__20 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__19 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__18 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__17 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__16 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__15 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__14 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__13 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__12 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__11 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__10 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__9 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__8 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__7 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__6 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__5 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__4 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__3 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__2 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__1 = ordered_img_data_0__31 ;
    assign ordered_img_data_24__0 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__15 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__14 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__13 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__12 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__11 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__10 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__9 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__8 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__7 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__6 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__5 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__4 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__3 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__2 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__1 = ordered_img_data_0__31 ;
    assign ordered_filter_data_0__0 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__15 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__14 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__13 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__12 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__11 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__10 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__9 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__8 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__7 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__6 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__5 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__4 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__3 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__2 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__1 = ordered_img_data_0__31 ;
    assign ordered_filter_data_1__0 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__15 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__14 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__13 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__12 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__11 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__10 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__9 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__8 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__7 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__6 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__5 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__4 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__3 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__2 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__1 = ordered_img_data_0__31 ;
    assign ordered_filter_data_2__0 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_3__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_4__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_5__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_6__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_7__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_8__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_9__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_10__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_11__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_12__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_13__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_14__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_15__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_16__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_17__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__15 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__14 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__13 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__12 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__11 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__10 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__9 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__8 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__7 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__6 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__5 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__4 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__3 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__2 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__1 = ordered_img_data_0__31 ;
    assign ordered_filter_data_18__0 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__15 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__14 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__13 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__12 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__11 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__10 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__9 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__8 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__7 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__6 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__5 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__4 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__3 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__2 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__1 = ordered_img_data_0__31 ;
    assign ordered_filter_data_19__0 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__15 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__14 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__13 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__12 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__11 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__10 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__9 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__8 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__7 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__6 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__5 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__4 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__3 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__2 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__1 = ordered_img_data_0__31 ;
    assign ordered_filter_data_20__0 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__15 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__14 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__13 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__12 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__11 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__10 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__9 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__8 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__7 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__6 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__5 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__4 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__3 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__2 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__1 = ordered_img_data_0__31 ;
    assign ordered_filter_data_21__0 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__15 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__14 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__13 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__12 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__11 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__10 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__9 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__8 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__7 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__6 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__5 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__4 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__3 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__2 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__1 = ordered_img_data_0__31 ;
    assign ordered_filter_data_22__0 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__15 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__14 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__13 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__12 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__11 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__10 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__9 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__8 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__7 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__6 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__5 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__4 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__3 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__2 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__1 = ordered_img_data_0__31 ;
    assign ordered_filter_data_23__0 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__31 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__30 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__29 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__28 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__27 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__26 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__25 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__24 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__23 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__22 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__21 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__20 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__19 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__18 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__17 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__16 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__15 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__14 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__13 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__12 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__11 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__10 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__9 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__8 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__7 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__6 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__5 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__4 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__3 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__2 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__1 = ordered_img_data_0__31 ;
    assign ordered_filter_data_24__0 = ordered_img_data_0__31 ;
    fake_gnd ix46 (.Y (ordered_img_data_0__31)) ;
    mux21_ni ix7 (.Y (ordered_filter_data_17__0), .A0 (filter_data_17__0), .A1 (
             filter_data_8__0), .S0 (nx1206)) ;
    mux21_ni ix15 (.Y (ordered_filter_data_17__1), .A0 (filter_data_17__1), .A1 (
             filter_data_8__1), .S0 (nx1206)) ;
    mux21_ni ix23 (.Y (ordered_filter_data_17__2), .A0 (filter_data_17__2), .A1 (
             filter_data_8__2), .S0 (nx1206)) ;
    mux21_ni ix31 (.Y (ordered_filter_data_17__3), .A0 (filter_data_17__3), .A1 (
             filter_data_8__3), .S0 (nx1206)) ;
    mux21_ni ix39 (.Y (ordered_filter_data_17__4), .A0 (filter_data_17__4), .A1 (
             filter_data_8__4), .S0 (nx1206)) ;
    mux21_ni ix47 (.Y (ordered_filter_data_17__5), .A0 (filter_data_17__5), .A1 (
             filter_data_8__5), .S0 (nx1206)) ;
    mux21_ni ix55 (.Y (ordered_filter_data_17__6), .A0 (filter_data_17__6), .A1 (
             filter_data_8__6), .S0 (nx1206)) ;
    mux21_ni ix63 (.Y (ordered_filter_data_17__7), .A0 (filter_data_17__7), .A1 (
             filter_data_8__7), .S0 (nx1209)) ;
    mux21_ni ix71 (.Y (ordered_filter_data_17__8), .A0 (filter_data_17__8), .A1 (
             filter_data_8__8), .S0 (nx1209)) ;
    mux21_ni ix79 (.Y (ordered_filter_data_17__9), .A0 (filter_data_17__9), .A1 (
             filter_data_8__9), .S0 (nx1209)) ;
    mux21_ni ix87 (.Y (ordered_filter_data_17__10), .A0 (filter_data_17__10), .A1 (
             filter_data_8__10), .S0 (nx1209)) ;
    mux21_ni ix95 (.Y (ordered_filter_data_17__11), .A0 (filter_data_17__11), .A1 (
             filter_data_8__11), .S0 (nx1209)) ;
    mux21_ni ix103 (.Y (ordered_filter_data_17__12), .A0 (filter_data_17__12), .A1 (
             filter_data_8__12), .S0 (nx1209)) ;
    mux21_ni ix111 (.Y (ordered_filter_data_17__13), .A0 (filter_data_17__13), .A1 (
             filter_data_8__13), .S0 (nx1209)) ;
    mux21_ni ix119 (.Y (ordered_filter_data_17__14), .A0 (filter_data_17__14), .A1 (
             filter_data_8__14), .S0 (nx1211)) ;
    mux21_ni ix127 (.Y (ordered_filter_data_17__15), .A0 (filter_data_17__31), .A1 (
             filter_data_8__31), .S0 (nx1211)) ;
    mux21_ni ix391 (.Y (ordered_filter_data_16__0), .A0 (filter_data_16__0), .A1 (
             filter_data_7__0), .S0 (nx1211)) ;
    mux21_ni ix399 (.Y (ordered_filter_data_16__1), .A0 (filter_data_16__1), .A1 (
             filter_data_7__1), .S0 (nx1211)) ;
    mux21_ni ix407 (.Y (ordered_filter_data_16__2), .A0 (filter_data_16__2), .A1 (
             filter_data_7__2), .S0 (nx1211)) ;
    mux21_ni ix415 (.Y (ordered_filter_data_16__3), .A0 (filter_data_16__3), .A1 (
             filter_data_7__3), .S0 (nx1211)) ;
    mux21_ni ix423 (.Y (ordered_filter_data_16__4), .A0 (filter_data_16__4), .A1 (
             filter_data_7__4), .S0 (nx1211)) ;
    mux21_ni ix431 (.Y (ordered_filter_data_16__5), .A0 (filter_data_16__5), .A1 (
             filter_data_7__5), .S0 (nx1213)) ;
    mux21_ni ix439 (.Y (ordered_filter_data_16__6), .A0 (filter_data_16__6), .A1 (
             filter_data_7__6), .S0 (nx1213)) ;
    mux21_ni ix447 (.Y (ordered_filter_data_16__7), .A0 (filter_data_16__7), .A1 (
             filter_data_7__7), .S0 (nx1213)) ;
    mux21_ni ix455 (.Y (ordered_filter_data_16__8), .A0 (filter_data_16__8), .A1 (
             filter_data_7__8), .S0 (nx1213)) ;
    mux21_ni ix463 (.Y (ordered_filter_data_16__9), .A0 (filter_data_16__9), .A1 (
             filter_data_7__9), .S0 (nx1213)) ;
    mux21_ni ix471 (.Y (ordered_filter_data_16__10), .A0 (filter_data_16__10), .A1 (
             filter_data_7__10), .S0 (nx1213)) ;
    mux21_ni ix479 (.Y (ordered_filter_data_16__11), .A0 (filter_data_16__11), .A1 (
             filter_data_7__11), .S0 (nx1213)) ;
    mux21_ni ix487 (.Y (ordered_filter_data_16__12), .A0 (filter_data_16__12), .A1 (
             filter_data_7__12), .S0 (nx1215)) ;
    mux21_ni ix495 (.Y (ordered_filter_data_16__13), .A0 (filter_data_16__13), .A1 (
             filter_data_7__13), .S0 (nx1215)) ;
    mux21_ni ix503 (.Y (ordered_filter_data_16__14), .A0 (filter_data_16__14), .A1 (
             filter_data_7__14), .S0 (nx1215)) ;
    mux21_ni ix511 (.Y (ordered_filter_data_16__15), .A0 (filter_data_16__31), .A1 (
             filter_data_7__31), .S0 (nx1215)) ;
    mux21_ni ix775 (.Y (ordered_filter_data_15__0), .A0 (filter_data_15__0), .A1 (
             filter_data_6__0), .S0 (nx1215)) ;
    mux21_ni ix783 (.Y (ordered_filter_data_15__1), .A0 (filter_data_15__1), .A1 (
             filter_data_6__1), .S0 (nx1215)) ;
    mux21_ni ix791 (.Y (ordered_filter_data_15__2), .A0 (filter_data_15__2), .A1 (
             filter_data_6__2), .S0 (nx1215)) ;
    mux21_ni ix799 (.Y (ordered_filter_data_15__3), .A0 (filter_data_15__3), .A1 (
             filter_data_6__3), .S0 (nx1217)) ;
    mux21_ni ix807 (.Y (ordered_filter_data_15__4), .A0 (filter_data_15__4), .A1 (
             filter_data_6__4), .S0 (nx1217)) ;
    mux21_ni ix815 (.Y (ordered_filter_data_15__5), .A0 (filter_data_15__5), .A1 (
             filter_data_6__5), .S0 (nx1217)) ;
    mux21_ni ix823 (.Y (ordered_filter_data_15__6), .A0 (filter_data_15__6), .A1 (
             filter_data_6__6), .S0 (nx1217)) ;
    mux21_ni ix831 (.Y (ordered_filter_data_15__7), .A0 (filter_data_15__7), .A1 (
             filter_data_6__7), .S0 (nx1217)) ;
    mux21_ni ix839 (.Y (ordered_filter_data_15__8), .A0 (filter_data_15__8), .A1 (
             filter_data_6__8), .S0 (nx1217)) ;
    mux21_ni ix847 (.Y (ordered_filter_data_15__9), .A0 (filter_data_15__9), .A1 (
             filter_data_6__9), .S0 (nx1217)) ;
    mux21_ni ix855 (.Y (ordered_filter_data_15__10), .A0 (filter_data_15__10), .A1 (
             filter_data_6__10), .S0 (nx1219)) ;
    mux21_ni ix863 (.Y (ordered_filter_data_15__11), .A0 (filter_data_15__11), .A1 (
             filter_data_6__11), .S0 (nx1219)) ;
    mux21_ni ix871 (.Y (ordered_filter_data_15__12), .A0 (filter_data_15__12), .A1 (
             filter_data_6__12), .S0 (nx1219)) ;
    mux21_ni ix879 (.Y (ordered_filter_data_15__13), .A0 (filter_data_15__13), .A1 (
             filter_data_6__13), .S0 (nx1219)) ;
    mux21_ni ix887 (.Y (ordered_filter_data_15__14), .A0 (filter_data_15__14), .A1 (
             filter_data_6__14), .S0 (nx1219)) ;
    mux21_ni ix895 (.Y (ordered_filter_data_15__15), .A0 (filter_data_15__31), .A1 (
             filter_data_6__31), .S0 (nx1219)) ;
    mux21_ni ix1159 (.Y (ordered_filter_data_14__0), .A0 (filter_data_14__0), .A1 (
             filter_data_5__0), .S0 (nx1219)) ;
    mux21_ni ix1167 (.Y (ordered_filter_data_14__1), .A0 (filter_data_14__1), .A1 (
             filter_data_5__1), .S0 (nx1221)) ;
    mux21_ni ix1175 (.Y (ordered_filter_data_14__2), .A0 (filter_data_14__2), .A1 (
             filter_data_5__2), .S0 (nx1221)) ;
    mux21_ni ix1183 (.Y (ordered_filter_data_14__3), .A0 (filter_data_14__3), .A1 (
             filter_data_5__3), .S0 (nx1221)) ;
    mux21_ni ix1191 (.Y (ordered_filter_data_14__4), .A0 (filter_data_14__4), .A1 (
             filter_data_5__4), .S0 (nx1221)) ;
    mux21_ni ix1199 (.Y (ordered_filter_data_14__5), .A0 (filter_data_14__5), .A1 (
             filter_data_5__5), .S0 (nx1221)) ;
    mux21_ni ix1207 (.Y (ordered_filter_data_14__6), .A0 (filter_data_14__6), .A1 (
             filter_data_5__6), .S0 (nx1221)) ;
    mux21_ni ix1215 (.Y (ordered_filter_data_14__7), .A0 (filter_data_14__7), .A1 (
             filter_data_5__7), .S0 (nx1221)) ;
    mux21_ni ix1223 (.Y (ordered_filter_data_14__8), .A0 (filter_data_14__8), .A1 (
             filter_data_5__8), .S0 (nx1223)) ;
    mux21_ni ix1231 (.Y (ordered_filter_data_14__9), .A0 (filter_data_14__9), .A1 (
             filter_data_5__9), .S0 (nx1223)) ;
    mux21_ni ix1239 (.Y (ordered_filter_data_14__10), .A0 (filter_data_14__10), 
             .A1 (filter_data_5__10), .S0 (nx1223)) ;
    mux21_ni ix1247 (.Y (ordered_filter_data_14__11), .A0 (filter_data_14__11), 
             .A1 (filter_data_5__11), .S0 (nx1223)) ;
    mux21_ni ix1255 (.Y (ordered_filter_data_14__12), .A0 (filter_data_14__12), 
             .A1 (filter_data_5__12), .S0 (nx1223)) ;
    mux21_ni ix1263 (.Y (ordered_filter_data_14__13), .A0 (filter_data_14__13), 
             .A1 (filter_data_5__13), .S0 (nx1223)) ;
    mux21_ni ix1271 (.Y (ordered_filter_data_14__14), .A0 (filter_data_14__14), 
             .A1 (filter_data_5__14), .S0 (nx1223)) ;
    mux21_ni ix1279 (.Y (ordered_filter_data_14__15), .A0 (filter_data_14__31), 
             .A1 (filter_data_5__31), .S0 (nx1225)) ;
    mux21_ni ix1543 (.Y (ordered_filter_data_13__0), .A0 (filter_data_9__0), .A1 (
             filter_data_4__0), .S0 (nx1225)) ;
    mux21_ni ix1551 (.Y (ordered_filter_data_13__1), .A0 (filter_data_9__1), .A1 (
             filter_data_4__1), .S0 (nx1225)) ;
    mux21_ni ix1559 (.Y (ordered_filter_data_13__2), .A0 (filter_data_9__2), .A1 (
             filter_data_4__2), .S0 (nx1225)) ;
    mux21_ni ix1567 (.Y (ordered_filter_data_13__3), .A0 (filter_data_9__3), .A1 (
             filter_data_4__3), .S0 (nx1225)) ;
    mux21_ni ix1575 (.Y (ordered_filter_data_13__4), .A0 (filter_data_9__4), .A1 (
             filter_data_4__4), .S0 (nx1225)) ;
    mux21_ni ix1583 (.Y (ordered_filter_data_13__5), .A0 (filter_data_9__5), .A1 (
             filter_data_4__5), .S0 (nx1225)) ;
    mux21_ni ix1591 (.Y (ordered_filter_data_13__6), .A0 (filter_data_9__6), .A1 (
             filter_data_4__6), .S0 (nx1227)) ;
    mux21_ni ix1599 (.Y (ordered_filter_data_13__7), .A0 (filter_data_9__7), .A1 (
             filter_data_4__7), .S0 (nx1227)) ;
    mux21_ni ix1607 (.Y (ordered_filter_data_13__8), .A0 (filter_data_9__8), .A1 (
             filter_data_4__8), .S0 (nx1227)) ;
    mux21_ni ix1615 (.Y (ordered_filter_data_13__9), .A0 (filter_data_9__9), .A1 (
             filter_data_4__9), .S0 (nx1227)) ;
    mux21_ni ix1623 (.Y (ordered_filter_data_13__10), .A0 (filter_data_9__10), .A1 (
             filter_data_4__10), .S0 (nx1227)) ;
    mux21_ni ix1631 (.Y (ordered_filter_data_13__11), .A0 (filter_data_9__11), .A1 (
             filter_data_4__11), .S0 (nx1227)) ;
    mux21_ni ix1639 (.Y (ordered_filter_data_13__12), .A0 (filter_data_9__12), .A1 (
             filter_data_4__12), .S0 (nx1227)) ;
    mux21_ni ix1647 (.Y (ordered_filter_data_13__13), .A0 (filter_data_9__13), .A1 (
             filter_data_4__13), .S0 (nx1229)) ;
    mux21_ni ix1655 (.Y (ordered_filter_data_13__14), .A0 (filter_data_9__14), .A1 (
             filter_data_4__14), .S0 (nx1229)) ;
    mux21_ni ix1663 (.Y (ordered_filter_data_13__15), .A0 (filter_data_9__31), .A1 (
             filter_data_4__31), .S0 (nx1229)) ;
    mux21_ni ix1927 (.Y (ordered_filter_data_12__0), .A0 (filter_data_4__0), .A1 (
             filter_data_3__0), .S0 (nx1229)) ;
    mux21_ni ix1935 (.Y (ordered_filter_data_12__1), .A0 (filter_data_4__1), .A1 (
             filter_data_3__1), .S0 (nx1229)) ;
    mux21_ni ix1943 (.Y (ordered_filter_data_12__2), .A0 (filter_data_4__2), .A1 (
             filter_data_3__2), .S0 (nx1229)) ;
    mux21_ni ix1951 (.Y (ordered_filter_data_12__3), .A0 (filter_data_4__3), .A1 (
             filter_data_3__3), .S0 (nx1229)) ;
    mux21_ni ix1959 (.Y (ordered_filter_data_12__4), .A0 (filter_data_4__4), .A1 (
             filter_data_3__4), .S0 (nx1231)) ;
    mux21_ni ix1967 (.Y (ordered_filter_data_12__5), .A0 (filter_data_4__5), .A1 (
             filter_data_3__5), .S0 (nx1231)) ;
    mux21_ni ix1975 (.Y (ordered_filter_data_12__6), .A0 (filter_data_4__6), .A1 (
             filter_data_3__6), .S0 (nx1231)) ;
    mux21_ni ix1983 (.Y (ordered_filter_data_12__7), .A0 (filter_data_4__7), .A1 (
             filter_data_3__7), .S0 (nx1231)) ;
    mux21_ni ix1991 (.Y (ordered_filter_data_12__8), .A0 (filter_data_4__8), .A1 (
             filter_data_3__8), .S0 (nx1231)) ;
    mux21_ni ix1999 (.Y (ordered_filter_data_12__9), .A0 (filter_data_4__9), .A1 (
             filter_data_3__9), .S0 (nx1231)) ;
    mux21_ni ix2007 (.Y (ordered_filter_data_12__10), .A0 (filter_data_4__10), .A1 (
             filter_data_3__10), .S0 (nx1231)) ;
    mux21_ni ix2015 (.Y (ordered_filter_data_12__11), .A0 (filter_data_4__11), .A1 (
             filter_data_3__11), .S0 (nx1233)) ;
    mux21_ni ix2023 (.Y (ordered_filter_data_12__12), .A0 (filter_data_4__12), .A1 (
             filter_data_3__12), .S0 (nx1233)) ;
    mux21_ni ix2031 (.Y (ordered_filter_data_12__13), .A0 (filter_data_4__13), .A1 (
             filter_data_3__13), .S0 (nx1233)) ;
    mux21_ni ix2039 (.Y (ordered_filter_data_12__14), .A0 (filter_data_4__14), .A1 (
             filter_data_3__14), .S0 (nx1233)) ;
    mux21_ni ix2047 (.Y (ordered_filter_data_12__15), .A0 (filter_data_4__31), .A1 (
             filter_data_3__31), .S0 (nx1233)) ;
    mux21_ni ix2311 (.Y (ordered_filter_data_11__0), .A0 (filter_data_13__0), .A1 (
             filter_data_2__0), .S0 (nx1233)) ;
    mux21_ni ix2319 (.Y (ordered_filter_data_11__1), .A0 (filter_data_13__1), .A1 (
             filter_data_2__1), .S0 (nx1233)) ;
    mux21_ni ix2327 (.Y (ordered_filter_data_11__2), .A0 (filter_data_13__2), .A1 (
             filter_data_2__2), .S0 (nx1235)) ;
    mux21_ni ix2335 (.Y (ordered_filter_data_11__3), .A0 (filter_data_13__3), .A1 (
             filter_data_2__3), .S0 (nx1235)) ;
    mux21_ni ix2343 (.Y (ordered_filter_data_11__4), .A0 (filter_data_13__4), .A1 (
             filter_data_2__4), .S0 (nx1235)) ;
    mux21_ni ix2351 (.Y (ordered_filter_data_11__5), .A0 (filter_data_13__5), .A1 (
             filter_data_2__5), .S0 (nx1235)) ;
    mux21_ni ix2359 (.Y (ordered_filter_data_11__6), .A0 (filter_data_13__6), .A1 (
             filter_data_2__6), .S0 (nx1235)) ;
    mux21_ni ix2367 (.Y (ordered_filter_data_11__7), .A0 (filter_data_13__7), .A1 (
             filter_data_2__7), .S0 (nx1235)) ;
    mux21_ni ix2375 (.Y (ordered_filter_data_11__8), .A0 (filter_data_13__8), .A1 (
             filter_data_2__8), .S0 (nx1235)) ;
    mux21_ni ix2383 (.Y (ordered_filter_data_11__9), .A0 (filter_data_13__9), .A1 (
             filter_data_2__9), .S0 (nx1237)) ;
    mux21_ni ix2391 (.Y (ordered_filter_data_11__10), .A0 (filter_data_13__10), 
             .A1 (filter_data_2__10), .S0 (nx1237)) ;
    mux21_ni ix2399 (.Y (ordered_filter_data_11__11), .A0 (filter_data_13__11), 
             .A1 (filter_data_2__11), .S0 (nx1237)) ;
    mux21_ni ix2407 (.Y (ordered_filter_data_11__12), .A0 (filter_data_13__12), 
             .A1 (filter_data_2__12), .S0 (nx1237)) ;
    mux21_ni ix2415 (.Y (ordered_filter_data_11__13), .A0 (filter_data_13__13), 
             .A1 (filter_data_2__13), .S0 (nx1237)) ;
    mux21_ni ix2423 (.Y (ordered_filter_data_11__14), .A0 (filter_data_13__14), 
             .A1 (filter_data_2__14), .S0 (nx1237)) ;
    mux21_ni ix2431 (.Y (ordered_filter_data_11__15), .A0 (filter_data_13__31), 
             .A1 (filter_data_2__31), .S0 (nx1237)) ;
    mux21_ni ix2567 (.Y (ordered_filter_data_10__0), .A0 (filter_data_8__0), .A1 (
             filter_data_1__0), .S0 (nx1239)) ;
    mux21_ni ix2575 (.Y (ordered_filter_data_10__1), .A0 (filter_data_8__1), .A1 (
             filter_data_1__1), .S0 (nx1239)) ;
    mux21_ni ix2583 (.Y (ordered_filter_data_10__2), .A0 (filter_data_8__2), .A1 (
             filter_data_1__2), .S0 (nx1239)) ;
    mux21_ni ix2591 (.Y (ordered_filter_data_10__3), .A0 (filter_data_8__3), .A1 (
             filter_data_1__3), .S0 (nx1239)) ;
    mux21_ni ix2599 (.Y (ordered_filter_data_10__4), .A0 (filter_data_8__4), .A1 (
             filter_data_1__4), .S0 (nx1239)) ;
    mux21_ni ix2607 (.Y (ordered_filter_data_10__5), .A0 (filter_data_8__5), .A1 (
             filter_data_1__5), .S0 (nx1239)) ;
    mux21_ni ix2615 (.Y (ordered_filter_data_10__6), .A0 (filter_data_8__6), .A1 (
             filter_data_1__6), .S0 (nx1239)) ;
    mux21_ni ix2623 (.Y (ordered_filter_data_10__7), .A0 (filter_data_8__7), .A1 (
             filter_data_1__7), .S0 (nx1241)) ;
    mux21_ni ix2631 (.Y (ordered_filter_data_10__8), .A0 (filter_data_8__8), .A1 (
             filter_data_1__8), .S0 (nx1241)) ;
    mux21_ni ix2639 (.Y (ordered_filter_data_10__9), .A0 (filter_data_8__9), .A1 (
             filter_data_1__9), .S0 (nx1241)) ;
    mux21_ni ix2647 (.Y (ordered_filter_data_10__10), .A0 (filter_data_8__10), .A1 (
             filter_data_1__10), .S0 (nx1241)) ;
    mux21_ni ix2655 (.Y (ordered_filter_data_10__11), .A0 (filter_data_8__11), .A1 (
             filter_data_1__11), .S0 (nx1241)) ;
    mux21_ni ix2663 (.Y (ordered_filter_data_10__12), .A0 (filter_data_8__12), .A1 (
             filter_data_1__12), .S0 (nx1241)) ;
    mux21_ni ix2671 (.Y (ordered_filter_data_10__13), .A0 (filter_data_8__13), .A1 (
             filter_data_1__13), .S0 (nx1241)) ;
    mux21_ni ix2679 (.Y (ordered_filter_data_10__14), .A0 (filter_data_8__14), .A1 (
             filter_data_1__14), .S0 (nx1243)) ;
    mux21_ni ix2687 (.Y (ordered_filter_data_10__15), .A0 (filter_data_8__31), .A1 (
             filter_data_1__31), .S0 (nx1243)) ;
    mux21_ni ix2823 (.Y (ordered_filter_data_9__0), .A0 (filter_data_3__0), .A1 (
             filter_data_0__0), .S0 (nx1243)) ;
    mux21_ni ix2831 (.Y (ordered_filter_data_9__1), .A0 (filter_data_3__1), .A1 (
             filter_data_0__1), .S0 (nx1243)) ;
    mux21_ni ix2839 (.Y (ordered_filter_data_9__2), .A0 (filter_data_3__2), .A1 (
             filter_data_0__2), .S0 (nx1243)) ;
    mux21_ni ix2847 (.Y (ordered_filter_data_9__3), .A0 (filter_data_3__3), .A1 (
             filter_data_0__3), .S0 (nx1243)) ;
    mux21_ni ix2855 (.Y (ordered_filter_data_9__4), .A0 (filter_data_3__4), .A1 (
             filter_data_0__4), .S0 (nx1243)) ;
    mux21_ni ix2863 (.Y (ordered_filter_data_9__5), .A0 (filter_data_3__5), .A1 (
             filter_data_0__5), .S0 (nx1245)) ;
    mux21_ni ix2871 (.Y (ordered_filter_data_9__6), .A0 (filter_data_3__6), .A1 (
             filter_data_0__6), .S0 (nx1245)) ;
    mux21_ni ix2879 (.Y (ordered_filter_data_9__7), .A0 (filter_data_3__7), .A1 (
             filter_data_0__7), .S0 (nx1245)) ;
    mux21_ni ix2887 (.Y (ordered_filter_data_9__8), .A0 (filter_data_3__8), .A1 (
             filter_data_0__8), .S0 (nx1245)) ;
    mux21_ni ix2895 (.Y (ordered_filter_data_9__9), .A0 (filter_data_3__9), .A1 (
             filter_data_0__9), .S0 (nx1245)) ;
    mux21_ni ix2903 (.Y (ordered_filter_data_9__10), .A0 (filter_data_3__10), .A1 (
             filter_data_0__10), .S0 (nx1245)) ;
    mux21_ni ix2911 (.Y (ordered_filter_data_9__11), .A0 (filter_data_3__11), .A1 (
             filter_data_0__11), .S0 (nx1245)) ;
    mux21_ni ix2919 (.Y (ordered_filter_data_9__12), .A0 (filter_data_3__12), .A1 (
             filter_data_0__12), .S0 (nx1247)) ;
    mux21_ni ix2927 (.Y (ordered_filter_data_9__13), .A0 (filter_data_3__13), .A1 (
             filter_data_0__13), .S0 (nx1247)) ;
    mux21_ni ix2935 (.Y (ordered_filter_data_9__14), .A0 (filter_data_3__14), .A1 (
             filter_data_0__14), .S0 (nx1247)) ;
    mux21_ni ix2943 (.Y (ordered_filter_data_9__15), .A0 (filter_data_3__31), .A1 (
             filter_data_0__31), .S0 (nx1247)) ;
    mux21_ni ix263 (.Y (ordered_filter_data_8__0), .A0 (filter_data_12__0), .A1 (
             filter_data_8__0), .S0 (nx1247)) ;
    mux21_ni ix271 (.Y (ordered_filter_data_8__1), .A0 (filter_data_12__1), .A1 (
             filter_data_8__1), .S0 (nx1247)) ;
    mux21_ni ix279 (.Y (ordered_filter_data_8__2), .A0 (filter_data_12__2), .A1 (
             filter_data_8__2), .S0 (nx1247)) ;
    mux21_ni ix287 (.Y (ordered_filter_data_8__3), .A0 (filter_data_12__3), .A1 (
             filter_data_8__3), .S0 (nx1249)) ;
    mux21_ni ix295 (.Y (ordered_filter_data_8__4), .A0 (filter_data_12__4), .A1 (
             filter_data_8__4), .S0 (nx1249)) ;
    mux21_ni ix303 (.Y (ordered_filter_data_8__5), .A0 (filter_data_12__5), .A1 (
             filter_data_8__5), .S0 (nx1249)) ;
    mux21_ni ix311 (.Y (ordered_filter_data_8__6), .A0 (filter_data_12__6), .A1 (
             filter_data_8__6), .S0 (nx1249)) ;
    mux21_ni ix319 (.Y (ordered_filter_data_8__7), .A0 (filter_data_12__7), .A1 (
             filter_data_8__7), .S0 (nx1249)) ;
    mux21_ni ix327 (.Y (ordered_filter_data_8__8), .A0 (filter_data_12__8), .A1 (
             filter_data_8__8), .S0 (nx1249)) ;
    mux21_ni ix335 (.Y (ordered_filter_data_8__9), .A0 (filter_data_12__9), .A1 (
             filter_data_8__9), .S0 (nx1249)) ;
    mux21_ni ix343 (.Y (ordered_filter_data_8__10), .A0 (filter_data_12__10), .A1 (
             filter_data_8__10), .S0 (nx1251)) ;
    mux21_ni ix351 (.Y (ordered_filter_data_8__11), .A0 (filter_data_12__11), .A1 (
             filter_data_8__11), .S0 (nx1251)) ;
    mux21_ni ix359 (.Y (ordered_filter_data_8__12), .A0 (filter_data_12__12), .A1 (
             filter_data_8__12), .S0 (nx1251)) ;
    mux21_ni ix367 (.Y (ordered_filter_data_8__13), .A0 (filter_data_12__13), .A1 (
             filter_data_8__13), .S0 (nx1251)) ;
    mux21_ni ix375 (.Y (ordered_filter_data_8__14), .A0 (filter_data_12__14), .A1 (
             filter_data_8__14), .S0 (nx1251)) ;
    mux21_ni ix383 (.Y (ordered_filter_data_8__15), .A0 (filter_data_12__31), .A1 (
             filter_data_8__31), .S0 (nx1251)) ;
    mux21_ni ix647 (.Y (ordered_filter_data_7__0), .A0 (filter_data_11__0), .A1 (
             filter_data_7__0), .S0 (nx1251)) ;
    mux21_ni ix655 (.Y (ordered_filter_data_7__1), .A0 (filter_data_11__1), .A1 (
             filter_data_7__1), .S0 (nx1253)) ;
    mux21_ni ix663 (.Y (ordered_filter_data_7__2), .A0 (filter_data_11__2), .A1 (
             filter_data_7__2), .S0 (nx1253)) ;
    mux21_ni ix671 (.Y (ordered_filter_data_7__3), .A0 (filter_data_11__3), .A1 (
             filter_data_7__3), .S0 (nx1253)) ;
    mux21_ni ix679 (.Y (ordered_filter_data_7__4), .A0 (filter_data_11__4), .A1 (
             filter_data_7__4), .S0 (nx1253)) ;
    mux21_ni ix687 (.Y (ordered_filter_data_7__5), .A0 (filter_data_11__5), .A1 (
             filter_data_7__5), .S0 (nx1253)) ;
    mux21_ni ix695 (.Y (ordered_filter_data_7__6), .A0 (filter_data_11__6), .A1 (
             filter_data_7__6), .S0 (nx1253)) ;
    mux21_ni ix703 (.Y (ordered_filter_data_7__7), .A0 (filter_data_11__7), .A1 (
             filter_data_7__7), .S0 (nx1253)) ;
    mux21_ni ix711 (.Y (ordered_filter_data_7__8), .A0 (filter_data_11__8), .A1 (
             filter_data_7__8), .S0 (nx1255)) ;
    mux21_ni ix719 (.Y (ordered_filter_data_7__9), .A0 (filter_data_11__9), .A1 (
             filter_data_7__9), .S0 (nx1255)) ;
    mux21_ni ix727 (.Y (ordered_filter_data_7__10), .A0 (filter_data_11__10), .A1 (
             filter_data_7__10), .S0 (nx1255)) ;
    mux21_ni ix735 (.Y (ordered_filter_data_7__11), .A0 (filter_data_11__11), .A1 (
             filter_data_7__11), .S0 (nx1255)) ;
    mux21_ni ix743 (.Y (ordered_filter_data_7__12), .A0 (filter_data_11__12), .A1 (
             filter_data_7__12), .S0 (nx1255)) ;
    mux21_ni ix751 (.Y (ordered_filter_data_7__13), .A0 (filter_data_11__13), .A1 (
             filter_data_7__13), .S0 (nx1255)) ;
    mux21_ni ix759 (.Y (ordered_filter_data_7__14), .A0 (filter_data_11__14), .A1 (
             filter_data_7__14), .S0 (nx1255)) ;
    mux21_ni ix767 (.Y (ordered_filter_data_7__15), .A0 (filter_data_11__31), .A1 (
             filter_data_7__31), .S0 (nx1257)) ;
    mux21_ni ix1031 (.Y (ordered_filter_data_6__0), .A0 (filter_data_10__0), .A1 (
             filter_data_6__0), .S0 (nx1257)) ;
    mux21_ni ix1039 (.Y (ordered_filter_data_6__1), .A0 (filter_data_10__1), .A1 (
             filter_data_6__1), .S0 (nx1257)) ;
    mux21_ni ix1047 (.Y (ordered_filter_data_6__2), .A0 (filter_data_10__2), .A1 (
             filter_data_6__2), .S0 (nx1257)) ;
    mux21_ni ix1055 (.Y (ordered_filter_data_6__3), .A0 (filter_data_10__3), .A1 (
             filter_data_6__3), .S0 (nx1257)) ;
    mux21_ni ix1063 (.Y (ordered_filter_data_6__4), .A0 (filter_data_10__4), .A1 (
             filter_data_6__4), .S0 (nx1257)) ;
    mux21_ni ix1071 (.Y (ordered_filter_data_6__5), .A0 (filter_data_10__5), .A1 (
             filter_data_6__5), .S0 (nx1257)) ;
    mux21_ni ix1079 (.Y (ordered_filter_data_6__6), .A0 (filter_data_10__6), .A1 (
             filter_data_6__6), .S0 (nx1259)) ;
    mux21_ni ix1087 (.Y (ordered_filter_data_6__7), .A0 (filter_data_10__7), .A1 (
             filter_data_6__7), .S0 (nx1259)) ;
    mux21_ni ix1095 (.Y (ordered_filter_data_6__8), .A0 (filter_data_10__8), .A1 (
             filter_data_6__8), .S0 (nx1259)) ;
    mux21_ni ix1103 (.Y (ordered_filter_data_6__9), .A0 (filter_data_10__9), .A1 (
             filter_data_6__9), .S0 (nx1259)) ;
    mux21_ni ix1111 (.Y (ordered_filter_data_6__10), .A0 (filter_data_10__10), .A1 (
             filter_data_6__10), .S0 (nx1259)) ;
    mux21_ni ix1119 (.Y (ordered_filter_data_6__11), .A0 (filter_data_10__11), .A1 (
             filter_data_6__11), .S0 (nx1259)) ;
    mux21_ni ix1127 (.Y (ordered_filter_data_6__12), .A0 (filter_data_10__12), .A1 (
             filter_data_6__12), .S0 (nx1259)) ;
    mux21_ni ix1135 (.Y (ordered_filter_data_6__13), .A0 (filter_data_10__13), .A1 (
             filter_data_6__13), .S0 (nx1261)) ;
    mux21_ni ix1143 (.Y (ordered_filter_data_6__14), .A0 (filter_data_10__14), .A1 (
             filter_data_6__14), .S0 (nx1261)) ;
    mux21_ni ix1151 (.Y (ordered_filter_data_6__15), .A0 (filter_data_10__31), .A1 (
             filter_data_6__31), .S0 (nx1261)) ;
    mux21_ni ix1415 (.Y (ordered_filter_data_5__0), .A0 (filter_data_7__0), .A1 (
             filter_data_5__0), .S0 (nx1261)) ;
    mux21_ni ix1423 (.Y (ordered_filter_data_5__1), .A0 (filter_data_7__1), .A1 (
             filter_data_5__1), .S0 (nx1261)) ;
    mux21_ni ix1431 (.Y (ordered_filter_data_5__2), .A0 (filter_data_7__2), .A1 (
             filter_data_5__2), .S0 (nx1261)) ;
    mux21_ni ix1439 (.Y (ordered_filter_data_5__3), .A0 (filter_data_7__3), .A1 (
             filter_data_5__3), .S0 (nx1261)) ;
    mux21_ni ix1447 (.Y (ordered_filter_data_5__4), .A0 (filter_data_7__4), .A1 (
             filter_data_5__4), .S0 (nx1263)) ;
    mux21_ni ix1455 (.Y (ordered_filter_data_5__5), .A0 (filter_data_7__5), .A1 (
             filter_data_5__5), .S0 (nx1263)) ;
    mux21_ni ix1463 (.Y (ordered_filter_data_5__6), .A0 (filter_data_7__6), .A1 (
             filter_data_5__6), .S0 (nx1263)) ;
    mux21_ni ix1471 (.Y (ordered_filter_data_5__7), .A0 (filter_data_7__7), .A1 (
             filter_data_5__7), .S0 (nx1263)) ;
    mux21_ni ix1479 (.Y (ordered_filter_data_5__8), .A0 (filter_data_7__8), .A1 (
             filter_data_5__8), .S0 (nx1263)) ;
    mux21_ni ix1487 (.Y (ordered_filter_data_5__9), .A0 (filter_data_7__9), .A1 (
             filter_data_5__9), .S0 (nx1263)) ;
    mux21_ni ix1495 (.Y (ordered_filter_data_5__10), .A0 (filter_data_7__10), .A1 (
             filter_data_5__10), .S0 (nx1263)) ;
    mux21_ni ix1503 (.Y (ordered_filter_data_5__11), .A0 (filter_data_7__11), .A1 (
             filter_data_5__11), .S0 (nx1265)) ;
    mux21_ni ix1511 (.Y (ordered_filter_data_5__12), .A0 (filter_data_7__12), .A1 (
             filter_data_5__12), .S0 (nx1265)) ;
    mux21_ni ix1519 (.Y (ordered_filter_data_5__13), .A0 (filter_data_7__13), .A1 (
             filter_data_5__13), .S0 (nx1265)) ;
    mux21_ni ix1527 (.Y (ordered_filter_data_5__14), .A0 (filter_data_7__14), .A1 (
             filter_data_5__14), .S0 (nx1265)) ;
    mux21_ni ix1535 (.Y (ordered_filter_data_5__15), .A0 (filter_data_7__31), .A1 (
             filter_data_5__31), .S0 (nx1265)) ;
    mux21_ni ix1799 (.Y (ordered_filter_data_4__0), .A0 (filter_data_6__0), .A1 (
             filter_data_4__0), .S0 (nx1265)) ;
    mux21_ni ix1807 (.Y (ordered_filter_data_4__1), .A0 (filter_data_6__1), .A1 (
             filter_data_4__1), .S0 (nx1265)) ;
    mux21_ni ix1815 (.Y (ordered_filter_data_4__2), .A0 (filter_data_6__2), .A1 (
             filter_data_4__2), .S0 (nx1267)) ;
    mux21_ni ix1823 (.Y (ordered_filter_data_4__3), .A0 (filter_data_6__3), .A1 (
             filter_data_4__3), .S0 (nx1267)) ;
    mux21_ni ix1831 (.Y (ordered_filter_data_4__4), .A0 (filter_data_6__4), .A1 (
             filter_data_4__4), .S0 (nx1267)) ;
    mux21_ni ix1839 (.Y (ordered_filter_data_4__5), .A0 (filter_data_6__5), .A1 (
             filter_data_4__5), .S0 (nx1267)) ;
    mux21_ni ix1847 (.Y (ordered_filter_data_4__6), .A0 (filter_data_6__6), .A1 (
             filter_data_4__6), .S0 (nx1267)) ;
    mux21_ni ix1855 (.Y (ordered_filter_data_4__7), .A0 (filter_data_6__7), .A1 (
             filter_data_4__7), .S0 (nx1267)) ;
    mux21_ni ix1863 (.Y (ordered_filter_data_4__8), .A0 (filter_data_6__8), .A1 (
             filter_data_4__8), .S0 (nx1267)) ;
    mux21_ni ix1871 (.Y (ordered_filter_data_4__9), .A0 (filter_data_6__9), .A1 (
             filter_data_4__9), .S0 (nx1269)) ;
    mux21_ni ix1879 (.Y (ordered_filter_data_4__10), .A0 (filter_data_6__10), .A1 (
             filter_data_4__10), .S0 (nx1269)) ;
    mux21_ni ix1887 (.Y (ordered_filter_data_4__11), .A0 (filter_data_6__11), .A1 (
             filter_data_4__11), .S0 (nx1269)) ;
    mux21_ni ix1895 (.Y (ordered_filter_data_4__12), .A0 (filter_data_6__12), .A1 (
             filter_data_4__12), .S0 (nx1269)) ;
    mux21_ni ix1903 (.Y (ordered_filter_data_4__13), .A0 (filter_data_6__13), .A1 (
             filter_data_4__13), .S0 (nx1269)) ;
    mux21_ni ix1911 (.Y (ordered_filter_data_4__14), .A0 (filter_data_6__14), .A1 (
             filter_data_4__14), .S0 (nx1269)) ;
    mux21_ni ix1919 (.Y (ordered_filter_data_4__15), .A0 (filter_data_6__31), .A1 (
             filter_data_4__31), .S0 (nx1269)) ;
    mux21_ni ix2183 (.Y (ordered_filter_data_3__0), .A0 (filter_data_5__0), .A1 (
             filter_data_3__0), .S0 (nx1271)) ;
    mux21_ni ix2191 (.Y (ordered_filter_data_3__1), .A0 (filter_data_5__1), .A1 (
             filter_data_3__1), .S0 (nx1271)) ;
    mux21_ni ix2199 (.Y (ordered_filter_data_3__2), .A0 (filter_data_5__2), .A1 (
             filter_data_3__2), .S0 (nx1271)) ;
    mux21_ni ix2207 (.Y (ordered_filter_data_3__3), .A0 (filter_data_5__3), .A1 (
             filter_data_3__3), .S0 (nx1271)) ;
    mux21_ni ix2215 (.Y (ordered_filter_data_3__4), .A0 (filter_data_5__4), .A1 (
             filter_data_3__4), .S0 (nx1271)) ;
    mux21_ni ix2223 (.Y (ordered_filter_data_3__5), .A0 (filter_data_5__5), .A1 (
             filter_data_3__5), .S0 (nx1271)) ;
    mux21_ni ix2231 (.Y (ordered_filter_data_3__6), .A0 (filter_data_5__6), .A1 (
             filter_data_3__6), .S0 (nx1271)) ;
    mux21_ni ix2239 (.Y (ordered_filter_data_3__7), .A0 (filter_data_5__7), .A1 (
             filter_data_3__7), .S0 (nx1273)) ;
    mux21_ni ix2247 (.Y (ordered_filter_data_3__8), .A0 (filter_data_5__8), .A1 (
             filter_data_3__8), .S0 (nx1273)) ;
    mux21_ni ix2255 (.Y (ordered_filter_data_3__9), .A0 (filter_data_5__9), .A1 (
             filter_data_3__9), .S0 (nx1273)) ;
    mux21_ni ix2263 (.Y (ordered_filter_data_3__10), .A0 (filter_data_5__10), .A1 (
             filter_data_3__10), .S0 (nx1273)) ;
    mux21_ni ix2271 (.Y (ordered_filter_data_3__11), .A0 (filter_data_5__11), .A1 (
             filter_data_3__11), .S0 (nx1273)) ;
    mux21_ni ix2279 (.Y (ordered_filter_data_3__12), .A0 (filter_data_5__12), .A1 (
             filter_data_3__12), .S0 (nx1273)) ;
    mux21_ni ix2287 (.Y (ordered_filter_data_3__13), .A0 (filter_data_5__13), .A1 (
             filter_data_3__13), .S0 (nx1273)) ;
    mux21_ni ix2295 (.Y (ordered_filter_data_3__14), .A0 (filter_data_5__14), .A1 (
             filter_data_3__14), .S0 (nx1354)) ;
    mux21_ni ix2303 (.Y (ordered_filter_data_3__15), .A0 (filter_data_5__31), .A1 (
             filter_data_3__31), .S0 (nx1354)) ;
    mux21_ni ix143 (.Y (ordered_img_data_17__1), .A0 (img_data_17__1), .A1 (
             img_data_13__1), .S0 (nx1354)) ;
    mux21_ni ix151 (.Y (ordered_img_data_17__2), .A0 (img_data_17__2), .A1 (
             img_data_13__2), .S0 (nx1354)) ;
    mux21_ni ix159 (.Y (ordered_img_data_17__3), .A0 (img_data_17__3), .A1 (
             img_data_13__3), .S0 (nx1354)) ;
    mux21_ni ix167 (.Y (ordered_img_data_17__4), .A0 (img_data_17__4), .A1 (
             img_data_13__4), .S0 (nx1354)) ;
    mux21_ni ix183 (.Y (ordered_img_data_17__6), .A0 (img_data_17__6), .A1 (
             img_data_13__6), .S0 (nx1354)) ;
    mux21_ni ix191 (.Y (ordered_img_data_17__7), .A0 (img_data_17__7), .A1 (
             img_data_13__7), .S0 (nx1356)) ;
    mux21_ni ix199 (.Y (ordered_img_data_17__8), .A0 (img_data_17__8), .A1 (
             img_data_13__8), .S0 (nx1356)) ;
    mux21_ni ix207 (.Y (ordered_img_data_17__9), .A0 (img_data_17__9), .A1 (
             img_data_13__9), .S0 (nx1356)) ;
    mux21_ni ix215 (.Y (ordered_img_data_17__10), .A0 (img_data_17__10), .A1 (
             img_data_13__10), .S0 (nx1356)) ;
    mux21_ni ix223 (.Y (ordered_img_data_17__11), .A0 (img_data_17__11), .A1 (
             img_data_13__11), .S0 (nx1356)) ;
    mux21_ni ix231 (.Y (ordered_img_data_17__12), .A0 (img_data_17__12), .A1 (
             img_data_13__12), .S0 (nx1356)) ;
    mux21_ni ix239 (.Y (ordered_img_data_17__13), .A0 (img_data_17__13), .A1 (
             img_data_13__13), .S0 (nx1356)) ;
    mux21_ni ix247 (.Y (ordered_img_data_17__14), .A0 (img_data_17__14), .A1 (
             img_data_13__14), .S0 (nx1358)) ;
    mux21_ni ix255 (.Y (ordered_img_data_17__31), .A0 (img_data_17__31), .A1 (
             img_data_13__31), .S0 (nx1358)) ;
    mux21_ni ix519 (.Y (ordered_img_data_16__0), .A0 (img_data_16__0), .A1 (
             img_data_12__0), .S0 (nx1358)) ;
    mux21_ni ix535 (.Y (ordered_img_data_16__2), .A0 (img_data_16__2), .A1 (
             img_data_12__2), .S0 (nx1358)) ;
    mux21_ni ix543 (.Y (ordered_img_data_16__3), .A0 (img_data_16__3), .A1 (
             img_data_12__3), .S0 (nx1358)) ;
    mux21_ni ix551 (.Y (ordered_img_data_16__4), .A0 (img_data_16__4), .A1 (
             img_data_12__4), .S0 (nx1358)) ;
    mux21_ni ix559 (.Y (ordered_img_data_16__5), .A0 (img_data_16__5), .A1 (
             img_data_12__5), .S0 (nx1358)) ;
    mux21_ni ix567 (.Y (ordered_img_data_16__6), .A0 (img_data_16__6), .A1 (
             img_data_12__6), .S0 (nx1361)) ;
    mux21_ni ix583 (.Y (ordered_img_data_16__8), .A0 (img_data_16__8), .A1 (
             img_data_12__8), .S0 (nx1361)) ;
    mux21_ni ix591 (.Y (ordered_img_data_16__9), .A0 (img_data_16__9), .A1 (
             img_data_12__9), .S0 (nx1361)) ;
    mux21_ni ix599 (.Y (ordered_img_data_16__10), .A0 (img_data_16__10), .A1 (
             img_data_12__10), .S0 (nx1361)) ;
    mux21_ni ix607 (.Y (ordered_img_data_16__11), .A0 (img_data_16__11), .A1 (
             img_data_12__11), .S0 (nx1361)) ;
    mux21_ni ix615 (.Y (ordered_img_data_16__12), .A0 (img_data_16__12), .A1 (
             img_data_12__12), .S0 (nx1361)) ;
    mux21_ni ix623 (.Y (ordered_img_data_16__13), .A0 (img_data_16__13), .A1 (
             img_data_12__13), .S0 (nx1361)) ;
    mux21_ni ix631 (.Y (ordered_img_data_16__14), .A0 (img_data_16__14), .A1 (
             img_data_12__14), .S0 (nx1363)) ;
    mux21_ni ix639 (.Y (ordered_img_data_16__31), .A0 (img_data_16__31), .A1 (
             img_data_12__31), .S0 (nx1363)) ;
    mux21_ni ix911 (.Y (ordered_img_data_15__1), .A0 (img_data_15__1), .A1 (
             img_data_11__1), .S0 (nx1363)) ;
    mux21_ni ix919 (.Y (ordered_img_data_15__2), .A0 (img_data_15__2), .A1 (
             img_data_11__2), .S0 (nx1363)) ;
    mux21_ni ix927 (.Y (ordered_img_data_15__3), .A0 (img_data_15__3), .A1 (
             img_data_11__3), .S0 (nx1363)) ;
    mux21_ni ix935 (.Y (ordered_img_data_15__4), .A0 (img_data_15__4), .A1 (
             img_data_11__4), .S0 (nx1363)) ;
    mux21_ni ix943 (.Y (ordered_img_data_15__5), .A0 (img_data_15__5), .A1 (
             img_data_11__5), .S0 (nx1363)) ;
    mux21_ni ix951 (.Y (ordered_img_data_15__6), .A0 (img_data_15__6), .A1 (
             img_data_11__6), .S0 (nx1365)) ;
    mux21_ni ix967 (.Y (ordered_img_data_15__8), .A0 (img_data_15__8), .A1 (
             img_data_11__8), .S0 (nx1287)) ;
    mux21_ni ix975 (.Y (ordered_img_data_15__9), .A0 (img_data_15__9), .A1 (
             img_data_11__9), .S0 (nx1287)) ;
    mux21_ni ix983 (.Y (ordered_img_data_15__10), .A0 (img_data_15__10), .A1 (
             img_data_11__10), .S0 (nx1287)) ;
    mux21_ni ix991 (.Y (ordered_img_data_15__11), .A0 (img_data_15__11), .A1 (
             img_data_11__11), .S0 (nx1287)) ;
    mux21_ni ix999 (.Y (ordered_img_data_15__12), .A0 (img_data_15__12), .A1 (
             img_data_11__12), .S0 (nx1287)) ;
    mux21_ni ix1007 (.Y (ordered_img_data_15__13), .A0 (img_data_15__13), .A1 (
             img_data_11__13), .S0 (nx1287)) ;
    mux21_ni ix1015 (.Y (ordered_img_data_15__14), .A0 (img_data_15__14), .A1 (
             img_data_11__14), .S0 (nx1287)) ;
    mux21_ni ix1023 (.Y (ordered_img_data_15__31), .A0 (img_data_15__31), .A1 (
             img_data_11__31), .S0 (nx1365)) ;
    mux21_ni ix1287 (.Y (ordered_img_data_14__0), .A0 (img_data_14__0), .A1 (
             img_data_8__0), .S0 (nx1365)) ;
    mux21_ni ix1295 (.Y (ordered_img_data_14__1), .A0 (img_data_14__1), .A1 (
             img_data_8__1), .S0 (nx1365)) ;
    mux21_ni ix1303 (.Y (ordered_img_data_14__2), .A0 (img_data_14__2), .A1 (
             img_data_8__2), .S0 (nx1365)) ;
    mux21_ni ix1319 (.Y (ordered_img_data_14__4), .A0 (img_data_14__4), .A1 (
             img_data_8__4), .S0 (nx1365)) ;
    mux21_ni ix1327 (.Y (ordered_img_data_14__5), .A0 (img_data_14__5), .A1 (
             img_data_8__5), .S0 (nx1365)) ;
    mux21_ni ix1335 (.Y (ordered_img_data_14__6), .A0 (img_data_14__6), .A1 (
             img_data_8__6), .S0 (nx1367)) ;
    mux21_ni ix1351 (.Y (ordered_img_data_14__8), .A0 (img_data_14__8), .A1 (
             img_data_8__8), .S0 (nx1367)) ;
    mux21_ni ix1359 (.Y (ordered_img_data_14__9), .A0 (img_data_14__9), .A1 (
             img_data_8__9), .S0 (nx1367)) ;
    mux21_ni ix1367 (.Y (ordered_img_data_14__10), .A0 (img_data_14__10), .A1 (
             img_data_8__10), .S0 (nx1367)) ;
    mux21_ni ix1375 (.Y (ordered_img_data_14__11), .A0 (img_data_14__11), .A1 (
             img_data_8__11), .S0 (nx1367)) ;
    mux21_ni ix1383 (.Y (ordered_img_data_14__12), .A0 (img_data_14__12), .A1 (
             img_data_8__12), .S0 (nx1367)) ;
    mux21_ni ix1391 (.Y (ordered_img_data_14__13), .A0 (img_data_14__13), .A1 (
             img_data_8__13), .S0 (nx1367)) ;
    mux21_ni ix1399 (.Y (ordered_img_data_14__14), .A0 (img_data_14__14), .A1 (
             img_data_8__14), .S0 (nx1369)) ;
    mux21_ni ix1407 (.Y (ordered_img_data_14__31), .A0 (img_data_14__31), .A1 (
             img_data_8__31), .S0 (nx1369)) ;
    mux21_ni ix1671 (.Y (ordered_img_data_13__0), .A0 (img_data_9__0), .A1 (
             img_data_7__0), .S0 (nx1369)) ;
    mux21_ni ix1679 (.Y (ordered_img_data_13__1), .A0 (img_data_9__1), .A1 (
             img_data_7__1), .S0 (nx1369)) ;
    mux21_ni ix1687 (.Y (ordered_img_data_13__2), .A0 (img_data_9__2), .A1 (
             img_data_7__2), .S0 (nx1369)) ;
    mux21_ni ix1703 (.Y (ordered_img_data_13__4), .A0 (img_data_9__4), .A1 (
             img_data_7__4), .S0 (nx1369)) ;
    mux21_ni ix1719 (.Y (ordered_img_data_13__6), .A0 (img_data_9__6), .A1 (
             img_data_7__6), .S0 (nx1369)) ;
    mux21_ni ix1727 (.Y (ordered_img_data_13__7), .A0 (img_data_9__7), .A1 (
             img_data_7__7), .S0 (nx1371)) ;
    mux21_ni ix1735 (.Y (ordered_img_data_13__8), .A0 (img_data_9__8), .A1 (
             img_data_7__8), .S0 (nx1371)) ;
    mux21_ni ix1743 (.Y (ordered_img_data_13__9), .A0 (img_data_9__9), .A1 (
             img_data_7__9), .S0 (nx1371)) ;
    mux21_ni ix1751 (.Y (ordered_img_data_13__10), .A0 (img_data_9__10), .A1 (
             img_data_7__10), .S0 (nx1371)) ;
    mux21_ni ix1759 (.Y (ordered_img_data_13__11), .A0 (img_data_9__11), .A1 (
             img_data_7__11), .S0 (nx1371)) ;
    mux21_ni ix1767 (.Y (ordered_img_data_13__12), .A0 (img_data_9__12), .A1 (
             img_data_7__12), .S0 (nx1371)) ;
    mux21_ni ix1775 (.Y (ordered_img_data_13__13), .A0 (img_data_9__13), .A1 (
             img_data_7__13), .S0 (nx1371)) ;
    mux21_ni ix1783 (.Y (ordered_img_data_13__14), .A0 (img_data_9__14), .A1 (
             img_data_7__14), .S0 (nx1373)) ;
    mux21_ni ix1791 (.Y (ordered_img_data_13__31), .A0 (img_data_9__31), .A1 (
             img_data_7__31), .S0 (nx1373)) ;
    mux21_ni ix2063 (.Y (ordered_img_data_12__1), .A0 (img_data_4__1), .A1 (
             img_data_6__1), .S0 (nx1373)) ;
    mux21_ni ix2071 (.Y (ordered_img_data_12__2), .A0 (img_data_4__2), .A1 (
             img_data_6__2), .S0 (nx1373)) ;
    mux21_ni ix2079 (.Y (ordered_img_data_12__3), .A0 (img_data_4__3), .A1 (
             img_data_6__3), .S0 (nx1373)) ;
    mux21_ni ix2095 (.Y (ordered_img_data_12__5), .A0 (img_data_4__5), .A1 (
             img_data_6__5), .S0 (nx1373)) ;
    mux21_ni ix2103 (.Y (ordered_img_data_12__6), .A0 (img_data_4__6), .A1 (
             img_data_6__6), .S0 (nx1373)) ;
    mux21_ni ix2111 (.Y (ordered_img_data_12__7), .A0 (img_data_4__7), .A1 (
             img_data_6__7), .S0 (nx1375)) ;
    mux21_ni ix2119 (.Y (ordered_img_data_12__8), .A0 (img_data_4__8), .A1 (
             img_data_6__8), .S0 (nx1375)) ;
    mux21_ni ix2127 (.Y (ordered_img_data_12__9), .A0 (img_data_4__9), .A1 (
             img_data_6__9), .S0 (nx1301)) ;
    mux21_ni ix2135 (.Y (ordered_img_data_12__10), .A0 (img_data_4__10), .A1 (
             img_data_6__10), .S0 (nx1301)) ;
    mux21_ni ix2143 (.Y (ordered_img_data_12__11), .A0 (img_data_4__11), .A1 (
             img_data_6__11), .S0 (nx1301)) ;
    mux21_ni ix2151 (.Y (ordered_img_data_12__12), .A0 (img_data_4__12), .A1 (
             img_data_6__12), .S0 (nx1301)) ;
    mux21_ni ix2159 (.Y (ordered_img_data_12__13), .A0 (img_data_4__13), .A1 (
             img_data_6__13), .S0 (nx1301)) ;
    mux21_ni ix2167 (.Y (ordered_img_data_12__14), .A0 (img_data_4__14), .A1 (
             img_data_6__14), .S0 (nx1301)) ;
    mux21_ni ix2175 (.Y (ordered_img_data_12__31), .A0 (img_data_4__31), .A1 (
             img_data_6__31), .S0 (nx1301)) ;
    mux21_ni ix2439 (.Y (ordered_img_data_11__0), .A0 (img_data_13__0), .A1 (
             img_data_3__0), .S0 (nx1375)) ;
    mux21_ni ix2447 (.Y (ordered_img_data_11__1), .A0 (img_data_13__1), .A1 (
             img_data_3__1), .S0 (nx1375)) ;
    mux21_ni ix2463 (.Y (ordered_img_data_11__3), .A0 (img_data_13__3), .A1 (
             img_data_3__3), .S0 (nx1375)) ;
    mux21_ni ix2471 (.Y (ordered_img_data_11__4), .A0 (img_data_13__4), .A1 (
             img_data_3__4), .S0 (nx1375)) ;
    mux21_ni ix2479 (.Y (ordered_img_data_11__5), .A0 (img_data_13__5), .A1 (
             img_data_3__5), .S0 (nx1375)) ;
    mux21_ni ix2487 (.Y (ordered_img_data_11__6), .A0 (img_data_13__6), .A1 (
             img_data_3__6), .S0 (nx1377)) ;
    mux21_ni ix2503 (.Y (ordered_img_data_11__8), .A0 (img_data_13__8), .A1 (
             img_data_3__8), .S0 (nx1377)) ;
    mux21_ni ix2511 (.Y (ordered_img_data_11__9), .A0 (img_data_13__9), .A1 (
             img_data_3__9), .S0 (nx1377)) ;
    mux21_ni ix2519 (.Y (ordered_img_data_11__10), .A0 (img_data_13__10), .A1 (
             img_data_3__10), .S0 (nx1377)) ;
    mux21_ni ix2527 (.Y (ordered_img_data_11__11), .A0 (img_data_13__11), .A1 (
             img_data_3__11), .S0 (nx1377)) ;
    mux21_ni ix2535 (.Y (ordered_img_data_11__12), .A0 (img_data_13__12), .A1 (
             img_data_3__12), .S0 (nx1377)) ;
    mux21_ni ix2543 (.Y (ordered_img_data_11__13), .A0 (img_data_13__13), .A1 (
             img_data_3__13), .S0 (nx1377)) ;
    mux21_ni ix2551 (.Y (ordered_img_data_11__14), .A0 (img_data_13__14), .A1 (
             img_data_3__14), .S0 (nx1379)) ;
    mux21_ni ix2559 (.Y (ordered_img_data_11__31), .A0 (img_data_13__31), .A1 (
             img_data_3__31), .S0 (nx1379)) ;
    mux21_ni ix2695 (.Y (ordered_img_data_10__0), .A0 (img_data_8__0), .A1 (
             img_data_2__0), .S0 (nx1379)) ;
    mux21_ni ix2711 (.Y (ordered_img_data_10__2), .A0 (img_data_8__2), .A1 (
             img_data_2__2), .S0 (nx1379)) ;
    mux21_ni ix2719 (.Y (ordered_img_data_10__3), .A0 (img_data_8__3), .A1 (
             img_data_2__3), .S0 (nx1379)) ;
    mux21_ni ix2727 (.Y (ordered_img_data_10__4), .A0 (img_data_8__4), .A1 (
             img_data_2__4), .S0 (nx1379)) ;
    mux21_ni ix2735 (.Y (ordered_img_data_10__5), .A0 (img_data_8__5), .A1 (
             img_data_2__5), .S0 (nx1379)) ;
    mux21_ni ix2743 (.Y (ordered_img_data_10__6), .A0 (img_data_8__6), .A1 (
             img_data_2__6), .S0 (nx1381)) ;
    mux21_ni ix2759 (.Y (ordered_img_data_10__8), .A0 (img_data_8__8), .A1 (
             img_data_2__8), .S0 (nx1381)) ;
    mux21_ni ix2767 (.Y (ordered_img_data_10__9), .A0 (img_data_8__9), .A1 (
             img_data_2__9), .S0 (nx1381)) ;
    mux21_ni ix2775 (.Y (ordered_img_data_10__10), .A0 (img_data_8__10), .A1 (
             img_data_2__10), .S0 (nx1381)) ;
    mux21_ni ix2783 (.Y (ordered_img_data_10__11), .A0 (img_data_8__11), .A1 (
             img_data_2__11), .S0 (nx1381)) ;
    mux21_ni ix2791 (.Y (ordered_img_data_10__12), .A0 (img_data_8__12), .A1 (
             img_data_2__12), .S0 (nx1381)) ;
    mux21_ni ix2799 (.Y (ordered_img_data_10__13), .A0 (img_data_8__13), .A1 (
             img_data_2__13), .S0 (nx1381)) ;
    mux21_ni ix2807 (.Y (ordered_img_data_10__14), .A0 (img_data_8__14), .A1 (
             img_data_2__14), .S0 (nx1383)) ;
    mux21_ni ix2815 (.Y (ordered_img_data_10__31), .A0 (img_data_8__31), .A1 (
             img_data_2__31), .S0 (nx1383)) ;
    mux21_ni ix2959 (.Y (ordered_img_data_9__1), .A0 (img_data_3__1), .A1 (
             img_data_1__1), .S0 (nx1383)) ;
    mux21_ni ix2967 (.Y (ordered_img_data_9__2), .A0 (img_data_3__2), .A1 (
             img_data_1__2), .S0 (nx1383)) ;
    mux21_ni ix2975 (.Y (ordered_img_data_9__3), .A0 (img_data_3__3), .A1 (
             img_data_1__3), .S0 (nx1383)) ;
    mux21_ni ix2983 (.Y (ordered_img_data_9__4), .A0 (img_data_3__4), .A1 (
             img_data_1__4), .S0 (nx1383)) ;
    mux21_ni ix2991 (.Y (ordered_img_data_9__5), .A0 (img_data_3__5), .A1 (
             img_data_1__5), .S0 (nx1383)) ;
    mux21_ni ix2999 (.Y (ordered_img_data_9__6), .A0 (img_data_3__6), .A1 (
             img_data_1__6), .S0 (nx1385)) ;
    mux21_ni ix3015 (.Y (ordered_img_data_9__8), .A0 (img_data_3__8), .A1 (
             img_data_1__8), .S0 (nx1385)) ;
    mux21_ni ix3023 (.Y (ordered_img_data_9__9), .A0 (img_data_3__9), .A1 (
             img_data_1__9), .S0 (nx1385)) ;
    mux21_ni ix3031 (.Y (ordered_img_data_9__10), .A0 (img_data_3__10), .A1 (
             img_data_1__10), .S0 (nx1315)) ;
    mux21_ni ix3039 (.Y (ordered_img_data_9__11), .A0 (img_data_3__11), .A1 (
             img_data_1__11), .S0 (nx1315)) ;
    mux21_ni ix3047 (.Y (ordered_img_data_9__12), .A0 (img_data_3__12), .A1 (
             img_data_1__12), .S0 (nx1315)) ;
    mux21_ni ix3055 (.Y (ordered_img_data_9__13), .A0 (img_data_3__13), .A1 (
             img_data_1__13), .S0 (nx1315)) ;
    mux21_ni ix3063 (.Y (ordered_img_data_9__14), .A0 (img_data_3__14), .A1 (
             img_data_1__14), .S0 (nx1315)) ;
    mux21_ni ix3071 (.Y (ordered_img_data_9__31), .A0 (img_data_3__31), .A1 (
             img_data_1__31), .S0 (nx1315)) ;
    inv02 ix1205 (.Y (nx1206), .A (nx1317)) ;
    inv02 ix1208 (.Y (nx1209), .A (nx1317)) ;
    inv02 ix1210 (.Y (nx1211), .A (nx1317)) ;
    inv02 ix1212 (.Y (nx1213), .A (nx1317)) ;
    inv02 ix1214 (.Y (nx1215), .A (nx1317)) ;
    inv02 ix1216 (.Y (nx1217), .A (nx1317)) ;
    inv02 ix1218 (.Y (nx1219), .A (nx1317)) ;
    inv02 ix1220 (.Y (nx1221), .A (nx1319)) ;
    inv02 ix1222 (.Y (nx1223), .A (nx1319)) ;
    inv02 ix1224 (.Y (nx1225), .A (nx1319)) ;
    inv02 ix1226 (.Y (nx1227), .A (nx1319)) ;
    inv02 ix1228 (.Y (nx1229), .A (nx1319)) ;
    inv02 ix1230 (.Y (nx1231), .A (nx1319)) ;
    inv02 ix1232 (.Y (nx1233), .A (nx1319)) ;
    inv02 ix1234 (.Y (nx1235), .A (nx1321)) ;
    inv02 ix1236 (.Y (nx1237), .A (nx1321)) ;
    inv02 ix1238 (.Y (nx1239), .A (nx1321)) ;
    inv02 ix1240 (.Y (nx1241), .A (nx1321)) ;
    inv02 ix1242 (.Y (nx1243), .A (nx1321)) ;
    inv02 ix1244 (.Y (nx1245), .A (nx1321)) ;
    inv02 ix1246 (.Y (nx1247), .A (nx1321)) ;
    inv02 ix1248 (.Y (nx1249), .A (nx1323)) ;
    inv02 ix1250 (.Y (nx1251), .A (nx1323)) ;
    inv02 ix1252 (.Y (nx1253), .A (nx1323)) ;
    inv02 ix1254 (.Y (nx1255), .A (nx1323)) ;
    inv02 ix1256 (.Y (nx1257), .A (nx1323)) ;
    inv02 ix1258 (.Y (nx1259), .A (nx1323)) ;
    inv02 ix1260 (.Y (nx1261), .A (nx1323)) ;
    inv02 ix1262 (.Y (nx1263), .A (nx1325)) ;
    inv02 ix1264 (.Y (nx1265), .A (nx1325)) ;
    inv02 ix1266 (.Y (nx1267), .A (nx1325)) ;
    inv02 ix1268 (.Y (nx1269), .A (nx1325)) ;
    inv02 ix1270 (.Y (nx1271), .A (nx1325)) ;
    inv02 ix1272 (.Y (nx1273), .A (nx1325)) ;
    inv02 ix1286 (.Y (nx1287), .A (nx1345)) ;
    inv02 ix1300 (.Y (nx1301), .A (nx1345)) ;
    inv02 ix1314 (.Y (nx1315), .A (nx1331)) ;
    inv02 ix1318 (.Y (nx1319), .A (filter_size)) ;
    inv02 ix1320 (.Y (nx1321), .A (nx1385)) ;
    inv02 ix1322 (.Y (nx1323), .A (nx1385)) ;
    inv02 ix1316 (.Y (nx1317), .A (nx1385)) ;
    ao22 reg_ordered_img_data_14__3 (.Y (ordered_img_data_14__3), .A0 (
         img_data_14__3), .A1 (nx1345), .B0 (img_data_8__3), .B1 (nx1385)) ;
    ao22 reg_ordered_img_data_12__4 (.Y (ordered_img_data_12__4), .A0 (
         img_data_4__4), .A1 (nx1345), .B0 (img_data_6__4), .B1 (nx1387)) ;
    ao22 reg_ordered_img_data_13__3 (.Y (ordered_img_data_13__3), .A0 (
         img_data_9__3), .A1 (nx1345), .B0 (img_data_7__3), .B1 (nx1387)) ;
    ao22 reg_ordered_img_data_13__5 (.Y (ordered_img_data_13__5), .A0 (
         img_data_9__5), .A1 (nx1345), .B0 (img_data_7__5), .B1 (nx1387)) ;
    ao22 reg_ordered_img_data_14__7 (.Y (ordered_img_data_14__7), .A0 (
         img_data_14__7), .A1 (nx1345), .B0 (img_data_8__7), .B1 (nx1387)) ;
    ao22 reg_ordered_img_data_12__0 (.Y (ordered_img_data_12__0), .A0 (
         img_data_4__0), .A1 (nx1346), .B0 (img_data_6__0), .B1 (nx1387)) ;
    ao22 reg_ordered_img_data_15__7 (.Y (ordered_img_data_15__7), .A0 (
         img_data_15__7), .A1 (nx1346), .B0 (img_data_11__7), .B1 (nx1387)) ;
    ao22 reg_ordered_img_data_11__2 (.Y (ordered_img_data_11__2), .A0 (
         img_data_13__2), .A1 (nx1346), .B0 (img_data_3__2), .B1 (nx1387)) ;
    ao22 reg_ordered_img_data_15__0 (.Y (ordered_img_data_15__0), .A0 (
         img_data_15__0), .A1 (nx1346), .B0 (img_data_11__0), .B1 (nx1389)) ;
    ao22 reg_ordered_img_data_16__7 (.Y (ordered_img_data_16__7), .A0 (
         img_data_16__7), .A1 (nx1346), .B0 (img_data_12__7), .B1 (nx1389)) ;
    ao22 reg_ordered_img_data_17__5 (.Y (ordered_img_data_17__5), .A0 (
         img_data_17__5), .A1 (nx1346), .B0 (img_data_13__5), .B1 (nx1389)) ;
    inv01 reg_nx1317_XX0_XREP32 (.Y (nx1317_XX0_XREP32), .A (nx1389)) ;
    ao22 reg_ordered_img_data_16__1 (.Y (ordered_img_data_16__1), .A0 (
         img_data_16__1), .A1 (nx1346), .B0 (img_data_12__1), .B1 (nx1389)) ;
    inv02 reg_nx1325 (.Y (nx1325), .A (nx1391)) ;
    ao22 reg_ordered_img_data_17__0 (.Y (ordered_img_data_17__0), .A0 (
         img_data_17__0), .A1 (nx1325), .B0 (img_data_13__0), .B1 (nx1389)) ;
    ao22 reg_ordered_img_data_9__7 (.Y (ordered_img_data_9__7), .A0 (
         img_data_3__7), .A1 (nx1331), .B0 (img_data_1__7), .B1 (nx1389)) ;
    ao22 reg_ordered_img_data_10__1 (.Y (ordered_img_data_10__1), .A0 (
         img_data_8__1), .A1 (nx1331), .B0 (img_data_2__1), .B1 (nx1391)) ;
    ao22 reg_ordered_img_data_10__7 (.Y (ordered_img_data_10__7), .A0 (
         img_data_8__7), .A1 (nx1331), .B0 (img_data_2__7), .B1 (nx1391)) ;
    ao22 reg_ordered_img_data_11__7 (.Y (ordered_img_data_11__7), .A0 (
         img_data_13__7), .A1 (nx1331), .B0 (img_data_3__7), .B1 (nx1391)) ;
    inv01 reg_nx1331 (.Y (nx1331), .A (nx1391)) ;
    ao22 reg_ordered_img_data_9__0 (.Y (ordered_img_data_9__0), .A0 (
         img_data_3__0), .A1 (nx1331), .B0 (img_data_1__0), .B1 (nx1391)) ;
    buf16 ix1347 (.Y (nx1345), .A (nx1317_XX0_XREP32)) ;
    buf16 ix1348 (.Y (nx1346), .A (nx1317_XX0_XREP32)) ;
    inv02 ix1353 (.Y (nx1354), .A (nx1319)) ;
    inv02 ix1355 (.Y (nx1356), .A (nx1319)) ;
    inv02 ix1357 (.Y (nx1358), .A (nx1319)) ;
    inv02 ix1360 (.Y (nx1361), .A (nx1319)) ;
    inv02 ix1362 (.Y (nx1363), .A (nx1319)) ;
    inv02 ix1364 (.Y (nx1365), .A (nx1319)) ;
    inv02 ix1366 (.Y (nx1367), .A (nx1319)) ;
    inv02 ix1368 (.Y (nx1369), .A (nx1319)) ;
    inv02 ix1370 (.Y (nx1371), .A (nx1319)) ;
    inv02 ix1372 (.Y (nx1373), .A (nx1319)) ;
    inv02 ix1374 (.Y (nx1375), .A (nx1319)) ;
    inv02 ix1376 (.Y (nx1377), .A (nx1319)) ;
    inv02 ix1378 (.Y (nx1379), .A (nx1319)) ;
    inv02 ix1380 (.Y (nx1381), .A (nx1319)) ;
    inv02 ix1382 (.Y (nx1383), .A (nx1319)) ;
    inv02 ix1384 (.Y (nx1385), .A (nx1319)) ;
    inv02 ix1386 (.Y (nx1387), .A (nx1319)) ;
    inv02 ix1388 (.Y (nx1389), .A (nx1319)) ;
    inv02 ix1390 (.Y (nx1391), .A (nx1319)) ;
endmodule


module CacheMuxer ( d_arr_mux_0__31, d_arr_mux_0__30, d_arr_mux_0__29, 
                    d_arr_mux_0__28, d_arr_mux_0__27, d_arr_mux_0__26, 
                    d_arr_mux_0__25, d_arr_mux_0__24, d_arr_mux_0__23, 
                    d_arr_mux_0__22, d_arr_mux_0__21, d_arr_mux_0__20, 
                    d_arr_mux_0__19, d_arr_mux_0__18, d_arr_mux_0__17, 
                    d_arr_mux_0__16, d_arr_mux_0__15, d_arr_mux_0__14, 
                    d_arr_mux_0__13, d_arr_mux_0__12, d_arr_mux_0__11, 
                    d_arr_mux_0__10, d_arr_mux_0__9, d_arr_mux_0__8, 
                    d_arr_mux_0__7, d_arr_mux_0__6, d_arr_mux_0__5, 
                    d_arr_mux_0__4, d_arr_mux_0__3, d_arr_mux_0__2, 
                    d_arr_mux_0__1, d_arr_mux_0__0, d_arr_mux_1__31, 
                    d_arr_mux_1__30, d_arr_mux_1__29, d_arr_mux_1__28, 
                    d_arr_mux_1__27, d_arr_mux_1__26, d_arr_mux_1__25, 
                    d_arr_mux_1__24, d_arr_mux_1__23, d_arr_mux_1__22, 
                    d_arr_mux_1__21, d_arr_mux_1__20, d_arr_mux_1__19, 
                    d_arr_mux_1__18, d_arr_mux_1__17, d_arr_mux_1__16, 
                    d_arr_mux_1__15, d_arr_mux_1__14, d_arr_mux_1__13, 
                    d_arr_mux_1__12, d_arr_mux_1__11, d_arr_mux_1__10, 
                    d_arr_mux_1__9, d_arr_mux_1__8, d_arr_mux_1__7, 
                    d_arr_mux_1__6, d_arr_mux_1__5, d_arr_mux_1__4, 
                    d_arr_mux_1__3, d_arr_mux_1__2, d_arr_mux_1__1, 
                    d_arr_mux_1__0, d_arr_mux_2__31, d_arr_mux_2__30, 
                    d_arr_mux_2__29, d_arr_mux_2__28, d_arr_mux_2__27, 
                    d_arr_mux_2__26, d_arr_mux_2__25, d_arr_mux_2__24, 
                    d_arr_mux_2__23, d_arr_mux_2__22, d_arr_mux_2__21, 
                    d_arr_mux_2__20, d_arr_mux_2__19, d_arr_mux_2__18, 
                    d_arr_mux_2__17, d_arr_mux_2__16, d_arr_mux_2__15, 
                    d_arr_mux_2__14, d_arr_mux_2__13, d_arr_mux_2__12, 
                    d_arr_mux_2__11, d_arr_mux_2__10, d_arr_mux_2__9, 
                    d_arr_mux_2__8, d_arr_mux_2__7, d_arr_mux_2__6, 
                    d_arr_mux_2__5, d_arr_mux_2__4, d_arr_mux_2__3, 
                    d_arr_mux_2__2, d_arr_mux_2__1, d_arr_mux_2__0, 
                    d_arr_mux_3__31, d_arr_mux_3__30, d_arr_mux_3__29, 
                    d_arr_mux_3__28, d_arr_mux_3__27, d_arr_mux_3__26, 
                    d_arr_mux_3__25, d_arr_mux_3__24, d_arr_mux_3__23, 
                    d_arr_mux_3__22, d_arr_mux_3__21, d_arr_mux_3__20, 
                    d_arr_mux_3__19, d_arr_mux_3__18, d_arr_mux_3__17, 
                    d_arr_mux_3__16, d_arr_mux_3__15, d_arr_mux_3__14, 
                    d_arr_mux_3__13, d_arr_mux_3__12, d_arr_mux_3__11, 
                    d_arr_mux_3__10, d_arr_mux_3__9, d_arr_mux_3__8, 
                    d_arr_mux_3__7, d_arr_mux_3__6, d_arr_mux_3__5, 
                    d_arr_mux_3__4, d_arr_mux_3__3, d_arr_mux_3__2, 
                    d_arr_mux_3__1, d_arr_mux_3__0, d_arr_mux_4__31, 
                    d_arr_mux_4__30, d_arr_mux_4__29, d_arr_mux_4__28, 
                    d_arr_mux_4__27, d_arr_mux_4__26, d_arr_mux_4__25, 
                    d_arr_mux_4__24, d_arr_mux_4__23, d_arr_mux_4__22, 
                    d_arr_mux_4__21, d_arr_mux_4__20, d_arr_mux_4__19, 
                    d_arr_mux_4__18, d_arr_mux_4__17, d_arr_mux_4__16, 
                    d_arr_mux_4__15, d_arr_mux_4__14, d_arr_mux_4__13, 
                    d_arr_mux_4__12, d_arr_mux_4__11, d_arr_mux_4__10, 
                    d_arr_mux_4__9, d_arr_mux_4__8, d_arr_mux_4__7, 
                    d_arr_mux_4__6, d_arr_mux_4__5, d_arr_mux_4__4, 
                    d_arr_mux_4__3, d_arr_mux_4__2, d_arr_mux_4__1, 
                    d_arr_mux_4__0, d_arr_mux_5__31, d_arr_mux_5__30, 
                    d_arr_mux_5__29, d_arr_mux_5__28, d_arr_mux_5__27, 
                    d_arr_mux_5__26, d_arr_mux_5__25, d_arr_mux_5__24, 
                    d_arr_mux_5__23, d_arr_mux_5__22, d_arr_mux_5__21, 
                    d_arr_mux_5__20, d_arr_mux_5__19, d_arr_mux_5__18, 
                    d_arr_mux_5__17, d_arr_mux_5__16, d_arr_mux_5__15, 
                    d_arr_mux_5__14, d_arr_mux_5__13, d_arr_mux_5__12, 
                    d_arr_mux_5__11, d_arr_mux_5__10, d_arr_mux_5__9, 
                    d_arr_mux_5__8, d_arr_mux_5__7, d_arr_mux_5__6, 
                    d_arr_mux_5__5, d_arr_mux_5__4, d_arr_mux_5__3, 
                    d_arr_mux_5__2, d_arr_mux_5__1, d_arr_mux_5__0, 
                    d_arr_mux_6__31, d_arr_mux_6__30, d_arr_mux_6__29, 
                    d_arr_mux_6__28, d_arr_mux_6__27, d_arr_mux_6__26, 
                    d_arr_mux_6__25, d_arr_mux_6__24, d_arr_mux_6__23, 
                    d_arr_mux_6__22, d_arr_mux_6__21, d_arr_mux_6__20, 
                    d_arr_mux_6__19, d_arr_mux_6__18, d_arr_mux_6__17, 
                    d_arr_mux_6__16, d_arr_mux_6__15, d_arr_mux_6__14, 
                    d_arr_mux_6__13, d_arr_mux_6__12, d_arr_mux_6__11, 
                    d_arr_mux_6__10, d_arr_mux_6__9, d_arr_mux_6__8, 
                    d_arr_mux_6__7, d_arr_mux_6__6, d_arr_mux_6__5, 
                    d_arr_mux_6__4, d_arr_mux_6__3, d_arr_mux_6__2, 
                    d_arr_mux_6__1, d_arr_mux_6__0, d_arr_mux_7__31, 
                    d_arr_mux_7__30, d_arr_mux_7__29, d_arr_mux_7__28, 
                    d_arr_mux_7__27, d_arr_mux_7__26, d_arr_mux_7__25, 
                    d_arr_mux_7__24, d_arr_mux_7__23, d_arr_mux_7__22, 
                    d_arr_mux_7__21, d_arr_mux_7__20, d_arr_mux_7__19, 
                    d_arr_mux_7__18, d_arr_mux_7__17, d_arr_mux_7__16, 
                    d_arr_mux_7__15, d_arr_mux_7__14, d_arr_mux_7__13, 
                    d_arr_mux_7__12, d_arr_mux_7__11, d_arr_mux_7__10, 
                    d_arr_mux_7__9, d_arr_mux_7__8, d_arr_mux_7__7, 
                    d_arr_mux_7__6, d_arr_mux_7__5, d_arr_mux_7__4, 
                    d_arr_mux_7__3, d_arr_mux_7__2, d_arr_mux_7__1, 
                    d_arr_mux_7__0, d_arr_mux_8__31, d_arr_mux_8__30, 
                    d_arr_mux_8__29, d_arr_mux_8__28, d_arr_mux_8__27, 
                    d_arr_mux_8__26, d_arr_mux_8__25, d_arr_mux_8__24, 
                    d_arr_mux_8__23, d_arr_mux_8__22, d_arr_mux_8__21, 
                    d_arr_mux_8__20, d_arr_mux_8__19, d_arr_mux_8__18, 
                    d_arr_mux_8__17, d_arr_mux_8__16, d_arr_mux_8__15, 
                    d_arr_mux_8__14, d_arr_mux_8__13, d_arr_mux_8__12, 
                    d_arr_mux_8__11, d_arr_mux_8__10, d_arr_mux_8__9, 
                    d_arr_mux_8__8, d_arr_mux_8__7, d_arr_mux_8__6, 
                    d_arr_mux_8__5, d_arr_mux_8__4, d_arr_mux_8__3, 
                    d_arr_mux_8__2, d_arr_mux_8__1, d_arr_mux_8__0, 
                    d_arr_mux_9__31, d_arr_mux_9__30, d_arr_mux_9__29, 
                    d_arr_mux_9__28, d_arr_mux_9__27, d_arr_mux_9__26, 
                    d_arr_mux_9__25, d_arr_mux_9__24, d_arr_mux_9__23, 
                    d_arr_mux_9__22, d_arr_mux_9__21, d_arr_mux_9__20, 
                    d_arr_mux_9__19, d_arr_mux_9__18, d_arr_mux_9__17, 
                    d_arr_mux_9__16, d_arr_mux_9__15, d_arr_mux_9__14, 
                    d_arr_mux_9__13, d_arr_mux_9__12, d_arr_mux_9__11, 
                    d_arr_mux_9__10, d_arr_mux_9__9, d_arr_mux_9__8, 
                    d_arr_mux_9__7, d_arr_mux_9__6, d_arr_mux_9__5, 
                    d_arr_mux_9__4, d_arr_mux_9__3, d_arr_mux_9__2, 
                    d_arr_mux_9__1, d_arr_mux_9__0, d_arr_mux_10__31, 
                    d_arr_mux_10__30, d_arr_mux_10__29, d_arr_mux_10__28, 
                    d_arr_mux_10__27, d_arr_mux_10__26, d_arr_mux_10__25, 
                    d_arr_mux_10__24, d_arr_mux_10__23, d_arr_mux_10__22, 
                    d_arr_mux_10__21, d_arr_mux_10__20, d_arr_mux_10__19, 
                    d_arr_mux_10__18, d_arr_mux_10__17, d_arr_mux_10__16, 
                    d_arr_mux_10__15, d_arr_mux_10__14, d_arr_mux_10__13, 
                    d_arr_mux_10__12, d_arr_mux_10__11, d_arr_mux_10__10, 
                    d_arr_mux_10__9, d_arr_mux_10__8, d_arr_mux_10__7, 
                    d_arr_mux_10__6, d_arr_mux_10__5, d_arr_mux_10__4, 
                    d_arr_mux_10__3, d_arr_mux_10__2, d_arr_mux_10__1, 
                    d_arr_mux_10__0, d_arr_mux_11__31, d_arr_mux_11__30, 
                    d_arr_mux_11__29, d_arr_mux_11__28, d_arr_mux_11__27, 
                    d_arr_mux_11__26, d_arr_mux_11__25, d_arr_mux_11__24, 
                    d_arr_mux_11__23, d_arr_mux_11__22, d_arr_mux_11__21, 
                    d_arr_mux_11__20, d_arr_mux_11__19, d_arr_mux_11__18, 
                    d_arr_mux_11__17, d_arr_mux_11__16, d_arr_mux_11__15, 
                    d_arr_mux_11__14, d_arr_mux_11__13, d_arr_mux_11__12, 
                    d_arr_mux_11__11, d_arr_mux_11__10, d_arr_mux_11__9, 
                    d_arr_mux_11__8, d_arr_mux_11__7, d_arr_mux_11__6, 
                    d_arr_mux_11__5, d_arr_mux_11__4, d_arr_mux_11__3, 
                    d_arr_mux_11__2, d_arr_mux_11__1, d_arr_mux_11__0, 
                    d_arr_mux_12__31, d_arr_mux_12__30, d_arr_mux_12__29, 
                    d_arr_mux_12__28, d_arr_mux_12__27, d_arr_mux_12__26, 
                    d_arr_mux_12__25, d_arr_mux_12__24, d_arr_mux_12__23, 
                    d_arr_mux_12__22, d_arr_mux_12__21, d_arr_mux_12__20, 
                    d_arr_mux_12__19, d_arr_mux_12__18, d_arr_mux_12__17, 
                    d_arr_mux_12__16, d_arr_mux_12__15, d_arr_mux_12__14, 
                    d_arr_mux_12__13, d_arr_mux_12__12, d_arr_mux_12__11, 
                    d_arr_mux_12__10, d_arr_mux_12__9, d_arr_mux_12__8, 
                    d_arr_mux_12__7, d_arr_mux_12__6, d_arr_mux_12__5, 
                    d_arr_mux_12__4, d_arr_mux_12__3, d_arr_mux_12__2, 
                    d_arr_mux_12__1, d_arr_mux_12__0, d_arr_mux_13__31, 
                    d_arr_mux_13__30, d_arr_mux_13__29, d_arr_mux_13__28, 
                    d_arr_mux_13__27, d_arr_mux_13__26, d_arr_mux_13__25, 
                    d_arr_mux_13__24, d_arr_mux_13__23, d_arr_mux_13__22, 
                    d_arr_mux_13__21, d_arr_mux_13__20, d_arr_mux_13__19, 
                    d_arr_mux_13__18, d_arr_mux_13__17, d_arr_mux_13__16, 
                    d_arr_mux_13__15, d_arr_mux_13__14, d_arr_mux_13__13, 
                    d_arr_mux_13__12, d_arr_mux_13__11, d_arr_mux_13__10, 
                    d_arr_mux_13__9, d_arr_mux_13__8, d_arr_mux_13__7, 
                    d_arr_mux_13__6, d_arr_mux_13__5, d_arr_mux_13__4, 
                    d_arr_mux_13__3, d_arr_mux_13__2, d_arr_mux_13__1, 
                    d_arr_mux_13__0, d_arr_mux_14__31, d_arr_mux_14__30, 
                    d_arr_mux_14__29, d_arr_mux_14__28, d_arr_mux_14__27, 
                    d_arr_mux_14__26, d_arr_mux_14__25, d_arr_mux_14__24, 
                    d_arr_mux_14__23, d_arr_mux_14__22, d_arr_mux_14__21, 
                    d_arr_mux_14__20, d_arr_mux_14__19, d_arr_mux_14__18, 
                    d_arr_mux_14__17, d_arr_mux_14__16, d_arr_mux_14__15, 
                    d_arr_mux_14__14, d_arr_mux_14__13, d_arr_mux_14__12, 
                    d_arr_mux_14__11, d_arr_mux_14__10, d_arr_mux_14__9, 
                    d_arr_mux_14__8, d_arr_mux_14__7, d_arr_mux_14__6, 
                    d_arr_mux_14__5, d_arr_mux_14__4, d_arr_mux_14__3, 
                    d_arr_mux_14__2, d_arr_mux_14__1, d_arr_mux_14__0, 
                    d_arr_mux_15__31, d_arr_mux_15__30, d_arr_mux_15__29, 
                    d_arr_mux_15__28, d_arr_mux_15__27, d_arr_mux_15__26, 
                    d_arr_mux_15__25, d_arr_mux_15__24, d_arr_mux_15__23, 
                    d_arr_mux_15__22, d_arr_mux_15__21, d_arr_mux_15__20, 
                    d_arr_mux_15__19, d_arr_mux_15__18, d_arr_mux_15__17, 
                    d_arr_mux_15__16, d_arr_mux_15__15, d_arr_mux_15__14, 
                    d_arr_mux_15__13, d_arr_mux_15__12, d_arr_mux_15__11, 
                    d_arr_mux_15__10, d_arr_mux_15__9, d_arr_mux_15__8, 
                    d_arr_mux_15__7, d_arr_mux_15__6, d_arr_mux_15__5, 
                    d_arr_mux_15__4, d_arr_mux_15__3, d_arr_mux_15__2, 
                    d_arr_mux_15__1, d_arr_mux_15__0, d_arr_mux_16__31, 
                    d_arr_mux_16__30, d_arr_mux_16__29, d_arr_mux_16__28, 
                    d_arr_mux_16__27, d_arr_mux_16__26, d_arr_mux_16__25, 
                    d_arr_mux_16__24, d_arr_mux_16__23, d_arr_mux_16__22, 
                    d_arr_mux_16__21, d_arr_mux_16__20, d_arr_mux_16__19, 
                    d_arr_mux_16__18, d_arr_mux_16__17, d_arr_mux_16__16, 
                    d_arr_mux_16__15, d_arr_mux_16__14, d_arr_mux_16__13, 
                    d_arr_mux_16__12, d_arr_mux_16__11, d_arr_mux_16__10, 
                    d_arr_mux_16__9, d_arr_mux_16__8, d_arr_mux_16__7, 
                    d_arr_mux_16__6, d_arr_mux_16__5, d_arr_mux_16__4, 
                    d_arr_mux_16__3, d_arr_mux_16__2, d_arr_mux_16__1, 
                    d_arr_mux_16__0, d_arr_mux_17__31, d_arr_mux_17__30, 
                    d_arr_mux_17__29, d_arr_mux_17__28, d_arr_mux_17__27, 
                    d_arr_mux_17__26, d_arr_mux_17__25, d_arr_mux_17__24, 
                    d_arr_mux_17__23, d_arr_mux_17__22, d_arr_mux_17__21, 
                    d_arr_mux_17__20, d_arr_mux_17__19, d_arr_mux_17__18, 
                    d_arr_mux_17__17, d_arr_mux_17__16, d_arr_mux_17__15, 
                    d_arr_mux_17__14, d_arr_mux_17__13, d_arr_mux_17__12, 
                    d_arr_mux_17__11, d_arr_mux_17__10, d_arr_mux_17__9, 
                    d_arr_mux_17__8, d_arr_mux_17__7, d_arr_mux_17__6, 
                    d_arr_mux_17__5, d_arr_mux_17__4, d_arr_mux_17__3, 
                    d_arr_mux_17__2, d_arr_mux_17__1, d_arr_mux_17__0, 
                    d_arr_mux_18__31, d_arr_mux_18__30, d_arr_mux_18__29, 
                    d_arr_mux_18__28, d_arr_mux_18__27, d_arr_mux_18__26, 
                    d_arr_mux_18__25, d_arr_mux_18__24, d_arr_mux_18__23, 
                    d_arr_mux_18__22, d_arr_mux_18__21, d_arr_mux_18__20, 
                    d_arr_mux_18__19, d_arr_mux_18__18, d_arr_mux_18__17, 
                    d_arr_mux_18__16, d_arr_mux_18__15, d_arr_mux_18__14, 
                    d_arr_mux_18__13, d_arr_mux_18__12, d_arr_mux_18__11, 
                    d_arr_mux_18__10, d_arr_mux_18__9, d_arr_mux_18__8, 
                    d_arr_mux_18__7, d_arr_mux_18__6, d_arr_mux_18__5, 
                    d_arr_mux_18__4, d_arr_mux_18__3, d_arr_mux_18__2, 
                    d_arr_mux_18__1, d_arr_mux_18__0, d_arr_mux_19__31, 
                    d_arr_mux_19__30, d_arr_mux_19__29, d_arr_mux_19__28, 
                    d_arr_mux_19__27, d_arr_mux_19__26, d_arr_mux_19__25, 
                    d_arr_mux_19__24, d_arr_mux_19__23, d_arr_mux_19__22, 
                    d_arr_mux_19__21, d_arr_mux_19__20, d_arr_mux_19__19, 
                    d_arr_mux_19__18, d_arr_mux_19__17, d_arr_mux_19__16, 
                    d_arr_mux_19__15, d_arr_mux_19__14, d_arr_mux_19__13, 
                    d_arr_mux_19__12, d_arr_mux_19__11, d_arr_mux_19__10, 
                    d_arr_mux_19__9, d_arr_mux_19__8, d_arr_mux_19__7, 
                    d_arr_mux_19__6, d_arr_mux_19__5, d_arr_mux_19__4, 
                    d_arr_mux_19__3, d_arr_mux_19__2, d_arr_mux_19__1, 
                    d_arr_mux_19__0, d_arr_mux_20__31, d_arr_mux_20__30, 
                    d_arr_mux_20__29, d_arr_mux_20__28, d_arr_mux_20__27, 
                    d_arr_mux_20__26, d_arr_mux_20__25, d_arr_mux_20__24, 
                    d_arr_mux_20__23, d_arr_mux_20__22, d_arr_mux_20__21, 
                    d_arr_mux_20__20, d_arr_mux_20__19, d_arr_mux_20__18, 
                    d_arr_mux_20__17, d_arr_mux_20__16, d_arr_mux_20__15, 
                    d_arr_mux_20__14, d_arr_mux_20__13, d_arr_mux_20__12, 
                    d_arr_mux_20__11, d_arr_mux_20__10, d_arr_mux_20__9, 
                    d_arr_mux_20__8, d_arr_mux_20__7, d_arr_mux_20__6, 
                    d_arr_mux_20__5, d_arr_mux_20__4, d_arr_mux_20__3, 
                    d_arr_mux_20__2, d_arr_mux_20__1, d_arr_mux_20__0, 
                    d_arr_mux_21__31, d_arr_mux_21__30, d_arr_mux_21__29, 
                    d_arr_mux_21__28, d_arr_mux_21__27, d_arr_mux_21__26, 
                    d_arr_mux_21__25, d_arr_mux_21__24, d_arr_mux_21__23, 
                    d_arr_mux_21__22, d_arr_mux_21__21, d_arr_mux_21__20, 
                    d_arr_mux_21__19, d_arr_mux_21__18, d_arr_mux_21__17, 
                    d_arr_mux_21__16, d_arr_mux_21__15, d_arr_mux_21__14, 
                    d_arr_mux_21__13, d_arr_mux_21__12, d_arr_mux_21__11, 
                    d_arr_mux_21__10, d_arr_mux_21__9, d_arr_mux_21__8, 
                    d_arr_mux_21__7, d_arr_mux_21__6, d_arr_mux_21__5, 
                    d_arr_mux_21__4, d_arr_mux_21__3, d_arr_mux_21__2, 
                    d_arr_mux_21__1, d_arr_mux_21__0, d_arr_mux_22__31, 
                    d_arr_mux_22__30, d_arr_mux_22__29, d_arr_mux_22__28, 
                    d_arr_mux_22__27, d_arr_mux_22__26, d_arr_mux_22__25, 
                    d_arr_mux_22__24, d_arr_mux_22__23, d_arr_mux_22__22, 
                    d_arr_mux_22__21, d_arr_mux_22__20, d_arr_mux_22__19, 
                    d_arr_mux_22__18, d_arr_mux_22__17, d_arr_mux_22__16, 
                    d_arr_mux_22__15, d_arr_mux_22__14, d_arr_mux_22__13, 
                    d_arr_mux_22__12, d_arr_mux_22__11, d_arr_mux_22__10, 
                    d_arr_mux_22__9, d_arr_mux_22__8, d_arr_mux_22__7, 
                    d_arr_mux_22__6, d_arr_mux_22__5, d_arr_mux_22__4, 
                    d_arr_mux_22__3, d_arr_mux_22__2, d_arr_mux_22__1, 
                    d_arr_mux_22__0, d_arr_mux_23__31, d_arr_mux_23__30, 
                    d_arr_mux_23__29, d_arr_mux_23__28, d_arr_mux_23__27, 
                    d_arr_mux_23__26, d_arr_mux_23__25, d_arr_mux_23__24, 
                    d_arr_mux_23__23, d_arr_mux_23__22, d_arr_mux_23__21, 
                    d_arr_mux_23__20, d_arr_mux_23__19, d_arr_mux_23__18, 
                    d_arr_mux_23__17, d_arr_mux_23__16, d_arr_mux_23__15, 
                    d_arr_mux_23__14, d_arr_mux_23__13, d_arr_mux_23__12, 
                    d_arr_mux_23__11, d_arr_mux_23__10, d_arr_mux_23__9, 
                    d_arr_mux_23__8, d_arr_mux_23__7, d_arr_mux_23__6, 
                    d_arr_mux_23__5, d_arr_mux_23__4, d_arr_mux_23__3, 
                    d_arr_mux_23__2, d_arr_mux_23__1, d_arr_mux_23__0, 
                    d_arr_mux_24__31, d_arr_mux_24__30, d_arr_mux_24__29, 
                    d_arr_mux_24__28, d_arr_mux_24__27, d_arr_mux_24__26, 
                    d_arr_mux_24__25, d_arr_mux_24__24, d_arr_mux_24__23, 
                    d_arr_mux_24__22, d_arr_mux_24__21, d_arr_mux_24__20, 
                    d_arr_mux_24__19, d_arr_mux_24__18, d_arr_mux_24__17, 
                    d_arr_mux_24__16, d_arr_mux_24__15, d_arr_mux_24__14, 
                    d_arr_mux_24__13, d_arr_mux_24__12, d_arr_mux_24__11, 
                    d_arr_mux_24__10, d_arr_mux_24__9, d_arr_mux_24__8, 
                    d_arr_mux_24__7, d_arr_mux_24__6, d_arr_mux_24__5, 
                    d_arr_mux_24__4, d_arr_mux_24__3, d_arr_mux_24__2, 
                    d_arr_mux_24__1, d_arr_mux_24__0, d_arr_mul_0__31, 
                    d_arr_mul_0__30, d_arr_mul_0__29, d_arr_mul_0__28, 
                    d_arr_mul_0__27, d_arr_mul_0__26, d_arr_mul_0__25, 
                    d_arr_mul_0__24, d_arr_mul_0__23, d_arr_mul_0__22, 
                    d_arr_mul_0__21, d_arr_mul_0__20, d_arr_mul_0__19, 
                    d_arr_mul_0__18, d_arr_mul_0__17, d_arr_mul_0__16, 
                    d_arr_mul_0__15, d_arr_mul_0__14, d_arr_mul_0__13, 
                    d_arr_mul_0__12, d_arr_mul_0__11, d_arr_mul_0__10, 
                    d_arr_mul_0__9, d_arr_mul_0__8, d_arr_mul_0__7, 
                    d_arr_mul_0__6, d_arr_mul_0__5, d_arr_mul_0__4, 
                    d_arr_mul_0__3, d_arr_mul_0__2, d_arr_mul_0__1, 
                    d_arr_mul_0__0, d_arr_mul_1__31, d_arr_mul_1__30, 
                    d_arr_mul_1__29, d_arr_mul_1__28, d_arr_mul_1__27, 
                    d_arr_mul_1__26, d_arr_mul_1__25, d_arr_mul_1__24, 
                    d_arr_mul_1__23, d_arr_mul_1__22, d_arr_mul_1__21, 
                    d_arr_mul_1__20, d_arr_mul_1__19, d_arr_mul_1__18, 
                    d_arr_mul_1__17, d_arr_mul_1__16, d_arr_mul_1__15, 
                    d_arr_mul_1__14, d_arr_mul_1__13, d_arr_mul_1__12, 
                    d_arr_mul_1__11, d_arr_mul_1__10, d_arr_mul_1__9, 
                    d_arr_mul_1__8, d_arr_mul_1__7, d_arr_mul_1__6, 
                    d_arr_mul_1__5, d_arr_mul_1__4, d_arr_mul_1__3, 
                    d_arr_mul_1__2, d_arr_mul_1__1, d_arr_mul_1__0, 
                    d_arr_mul_2__31, d_arr_mul_2__30, d_arr_mul_2__29, 
                    d_arr_mul_2__28, d_arr_mul_2__27, d_arr_mul_2__26, 
                    d_arr_mul_2__25, d_arr_mul_2__24, d_arr_mul_2__23, 
                    d_arr_mul_2__22, d_arr_mul_2__21, d_arr_mul_2__20, 
                    d_arr_mul_2__19, d_arr_mul_2__18, d_arr_mul_2__17, 
                    d_arr_mul_2__16, d_arr_mul_2__15, d_arr_mul_2__14, 
                    d_arr_mul_2__13, d_arr_mul_2__12, d_arr_mul_2__11, 
                    d_arr_mul_2__10, d_arr_mul_2__9, d_arr_mul_2__8, 
                    d_arr_mul_2__7, d_arr_mul_2__6, d_arr_mul_2__5, 
                    d_arr_mul_2__4, d_arr_mul_2__3, d_arr_mul_2__2, 
                    d_arr_mul_2__1, d_arr_mul_2__0, d_arr_mul_3__31, 
                    d_arr_mul_3__30, d_arr_mul_3__29, d_arr_mul_3__28, 
                    d_arr_mul_3__27, d_arr_mul_3__26, d_arr_mul_3__25, 
                    d_arr_mul_3__24, d_arr_mul_3__23, d_arr_mul_3__22, 
                    d_arr_mul_3__21, d_arr_mul_3__20, d_arr_mul_3__19, 
                    d_arr_mul_3__18, d_arr_mul_3__17, d_arr_mul_3__16, 
                    d_arr_mul_3__15, d_arr_mul_3__14, d_arr_mul_3__13, 
                    d_arr_mul_3__12, d_arr_mul_3__11, d_arr_mul_3__10, 
                    d_arr_mul_3__9, d_arr_mul_3__8, d_arr_mul_3__7, 
                    d_arr_mul_3__6, d_arr_mul_3__5, d_arr_mul_3__4, 
                    d_arr_mul_3__3, d_arr_mul_3__2, d_arr_mul_3__1, 
                    d_arr_mul_3__0, d_arr_mul_4__31, d_arr_mul_4__30, 
                    d_arr_mul_4__29, d_arr_mul_4__28, d_arr_mul_4__27, 
                    d_arr_mul_4__26, d_arr_mul_4__25, d_arr_mul_4__24, 
                    d_arr_mul_4__23, d_arr_mul_4__22, d_arr_mul_4__21, 
                    d_arr_mul_4__20, d_arr_mul_4__19, d_arr_mul_4__18, 
                    d_arr_mul_4__17, d_arr_mul_4__16, d_arr_mul_4__15, 
                    d_arr_mul_4__14, d_arr_mul_4__13, d_arr_mul_4__12, 
                    d_arr_mul_4__11, d_arr_mul_4__10, d_arr_mul_4__9, 
                    d_arr_mul_4__8, d_arr_mul_4__7, d_arr_mul_4__6, 
                    d_arr_mul_4__5, d_arr_mul_4__4, d_arr_mul_4__3, 
                    d_arr_mul_4__2, d_arr_mul_4__1, d_arr_mul_4__0, 
                    d_arr_mul_5__31, d_arr_mul_5__30, d_arr_mul_5__29, 
                    d_arr_mul_5__28, d_arr_mul_5__27, d_arr_mul_5__26, 
                    d_arr_mul_5__25, d_arr_mul_5__24, d_arr_mul_5__23, 
                    d_arr_mul_5__22, d_arr_mul_5__21, d_arr_mul_5__20, 
                    d_arr_mul_5__19, d_arr_mul_5__18, d_arr_mul_5__17, 
                    d_arr_mul_5__16, d_arr_mul_5__15, d_arr_mul_5__14, 
                    d_arr_mul_5__13, d_arr_mul_5__12, d_arr_mul_5__11, 
                    d_arr_mul_5__10, d_arr_mul_5__9, d_arr_mul_5__8, 
                    d_arr_mul_5__7, d_arr_mul_5__6, d_arr_mul_5__5, 
                    d_arr_mul_5__4, d_arr_mul_5__3, d_arr_mul_5__2, 
                    d_arr_mul_5__1, d_arr_mul_5__0, d_arr_mul_6__31, 
                    d_arr_mul_6__30, d_arr_mul_6__29, d_arr_mul_6__28, 
                    d_arr_mul_6__27, d_arr_mul_6__26, d_arr_mul_6__25, 
                    d_arr_mul_6__24, d_arr_mul_6__23, d_arr_mul_6__22, 
                    d_arr_mul_6__21, d_arr_mul_6__20, d_arr_mul_6__19, 
                    d_arr_mul_6__18, d_arr_mul_6__17, d_arr_mul_6__16, 
                    d_arr_mul_6__15, d_arr_mul_6__14, d_arr_mul_6__13, 
                    d_arr_mul_6__12, d_arr_mul_6__11, d_arr_mul_6__10, 
                    d_arr_mul_6__9, d_arr_mul_6__8, d_arr_mul_6__7, 
                    d_arr_mul_6__6, d_arr_mul_6__5, d_arr_mul_6__4, 
                    d_arr_mul_6__3, d_arr_mul_6__2, d_arr_mul_6__1, 
                    d_arr_mul_6__0, d_arr_mul_7__31, d_arr_mul_7__30, 
                    d_arr_mul_7__29, d_arr_mul_7__28, d_arr_mul_7__27, 
                    d_arr_mul_7__26, d_arr_mul_7__25, d_arr_mul_7__24, 
                    d_arr_mul_7__23, d_arr_mul_7__22, d_arr_mul_7__21, 
                    d_arr_mul_7__20, d_arr_mul_7__19, d_arr_mul_7__18, 
                    d_arr_mul_7__17, d_arr_mul_7__16, d_arr_mul_7__15, 
                    d_arr_mul_7__14, d_arr_mul_7__13, d_arr_mul_7__12, 
                    d_arr_mul_7__11, d_arr_mul_7__10, d_arr_mul_7__9, 
                    d_arr_mul_7__8, d_arr_mul_7__7, d_arr_mul_7__6, 
                    d_arr_mul_7__5, d_arr_mul_7__4, d_arr_mul_7__3, 
                    d_arr_mul_7__2, d_arr_mul_7__1, d_arr_mul_7__0, 
                    d_arr_mul_8__31, d_arr_mul_8__30, d_arr_mul_8__29, 
                    d_arr_mul_8__28, d_arr_mul_8__27, d_arr_mul_8__26, 
                    d_arr_mul_8__25, d_arr_mul_8__24, d_arr_mul_8__23, 
                    d_arr_mul_8__22, d_arr_mul_8__21, d_arr_mul_8__20, 
                    d_arr_mul_8__19, d_arr_mul_8__18, d_arr_mul_8__17, 
                    d_arr_mul_8__16, d_arr_mul_8__15, d_arr_mul_8__14, 
                    d_arr_mul_8__13, d_arr_mul_8__12, d_arr_mul_8__11, 
                    d_arr_mul_8__10, d_arr_mul_8__9, d_arr_mul_8__8, 
                    d_arr_mul_8__7, d_arr_mul_8__6, d_arr_mul_8__5, 
                    d_arr_mul_8__4, d_arr_mul_8__3, d_arr_mul_8__2, 
                    d_arr_mul_8__1, d_arr_mul_8__0, d_arr_mul_9__31, 
                    d_arr_mul_9__30, d_arr_mul_9__29, d_arr_mul_9__28, 
                    d_arr_mul_9__27, d_arr_mul_9__26, d_arr_mul_9__25, 
                    d_arr_mul_9__24, d_arr_mul_9__23, d_arr_mul_9__22, 
                    d_arr_mul_9__21, d_arr_mul_9__20, d_arr_mul_9__19, 
                    d_arr_mul_9__18, d_arr_mul_9__17, d_arr_mul_9__16, 
                    d_arr_mul_9__15, d_arr_mul_9__14, d_arr_mul_9__13, 
                    d_arr_mul_9__12, d_arr_mul_9__11, d_arr_mul_9__10, 
                    d_arr_mul_9__9, d_arr_mul_9__8, d_arr_mul_9__7, 
                    d_arr_mul_9__6, d_arr_mul_9__5, d_arr_mul_9__4, 
                    d_arr_mul_9__3, d_arr_mul_9__2, d_arr_mul_9__1, 
                    d_arr_mul_9__0, d_arr_mul_10__31, d_arr_mul_10__30, 
                    d_arr_mul_10__29, d_arr_mul_10__28, d_arr_mul_10__27, 
                    d_arr_mul_10__26, d_arr_mul_10__25, d_arr_mul_10__24, 
                    d_arr_mul_10__23, d_arr_mul_10__22, d_arr_mul_10__21, 
                    d_arr_mul_10__20, d_arr_mul_10__19, d_arr_mul_10__18, 
                    d_arr_mul_10__17, d_arr_mul_10__16, d_arr_mul_10__15, 
                    d_arr_mul_10__14, d_arr_mul_10__13, d_arr_mul_10__12, 
                    d_arr_mul_10__11, d_arr_mul_10__10, d_arr_mul_10__9, 
                    d_arr_mul_10__8, d_arr_mul_10__7, d_arr_mul_10__6, 
                    d_arr_mul_10__5, d_arr_mul_10__4, d_arr_mul_10__3, 
                    d_arr_mul_10__2, d_arr_mul_10__1, d_arr_mul_10__0, 
                    d_arr_mul_11__31, d_arr_mul_11__30, d_arr_mul_11__29, 
                    d_arr_mul_11__28, d_arr_mul_11__27, d_arr_mul_11__26, 
                    d_arr_mul_11__25, d_arr_mul_11__24, d_arr_mul_11__23, 
                    d_arr_mul_11__22, d_arr_mul_11__21, d_arr_mul_11__20, 
                    d_arr_mul_11__19, d_arr_mul_11__18, d_arr_mul_11__17, 
                    d_arr_mul_11__16, d_arr_mul_11__15, d_arr_mul_11__14, 
                    d_arr_mul_11__13, d_arr_mul_11__12, d_arr_mul_11__11, 
                    d_arr_mul_11__10, d_arr_mul_11__9, d_arr_mul_11__8, 
                    d_arr_mul_11__7, d_arr_mul_11__6, d_arr_mul_11__5, 
                    d_arr_mul_11__4, d_arr_mul_11__3, d_arr_mul_11__2, 
                    d_arr_mul_11__1, d_arr_mul_11__0, d_arr_mul_12__31, 
                    d_arr_mul_12__30, d_arr_mul_12__29, d_arr_mul_12__28, 
                    d_arr_mul_12__27, d_arr_mul_12__26, d_arr_mul_12__25, 
                    d_arr_mul_12__24, d_arr_mul_12__23, d_arr_mul_12__22, 
                    d_arr_mul_12__21, d_arr_mul_12__20, d_arr_mul_12__19, 
                    d_arr_mul_12__18, d_arr_mul_12__17, d_arr_mul_12__16, 
                    d_arr_mul_12__15, d_arr_mul_12__14, d_arr_mul_12__13, 
                    d_arr_mul_12__12, d_arr_mul_12__11, d_arr_mul_12__10, 
                    d_arr_mul_12__9, d_arr_mul_12__8, d_arr_mul_12__7, 
                    d_arr_mul_12__6, d_arr_mul_12__5, d_arr_mul_12__4, 
                    d_arr_mul_12__3, d_arr_mul_12__2, d_arr_mul_12__1, 
                    d_arr_mul_12__0, d_arr_mul_13__31, d_arr_mul_13__30, 
                    d_arr_mul_13__29, d_arr_mul_13__28, d_arr_mul_13__27, 
                    d_arr_mul_13__26, d_arr_mul_13__25, d_arr_mul_13__24, 
                    d_arr_mul_13__23, d_arr_mul_13__22, d_arr_mul_13__21, 
                    d_arr_mul_13__20, d_arr_mul_13__19, d_arr_mul_13__18, 
                    d_arr_mul_13__17, d_arr_mul_13__16, d_arr_mul_13__15, 
                    d_arr_mul_13__14, d_arr_mul_13__13, d_arr_mul_13__12, 
                    d_arr_mul_13__11, d_arr_mul_13__10, d_arr_mul_13__9, 
                    d_arr_mul_13__8, d_arr_mul_13__7, d_arr_mul_13__6, 
                    d_arr_mul_13__5, d_arr_mul_13__4, d_arr_mul_13__3, 
                    d_arr_mul_13__2, d_arr_mul_13__1, d_arr_mul_13__0, 
                    d_arr_mul_14__31, d_arr_mul_14__30, d_arr_mul_14__29, 
                    d_arr_mul_14__28, d_arr_mul_14__27, d_arr_mul_14__26, 
                    d_arr_mul_14__25, d_arr_mul_14__24, d_arr_mul_14__23, 
                    d_arr_mul_14__22, d_arr_mul_14__21, d_arr_mul_14__20, 
                    d_arr_mul_14__19, d_arr_mul_14__18, d_arr_mul_14__17, 
                    d_arr_mul_14__16, d_arr_mul_14__15, d_arr_mul_14__14, 
                    d_arr_mul_14__13, d_arr_mul_14__12, d_arr_mul_14__11, 
                    d_arr_mul_14__10, d_arr_mul_14__9, d_arr_mul_14__8, 
                    d_arr_mul_14__7, d_arr_mul_14__6, d_arr_mul_14__5, 
                    d_arr_mul_14__4, d_arr_mul_14__3, d_arr_mul_14__2, 
                    d_arr_mul_14__1, d_arr_mul_14__0, d_arr_mul_15__31, 
                    d_arr_mul_15__30, d_arr_mul_15__29, d_arr_mul_15__28, 
                    d_arr_mul_15__27, d_arr_mul_15__26, d_arr_mul_15__25, 
                    d_arr_mul_15__24, d_arr_mul_15__23, d_arr_mul_15__22, 
                    d_arr_mul_15__21, d_arr_mul_15__20, d_arr_mul_15__19, 
                    d_arr_mul_15__18, d_arr_mul_15__17, d_arr_mul_15__16, 
                    d_arr_mul_15__15, d_arr_mul_15__14, d_arr_mul_15__13, 
                    d_arr_mul_15__12, d_arr_mul_15__11, d_arr_mul_15__10, 
                    d_arr_mul_15__9, d_arr_mul_15__8, d_arr_mul_15__7, 
                    d_arr_mul_15__6, d_arr_mul_15__5, d_arr_mul_15__4, 
                    d_arr_mul_15__3, d_arr_mul_15__2, d_arr_mul_15__1, 
                    d_arr_mul_15__0, d_arr_mul_16__31, d_arr_mul_16__30, 
                    d_arr_mul_16__29, d_arr_mul_16__28, d_arr_mul_16__27, 
                    d_arr_mul_16__26, d_arr_mul_16__25, d_arr_mul_16__24, 
                    d_arr_mul_16__23, d_arr_mul_16__22, d_arr_mul_16__21, 
                    d_arr_mul_16__20, d_arr_mul_16__19, d_arr_mul_16__18, 
                    d_arr_mul_16__17, d_arr_mul_16__16, d_arr_mul_16__15, 
                    d_arr_mul_16__14, d_arr_mul_16__13, d_arr_mul_16__12, 
                    d_arr_mul_16__11, d_arr_mul_16__10, d_arr_mul_16__9, 
                    d_arr_mul_16__8, d_arr_mul_16__7, d_arr_mul_16__6, 
                    d_arr_mul_16__5, d_arr_mul_16__4, d_arr_mul_16__3, 
                    d_arr_mul_16__2, d_arr_mul_16__1, d_arr_mul_16__0, 
                    d_arr_mul_17__31, d_arr_mul_17__30, d_arr_mul_17__29, 
                    d_arr_mul_17__28, d_arr_mul_17__27, d_arr_mul_17__26, 
                    d_arr_mul_17__25, d_arr_mul_17__24, d_arr_mul_17__23, 
                    d_arr_mul_17__22, d_arr_mul_17__21, d_arr_mul_17__20, 
                    d_arr_mul_17__19, d_arr_mul_17__18, d_arr_mul_17__17, 
                    d_arr_mul_17__16, d_arr_mul_17__15, d_arr_mul_17__14, 
                    d_arr_mul_17__13, d_arr_mul_17__12, d_arr_mul_17__11, 
                    d_arr_mul_17__10, d_arr_mul_17__9, d_arr_mul_17__8, 
                    d_arr_mul_17__7, d_arr_mul_17__6, d_arr_mul_17__5, 
                    d_arr_mul_17__4, d_arr_mul_17__3, d_arr_mul_17__2, 
                    d_arr_mul_17__1, d_arr_mul_17__0, d_arr_mul_18__31, 
                    d_arr_mul_18__30, d_arr_mul_18__29, d_arr_mul_18__28, 
                    d_arr_mul_18__27, d_arr_mul_18__26, d_arr_mul_18__25, 
                    d_arr_mul_18__24, d_arr_mul_18__23, d_arr_mul_18__22, 
                    d_arr_mul_18__21, d_arr_mul_18__20, d_arr_mul_18__19, 
                    d_arr_mul_18__18, d_arr_mul_18__17, d_arr_mul_18__16, 
                    d_arr_mul_18__15, d_arr_mul_18__14, d_arr_mul_18__13, 
                    d_arr_mul_18__12, d_arr_mul_18__11, d_arr_mul_18__10, 
                    d_arr_mul_18__9, d_arr_mul_18__8, d_arr_mul_18__7, 
                    d_arr_mul_18__6, d_arr_mul_18__5, d_arr_mul_18__4, 
                    d_arr_mul_18__3, d_arr_mul_18__2, d_arr_mul_18__1, 
                    d_arr_mul_18__0, d_arr_mul_19__31, d_arr_mul_19__30, 
                    d_arr_mul_19__29, d_arr_mul_19__28, d_arr_mul_19__27, 
                    d_arr_mul_19__26, d_arr_mul_19__25, d_arr_mul_19__24, 
                    d_arr_mul_19__23, d_arr_mul_19__22, d_arr_mul_19__21, 
                    d_arr_mul_19__20, d_arr_mul_19__19, d_arr_mul_19__18, 
                    d_arr_mul_19__17, d_arr_mul_19__16, d_arr_mul_19__15, 
                    d_arr_mul_19__14, d_arr_mul_19__13, d_arr_mul_19__12, 
                    d_arr_mul_19__11, d_arr_mul_19__10, d_arr_mul_19__9, 
                    d_arr_mul_19__8, d_arr_mul_19__7, d_arr_mul_19__6, 
                    d_arr_mul_19__5, d_arr_mul_19__4, d_arr_mul_19__3, 
                    d_arr_mul_19__2, d_arr_mul_19__1, d_arr_mul_19__0, 
                    d_arr_mul_20__31, d_arr_mul_20__30, d_arr_mul_20__29, 
                    d_arr_mul_20__28, d_arr_mul_20__27, d_arr_mul_20__26, 
                    d_arr_mul_20__25, d_arr_mul_20__24, d_arr_mul_20__23, 
                    d_arr_mul_20__22, d_arr_mul_20__21, d_arr_mul_20__20, 
                    d_arr_mul_20__19, d_arr_mul_20__18, d_arr_mul_20__17, 
                    d_arr_mul_20__16, d_arr_mul_20__15, d_arr_mul_20__14, 
                    d_arr_mul_20__13, d_arr_mul_20__12, d_arr_mul_20__11, 
                    d_arr_mul_20__10, d_arr_mul_20__9, d_arr_mul_20__8, 
                    d_arr_mul_20__7, d_arr_mul_20__6, d_arr_mul_20__5, 
                    d_arr_mul_20__4, d_arr_mul_20__3, d_arr_mul_20__2, 
                    d_arr_mul_20__1, d_arr_mul_20__0, d_arr_mul_21__31, 
                    d_arr_mul_21__30, d_arr_mul_21__29, d_arr_mul_21__28, 
                    d_arr_mul_21__27, d_arr_mul_21__26, d_arr_mul_21__25, 
                    d_arr_mul_21__24, d_arr_mul_21__23, d_arr_mul_21__22, 
                    d_arr_mul_21__21, d_arr_mul_21__20, d_arr_mul_21__19, 
                    d_arr_mul_21__18, d_arr_mul_21__17, d_arr_mul_21__16, 
                    d_arr_mul_21__15, d_arr_mul_21__14, d_arr_mul_21__13, 
                    d_arr_mul_21__12, d_arr_mul_21__11, d_arr_mul_21__10, 
                    d_arr_mul_21__9, d_arr_mul_21__8, d_arr_mul_21__7, 
                    d_arr_mul_21__6, d_arr_mul_21__5, d_arr_mul_21__4, 
                    d_arr_mul_21__3, d_arr_mul_21__2, d_arr_mul_21__1, 
                    d_arr_mul_21__0, d_arr_mul_22__31, d_arr_mul_22__30, 
                    d_arr_mul_22__29, d_arr_mul_22__28, d_arr_mul_22__27, 
                    d_arr_mul_22__26, d_arr_mul_22__25, d_arr_mul_22__24, 
                    d_arr_mul_22__23, d_arr_mul_22__22, d_arr_mul_22__21, 
                    d_arr_mul_22__20, d_arr_mul_22__19, d_arr_mul_22__18, 
                    d_arr_mul_22__17, d_arr_mul_22__16, d_arr_mul_22__15, 
                    d_arr_mul_22__14, d_arr_mul_22__13, d_arr_mul_22__12, 
                    d_arr_mul_22__11, d_arr_mul_22__10, d_arr_mul_22__9, 
                    d_arr_mul_22__8, d_arr_mul_22__7, d_arr_mul_22__6, 
                    d_arr_mul_22__5, d_arr_mul_22__4, d_arr_mul_22__3, 
                    d_arr_mul_22__2, d_arr_mul_22__1, d_arr_mul_22__0, 
                    d_arr_mul_23__31, d_arr_mul_23__30, d_arr_mul_23__29, 
                    d_arr_mul_23__28, d_arr_mul_23__27, d_arr_mul_23__26, 
                    d_arr_mul_23__25, d_arr_mul_23__24, d_arr_mul_23__23, 
                    d_arr_mul_23__22, d_arr_mul_23__21, d_arr_mul_23__20, 
                    d_arr_mul_23__19, d_arr_mul_23__18, d_arr_mul_23__17, 
                    d_arr_mul_23__16, d_arr_mul_23__15, d_arr_mul_23__14, 
                    d_arr_mul_23__13, d_arr_mul_23__12, d_arr_mul_23__11, 
                    d_arr_mul_23__10, d_arr_mul_23__9, d_arr_mul_23__8, 
                    d_arr_mul_23__7, d_arr_mul_23__6, d_arr_mul_23__5, 
                    d_arr_mul_23__4, d_arr_mul_23__3, d_arr_mul_23__2, 
                    d_arr_mul_23__1, d_arr_mul_23__0, d_arr_mul_24__31, 
                    d_arr_mul_24__30, d_arr_mul_24__29, d_arr_mul_24__28, 
                    d_arr_mul_24__27, d_arr_mul_24__26, d_arr_mul_24__25, 
                    d_arr_mul_24__24, d_arr_mul_24__23, d_arr_mul_24__22, 
                    d_arr_mul_24__21, d_arr_mul_24__20, d_arr_mul_24__19, 
                    d_arr_mul_24__18, d_arr_mul_24__17, d_arr_mul_24__16, 
                    d_arr_mul_24__15, d_arr_mul_24__14, d_arr_mul_24__13, 
                    d_arr_mul_24__12, d_arr_mul_24__11, d_arr_mul_24__10, 
                    d_arr_mul_24__9, d_arr_mul_24__8, d_arr_mul_24__7, 
                    d_arr_mul_24__6, d_arr_mul_24__5, d_arr_mul_24__4, 
                    d_arr_mul_24__3, d_arr_mul_24__2, d_arr_mul_24__1, 
                    d_arr_mul_24__0, d_arr_add_0__31, d_arr_add_0__30, 
                    d_arr_add_0__29, d_arr_add_0__28, d_arr_add_0__27, 
                    d_arr_add_0__26, d_arr_add_0__25, d_arr_add_0__24, 
                    d_arr_add_0__23, d_arr_add_0__22, d_arr_add_0__21, 
                    d_arr_add_0__20, d_arr_add_0__19, d_arr_add_0__18, 
                    d_arr_add_0__17, d_arr_add_0__16, d_arr_add_0__15, 
                    d_arr_add_0__14, d_arr_add_0__13, d_arr_add_0__12, 
                    d_arr_add_0__11, d_arr_add_0__10, d_arr_add_0__9, 
                    d_arr_add_0__8, d_arr_add_0__7, d_arr_add_0__6, 
                    d_arr_add_0__5, d_arr_add_0__4, d_arr_add_0__3, 
                    d_arr_add_0__2, d_arr_add_0__1, d_arr_add_0__0, 
                    d_arr_add_1__31, d_arr_add_1__30, d_arr_add_1__29, 
                    d_arr_add_1__28, d_arr_add_1__27, d_arr_add_1__26, 
                    d_arr_add_1__25, d_arr_add_1__24, d_arr_add_1__23, 
                    d_arr_add_1__22, d_arr_add_1__21, d_arr_add_1__20, 
                    d_arr_add_1__19, d_arr_add_1__18, d_arr_add_1__17, 
                    d_arr_add_1__16, d_arr_add_1__15, d_arr_add_1__14, 
                    d_arr_add_1__13, d_arr_add_1__12, d_arr_add_1__11, 
                    d_arr_add_1__10, d_arr_add_1__9, d_arr_add_1__8, 
                    d_arr_add_1__7, d_arr_add_1__6, d_arr_add_1__5, 
                    d_arr_add_1__4, d_arr_add_1__3, d_arr_add_1__2, 
                    d_arr_add_1__1, d_arr_add_1__0, d_arr_add_2__31, 
                    d_arr_add_2__30, d_arr_add_2__29, d_arr_add_2__28, 
                    d_arr_add_2__27, d_arr_add_2__26, d_arr_add_2__25, 
                    d_arr_add_2__24, d_arr_add_2__23, d_arr_add_2__22, 
                    d_arr_add_2__21, d_arr_add_2__20, d_arr_add_2__19, 
                    d_arr_add_2__18, d_arr_add_2__17, d_arr_add_2__16, 
                    d_arr_add_2__15, d_arr_add_2__14, d_arr_add_2__13, 
                    d_arr_add_2__12, d_arr_add_2__11, d_arr_add_2__10, 
                    d_arr_add_2__9, d_arr_add_2__8, d_arr_add_2__7, 
                    d_arr_add_2__6, d_arr_add_2__5, d_arr_add_2__4, 
                    d_arr_add_2__3, d_arr_add_2__2, d_arr_add_2__1, 
                    d_arr_add_2__0, d_arr_add_3__31, d_arr_add_3__30, 
                    d_arr_add_3__29, d_arr_add_3__28, d_arr_add_3__27, 
                    d_arr_add_3__26, d_arr_add_3__25, d_arr_add_3__24, 
                    d_arr_add_3__23, d_arr_add_3__22, d_arr_add_3__21, 
                    d_arr_add_3__20, d_arr_add_3__19, d_arr_add_3__18, 
                    d_arr_add_3__17, d_arr_add_3__16, d_arr_add_3__15, 
                    d_arr_add_3__14, d_arr_add_3__13, d_arr_add_3__12, 
                    d_arr_add_3__11, d_arr_add_3__10, d_arr_add_3__9, 
                    d_arr_add_3__8, d_arr_add_3__7, d_arr_add_3__6, 
                    d_arr_add_3__5, d_arr_add_3__4, d_arr_add_3__3, 
                    d_arr_add_3__2, d_arr_add_3__1, d_arr_add_3__0, 
                    d_arr_add_4__31, d_arr_add_4__30, d_arr_add_4__29, 
                    d_arr_add_4__28, d_arr_add_4__27, d_arr_add_4__26, 
                    d_arr_add_4__25, d_arr_add_4__24, d_arr_add_4__23, 
                    d_arr_add_4__22, d_arr_add_4__21, d_arr_add_4__20, 
                    d_arr_add_4__19, d_arr_add_4__18, d_arr_add_4__17, 
                    d_arr_add_4__16, d_arr_add_4__15, d_arr_add_4__14, 
                    d_arr_add_4__13, d_arr_add_4__12, d_arr_add_4__11, 
                    d_arr_add_4__10, d_arr_add_4__9, d_arr_add_4__8, 
                    d_arr_add_4__7, d_arr_add_4__6, d_arr_add_4__5, 
                    d_arr_add_4__4, d_arr_add_4__3, d_arr_add_4__2, 
                    d_arr_add_4__1, d_arr_add_4__0, d_arr_add_5__31, 
                    d_arr_add_5__30, d_arr_add_5__29, d_arr_add_5__28, 
                    d_arr_add_5__27, d_arr_add_5__26, d_arr_add_5__25, 
                    d_arr_add_5__24, d_arr_add_5__23, d_arr_add_5__22, 
                    d_arr_add_5__21, d_arr_add_5__20, d_arr_add_5__19, 
                    d_arr_add_5__18, d_arr_add_5__17, d_arr_add_5__16, 
                    d_arr_add_5__15, d_arr_add_5__14, d_arr_add_5__13, 
                    d_arr_add_5__12, d_arr_add_5__11, d_arr_add_5__10, 
                    d_arr_add_5__9, d_arr_add_5__8, d_arr_add_5__7, 
                    d_arr_add_5__6, d_arr_add_5__5, d_arr_add_5__4, 
                    d_arr_add_5__3, d_arr_add_5__2, d_arr_add_5__1, 
                    d_arr_add_5__0, d_arr_add_6__31, d_arr_add_6__30, 
                    d_arr_add_6__29, d_arr_add_6__28, d_arr_add_6__27, 
                    d_arr_add_6__26, d_arr_add_6__25, d_arr_add_6__24, 
                    d_arr_add_6__23, d_arr_add_6__22, d_arr_add_6__21, 
                    d_arr_add_6__20, d_arr_add_6__19, d_arr_add_6__18, 
                    d_arr_add_6__17, d_arr_add_6__16, d_arr_add_6__15, 
                    d_arr_add_6__14, d_arr_add_6__13, d_arr_add_6__12, 
                    d_arr_add_6__11, d_arr_add_6__10, d_arr_add_6__9, 
                    d_arr_add_6__8, d_arr_add_6__7, d_arr_add_6__6, 
                    d_arr_add_6__5, d_arr_add_6__4, d_arr_add_6__3, 
                    d_arr_add_6__2, d_arr_add_6__1, d_arr_add_6__0, 
                    d_arr_add_7__31, d_arr_add_7__30, d_arr_add_7__29, 
                    d_arr_add_7__28, d_arr_add_7__27, d_arr_add_7__26, 
                    d_arr_add_7__25, d_arr_add_7__24, d_arr_add_7__23, 
                    d_arr_add_7__22, d_arr_add_7__21, d_arr_add_7__20, 
                    d_arr_add_7__19, d_arr_add_7__18, d_arr_add_7__17, 
                    d_arr_add_7__16, d_arr_add_7__15, d_arr_add_7__14, 
                    d_arr_add_7__13, d_arr_add_7__12, d_arr_add_7__11, 
                    d_arr_add_7__10, d_arr_add_7__9, d_arr_add_7__8, 
                    d_arr_add_7__7, d_arr_add_7__6, d_arr_add_7__5, 
                    d_arr_add_7__4, d_arr_add_7__3, d_arr_add_7__2, 
                    d_arr_add_7__1, d_arr_add_7__0, d_arr_add_8__31, 
                    d_arr_add_8__30, d_arr_add_8__29, d_arr_add_8__28, 
                    d_arr_add_8__27, d_arr_add_8__26, d_arr_add_8__25, 
                    d_arr_add_8__24, d_arr_add_8__23, d_arr_add_8__22, 
                    d_arr_add_8__21, d_arr_add_8__20, d_arr_add_8__19, 
                    d_arr_add_8__18, d_arr_add_8__17, d_arr_add_8__16, 
                    d_arr_add_8__15, d_arr_add_8__14, d_arr_add_8__13, 
                    d_arr_add_8__12, d_arr_add_8__11, d_arr_add_8__10, 
                    d_arr_add_8__9, d_arr_add_8__8, d_arr_add_8__7, 
                    d_arr_add_8__6, d_arr_add_8__5, d_arr_add_8__4, 
                    d_arr_add_8__3, d_arr_add_8__2, d_arr_add_8__1, 
                    d_arr_add_8__0, d_arr_add_9__31, d_arr_add_9__30, 
                    d_arr_add_9__29, d_arr_add_9__28, d_arr_add_9__27, 
                    d_arr_add_9__26, d_arr_add_9__25, d_arr_add_9__24, 
                    d_arr_add_9__23, d_arr_add_9__22, d_arr_add_9__21, 
                    d_arr_add_9__20, d_arr_add_9__19, d_arr_add_9__18, 
                    d_arr_add_9__17, d_arr_add_9__16, d_arr_add_9__15, 
                    d_arr_add_9__14, d_arr_add_9__13, d_arr_add_9__12, 
                    d_arr_add_9__11, d_arr_add_9__10, d_arr_add_9__9, 
                    d_arr_add_9__8, d_arr_add_9__7, d_arr_add_9__6, 
                    d_arr_add_9__5, d_arr_add_9__4, d_arr_add_9__3, 
                    d_arr_add_9__2, d_arr_add_9__1, d_arr_add_9__0, 
                    d_arr_add_10__31, d_arr_add_10__30, d_arr_add_10__29, 
                    d_arr_add_10__28, d_arr_add_10__27, d_arr_add_10__26, 
                    d_arr_add_10__25, d_arr_add_10__24, d_arr_add_10__23, 
                    d_arr_add_10__22, d_arr_add_10__21, d_arr_add_10__20, 
                    d_arr_add_10__19, d_arr_add_10__18, d_arr_add_10__17, 
                    d_arr_add_10__16, d_arr_add_10__15, d_arr_add_10__14, 
                    d_arr_add_10__13, d_arr_add_10__12, d_arr_add_10__11, 
                    d_arr_add_10__10, d_arr_add_10__9, d_arr_add_10__8, 
                    d_arr_add_10__7, d_arr_add_10__6, d_arr_add_10__5, 
                    d_arr_add_10__4, d_arr_add_10__3, d_arr_add_10__2, 
                    d_arr_add_10__1, d_arr_add_10__0, d_arr_add_11__31, 
                    d_arr_add_11__30, d_arr_add_11__29, d_arr_add_11__28, 
                    d_arr_add_11__27, d_arr_add_11__26, d_arr_add_11__25, 
                    d_arr_add_11__24, d_arr_add_11__23, d_arr_add_11__22, 
                    d_arr_add_11__21, d_arr_add_11__20, d_arr_add_11__19, 
                    d_arr_add_11__18, d_arr_add_11__17, d_arr_add_11__16, 
                    d_arr_add_11__15, d_arr_add_11__14, d_arr_add_11__13, 
                    d_arr_add_11__12, d_arr_add_11__11, d_arr_add_11__10, 
                    d_arr_add_11__9, d_arr_add_11__8, d_arr_add_11__7, 
                    d_arr_add_11__6, d_arr_add_11__5, d_arr_add_11__4, 
                    d_arr_add_11__3, d_arr_add_11__2, d_arr_add_11__1, 
                    d_arr_add_11__0, d_arr_add_12__31, d_arr_add_12__30, 
                    d_arr_add_12__29, d_arr_add_12__28, d_arr_add_12__27, 
                    d_arr_add_12__26, d_arr_add_12__25, d_arr_add_12__24, 
                    d_arr_add_12__23, d_arr_add_12__22, d_arr_add_12__21, 
                    d_arr_add_12__20, d_arr_add_12__19, d_arr_add_12__18, 
                    d_arr_add_12__17, d_arr_add_12__16, d_arr_add_12__15, 
                    d_arr_add_12__14, d_arr_add_12__13, d_arr_add_12__12, 
                    d_arr_add_12__11, d_arr_add_12__10, d_arr_add_12__9, 
                    d_arr_add_12__8, d_arr_add_12__7, d_arr_add_12__6, 
                    d_arr_add_12__5, d_arr_add_12__4, d_arr_add_12__3, 
                    d_arr_add_12__2, d_arr_add_12__1, d_arr_add_12__0, 
                    d_arr_add_13__31, d_arr_add_13__30, d_arr_add_13__29, 
                    d_arr_add_13__28, d_arr_add_13__27, d_arr_add_13__26, 
                    d_arr_add_13__25, d_arr_add_13__24, d_arr_add_13__23, 
                    d_arr_add_13__22, d_arr_add_13__21, d_arr_add_13__20, 
                    d_arr_add_13__19, d_arr_add_13__18, d_arr_add_13__17, 
                    d_arr_add_13__16, d_arr_add_13__15, d_arr_add_13__14, 
                    d_arr_add_13__13, d_arr_add_13__12, d_arr_add_13__11, 
                    d_arr_add_13__10, d_arr_add_13__9, d_arr_add_13__8, 
                    d_arr_add_13__7, d_arr_add_13__6, d_arr_add_13__5, 
                    d_arr_add_13__4, d_arr_add_13__3, d_arr_add_13__2, 
                    d_arr_add_13__1, d_arr_add_13__0, d_arr_add_14__31, 
                    d_arr_add_14__30, d_arr_add_14__29, d_arr_add_14__28, 
                    d_arr_add_14__27, d_arr_add_14__26, d_arr_add_14__25, 
                    d_arr_add_14__24, d_arr_add_14__23, d_arr_add_14__22, 
                    d_arr_add_14__21, d_arr_add_14__20, d_arr_add_14__19, 
                    d_arr_add_14__18, d_arr_add_14__17, d_arr_add_14__16, 
                    d_arr_add_14__15, d_arr_add_14__14, d_arr_add_14__13, 
                    d_arr_add_14__12, d_arr_add_14__11, d_arr_add_14__10, 
                    d_arr_add_14__9, d_arr_add_14__8, d_arr_add_14__7, 
                    d_arr_add_14__6, d_arr_add_14__5, d_arr_add_14__4, 
                    d_arr_add_14__3, d_arr_add_14__2, d_arr_add_14__1, 
                    d_arr_add_14__0, d_arr_add_15__31, d_arr_add_15__30, 
                    d_arr_add_15__29, d_arr_add_15__28, d_arr_add_15__27, 
                    d_arr_add_15__26, d_arr_add_15__25, d_arr_add_15__24, 
                    d_arr_add_15__23, d_arr_add_15__22, d_arr_add_15__21, 
                    d_arr_add_15__20, d_arr_add_15__19, d_arr_add_15__18, 
                    d_arr_add_15__17, d_arr_add_15__16, d_arr_add_15__15, 
                    d_arr_add_15__14, d_arr_add_15__13, d_arr_add_15__12, 
                    d_arr_add_15__11, d_arr_add_15__10, d_arr_add_15__9, 
                    d_arr_add_15__8, d_arr_add_15__7, d_arr_add_15__6, 
                    d_arr_add_15__5, d_arr_add_15__4, d_arr_add_15__3, 
                    d_arr_add_15__2, d_arr_add_15__1, d_arr_add_15__0, 
                    d_arr_add_16__31, d_arr_add_16__30, d_arr_add_16__29, 
                    d_arr_add_16__28, d_arr_add_16__27, d_arr_add_16__26, 
                    d_arr_add_16__25, d_arr_add_16__24, d_arr_add_16__23, 
                    d_arr_add_16__22, d_arr_add_16__21, d_arr_add_16__20, 
                    d_arr_add_16__19, d_arr_add_16__18, d_arr_add_16__17, 
                    d_arr_add_16__16, d_arr_add_16__15, d_arr_add_16__14, 
                    d_arr_add_16__13, d_arr_add_16__12, d_arr_add_16__11, 
                    d_arr_add_16__10, d_arr_add_16__9, d_arr_add_16__8, 
                    d_arr_add_16__7, d_arr_add_16__6, d_arr_add_16__5, 
                    d_arr_add_16__4, d_arr_add_16__3, d_arr_add_16__2, 
                    d_arr_add_16__1, d_arr_add_16__0, d_arr_add_17__31, 
                    d_arr_add_17__30, d_arr_add_17__29, d_arr_add_17__28, 
                    d_arr_add_17__27, d_arr_add_17__26, d_arr_add_17__25, 
                    d_arr_add_17__24, d_arr_add_17__23, d_arr_add_17__22, 
                    d_arr_add_17__21, d_arr_add_17__20, d_arr_add_17__19, 
                    d_arr_add_17__18, d_arr_add_17__17, d_arr_add_17__16, 
                    d_arr_add_17__15, d_arr_add_17__14, d_arr_add_17__13, 
                    d_arr_add_17__12, d_arr_add_17__11, d_arr_add_17__10, 
                    d_arr_add_17__9, d_arr_add_17__8, d_arr_add_17__7, 
                    d_arr_add_17__6, d_arr_add_17__5, d_arr_add_17__4, 
                    d_arr_add_17__3, d_arr_add_17__2, d_arr_add_17__1, 
                    d_arr_add_17__0, d_arr_add_18__31, d_arr_add_18__30, 
                    d_arr_add_18__29, d_arr_add_18__28, d_arr_add_18__27, 
                    d_arr_add_18__26, d_arr_add_18__25, d_arr_add_18__24, 
                    d_arr_add_18__23, d_arr_add_18__22, d_arr_add_18__21, 
                    d_arr_add_18__20, d_arr_add_18__19, d_arr_add_18__18, 
                    d_arr_add_18__17, d_arr_add_18__16, d_arr_add_18__15, 
                    d_arr_add_18__14, d_arr_add_18__13, d_arr_add_18__12, 
                    d_arr_add_18__11, d_arr_add_18__10, d_arr_add_18__9, 
                    d_arr_add_18__8, d_arr_add_18__7, d_arr_add_18__6, 
                    d_arr_add_18__5, d_arr_add_18__4, d_arr_add_18__3, 
                    d_arr_add_18__2, d_arr_add_18__1, d_arr_add_18__0, 
                    d_arr_add_19__31, d_arr_add_19__30, d_arr_add_19__29, 
                    d_arr_add_19__28, d_arr_add_19__27, d_arr_add_19__26, 
                    d_arr_add_19__25, d_arr_add_19__24, d_arr_add_19__23, 
                    d_arr_add_19__22, d_arr_add_19__21, d_arr_add_19__20, 
                    d_arr_add_19__19, d_arr_add_19__18, d_arr_add_19__17, 
                    d_arr_add_19__16, d_arr_add_19__15, d_arr_add_19__14, 
                    d_arr_add_19__13, d_arr_add_19__12, d_arr_add_19__11, 
                    d_arr_add_19__10, d_arr_add_19__9, d_arr_add_19__8, 
                    d_arr_add_19__7, d_arr_add_19__6, d_arr_add_19__5, 
                    d_arr_add_19__4, d_arr_add_19__3, d_arr_add_19__2, 
                    d_arr_add_19__1, d_arr_add_19__0, d_arr_add_20__31, 
                    d_arr_add_20__30, d_arr_add_20__29, d_arr_add_20__28, 
                    d_arr_add_20__27, d_arr_add_20__26, d_arr_add_20__25, 
                    d_arr_add_20__24, d_arr_add_20__23, d_arr_add_20__22, 
                    d_arr_add_20__21, d_arr_add_20__20, d_arr_add_20__19, 
                    d_arr_add_20__18, d_arr_add_20__17, d_arr_add_20__16, 
                    d_arr_add_20__15, d_arr_add_20__14, d_arr_add_20__13, 
                    d_arr_add_20__12, d_arr_add_20__11, d_arr_add_20__10, 
                    d_arr_add_20__9, d_arr_add_20__8, d_arr_add_20__7, 
                    d_arr_add_20__6, d_arr_add_20__5, d_arr_add_20__4, 
                    d_arr_add_20__3, d_arr_add_20__2, d_arr_add_20__1, 
                    d_arr_add_20__0, d_arr_add_21__31, d_arr_add_21__30, 
                    d_arr_add_21__29, d_arr_add_21__28, d_arr_add_21__27, 
                    d_arr_add_21__26, d_arr_add_21__25, d_arr_add_21__24, 
                    d_arr_add_21__23, d_arr_add_21__22, d_arr_add_21__21, 
                    d_arr_add_21__20, d_arr_add_21__19, d_arr_add_21__18, 
                    d_arr_add_21__17, d_arr_add_21__16, d_arr_add_21__15, 
                    d_arr_add_21__14, d_arr_add_21__13, d_arr_add_21__12, 
                    d_arr_add_21__11, d_arr_add_21__10, d_arr_add_21__9, 
                    d_arr_add_21__8, d_arr_add_21__7, d_arr_add_21__6, 
                    d_arr_add_21__5, d_arr_add_21__4, d_arr_add_21__3, 
                    d_arr_add_21__2, d_arr_add_21__1, d_arr_add_21__0, 
                    d_arr_add_22__31, d_arr_add_22__30, d_arr_add_22__29, 
                    d_arr_add_22__28, d_arr_add_22__27, d_arr_add_22__26, 
                    d_arr_add_22__25, d_arr_add_22__24, d_arr_add_22__23, 
                    d_arr_add_22__22, d_arr_add_22__21, d_arr_add_22__20, 
                    d_arr_add_22__19, d_arr_add_22__18, d_arr_add_22__17, 
                    d_arr_add_22__16, d_arr_add_22__15, d_arr_add_22__14, 
                    d_arr_add_22__13, d_arr_add_22__12, d_arr_add_22__11, 
                    d_arr_add_22__10, d_arr_add_22__9, d_arr_add_22__8, 
                    d_arr_add_22__7, d_arr_add_22__6, d_arr_add_22__5, 
                    d_arr_add_22__4, d_arr_add_22__3, d_arr_add_22__2, 
                    d_arr_add_22__1, d_arr_add_22__0, d_arr_add_23__31, 
                    d_arr_add_23__30, d_arr_add_23__29, d_arr_add_23__28, 
                    d_arr_add_23__27, d_arr_add_23__26, d_arr_add_23__25, 
                    d_arr_add_23__24, d_arr_add_23__23, d_arr_add_23__22, 
                    d_arr_add_23__21, d_arr_add_23__20, d_arr_add_23__19, 
                    d_arr_add_23__18, d_arr_add_23__17, d_arr_add_23__16, 
                    d_arr_add_23__15, d_arr_add_23__14, d_arr_add_23__13, 
                    d_arr_add_23__12, d_arr_add_23__11, d_arr_add_23__10, 
                    d_arr_add_23__9, d_arr_add_23__8, d_arr_add_23__7, 
                    d_arr_add_23__6, d_arr_add_23__5, d_arr_add_23__4, 
                    d_arr_add_23__3, d_arr_add_23__2, d_arr_add_23__1, 
                    d_arr_add_23__0, d_arr_add_24__31, d_arr_add_24__30, 
                    d_arr_add_24__29, d_arr_add_24__28, d_arr_add_24__27, 
                    d_arr_add_24__26, d_arr_add_24__25, d_arr_add_24__24, 
                    d_arr_add_24__23, d_arr_add_24__22, d_arr_add_24__21, 
                    d_arr_add_24__20, d_arr_add_24__19, d_arr_add_24__18, 
                    d_arr_add_24__17, d_arr_add_24__16, d_arr_add_24__15, 
                    d_arr_add_24__14, d_arr_add_24__13, d_arr_add_24__12, 
                    d_arr_add_24__11, d_arr_add_24__10, d_arr_add_24__9, 
                    d_arr_add_24__8, d_arr_add_24__7, d_arr_add_24__6, 
                    d_arr_add_24__5, d_arr_add_24__4, d_arr_add_24__3, 
                    d_arr_add_24__2, d_arr_add_24__1, d_arr_add_24__0, 
                    d_arr_merge1_0__31, d_arr_merge1_0__30, d_arr_merge1_0__29, 
                    d_arr_merge1_0__28, d_arr_merge1_0__27, d_arr_merge1_0__26, 
                    d_arr_merge1_0__25, d_arr_merge1_0__24, d_arr_merge1_0__23, 
                    d_arr_merge1_0__22, d_arr_merge1_0__21, d_arr_merge1_0__20, 
                    d_arr_merge1_0__19, d_arr_merge1_0__18, d_arr_merge1_0__17, 
                    d_arr_merge1_0__16, d_arr_merge1_0__15, d_arr_merge1_0__14, 
                    d_arr_merge1_0__13, d_arr_merge1_0__12, d_arr_merge1_0__11, 
                    d_arr_merge1_0__10, d_arr_merge1_0__9, d_arr_merge1_0__8, 
                    d_arr_merge1_0__7, d_arr_merge1_0__6, d_arr_merge1_0__5, 
                    d_arr_merge1_0__4, d_arr_merge1_0__3, d_arr_merge1_0__2, 
                    d_arr_merge1_0__1, d_arr_merge1_0__0, d_arr_merge1_1__31, 
                    d_arr_merge1_1__30, d_arr_merge1_1__29, d_arr_merge1_1__28, 
                    d_arr_merge1_1__27, d_arr_merge1_1__26, d_arr_merge1_1__25, 
                    d_arr_merge1_1__24, d_arr_merge1_1__23, d_arr_merge1_1__22, 
                    d_arr_merge1_1__21, d_arr_merge1_1__20, d_arr_merge1_1__19, 
                    d_arr_merge1_1__18, d_arr_merge1_1__17, d_arr_merge1_1__16, 
                    d_arr_merge1_1__15, d_arr_merge1_1__14, d_arr_merge1_1__13, 
                    d_arr_merge1_1__12, d_arr_merge1_1__11, d_arr_merge1_1__10, 
                    d_arr_merge1_1__9, d_arr_merge1_1__8, d_arr_merge1_1__7, 
                    d_arr_merge1_1__6, d_arr_merge1_1__5, d_arr_merge1_1__4, 
                    d_arr_merge1_1__3, d_arr_merge1_1__2, d_arr_merge1_1__1, 
                    d_arr_merge1_1__0, d_arr_merge1_2__31, d_arr_merge1_2__30, 
                    d_arr_merge1_2__29, d_arr_merge1_2__28, d_arr_merge1_2__27, 
                    d_arr_merge1_2__26, d_arr_merge1_2__25, d_arr_merge1_2__24, 
                    d_arr_merge1_2__23, d_arr_merge1_2__22, d_arr_merge1_2__21, 
                    d_arr_merge1_2__20, d_arr_merge1_2__19, d_arr_merge1_2__18, 
                    d_arr_merge1_2__17, d_arr_merge1_2__16, d_arr_merge1_2__15, 
                    d_arr_merge1_2__14, d_arr_merge1_2__13, d_arr_merge1_2__12, 
                    d_arr_merge1_2__11, d_arr_merge1_2__10, d_arr_merge1_2__9, 
                    d_arr_merge1_2__8, d_arr_merge1_2__7, d_arr_merge1_2__6, 
                    d_arr_merge1_2__5, d_arr_merge1_2__4, d_arr_merge1_2__3, 
                    d_arr_merge1_2__2, d_arr_merge1_2__1, d_arr_merge1_2__0, 
                    d_arr_merge1_3__31, d_arr_merge1_3__30, d_arr_merge1_3__29, 
                    d_arr_merge1_3__28, d_arr_merge1_3__27, d_arr_merge1_3__26, 
                    d_arr_merge1_3__25, d_arr_merge1_3__24, d_arr_merge1_3__23, 
                    d_arr_merge1_3__22, d_arr_merge1_3__21, d_arr_merge1_3__20, 
                    d_arr_merge1_3__19, d_arr_merge1_3__18, d_arr_merge1_3__17, 
                    d_arr_merge1_3__16, d_arr_merge1_3__15, d_arr_merge1_3__14, 
                    d_arr_merge1_3__13, d_arr_merge1_3__12, d_arr_merge1_3__11, 
                    d_arr_merge1_3__10, d_arr_merge1_3__9, d_arr_merge1_3__8, 
                    d_arr_merge1_3__7, d_arr_merge1_3__6, d_arr_merge1_3__5, 
                    d_arr_merge1_3__4, d_arr_merge1_3__3, d_arr_merge1_3__2, 
                    d_arr_merge1_3__1, d_arr_merge1_3__0, d_arr_merge1_4__31, 
                    d_arr_merge1_4__30, d_arr_merge1_4__29, d_arr_merge1_4__28, 
                    d_arr_merge1_4__27, d_arr_merge1_4__26, d_arr_merge1_4__25, 
                    d_arr_merge1_4__24, d_arr_merge1_4__23, d_arr_merge1_4__22, 
                    d_arr_merge1_4__21, d_arr_merge1_4__20, d_arr_merge1_4__19, 
                    d_arr_merge1_4__18, d_arr_merge1_4__17, d_arr_merge1_4__16, 
                    d_arr_merge1_4__15, d_arr_merge1_4__14, d_arr_merge1_4__13, 
                    d_arr_merge1_4__12, d_arr_merge1_4__11, d_arr_merge1_4__10, 
                    d_arr_merge1_4__9, d_arr_merge1_4__8, d_arr_merge1_4__7, 
                    d_arr_merge1_4__6, d_arr_merge1_4__5, d_arr_merge1_4__4, 
                    d_arr_merge1_4__3, d_arr_merge1_4__2, d_arr_merge1_4__1, 
                    d_arr_merge1_4__0, d_arr_merge1_5__31, d_arr_merge1_5__30, 
                    d_arr_merge1_5__29, d_arr_merge1_5__28, d_arr_merge1_5__27, 
                    d_arr_merge1_5__26, d_arr_merge1_5__25, d_arr_merge1_5__24, 
                    d_arr_merge1_5__23, d_arr_merge1_5__22, d_arr_merge1_5__21, 
                    d_arr_merge1_5__20, d_arr_merge1_5__19, d_arr_merge1_5__18, 
                    d_arr_merge1_5__17, d_arr_merge1_5__16, d_arr_merge1_5__15, 
                    d_arr_merge1_5__14, d_arr_merge1_5__13, d_arr_merge1_5__12, 
                    d_arr_merge1_5__11, d_arr_merge1_5__10, d_arr_merge1_5__9, 
                    d_arr_merge1_5__8, d_arr_merge1_5__7, d_arr_merge1_5__6, 
                    d_arr_merge1_5__5, d_arr_merge1_5__4, d_arr_merge1_5__3, 
                    d_arr_merge1_5__2, d_arr_merge1_5__1, d_arr_merge1_5__0, 
                    d_arr_merge1_6__31, d_arr_merge1_6__30, d_arr_merge1_6__29, 
                    d_arr_merge1_6__28, d_arr_merge1_6__27, d_arr_merge1_6__26, 
                    d_arr_merge1_6__25, d_arr_merge1_6__24, d_arr_merge1_6__23, 
                    d_arr_merge1_6__22, d_arr_merge1_6__21, d_arr_merge1_6__20, 
                    d_arr_merge1_6__19, d_arr_merge1_6__18, d_arr_merge1_6__17, 
                    d_arr_merge1_6__16, d_arr_merge1_6__15, d_arr_merge1_6__14, 
                    d_arr_merge1_6__13, d_arr_merge1_6__12, d_arr_merge1_6__11, 
                    d_arr_merge1_6__10, d_arr_merge1_6__9, d_arr_merge1_6__8, 
                    d_arr_merge1_6__7, d_arr_merge1_6__6, d_arr_merge1_6__5, 
                    d_arr_merge1_6__4, d_arr_merge1_6__3, d_arr_merge1_6__2, 
                    d_arr_merge1_6__1, d_arr_merge1_6__0, d_arr_merge1_7__31, 
                    d_arr_merge1_7__30, d_arr_merge1_7__29, d_arr_merge1_7__28, 
                    d_arr_merge1_7__27, d_arr_merge1_7__26, d_arr_merge1_7__25, 
                    d_arr_merge1_7__24, d_arr_merge1_7__23, d_arr_merge1_7__22, 
                    d_arr_merge1_7__21, d_arr_merge1_7__20, d_arr_merge1_7__19, 
                    d_arr_merge1_7__18, d_arr_merge1_7__17, d_arr_merge1_7__16, 
                    d_arr_merge1_7__15, d_arr_merge1_7__14, d_arr_merge1_7__13, 
                    d_arr_merge1_7__12, d_arr_merge1_7__11, d_arr_merge1_7__10, 
                    d_arr_merge1_7__9, d_arr_merge1_7__8, d_arr_merge1_7__7, 
                    d_arr_merge1_7__6, d_arr_merge1_7__5, d_arr_merge1_7__4, 
                    d_arr_merge1_7__3, d_arr_merge1_7__2, d_arr_merge1_7__1, 
                    d_arr_merge1_7__0, d_arr_merge1_8__31, d_arr_merge1_8__30, 
                    d_arr_merge1_8__29, d_arr_merge1_8__28, d_arr_merge1_8__27, 
                    d_arr_merge1_8__26, d_arr_merge1_8__25, d_arr_merge1_8__24, 
                    d_arr_merge1_8__23, d_arr_merge1_8__22, d_arr_merge1_8__21, 
                    d_arr_merge1_8__20, d_arr_merge1_8__19, d_arr_merge1_8__18, 
                    d_arr_merge1_8__17, d_arr_merge1_8__16, d_arr_merge1_8__15, 
                    d_arr_merge1_8__14, d_arr_merge1_8__13, d_arr_merge1_8__12, 
                    d_arr_merge1_8__11, d_arr_merge1_8__10, d_arr_merge1_8__9, 
                    d_arr_merge1_8__8, d_arr_merge1_8__7, d_arr_merge1_8__6, 
                    d_arr_merge1_8__5, d_arr_merge1_8__4, d_arr_merge1_8__3, 
                    d_arr_merge1_8__2, d_arr_merge1_8__1, d_arr_merge1_8__0, 
                    d_arr_merge1_9__31, d_arr_merge1_9__30, d_arr_merge1_9__29, 
                    d_arr_merge1_9__28, d_arr_merge1_9__27, d_arr_merge1_9__26, 
                    d_arr_merge1_9__25, d_arr_merge1_9__24, d_arr_merge1_9__23, 
                    d_arr_merge1_9__22, d_arr_merge1_9__21, d_arr_merge1_9__20, 
                    d_arr_merge1_9__19, d_arr_merge1_9__18, d_arr_merge1_9__17, 
                    d_arr_merge1_9__16, d_arr_merge1_9__15, d_arr_merge1_9__14, 
                    d_arr_merge1_9__13, d_arr_merge1_9__12, d_arr_merge1_9__11, 
                    d_arr_merge1_9__10, d_arr_merge1_9__9, d_arr_merge1_9__8, 
                    d_arr_merge1_9__7, d_arr_merge1_9__6, d_arr_merge1_9__5, 
                    d_arr_merge1_9__4, d_arr_merge1_9__3, d_arr_merge1_9__2, 
                    d_arr_merge1_9__1, d_arr_merge1_9__0, d_arr_merge1_10__31, 
                    d_arr_merge1_10__30, d_arr_merge1_10__29, 
                    d_arr_merge1_10__28, d_arr_merge1_10__27, 
                    d_arr_merge1_10__26, d_arr_merge1_10__25, 
                    d_arr_merge1_10__24, d_arr_merge1_10__23, 
                    d_arr_merge1_10__22, d_arr_merge1_10__21, 
                    d_arr_merge1_10__20, d_arr_merge1_10__19, 
                    d_arr_merge1_10__18, d_arr_merge1_10__17, 
                    d_arr_merge1_10__16, d_arr_merge1_10__15, 
                    d_arr_merge1_10__14, d_arr_merge1_10__13, 
                    d_arr_merge1_10__12, d_arr_merge1_10__11, 
                    d_arr_merge1_10__10, d_arr_merge1_10__9, d_arr_merge1_10__8, 
                    d_arr_merge1_10__7, d_arr_merge1_10__6, d_arr_merge1_10__5, 
                    d_arr_merge1_10__4, d_arr_merge1_10__3, d_arr_merge1_10__2, 
                    d_arr_merge1_10__1, d_arr_merge1_10__0, d_arr_merge1_11__31, 
                    d_arr_merge1_11__30, d_arr_merge1_11__29, 
                    d_arr_merge1_11__28, d_arr_merge1_11__27, 
                    d_arr_merge1_11__26, d_arr_merge1_11__25, 
                    d_arr_merge1_11__24, d_arr_merge1_11__23, 
                    d_arr_merge1_11__22, d_arr_merge1_11__21, 
                    d_arr_merge1_11__20, d_arr_merge1_11__19, 
                    d_arr_merge1_11__18, d_arr_merge1_11__17, 
                    d_arr_merge1_11__16, d_arr_merge1_11__15, 
                    d_arr_merge1_11__14, d_arr_merge1_11__13, 
                    d_arr_merge1_11__12, d_arr_merge1_11__11, 
                    d_arr_merge1_11__10, d_arr_merge1_11__9, d_arr_merge1_11__8, 
                    d_arr_merge1_11__7, d_arr_merge1_11__6, d_arr_merge1_11__5, 
                    d_arr_merge1_11__4, d_arr_merge1_11__3, d_arr_merge1_11__2, 
                    d_arr_merge1_11__1, d_arr_merge1_11__0, d_arr_merge1_12__31, 
                    d_arr_merge1_12__30, d_arr_merge1_12__29, 
                    d_arr_merge1_12__28, d_arr_merge1_12__27, 
                    d_arr_merge1_12__26, d_arr_merge1_12__25, 
                    d_arr_merge1_12__24, d_arr_merge1_12__23, 
                    d_arr_merge1_12__22, d_arr_merge1_12__21, 
                    d_arr_merge1_12__20, d_arr_merge1_12__19, 
                    d_arr_merge1_12__18, d_arr_merge1_12__17, 
                    d_arr_merge1_12__16, d_arr_merge1_12__15, 
                    d_arr_merge1_12__14, d_arr_merge1_12__13, 
                    d_arr_merge1_12__12, d_arr_merge1_12__11, 
                    d_arr_merge1_12__10, d_arr_merge1_12__9, d_arr_merge1_12__8, 
                    d_arr_merge1_12__7, d_arr_merge1_12__6, d_arr_merge1_12__5, 
                    d_arr_merge1_12__4, d_arr_merge1_12__3, d_arr_merge1_12__2, 
                    d_arr_merge1_12__1, d_arr_merge1_12__0, d_arr_merge1_13__31, 
                    d_arr_merge1_13__30, d_arr_merge1_13__29, 
                    d_arr_merge1_13__28, d_arr_merge1_13__27, 
                    d_arr_merge1_13__26, d_arr_merge1_13__25, 
                    d_arr_merge1_13__24, d_arr_merge1_13__23, 
                    d_arr_merge1_13__22, d_arr_merge1_13__21, 
                    d_arr_merge1_13__20, d_arr_merge1_13__19, 
                    d_arr_merge1_13__18, d_arr_merge1_13__17, 
                    d_arr_merge1_13__16, d_arr_merge1_13__15, 
                    d_arr_merge1_13__14, d_arr_merge1_13__13, 
                    d_arr_merge1_13__12, d_arr_merge1_13__11, 
                    d_arr_merge1_13__10, d_arr_merge1_13__9, d_arr_merge1_13__8, 
                    d_arr_merge1_13__7, d_arr_merge1_13__6, d_arr_merge1_13__5, 
                    d_arr_merge1_13__4, d_arr_merge1_13__3, d_arr_merge1_13__2, 
                    d_arr_merge1_13__1, d_arr_merge1_13__0, d_arr_merge1_14__31, 
                    d_arr_merge1_14__30, d_arr_merge1_14__29, 
                    d_arr_merge1_14__28, d_arr_merge1_14__27, 
                    d_arr_merge1_14__26, d_arr_merge1_14__25, 
                    d_arr_merge1_14__24, d_arr_merge1_14__23, 
                    d_arr_merge1_14__22, d_arr_merge1_14__21, 
                    d_arr_merge1_14__20, d_arr_merge1_14__19, 
                    d_arr_merge1_14__18, d_arr_merge1_14__17, 
                    d_arr_merge1_14__16, d_arr_merge1_14__15, 
                    d_arr_merge1_14__14, d_arr_merge1_14__13, 
                    d_arr_merge1_14__12, d_arr_merge1_14__11, 
                    d_arr_merge1_14__10, d_arr_merge1_14__9, d_arr_merge1_14__8, 
                    d_arr_merge1_14__7, d_arr_merge1_14__6, d_arr_merge1_14__5, 
                    d_arr_merge1_14__4, d_arr_merge1_14__3, d_arr_merge1_14__2, 
                    d_arr_merge1_14__1, d_arr_merge1_14__0, d_arr_merge1_15__31, 
                    d_arr_merge1_15__30, d_arr_merge1_15__29, 
                    d_arr_merge1_15__28, d_arr_merge1_15__27, 
                    d_arr_merge1_15__26, d_arr_merge1_15__25, 
                    d_arr_merge1_15__24, d_arr_merge1_15__23, 
                    d_arr_merge1_15__22, d_arr_merge1_15__21, 
                    d_arr_merge1_15__20, d_arr_merge1_15__19, 
                    d_arr_merge1_15__18, d_arr_merge1_15__17, 
                    d_arr_merge1_15__16, d_arr_merge1_15__15, 
                    d_arr_merge1_15__14, d_arr_merge1_15__13, 
                    d_arr_merge1_15__12, d_arr_merge1_15__11, 
                    d_arr_merge1_15__10, d_arr_merge1_15__9, d_arr_merge1_15__8, 
                    d_arr_merge1_15__7, d_arr_merge1_15__6, d_arr_merge1_15__5, 
                    d_arr_merge1_15__4, d_arr_merge1_15__3, d_arr_merge1_15__2, 
                    d_arr_merge1_15__1, d_arr_merge1_15__0, d_arr_merge1_16__31, 
                    d_arr_merge1_16__30, d_arr_merge1_16__29, 
                    d_arr_merge1_16__28, d_arr_merge1_16__27, 
                    d_arr_merge1_16__26, d_arr_merge1_16__25, 
                    d_arr_merge1_16__24, d_arr_merge1_16__23, 
                    d_arr_merge1_16__22, d_arr_merge1_16__21, 
                    d_arr_merge1_16__20, d_arr_merge1_16__19, 
                    d_arr_merge1_16__18, d_arr_merge1_16__17, 
                    d_arr_merge1_16__16, d_arr_merge1_16__15, 
                    d_arr_merge1_16__14, d_arr_merge1_16__13, 
                    d_arr_merge1_16__12, d_arr_merge1_16__11, 
                    d_arr_merge1_16__10, d_arr_merge1_16__9, d_arr_merge1_16__8, 
                    d_arr_merge1_16__7, d_arr_merge1_16__6, d_arr_merge1_16__5, 
                    d_arr_merge1_16__4, d_arr_merge1_16__3, d_arr_merge1_16__2, 
                    d_arr_merge1_16__1, d_arr_merge1_16__0, d_arr_merge1_17__31, 
                    d_arr_merge1_17__30, d_arr_merge1_17__29, 
                    d_arr_merge1_17__28, d_arr_merge1_17__27, 
                    d_arr_merge1_17__26, d_arr_merge1_17__25, 
                    d_arr_merge1_17__24, d_arr_merge1_17__23, 
                    d_arr_merge1_17__22, d_arr_merge1_17__21, 
                    d_arr_merge1_17__20, d_arr_merge1_17__19, 
                    d_arr_merge1_17__18, d_arr_merge1_17__17, 
                    d_arr_merge1_17__16, d_arr_merge1_17__15, 
                    d_arr_merge1_17__14, d_arr_merge1_17__13, 
                    d_arr_merge1_17__12, d_arr_merge1_17__11, 
                    d_arr_merge1_17__10, d_arr_merge1_17__9, d_arr_merge1_17__8, 
                    d_arr_merge1_17__7, d_arr_merge1_17__6, d_arr_merge1_17__5, 
                    d_arr_merge1_17__4, d_arr_merge1_17__3, d_arr_merge1_17__2, 
                    d_arr_merge1_17__1, d_arr_merge1_17__0, d_arr_merge1_18__31, 
                    d_arr_merge1_18__30, d_arr_merge1_18__29, 
                    d_arr_merge1_18__28, d_arr_merge1_18__27, 
                    d_arr_merge1_18__26, d_arr_merge1_18__25, 
                    d_arr_merge1_18__24, d_arr_merge1_18__23, 
                    d_arr_merge1_18__22, d_arr_merge1_18__21, 
                    d_arr_merge1_18__20, d_arr_merge1_18__19, 
                    d_arr_merge1_18__18, d_arr_merge1_18__17, 
                    d_arr_merge1_18__16, d_arr_merge1_18__15, 
                    d_arr_merge1_18__14, d_arr_merge1_18__13, 
                    d_arr_merge1_18__12, d_arr_merge1_18__11, 
                    d_arr_merge1_18__10, d_arr_merge1_18__9, d_arr_merge1_18__8, 
                    d_arr_merge1_18__7, d_arr_merge1_18__6, d_arr_merge1_18__5, 
                    d_arr_merge1_18__4, d_arr_merge1_18__3, d_arr_merge1_18__2, 
                    d_arr_merge1_18__1, d_arr_merge1_18__0, d_arr_merge1_19__31, 
                    d_arr_merge1_19__30, d_arr_merge1_19__29, 
                    d_arr_merge1_19__28, d_arr_merge1_19__27, 
                    d_arr_merge1_19__26, d_arr_merge1_19__25, 
                    d_arr_merge1_19__24, d_arr_merge1_19__23, 
                    d_arr_merge1_19__22, d_arr_merge1_19__21, 
                    d_arr_merge1_19__20, d_arr_merge1_19__19, 
                    d_arr_merge1_19__18, d_arr_merge1_19__17, 
                    d_arr_merge1_19__16, d_arr_merge1_19__15, 
                    d_arr_merge1_19__14, d_arr_merge1_19__13, 
                    d_arr_merge1_19__12, d_arr_merge1_19__11, 
                    d_arr_merge1_19__10, d_arr_merge1_19__9, d_arr_merge1_19__8, 
                    d_arr_merge1_19__7, d_arr_merge1_19__6, d_arr_merge1_19__5, 
                    d_arr_merge1_19__4, d_arr_merge1_19__3, d_arr_merge1_19__2, 
                    d_arr_merge1_19__1, d_arr_merge1_19__0, d_arr_merge1_20__31, 
                    d_arr_merge1_20__30, d_arr_merge1_20__29, 
                    d_arr_merge1_20__28, d_arr_merge1_20__27, 
                    d_arr_merge1_20__26, d_arr_merge1_20__25, 
                    d_arr_merge1_20__24, d_arr_merge1_20__23, 
                    d_arr_merge1_20__22, d_arr_merge1_20__21, 
                    d_arr_merge1_20__20, d_arr_merge1_20__19, 
                    d_arr_merge1_20__18, d_arr_merge1_20__17, 
                    d_arr_merge1_20__16, d_arr_merge1_20__15, 
                    d_arr_merge1_20__14, d_arr_merge1_20__13, 
                    d_arr_merge1_20__12, d_arr_merge1_20__11, 
                    d_arr_merge1_20__10, d_arr_merge1_20__9, d_arr_merge1_20__8, 
                    d_arr_merge1_20__7, d_arr_merge1_20__6, d_arr_merge1_20__5, 
                    d_arr_merge1_20__4, d_arr_merge1_20__3, d_arr_merge1_20__2, 
                    d_arr_merge1_20__1, d_arr_merge1_20__0, d_arr_merge1_21__31, 
                    d_arr_merge1_21__30, d_arr_merge1_21__29, 
                    d_arr_merge1_21__28, d_arr_merge1_21__27, 
                    d_arr_merge1_21__26, d_arr_merge1_21__25, 
                    d_arr_merge1_21__24, d_arr_merge1_21__23, 
                    d_arr_merge1_21__22, d_arr_merge1_21__21, 
                    d_arr_merge1_21__20, d_arr_merge1_21__19, 
                    d_arr_merge1_21__18, d_arr_merge1_21__17, 
                    d_arr_merge1_21__16, d_arr_merge1_21__15, 
                    d_arr_merge1_21__14, d_arr_merge1_21__13, 
                    d_arr_merge1_21__12, d_arr_merge1_21__11, 
                    d_arr_merge1_21__10, d_arr_merge1_21__9, d_arr_merge1_21__8, 
                    d_arr_merge1_21__7, d_arr_merge1_21__6, d_arr_merge1_21__5, 
                    d_arr_merge1_21__4, d_arr_merge1_21__3, d_arr_merge1_21__2, 
                    d_arr_merge1_21__1, d_arr_merge1_21__0, d_arr_merge1_22__31, 
                    d_arr_merge1_22__30, d_arr_merge1_22__29, 
                    d_arr_merge1_22__28, d_arr_merge1_22__27, 
                    d_arr_merge1_22__26, d_arr_merge1_22__25, 
                    d_arr_merge1_22__24, d_arr_merge1_22__23, 
                    d_arr_merge1_22__22, d_arr_merge1_22__21, 
                    d_arr_merge1_22__20, d_arr_merge1_22__19, 
                    d_arr_merge1_22__18, d_arr_merge1_22__17, 
                    d_arr_merge1_22__16, d_arr_merge1_22__15, 
                    d_arr_merge1_22__14, d_arr_merge1_22__13, 
                    d_arr_merge1_22__12, d_arr_merge1_22__11, 
                    d_arr_merge1_22__10, d_arr_merge1_22__9, d_arr_merge1_22__8, 
                    d_arr_merge1_22__7, d_arr_merge1_22__6, d_arr_merge1_22__5, 
                    d_arr_merge1_22__4, d_arr_merge1_22__3, d_arr_merge1_22__2, 
                    d_arr_merge1_22__1, d_arr_merge1_22__0, d_arr_merge1_23__31, 
                    d_arr_merge1_23__30, d_arr_merge1_23__29, 
                    d_arr_merge1_23__28, d_arr_merge1_23__27, 
                    d_arr_merge1_23__26, d_arr_merge1_23__25, 
                    d_arr_merge1_23__24, d_arr_merge1_23__23, 
                    d_arr_merge1_23__22, d_arr_merge1_23__21, 
                    d_arr_merge1_23__20, d_arr_merge1_23__19, 
                    d_arr_merge1_23__18, d_arr_merge1_23__17, 
                    d_arr_merge1_23__16, d_arr_merge1_23__15, 
                    d_arr_merge1_23__14, d_arr_merge1_23__13, 
                    d_arr_merge1_23__12, d_arr_merge1_23__11, 
                    d_arr_merge1_23__10, d_arr_merge1_23__9, d_arr_merge1_23__8, 
                    d_arr_merge1_23__7, d_arr_merge1_23__6, d_arr_merge1_23__5, 
                    d_arr_merge1_23__4, d_arr_merge1_23__3, d_arr_merge1_23__2, 
                    d_arr_merge1_23__1, d_arr_merge1_23__0, d_arr_merge1_24__31, 
                    d_arr_merge1_24__30, d_arr_merge1_24__29, 
                    d_arr_merge1_24__28, d_arr_merge1_24__27, 
                    d_arr_merge1_24__26, d_arr_merge1_24__25, 
                    d_arr_merge1_24__24, d_arr_merge1_24__23, 
                    d_arr_merge1_24__22, d_arr_merge1_24__21, 
                    d_arr_merge1_24__20, d_arr_merge1_24__19, 
                    d_arr_merge1_24__18, d_arr_merge1_24__17, 
                    d_arr_merge1_24__16, d_arr_merge1_24__15, 
                    d_arr_merge1_24__14, d_arr_merge1_24__13, 
                    d_arr_merge1_24__12, d_arr_merge1_24__11, 
                    d_arr_merge1_24__10, d_arr_merge1_24__9, d_arr_merge1_24__8, 
                    d_arr_merge1_24__7, d_arr_merge1_24__6, d_arr_merge1_24__5, 
                    d_arr_merge1_24__4, d_arr_merge1_24__3, d_arr_merge1_24__2, 
                    d_arr_merge1_24__1, d_arr_merge1_24__0, d_arr_merge2_0__31, 
                    d_arr_merge2_0__30, d_arr_merge2_0__29, d_arr_merge2_0__28, 
                    d_arr_merge2_0__27, d_arr_merge2_0__26, d_arr_merge2_0__25, 
                    d_arr_merge2_0__24, d_arr_merge2_0__23, d_arr_merge2_0__22, 
                    d_arr_merge2_0__21, d_arr_merge2_0__20, d_arr_merge2_0__19, 
                    d_arr_merge2_0__18, d_arr_merge2_0__17, d_arr_merge2_0__16, 
                    d_arr_merge2_0__15, d_arr_merge2_0__14, d_arr_merge2_0__13, 
                    d_arr_merge2_0__12, d_arr_merge2_0__11, d_arr_merge2_0__10, 
                    d_arr_merge2_0__9, d_arr_merge2_0__8, d_arr_merge2_0__7, 
                    d_arr_merge2_0__6, d_arr_merge2_0__5, d_arr_merge2_0__4, 
                    d_arr_merge2_0__3, d_arr_merge2_0__2, d_arr_merge2_0__1, 
                    d_arr_merge2_0__0, d_arr_merge2_1__31, d_arr_merge2_1__30, 
                    d_arr_merge2_1__29, d_arr_merge2_1__28, d_arr_merge2_1__27, 
                    d_arr_merge2_1__26, d_arr_merge2_1__25, d_arr_merge2_1__24, 
                    d_arr_merge2_1__23, d_arr_merge2_1__22, d_arr_merge2_1__21, 
                    d_arr_merge2_1__20, d_arr_merge2_1__19, d_arr_merge2_1__18, 
                    d_arr_merge2_1__17, d_arr_merge2_1__16, d_arr_merge2_1__15, 
                    d_arr_merge2_1__14, d_arr_merge2_1__13, d_arr_merge2_1__12, 
                    d_arr_merge2_1__11, d_arr_merge2_1__10, d_arr_merge2_1__9, 
                    d_arr_merge2_1__8, d_arr_merge2_1__7, d_arr_merge2_1__6, 
                    d_arr_merge2_1__5, d_arr_merge2_1__4, d_arr_merge2_1__3, 
                    d_arr_merge2_1__2, d_arr_merge2_1__1, d_arr_merge2_1__0, 
                    d_arr_merge2_2__31, d_arr_merge2_2__30, d_arr_merge2_2__29, 
                    d_arr_merge2_2__28, d_arr_merge2_2__27, d_arr_merge2_2__26, 
                    d_arr_merge2_2__25, d_arr_merge2_2__24, d_arr_merge2_2__23, 
                    d_arr_merge2_2__22, d_arr_merge2_2__21, d_arr_merge2_2__20, 
                    d_arr_merge2_2__19, d_arr_merge2_2__18, d_arr_merge2_2__17, 
                    d_arr_merge2_2__16, d_arr_merge2_2__15, d_arr_merge2_2__14, 
                    d_arr_merge2_2__13, d_arr_merge2_2__12, d_arr_merge2_2__11, 
                    d_arr_merge2_2__10, d_arr_merge2_2__9, d_arr_merge2_2__8, 
                    d_arr_merge2_2__7, d_arr_merge2_2__6, d_arr_merge2_2__5, 
                    d_arr_merge2_2__4, d_arr_merge2_2__3, d_arr_merge2_2__2, 
                    d_arr_merge2_2__1, d_arr_merge2_2__0, d_arr_merge2_3__31, 
                    d_arr_merge2_3__30, d_arr_merge2_3__29, d_arr_merge2_3__28, 
                    d_arr_merge2_3__27, d_arr_merge2_3__26, d_arr_merge2_3__25, 
                    d_arr_merge2_3__24, d_arr_merge2_3__23, d_arr_merge2_3__22, 
                    d_arr_merge2_3__21, d_arr_merge2_3__20, d_arr_merge2_3__19, 
                    d_arr_merge2_3__18, d_arr_merge2_3__17, d_arr_merge2_3__16, 
                    d_arr_merge2_3__15, d_arr_merge2_3__14, d_arr_merge2_3__13, 
                    d_arr_merge2_3__12, d_arr_merge2_3__11, d_arr_merge2_3__10, 
                    d_arr_merge2_3__9, d_arr_merge2_3__8, d_arr_merge2_3__7, 
                    d_arr_merge2_3__6, d_arr_merge2_3__5, d_arr_merge2_3__4, 
                    d_arr_merge2_3__3, d_arr_merge2_3__2, d_arr_merge2_3__1, 
                    d_arr_merge2_3__0, d_arr_merge2_4__31, d_arr_merge2_4__30, 
                    d_arr_merge2_4__29, d_arr_merge2_4__28, d_arr_merge2_4__27, 
                    d_arr_merge2_4__26, d_arr_merge2_4__25, d_arr_merge2_4__24, 
                    d_arr_merge2_4__23, d_arr_merge2_4__22, d_arr_merge2_4__21, 
                    d_arr_merge2_4__20, d_arr_merge2_4__19, d_arr_merge2_4__18, 
                    d_arr_merge2_4__17, d_arr_merge2_4__16, d_arr_merge2_4__15, 
                    d_arr_merge2_4__14, d_arr_merge2_4__13, d_arr_merge2_4__12, 
                    d_arr_merge2_4__11, d_arr_merge2_4__10, d_arr_merge2_4__9, 
                    d_arr_merge2_4__8, d_arr_merge2_4__7, d_arr_merge2_4__6, 
                    d_arr_merge2_4__5, d_arr_merge2_4__4, d_arr_merge2_4__3, 
                    d_arr_merge2_4__2, d_arr_merge2_4__1, d_arr_merge2_4__0, 
                    d_arr_merge2_5__31, d_arr_merge2_5__30, d_arr_merge2_5__29, 
                    d_arr_merge2_5__28, d_arr_merge2_5__27, d_arr_merge2_5__26, 
                    d_arr_merge2_5__25, d_arr_merge2_5__24, d_arr_merge2_5__23, 
                    d_arr_merge2_5__22, d_arr_merge2_5__21, d_arr_merge2_5__20, 
                    d_arr_merge2_5__19, d_arr_merge2_5__18, d_arr_merge2_5__17, 
                    d_arr_merge2_5__16, d_arr_merge2_5__15, d_arr_merge2_5__14, 
                    d_arr_merge2_5__13, d_arr_merge2_5__12, d_arr_merge2_5__11, 
                    d_arr_merge2_5__10, d_arr_merge2_5__9, d_arr_merge2_5__8, 
                    d_arr_merge2_5__7, d_arr_merge2_5__6, d_arr_merge2_5__5, 
                    d_arr_merge2_5__4, d_arr_merge2_5__3, d_arr_merge2_5__2, 
                    d_arr_merge2_5__1, d_arr_merge2_5__0, d_arr_merge2_6__31, 
                    d_arr_merge2_6__30, d_arr_merge2_6__29, d_arr_merge2_6__28, 
                    d_arr_merge2_6__27, d_arr_merge2_6__26, d_arr_merge2_6__25, 
                    d_arr_merge2_6__24, d_arr_merge2_6__23, d_arr_merge2_6__22, 
                    d_arr_merge2_6__21, d_arr_merge2_6__20, d_arr_merge2_6__19, 
                    d_arr_merge2_6__18, d_arr_merge2_6__17, d_arr_merge2_6__16, 
                    d_arr_merge2_6__15, d_arr_merge2_6__14, d_arr_merge2_6__13, 
                    d_arr_merge2_6__12, d_arr_merge2_6__11, d_arr_merge2_6__10, 
                    d_arr_merge2_6__9, d_arr_merge2_6__8, d_arr_merge2_6__7, 
                    d_arr_merge2_6__6, d_arr_merge2_6__5, d_arr_merge2_6__4, 
                    d_arr_merge2_6__3, d_arr_merge2_6__2, d_arr_merge2_6__1, 
                    d_arr_merge2_6__0, d_arr_merge2_7__31, d_arr_merge2_7__30, 
                    d_arr_merge2_7__29, d_arr_merge2_7__28, d_arr_merge2_7__27, 
                    d_arr_merge2_7__26, d_arr_merge2_7__25, d_arr_merge2_7__24, 
                    d_arr_merge2_7__23, d_arr_merge2_7__22, d_arr_merge2_7__21, 
                    d_arr_merge2_7__20, d_arr_merge2_7__19, d_arr_merge2_7__18, 
                    d_arr_merge2_7__17, d_arr_merge2_7__16, d_arr_merge2_7__15, 
                    d_arr_merge2_7__14, d_arr_merge2_7__13, d_arr_merge2_7__12, 
                    d_arr_merge2_7__11, d_arr_merge2_7__10, d_arr_merge2_7__9, 
                    d_arr_merge2_7__8, d_arr_merge2_7__7, d_arr_merge2_7__6, 
                    d_arr_merge2_7__5, d_arr_merge2_7__4, d_arr_merge2_7__3, 
                    d_arr_merge2_7__2, d_arr_merge2_7__1, d_arr_merge2_7__0, 
                    d_arr_merge2_8__31, d_arr_merge2_8__30, d_arr_merge2_8__29, 
                    d_arr_merge2_8__28, d_arr_merge2_8__27, d_arr_merge2_8__26, 
                    d_arr_merge2_8__25, d_arr_merge2_8__24, d_arr_merge2_8__23, 
                    d_arr_merge2_8__22, d_arr_merge2_8__21, d_arr_merge2_8__20, 
                    d_arr_merge2_8__19, d_arr_merge2_8__18, d_arr_merge2_8__17, 
                    d_arr_merge2_8__16, d_arr_merge2_8__15, d_arr_merge2_8__14, 
                    d_arr_merge2_8__13, d_arr_merge2_8__12, d_arr_merge2_8__11, 
                    d_arr_merge2_8__10, d_arr_merge2_8__9, d_arr_merge2_8__8, 
                    d_arr_merge2_8__7, d_arr_merge2_8__6, d_arr_merge2_8__5, 
                    d_arr_merge2_8__4, d_arr_merge2_8__3, d_arr_merge2_8__2, 
                    d_arr_merge2_8__1, d_arr_merge2_8__0, d_arr_merge2_9__31, 
                    d_arr_merge2_9__30, d_arr_merge2_9__29, d_arr_merge2_9__28, 
                    d_arr_merge2_9__27, d_arr_merge2_9__26, d_arr_merge2_9__25, 
                    d_arr_merge2_9__24, d_arr_merge2_9__23, d_arr_merge2_9__22, 
                    d_arr_merge2_9__21, d_arr_merge2_9__20, d_arr_merge2_9__19, 
                    d_arr_merge2_9__18, d_arr_merge2_9__17, d_arr_merge2_9__16, 
                    d_arr_merge2_9__15, d_arr_merge2_9__14, d_arr_merge2_9__13, 
                    d_arr_merge2_9__12, d_arr_merge2_9__11, d_arr_merge2_9__10, 
                    d_arr_merge2_9__9, d_arr_merge2_9__8, d_arr_merge2_9__7, 
                    d_arr_merge2_9__6, d_arr_merge2_9__5, d_arr_merge2_9__4, 
                    d_arr_merge2_9__3, d_arr_merge2_9__2, d_arr_merge2_9__1, 
                    d_arr_merge2_9__0, d_arr_merge2_10__31, d_arr_merge2_10__30, 
                    d_arr_merge2_10__29, d_arr_merge2_10__28, 
                    d_arr_merge2_10__27, d_arr_merge2_10__26, 
                    d_arr_merge2_10__25, d_arr_merge2_10__24, 
                    d_arr_merge2_10__23, d_arr_merge2_10__22, 
                    d_arr_merge2_10__21, d_arr_merge2_10__20, 
                    d_arr_merge2_10__19, d_arr_merge2_10__18, 
                    d_arr_merge2_10__17, d_arr_merge2_10__16, 
                    d_arr_merge2_10__15, d_arr_merge2_10__14, 
                    d_arr_merge2_10__13, d_arr_merge2_10__12, 
                    d_arr_merge2_10__11, d_arr_merge2_10__10, d_arr_merge2_10__9, 
                    d_arr_merge2_10__8, d_arr_merge2_10__7, d_arr_merge2_10__6, 
                    d_arr_merge2_10__5, d_arr_merge2_10__4, d_arr_merge2_10__3, 
                    d_arr_merge2_10__2, d_arr_merge2_10__1, d_arr_merge2_10__0, 
                    d_arr_merge2_11__31, d_arr_merge2_11__30, 
                    d_arr_merge2_11__29, d_arr_merge2_11__28, 
                    d_arr_merge2_11__27, d_arr_merge2_11__26, 
                    d_arr_merge2_11__25, d_arr_merge2_11__24, 
                    d_arr_merge2_11__23, d_arr_merge2_11__22, 
                    d_arr_merge2_11__21, d_arr_merge2_11__20, 
                    d_arr_merge2_11__19, d_arr_merge2_11__18, 
                    d_arr_merge2_11__17, d_arr_merge2_11__16, 
                    d_arr_merge2_11__15, d_arr_merge2_11__14, 
                    d_arr_merge2_11__13, d_arr_merge2_11__12, 
                    d_arr_merge2_11__11, d_arr_merge2_11__10, d_arr_merge2_11__9, 
                    d_arr_merge2_11__8, d_arr_merge2_11__7, d_arr_merge2_11__6, 
                    d_arr_merge2_11__5, d_arr_merge2_11__4, d_arr_merge2_11__3, 
                    d_arr_merge2_11__2, d_arr_merge2_11__1, d_arr_merge2_11__0, 
                    d_arr_merge2_12__31, d_arr_merge2_12__30, 
                    d_arr_merge2_12__29, d_arr_merge2_12__28, 
                    d_arr_merge2_12__27, d_arr_merge2_12__26, 
                    d_arr_merge2_12__25, d_arr_merge2_12__24, 
                    d_arr_merge2_12__23, d_arr_merge2_12__22, 
                    d_arr_merge2_12__21, d_arr_merge2_12__20, 
                    d_arr_merge2_12__19, d_arr_merge2_12__18, 
                    d_arr_merge2_12__17, d_arr_merge2_12__16, 
                    d_arr_merge2_12__15, d_arr_merge2_12__14, 
                    d_arr_merge2_12__13, d_arr_merge2_12__12, 
                    d_arr_merge2_12__11, d_arr_merge2_12__10, d_arr_merge2_12__9, 
                    d_arr_merge2_12__8, d_arr_merge2_12__7, d_arr_merge2_12__6, 
                    d_arr_merge2_12__5, d_arr_merge2_12__4, d_arr_merge2_12__3, 
                    d_arr_merge2_12__2, d_arr_merge2_12__1, d_arr_merge2_12__0, 
                    d_arr_merge2_13__31, d_arr_merge2_13__30, 
                    d_arr_merge2_13__29, d_arr_merge2_13__28, 
                    d_arr_merge2_13__27, d_arr_merge2_13__26, 
                    d_arr_merge2_13__25, d_arr_merge2_13__24, 
                    d_arr_merge2_13__23, d_arr_merge2_13__22, 
                    d_arr_merge2_13__21, d_arr_merge2_13__20, 
                    d_arr_merge2_13__19, d_arr_merge2_13__18, 
                    d_arr_merge2_13__17, d_arr_merge2_13__16, 
                    d_arr_merge2_13__15, d_arr_merge2_13__14, 
                    d_arr_merge2_13__13, d_arr_merge2_13__12, 
                    d_arr_merge2_13__11, d_arr_merge2_13__10, d_arr_merge2_13__9, 
                    d_arr_merge2_13__8, d_arr_merge2_13__7, d_arr_merge2_13__6, 
                    d_arr_merge2_13__5, d_arr_merge2_13__4, d_arr_merge2_13__3, 
                    d_arr_merge2_13__2, d_arr_merge2_13__1, d_arr_merge2_13__0, 
                    d_arr_merge2_14__31, d_arr_merge2_14__30, 
                    d_arr_merge2_14__29, d_arr_merge2_14__28, 
                    d_arr_merge2_14__27, d_arr_merge2_14__26, 
                    d_arr_merge2_14__25, d_arr_merge2_14__24, 
                    d_arr_merge2_14__23, d_arr_merge2_14__22, 
                    d_arr_merge2_14__21, d_arr_merge2_14__20, 
                    d_arr_merge2_14__19, d_arr_merge2_14__18, 
                    d_arr_merge2_14__17, d_arr_merge2_14__16, 
                    d_arr_merge2_14__15, d_arr_merge2_14__14, 
                    d_arr_merge2_14__13, d_arr_merge2_14__12, 
                    d_arr_merge2_14__11, d_arr_merge2_14__10, d_arr_merge2_14__9, 
                    d_arr_merge2_14__8, d_arr_merge2_14__7, d_arr_merge2_14__6, 
                    d_arr_merge2_14__5, d_arr_merge2_14__4, d_arr_merge2_14__3, 
                    d_arr_merge2_14__2, d_arr_merge2_14__1, d_arr_merge2_14__0, 
                    d_arr_merge2_15__31, d_arr_merge2_15__30, 
                    d_arr_merge2_15__29, d_arr_merge2_15__28, 
                    d_arr_merge2_15__27, d_arr_merge2_15__26, 
                    d_arr_merge2_15__25, d_arr_merge2_15__24, 
                    d_arr_merge2_15__23, d_arr_merge2_15__22, 
                    d_arr_merge2_15__21, d_arr_merge2_15__20, 
                    d_arr_merge2_15__19, d_arr_merge2_15__18, 
                    d_arr_merge2_15__17, d_arr_merge2_15__16, 
                    d_arr_merge2_15__15, d_arr_merge2_15__14, 
                    d_arr_merge2_15__13, d_arr_merge2_15__12, 
                    d_arr_merge2_15__11, d_arr_merge2_15__10, d_arr_merge2_15__9, 
                    d_arr_merge2_15__8, d_arr_merge2_15__7, d_arr_merge2_15__6, 
                    d_arr_merge2_15__5, d_arr_merge2_15__4, d_arr_merge2_15__3, 
                    d_arr_merge2_15__2, d_arr_merge2_15__1, d_arr_merge2_15__0, 
                    d_arr_merge2_16__31, d_arr_merge2_16__30, 
                    d_arr_merge2_16__29, d_arr_merge2_16__28, 
                    d_arr_merge2_16__27, d_arr_merge2_16__26, 
                    d_arr_merge2_16__25, d_arr_merge2_16__24, 
                    d_arr_merge2_16__23, d_arr_merge2_16__22, 
                    d_arr_merge2_16__21, d_arr_merge2_16__20, 
                    d_arr_merge2_16__19, d_arr_merge2_16__18, 
                    d_arr_merge2_16__17, d_arr_merge2_16__16, 
                    d_arr_merge2_16__15, d_arr_merge2_16__14, 
                    d_arr_merge2_16__13, d_arr_merge2_16__12, 
                    d_arr_merge2_16__11, d_arr_merge2_16__10, d_arr_merge2_16__9, 
                    d_arr_merge2_16__8, d_arr_merge2_16__7, d_arr_merge2_16__6, 
                    d_arr_merge2_16__5, d_arr_merge2_16__4, d_arr_merge2_16__3, 
                    d_arr_merge2_16__2, d_arr_merge2_16__1, d_arr_merge2_16__0, 
                    d_arr_merge2_17__31, d_arr_merge2_17__30, 
                    d_arr_merge2_17__29, d_arr_merge2_17__28, 
                    d_arr_merge2_17__27, d_arr_merge2_17__26, 
                    d_arr_merge2_17__25, d_arr_merge2_17__24, 
                    d_arr_merge2_17__23, d_arr_merge2_17__22, 
                    d_arr_merge2_17__21, d_arr_merge2_17__20, 
                    d_arr_merge2_17__19, d_arr_merge2_17__18, 
                    d_arr_merge2_17__17, d_arr_merge2_17__16, 
                    d_arr_merge2_17__15, d_arr_merge2_17__14, 
                    d_arr_merge2_17__13, d_arr_merge2_17__12, 
                    d_arr_merge2_17__11, d_arr_merge2_17__10, d_arr_merge2_17__9, 
                    d_arr_merge2_17__8, d_arr_merge2_17__7, d_arr_merge2_17__6, 
                    d_arr_merge2_17__5, d_arr_merge2_17__4, d_arr_merge2_17__3, 
                    d_arr_merge2_17__2, d_arr_merge2_17__1, d_arr_merge2_17__0, 
                    d_arr_merge2_18__31, d_arr_merge2_18__30, 
                    d_arr_merge2_18__29, d_arr_merge2_18__28, 
                    d_arr_merge2_18__27, d_arr_merge2_18__26, 
                    d_arr_merge2_18__25, d_arr_merge2_18__24, 
                    d_arr_merge2_18__23, d_arr_merge2_18__22, 
                    d_arr_merge2_18__21, d_arr_merge2_18__20, 
                    d_arr_merge2_18__19, d_arr_merge2_18__18, 
                    d_arr_merge2_18__17, d_arr_merge2_18__16, 
                    d_arr_merge2_18__15, d_arr_merge2_18__14, 
                    d_arr_merge2_18__13, d_arr_merge2_18__12, 
                    d_arr_merge2_18__11, d_arr_merge2_18__10, d_arr_merge2_18__9, 
                    d_arr_merge2_18__8, d_arr_merge2_18__7, d_arr_merge2_18__6, 
                    d_arr_merge2_18__5, d_arr_merge2_18__4, d_arr_merge2_18__3, 
                    d_arr_merge2_18__2, d_arr_merge2_18__1, d_arr_merge2_18__0, 
                    d_arr_merge2_19__31, d_arr_merge2_19__30, 
                    d_arr_merge2_19__29, d_arr_merge2_19__28, 
                    d_arr_merge2_19__27, d_arr_merge2_19__26, 
                    d_arr_merge2_19__25, d_arr_merge2_19__24, 
                    d_arr_merge2_19__23, d_arr_merge2_19__22, 
                    d_arr_merge2_19__21, d_arr_merge2_19__20, 
                    d_arr_merge2_19__19, d_arr_merge2_19__18, 
                    d_arr_merge2_19__17, d_arr_merge2_19__16, 
                    d_arr_merge2_19__15, d_arr_merge2_19__14, 
                    d_arr_merge2_19__13, d_arr_merge2_19__12, 
                    d_arr_merge2_19__11, d_arr_merge2_19__10, d_arr_merge2_19__9, 
                    d_arr_merge2_19__8, d_arr_merge2_19__7, d_arr_merge2_19__6, 
                    d_arr_merge2_19__5, d_arr_merge2_19__4, d_arr_merge2_19__3, 
                    d_arr_merge2_19__2, d_arr_merge2_19__1, d_arr_merge2_19__0, 
                    d_arr_merge2_20__31, d_arr_merge2_20__30, 
                    d_arr_merge2_20__29, d_arr_merge2_20__28, 
                    d_arr_merge2_20__27, d_arr_merge2_20__26, 
                    d_arr_merge2_20__25, d_arr_merge2_20__24, 
                    d_arr_merge2_20__23, d_arr_merge2_20__22, 
                    d_arr_merge2_20__21, d_arr_merge2_20__20, 
                    d_arr_merge2_20__19, d_arr_merge2_20__18, 
                    d_arr_merge2_20__17, d_arr_merge2_20__16, 
                    d_arr_merge2_20__15, d_arr_merge2_20__14, 
                    d_arr_merge2_20__13, d_arr_merge2_20__12, 
                    d_arr_merge2_20__11, d_arr_merge2_20__10, d_arr_merge2_20__9, 
                    d_arr_merge2_20__8, d_arr_merge2_20__7, d_arr_merge2_20__6, 
                    d_arr_merge2_20__5, d_arr_merge2_20__4, d_arr_merge2_20__3, 
                    d_arr_merge2_20__2, d_arr_merge2_20__1, d_arr_merge2_20__0, 
                    d_arr_merge2_21__31, d_arr_merge2_21__30, 
                    d_arr_merge2_21__29, d_arr_merge2_21__28, 
                    d_arr_merge2_21__27, d_arr_merge2_21__26, 
                    d_arr_merge2_21__25, d_arr_merge2_21__24, 
                    d_arr_merge2_21__23, d_arr_merge2_21__22, 
                    d_arr_merge2_21__21, d_arr_merge2_21__20, 
                    d_arr_merge2_21__19, d_arr_merge2_21__18, 
                    d_arr_merge2_21__17, d_arr_merge2_21__16, 
                    d_arr_merge2_21__15, d_arr_merge2_21__14, 
                    d_arr_merge2_21__13, d_arr_merge2_21__12, 
                    d_arr_merge2_21__11, d_arr_merge2_21__10, d_arr_merge2_21__9, 
                    d_arr_merge2_21__8, d_arr_merge2_21__7, d_arr_merge2_21__6, 
                    d_arr_merge2_21__5, d_arr_merge2_21__4, d_arr_merge2_21__3, 
                    d_arr_merge2_21__2, d_arr_merge2_21__1, d_arr_merge2_21__0, 
                    d_arr_merge2_22__31, d_arr_merge2_22__30, 
                    d_arr_merge2_22__29, d_arr_merge2_22__28, 
                    d_arr_merge2_22__27, d_arr_merge2_22__26, 
                    d_arr_merge2_22__25, d_arr_merge2_22__24, 
                    d_arr_merge2_22__23, d_arr_merge2_22__22, 
                    d_arr_merge2_22__21, d_arr_merge2_22__20, 
                    d_arr_merge2_22__19, d_arr_merge2_22__18, 
                    d_arr_merge2_22__17, d_arr_merge2_22__16, 
                    d_arr_merge2_22__15, d_arr_merge2_22__14, 
                    d_arr_merge2_22__13, d_arr_merge2_22__12, 
                    d_arr_merge2_22__11, d_arr_merge2_22__10, d_arr_merge2_22__9, 
                    d_arr_merge2_22__8, d_arr_merge2_22__7, d_arr_merge2_22__6, 
                    d_arr_merge2_22__5, d_arr_merge2_22__4, d_arr_merge2_22__3, 
                    d_arr_merge2_22__2, d_arr_merge2_22__1, d_arr_merge2_22__0, 
                    d_arr_merge2_23__31, d_arr_merge2_23__30, 
                    d_arr_merge2_23__29, d_arr_merge2_23__28, 
                    d_arr_merge2_23__27, d_arr_merge2_23__26, 
                    d_arr_merge2_23__25, d_arr_merge2_23__24, 
                    d_arr_merge2_23__23, d_arr_merge2_23__22, 
                    d_arr_merge2_23__21, d_arr_merge2_23__20, 
                    d_arr_merge2_23__19, d_arr_merge2_23__18, 
                    d_arr_merge2_23__17, d_arr_merge2_23__16, 
                    d_arr_merge2_23__15, d_arr_merge2_23__14, 
                    d_arr_merge2_23__13, d_arr_merge2_23__12, 
                    d_arr_merge2_23__11, d_arr_merge2_23__10, d_arr_merge2_23__9, 
                    d_arr_merge2_23__8, d_arr_merge2_23__7, d_arr_merge2_23__6, 
                    d_arr_merge2_23__5, d_arr_merge2_23__4, d_arr_merge2_23__3, 
                    d_arr_merge2_23__2, d_arr_merge2_23__1, d_arr_merge2_23__0, 
                    d_arr_merge2_24__31, d_arr_merge2_24__30, 
                    d_arr_merge2_24__29, d_arr_merge2_24__28, 
                    d_arr_merge2_24__27, d_arr_merge2_24__26, 
                    d_arr_merge2_24__25, d_arr_merge2_24__24, 
                    d_arr_merge2_24__23, d_arr_merge2_24__22, 
                    d_arr_merge2_24__21, d_arr_merge2_24__20, 
                    d_arr_merge2_24__19, d_arr_merge2_24__18, 
                    d_arr_merge2_24__17, d_arr_merge2_24__16, 
                    d_arr_merge2_24__15, d_arr_merge2_24__14, 
                    d_arr_merge2_24__13, d_arr_merge2_24__12, 
                    d_arr_merge2_24__11, d_arr_merge2_24__10, d_arr_merge2_24__9, 
                    d_arr_merge2_24__8, d_arr_merge2_24__7, d_arr_merge2_24__6, 
                    d_arr_merge2_24__5, d_arr_merge2_24__4, d_arr_merge2_24__3, 
                    d_arr_merge2_24__2, d_arr_merge2_24__1, d_arr_merge2_24__0, 
                    d_arr_relu_0__31, d_arr_relu_0__30, d_arr_relu_0__29, 
                    d_arr_relu_0__28, d_arr_relu_0__27, d_arr_relu_0__26, 
                    d_arr_relu_0__25, d_arr_relu_0__24, d_arr_relu_0__23, 
                    d_arr_relu_0__22, d_arr_relu_0__21, d_arr_relu_0__20, 
                    d_arr_relu_0__19, d_arr_relu_0__18, d_arr_relu_0__17, 
                    d_arr_relu_0__16, d_arr_relu_0__15, d_arr_relu_0__14, 
                    d_arr_relu_0__13, d_arr_relu_0__12, d_arr_relu_0__11, 
                    d_arr_relu_0__10, d_arr_relu_0__9, d_arr_relu_0__8, 
                    d_arr_relu_0__7, d_arr_relu_0__6, d_arr_relu_0__5, 
                    d_arr_relu_0__4, d_arr_relu_0__3, d_arr_relu_0__2, 
                    d_arr_relu_0__1, d_arr_relu_0__0, d_arr_relu_1__31, 
                    d_arr_relu_1__30, d_arr_relu_1__29, d_arr_relu_1__28, 
                    d_arr_relu_1__27, d_arr_relu_1__26, d_arr_relu_1__25, 
                    d_arr_relu_1__24, d_arr_relu_1__23, d_arr_relu_1__22, 
                    d_arr_relu_1__21, d_arr_relu_1__20, d_arr_relu_1__19, 
                    d_arr_relu_1__18, d_arr_relu_1__17, d_arr_relu_1__16, 
                    d_arr_relu_1__15, d_arr_relu_1__14, d_arr_relu_1__13, 
                    d_arr_relu_1__12, d_arr_relu_1__11, d_arr_relu_1__10, 
                    d_arr_relu_1__9, d_arr_relu_1__8, d_arr_relu_1__7, 
                    d_arr_relu_1__6, d_arr_relu_1__5, d_arr_relu_1__4, 
                    d_arr_relu_1__3, d_arr_relu_1__2, d_arr_relu_1__1, 
                    d_arr_relu_1__0, d_arr_relu_2__31, d_arr_relu_2__30, 
                    d_arr_relu_2__29, d_arr_relu_2__28, d_arr_relu_2__27, 
                    d_arr_relu_2__26, d_arr_relu_2__25, d_arr_relu_2__24, 
                    d_arr_relu_2__23, d_arr_relu_2__22, d_arr_relu_2__21, 
                    d_arr_relu_2__20, d_arr_relu_2__19, d_arr_relu_2__18, 
                    d_arr_relu_2__17, d_arr_relu_2__16, d_arr_relu_2__15, 
                    d_arr_relu_2__14, d_arr_relu_2__13, d_arr_relu_2__12, 
                    d_arr_relu_2__11, d_arr_relu_2__10, d_arr_relu_2__9, 
                    d_arr_relu_2__8, d_arr_relu_2__7, d_arr_relu_2__6, 
                    d_arr_relu_2__5, d_arr_relu_2__4, d_arr_relu_2__3, 
                    d_arr_relu_2__2, d_arr_relu_2__1, d_arr_relu_2__0, 
                    d_arr_relu_3__31, d_arr_relu_3__30, d_arr_relu_3__29, 
                    d_arr_relu_3__28, d_arr_relu_3__27, d_arr_relu_3__26, 
                    d_arr_relu_3__25, d_arr_relu_3__24, d_arr_relu_3__23, 
                    d_arr_relu_3__22, d_arr_relu_3__21, d_arr_relu_3__20, 
                    d_arr_relu_3__19, d_arr_relu_3__18, d_arr_relu_3__17, 
                    d_arr_relu_3__16, d_arr_relu_3__15, d_arr_relu_3__14, 
                    d_arr_relu_3__13, d_arr_relu_3__12, d_arr_relu_3__11, 
                    d_arr_relu_3__10, d_arr_relu_3__9, d_arr_relu_3__8, 
                    d_arr_relu_3__7, d_arr_relu_3__6, d_arr_relu_3__5, 
                    d_arr_relu_3__4, d_arr_relu_3__3, d_arr_relu_3__2, 
                    d_arr_relu_3__1, d_arr_relu_3__0, d_arr_relu_4__31, 
                    d_arr_relu_4__30, d_arr_relu_4__29, d_arr_relu_4__28, 
                    d_arr_relu_4__27, d_arr_relu_4__26, d_arr_relu_4__25, 
                    d_arr_relu_4__24, d_arr_relu_4__23, d_arr_relu_4__22, 
                    d_arr_relu_4__21, d_arr_relu_4__20, d_arr_relu_4__19, 
                    d_arr_relu_4__18, d_arr_relu_4__17, d_arr_relu_4__16, 
                    d_arr_relu_4__15, d_arr_relu_4__14, d_arr_relu_4__13, 
                    d_arr_relu_4__12, d_arr_relu_4__11, d_arr_relu_4__10, 
                    d_arr_relu_4__9, d_arr_relu_4__8, d_arr_relu_4__7, 
                    d_arr_relu_4__6, d_arr_relu_4__5, d_arr_relu_4__4, 
                    d_arr_relu_4__3, d_arr_relu_4__2, d_arr_relu_4__1, 
                    d_arr_relu_4__0, d_arr_relu_5__31, d_arr_relu_5__30, 
                    d_arr_relu_5__29, d_arr_relu_5__28, d_arr_relu_5__27, 
                    d_arr_relu_5__26, d_arr_relu_5__25, d_arr_relu_5__24, 
                    d_arr_relu_5__23, d_arr_relu_5__22, d_arr_relu_5__21, 
                    d_arr_relu_5__20, d_arr_relu_5__19, d_arr_relu_5__18, 
                    d_arr_relu_5__17, d_arr_relu_5__16, d_arr_relu_5__15, 
                    d_arr_relu_5__14, d_arr_relu_5__13, d_arr_relu_5__12, 
                    d_arr_relu_5__11, d_arr_relu_5__10, d_arr_relu_5__9, 
                    d_arr_relu_5__8, d_arr_relu_5__7, d_arr_relu_5__6, 
                    d_arr_relu_5__5, d_arr_relu_5__4, d_arr_relu_5__3, 
                    d_arr_relu_5__2, d_arr_relu_5__1, d_arr_relu_5__0, 
                    d_arr_relu_6__31, d_arr_relu_6__30, d_arr_relu_6__29, 
                    d_arr_relu_6__28, d_arr_relu_6__27, d_arr_relu_6__26, 
                    d_arr_relu_6__25, d_arr_relu_6__24, d_arr_relu_6__23, 
                    d_arr_relu_6__22, d_arr_relu_6__21, d_arr_relu_6__20, 
                    d_arr_relu_6__19, d_arr_relu_6__18, d_arr_relu_6__17, 
                    d_arr_relu_6__16, d_arr_relu_6__15, d_arr_relu_6__14, 
                    d_arr_relu_6__13, d_arr_relu_6__12, d_arr_relu_6__11, 
                    d_arr_relu_6__10, d_arr_relu_6__9, d_arr_relu_6__8, 
                    d_arr_relu_6__7, d_arr_relu_6__6, d_arr_relu_6__5, 
                    d_arr_relu_6__4, d_arr_relu_6__3, d_arr_relu_6__2, 
                    d_arr_relu_6__1, d_arr_relu_6__0, d_arr_relu_7__31, 
                    d_arr_relu_7__30, d_arr_relu_7__29, d_arr_relu_7__28, 
                    d_arr_relu_7__27, d_arr_relu_7__26, d_arr_relu_7__25, 
                    d_arr_relu_7__24, d_arr_relu_7__23, d_arr_relu_7__22, 
                    d_arr_relu_7__21, d_arr_relu_7__20, d_arr_relu_7__19, 
                    d_arr_relu_7__18, d_arr_relu_7__17, d_arr_relu_7__16, 
                    d_arr_relu_7__15, d_arr_relu_7__14, d_arr_relu_7__13, 
                    d_arr_relu_7__12, d_arr_relu_7__11, d_arr_relu_7__10, 
                    d_arr_relu_7__9, d_arr_relu_7__8, d_arr_relu_7__7, 
                    d_arr_relu_7__6, d_arr_relu_7__5, d_arr_relu_7__4, 
                    d_arr_relu_7__3, d_arr_relu_7__2, d_arr_relu_7__1, 
                    d_arr_relu_7__0, d_arr_relu_8__31, d_arr_relu_8__30, 
                    d_arr_relu_8__29, d_arr_relu_8__28, d_arr_relu_8__27, 
                    d_arr_relu_8__26, d_arr_relu_8__25, d_arr_relu_8__24, 
                    d_arr_relu_8__23, d_arr_relu_8__22, d_arr_relu_8__21, 
                    d_arr_relu_8__20, d_arr_relu_8__19, d_arr_relu_8__18, 
                    d_arr_relu_8__17, d_arr_relu_8__16, d_arr_relu_8__15, 
                    d_arr_relu_8__14, d_arr_relu_8__13, d_arr_relu_8__12, 
                    d_arr_relu_8__11, d_arr_relu_8__10, d_arr_relu_8__9, 
                    d_arr_relu_8__8, d_arr_relu_8__7, d_arr_relu_8__6, 
                    d_arr_relu_8__5, d_arr_relu_8__4, d_arr_relu_8__3, 
                    d_arr_relu_8__2, d_arr_relu_8__1, d_arr_relu_8__0, 
                    d_arr_relu_9__31, d_arr_relu_9__30, d_arr_relu_9__29, 
                    d_arr_relu_9__28, d_arr_relu_9__27, d_arr_relu_9__26, 
                    d_arr_relu_9__25, d_arr_relu_9__24, d_arr_relu_9__23, 
                    d_arr_relu_9__22, d_arr_relu_9__21, d_arr_relu_9__20, 
                    d_arr_relu_9__19, d_arr_relu_9__18, d_arr_relu_9__17, 
                    d_arr_relu_9__16, d_arr_relu_9__15, d_arr_relu_9__14, 
                    d_arr_relu_9__13, d_arr_relu_9__12, d_arr_relu_9__11, 
                    d_arr_relu_9__10, d_arr_relu_9__9, d_arr_relu_9__8, 
                    d_arr_relu_9__7, d_arr_relu_9__6, d_arr_relu_9__5, 
                    d_arr_relu_9__4, d_arr_relu_9__3, d_arr_relu_9__2, 
                    d_arr_relu_9__1, d_arr_relu_9__0, d_arr_relu_10__31, 
                    d_arr_relu_10__30, d_arr_relu_10__29, d_arr_relu_10__28, 
                    d_arr_relu_10__27, d_arr_relu_10__26, d_arr_relu_10__25, 
                    d_arr_relu_10__24, d_arr_relu_10__23, d_arr_relu_10__22, 
                    d_arr_relu_10__21, d_arr_relu_10__20, d_arr_relu_10__19, 
                    d_arr_relu_10__18, d_arr_relu_10__17, d_arr_relu_10__16, 
                    d_arr_relu_10__15, d_arr_relu_10__14, d_arr_relu_10__13, 
                    d_arr_relu_10__12, d_arr_relu_10__11, d_arr_relu_10__10, 
                    d_arr_relu_10__9, d_arr_relu_10__8, d_arr_relu_10__7, 
                    d_arr_relu_10__6, d_arr_relu_10__5, d_arr_relu_10__4, 
                    d_arr_relu_10__3, d_arr_relu_10__2, d_arr_relu_10__1, 
                    d_arr_relu_10__0, d_arr_relu_11__31, d_arr_relu_11__30, 
                    d_arr_relu_11__29, d_arr_relu_11__28, d_arr_relu_11__27, 
                    d_arr_relu_11__26, d_arr_relu_11__25, d_arr_relu_11__24, 
                    d_arr_relu_11__23, d_arr_relu_11__22, d_arr_relu_11__21, 
                    d_arr_relu_11__20, d_arr_relu_11__19, d_arr_relu_11__18, 
                    d_arr_relu_11__17, d_arr_relu_11__16, d_arr_relu_11__15, 
                    d_arr_relu_11__14, d_arr_relu_11__13, d_arr_relu_11__12, 
                    d_arr_relu_11__11, d_arr_relu_11__10, d_arr_relu_11__9, 
                    d_arr_relu_11__8, d_arr_relu_11__7, d_arr_relu_11__6, 
                    d_arr_relu_11__5, d_arr_relu_11__4, d_arr_relu_11__3, 
                    d_arr_relu_11__2, d_arr_relu_11__1, d_arr_relu_11__0, 
                    d_arr_relu_12__31, d_arr_relu_12__30, d_arr_relu_12__29, 
                    d_arr_relu_12__28, d_arr_relu_12__27, d_arr_relu_12__26, 
                    d_arr_relu_12__25, d_arr_relu_12__24, d_arr_relu_12__23, 
                    d_arr_relu_12__22, d_arr_relu_12__21, d_arr_relu_12__20, 
                    d_arr_relu_12__19, d_arr_relu_12__18, d_arr_relu_12__17, 
                    d_arr_relu_12__16, d_arr_relu_12__15, d_arr_relu_12__14, 
                    d_arr_relu_12__13, d_arr_relu_12__12, d_arr_relu_12__11, 
                    d_arr_relu_12__10, d_arr_relu_12__9, d_arr_relu_12__8, 
                    d_arr_relu_12__7, d_arr_relu_12__6, d_arr_relu_12__5, 
                    d_arr_relu_12__4, d_arr_relu_12__3, d_arr_relu_12__2, 
                    d_arr_relu_12__1, d_arr_relu_12__0, d_arr_relu_13__31, 
                    d_arr_relu_13__30, d_arr_relu_13__29, d_arr_relu_13__28, 
                    d_arr_relu_13__27, d_arr_relu_13__26, d_arr_relu_13__25, 
                    d_arr_relu_13__24, d_arr_relu_13__23, d_arr_relu_13__22, 
                    d_arr_relu_13__21, d_arr_relu_13__20, d_arr_relu_13__19, 
                    d_arr_relu_13__18, d_arr_relu_13__17, d_arr_relu_13__16, 
                    d_arr_relu_13__15, d_arr_relu_13__14, d_arr_relu_13__13, 
                    d_arr_relu_13__12, d_arr_relu_13__11, d_arr_relu_13__10, 
                    d_arr_relu_13__9, d_arr_relu_13__8, d_arr_relu_13__7, 
                    d_arr_relu_13__6, d_arr_relu_13__5, d_arr_relu_13__4, 
                    d_arr_relu_13__3, d_arr_relu_13__2, d_arr_relu_13__1, 
                    d_arr_relu_13__0, d_arr_relu_14__31, d_arr_relu_14__30, 
                    d_arr_relu_14__29, d_arr_relu_14__28, d_arr_relu_14__27, 
                    d_arr_relu_14__26, d_arr_relu_14__25, d_arr_relu_14__24, 
                    d_arr_relu_14__23, d_arr_relu_14__22, d_arr_relu_14__21, 
                    d_arr_relu_14__20, d_arr_relu_14__19, d_arr_relu_14__18, 
                    d_arr_relu_14__17, d_arr_relu_14__16, d_arr_relu_14__15, 
                    d_arr_relu_14__14, d_arr_relu_14__13, d_arr_relu_14__12, 
                    d_arr_relu_14__11, d_arr_relu_14__10, d_arr_relu_14__9, 
                    d_arr_relu_14__8, d_arr_relu_14__7, d_arr_relu_14__6, 
                    d_arr_relu_14__5, d_arr_relu_14__4, d_arr_relu_14__3, 
                    d_arr_relu_14__2, d_arr_relu_14__1, d_arr_relu_14__0, 
                    d_arr_relu_15__31, d_arr_relu_15__30, d_arr_relu_15__29, 
                    d_arr_relu_15__28, d_arr_relu_15__27, d_arr_relu_15__26, 
                    d_arr_relu_15__25, d_arr_relu_15__24, d_arr_relu_15__23, 
                    d_arr_relu_15__22, d_arr_relu_15__21, d_arr_relu_15__20, 
                    d_arr_relu_15__19, d_arr_relu_15__18, d_arr_relu_15__17, 
                    d_arr_relu_15__16, d_arr_relu_15__15, d_arr_relu_15__14, 
                    d_arr_relu_15__13, d_arr_relu_15__12, d_arr_relu_15__11, 
                    d_arr_relu_15__10, d_arr_relu_15__9, d_arr_relu_15__8, 
                    d_arr_relu_15__7, d_arr_relu_15__6, d_arr_relu_15__5, 
                    d_arr_relu_15__4, d_arr_relu_15__3, d_arr_relu_15__2, 
                    d_arr_relu_15__1, d_arr_relu_15__0, d_arr_relu_16__31, 
                    d_arr_relu_16__30, d_arr_relu_16__29, d_arr_relu_16__28, 
                    d_arr_relu_16__27, d_arr_relu_16__26, d_arr_relu_16__25, 
                    d_arr_relu_16__24, d_arr_relu_16__23, d_arr_relu_16__22, 
                    d_arr_relu_16__21, d_arr_relu_16__20, d_arr_relu_16__19, 
                    d_arr_relu_16__18, d_arr_relu_16__17, d_arr_relu_16__16, 
                    d_arr_relu_16__15, d_arr_relu_16__14, d_arr_relu_16__13, 
                    d_arr_relu_16__12, d_arr_relu_16__11, d_arr_relu_16__10, 
                    d_arr_relu_16__9, d_arr_relu_16__8, d_arr_relu_16__7, 
                    d_arr_relu_16__6, d_arr_relu_16__5, d_arr_relu_16__4, 
                    d_arr_relu_16__3, d_arr_relu_16__2, d_arr_relu_16__1, 
                    d_arr_relu_16__0, d_arr_relu_17__31, d_arr_relu_17__30, 
                    d_arr_relu_17__29, d_arr_relu_17__28, d_arr_relu_17__27, 
                    d_arr_relu_17__26, d_arr_relu_17__25, d_arr_relu_17__24, 
                    d_arr_relu_17__23, d_arr_relu_17__22, d_arr_relu_17__21, 
                    d_arr_relu_17__20, d_arr_relu_17__19, d_arr_relu_17__18, 
                    d_arr_relu_17__17, d_arr_relu_17__16, d_arr_relu_17__15, 
                    d_arr_relu_17__14, d_arr_relu_17__13, d_arr_relu_17__12, 
                    d_arr_relu_17__11, d_arr_relu_17__10, d_arr_relu_17__9, 
                    d_arr_relu_17__8, d_arr_relu_17__7, d_arr_relu_17__6, 
                    d_arr_relu_17__5, d_arr_relu_17__4, d_arr_relu_17__3, 
                    d_arr_relu_17__2, d_arr_relu_17__1, d_arr_relu_17__0, 
                    d_arr_relu_18__31, d_arr_relu_18__30, d_arr_relu_18__29, 
                    d_arr_relu_18__28, d_arr_relu_18__27, d_arr_relu_18__26, 
                    d_arr_relu_18__25, d_arr_relu_18__24, d_arr_relu_18__23, 
                    d_arr_relu_18__22, d_arr_relu_18__21, d_arr_relu_18__20, 
                    d_arr_relu_18__19, d_arr_relu_18__18, d_arr_relu_18__17, 
                    d_arr_relu_18__16, d_arr_relu_18__15, d_arr_relu_18__14, 
                    d_arr_relu_18__13, d_arr_relu_18__12, d_arr_relu_18__11, 
                    d_arr_relu_18__10, d_arr_relu_18__9, d_arr_relu_18__8, 
                    d_arr_relu_18__7, d_arr_relu_18__6, d_arr_relu_18__5, 
                    d_arr_relu_18__4, d_arr_relu_18__3, d_arr_relu_18__2, 
                    d_arr_relu_18__1, d_arr_relu_18__0, d_arr_relu_19__31, 
                    d_arr_relu_19__30, d_arr_relu_19__29, d_arr_relu_19__28, 
                    d_arr_relu_19__27, d_arr_relu_19__26, d_arr_relu_19__25, 
                    d_arr_relu_19__24, d_arr_relu_19__23, d_arr_relu_19__22, 
                    d_arr_relu_19__21, d_arr_relu_19__20, d_arr_relu_19__19, 
                    d_arr_relu_19__18, d_arr_relu_19__17, d_arr_relu_19__16, 
                    d_arr_relu_19__15, d_arr_relu_19__14, d_arr_relu_19__13, 
                    d_arr_relu_19__12, d_arr_relu_19__11, d_arr_relu_19__10, 
                    d_arr_relu_19__9, d_arr_relu_19__8, d_arr_relu_19__7, 
                    d_arr_relu_19__6, d_arr_relu_19__5, d_arr_relu_19__4, 
                    d_arr_relu_19__3, d_arr_relu_19__2, d_arr_relu_19__1, 
                    d_arr_relu_19__0, d_arr_relu_20__31, d_arr_relu_20__30, 
                    d_arr_relu_20__29, d_arr_relu_20__28, d_arr_relu_20__27, 
                    d_arr_relu_20__26, d_arr_relu_20__25, d_arr_relu_20__24, 
                    d_arr_relu_20__23, d_arr_relu_20__22, d_arr_relu_20__21, 
                    d_arr_relu_20__20, d_arr_relu_20__19, d_arr_relu_20__18, 
                    d_arr_relu_20__17, d_arr_relu_20__16, d_arr_relu_20__15, 
                    d_arr_relu_20__14, d_arr_relu_20__13, d_arr_relu_20__12, 
                    d_arr_relu_20__11, d_arr_relu_20__10, d_arr_relu_20__9, 
                    d_arr_relu_20__8, d_arr_relu_20__7, d_arr_relu_20__6, 
                    d_arr_relu_20__5, d_arr_relu_20__4, d_arr_relu_20__3, 
                    d_arr_relu_20__2, d_arr_relu_20__1, d_arr_relu_20__0, 
                    d_arr_relu_21__31, d_arr_relu_21__30, d_arr_relu_21__29, 
                    d_arr_relu_21__28, d_arr_relu_21__27, d_arr_relu_21__26, 
                    d_arr_relu_21__25, d_arr_relu_21__24, d_arr_relu_21__23, 
                    d_arr_relu_21__22, d_arr_relu_21__21, d_arr_relu_21__20, 
                    d_arr_relu_21__19, d_arr_relu_21__18, d_arr_relu_21__17, 
                    d_arr_relu_21__16, d_arr_relu_21__15, d_arr_relu_21__14, 
                    d_arr_relu_21__13, d_arr_relu_21__12, d_arr_relu_21__11, 
                    d_arr_relu_21__10, d_arr_relu_21__9, d_arr_relu_21__8, 
                    d_arr_relu_21__7, d_arr_relu_21__6, d_arr_relu_21__5, 
                    d_arr_relu_21__4, d_arr_relu_21__3, d_arr_relu_21__2, 
                    d_arr_relu_21__1, d_arr_relu_21__0, d_arr_relu_22__31, 
                    d_arr_relu_22__30, d_arr_relu_22__29, d_arr_relu_22__28, 
                    d_arr_relu_22__27, d_arr_relu_22__26, d_arr_relu_22__25, 
                    d_arr_relu_22__24, d_arr_relu_22__23, d_arr_relu_22__22, 
                    d_arr_relu_22__21, d_arr_relu_22__20, d_arr_relu_22__19, 
                    d_arr_relu_22__18, d_arr_relu_22__17, d_arr_relu_22__16, 
                    d_arr_relu_22__15, d_arr_relu_22__14, d_arr_relu_22__13, 
                    d_arr_relu_22__12, d_arr_relu_22__11, d_arr_relu_22__10, 
                    d_arr_relu_22__9, d_arr_relu_22__8, d_arr_relu_22__7, 
                    d_arr_relu_22__6, d_arr_relu_22__5, d_arr_relu_22__4, 
                    d_arr_relu_22__3, d_arr_relu_22__2, d_arr_relu_22__1, 
                    d_arr_relu_22__0, d_arr_relu_23__31, d_arr_relu_23__30, 
                    d_arr_relu_23__29, d_arr_relu_23__28, d_arr_relu_23__27, 
                    d_arr_relu_23__26, d_arr_relu_23__25, d_arr_relu_23__24, 
                    d_arr_relu_23__23, d_arr_relu_23__22, d_arr_relu_23__21, 
                    d_arr_relu_23__20, d_arr_relu_23__19, d_arr_relu_23__18, 
                    d_arr_relu_23__17, d_arr_relu_23__16, d_arr_relu_23__15, 
                    d_arr_relu_23__14, d_arr_relu_23__13, d_arr_relu_23__12, 
                    d_arr_relu_23__11, d_arr_relu_23__10, d_arr_relu_23__9, 
                    d_arr_relu_23__8, d_arr_relu_23__7, d_arr_relu_23__6, 
                    d_arr_relu_23__5, d_arr_relu_23__4, d_arr_relu_23__3, 
                    d_arr_relu_23__2, d_arr_relu_23__1, d_arr_relu_23__0, 
                    d_arr_relu_24__31, d_arr_relu_24__30, d_arr_relu_24__29, 
                    d_arr_relu_24__28, d_arr_relu_24__27, d_arr_relu_24__26, 
                    d_arr_relu_24__25, d_arr_relu_24__24, d_arr_relu_24__23, 
                    d_arr_relu_24__22, d_arr_relu_24__21, d_arr_relu_24__20, 
                    d_arr_relu_24__19, d_arr_relu_24__18, d_arr_relu_24__17, 
                    d_arr_relu_24__16, d_arr_relu_24__15, d_arr_relu_24__14, 
                    d_arr_relu_24__13, d_arr_relu_24__12, d_arr_relu_24__11, 
                    d_arr_relu_24__10, d_arr_relu_24__9, d_arr_relu_24__8, 
                    d_arr_relu_24__7, d_arr_relu_24__6, d_arr_relu_24__5, 
                    d_arr_relu_24__4, d_arr_relu_24__3, d_arr_relu_24__2, 
                    d_arr_relu_24__1, d_arr_relu_24__0, sel_mux, sel_mul, 
                    sel_add, sel_merge1, sel_merge2, sel_relu, d_arr_0__31, 
                    d_arr_0__30, d_arr_0__29, d_arr_0__28, d_arr_0__27, 
                    d_arr_0__26, d_arr_0__25, d_arr_0__24, d_arr_0__23, 
                    d_arr_0__22, d_arr_0__21, d_arr_0__20, d_arr_0__19, 
                    d_arr_0__18, d_arr_0__17, d_arr_0__16, d_arr_0__15, 
                    d_arr_0__14, d_arr_0__13, d_arr_0__12, d_arr_0__11, 
                    d_arr_0__10, d_arr_0__9, d_arr_0__8, d_arr_0__7, d_arr_0__6, 
                    d_arr_0__5, d_arr_0__4, d_arr_0__3, d_arr_0__2, d_arr_0__1, 
                    d_arr_0__0, d_arr_1__31, d_arr_1__30, d_arr_1__29, 
                    d_arr_1__28, d_arr_1__27, d_arr_1__26, d_arr_1__25, 
                    d_arr_1__24, d_arr_1__23, d_arr_1__22, d_arr_1__21, 
                    d_arr_1__20, d_arr_1__19, d_arr_1__18, d_arr_1__17, 
                    d_arr_1__16, d_arr_1__15, d_arr_1__14, d_arr_1__13, 
                    d_arr_1__12, d_arr_1__11, d_arr_1__10, d_arr_1__9, 
                    d_arr_1__8, d_arr_1__7, d_arr_1__6, d_arr_1__5, d_arr_1__4, 
                    d_arr_1__3, d_arr_1__2, d_arr_1__1, d_arr_1__0, d_arr_2__31, 
                    d_arr_2__30, d_arr_2__29, d_arr_2__28, d_arr_2__27, 
                    d_arr_2__26, d_arr_2__25, d_arr_2__24, d_arr_2__23, 
                    d_arr_2__22, d_arr_2__21, d_arr_2__20, d_arr_2__19, 
                    d_arr_2__18, d_arr_2__17, d_arr_2__16, d_arr_2__15, 
                    d_arr_2__14, d_arr_2__13, d_arr_2__12, d_arr_2__11, 
                    d_arr_2__10, d_arr_2__9, d_arr_2__8, d_arr_2__7, d_arr_2__6, 
                    d_arr_2__5, d_arr_2__4, d_arr_2__3, d_arr_2__2, d_arr_2__1, 
                    d_arr_2__0, d_arr_3__31, d_arr_3__30, d_arr_3__29, 
                    d_arr_3__28, d_arr_3__27, d_arr_3__26, d_arr_3__25, 
                    d_arr_3__24, d_arr_3__23, d_arr_3__22, d_arr_3__21, 
                    d_arr_3__20, d_arr_3__19, d_arr_3__18, d_arr_3__17, 
                    d_arr_3__16, d_arr_3__15, d_arr_3__14, d_arr_3__13, 
                    d_arr_3__12, d_arr_3__11, d_arr_3__10, d_arr_3__9, 
                    d_arr_3__8, d_arr_3__7, d_arr_3__6, d_arr_3__5, d_arr_3__4, 
                    d_arr_3__3, d_arr_3__2, d_arr_3__1, d_arr_3__0, d_arr_4__31, 
                    d_arr_4__30, d_arr_4__29, d_arr_4__28, d_arr_4__27, 
                    d_arr_4__26, d_arr_4__25, d_arr_4__24, d_arr_4__23, 
                    d_arr_4__22, d_arr_4__21, d_arr_4__20, d_arr_4__19, 
                    d_arr_4__18, d_arr_4__17, d_arr_4__16, d_arr_4__15, 
                    d_arr_4__14, d_arr_4__13, d_arr_4__12, d_arr_4__11, 
                    d_arr_4__10, d_arr_4__9, d_arr_4__8, d_arr_4__7, d_arr_4__6, 
                    d_arr_4__5, d_arr_4__4, d_arr_4__3, d_arr_4__2, d_arr_4__1, 
                    d_arr_4__0, d_arr_5__31, d_arr_5__30, d_arr_5__29, 
                    d_arr_5__28, d_arr_5__27, d_arr_5__26, d_arr_5__25, 
                    d_arr_5__24, d_arr_5__23, d_arr_5__22, d_arr_5__21, 
                    d_arr_5__20, d_arr_5__19, d_arr_5__18, d_arr_5__17, 
                    d_arr_5__16, d_arr_5__15, d_arr_5__14, d_arr_5__13, 
                    d_arr_5__12, d_arr_5__11, d_arr_5__10, d_arr_5__9, 
                    d_arr_5__8, d_arr_5__7, d_arr_5__6, d_arr_5__5, d_arr_5__4, 
                    d_arr_5__3, d_arr_5__2, d_arr_5__1, d_arr_5__0, d_arr_6__31, 
                    d_arr_6__30, d_arr_6__29, d_arr_6__28, d_arr_6__27, 
                    d_arr_6__26, d_arr_6__25, d_arr_6__24, d_arr_6__23, 
                    d_arr_6__22, d_arr_6__21, d_arr_6__20, d_arr_6__19, 
                    d_arr_6__18, d_arr_6__17, d_arr_6__16, d_arr_6__15, 
                    d_arr_6__14, d_arr_6__13, d_arr_6__12, d_arr_6__11, 
                    d_arr_6__10, d_arr_6__9, d_arr_6__8, d_arr_6__7, d_arr_6__6, 
                    d_arr_6__5, d_arr_6__4, d_arr_6__3, d_arr_6__2, d_arr_6__1, 
                    d_arr_6__0, d_arr_7__31, d_arr_7__30, d_arr_7__29, 
                    d_arr_7__28, d_arr_7__27, d_arr_7__26, d_arr_7__25, 
                    d_arr_7__24, d_arr_7__23, d_arr_7__22, d_arr_7__21, 
                    d_arr_7__20, d_arr_7__19, d_arr_7__18, d_arr_7__17, 
                    d_arr_7__16, d_arr_7__15, d_arr_7__14, d_arr_7__13, 
                    d_arr_7__12, d_arr_7__11, d_arr_7__10, d_arr_7__9, 
                    d_arr_7__8, d_arr_7__7, d_arr_7__6, d_arr_7__5, d_arr_7__4, 
                    d_arr_7__3, d_arr_7__2, d_arr_7__1, d_arr_7__0, d_arr_8__31, 
                    d_arr_8__30, d_arr_8__29, d_arr_8__28, d_arr_8__27, 
                    d_arr_8__26, d_arr_8__25, d_arr_8__24, d_arr_8__23, 
                    d_arr_8__22, d_arr_8__21, d_arr_8__20, d_arr_8__19, 
                    d_arr_8__18, d_arr_8__17, d_arr_8__16, d_arr_8__15, 
                    d_arr_8__14, d_arr_8__13, d_arr_8__12, d_arr_8__11, 
                    d_arr_8__10, d_arr_8__9, d_arr_8__8, d_arr_8__7, d_arr_8__6, 
                    d_arr_8__5, d_arr_8__4, d_arr_8__3, d_arr_8__2, d_arr_8__1, 
                    d_arr_8__0, d_arr_9__31, d_arr_9__30, d_arr_9__29, 
                    d_arr_9__28, d_arr_9__27, d_arr_9__26, d_arr_9__25, 
                    d_arr_9__24, d_arr_9__23, d_arr_9__22, d_arr_9__21, 
                    d_arr_9__20, d_arr_9__19, d_arr_9__18, d_arr_9__17, 
                    d_arr_9__16, d_arr_9__15, d_arr_9__14, d_arr_9__13, 
                    d_arr_9__12, d_arr_9__11, d_arr_9__10, d_arr_9__9, 
                    d_arr_9__8, d_arr_9__7, d_arr_9__6, d_arr_9__5, d_arr_9__4, 
                    d_arr_9__3, d_arr_9__2, d_arr_9__1, d_arr_9__0, d_arr_10__31, 
                    d_arr_10__30, d_arr_10__29, d_arr_10__28, d_arr_10__27, 
                    d_arr_10__26, d_arr_10__25, d_arr_10__24, d_arr_10__23, 
                    d_arr_10__22, d_arr_10__21, d_arr_10__20, d_arr_10__19, 
                    d_arr_10__18, d_arr_10__17, d_arr_10__16, d_arr_10__15, 
                    d_arr_10__14, d_arr_10__13, d_arr_10__12, d_arr_10__11, 
                    d_arr_10__10, d_arr_10__9, d_arr_10__8, d_arr_10__7, 
                    d_arr_10__6, d_arr_10__5, d_arr_10__4, d_arr_10__3, 
                    d_arr_10__2, d_arr_10__1, d_arr_10__0, d_arr_11__31, 
                    d_arr_11__30, d_arr_11__29, d_arr_11__28, d_arr_11__27, 
                    d_arr_11__26, d_arr_11__25, d_arr_11__24, d_arr_11__23, 
                    d_arr_11__22, d_arr_11__21, d_arr_11__20, d_arr_11__19, 
                    d_arr_11__18, d_arr_11__17, d_arr_11__16, d_arr_11__15, 
                    d_arr_11__14, d_arr_11__13, d_arr_11__12, d_arr_11__11, 
                    d_arr_11__10, d_arr_11__9, d_arr_11__8, d_arr_11__7, 
                    d_arr_11__6, d_arr_11__5, d_arr_11__4, d_arr_11__3, 
                    d_arr_11__2, d_arr_11__1, d_arr_11__0, d_arr_12__31, 
                    d_arr_12__30, d_arr_12__29, d_arr_12__28, d_arr_12__27, 
                    d_arr_12__26, d_arr_12__25, d_arr_12__24, d_arr_12__23, 
                    d_arr_12__22, d_arr_12__21, d_arr_12__20, d_arr_12__19, 
                    d_arr_12__18, d_arr_12__17, d_arr_12__16, d_arr_12__15, 
                    d_arr_12__14, d_arr_12__13, d_arr_12__12, d_arr_12__11, 
                    d_arr_12__10, d_arr_12__9, d_arr_12__8, d_arr_12__7, 
                    d_arr_12__6, d_arr_12__5, d_arr_12__4, d_arr_12__3, 
                    d_arr_12__2, d_arr_12__1, d_arr_12__0, d_arr_13__31, 
                    d_arr_13__30, d_arr_13__29, d_arr_13__28, d_arr_13__27, 
                    d_arr_13__26, d_arr_13__25, d_arr_13__24, d_arr_13__23, 
                    d_arr_13__22, d_arr_13__21, d_arr_13__20, d_arr_13__19, 
                    d_arr_13__18, d_arr_13__17, d_arr_13__16, d_arr_13__15, 
                    d_arr_13__14, d_arr_13__13, d_arr_13__12, d_arr_13__11, 
                    d_arr_13__10, d_arr_13__9, d_arr_13__8, d_arr_13__7, 
                    d_arr_13__6, d_arr_13__5, d_arr_13__4, d_arr_13__3, 
                    d_arr_13__2, d_arr_13__1, d_arr_13__0, d_arr_14__31, 
                    d_arr_14__30, d_arr_14__29, d_arr_14__28, d_arr_14__27, 
                    d_arr_14__26, d_arr_14__25, d_arr_14__24, d_arr_14__23, 
                    d_arr_14__22, d_arr_14__21, d_arr_14__20, d_arr_14__19, 
                    d_arr_14__18, d_arr_14__17, d_arr_14__16, d_arr_14__15, 
                    d_arr_14__14, d_arr_14__13, d_arr_14__12, d_arr_14__11, 
                    d_arr_14__10, d_arr_14__9, d_arr_14__8, d_arr_14__7, 
                    d_arr_14__6, d_arr_14__5, d_arr_14__4, d_arr_14__3, 
                    d_arr_14__2, d_arr_14__1, d_arr_14__0, d_arr_15__31, 
                    d_arr_15__30, d_arr_15__29, d_arr_15__28, d_arr_15__27, 
                    d_arr_15__26, d_arr_15__25, d_arr_15__24, d_arr_15__23, 
                    d_arr_15__22, d_arr_15__21, d_arr_15__20, d_arr_15__19, 
                    d_arr_15__18, d_arr_15__17, d_arr_15__16, d_arr_15__15, 
                    d_arr_15__14, d_arr_15__13, d_arr_15__12, d_arr_15__11, 
                    d_arr_15__10, d_arr_15__9, d_arr_15__8, d_arr_15__7, 
                    d_arr_15__6, d_arr_15__5, d_arr_15__4, d_arr_15__3, 
                    d_arr_15__2, d_arr_15__1, d_arr_15__0, d_arr_16__31, 
                    d_arr_16__30, d_arr_16__29, d_arr_16__28, d_arr_16__27, 
                    d_arr_16__26, d_arr_16__25, d_arr_16__24, d_arr_16__23, 
                    d_arr_16__22, d_arr_16__21, d_arr_16__20, d_arr_16__19, 
                    d_arr_16__18, d_arr_16__17, d_arr_16__16, d_arr_16__15, 
                    d_arr_16__14, d_arr_16__13, d_arr_16__12, d_arr_16__11, 
                    d_arr_16__10, d_arr_16__9, d_arr_16__8, d_arr_16__7, 
                    d_arr_16__6, d_arr_16__5, d_arr_16__4, d_arr_16__3, 
                    d_arr_16__2, d_arr_16__1, d_arr_16__0, d_arr_17__31, 
                    d_arr_17__30, d_arr_17__29, d_arr_17__28, d_arr_17__27, 
                    d_arr_17__26, d_arr_17__25, d_arr_17__24, d_arr_17__23, 
                    d_arr_17__22, d_arr_17__21, d_arr_17__20, d_arr_17__19, 
                    d_arr_17__18, d_arr_17__17, d_arr_17__16, d_arr_17__15, 
                    d_arr_17__14, d_arr_17__13, d_arr_17__12, d_arr_17__11, 
                    d_arr_17__10, d_arr_17__9, d_arr_17__8, d_arr_17__7, 
                    d_arr_17__6, d_arr_17__5, d_arr_17__4, d_arr_17__3, 
                    d_arr_17__2, d_arr_17__1, d_arr_17__0, d_arr_18__31, 
                    d_arr_18__30, d_arr_18__29, d_arr_18__28, d_arr_18__27, 
                    d_arr_18__26, d_arr_18__25, d_arr_18__24, d_arr_18__23, 
                    d_arr_18__22, d_arr_18__21, d_arr_18__20, d_arr_18__19, 
                    d_arr_18__18, d_arr_18__17, d_arr_18__16, d_arr_18__15, 
                    d_arr_18__14, d_arr_18__13, d_arr_18__12, d_arr_18__11, 
                    d_arr_18__10, d_arr_18__9, d_arr_18__8, d_arr_18__7, 
                    d_arr_18__6, d_arr_18__5, d_arr_18__4, d_arr_18__3, 
                    d_arr_18__2, d_arr_18__1, d_arr_18__0, d_arr_19__31, 
                    d_arr_19__30, d_arr_19__29, d_arr_19__28, d_arr_19__27, 
                    d_arr_19__26, d_arr_19__25, d_arr_19__24, d_arr_19__23, 
                    d_arr_19__22, d_arr_19__21, d_arr_19__20, d_arr_19__19, 
                    d_arr_19__18, d_arr_19__17, d_arr_19__16, d_arr_19__15, 
                    d_arr_19__14, d_arr_19__13, d_arr_19__12, d_arr_19__11, 
                    d_arr_19__10, d_arr_19__9, d_arr_19__8, d_arr_19__7, 
                    d_arr_19__6, d_arr_19__5, d_arr_19__4, d_arr_19__3, 
                    d_arr_19__2, d_arr_19__1, d_arr_19__0, d_arr_20__31, 
                    d_arr_20__30, d_arr_20__29, d_arr_20__28, d_arr_20__27, 
                    d_arr_20__26, d_arr_20__25, d_arr_20__24, d_arr_20__23, 
                    d_arr_20__22, d_arr_20__21, d_arr_20__20, d_arr_20__19, 
                    d_arr_20__18, d_arr_20__17, d_arr_20__16, d_arr_20__15, 
                    d_arr_20__14, d_arr_20__13, d_arr_20__12, d_arr_20__11, 
                    d_arr_20__10, d_arr_20__9, d_arr_20__8, d_arr_20__7, 
                    d_arr_20__6, d_arr_20__5, d_arr_20__4, d_arr_20__3, 
                    d_arr_20__2, d_arr_20__1, d_arr_20__0, d_arr_21__31, 
                    d_arr_21__30, d_arr_21__29, d_arr_21__28, d_arr_21__27, 
                    d_arr_21__26, d_arr_21__25, d_arr_21__24, d_arr_21__23, 
                    d_arr_21__22, d_arr_21__21, d_arr_21__20, d_arr_21__19, 
                    d_arr_21__18, d_arr_21__17, d_arr_21__16, d_arr_21__15, 
                    d_arr_21__14, d_arr_21__13, d_arr_21__12, d_arr_21__11, 
                    d_arr_21__10, d_arr_21__9, d_arr_21__8, d_arr_21__7, 
                    d_arr_21__6, d_arr_21__5, d_arr_21__4, d_arr_21__3, 
                    d_arr_21__2, d_arr_21__1, d_arr_21__0, d_arr_22__31, 
                    d_arr_22__30, d_arr_22__29, d_arr_22__28, d_arr_22__27, 
                    d_arr_22__26, d_arr_22__25, d_arr_22__24, d_arr_22__23, 
                    d_arr_22__22, d_arr_22__21, d_arr_22__20, d_arr_22__19, 
                    d_arr_22__18, d_arr_22__17, d_arr_22__16, d_arr_22__15, 
                    d_arr_22__14, d_arr_22__13, d_arr_22__12, d_arr_22__11, 
                    d_arr_22__10, d_arr_22__9, d_arr_22__8, d_arr_22__7, 
                    d_arr_22__6, d_arr_22__5, d_arr_22__4, d_arr_22__3, 
                    d_arr_22__2, d_arr_22__1, d_arr_22__0, d_arr_23__31, 
                    d_arr_23__30, d_arr_23__29, d_arr_23__28, d_arr_23__27, 
                    d_arr_23__26, d_arr_23__25, d_arr_23__24, d_arr_23__23, 
                    d_arr_23__22, d_arr_23__21, d_arr_23__20, d_arr_23__19, 
                    d_arr_23__18, d_arr_23__17, d_arr_23__16, d_arr_23__15, 
                    d_arr_23__14, d_arr_23__13, d_arr_23__12, d_arr_23__11, 
                    d_arr_23__10, d_arr_23__9, d_arr_23__8, d_arr_23__7, 
                    d_arr_23__6, d_arr_23__5, d_arr_23__4, d_arr_23__3, 
                    d_arr_23__2, d_arr_23__1, d_arr_23__0, d_arr_24__31, 
                    d_arr_24__30, d_arr_24__29, d_arr_24__28, d_arr_24__27, 
                    d_arr_24__26, d_arr_24__25, d_arr_24__24, d_arr_24__23, 
                    d_arr_24__22, d_arr_24__21, d_arr_24__20, d_arr_24__19, 
                    d_arr_24__18, d_arr_24__17, d_arr_24__16, d_arr_24__15, 
                    d_arr_24__14, d_arr_24__13, d_arr_24__12, d_arr_24__11, 
                    d_arr_24__10, d_arr_24__9, d_arr_24__8, d_arr_24__7, 
                    d_arr_24__6, d_arr_24__5, d_arr_24__4, d_arr_24__3, 
                    d_arr_24__2, d_arr_24__1, d_arr_24__0 ) ;

    input d_arr_mux_0__31 ;
    input d_arr_mux_0__30 ;
    input d_arr_mux_0__29 ;
    input d_arr_mux_0__28 ;
    input d_arr_mux_0__27 ;
    input d_arr_mux_0__26 ;
    input d_arr_mux_0__25 ;
    input d_arr_mux_0__24 ;
    input d_arr_mux_0__23 ;
    input d_arr_mux_0__22 ;
    input d_arr_mux_0__21 ;
    input d_arr_mux_0__20 ;
    input d_arr_mux_0__19 ;
    input d_arr_mux_0__18 ;
    input d_arr_mux_0__17 ;
    input d_arr_mux_0__16 ;
    input d_arr_mux_0__15 ;
    input d_arr_mux_0__14 ;
    input d_arr_mux_0__13 ;
    input d_arr_mux_0__12 ;
    input d_arr_mux_0__11 ;
    input d_arr_mux_0__10 ;
    input d_arr_mux_0__9 ;
    input d_arr_mux_0__8 ;
    input d_arr_mux_0__7 ;
    input d_arr_mux_0__6 ;
    input d_arr_mux_0__5 ;
    input d_arr_mux_0__4 ;
    input d_arr_mux_0__3 ;
    input d_arr_mux_0__2 ;
    input d_arr_mux_0__1 ;
    input d_arr_mux_0__0 ;
    input d_arr_mux_1__31 ;
    input d_arr_mux_1__30 ;
    input d_arr_mux_1__29 ;
    input d_arr_mux_1__28 ;
    input d_arr_mux_1__27 ;
    input d_arr_mux_1__26 ;
    input d_arr_mux_1__25 ;
    input d_arr_mux_1__24 ;
    input d_arr_mux_1__23 ;
    input d_arr_mux_1__22 ;
    input d_arr_mux_1__21 ;
    input d_arr_mux_1__20 ;
    input d_arr_mux_1__19 ;
    input d_arr_mux_1__18 ;
    input d_arr_mux_1__17 ;
    input d_arr_mux_1__16 ;
    input d_arr_mux_1__15 ;
    input d_arr_mux_1__14 ;
    input d_arr_mux_1__13 ;
    input d_arr_mux_1__12 ;
    input d_arr_mux_1__11 ;
    input d_arr_mux_1__10 ;
    input d_arr_mux_1__9 ;
    input d_arr_mux_1__8 ;
    input d_arr_mux_1__7 ;
    input d_arr_mux_1__6 ;
    input d_arr_mux_1__5 ;
    input d_arr_mux_1__4 ;
    input d_arr_mux_1__3 ;
    input d_arr_mux_1__2 ;
    input d_arr_mux_1__1 ;
    input d_arr_mux_1__0 ;
    input d_arr_mux_2__31 ;
    input d_arr_mux_2__30 ;
    input d_arr_mux_2__29 ;
    input d_arr_mux_2__28 ;
    input d_arr_mux_2__27 ;
    input d_arr_mux_2__26 ;
    input d_arr_mux_2__25 ;
    input d_arr_mux_2__24 ;
    input d_arr_mux_2__23 ;
    input d_arr_mux_2__22 ;
    input d_arr_mux_2__21 ;
    input d_arr_mux_2__20 ;
    input d_arr_mux_2__19 ;
    input d_arr_mux_2__18 ;
    input d_arr_mux_2__17 ;
    input d_arr_mux_2__16 ;
    input d_arr_mux_2__15 ;
    input d_arr_mux_2__14 ;
    input d_arr_mux_2__13 ;
    input d_arr_mux_2__12 ;
    input d_arr_mux_2__11 ;
    input d_arr_mux_2__10 ;
    input d_arr_mux_2__9 ;
    input d_arr_mux_2__8 ;
    input d_arr_mux_2__7 ;
    input d_arr_mux_2__6 ;
    input d_arr_mux_2__5 ;
    input d_arr_mux_2__4 ;
    input d_arr_mux_2__3 ;
    input d_arr_mux_2__2 ;
    input d_arr_mux_2__1 ;
    input d_arr_mux_2__0 ;
    input d_arr_mux_3__31 ;
    input d_arr_mux_3__30 ;
    input d_arr_mux_3__29 ;
    input d_arr_mux_3__28 ;
    input d_arr_mux_3__27 ;
    input d_arr_mux_3__26 ;
    input d_arr_mux_3__25 ;
    input d_arr_mux_3__24 ;
    input d_arr_mux_3__23 ;
    input d_arr_mux_3__22 ;
    input d_arr_mux_3__21 ;
    input d_arr_mux_3__20 ;
    input d_arr_mux_3__19 ;
    input d_arr_mux_3__18 ;
    input d_arr_mux_3__17 ;
    input d_arr_mux_3__16 ;
    input d_arr_mux_3__15 ;
    input d_arr_mux_3__14 ;
    input d_arr_mux_3__13 ;
    input d_arr_mux_3__12 ;
    input d_arr_mux_3__11 ;
    input d_arr_mux_3__10 ;
    input d_arr_mux_3__9 ;
    input d_arr_mux_3__8 ;
    input d_arr_mux_3__7 ;
    input d_arr_mux_3__6 ;
    input d_arr_mux_3__5 ;
    input d_arr_mux_3__4 ;
    input d_arr_mux_3__3 ;
    input d_arr_mux_3__2 ;
    input d_arr_mux_3__1 ;
    input d_arr_mux_3__0 ;
    input d_arr_mux_4__31 ;
    input d_arr_mux_4__30 ;
    input d_arr_mux_4__29 ;
    input d_arr_mux_4__28 ;
    input d_arr_mux_4__27 ;
    input d_arr_mux_4__26 ;
    input d_arr_mux_4__25 ;
    input d_arr_mux_4__24 ;
    input d_arr_mux_4__23 ;
    input d_arr_mux_4__22 ;
    input d_arr_mux_4__21 ;
    input d_arr_mux_4__20 ;
    input d_arr_mux_4__19 ;
    input d_arr_mux_4__18 ;
    input d_arr_mux_4__17 ;
    input d_arr_mux_4__16 ;
    input d_arr_mux_4__15 ;
    input d_arr_mux_4__14 ;
    input d_arr_mux_4__13 ;
    input d_arr_mux_4__12 ;
    input d_arr_mux_4__11 ;
    input d_arr_mux_4__10 ;
    input d_arr_mux_4__9 ;
    input d_arr_mux_4__8 ;
    input d_arr_mux_4__7 ;
    input d_arr_mux_4__6 ;
    input d_arr_mux_4__5 ;
    input d_arr_mux_4__4 ;
    input d_arr_mux_4__3 ;
    input d_arr_mux_4__2 ;
    input d_arr_mux_4__1 ;
    input d_arr_mux_4__0 ;
    input d_arr_mux_5__31 ;
    input d_arr_mux_5__30 ;
    input d_arr_mux_5__29 ;
    input d_arr_mux_5__28 ;
    input d_arr_mux_5__27 ;
    input d_arr_mux_5__26 ;
    input d_arr_mux_5__25 ;
    input d_arr_mux_5__24 ;
    input d_arr_mux_5__23 ;
    input d_arr_mux_5__22 ;
    input d_arr_mux_5__21 ;
    input d_arr_mux_5__20 ;
    input d_arr_mux_5__19 ;
    input d_arr_mux_5__18 ;
    input d_arr_mux_5__17 ;
    input d_arr_mux_5__16 ;
    input d_arr_mux_5__15 ;
    input d_arr_mux_5__14 ;
    input d_arr_mux_5__13 ;
    input d_arr_mux_5__12 ;
    input d_arr_mux_5__11 ;
    input d_arr_mux_5__10 ;
    input d_arr_mux_5__9 ;
    input d_arr_mux_5__8 ;
    input d_arr_mux_5__7 ;
    input d_arr_mux_5__6 ;
    input d_arr_mux_5__5 ;
    input d_arr_mux_5__4 ;
    input d_arr_mux_5__3 ;
    input d_arr_mux_5__2 ;
    input d_arr_mux_5__1 ;
    input d_arr_mux_5__0 ;
    input d_arr_mux_6__31 ;
    input d_arr_mux_6__30 ;
    input d_arr_mux_6__29 ;
    input d_arr_mux_6__28 ;
    input d_arr_mux_6__27 ;
    input d_arr_mux_6__26 ;
    input d_arr_mux_6__25 ;
    input d_arr_mux_6__24 ;
    input d_arr_mux_6__23 ;
    input d_arr_mux_6__22 ;
    input d_arr_mux_6__21 ;
    input d_arr_mux_6__20 ;
    input d_arr_mux_6__19 ;
    input d_arr_mux_6__18 ;
    input d_arr_mux_6__17 ;
    input d_arr_mux_6__16 ;
    input d_arr_mux_6__15 ;
    input d_arr_mux_6__14 ;
    input d_arr_mux_6__13 ;
    input d_arr_mux_6__12 ;
    input d_arr_mux_6__11 ;
    input d_arr_mux_6__10 ;
    input d_arr_mux_6__9 ;
    input d_arr_mux_6__8 ;
    input d_arr_mux_6__7 ;
    input d_arr_mux_6__6 ;
    input d_arr_mux_6__5 ;
    input d_arr_mux_6__4 ;
    input d_arr_mux_6__3 ;
    input d_arr_mux_6__2 ;
    input d_arr_mux_6__1 ;
    input d_arr_mux_6__0 ;
    input d_arr_mux_7__31 ;
    input d_arr_mux_7__30 ;
    input d_arr_mux_7__29 ;
    input d_arr_mux_7__28 ;
    input d_arr_mux_7__27 ;
    input d_arr_mux_7__26 ;
    input d_arr_mux_7__25 ;
    input d_arr_mux_7__24 ;
    input d_arr_mux_7__23 ;
    input d_arr_mux_7__22 ;
    input d_arr_mux_7__21 ;
    input d_arr_mux_7__20 ;
    input d_arr_mux_7__19 ;
    input d_arr_mux_7__18 ;
    input d_arr_mux_7__17 ;
    input d_arr_mux_7__16 ;
    input d_arr_mux_7__15 ;
    input d_arr_mux_7__14 ;
    input d_arr_mux_7__13 ;
    input d_arr_mux_7__12 ;
    input d_arr_mux_7__11 ;
    input d_arr_mux_7__10 ;
    input d_arr_mux_7__9 ;
    input d_arr_mux_7__8 ;
    input d_arr_mux_7__7 ;
    input d_arr_mux_7__6 ;
    input d_arr_mux_7__5 ;
    input d_arr_mux_7__4 ;
    input d_arr_mux_7__3 ;
    input d_arr_mux_7__2 ;
    input d_arr_mux_7__1 ;
    input d_arr_mux_7__0 ;
    input d_arr_mux_8__31 ;
    input d_arr_mux_8__30 ;
    input d_arr_mux_8__29 ;
    input d_arr_mux_8__28 ;
    input d_arr_mux_8__27 ;
    input d_arr_mux_8__26 ;
    input d_arr_mux_8__25 ;
    input d_arr_mux_8__24 ;
    input d_arr_mux_8__23 ;
    input d_arr_mux_8__22 ;
    input d_arr_mux_8__21 ;
    input d_arr_mux_8__20 ;
    input d_arr_mux_8__19 ;
    input d_arr_mux_8__18 ;
    input d_arr_mux_8__17 ;
    input d_arr_mux_8__16 ;
    input d_arr_mux_8__15 ;
    input d_arr_mux_8__14 ;
    input d_arr_mux_8__13 ;
    input d_arr_mux_8__12 ;
    input d_arr_mux_8__11 ;
    input d_arr_mux_8__10 ;
    input d_arr_mux_8__9 ;
    input d_arr_mux_8__8 ;
    input d_arr_mux_8__7 ;
    input d_arr_mux_8__6 ;
    input d_arr_mux_8__5 ;
    input d_arr_mux_8__4 ;
    input d_arr_mux_8__3 ;
    input d_arr_mux_8__2 ;
    input d_arr_mux_8__1 ;
    input d_arr_mux_8__0 ;
    input d_arr_mux_9__31 ;
    input d_arr_mux_9__30 ;
    input d_arr_mux_9__29 ;
    input d_arr_mux_9__28 ;
    input d_arr_mux_9__27 ;
    input d_arr_mux_9__26 ;
    input d_arr_mux_9__25 ;
    input d_arr_mux_9__24 ;
    input d_arr_mux_9__23 ;
    input d_arr_mux_9__22 ;
    input d_arr_mux_9__21 ;
    input d_arr_mux_9__20 ;
    input d_arr_mux_9__19 ;
    input d_arr_mux_9__18 ;
    input d_arr_mux_9__17 ;
    input d_arr_mux_9__16 ;
    input d_arr_mux_9__15 ;
    input d_arr_mux_9__14 ;
    input d_arr_mux_9__13 ;
    input d_arr_mux_9__12 ;
    input d_arr_mux_9__11 ;
    input d_arr_mux_9__10 ;
    input d_arr_mux_9__9 ;
    input d_arr_mux_9__8 ;
    input d_arr_mux_9__7 ;
    input d_arr_mux_9__6 ;
    input d_arr_mux_9__5 ;
    input d_arr_mux_9__4 ;
    input d_arr_mux_9__3 ;
    input d_arr_mux_9__2 ;
    input d_arr_mux_9__1 ;
    input d_arr_mux_9__0 ;
    input d_arr_mux_10__31 ;
    input d_arr_mux_10__30 ;
    input d_arr_mux_10__29 ;
    input d_arr_mux_10__28 ;
    input d_arr_mux_10__27 ;
    input d_arr_mux_10__26 ;
    input d_arr_mux_10__25 ;
    input d_arr_mux_10__24 ;
    input d_arr_mux_10__23 ;
    input d_arr_mux_10__22 ;
    input d_arr_mux_10__21 ;
    input d_arr_mux_10__20 ;
    input d_arr_mux_10__19 ;
    input d_arr_mux_10__18 ;
    input d_arr_mux_10__17 ;
    input d_arr_mux_10__16 ;
    input d_arr_mux_10__15 ;
    input d_arr_mux_10__14 ;
    input d_arr_mux_10__13 ;
    input d_arr_mux_10__12 ;
    input d_arr_mux_10__11 ;
    input d_arr_mux_10__10 ;
    input d_arr_mux_10__9 ;
    input d_arr_mux_10__8 ;
    input d_arr_mux_10__7 ;
    input d_arr_mux_10__6 ;
    input d_arr_mux_10__5 ;
    input d_arr_mux_10__4 ;
    input d_arr_mux_10__3 ;
    input d_arr_mux_10__2 ;
    input d_arr_mux_10__1 ;
    input d_arr_mux_10__0 ;
    input d_arr_mux_11__31 ;
    input d_arr_mux_11__30 ;
    input d_arr_mux_11__29 ;
    input d_arr_mux_11__28 ;
    input d_arr_mux_11__27 ;
    input d_arr_mux_11__26 ;
    input d_arr_mux_11__25 ;
    input d_arr_mux_11__24 ;
    input d_arr_mux_11__23 ;
    input d_arr_mux_11__22 ;
    input d_arr_mux_11__21 ;
    input d_arr_mux_11__20 ;
    input d_arr_mux_11__19 ;
    input d_arr_mux_11__18 ;
    input d_arr_mux_11__17 ;
    input d_arr_mux_11__16 ;
    input d_arr_mux_11__15 ;
    input d_arr_mux_11__14 ;
    input d_arr_mux_11__13 ;
    input d_arr_mux_11__12 ;
    input d_arr_mux_11__11 ;
    input d_arr_mux_11__10 ;
    input d_arr_mux_11__9 ;
    input d_arr_mux_11__8 ;
    input d_arr_mux_11__7 ;
    input d_arr_mux_11__6 ;
    input d_arr_mux_11__5 ;
    input d_arr_mux_11__4 ;
    input d_arr_mux_11__3 ;
    input d_arr_mux_11__2 ;
    input d_arr_mux_11__1 ;
    input d_arr_mux_11__0 ;
    input d_arr_mux_12__31 ;
    input d_arr_mux_12__30 ;
    input d_arr_mux_12__29 ;
    input d_arr_mux_12__28 ;
    input d_arr_mux_12__27 ;
    input d_arr_mux_12__26 ;
    input d_arr_mux_12__25 ;
    input d_arr_mux_12__24 ;
    input d_arr_mux_12__23 ;
    input d_arr_mux_12__22 ;
    input d_arr_mux_12__21 ;
    input d_arr_mux_12__20 ;
    input d_arr_mux_12__19 ;
    input d_arr_mux_12__18 ;
    input d_arr_mux_12__17 ;
    input d_arr_mux_12__16 ;
    input d_arr_mux_12__15 ;
    input d_arr_mux_12__14 ;
    input d_arr_mux_12__13 ;
    input d_arr_mux_12__12 ;
    input d_arr_mux_12__11 ;
    input d_arr_mux_12__10 ;
    input d_arr_mux_12__9 ;
    input d_arr_mux_12__8 ;
    input d_arr_mux_12__7 ;
    input d_arr_mux_12__6 ;
    input d_arr_mux_12__5 ;
    input d_arr_mux_12__4 ;
    input d_arr_mux_12__3 ;
    input d_arr_mux_12__2 ;
    input d_arr_mux_12__1 ;
    input d_arr_mux_12__0 ;
    input d_arr_mux_13__31 ;
    input d_arr_mux_13__30 ;
    input d_arr_mux_13__29 ;
    input d_arr_mux_13__28 ;
    input d_arr_mux_13__27 ;
    input d_arr_mux_13__26 ;
    input d_arr_mux_13__25 ;
    input d_arr_mux_13__24 ;
    input d_arr_mux_13__23 ;
    input d_arr_mux_13__22 ;
    input d_arr_mux_13__21 ;
    input d_arr_mux_13__20 ;
    input d_arr_mux_13__19 ;
    input d_arr_mux_13__18 ;
    input d_arr_mux_13__17 ;
    input d_arr_mux_13__16 ;
    input d_arr_mux_13__15 ;
    input d_arr_mux_13__14 ;
    input d_arr_mux_13__13 ;
    input d_arr_mux_13__12 ;
    input d_arr_mux_13__11 ;
    input d_arr_mux_13__10 ;
    input d_arr_mux_13__9 ;
    input d_arr_mux_13__8 ;
    input d_arr_mux_13__7 ;
    input d_arr_mux_13__6 ;
    input d_arr_mux_13__5 ;
    input d_arr_mux_13__4 ;
    input d_arr_mux_13__3 ;
    input d_arr_mux_13__2 ;
    input d_arr_mux_13__1 ;
    input d_arr_mux_13__0 ;
    input d_arr_mux_14__31 ;
    input d_arr_mux_14__30 ;
    input d_arr_mux_14__29 ;
    input d_arr_mux_14__28 ;
    input d_arr_mux_14__27 ;
    input d_arr_mux_14__26 ;
    input d_arr_mux_14__25 ;
    input d_arr_mux_14__24 ;
    input d_arr_mux_14__23 ;
    input d_arr_mux_14__22 ;
    input d_arr_mux_14__21 ;
    input d_arr_mux_14__20 ;
    input d_arr_mux_14__19 ;
    input d_arr_mux_14__18 ;
    input d_arr_mux_14__17 ;
    input d_arr_mux_14__16 ;
    input d_arr_mux_14__15 ;
    input d_arr_mux_14__14 ;
    input d_arr_mux_14__13 ;
    input d_arr_mux_14__12 ;
    input d_arr_mux_14__11 ;
    input d_arr_mux_14__10 ;
    input d_arr_mux_14__9 ;
    input d_arr_mux_14__8 ;
    input d_arr_mux_14__7 ;
    input d_arr_mux_14__6 ;
    input d_arr_mux_14__5 ;
    input d_arr_mux_14__4 ;
    input d_arr_mux_14__3 ;
    input d_arr_mux_14__2 ;
    input d_arr_mux_14__1 ;
    input d_arr_mux_14__0 ;
    input d_arr_mux_15__31 ;
    input d_arr_mux_15__30 ;
    input d_arr_mux_15__29 ;
    input d_arr_mux_15__28 ;
    input d_arr_mux_15__27 ;
    input d_arr_mux_15__26 ;
    input d_arr_mux_15__25 ;
    input d_arr_mux_15__24 ;
    input d_arr_mux_15__23 ;
    input d_arr_mux_15__22 ;
    input d_arr_mux_15__21 ;
    input d_arr_mux_15__20 ;
    input d_arr_mux_15__19 ;
    input d_arr_mux_15__18 ;
    input d_arr_mux_15__17 ;
    input d_arr_mux_15__16 ;
    input d_arr_mux_15__15 ;
    input d_arr_mux_15__14 ;
    input d_arr_mux_15__13 ;
    input d_arr_mux_15__12 ;
    input d_arr_mux_15__11 ;
    input d_arr_mux_15__10 ;
    input d_arr_mux_15__9 ;
    input d_arr_mux_15__8 ;
    input d_arr_mux_15__7 ;
    input d_arr_mux_15__6 ;
    input d_arr_mux_15__5 ;
    input d_arr_mux_15__4 ;
    input d_arr_mux_15__3 ;
    input d_arr_mux_15__2 ;
    input d_arr_mux_15__1 ;
    input d_arr_mux_15__0 ;
    input d_arr_mux_16__31 ;
    input d_arr_mux_16__30 ;
    input d_arr_mux_16__29 ;
    input d_arr_mux_16__28 ;
    input d_arr_mux_16__27 ;
    input d_arr_mux_16__26 ;
    input d_arr_mux_16__25 ;
    input d_arr_mux_16__24 ;
    input d_arr_mux_16__23 ;
    input d_arr_mux_16__22 ;
    input d_arr_mux_16__21 ;
    input d_arr_mux_16__20 ;
    input d_arr_mux_16__19 ;
    input d_arr_mux_16__18 ;
    input d_arr_mux_16__17 ;
    input d_arr_mux_16__16 ;
    input d_arr_mux_16__15 ;
    input d_arr_mux_16__14 ;
    input d_arr_mux_16__13 ;
    input d_arr_mux_16__12 ;
    input d_arr_mux_16__11 ;
    input d_arr_mux_16__10 ;
    input d_arr_mux_16__9 ;
    input d_arr_mux_16__8 ;
    input d_arr_mux_16__7 ;
    input d_arr_mux_16__6 ;
    input d_arr_mux_16__5 ;
    input d_arr_mux_16__4 ;
    input d_arr_mux_16__3 ;
    input d_arr_mux_16__2 ;
    input d_arr_mux_16__1 ;
    input d_arr_mux_16__0 ;
    input d_arr_mux_17__31 ;
    input d_arr_mux_17__30 ;
    input d_arr_mux_17__29 ;
    input d_arr_mux_17__28 ;
    input d_arr_mux_17__27 ;
    input d_arr_mux_17__26 ;
    input d_arr_mux_17__25 ;
    input d_arr_mux_17__24 ;
    input d_arr_mux_17__23 ;
    input d_arr_mux_17__22 ;
    input d_arr_mux_17__21 ;
    input d_arr_mux_17__20 ;
    input d_arr_mux_17__19 ;
    input d_arr_mux_17__18 ;
    input d_arr_mux_17__17 ;
    input d_arr_mux_17__16 ;
    input d_arr_mux_17__15 ;
    input d_arr_mux_17__14 ;
    input d_arr_mux_17__13 ;
    input d_arr_mux_17__12 ;
    input d_arr_mux_17__11 ;
    input d_arr_mux_17__10 ;
    input d_arr_mux_17__9 ;
    input d_arr_mux_17__8 ;
    input d_arr_mux_17__7 ;
    input d_arr_mux_17__6 ;
    input d_arr_mux_17__5 ;
    input d_arr_mux_17__4 ;
    input d_arr_mux_17__3 ;
    input d_arr_mux_17__2 ;
    input d_arr_mux_17__1 ;
    input d_arr_mux_17__0 ;
    input d_arr_mux_18__31 ;
    input d_arr_mux_18__30 ;
    input d_arr_mux_18__29 ;
    input d_arr_mux_18__28 ;
    input d_arr_mux_18__27 ;
    input d_arr_mux_18__26 ;
    input d_arr_mux_18__25 ;
    input d_arr_mux_18__24 ;
    input d_arr_mux_18__23 ;
    input d_arr_mux_18__22 ;
    input d_arr_mux_18__21 ;
    input d_arr_mux_18__20 ;
    input d_arr_mux_18__19 ;
    input d_arr_mux_18__18 ;
    input d_arr_mux_18__17 ;
    input d_arr_mux_18__16 ;
    input d_arr_mux_18__15 ;
    input d_arr_mux_18__14 ;
    input d_arr_mux_18__13 ;
    input d_arr_mux_18__12 ;
    input d_arr_mux_18__11 ;
    input d_arr_mux_18__10 ;
    input d_arr_mux_18__9 ;
    input d_arr_mux_18__8 ;
    input d_arr_mux_18__7 ;
    input d_arr_mux_18__6 ;
    input d_arr_mux_18__5 ;
    input d_arr_mux_18__4 ;
    input d_arr_mux_18__3 ;
    input d_arr_mux_18__2 ;
    input d_arr_mux_18__1 ;
    input d_arr_mux_18__0 ;
    input d_arr_mux_19__31 ;
    input d_arr_mux_19__30 ;
    input d_arr_mux_19__29 ;
    input d_arr_mux_19__28 ;
    input d_arr_mux_19__27 ;
    input d_arr_mux_19__26 ;
    input d_arr_mux_19__25 ;
    input d_arr_mux_19__24 ;
    input d_arr_mux_19__23 ;
    input d_arr_mux_19__22 ;
    input d_arr_mux_19__21 ;
    input d_arr_mux_19__20 ;
    input d_arr_mux_19__19 ;
    input d_arr_mux_19__18 ;
    input d_arr_mux_19__17 ;
    input d_arr_mux_19__16 ;
    input d_arr_mux_19__15 ;
    input d_arr_mux_19__14 ;
    input d_arr_mux_19__13 ;
    input d_arr_mux_19__12 ;
    input d_arr_mux_19__11 ;
    input d_arr_mux_19__10 ;
    input d_arr_mux_19__9 ;
    input d_arr_mux_19__8 ;
    input d_arr_mux_19__7 ;
    input d_arr_mux_19__6 ;
    input d_arr_mux_19__5 ;
    input d_arr_mux_19__4 ;
    input d_arr_mux_19__3 ;
    input d_arr_mux_19__2 ;
    input d_arr_mux_19__1 ;
    input d_arr_mux_19__0 ;
    input d_arr_mux_20__31 ;
    input d_arr_mux_20__30 ;
    input d_arr_mux_20__29 ;
    input d_arr_mux_20__28 ;
    input d_arr_mux_20__27 ;
    input d_arr_mux_20__26 ;
    input d_arr_mux_20__25 ;
    input d_arr_mux_20__24 ;
    input d_arr_mux_20__23 ;
    input d_arr_mux_20__22 ;
    input d_arr_mux_20__21 ;
    input d_arr_mux_20__20 ;
    input d_arr_mux_20__19 ;
    input d_arr_mux_20__18 ;
    input d_arr_mux_20__17 ;
    input d_arr_mux_20__16 ;
    input d_arr_mux_20__15 ;
    input d_arr_mux_20__14 ;
    input d_arr_mux_20__13 ;
    input d_arr_mux_20__12 ;
    input d_arr_mux_20__11 ;
    input d_arr_mux_20__10 ;
    input d_arr_mux_20__9 ;
    input d_arr_mux_20__8 ;
    input d_arr_mux_20__7 ;
    input d_arr_mux_20__6 ;
    input d_arr_mux_20__5 ;
    input d_arr_mux_20__4 ;
    input d_arr_mux_20__3 ;
    input d_arr_mux_20__2 ;
    input d_arr_mux_20__1 ;
    input d_arr_mux_20__0 ;
    input d_arr_mux_21__31 ;
    input d_arr_mux_21__30 ;
    input d_arr_mux_21__29 ;
    input d_arr_mux_21__28 ;
    input d_arr_mux_21__27 ;
    input d_arr_mux_21__26 ;
    input d_arr_mux_21__25 ;
    input d_arr_mux_21__24 ;
    input d_arr_mux_21__23 ;
    input d_arr_mux_21__22 ;
    input d_arr_mux_21__21 ;
    input d_arr_mux_21__20 ;
    input d_arr_mux_21__19 ;
    input d_arr_mux_21__18 ;
    input d_arr_mux_21__17 ;
    input d_arr_mux_21__16 ;
    input d_arr_mux_21__15 ;
    input d_arr_mux_21__14 ;
    input d_arr_mux_21__13 ;
    input d_arr_mux_21__12 ;
    input d_arr_mux_21__11 ;
    input d_arr_mux_21__10 ;
    input d_arr_mux_21__9 ;
    input d_arr_mux_21__8 ;
    input d_arr_mux_21__7 ;
    input d_arr_mux_21__6 ;
    input d_arr_mux_21__5 ;
    input d_arr_mux_21__4 ;
    input d_arr_mux_21__3 ;
    input d_arr_mux_21__2 ;
    input d_arr_mux_21__1 ;
    input d_arr_mux_21__0 ;
    input d_arr_mux_22__31 ;
    input d_arr_mux_22__30 ;
    input d_arr_mux_22__29 ;
    input d_arr_mux_22__28 ;
    input d_arr_mux_22__27 ;
    input d_arr_mux_22__26 ;
    input d_arr_mux_22__25 ;
    input d_arr_mux_22__24 ;
    input d_arr_mux_22__23 ;
    input d_arr_mux_22__22 ;
    input d_arr_mux_22__21 ;
    input d_arr_mux_22__20 ;
    input d_arr_mux_22__19 ;
    input d_arr_mux_22__18 ;
    input d_arr_mux_22__17 ;
    input d_arr_mux_22__16 ;
    input d_arr_mux_22__15 ;
    input d_arr_mux_22__14 ;
    input d_arr_mux_22__13 ;
    input d_arr_mux_22__12 ;
    input d_arr_mux_22__11 ;
    input d_arr_mux_22__10 ;
    input d_arr_mux_22__9 ;
    input d_arr_mux_22__8 ;
    input d_arr_mux_22__7 ;
    input d_arr_mux_22__6 ;
    input d_arr_mux_22__5 ;
    input d_arr_mux_22__4 ;
    input d_arr_mux_22__3 ;
    input d_arr_mux_22__2 ;
    input d_arr_mux_22__1 ;
    input d_arr_mux_22__0 ;
    input d_arr_mux_23__31 ;
    input d_arr_mux_23__30 ;
    input d_arr_mux_23__29 ;
    input d_arr_mux_23__28 ;
    input d_arr_mux_23__27 ;
    input d_arr_mux_23__26 ;
    input d_arr_mux_23__25 ;
    input d_arr_mux_23__24 ;
    input d_arr_mux_23__23 ;
    input d_arr_mux_23__22 ;
    input d_arr_mux_23__21 ;
    input d_arr_mux_23__20 ;
    input d_arr_mux_23__19 ;
    input d_arr_mux_23__18 ;
    input d_arr_mux_23__17 ;
    input d_arr_mux_23__16 ;
    input d_arr_mux_23__15 ;
    input d_arr_mux_23__14 ;
    input d_arr_mux_23__13 ;
    input d_arr_mux_23__12 ;
    input d_arr_mux_23__11 ;
    input d_arr_mux_23__10 ;
    input d_arr_mux_23__9 ;
    input d_arr_mux_23__8 ;
    input d_arr_mux_23__7 ;
    input d_arr_mux_23__6 ;
    input d_arr_mux_23__5 ;
    input d_arr_mux_23__4 ;
    input d_arr_mux_23__3 ;
    input d_arr_mux_23__2 ;
    input d_arr_mux_23__1 ;
    input d_arr_mux_23__0 ;
    input d_arr_mux_24__31 ;
    input d_arr_mux_24__30 ;
    input d_arr_mux_24__29 ;
    input d_arr_mux_24__28 ;
    input d_arr_mux_24__27 ;
    input d_arr_mux_24__26 ;
    input d_arr_mux_24__25 ;
    input d_arr_mux_24__24 ;
    input d_arr_mux_24__23 ;
    input d_arr_mux_24__22 ;
    input d_arr_mux_24__21 ;
    input d_arr_mux_24__20 ;
    input d_arr_mux_24__19 ;
    input d_arr_mux_24__18 ;
    input d_arr_mux_24__17 ;
    input d_arr_mux_24__16 ;
    input d_arr_mux_24__15 ;
    input d_arr_mux_24__14 ;
    input d_arr_mux_24__13 ;
    input d_arr_mux_24__12 ;
    input d_arr_mux_24__11 ;
    input d_arr_mux_24__10 ;
    input d_arr_mux_24__9 ;
    input d_arr_mux_24__8 ;
    input d_arr_mux_24__7 ;
    input d_arr_mux_24__6 ;
    input d_arr_mux_24__5 ;
    input d_arr_mux_24__4 ;
    input d_arr_mux_24__3 ;
    input d_arr_mux_24__2 ;
    input d_arr_mux_24__1 ;
    input d_arr_mux_24__0 ;
    input d_arr_mul_0__31 ;
    input d_arr_mul_0__30 ;
    input d_arr_mul_0__29 ;
    input d_arr_mul_0__28 ;
    input d_arr_mul_0__27 ;
    input d_arr_mul_0__26 ;
    input d_arr_mul_0__25 ;
    input d_arr_mul_0__24 ;
    input d_arr_mul_0__23 ;
    input d_arr_mul_0__22 ;
    input d_arr_mul_0__21 ;
    input d_arr_mul_0__20 ;
    input d_arr_mul_0__19 ;
    input d_arr_mul_0__18 ;
    input d_arr_mul_0__17 ;
    input d_arr_mul_0__16 ;
    input d_arr_mul_0__15 ;
    input d_arr_mul_0__14 ;
    input d_arr_mul_0__13 ;
    input d_arr_mul_0__12 ;
    input d_arr_mul_0__11 ;
    input d_arr_mul_0__10 ;
    input d_arr_mul_0__9 ;
    input d_arr_mul_0__8 ;
    input d_arr_mul_0__7 ;
    input d_arr_mul_0__6 ;
    input d_arr_mul_0__5 ;
    input d_arr_mul_0__4 ;
    input d_arr_mul_0__3 ;
    input d_arr_mul_0__2 ;
    input d_arr_mul_0__1 ;
    input d_arr_mul_0__0 ;
    input d_arr_mul_1__31 ;
    input d_arr_mul_1__30 ;
    input d_arr_mul_1__29 ;
    input d_arr_mul_1__28 ;
    input d_arr_mul_1__27 ;
    input d_arr_mul_1__26 ;
    input d_arr_mul_1__25 ;
    input d_arr_mul_1__24 ;
    input d_arr_mul_1__23 ;
    input d_arr_mul_1__22 ;
    input d_arr_mul_1__21 ;
    input d_arr_mul_1__20 ;
    input d_arr_mul_1__19 ;
    input d_arr_mul_1__18 ;
    input d_arr_mul_1__17 ;
    input d_arr_mul_1__16 ;
    input d_arr_mul_1__15 ;
    input d_arr_mul_1__14 ;
    input d_arr_mul_1__13 ;
    input d_arr_mul_1__12 ;
    input d_arr_mul_1__11 ;
    input d_arr_mul_1__10 ;
    input d_arr_mul_1__9 ;
    input d_arr_mul_1__8 ;
    input d_arr_mul_1__7 ;
    input d_arr_mul_1__6 ;
    input d_arr_mul_1__5 ;
    input d_arr_mul_1__4 ;
    input d_arr_mul_1__3 ;
    input d_arr_mul_1__2 ;
    input d_arr_mul_1__1 ;
    input d_arr_mul_1__0 ;
    input d_arr_mul_2__31 ;
    input d_arr_mul_2__30 ;
    input d_arr_mul_2__29 ;
    input d_arr_mul_2__28 ;
    input d_arr_mul_2__27 ;
    input d_arr_mul_2__26 ;
    input d_arr_mul_2__25 ;
    input d_arr_mul_2__24 ;
    input d_arr_mul_2__23 ;
    input d_arr_mul_2__22 ;
    input d_arr_mul_2__21 ;
    input d_arr_mul_2__20 ;
    input d_arr_mul_2__19 ;
    input d_arr_mul_2__18 ;
    input d_arr_mul_2__17 ;
    input d_arr_mul_2__16 ;
    input d_arr_mul_2__15 ;
    input d_arr_mul_2__14 ;
    input d_arr_mul_2__13 ;
    input d_arr_mul_2__12 ;
    input d_arr_mul_2__11 ;
    input d_arr_mul_2__10 ;
    input d_arr_mul_2__9 ;
    input d_arr_mul_2__8 ;
    input d_arr_mul_2__7 ;
    input d_arr_mul_2__6 ;
    input d_arr_mul_2__5 ;
    input d_arr_mul_2__4 ;
    input d_arr_mul_2__3 ;
    input d_arr_mul_2__2 ;
    input d_arr_mul_2__1 ;
    input d_arr_mul_2__0 ;
    input d_arr_mul_3__31 ;
    input d_arr_mul_3__30 ;
    input d_arr_mul_3__29 ;
    input d_arr_mul_3__28 ;
    input d_arr_mul_3__27 ;
    input d_arr_mul_3__26 ;
    input d_arr_mul_3__25 ;
    input d_arr_mul_3__24 ;
    input d_arr_mul_3__23 ;
    input d_arr_mul_3__22 ;
    input d_arr_mul_3__21 ;
    input d_arr_mul_3__20 ;
    input d_arr_mul_3__19 ;
    input d_arr_mul_3__18 ;
    input d_arr_mul_3__17 ;
    input d_arr_mul_3__16 ;
    input d_arr_mul_3__15 ;
    input d_arr_mul_3__14 ;
    input d_arr_mul_3__13 ;
    input d_arr_mul_3__12 ;
    input d_arr_mul_3__11 ;
    input d_arr_mul_3__10 ;
    input d_arr_mul_3__9 ;
    input d_arr_mul_3__8 ;
    input d_arr_mul_3__7 ;
    input d_arr_mul_3__6 ;
    input d_arr_mul_3__5 ;
    input d_arr_mul_3__4 ;
    input d_arr_mul_3__3 ;
    input d_arr_mul_3__2 ;
    input d_arr_mul_3__1 ;
    input d_arr_mul_3__0 ;
    input d_arr_mul_4__31 ;
    input d_arr_mul_4__30 ;
    input d_arr_mul_4__29 ;
    input d_arr_mul_4__28 ;
    input d_arr_mul_4__27 ;
    input d_arr_mul_4__26 ;
    input d_arr_mul_4__25 ;
    input d_arr_mul_4__24 ;
    input d_arr_mul_4__23 ;
    input d_arr_mul_4__22 ;
    input d_arr_mul_4__21 ;
    input d_arr_mul_4__20 ;
    input d_arr_mul_4__19 ;
    input d_arr_mul_4__18 ;
    input d_arr_mul_4__17 ;
    input d_arr_mul_4__16 ;
    input d_arr_mul_4__15 ;
    input d_arr_mul_4__14 ;
    input d_arr_mul_4__13 ;
    input d_arr_mul_4__12 ;
    input d_arr_mul_4__11 ;
    input d_arr_mul_4__10 ;
    input d_arr_mul_4__9 ;
    input d_arr_mul_4__8 ;
    input d_arr_mul_4__7 ;
    input d_arr_mul_4__6 ;
    input d_arr_mul_4__5 ;
    input d_arr_mul_4__4 ;
    input d_arr_mul_4__3 ;
    input d_arr_mul_4__2 ;
    input d_arr_mul_4__1 ;
    input d_arr_mul_4__0 ;
    input d_arr_mul_5__31 ;
    input d_arr_mul_5__30 ;
    input d_arr_mul_5__29 ;
    input d_arr_mul_5__28 ;
    input d_arr_mul_5__27 ;
    input d_arr_mul_5__26 ;
    input d_arr_mul_5__25 ;
    input d_arr_mul_5__24 ;
    input d_arr_mul_5__23 ;
    input d_arr_mul_5__22 ;
    input d_arr_mul_5__21 ;
    input d_arr_mul_5__20 ;
    input d_arr_mul_5__19 ;
    input d_arr_mul_5__18 ;
    input d_arr_mul_5__17 ;
    input d_arr_mul_5__16 ;
    input d_arr_mul_5__15 ;
    input d_arr_mul_5__14 ;
    input d_arr_mul_5__13 ;
    input d_arr_mul_5__12 ;
    input d_arr_mul_5__11 ;
    input d_arr_mul_5__10 ;
    input d_arr_mul_5__9 ;
    input d_arr_mul_5__8 ;
    input d_arr_mul_5__7 ;
    input d_arr_mul_5__6 ;
    input d_arr_mul_5__5 ;
    input d_arr_mul_5__4 ;
    input d_arr_mul_5__3 ;
    input d_arr_mul_5__2 ;
    input d_arr_mul_5__1 ;
    input d_arr_mul_5__0 ;
    input d_arr_mul_6__31 ;
    input d_arr_mul_6__30 ;
    input d_arr_mul_6__29 ;
    input d_arr_mul_6__28 ;
    input d_arr_mul_6__27 ;
    input d_arr_mul_6__26 ;
    input d_arr_mul_6__25 ;
    input d_arr_mul_6__24 ;
    input d_arr_mul_6__23 ;
    input d_arr_mul_6__22 ;
    input d_arr_mul_6__21 ;
    input d_arr_mul_6__20 ;
    input d_arr_mul_6__19 ;
    input d_arr_mul_6__18 ;
    input d_arr_mul_6__17 ;
    input d_arr_mul_6__16 ;
    input d_arr_mul_6__15 ;
    input d_arr_mul_6__14 ;
    input d_arr_mul_6__13 ;
    input d_arr_mul_6__12 ;
    input d_arr_mul_6__11 ;
    input d_arr_mul_6__10 ;
    input d_arr_mul_6__9 ;
    input d_arr_mul_6__8 ;
    input d_arr_mul_6__7 ;
    input d_arr_mul_6__6 ;
    input d_arr_mul_6__5 ;
    input d_arr_mul_6__4 ;
    input d_arr_mul_6__3 ;
    input d_arr_mul_6__2 ;
    input d_arr_mul_6__1 ;
    input d_arr_mul_6__0 ;
    input d_arr_mul_7__31 ;
    input d_arr_mul_7__30 ;
    input d_arr_mul_7__29 ;
    input d_arr_mul_7__28 ;
    input d_arr_mul_7__27 ;
    input d_arr_mul_7__26 ;
    input d_arr_mul_7__25 ;
    input d_arr_mul_7__24 ;
    input d_arr_mul_7__23 ;
    input d_arr_mul_7__22 ;
    input d_arr_mul_7__21 ;
    input d_arr_mul_7__20 ;
    input d_arr_mul_7__19 ;
    input d_arr_mul_7__18 ;
    input d_arr_mul_7__17 ;
    input d_arr_mul_7__16 ;
    input d_arr_mul_7__15 ;
    input d_arr_mul_7__14 ;
    input d_arr_mul_7__13 ;
    input d_arr_mul_7__12 ;
    input d_arr_mul_7__11 ;
    input d_arr_mul_7__10 ;
    input d_arr_mul_7__9 ;
    input d_arr_mul_7__8 ;
    input d_arr_mul_7__7 ;
    input d_arr_mul_7__6 ;
    input d_arr_mul_7__5 ;
    input d_arr_mul_7__4 ;
    input d_arr_mul_7__3 ;
    input d_arr_mul_7__2 ;
    input d_arr_mul_7__1 ;
    input d_arr_mul_7__0 ;
    input d_arr_mul_8__31 ;
    input d_arr_mul_8__30 ;
    input d_arr_mul_8__29 ;
    input d_arr_mul_8__28 ;
    input d_arr_mul_8__27 ;
    input d_arr_mul_8__26 ;
    input d_arr_mul_8__25 ;
    input d_arr_mul_8__24 ;
    input d_arr_mul_8__23 ;
    input d_arr_mul_8__22 ;
    input d_arr_mul_8__21 ;
    input d_arr_mul_8__20 ;
    input d_arr_mul_8__19 ;
    input d_arr_mul_8__18 ;
    input d_arr_mul_8__17 ;
    input d_arr_mul_8__16 ;
    input d_arr_mul_8__15 ;
    input d_arr_mul_8__14 ;
    input d_arr_mul_8__13 ;
    input d_arr_mul_8__12 ;
    input d_arr_mul_8__11 ;
    input d_arr_mul_8__10 ;
    input d_arr_mul_8__9 ;
    input d_arr_mul_8__8 ;
    input d_arr_mul_8__7 ;
    input d_arr_mul_8__6 ;
    input d_arr_mul_8__5 ;
    input d_arr_mul_8__4 ;
    input d_arr_mul_8__3 ;
    input d_arr_mul_8__2 ;
    input d_arr_mul_8__1 ;
    input d_arr_mul_8__0 ;
    input d_arr_mul_9__31 ;
    input d_arr_mul_9__30 ;
    input d_arr_mul_9__29 ;
    input d_arr_mul_9__28 ;
    input d_arr_mul_9__27 ;
    input d_arr_mul_9__26 ;
    input d_arr_mul_9__25 ;
    input d_arr_mul_9__24 ;
    input d_arr_mul_9__23 ;
    input d_arr_mul_9__22 ;
    input d_arr_mul_9__21 ;
    input d_arr_mul_9__20 ;
    input d_arr_mul_9__19 ;
    input d_arr_mul_9__18 ;
    input d_arr_mul_9__17 ;
    input d_arr_mul_9__16 ;
    input d_arr_mul_9__15 ;
    input d_arr_mul_9__14 ;
    input d_arr_mul_9__13 ;
    input d_arr_mul_9__12 ;
    input d_arr_mul_9__11 ;
    input d_arr_mul_9__10 ;
    input d_arr_mul_9__9 ;
    input d_arr_mul_9__8 ;
    input d_arr_mul_9__7 ;
    input d_arr_mul_9__6 ;
    input d_arr_mul_9__5 ;
    input d_arr_mul_9__4 ;
    input d_arr_mul_9__3 ;
    input d_arr_mul_9__2 ;
    input d_arr_mul_9__1 ;
    input d_arr_mul_9__0 ;
    input d_arr_mul_10__31 ;
    input d_arr_mul_10__30 ;
    input d_arr_mul_10__29 ;
    input d_arr_mul_10__28 ;
    input d_arr_mul_10__27 ;
    input d_arr_mul_10__26 ;
    input d_arr_mul_10__25 ;
    input d_arr_mul_10__24 ;
    input d_arr_mul_10__23 ;
    input d_arr_mul_10__22 ;
    input d_arr_mul_10__21 ;
    input d_arr_mul_10__20 ;
    input d_arr_mul_10__19 ;
    input d_arr_mul_10__18 ;
    input d_arr_mul_10__17 ;
    input d_arr_mul_10__16 ;
    input d_arr_mul_10__15 ;
    input d_arr_mul_10__14 ;
    input d_arr_mul_10__13 ;
    input d_arr_mul_10__12 ;
    input d_arr_mul_10__11 ;
    input d_arr_mul_10__10 ;
    input d_arr_mul_10__9 ;
    input d_arr_mul_10__8 ;
    input d_arr_mul_10__7 ;
    input d_arr_mul_10__6 ;
    input d_arr_mul_10__5 ;
    input d_arr_mul_10__4 ;
    input d_arr_mul_10__3 ;
    input d_arr_mul_10__2 ;
    input d_arr_mul_10__1 ;
    input d_arr_mul_10__0 ;
    input d_arr_mul_11__31 ;
    input d_arr_mul_11__30 ;
    input d_arr_mul_11__29 ;
    input d_arr_mul_11__28 ;
    input d_arr_mul_11__27 ;
    input d_arr_mul_11__26 ;
    input d_arr_mul_11__25 ;
    input d_arr_mul_11__24 ;
    input d_arr_mul_11__23 ;
    input d_arr_mul_11__22 ;
    input d_arr_mul_11__21 ;
    input d_arr_mul_11__20 ;
    input d_arr_mul_11__19 ;
    input d_arr_mul_11__18 ;
    input d_arr_mul_11__17 ;
    input d_arr_mul_11__16 ;
    input d_arr_mul_11__15 ;
    input d_arr_mul_11__14 ;
    input d_arr_mul_11__13 ;
    input d_arr_mul_11__12 ;
    input d_arr_mul_11__11 ;
    input d_arr_mul_11__10 ;
    input d_arr_mul_11__9 ;
    input d_arr_mul_11__8 ;
    input d_arr_mul_11__7 ;
    input d_arr_mul_11__6 ;
    input d_arr_mul_11__5 ;
    input d_arr_mul_11__4 ;
    input d_arr_mul_11__3 ;
    input d_arr_mul_11__2 ;
    input d_arr_mul_11__1 ;
    input d_arr_mul_11__0 ;
    input d_arr_mul_12__31 ;
    input d_arr_mul_12__30 ;
    input d_arr_mul_12__29 ;
    input d_arr_mul_12__28 ;
    input d_arr_mul_12__27 ;
    input d_arr_mul_12__26 ;
    input d_arr_mul_12__25 ;
    input d_arr_mul_12__24 ;
    input d_arr_mul_12__23 ;
    input d_arr_mul_12__22 ;
    input d_arr_mul_12__21 ;
    input d_arr_mul_12__20 ;
    input d_arr_mul_12__19 ;
    input d_arr_mul_12__18 ;
    input d_arr_mul_12__17 ;
    input d_arr_mul_12__16 ;
    input d_arr_mul_12__15 ;
    input d_arr_mul_12__14 ;
    input d_arr_mul_12__13 ;
    input d_arr_mul_12__12 ;
    input d_arr_mul_12__11 ;
    input d_arr_mul_12__10 ;
    input d_arr_mul_12__9 ;
    input d_arr_mul_12__8 ;
    input d_arr_mul_12__7 ;
    input d_arr_mul_12__6 ;
    input d_arr_mul_12__5 ;
    input d_arr_mul_12__4 ;
    input d_arr_mul_12__3 ;
    input d_arr_mul_12__2 ;
    input d_arr_mul_12__1 ;
    input d_arr_mul_12__0 ;
    input d_arr_mul_13__31 ;
    input d_arr_mul_13__30 ;
    input d_arr_mul_13__29 ;
    input d_arr_mul_13__28 ;
    input d_arr_mul_13__27 ;
    input d_arr_mul_13__26 ;
    input d_arr_mul_13__25 ;
    input d_arr_mul_13__24 ;
    input d_arr_mul_13__23 ;
    input d_arr_mul_13__22 ;
    input d_arr_mul_13__21 ;
    input d_arr_mul_13__20 ;
    input d_arr_mul_13__19 ;
    input d_arr_mul_13__18 ;
    input d_arr_mul_13__17 ;
    input d_arr_mul_13__16 ;
    input d_arr_mul_13__15 ;
    input d_arr_mul_13__14 ;
    input d_arr_mul_13__13 ;
    input d_arr_mul_13__12 ;
    input d_arr_mul_13__11 ;
    input d_arr_mul_13__10 ;
    input d_arr_mul_13__9 ;
    input d_arr_mul_13__8 ;
    input d_arr_mul_13__7 ;
    input d_arr_mul_13__6 ;
    input d_arr_mul_13__5 ;
    input d_arr_mul_13__4 ;
    input d_arr_mul_13__3 ;
    input d_arr_mul_13__2 ;
    input d_arr_mul_13__1 ;
    input d_arr_mul_13__0 ;
    input d_arr_mul_14__31 ;
    input d_arr_mul_14__30 ;
    input d_arr_mul_14__29 ;
    input d_arr_mul_14__28 ;
    input d_arr_mul_14__27 ;
    input d_arr_mul_14__26 ;
    input d_arr_mul_14__25 ;
    input d_arr_mul_14__24 ;
    input d_arr_mul_14__23 ;
    input d_arr_mul_14__22 ;
    input d_arr_mul_14__21 ;
    input d_arr_mul_14__20 ;
    input d_arr_mul_14__19 ;
    input d_arr_mul_14__18 ;
    input d_arr_mul_14__17 ;
    input d_arr_mul_14__16 ;
    input d_arr_mul_14__15 ;
    input d_arr_mul_14__14 ;
    input d_arr_mul_14__13 ;
    input d_arr_mul_14__12 ;
    input d_arr_mul_14__11 ;
    input d_arr_mul_14__10 ;
    input d_arr_mul_14__9 ;
    input d_arr_mul_14__8 ;
    input d_arr_mul_14__7 ;
    input d_arr_mul_14__6 ;
    input d_arr_mul_14__5 ;
    input d_arr_mul_14__4 ;
    input d_arr_mul_14__3 ;
    input d_arr_mul_14__2 ;
    input d_arr_mul_14__1 ;
    input d_arr_mul_14__0 ;
    input d_arr_mul_15__31 ;
    input d_arr_mul_15__30 ;
    input d_arr_mul_15__29 ;
    input d_arr_mul_15__28 ;
    input d_arr_mul_15__27 ;
    input d_arr_mul_15__26 ;
    input d_arr_mul_15__25 ;
    input d_arr_mul_15__24 ;
    input d_arr_mul_15__23 ;
    input d_arr_mul_15__22 ;
    input d_arr_mul_15__21 ;
    input d_arr_mul_15__20 ;
    input d_arr_mul_15__19 ;
    input d_arr_mul_15__18 ;
    input d_arr_mul_15__17 ;
    input d_arr_mul_15__16 ;
    input d_arr_mul_15__15 ;
    input d_arr_mul_15__14 ;
    input d_arr_mul_15__13 ;
    input d_arr_mul_15__12 ;
    input d_arr_mul_15__11 ;
    input d_arr_mul_15__10 ;
    input d_arr_mul_15__9 ;
    input d_arr_mul_15__8 ;
    input d_arr_mul_15__7 ;
    input d_arr_mul_15__6 ;
    input d_arr_mul_15__5 ;
    input d_arr_mul_15__4 ;
    input d_arr_mul_15__3 ;
    input d_arr_mul_15__2 ;
    input d_arr_mul_15__1 ;
    input d_arr_mul_15__0 ;
    input d_arr_mul_16__31 ;
    input d_arr_mul_16__30 ;
    input d_arr_mul_16__29 ;
    input d_arr_mul_16__28 ;
    input d_arr_mul_16__27 ;
    input d_arr_mul_16__26 ;
    input d_arr_mul_16__25 ;
    input d_arr_mul_16__24 ;
    input d_arr_mul_16__23 ;
    input d_arr_mul_16__22 ;
    input d_arr_mul_16__21 ;
    input d_arr_mul_16__20 ;
    input d_arr_mul_16__19 ;
    input d_arr_mul_16__18 ;
    input d_arr_mul_16__17 ;
    input d_arr_mul_16__16 ;
    input d_arr_mul_16__15 ;
    input d_arr_mul_16__14 ;
    input d_arr_mul_16__13 ;
    input d_arr_mul_16__12 ;
    input d_arr_mul_16__11 ;
    input d_arr_mul_16__10 ;
    input d_arr_mul_16__9 ;
    input d_arr_mul_16__8 ;
    input d_arr_mul_16__7 ;
    input d_arr_mul_16__6 ;
    input d_arr_mul_16__5 ;
    input d_arr_mul_16__4 ;
    input d_arr_mul_16__3 ;
    input d_arr_mul_16__2 ;
    input d_arr_mul_16__1 ;
    input d_arr_mul_16__0 ;
    input d_arr_mul_17__31 ;
    input d_arr_mul_17__30 ;
    input d_arr_mul_17__29 ;
    input d_arr_mul_17__28 ;
    input d_arr_mul_17__27 ;
    input d_arr_mul_17__26 ;
    input d_arr_mul_17__25 ;
    input d_arr_mul_17__24 ;
    input d_arr_mul_17__23 ;
    input d_arr_mul_17__22 ;
    input d_arr_mul_17__21 ;
    input d_arr_mul_17__20 ;
    input d_arr_mul_17__19 ;
    input d_arr_mul_17__18 ;
    input d_arr_mul_17__17 ;
    input d_arr_mul_17__16 ;
    input d_arr_mul_17__15 ;
    input d_arr_mul_17__14 ;
    input d_arr_mul_17__13 ;
    input d_arr_mul_17__12 ;
    input d_arr_mul_17__11 ;
    input d_arr_mul_17__10 ;
    input d_arr_mul_17__9 ;
    input d_arr_mul_17__8 ;
    input d_arr_mul_17__7 ;
    input d_arr_mul_17__6 ;
    input d_arr_mul_17__5 ;
    input d_arr_mul_17__4 ;
    input d_arr_mul_17__3 ;
    input d_arr_mul_17__2 ;
    input d_arr_mul_17__1 ;
    input d_arr_mul_17__0 ;
    input d_arr_mul_18__31 ;
    input d_arr_mul_18__30 ;
    input d_arr_mul_18__29 ;
    input d_arr_mul_18__28 ;
    input d_arr_mul_18__27 ;
    input d_arr_mul_18__26 ;
    input d_arr_mul_18__25 ;
    input d_arr_mul_18__24 ;
    input d_arr_mul_18__23 ;
    input d_arr_mul_18__22 ;
    input d_arr_mul_18__21 ;
    input d_arr_mul_18__20 ;
    input d_arr_mul_18__19 ;
    input d_arr_mul_18__18 ;
    input d_arr_mul_18__17 ;
    input d_arr_mul_18__16 ;
    input d_arr_mul_18__15 ;
    input d_arr_mul_18__14 ;
    input d_arr_mul_18__13 ;
    input d_arr_mul_18__12 ;
    input d_arr_mul_18__11 ;
    input d_arr_mul_18__10 ;
    input d_arr_mul_18__9 ;
    input d_arr_mul_18__8 ;
    input d_arr_mul_18__7 ;
    input d_arr_mul_18__6 ;
    input d_arr_mul_18__5 ;
    input d_arr_mul_18__4 ;
    input d_arr_mul_18__3 ;
    input d_arr_mul_18__2 ;
    input d_arr_mul_18__1 ;
    input d_arr_mul_18__0 ;
    input d_arr_mul_19__31 ;
    input d_arr_mul_19__30 ;
    input d_arr_mul_19__29 ;
    input d_arr_mul_19__28 ;
    input d_arr_mul_19__27 ;
    input d_arr_mul_19__26 ;
    input d_arr_mul_19__25 ;
    input d_arr_mul_19__24 ;
    input d_arr_mul_19__23 ;
    input d_arr_mul_19__22 ;
    input d_arr_mul_19__21 ;
    input d_arr_mul_19__20 ;
    input d_arr_mul_19__19 ;
    input d_arr_mul_19__18 ;
    input d_arr_mul_19__17 ;
    input d_arr_mul_19__16 ;
    input d_arr_mul_19__15 ;
    input d_arr_mul_19__14 ;
    input d_arr_mul_19__13 ;
    input d_arr_mul_19__12 ;
    input d_arr_mul_19__11 ;
    input d_arr_mul_19__10 ;
    input d_arr_mul_19__9 ;
    input d_arr_mul_19__8 ;
    input d_arr_mul_19__7 ;
    input d_arr_mul_19__6 ;
    input d_arr_mul_19__5 ;
    input d_arr_mul_19__4 ;
    input d_arr_mul_19__3 ;
    input d_arr_mul_19__2 ;
    input d_arr_mul_19__1 ;
    input d_arr_mul_19__0 ;
    input d_arr_mul_20__31 ;
    input d_arr_mul_20__30 ;
    input d_arr_mul_20__29 ;
    input d_arr_mul_20__28 ;
    input d_arr_mul_20__27 ;
    input d_arr_mul_20__26 ;
    input d_arr_mul_20__25 ;
    input d_arr_mul_20__24 ;
    input d_arr_mul_20__23 ;
    input d_arr_mul_20__22 ;
    input d_arr_mul_20__21 ;
    input d_arr_mul_20__20 ;
    input d_arr_mul_20__19 ;
    input d_arr_mul_20__18 ;
    input d_arr_mul_20__17 ;
    input d_arr_mul_20__16 ;
    input d_arr_mul_20__15 ;
    input d_arr_mul_20__14 ;
    input d_arr_mul_20__13 ;
    input d_arr_mul_20__12 ;
    input d_arr_mul_20__11 ;
    input d_arr_mul_20__10 ;
    input d_arr_mul_20__9 ;
    input d_arr_mul_20__8 ;
    input d_arr_mul_20__7 ;
    input d_arr_mul_20__6 ;
    input d_arr_mul_20__5 ;
    input d_arr_mul_20__4 ;
    input d_arr_mul_20__3 ;
    input d_arr_mul_20__2 ;
    input d_arr_mul_20__1 ;
    input d_arr_mul_20__0 ;
    input d_arr_mul_21__31 ;
    input d_arr_mul_21__30 ;
    input d_arr_mul_21__29 ;
    input d_arr_mul_21__28 ;
    input d_arr_mul_21__27 ;
    input d_arr_mul_21__26 ;
    input d_arr_mul_21__25 ;
    input d_arr_mul_21__24 ;
    input d_arr_mul_21__23 ;
    input d_arr_mul_21__22 ;
    input d_arr_mul_21__21 ;
    input d_arr_mul_21__20 ;
    input d_arr_mul_21__19 ;
    input d_arr_mul_21__18 ;
    input d_arr_mul_21__17 ;
    input d_arr_mul_21__16 ;
    input d_arr_mul_21__15 ;
    input d_arr_mul_21__14 ;
    input d_arr_mul_21__13 ;
    input d_arr_mul_21__12 ;
    input d_arr_mul_21__11 ;
    input d_arr_mul_21__10 ;
    input d_arr_mul_21__9 ;
    input d_arr_mul_21__8 ;
    input d_arr_mul_21__7 ;
    input d_arr_mul_21__6 ;
    input d_arr_mul_21__5 ;
    input d_arr_mul_21__4 ;
    input d_arr_mul_21__3 ;
    input d_arr_mul_21__2 ;
    input d_arr_mul_21__1 ;
    input d_arr_mul_21__0 ;
    input d_arr_mul_22__31 ;
    input d_arr_mul_22__30 ;
    input d_arr_mul_22__29 ;
    input d_arr_mul_22__28 ;
    input d_arr_mul_22__27 ;
    input d_arr_mul_22__26 ;
    input d_arr_mul_22__25 ;
    input d_arr_mul_22__24 ;
    input d_arr_mul_22__23 ;
    input d_arr_mul_22__22 ;
    input d_arr_mul_22__21 ;
    input d_arr_mul_22__20 ;
    input d_arr_mul_22__19 ;
    input d_arr_mul_22__18 ;
    input d_arr_mul_22__17 ;
    input d_arr_mul_22__16 ;
    input d_arr_mul_22__15 ;
    input d_arr_mul_22__14 ;
    input d_arr_mul_22__13 ;
    input d_arr_mul_22__12 ;
    input d_arr_mul_22__11 ;
    input d_arr_mul_22__10 ;
    input d_arr_mul_22__9 ;
    input d_arr_mul_22__8 ;
    input d_arr_mul_22__7 ;
    input d_arr_mul_22__6 ;
    input d_arr_mul_22__5 ;
    input d_arr_mul_22__4 ;
    input d_arr_mul_22__3 ;
    input d_arr_mul_22__2 ;
    input d_arr_mul_22__1 ;
    input d_arr_mul_22__0 ;
    input d_arr_mul_23__31 ;
    input d_arr_mul_23__30 ;
    input d_arr_mul_23__29 ;
    input d_arr_mul_23__28 ;
    input d_arr_mul_23__27 ;
    input d_arr_mul_23__26 ;
    input d_arr_mul_23__25 ;
    input d_arr_mul_23__24 ;
    input d_arr_mul_23__23 ;
    input d_arr_mul_23__22 ;
    input d_arr_mul_23__21 ;
    input d_arr_mul_23__20 ;
    input d_arr_mul_23__19 ;
    input d_arr_mul_23__18 ;
    input d_arr_mul_23__17 ;
    input d_arr_mul_23__16 ;
    input d_arr_mul_23__15 ;
    input d_arr_mul_23__14 ;
    input d_arr_mul_23__13 ;
    input d_arr_mul_23__12 ;
    input d_arr_mul_23__11 ;
    input d_arr_mul_23__10 ;
    input d_arr_mul_23__9 ;
    input d_arr_mul_23__8 ;
    input d_arr_mul_23__7 ;
    input d_arr_mul_23__6 ;
    input d_arr_mul_23__5 ;
    input d_arr_mul_23__4 ;
    input d_arr_mul_23__3 ;
    input d_arr_mul_23__2 ;
    input d_arr_mul_23__1 ;
    input d_arr_mul_23__0 ;
    input d_arr_mul_24__31 ;
    input d_arr_mul_24__30 ;
    input d_arr_mul_24__29 ;
    input d_arr_mul_24__28 ;
    input d_arr_mul_24__27 ;
    input d_arr_mul_24__26 ;
    input d_arr_mul_24__25 ;
    input d_arr_mul_24__24 ;
    input d_arr_mul_24__23 ;
    input d_arr_mul_24__22 ;
    input d_arr_mul_24__21 ;
    input d_arr_mul_24__20 ;
    input d_arr_mul_24__19 ;
    input d_arr_mul_24__18 ;
    input d_arr_mul_24__17 ;
    input d_arr_mul_24__16 ;
    input d_arr_mul_24__15 ;
    input d_arr_mul_24__14 ;
    input d_arr_mul_24__13 ;
    input d_arr_mul_24__12 ;
    input d_arr_mul_24__11 ;
    input d_arr_mul_24__10 ;
    input d_arr_mul_24__9 ;
    input d_arr_mul_24__8 ;
    input d_arr_mul_24__7 ;
    input d_arr_mul_24__6 ;
    input d_arr_mul_24__5 ;
    input d_arr_mul_24__4 ;
    input d_arr_mul_24__3 ;
    input d_arr_mul_24__2 ;
    input d_arr_mul_24__1 ;
    input d_arr_mul_24__0 ;
    input d_arr_add_0__31 ;
    input d_arr_add_0__30 ;
    input d_arr_add_0__29 ;
    input d_arr_add_0__28 ;
    input d_arr_add_0__27 ;
    input d_arr_add_0__26 ;
    input d_arr_add_0__25 ;
    input d_arr_add_0__24 ;
    input d_arr_add_0__23 ;
    input d_arr_add_0__22 ;
    input d_arr_add_0__21 ;
    input d_arr_add_0__20 ;
    input d_arr_add_0__19 ;
    input d_arr_add_0__18 ;
    input d_arr_add_0__17 ;
    input d_arr_add_0__16 ;
    input d_arr_add_0__15 ;
    input d_arr_add_0__14 ;
    input d_arr_add_0__13 ;
    input d_arr_add_0__12 ;
    input d_arr_add_0__11 ;
    input d_arr_add_0__10 ;
    input d_arr_add_0__9 ;
    input d_arr_add_0__8 ;
    input d_arr_add_0__7 ;
    input d_arr_add_0__6 ;
    input d_arr_add_0__5 ;
    input d_arr_add_0__4 ;
    input d_arr_add_0__3 ;
    input d_arr_add_0__2 ;
    input d_arr_add_0__1 ;
    input d_arr_add_0__0 ;
    input d_arr_add_1__31 ;
    input d_arr_add_1__30 ;
    input d_arr_add_1__29 ;
    input d_arr_add_1__28 ;
    input d_arr_add_1__27 ;
    input d_arr_add_1__26 ;
    input d_arr_add_1__25 ;
    input d_arr_add_1__24 ;
    input d_arr_add_1__23 ;
    input d_arr_add_1__22 ;
    input d_arr_add_1__21 ;
    input d_arr_add_1__20 ;
    input d_arr_add_1__19 ;
    input d_arr_add_1__18 ;
    input d_arr_add_1__17 ;
    input d_arr_add_1__16 ;
    input d_arr_add_1__15 ;
    input d_arr_add_1__14 ;
    input d_arr_add_1__13 ;
    input d_arr_add_1__12 ;
    input d_arr_add_1__11 ;
    input d_arr_add_1__10 ;
    input d_arr_add_1__9 ;
    input d_arr_add_1__8 ;
    input d_arr_add_1__7 ;
    input d_arr_add_1__6 ;
    input d_arr_add_1__5 ;
    input d_arr_add_1__4 ;
    input d_arr_add_1__3 ;
    input d_arr_add_1__2 ;
    input d_arr_add_1__1 ;
    input d_arr_add_1__0 ;
    input d_arr_add_2__31 ;
    input d_arr_add_2__30 ;
    input d_arr_add_2__29 ;
    input d_arr_add_2__28 ;
    input d_arr_add_2__27 ;
    input d_arr_add_2__26 ;
    input d_arr_add_2__25 ;
    input d_arr_add_2__24 ;
    input d_arr_add_2__23 ;
    input d_arr_add_2__22 ;
    input d_arr_add_2__21 ;
    input d_arr_add_2__20 ;
    input d_arr_add_2__19 ;
    input d_arr_add_2__18 ;
    input d_arr_add_2__17 ;
    input d_arr_add_2__16 ;
    input d_arr_add_2__15 ;
    input d_arr_add_2__14 ;
    input d_arr_add_2__13 ;
    input d_arr_add_2__12 ;
    input d_arr_add_2__11 ;
    input d_arr_add_2__10 ;
    input d_arr_add_2__9 ;
    input d_arr_add_2__8 ;
    input d_arr_add_2__7 ;
    input d_arr_add_2__6 ;
    input d_arr_add_2__5 ;
    input d_arr_add_2__4 ;
    input d_arr_add_2__3 ;
    input d_arr_add_2__2 ;
    input d_arr_add_2__1 ;
    input d_arr_add_2__0 ;
    input d_arr_add_3__31 ;
    input d_arr_add_3__30 ;
    input d_arr_add_3__29 ;
    input d_arr_add_3__28 ;
    input d_arr_add_3__27 ;
    input d_arr_add_3__26 ;
    input d_arr_add_3__25 ;
    input d_arr_add_3__24 ;
    input d_arr_add_3__23 ;
    input d_arr_add_3__22 ;
    input d_arr_add_3__21 ;
    input d_arr_add_3__20 ;
    input d_arr_add_3__19 ;
    input d_arr_add_3__18 ;
    input d_arr_add_3__17 ;
    input d_arr_add_3__16 ;
    input d_arr_add_3__15 ;
    input d_arr_add_3__14 ;
    input d_arr_add_3__13 ;
    input d_arr_add_3__12 ;
    input d_arr_add_3__11 ;
    input d_arr_add_3__10 ;
    input d_arr_add_3__9 ;
    input d_arr_add_3__8 ;
    input d_arr_add_3__7 ;
    input d_arr_add_3__6 ;
    input d_arr_add_3__5 ;
    input d_arr_add_3__4 ;
    input d_arr_add_3__3 ;
    input d_arr_add_3__2 ;
    input d_arr_add_3__1 ;
    input d_arr_add_3__0 ;
    input d_arr_add_4__31 ;
    input d_arr_add_4__30 ;
    input d_arr_add_4__29 ;
    input d_arr_add_4__28 ;
    input d_arr_add_4__27 ;
    input d_arr_add_4__26 ;
    input d_arr_add_4__25 ;
    input d_arr_add_4__24 ;
    input d_arr_add_4__23 ;
    input d_arr_add_4__22 ;
    input d_arr_add_4__21 ;
    input d_arr_add_4__20 ;
    input d_arr_add_4__19 ;
    input d_arr_add_4__18 ;
    input d_arr_add_4__17 ;
    input d_arr_add_4__16 ;
    input d_arr_add_4__15 ;
    input d_arr_add_4__14 ;
    input d_arr_add_4__13 ;
    input d_arr_add_4__12 ;
    input d_arr_add_4__11 ;
    input d_arr_add_4__10 ;
    input d_arr_add_4__9 ;
    input d_arr_add_4__8 ;
    input d_arr_add_4__7 ;
    input d_arr_add_4__6 ;
    input d_arr_add_4__5 ;
    input d_arr_add_4__4 ;
    input d_arr_add_4__3 ;
    input d_arr_add_4__2 ;
    input d_arr_add_4__1 ;
    input d_arr_add_4__0 ;
    input d_arr_add_5__31 ;
    input d_arr_add_5__30 ;
    input d_arr_add_5__29 ;
    input d_arr_add_5__28 ;
    input d_arr_add_5__27 ;
    input d_arr_add_5__26 ;
    input d_arr_add_5__25 ;
    input d_arr_add_5__24 ;
    input d_arr_add_5__23 ;
    input d_arr_add_5__22 ;
    input d_arr_add_5__21 ;
    input d_arr_add_5__20 ;
    input d_arr_add_5__19 ;
    input d_arr_add_5__18 ;
    input d_arr_add_5__17 ;
    input d_arr_add_5__16 ;
    input d_arr_add_5__15 ;
    input d_arr_add_5__14 ;
    input d_arr_add_5__13 ;
    input d_arr_add_5__12 ;
    input d_arr_add_5__11 ;
    input d_arr_add_5__10 ;
    input d_arr_add_5__9 ;
    input d_arr_add_5__8 ;
    input d_arr_add_5__7 ;
    input d_arr_add_5__6 ;
    input d_arr_add_5__5 ;
    input d_arr_add_5__4 ;
    input d_arr_add_5__3 ;
    input d_arr_add_5__2 ;
    input d_arr_add_5__1 ;
    input d_arr_add_5__0 ;
    input d_arr_add_6__31 ;
    input d_arr_add_6__30 ;
    input d_arr_add_6__29 ;
    input d_arr_add_6__28 ;
    input d_arr_add_6__27 ;
    input d_arr_add_6__26 ;
    input d_arr_add_6__25 ;
    input d_arr_add_6__24 ;
    input d_arr_add_6__23 ;
    input d_arr_add_6__22 ;
    input d_arr_add_6__21 ;
    input d_arr_add_6__20 ;
    input d_arr_add_6__19 ;
    input d_arr_add_6__18 ;
    input d_arr_add_6__17 ;
    input d_arr_add_6__16 ;
    input d_arr_add_6__15 ;
    input d_arr_add_6__14 ;
    input d_arr_add_6__13 ;
    input d_arr_add_6__12 ;
    input d_arr_add_6__11 ;
    input d_arr_add_6__10 ;
    input d_arr_add_6__9 ;
    input d_arr_add_6__8 ;
    input d_arr_add_6__7 ;
    input d_arr_add_6__6 ;
    input d_arr_add_6__5 ;
    input d_arr_add_6__4 ;
    input d_arr_add_6__3 ;
    input d_arr_add_6__2 ;
    input d_arr_add_6__1 ;
    input d_arr_add_6__0 ;
    input d_arr_add_7__31 ;
    input d_arr_add_7__30 ;
    input d_arr_add_7__29 ;
    input d_arr_add_7__28 ;
    input d_arr_add_7__27 ;
    input d_arr_add_7__26 ;
    input d_arr_add_7__25 ;
    input d_arr_add_7__24 ;
    input d_arr_add_7__23 ;
    input d_arr_add_7__22 ;
    input d_arr_add_7__21 ;
    input d_arr_add_7__20 ;
    input d_arr_add_7__19 ;
    input d_arr_add_7__18 ;
    input d_arr_add_7__17 ;
    input d_arr_add_7__16 ;
    input d_arr_add_7__15 ;
    input d_arr_add_7__14 ;
    input d_arr_add_7__13 ;
    input d_arr_add_7__12 ;
    input d_arr_add_7__11 ;
    input d_arr_add_7__10 ;
    input d_arr_add_7__9 ;
    input d_arr_add_7__8 ;
    input d_arr_add_7__7 ;
    input d_arr_add_7__6 ;
    input d_arr_add_7__5 ;
    input d_arr_add_7__4 ;
    input d_arr_add_7__3 ;
    input d_arr_add_7__2 ;
    input d_arr_add_7__1 ;
    input d_arr_add_7__0 ;
    input d_arr_add_8__31 ;
    input d_arr_add_8__30 ;
    input d_arr_add_8__29 ;
    input d_arr_add_8__28 ;
    input d_arr_add_8__27 ;
    input d_arr_add_8__26 ;
    input d_arr_add_8__25 ;
    input d_arr_add_8__24 ;
    input d_arr_add_8__23 ;
    input d_arr_add_8__22 ;
    input d_arr_add_8__21 ;
    input d_arr_add_8__20 ;
    input d_arr_add_8__19 ;
    input d_arr_add_8__18 ;
    input d_arr_add_8__17 ;
    input d_arr_add_8__16 ;
    input d_arr_add_8__15 ;
    input d_arr_add_8__14 ;
    input d_arr_add_8__13 ;
    input d_arr_add_8__12 ;
    input d_arr_add_8__11 ;
    input d_arr_add_8__10 ;
    input d_arr_add_8__9 ;
    input d_arr_add_8__8 ;
    input d_arr_add_8__7 ;
    input d_arr_add_8__6 ;
    input d_arr_add_8__5 ;
    input d_arr_add_8__4 ;
    input d_arr_add_8__3 ;
    input d_arr_add_8__2 ;
    input d_arr_add_8__1 ;
    input d_arr_add_8__0 ;
    input d_arr_add_9__31 ;
    input d_arr_add_9__30 ;
    input d_arr_add_9__29 ;
    input d_arr_add_9__28 ;
    input d_arr_add_9__27 ;
    input d_arr_add_9__26 ;
    input d_arr_add_9__25 ;
    input d_arr_add_9__24 ;
    input d_arr_add_9__23 ;
    input d_arr_add_9__22 ;
    input d_arr_add_9__21 ;
    input d_arr_add_9__20 ;
    input d_arr_add_9__19 ;
    input d_arr_add_9__18 ;
    input d_arr_add_9__17 ;
    input d_arr_add_9__16 ;
    input d_arr_add_9__15 ;
    input d_arr_add_9__14 ;
    input d_arr_add_9__13 ;
    input d_arr_add_9__12 ;
    input d_arr_add_9__11 ;
    input d_arr_add_9__10 ;
    input d_arr_add_9__9 ;
    input d_arr_add_9__8 ;
    input d_arr_add_9__7 ;
    input d_arr_add_9__6 ;
    input d_arr_add_9__5 ;
    input d_arr_add_9__4 ;
    input d_arr_add_9__3 ;
    input d_arr_add_9__2 ;
    input d_arr_add_9__1 ;
    input d_arr_add_9__0 ;
    input d_arr_add_10__31 ;
    input d_arr_add_10__30 ;
    input d_arr_add_10__29 ;
    input d_arr_add_10__28 ;
    input d_arr_add_10__27 ;
    input d_arr_add_10__26 ;
    input d_arr_add_10__25 ;
    input d_arr_add_10__24 ;
    input d_arr_add_10__23 ;
    input d_arr_add_10__22 ;
    input d_arr_add_10__21 ;
    input d_arr_add_10__20 ;
    input d_arr_add_10__19 ;
    input d_arr_add_10__18 ;
    input d_arr_add_10__17 ;
    input d_arr_add_10__16 ;
    input d_arr_add_10__15 ;
    input d_arr_add_10__14 ;
    input d_arr_add_10__13 ;
    input d_arr_add_10__12 ;
    input d_arr_add_10__11 ;
    input d_arr_add_10__10 ;
    input d_arr_add_10__9 ;
    input d_arr_add_10__8 ;
    input d_arr_add_10__7 ;
    input d_arr_add_10__6 ;
    input d_arr_add_10__5 ;
    input d_arr_add_10__4 ;
    input d_arr_add_10__3 ;
    input d_arr_add_10__2 ;
    input d_arr_add_10__1 ;
    input d_arr_add_10__0 ;
    input d_arr_add_11__31 ;
    input d_arr_add_11__30 ;
    input d_arr_add_11__29 ;
    input d_arr_add_11__28 ;
    input d_arr_add_11__27 ;
    input d_arr_add_11__26 ;
    input d_arr_add_11__25 ;
    input d_arr_add_11__24 ;
    input d_arr_add_11__23 ;
    input d_arr_add_11__22 ;
    input d_arr_add_11__21 ;
    input d_arr_add_11__20 ;
    input d_arr_add_11__19 ;
    input d_arr_add_11__18 ;
    input d_arr_add_11__17 ;
    input d_arr_add_11__16 ;
    input d_arr_add_11__15 ;
    input d_arr_add_11__14 ;
    input d_arr_add_11__13 ;
    input d_arr_add_11__12 ;
    input d_arr_add_11__11 ;
    input d_arr_add_11__10 ;
    input d_arr_add_11__9 ;
    input d_arr_add_11__8 ;
    input d_arr_add_11__7 ;
    input d_arr_add_11__6 ;
    input d_arr_add_11__5 ;
    input d_arr_add_11__4 ;
    input d_arr_add_11__3 ;
    input d_arr_add_11__2 ;
    input d_arr_add_11__1 ;
    input d_arr_add_11__0 ;
    input d_arr_add_12__31 ;
    input d_arr_add_12__30 ;
    input d_arr_add_12__29 ;
    input d_arr_add_12__28 ;
    input d_arr_add_12__27 ;
    input d_arr_add_12__26 ;
    input d_arr_add_12__25 ;
    input d_arr_add_12__24 ;
    input d_arr_add_12__23 ;
    input d_arr_add_12__22 ;
    input d_arr_add_12__21 ;
    input d_arr_add_12__20 ;
    input d_arr_add_12__19 ;
    input d_arr_add_12__18 ;
    input d_arr_add_12__17 ;
    input d_arr_add_12__16 ;
    input d_arr_add_12__15 ;
    input d_arr_add_12__14 ;
    input d_arr_add_12__13 ;
    input d_arr_add_12__12 ;
    input d_arr_add_12__11 ;
    input d_arr_add_12__10 ;
    input d_arr_add_12__9 ;
    input d_arr_add_12__8 ;
    input d_arr_add_12__7 ;
    input d_arr_add_12__6 ;
    input d_arr_add_12__5 ;
    input d_arr_add_12__4 ;
    input d_arr_add_12__3 ;
    input d_arr_add_12__2 ;
    input d_arr_add_12__1 ;
    input d_arr_add_12__0 ;
    input d_arr_add_13__31 ;
    input d_arr_add_13__30 ;
    input d_arr_add_13__29 ;
    input d_arr_add_13__28 ;
    input d_arr_add_13__27 ;
    input d_arr_add_13__26 ;
    input d_arr_add_13__25 ;
    input d_arr_add_13__24 ;
    input d_arr_add_13__23 ;
    input d_arr_add_13__22 ;
    input d_arr_add_13__21 ;
    input d_arr_add_13__20 ;
    input d_arr_add_13__19 ;
    input d_arr_add_13__18 ;
    input d_arr_add_13__17 ;
    input d_arr_add_13__16 ;
    input d_arr_add_13__15 ;
    input d_arr_add_13__14 ;
    input d_arr_add_13__13 ;
    input d_arr_add_13__12 ;
    input d_arr_add_13__11 ;
    input d_arr_add_13__10 ;
    input d_arr_add_13__9 ;
    input d_arr_add_13__8 ;
    input d_arr_add_13__7 ;
    input d_arr_add_13__6 ;
    input d_arr_add_13__5 ;
    input d_arr_add_13__4 ;
    input d_arr_add_13__3 ;
    input d_arr_add_13__2 ;
    input d_arr_add_13__1 ;
    input d_arr_add_13__0 ;
    input d_arr_add_14__31 ;
    input d_arr_add_14__30 ;
    input d_arr_add_14__29 ;
    input d_arr_add_14__28 ;
    input d_arr_add_14__27 ;
    input d_arr_add_14__26 ;
    input d_arr_add_14__25 ;
    input d_arr_add_14__24 ;
    input d_arr_add_14__23 ;
    input d_arr_add_14__22 ;
    input d_arr_add_14__21 ;
    input d_arr_add_14__20 ;
    input d_arr_add_14__19 ;
    input d_arr_add_14__18 ;
    input d_arr_add_14__17 ;
    input d_arr_add_14__16 ;
    input d_arr_add_14__15 ;
    input d_arr_add_14__14 ;
    input d_arr_add_14__13 ;
    input d_arr_add_14__12 ;
    input d_arr_add_14__11 ;
    input d_arr_add_14__10 ;
    input d_arr_add_14__9 ;
    input d_arr_add_14__8 ;
    input d_arr_add_14__7 ;
    input d_arr_add_14__6 ;
    input d_arr_add_14__5 ;
    input d_arr_add_14__4 ;
    input d_arr_add_14__3 ;
    input d_arr_add_14__2 ;
    input d_arr_add_14__1 ;
    input d_arr_add_14__0 ;
    input d_arr_add_15__31 ;
    input d_arr_add_15__30 ;
    input d_arr_add_15__29 ;
    input d_arr_add_15__28 ;
    input d_arr_add_15__27 ;
    input d_arr_add_15__26 ;
    input d_arr_add_15__25 ;
    input d_arr_add_15__24 ;
    input d_arr_add_15__23 ;
    input d_arr_add_15__22 ;
    input d_arr_add_15__21 ;
    input d_arr_add_15__20 ;
    input d_arr_add_15__19 ;
    input d_arr_add_15__18 ;
    input d_arr_add_15__17 ;
    input d_arr_add_15__16 ;
    input d_arr_add_15__15 ;
    input d_arr_add_15__14 ;
    input d_arr_add_15__13 ;
    input d_arr_add_15__12 ;
    input d_arr_add_15__11 ;
    input d_arr_add_15__10 ;
    input d_arr_add_15__9 ;
    input d_arr_add_15__8 ;
    input d_arr_add_15__7 ;
    input d_arr_add_15__6 ;
    input d_arr_add_15__5 ;
    input d_arr_add_15__4 ;
    input d_arr_add_15__3 ;
    input d_arr_add_15__2 ;
    input d_arr_add_15__1 ;
    input d_arr_add_15__0 ;
    input d_arr_add_16__31 ;
    input d_arr_add_16__30 ;
    input d_arr_add_16__29 ;
    input d_arr_add_16__28 ;
    input d_arr_add_16__27 ;
    input d_arr_add_16__26 ;
    input d_arr_add_16__25 ;
    input d_arr_add_16__24 ;
    input d_arr_add_16__23 ;
    input d_arr_add_16__22 ;
    input d_arr_add_16__21 ;
    input d_arr_add_16__20 ;
    input d_arr_add_16__19 ;
    input d_arr_add_16__18 ;
    input d_arr_add_16__17 ;
    input d_arr_add_16__16 ;
    input d_arr_add_16__15 ;
    input d_arr_add_16__14 ;
    input d_arr_add_16__13 ;
    input d_arr_add_16__12 ;
    input d_arr_add_16__11 ;
    input d_arr_add_16__10 ;
    input d_arr_add_16__9 ;
    input d_arr_add_16__8 ;
    input d_arr_add_16__7 ;
    input d_arr_add_16__6 ;
    input d_arr_add_16__5 ;
    input d_arr_add_16__4 ;
    input d_arr_add_16__3 ;
    input d_arr_add_16__2 ;
    input d_arr_add_16__1 ;
    input d_arr_add_16__0 ;
    input d_arr_add_17__31 ;
    input d_arr_add_17__30 ;
    input d_arr_add_17__29 ;
    input d_arr_add_17__28 ;
    input d_arr_add_17__27 ;
    input d_arr_add_17__26 ;
    input d_arr_add_17__25 ;
    input d_arr_add_17__24 ;
    input d_arr_add_17__23 ;
    input d_arr_add_17__22 ;
    input d_arr_add_17__21 ;
    input d_arr_add_17__20 ;
    input d_arr_add_17__19 ;
    input d_arr_add_17__18 ;
    input d_arr_add_17__17 ;
    input d_arr_add_17__16 ;
    input d_arr_add_17__15 ;
    input d_arr_add_17__14 ;
    input d_arr_add_17__13 ;
    input d_arr_add_17__12 ;
    input d_arr_add_17__11 ;
    input d_arr_add_17__10 ;
    input d_arr_add_17__9 ;
    input d_arr_add_17__8 ;
    input d_arr_add_17__7 ;
    input d_arr_add_17__6 ;
    input d_arr_add_17__5 ;
    input d_arr_add_17__4 ;
    input d_arr_add_17__3 ;
    input d_arr_add_17__2 ;
    input d_arr_add_17__1 ;
    input d_arr_add_17__0 ;
    input d_arr_add_18__31 ;
    input d_arr_add_18__30 ;
    input d_arr_add_18__29 ;
    input d_arr_add_18__28 ;
    input d_arr_add_18__27 ;
    input d_arr_add_18__26 ;
    input d_arr_add_18__25 ;
    input d_arr_add_18__24 ;
    input d_arr_add_18__23 ;
    input d_arr_add_18__22 ;
    input d_arr_add_18__21 ;
    input d_arr_add_18__20 ;
    input d_arr_add_18__19 ;
    input d_arr_add_18__18 ;
    input d_arr_add_18__17 ;
    input d_arr_add_18__16 ;
    input d_arr_add_18__15 ;
    input d_arr_add_18__14 ;
    input d_arr_add_18__13 ;
    input d_arr_add_18__12 ;
    input d_arr_add_18__11 ;
    input d_arr_add_18__10 ;
    input d_arr_add_18__9 ;
    input d_arr_add_18__8 ;
    input d_arr_add_18__7 ;
    input d_arr_add_18__6 ;
    input d_arr_add_18__5 ;
    input d_arr_add_18__4 ;
    input d_arr_add_18__3 ;
    input d_arr_add_18__2 ;
    input d_arr_add_18__1 ;
    input d_arr_add_18__0 ;
    input d_arr_add_19__31 ;
    input d_arr_add_19__30 ;
    input d_arr_add_19__29 ;
    input d_arr_add_19__28 ;
    input d_arr_add_19__27 ;
    input d_arr_add_19__26 ;
    input d_arr_add_19__25 ;
    input d_arr_add_19__24 ;
    input d_arr_add_19__23 ;
    input d_arr_add_19__22 ;
    input d_arr_add_19__21 ;
    input d_arr_add_19__20 ;
    input d_arr_add_19__19 ;
    input d_arr_add_19__18 ;
    input d_arr_add_19__17 ;
    input d_arr_add_19__16 ;
    input d_arr_add_19__15 ;
    input d_arr_add_19__14 ;
    input d_arr_add_19__13 ;
    input d_arr_add_19__12 ;
    input d_arr_add_19__11 ;
    input d_arr_add_19__10 ;
    input d_arr_add_19__9 ;
    input d_arr_add_19__8 ;
    input d_arr_add_19__7 ;
    input d_arr_add_19__6 ;
    input d_arr_add_19__5 ;
    input d_arr_add_19__4 ;
    input d_arr_add_19__3 ;
    input d_arr_add_19__2 ;
    input d_arr_add_19__1 ;
    input d_arr_add_19__0 ;
    input d_arr_add_20__31 ;
    input d_arr_add_20__30 ;
    input d_arr_add_20__29 ;
    input d_arr_add_20__28 ;
    input d_arr_add_20__27 ;
    input d_arr_add_20__26 ;
    input d_arr_add_20__25 ;
    input d_arr_add_20__24 ;
    input d_arr_add_20__23 ;
    input d_arr_add_20__22 ;
    input d_arr_add_20__21 ;
    input d_arr_add_20__20 ;
    input d_arr_add_20__19 ;
    input d_arr_add_20__18 ;
    input d_arr_add_20__17 ;
    input d_arr_add_20__16 ;
    input d_arr_add_20__15 ;
    input d_arr_add_20__14 ;
    input d_arr_add_20__13 ;
    input d_arr_add_20__12 ;
    input d_arr_add_20__11 ;
    input d_arr_add_20__10 ;
    input d_arr_add_20__9 ;
    input d_arr_add_20__8 ;
    input d_arr_add_20__7 ;
    input d_arr_add_20__6 ;
    input d_arr_add_20__5 ;
    input d_arr_add_20__4 ;
    input d_arr_add_20__3 ;
    input d_arr_add_20__2 ;
    input d_arr_add_20__1 ;
    input d_arr_add_20__0 ;
    input d_arr_add_21__31 ;
    input d_arr_add_21__30 ;
    input d_arr_add_21__29 ;
    input d_arr_add_21__28 ;
    input d_arr_add_21__27 ;
    input d_arr_add_21__26 ;
    input d_arr_add_21__25 ;
    input d_arr_add_21__24 ;
    input d_arr_add_21__23 ;
    input d_arr_add_21__22 ;
    input d_arr_add_21__21 ;
    input d_arr_add_21__20 ;
    input d_arr_add_21__19 ;
    input d_arr_add_21__18 ;
    input d_arr_add_21__17 ;
    input d_arr_add_21__16 ;
    input d_arr_add_21__15 ;
    input d_arr_add_21__14 ;
    input d_arr_add_21__13 ;
    input d_arr_add_21__12 ;
    input d_arr_add_21__11 ;
    input d_arr_add_21__10 ;
    input d_arr_add_21__9 ;
    input d_arr_add_21__8 ;
    input d_arr_add_21__7 ;
    input d_arr_add_21__6 ;
    input d_arr_add_21__5 ;
    input d_arr_add_21__4 ;
    input d_arr_add_21__3 ;
    input d_arr_add_21__2 ;
    input d_arr_add_21__1 ;
    input d_arr_add_21__0 ;
    input d_arr_add_22__31 ;
    input d_arr_add_22__30 ;
    input d_arr_add_22__29 ;
    input d_arr_add_22__28 ;
    input d_arr_add_22__27 ;
    input d_arr_add_22__26 ;
    input d_arr_add_22__25 ;
    input d_arr_add_22__24 ;
    input d_arr_add_22__23 ;
    input d_arr_add_22__22 ;
    input d_arr_add_22__21 ;
    input d_arr_add_22__20 ;
    input d_arr_add_22__19 ;
    input d_arr_add_22__18 ;
    input d_arr_add_22__17 ;
    input d_arr_add_22__16 ;
    input d_arr_add_22__15 ;
    input d_arr_add_22__14 ;
    input d_arr_add_22__13 ;
    input d_arr_add_22__12 ;
    input d_arr_add_22__11 ;
    input d_arr_add_22__10 ;
    input d_arr_add_22__9 ;
    input d_arr_add_22__8 ;
    input d_arr_add_22__7 ;
    input d_arr_add_22__6 ;
    input d_arr_add_22__5 ;
    input d_arr_add_22__4 ;
    input d_arr_add_22__3 ;
    input d_arr_add_22__2 ;
    input d_arr_add_22__1 ;
    input d_arr_add_22__0 ;
    input d_arr_add_23__31 ;
    input d_arr_add_23__30 ;
    input d_arr_add_23__29 ;
    input d_arr_add_23__28 ;
    input d_arr_add_23__27 ;
    input d_arr_add_23__26 ;
    input d_arr_add_23__25 ;
    input d_arr_add_23__24 ;
    input d_arr_add_23__23 ;
    input d_arr_add_23__22 ;
    input d_arr_add_23__21 ;
    input d_arr_add_23__20 ;
    input d_arr_add_23__19 ;
    input d_arr_add_23__18 ;
    input d_arr_add_23__17 ;
    input d_arr_add_23__16 ;
    input d_arr_add_23__15 ;
    input d_arr_add_23__14 ;
    input d_arr_add_23__13 ;
    input d_arr_add_23__12 ;
    input d_arr_add_23__11 ;
    input d_arr_add_23__10 ;
    input d_arr_add_23__9 ;
    input d_arr_add_23__8 ;
    input d_arr_add_23__7 ;
    input d_arr_add_23__6 ;
    input d_arr_add_23__5 ;
    input d_arr_add_23__4 ;
    input d_arr_add_23__3 ;
    input d_arr_add_23__2 ;
    input d_arr_add_23__1 ;
    input d_arr_add_23__0 ;
    input d_arr_add_24__31 ;
    input d_arr_add_24__30 ;
    input d_arr_add_24__29 ;
    input d_arr_add_24__28 ;
    input d_arr_add_24__27 ;
    input d_arr_add_24__26 ;
    input d_arr_add_24__25 ;
    input d_arr_add_24__24 ;
    input d_arr_add_24__23 ;
    input d_arr_add_24__22 ;
    input d_arr_add_24__21 ;
    input d_arr_add_24__20 ;
    input d_arr_add_24__19 ;
    input d_arr_add_24__18 ;
    input d_arr_add_24__17 ;
    input d_arr_add_24__16 ;
    input d_arr_add_24__15 ;
    input d_arr_add_24__14 ;
    input d_arr_add_24__13 ;
    input d_arr_add_24__12 ;
    input d_arr_add_24__11 ;
    input d_arr_add_24__10 ;
    input d_arr_add_24__9 ;
    input d_arr_add_24__8 ;
    input d_arr_add_24__7 ;
    input d_arr_add_24__6 ;
    input d_arr_add_24__5 ;
    input d_arr_add_24__4 ;
    input d_arr_add_24__3 ;
    input d_arr_add_24__2 ;
    input d_arr_add_24__1 ;
    input d_arr_add_24__0 ;
    input d_arr_merge1_0__31 ;
    input d_arr_merge1_0__30 ;
    input d_arr_merge1_0__29 ;
    input d_arr_merge1_0__28 ;
    input d_arr_merge1_0__27 ;
    input d_arr_merge1_0__26 ;
    input d_arr_merge1_0__25 ;
    input d_arr_merge1_0__24 ;
    input d_arr_merge1_0__23 ;
    input d_arr_merge1_0__22 ;
    input d_arr_merge1_0__21 ;
    input d_arr_merge1_0__20 ;
    input d_arr_merge1_0__19 ;
    input d_arr_merge1_0__18 ;
    input d_arr_merge1_0__17 ;
    input d_arr_merge1_0__16 ;
    input d_arr_merge1_0__15 ;
    input d_arr_merge1_0__14 ;
    input d_arr_merge1_0__13 ;
    input d_arr_merge1_0__12 ;
    input d_arr_merge1_0__11 ;
    input d_arr_merge1_0__10 ;
    input d_arr_merge1_0__9 ;
    input d_arr_merge1_0__8 ;
    input d_arr_merge1_0__7 ;
    input d_arr_merge1_0__6 ;
    input d_arr_merge1_0__5 ;
    input d_arr_merge1_0__4 ;
    input d_arr_merge1_0__3 ;
    input d_arr_merge1_0__2 ;
    input d_arr_merge1_0__1 ;
    input d_arr_merge1_0__0 ;
    input d_arr_merge1_1__31 ;
    input d_arr_merge1_1__30 ;
    input d_arr_merge1_1__29 ;
    input d_arr_merge1_1__28 ;
    input d_arr_merge1_1__27 ;
    input d_arr_merge1_1__26 ;
    input d_arr_merge1_1__25 ;
    input d_arr_merge1_1__24 ;
    input d_arr_merge1_1__23 ;
    input d_arr_merge1_1__22 ;
    input d_arr_merge1_1__21 ;
    input d_arr_merge1_1__20 ;
    input d_arr_merge1_1__19 ;
    input d_arr_merge1_1__18 ;
    input d_arr_merge1_1__17 ;
    input d_arr_merge1_1__16 ;
    input d_arr_merge1_1__15 ;
    input d_arr_merge1_1__14 ;
    input d_arr_merge1_1__13 ;
    input d_arr_merge1_1__12 ;
    input d_arr_merge1_1__11 ;
    input d_arr_merge1_1__10 ;
    input d_arr_merge1_1__9 ;
    input d_arr_merge1_1__8 ;
    input d_arr_merge1_1__7 ;
    input d_arr_merge1_1__6 ;
    input d_arr_merge1_1__5 ;
    input d_arr_merge1_1__4 ;
    input d_arr_merge1_1__3 ;
    input d_arr_merge1_1__2 ;
    input d_arr_merge1_1__1 ;
    input d_arr_merge1_1__0 ;
    input d_arr_merge1_2__31 ;
    input d_arr_merge1_2__30 ;
    input d_arr_merge1_2__29 ;
    input d_arr_merge1_2__28 ;
    input d_arr_merge1_2__27 ;
    input d_arr_merge1_2__26 ;
    input d_arr_merge1_2__25 ;
    input d_arr_merge1_2__24 ;
    input d_arr_merge1_2__23 ;
    input d_arr_merge1_2__22 ;
    input d_arr_merge1_2__21 ;
    input d_arr_merge1_2__20 ;
    input d_arr_merge1_2__19 ;
    input d_arr_merge1_2__18 ;
    input d_arr_merge1_2__17 ;
    input d_arr_merge1_2__16 ;
    input d_arr_merge1_2__15 ;
    input d_arr_merge1_2__14 ;
    input d_arr_merge1_2__13 ;
    input d_arr_merge1_2__12 ;
    input d_arr_merge1_2__11 ;
    input d_arr_merge1_2__10 ;
    input d_arr_merge1_2__9 ;
    input d_arr_merge1_2__8 ;
    input d_arr_merge1_2__7 ;
    input d_arr_merge1_2__6 ;
    input d_arr_merge1_2__5 ;
    input d_arr_merge1_2__4 ;
    input d_arr_merge1_2__3 ;
    input d_arr_merge1_2__2 ;
    input d_arr_merge1_2__1 ;
    input d_arr_merge1_2__0 ;
    input d_arr_merge1_3__31 ;
    input d_arr_merge1_3__30 ;
    input d_arr_merge1_3__29 ;
    input d_arr_merge1_3__28 ;
    input d_arr_merge1_3__27 ;
    input d_arr_merge1_3__26 ;
    input d_arr_merge1_3__25 ;
    input d_arr_merge1_3__24 ;
    input d_arr_merge1_3__23 ;
    input d_arr_merge1_3__22 ;
    input d_arr_merge1_3__21 ;
    input d_arr_merge1_3__20 ;
    input d_arr_merge1_3__19 ;
    input d_arr_merge1_3__18 ;
    input d_arr_merge1_3__17 ;
    input d_arr_merge1_3__16 ;
    input d_arr_merge1_3__15 ;
    input d_arr_merge1_3__14 ;
    input d_arr_merge1_3__13 ;
    input d_arr_merge1_3__12 ;
    input d_arr_merge1_3__11 ;
    input d_arr_merge1_3__10 ;
    input d_arr_merge1_3__9 ;
    input d_arr_merge1_3__8 ;
    input d_arr_merge1_3__7 ;
    input d_arr_merge1_3__6 ;
    input d_arr_merge1_3__5 ;
    input d_arr_merge1_3__4 ;
    input d_arr_merge1_3__3 ;
    input d_arr_merge1_3__2 ;
    input d_arr_merge1_3__1 ;
    input d_arr_merge1_3__0 ;
    input d_arr_merge1_4__31 ;
    input d_arr_merge1_4__30 ;
    input d_arr_merge1_4__29 ;
    input d_arr_merge1_4__28 ;
    input d_arr_merge1_4__27 ;
    input d_arr_merge1_4__26 ;
    input d_arr_merge1_4__25 ;
    input d_arr_merge1_4__24 ;
    input d_arr_merge1_4__23 ;
    input d_arr_merge1_4__22 ;
    input d_arr_merge1_4__21 ;
    input d_arr_merge1_4__20 ;
    input d_arr_merge1_4__19 ;
    input d_arr_merge1_4__18 ;
    input d_arr_merge1_4__17 ;
    input d_arr_merge1_4__16 ;
    input d_arr_merge1_4__15 ;
    input d_arr_merge1_4__14 ;
    input d_arr_merge1_4__13 ;
    input d_arr_merge1_4__12 ;
    input d_arr_merge1_4__11 ;
    input d_arr_merge1_4__10 ;
    input d_arr_merge1_4__9 ;
    input d_arr_merge1_4__8 ;
    input d_arr_merge1_4__7 ;
    input d_arr_merge1_4__6 ;
    input d_arr_merge1_4__5 ;
    input d_arr_merge1_4__4 ;
    input d_arr_merge1_4__3 ;
    input d_arr_merge1_4__2 ;
    input d_arr_merge1_4__1 ;
    input d_arr_merge1_4__0 ;
    input d_arr_merge1_5__31 ;
    input d_arr_merge1_5__30 ;
    input d_arr_merge1_5__29 ;
    input d_arr_merge1_5__28 ;
    input d_arr_merge1_5__27 ;
    input d_arr_merge1_5__26 ;
    input d_arr_merge1_5__25 ;
    input d_arr_merge1_5__24 ;
    input d_arr_merge1_5__23 ;
    input d_arr_merge1_5__22 ;
    input d_arr_merge1_5__21 ;
    input d_arr_merge1_5__20 ;
    input d_arr_merge1_5__19 ;
    input d_arr_merge1_5__18 ;
    input d_arr_merge1_5__17 ;
    input d_arr_merge1_5__16 ;
    input d_arr_merge1_5__15 ;
    input d_arr_merge1_5__14 ;
    input d_arr_merge1_5__13 ;
    input d_arr_merge1_5__12 ;
    input d_arr_merge1_5__11 ;
    input d_arr_merge1_5__10 ;
    input d_arr_merge1_5__9 ;
    input d_arr_merge1_5__8 ;
    input d_arr_merge1_5__7 ;
    input d_arr_merge1_5__6 ;
    input d_arr_merge1_5__5 ;
    input d_arr_merge1_5__4 ;
    input d_arr_merge1_5__3 ;
    input d_arr_merge1_5__2 ;
    input d_arr_merge1_5__1 ;
    input d_arr_merge1_5__0 ;
    input d_arr_merge1_6__31 ;
    input d_arr_merge1_6__30 ;
    input d_arr_merge1_6__29 ;
    input d_arr_merge1_6__28 ;
    input d_arr_merge1_6__27 ;
    input d_arr_merge1_6__26 ;
    input d_arr_merge1_6__25 ;
    input d_arr_merge1_6__24 ;
    input d_arr_merge1_6__23 ;
    input d_arr_merge1_6__22 ;
    input d_arr_merge1_6__21 ;
    input d_arr_merge1_6__20 ;
    input d_arr_merge1_6__19 ;
    input d_arr_merge1_6__18 ;
    input d_arr_merge1_6__17 ;
    input d_arr_merge1_6__16 ;
    input d_arr_merge1_6__15 ;
    input d_arr_merge1_6__14 ;
    input d_arr_merge1_6__13 ;
    input d_arr_merge1_6__12 ;
    input d_arr_merge1_6__11 ;
    input d_arr_merge1_6__10 ;
    input d_arr_merge1_6__9 ;
    input d_arr_merge1_6__8 ;
    input d_arr_merge1_6__7 ;
    input d_arr_merge1_6__6 ;
    input d_arr_merge1_6__5 ;
    input d_arr_merge1_6__4 ;
    input d_arr_merge1_6__3 ;
    input d_arr_merge1_6__2 ;
    input d_arr_merge1_6__1 ;
    input d_arr_merge1_6__0 ;
    input d_arr_merge1_7__31 ;
    input d_arr_merge1_7__30 ;
    input d_arr_merge1_7__29 ;
    input d_arr_merge1_7__28 ;
    input d_arr_merge1_7__27 ;
    input d_arr_merge1_7__26 ;
    input d_arr_merge1_7__25 ;
    input d_arr_merge1_7__24 ;
    input d_arr_merge1_7__23 ;
    input d_arr_merge1_7__22 ;
    input d_arr_merge1_7__21 ;
    input d_arr_merge1_7__20 ;
    input d_arr_merge1_7__19 ;
    input d_arr_merge1_7__18 ;
    input d_arr_merge1_7__17 ;
    input d_arr_merge1_7__16 ;
    input d_arr_merge1_7__15 ;
    input d_arr_merge1_7__14 ;
    input d_arr_merge1_7__13 ;
    input d_arr_merge1_7__12 ;
    input d_arr_merge1_7__11 ;
    input d_arr_merge1_7__10 ;
    input d_arr_merge1_7__9 ;
    input d_arr_merge1_7__8 ;
    input d_arr_merge1_7__7 ;
    input d_arr_merge1_7__6 ;
    input d_arr_merge1_7__5 ;
    input d_arr_merge1_7__4 ;
    input d_arr_merge1_7__3 ;
    input d_arr_merge1_7__2 ;
    input d_arr_merge1_7__1 ;
    input d_arr_merge1_7__0 ;
    input d_arr_merge1_8__31 ;
    input d_arr_merge1_8__30 ;
    input d_arr_merge1_8__29 ;
    input d_arr_merge1_8__28 ;
    input d_arr_merge1_8__27 ;
    input d_arr_merge1_8__26 ;
    input d_arr_merge1_8__25 ;
    input d_arr_merge1_8__24 ;
    input d_arr_merge1_8__23 ;
    input d_arr_merge1_8__22 ;
    input d_arr_merge1_8__21 ;
    input d_arr_merge1_8__20 ;
    input d_arr_merge1_8__19 ;
    input d_arr_merge1_8__18 ;
    input d_arr_merge1_8__17 ;
    input d_arr_merge1_8__16 ;
    input d_arr_merge1_8__15 ;
    input d_arr_merge1_8__14 ;
    input d_arr_merge1_8__13 ;
    input d_arr_merge1_8__12 ;
    input d_arr_merge1_8__11 ;
    input d_arr_merge1_8__10 ;
    input d_arr_merge1_8__9 ;
    input d_arr_merge1_8__8 ;
    input d_arr_merge1_8__7 ;
    input d_arr_merge1_8__6 ;
    input d_arr_merge1_8__5 ;
    input d_arr_merge1_8__4 ;
    input d_arr_merge1_8__3 ;
    input d_arr_merge1_8__2 ;
    input d_arr_merge1_8__1 ;
    input d_arr_merge1_8__0 ;
    input d_arr_merge1_9__31 ;
    input d_arr_merge1_9__30 ;
    input d_arr_merge1_9__29 ;
    input d_arr_merge1_9__28 ;
    input d_arr_merge1_9__27 ;
    input d_arr_merge1_9__26 ;
    input d_arr_merge1_9__25 ;
    input d_arr_merge1_9__24 ;
    input d_arr_merge1_9__23 ;
    input d_arr_merge1_9__22 ;
    input d_arr_merge1_9__21 ;
    input d_arr_merge1_9__20 ;
    input d_arr_merge1_9__19 ;
    input d_arr_merge1_9__18 ;
    input d_arr_merge1_9__17 ;
    input d_arr_merge1_9__16 ;
    input d_arr_merge1_9__15 ;
    input d_arr_merge1_9__14 ;
    input d_arr_merge1_9__13 ;
    input d_arr_merge1_9__12 ;
    input d_arr_merge1_9__11 ;
    input d_arr_merge1_9__10 ;
    input d_arr_merge1_9__9 ;
    input d_arr_merge1_9__8 ;
    input d_arr_merge1_9__7 ;
    input d_arr_merge1_9__6 ;
    input d_arr_merge1_9__5 ;
    input d_arr_merge1_9__4 ;
    input d_arr_merge1_9__3 ;
    input d_arr_merge1_9__2 ;
    input d_arr_merge1_9__1 ;
    input d_arr_merge1_9__0 ;
    input d_arr_merge1_10__31 ;
    input d_arr_merge1_10__30 ;
    input d_arr_merge1_10__29 ;
    input d_arr_merge1_10__28 ;
    input d_arr_merge1_10__27 ;
    input d_arr_merge1_10__26 ;
    input d_arr_merge1_10__25 ;
    input d_arr_merge1_10__24 ;
    input d_arr_merge1_10__23 ;
    input d_arr_merge1_10__22 ;
    input d_arr_merge1_10__21 ;
    input d_arr_merge1_10__20 ;
    input d_arr_merge1_10__19 ;
    input d_arr_merge1_10__18 ;
    input d_arr_merge1_10__17 ;
    input d_arr_merge1_10__16 ;
    input d_arr_merge1_10__15 ;
    input d_arr_merge1_10__14 ;
    input d_arr_merge1_10__13 ;
    input d_arr_merge1_10__12 ;
    input d_arr_merge1_10__11 ;
    input d_arr_merge1_10__10 ;
    input d_arr_merge1_10__9 ;
    input d_arr_merge1_10__8 ;
    input d_arr_merge1_10__7 ;
    input d_arr_merge1_10__6 ;
    input d_arr_merge1_10__5 ;
    input d_arr_merge1_10__4 ;
    input d_arr_merge1_10__3 ;
    input d_arr_merge1_10__2 ;
    input d_arr_merge1_10__1 ;
    input d_arr_merge1_10__0 ;
    input d_arr_merge1_11__31 ;
    input d_arr_merge1_11__30 ;
    input d_arr_merge1_11__29 ;
    input d_arr_merge1_11__28 ;
    input d_arr_merge1_11__27 ;
    input d_arr_merge1_11__26 ;
    input d_arr_merge1_11__25 ;
    input d_arr_merge1_11__24 ;
    input d_arr_merge1_11__23 ;
    input d_arr_merge1_11__22 ;
    input d_arr_merge1_11__21 ;
    input d_arr_merge1_11__20 ;
    input d_arr_merge1_11__19 ;
    input d_arr_merge1_11__18 ;
    input d_arr_merge1_11__17 ;
    input d_arr_merge1_11__16 ;
    input d_arr_merge1_11__15 ;
    input d_arr_merge1_11__14 ;
    input d_arr_merge1_11__13 ;
    input d_arr_merge1_11__12 ;
    input d_arr_merge1_11__11 ;
    input d_arr_merge1_11__10 ;
    input d_arr_merge1_11__9 ;
    input d_arr_merge1_11__8 ;
    input d_arr_merge1_11__7 ;
    input d_arr_merge1_11__6 ;
    input d_arr_merge1_11__5 ;
    input d_arr_merge1_11__4 ;
    input d_arr_merge1_11__3 ;
    input d_arr_merge1_11__2 ;
    input d_arr_merge1_11__1 ;
    input d_arr_merge1_11__0 ;
    input d_arr_merge1_12__31 ;
    input d_arr_merge1_12__30 ;
    input d_arr_merge1_12__29 ;
    input d_arr_merge1_12__28 ;
    input d_arr_merge1_12__27 ;
    input d_arr_merge1_12__26 ;
    input d_arr_merge1_12__25 ;
    input d_arr_merge1_12__24 ;
    input d_arr_merge1_12__23 ;
    input d_arr_merge1_12__22 ;
    input d_arr_merge1_12__21 ;
    input d_arr_merge1_12__20 ;
    input d_arr_merge1_12__19 ;
    input d_arr_merge1_12__18 ;
    input d_arr_merge1_12__17 ;
    input d_arr_merge1_12__16 ;
    input d_arr_merge1_12__15 ;
    input d_arr_merge1_12__14 ;
    input d_arr_merge1_12__13 ;
    input d_arr_merge1_12__12 ;
    input d_arr_merge1_12__11 ;
    input d_arr_merge1_12__10 ;
    input d_arr_merge1_12__9 ;
    input d_arr_merge1_12__8 ;
    input d_arr_merge1_12__7 ;
    input d_arr_merge1_12__6 ;
    input d_arr_merge1_12__5 ;
    input d_arr_merge1_12__4 ;
    input d_arr_merge1_12__3 ;
    input d_arr_merge1_12__2 ;
    input d_arr_merge1_12__1 ;
    input d_arr_merge1_12__0 ;
    input d_arr_merge1_13__31 ;
    input d_arr_merge1_13__30 ;
    input d_arr_merge1_13__29 ;
    input d_arr_merge1_13__28 ;
    input d_arr_merge1_13__27 ;
    input d_arr_merge1_13__26 ;
    input d_arr_merge1_13__25 ;
    input d_arr_merge1_13__24 ;
    input d_arr_merge1_13__23 ;
    input d_arr_merge1_13__22 ;
    input d_arr_merge1_13__21 ;
    input d_arr_merge1_13__20 ;
    input d_arr_merge1_13__19 ;
    input d_arr_merge1_13__18 ;
    input d_arr_merge1_13__17 ;
    input d_arr_merge1_13__16 ;
    input d_arr_merge1_13__15 ;
    input d_arr_merge1_13__14 ;
    input d_arr_merge1_13__13 ;
    input d_arr_merge1_13__12 ;
    input d_arr_merge1_13__11 ;
    input d_arr_merge1_13__10 ;
    input d_arr_merge1_13__9 ;
    input d_arr_merge1_13__8 ;
    input d_arr_merge1_13__7 ;
    input d_arr_merge1_13__6 ;
    input d_arr_merge1_13__5 ;
    input d_arr_merge1_13__4 ;
    input d_arr_merge1_13__3 ;
    input d_arr_merge1_13__2 ;
    input d_arr_merge1_13__1 ;
    input d_arr_merge1_13__0 ;
    input d_arr_merge1_14__31 ;
    input d_arr_merge1_14__30 ;
    input d_arr_merge1_14__29 ;
    input d_arr_merge1_14__28 ;
    input d_arr_merge1_14__27 ;
    input d_arr_merge1_14__26 ;
    input d_arr_merge1_14__25 ;
    input d_arr_merge1_14__24 ;
    input d_arr_merge1_14__23 ;
    input d_arr_merge1_14__22 ;
    input d_arr_merge1_14__21 ;
    input d_arr_merge1_14__20 ;
    input d_arr_merge1_14__19 ;
    input d_arr_merge1_14__18 ;
    input d_arr_merge1_14__17 ;
    input d_arr_merge1_14__16 ;
    input d_arr_merge1_14__15 ;
    input d_arr_merge1_14__14 ;
    input d_arr_merge1_14__13 ;
    input d_arr_merge1_14__12 ;
    input d_arr_merge1_14__11 ;
    input d_arr_merge1_14__10 ;
    input d_arr_merge1_14__9 ;
    input d_arr_merge1_14__8 ;
    input d_arr_merge1_14__7 ;
    input d_arr_merge1_14__6 ;
    input d_arr_merge1_14__5 ;
    input d_arr_merge1_14__4 ;
    input d_arr_merge1_14__3 ;
    input d_arr_merge1_14__2 ;
    input d_arr_merge1_14__1 ;
    input d_arr_merge1_14__0 ;
    input d_arr_merge1_15__31 ;
    input d_arr_merge1_15__30 ;
    input d_arr_merge1_15__29 ;
    input d_arr_merge1_15__28 ;
    input d_arr_merge1_15__27 ;
    input d_arr_merge1_15__26 ;
    input d_arr_merge1_15__25 ;
    input d_arr_merge1_15__24 ;
    input d_arr_merge1_15__23 ;
    input d_arr_merge1_15__22 ;
    input d_arr_merge1_15__21 ;
    input d_arr_merge1_15__20 ;
    input d_arr_merge1_15__19 ;
    input d_arr_merge1_15__18 ;
    input d_arr_merge1_15__17 ;
    input d_arr_merge1_15__16 ;
    input d_arr_merge1_15__15 ;
    input d_arr_merge1_15__14 ;
    input d_arr_merge1_15__13 ;
    input d_arr_merge1_15__12 ;
    input d_arr_merge1_15__11 ;
    input d_arr_merge1_15__10 ;
    input d_arr_merge1_15__9 ;
    input d_arr_merge1_15__8 ;
    input d_arr_merge1_15__7 ;
    input d_arr_merge1_15__6 ;
    input d_arr_merge1_15__5 ;
    input d_arr_merge1_15__4 ;
    input d_arr_merge1_15__3 ;
    input d_arr_merge1_15__2 ;
    input d_arr_merge1_15__1 ;
    input d_arr_merge1_15__0 ;
    input d_arr_merge1_16__31 ;
    input d_arr_merge1_16__30 ;
    input d_arr_merge1_16__29 ;
    input d_arr_merge1_16__28 ;
    input d_arr_merge1_16__27 ;
    input d_arr_merge1_16__26 ;
    input d_arr_merge1_16__25 ;
    input d_arr_merge1_16__24 ;
    input d_arr_merge1_16__23 ;
    input d_arr_merge1_16__22 ;
    input d_arr_merge1_16__21 ;
    input d_arr_merge1_16__20 ;
    input d_arr_merge1_16__19 ;
    input d_arr_merge1_16__18 ;
    input d_arr_merge1_16__17 ;
    input d_arr_merge1_16__16 ;
    input d_arr_merge1_16__15 ;
    input d_arr_merge1_16__14 ;
    input d_arr_merge1_16__13 ;
    input d_arr_merge1_16__12 ;
    input d_arr_merge1_16__11 ;
    input d_arr_merge1_16__10 ;
    input d_arr_merge1_16__9 ;
    input d_arr_merge1_16__8 ;
    input d_arr_merge1_16__7 ;
    input d_arr_merge1_16__6 ;
    input d_arr_merge1_16__5 ;
    input d_arr_merge1_16__4 ;
    input d_arr_merge1_16__3 ;
    input d_arr_merge1_16__2 ;
    input d_arr_merge1_16__1 ;
    input d_arr_merge1_16__0 ;
    input d_arr_merge1_17__31 ;
    input d_arr_merge1_17__30 ;
    input d_arr_merge1_17__29 ;
    input d_arr_merge1_17__28 ;
    input d_arr_merge1_17__27 ;
    input d_arr_merge1_17__26 ;
    input d_arr_merge1_17__25 ;
    input d_arr_merge1_17__24 ;
    input d_arr_merge1_17__23 ;
    input d_arr_merge1_17__22 ;
    input d_arr_merge1_17__21 ;
    input d_arr_merge1_17__20 ;
    input d_arr_merge1_17__19 ;
    input d_arr_merge1_17__18 ;
    input d_arr_merge1_17__17 ;
    input d_arr_merge1_17__16 ;
    input d_arr_merge1_17__15 ;
    input d_arr_merge1_17__14 ;
    input d_arr_merge1_17__13 ;
    input d_arr_merge1_17__12 ;
    input d_arr_merge1_17__11 ;
    input d_arr_merge1_17__10 ;
    input d_arr_merge1_17__9 ;
    input d_arr_merge1_17__8 ;
    input d_arr_merge1_17__7 ;
    input d_arr_merge1_17__6 ;
    input d_arr_merge1_17__5 ;
    input d_arr_merge1_17__4 ;
    input d_arr_merge1_17__3 ;
    input d_arr_merge1_17__2 ;
    input d_arr_merge1_17__1 ;
    input d_arr_merge1_17__0 ;
    input d_arr_merge1_18__31 ;
    input d_arr_merge1_18__30 ;
    input d_arr_merge1_18__29 ;
    input d_arr_merge1_18__28 ;
    input d_arr_merge1_18__27 ;
    input d_arr_merge1_18__26 ;
    input d_arr_merge1_18__25 ;
    input d_arr_merge1_18__24 ;
    input d_arr_merge1_18__23 ;
    input d_arr_merge1_18__22 ;
    input d_arr_merge1_18__21 ;
    input d_arr_merge1_18__20 ;
    input d_arr_merge1_18__19 ;
    input d_arr_merge1_18__18 ;
    input d_arr_merge1_18__17 ;
    input d_arr_merge1_18__16 ;
    input d_arr_merge1_18__15 ;
    input d_arr_merge1_18__14 ;
    input d_arr_merge1_18__13 ;
    input d_arr_merge1_18__12 ;
    input d_arr_merge1_18__11 ;
    input d_arr_merge1_18__10 ;
    input d_arr_merge1_18__9 ;
    input d_arr_merge1_18__8 ;
    input d_arr_merge1_18__7 ;
    input d_arr_merge1_18__6 ;
    input d_arr_merge1_18__5 ;
    input d_arr_merge1_18__4 ;
    input d_arr_merge1_18__3 ;
    input d_arr_merge1_18__2 ;
    input d_arr_merge1_18__1 ;
    input d_arr_merge1_18__0 ;
    input d_arr_merge1_19__31 ;
    input d_arr_merge1_19__30 ;
    input d_arr_merge1_19__29 ;
    input d_arr_merge1_19__28 ;
    input d_arr_merge1_19__27 ;
    input d_arr_merge1_19__26 ;
    input d_arr_merge1_19__25 ;
    input d_arr_merge1_19__24 ;
    input d_arr_merge1_19__23 ;
    input d_arr_merge1_19__22 ;
    input d_arr_merge1_19__21 ;
    input d_arr_merge1_19__20 ;
    input d_arr_merge1_19__19 ;
    input d_arr_merge1_19__18 ;
    input d_arr_merge1_19__17 ;
    input d_arr_merge1_19__16 ;
    input d_arr_merge1_19__15 ;
    input d_arr_merge1_19__14 ;
    input d_arr_merge1_19__13 ;
    input d_arr_merge1_19__12 ;
    input d_arr_merge1_19__11 ;
    input d_arr_merge1_19__10 ;
    input d_arr_merge1_19__9 ;
    input d_arr_merge1_19__8 ;
    input d_arr_merge1_19__7 ;
    input d_arr_merge1_19__6 ;
    input d_arr_merge1_19__5 ;
    input d_arr_merge1_19__4 ;
    input d_arr_merge1_19__3 ;
    input d_arr_merge1_19__2 ;
    input d_arr_merge1_19__1 ;
    input d_arr_merge1_19__0 ;
    input d_arr_merge1_20__31 ;
    input d_arr_merge1_20__30 ;
    input d_arr_merge1_20__29 ;
    input d_arr_merge1_20__28 ;
    input d_arr_merge1_20__27 ;
    input d_arr_merge1_20__26 ;
    input d_arr_merge1_20__25 ;
    input d_arr_merge1_20__24 ;
    input d_arr_merge1_20__23 ;
    input d_arr_merge1_20__22 ;
    input d_arr_merge1_20__21 ;
    input d_arr_merge1_20__20 ;
    input d_arr_merge1_20__19 ;
    input d_arr_merge1_20__18 ;
    input d_arr_merge1_20__17 ;
    input d_arr_merge1_20__16 ;
    input d_arr_merge1_20__15 ;
    input d_arr_merge1_20__14 ;
    input d_arr_merge1_20__13 ;
    input d_arr_merge1_20__12 ;
    input d_arr_merge1_20__11 ;
    input d_arr_merge1_20__10 ;
    input d_arr_merge1_20__9 ;
    input d_arr_merge1_20__8 ;
    input d_arr_merge1_20__7 ;
    input d_arr_merge1_20__6 ;
    input d_arr_merge1_20__5 ;
    input d_arr_merge1_20__4 ;
    input d_arr_merge1_20__3 ;
    input d_arr_merge1_20__2 ;
    input d_arr_merge1_20__1 ;
    input d_arr_merge1_20__0 ;
    input d_arr_merge1_21__31 ;
    input d_arr_merge1_21__30 ;
    input d_arr_merge1_21__29 ;
    input d_arr_merge1_21__28 ;
    input d_arr_merge1_21__27 ;
    input d_arr_merge1_21__26 ;
    input d_arr_merge1_21__25 ;
    input d_arr_merge1_21__24 ;
    input d_arr_merge1_21__23 ;
    input d_arr_merge1_21__22 ;
    input d_arr_merge1_21__21 ;
    input d_arr_merge1_21__20 ;
    input d_arr_merge1_21__19 ;
    input d_arr_merge1_21__18 ;
    input d_arr_merge1_21__17 ;
    input d_arr_merge1_21__16 ;
    input d_arr_merge1_21__15 ;
    input d_arr_merge1_21__14 ;
    input d_arr_merge1_21__13 ;
    input d_arr_merge1_21__12 ;
    input d_arr_merge1_21__11 ;
    input d_arr_merge1_21__10 ;
    input d_arr_merge1_21__9 ;
    input d_arr_merge1_21__8 ;
    input d_arr_merge1_21__7 ;
    input d_arr_merge1_21__6 ;
    input d_arr_merge1_21__5 ;
    input d_arr_merge1_21__4 ;
    input d_arr_merge1_21__3 ;
    input d_arr_merge1_21__2 ;
    input d_arr_merge1_21__1 ;
    input d_arr_merge1_21__0 ;
    input d_arr_merge1_22__31 ;
    input d_arr_merge1_22__30 ;
    input d_arr_merge1_22__29 ;
    input d_arr_merge1_22__28 ;
    input d_arr_merge1_22__27 ;
    input d_arr_merge1_22__26 ;
    input d_arr_merge1_22__25 ;
    input d_arr_merge1_22__24 ;
    input d_arr_merge1_22__23 ;
    input d_arr_merge1_22__22 ;
    input d_arr_merge1_22__21 ;
    input d_arr_merge1_22__20 ;
    input d_arr_merge1_22__19 ;
    input d_arr_merge1_22__18 ;
    input d_arr_merge1_22__17 ;
    input d_arr_merge1_22__16 ;
    input d_arr_merge1_22__15 ;
    input d_arr_merge1_22__14 ;
    input d_arr_merge1_22__13 ;
    input d_arr_merge1_22__12 ;
    input d_arr_merge1_22__11 ;
    input d_arr_merge1_22__10 ;
    input d_arr_merge1_22__9 ;
    input d_arr_merge1_22__8 ;
    input d_arr_merge1_22__7 ;
    input d_arr_merge1_22__6 ;
    input d_arr_merge1_22__5 ;
    input d_arr_merge1_22__4 ;
    input d_arr_merge1_22__3 ;
    input d_arr_merge1_22__2 ;
    input d_arr_merge1_22__1 ;
    input d_arr_merge1_22__0 ;
    input d_arr_merge1_23__31 ;
    input d_arr_merge1_23__30 ;
    input d_arr_merge1_23__29 ;
    input d_arr_merge1_23__28 ;
    input d_arr_merge1_23__27 ;
    input d_arr_merge1_23__26 ;
    input d_arr_merge1_23__25 ;
    input d_arr_merge1_23__24 ;
    input d_arr_merge1_23__23 ;
    input d_arr_merge1_23__22 ;
    input d_arr_merge1_23__21 ;
    input d_arr_merge1_23__20 ;
    input d_arr_merge1_23__19 ;
    input d_arr_merge1_23__18 ;
    input d_arr_merge1_23__17 ;
    input d_arr_merge1_23__16 ;
    input d_arr_merge1_23__15 ;
    input d_arr_merge1_23__14 ;
    input d_arr_merge1_23__13 ;
    input d_arr_merge1_23__12 ;
    input d_arr_merge1_23__11 ;
    input d_arr_merge1_23__10 ;
    input d_arr_merge1_23__9 ;
    input d_arr_merge1_23__8 ;
    input d_arr_merge1_23__7 ;
    input d_arr_merge1_23__6 ;
    input d_arr_merge1_23__5 ;
    input d_arr_merge1_23__4 ;
    input d_arr_merge1_23__3 ;
    input d_arr_merge1_23__2 ;
    input d_arr_merge1_23__1 ;
    input d_arr_merge1_23__0 ;
    input d_arr_merge1_24__31 ;
    input d_arr_merge1_24__30 ;
    input d_arr_merge1_24__29 ;
    input d_arr_merge1_24__28 ;
    input d_arr_merge1_24__27 ;
    input d_arr_merge1_24__26 ;
    input d_arr_merge1_24__25 ;
    input d_arr_merge1_24__24 ;
    input d_arr_merge1_24__23 ;
    input d_arr_merge1_24__22 ;
    input d_arr_merge1_24__21 ;
    input d_arr_merge1_24__20 ;
    input d_arr_merge1_24__19 ;
    input d_arr_merge1_24__18 ;
    input d_arr_merge1_24__17 ;
    input d_arr_merge1_24__16 ;
    input d_arr_merge1_24__15 ;
    input d_arr_merge1_24__14 ;
    input d_arr_merge1_24__13 ;
    input d_arr_merge1_24__12 ;
    input d_arr_merge1_24__11 ;
    input d_arr_merge1_24__10 ;
    input d_arr_merge1_24__9 ;
    input d_arr_merge1_24__8 ;
    input d_arr_merge1_24__7 ;
    input d_arr_merge1_24__6 ;
    input d_arr_merge1_24__5 ;
    input d_arr_merge1_24__4 ;
    input d_arr_merge1_24__3 ;
    input d_arr_merge1_24__2 ;
    input d_arr_merge1_24__1 ;
    input d_arr_merge1_24__0 ;
    input d_arr_merge2_0__31 ;
    input d_arr_merge2_0__30 ;
    input d_arr_merge2_0__29 ;
    input d_arr_merge2_0__28 ;
    input d_arr_merge2_0__27 ;
    input d_arr_merge2_0__26 ;
    input d_arr_merge2_0__25 ;
    input d_arr_merge2_0__24 ;
    input d_arr_merge2_0__23 ;
    input d_arr_merge2_0__22 ;
    input d_arr_merge2_0__21 ;
    input d_arr_merge2_0__20 ;
    input d_arr_merge2_0__19 ;
    input d_arr_merge2_0__18 ;
    input d_arr_merge2_0__17 ;
    input d_arr_merge2_0__16 ;
    input d_arr_merge2_0__15 ;
    input d_arr_merge2_0__14 ;
    input d_arr_merge2_0__13 ;
    input d_arr_merge2_0__12 ;
    input d_arr_merge2_0__11 ;
    input d_arr_merge2_0__10 ;
    input d_arr_merge2_0__9 ;
    input d_arr_merge2_0__8 ;
    input d_arr_merge2_0__7 ;
    input d_arr_merge2_0__6 ;
    input d_arr_merge2_0__5 ;
    input d_arr_merge2_0__4 ;
    input d_arr_merge2_0__3 ;
    input d_arr_merge2_0__2 ;
    input d_arr_merge2_0__1 ;
    input d_arr_merge2_0__0 ;
    input d_arr_merge2_1__31 ;
    input d_arr_merge2_1__30 ;
    input d_arr_merge2_1__29 ;
    input d_arr_merge2_1__28 ;
    input d_arr_merge2_1__27 ;
    input d_arr_merge2_1__26 ;
    input d_arr_merge2_1__25 ;
    input d_arr_merge2_1__24 ;
    input d_arr_merge2_1__23 ;
    input d_arr_merge2_1__22 ;
    input d_arr_merge2_1__21 ;
    input d_arr_merge2_1__20 ;
    input d_arr_merge2_1__19 ;
    input d_arr_merge2_1__18 ;
    input d_arr_merge2_1__17 ;
    input d_arr_merge2_1__16 ;
    input d_arr_merge2_1__15 ;
    input d_arr_merge2_1__14 ;
    input d_arr_merge2_1__13 ;
    input d_arr_merge2_1__12 ;
    input d_arr_merge2_1__11 ;
    input d_arr_merge2_1__10 ;
    input d_arr_merge2_1__9 ;
    input d_arr_merge2_1__8 ;
    input d_arr_merge2_1__7 ;
    input d_arr_merge2_1__6 ;
    input d_arr_merge2_1__5 ;
    input d_arr_merge2_1__4 ;
    input d_arr_merge2_1__3 ;
    input d_arr_merge2_1__2 ;
    input d_arr_merge2_1__1 ;
    input d_arr_merge2_1__0 ;
    input d_arr_merge2_2__31 ;
    input d_arr_merge2_2__30 ;
    input d_arr_merge2_2__29 ;
    input d_arr_merge2_2__28 ;
    input d_arr_merge2_2__27 ;
    input d_arr_merge2_2__26 ;
    input d_arr_merge2_2__25 ;
    input d_arr_merge2_2__24 ;
    input d_arr_merge2_2__23 ;
    input d_arr_merge2_2__22 ;
    input d_arr_merge2_2__21 ;
    input d_arr_merge2_2__20 ;
    input d_arr_merge2_2__19 ;
    input d_arr_merge2_2__18 ;
    input d_arr_merge2_2__17 ;
    input d_arr_merge2_2__16 ;
    input d_arr_merge2_2__15 ;
    input d_arr_merge2_2__14 ;
    input d_arr_merge2_2__13 ;
    input d_arr_merge2_2__12 ;
    input d_arr_merge2_2__11 ;
    input d_arr_merge2_2__10 ;
    input d_arr_merge2_2__9 ;
    input d_arr_merge2_2__8 ;
    input d_arr_merge2_2__7 ;
    input d_arr_merge2_2__6 ;
    input d_arr_merge2_2__5 ;
    input d_arr_merge2_2__4 ;
    input d_arr_merge2_2__3 ;
    input d_arr_merge2_2__2 ;
    input d_arr_merge2_2__1 ;
    input d_arr_merge2_2__0 ;
    input d_arr_merge2_3__31 ;
    input d_arr_merge2_3__30 ;
    input d_arr_merge2_3__29 ;
    input d_arr_merge2_3__28 ;
    input d_arr_merge2_3__27 ;
    input d_arr_merge2_3__26 ;
    input d_arr_merge2_3__25 ;
    input d_arr_merge2_3__24 ;
    input d_arr_merge2_3__23 ;
    input d_arr_merge2_3__22 ;
    input d_arr_merge2_3__21 ;
    input d_arr_merge2_3__20 ;
    input d_arr_merge2_3__19 ;
    input d_arr_merge2_3__18 ;
    input d_arr_merge2_3__17 ;
    input d_arr_merge2_3__16 ;
    input d_arr_merge2_3__15 ;
    input d_arr_merge2_3__14 ;
    input d_arr_merge2_3__13 ;
    input d_arr_merge2_3__12 ;
    input d_arr_merge2_3__11 ;
    input d_arr_merge2_3__10 ;
    input d_arr_merge2_3__9 ;
    input d_arr_merge2_3__8 ;
    input d_arr_merge2_3__7 ;
    input d_arr_merge2_3__6 ;
    input d_arr_merge2_3__5 ;
    input d_arr_merge2_3__4 ;
    input d_arr_merge2_3__3 ;
    input d_arr_merge2_3__2 ;
    input d_arr_merge2_3__1 ;
    input d_arr_merge2_3__0 ;
    input d_arr_merge2_4__31 ;
    input d_arr_merge2_4__30 ;
    input d_arr_merge2_4__29 ;
    input d_arr_merge2_4__28 ;
    input d_arr_merge2_4__27 ;
    input d_arr_merge2_4__26 ;
    input d_arr_merge2_4__25 ;
    input d_arr_merge2_4__24 ;
    input d_arr_merge2_4__23 ;
    input d_arr_merge2_4__22 ;
    input d_arr_merge2_4__21 ;
    input d_arr_merge2_4__20 ;
    input d_arr_merge2_4__19 ;
    input d_arr_merge2_4__18 ;
    input d_arr_merge2_4__17 ;
    input d_arr_merge2_4__16 ;
    input d_arr_merge2_4__15 ;
    input d_arr_merge2_4__14 ;
    input d_arr_merge2_4__13 ;
    input d_arr_merge2_4__12 ;
    input d_arr_merge2_4__11 ;
    input d_arr_merge2_4__10 ;
    input d_arr_merge2_4__9 ;
    input d_arr_merge2_4__8 ;
    input d_arr_merge2_4__7 ;
    input d_arr_merge2_4__6 ;
    input d_arr_merge2_4__5 ;
    input d_arr_merge2_4__4 ;
    input d_arr_merge2_4__3 ;
    input d_arr_merge2_4__2 ;
    input d_arr_merge2_4__1 ;
    input d_arr_merge2_4__0 ;
    input d_arr_merge2_5__31 ;
    input d_arr_merge2_5__30 ;
    input d_arr_merge2_5__29 ;
    input d_arr_merge2_5__28 ;
    input d_arr_merge2_5__27 ;
    input d_arr_merge2_5__26 ;
    input d_arr_merge2_5__25 ;
    input d_arr_merge2_5__24 ;
    input d_arr_merge2_5__23 ;
    input d_arr_merge2_5__22 ;
    input d_arr_merge2_5__21 ;
    input d_arr_merge2_5__20 ;
    input d_arr_merge2_5__19 ;
    input d_arr_merge2_5__18 ;
    input d_arr_merge2_5__17 ;
    input d_arr_merge2_5__16 ;
    input d_arr_merge2_5__15 ;
    input d_arr_merge2_5__14 ;
    input d_arr_merge2_5__13 ;
    input d_arr_merge2_5__12 ;
    input d_arr_merge2_5__11 ;
    input d_arr_merge2_5__10 ;
    input d_arr_merge2_5__9 ;
    input d_arr_merge2_5__8 ;
    input d_arr_merge2_5__7 ;
    input d_arr_merge2_5__6 ;
    input d_arr_merge2_5__5 ;
    input d_arr_merge2_5__4 ;
    input d_arr_merge2_5__3 ;
    input d_arr_merge2_5__2 ;
    input d_arr_merge2_5__1 ;
    input d_arr_merge2_5__0 ;
    input d_arr_merge2_6__31 ;
    input d_arr_merge2_6__30 ;
    input d_arr_merge2_6__29 ;
    input d_arr_merge2_6__28 ;
    input d_arr_merge2_6__27 ;
    input d_arr_merge2_6__26 ;
    input d_arr_merge2_6__25 ;
    input d_arr_merge2_6__24 ;
    input d_arr_merge2_6__23 ;
    input d_arr_merge2_6__22 ;
    input d_arr_merge2_6__21 ;
    input d_arr_merge2_6__20 ;
    input d_arr_merge2_6__19 ;
    input d_arr_merge2_6__18 ;
    input d_arr_merge2_6__17 ;
    input d_arr_merge2_6__16 ;
    input d_arr_merge2_6__15 ;
    input d_arr_merge2_6__14 ;
    input d_arr_merge2_6__13 ;
    input d_arr_merge2_6__12 ;
    input d_arr_merge2_6__11 ;
    input d_arr_merge2_6__10 ;
    input d_arr_merge2_6__9 ;
    input d_arr_merge2_6__8 ;
    input d_arr_merge2_6__7 ;
    input d_arr_merge2_6__6 ;
    input d_arr_merge2_6__5 ;
    input d_arr_merge2_6__4 ;
    input d_arr_merge2_6__3 ;
    input d_arr_merge2_6__2 ;
    input d_arr_merge2_6__1 ;
    input d_arr_merge2_6__0 ;
    input d_arr_merge2_7__31 ;
    input d_arr_merge2_7__30 ;
    input d_arr_merge2_7__29 ;
    input d_arr_merge2_7__28 ;
    input d_arr_merge2_7__27 ;
    input d_arr_merge2_7__26 ;
    input d_arr_merge2_7__25 ;
    input d_arr_merge2_7__24 ;
    input d_arr_merge2_7__23 ;
    input d_arr_merge2_7__22 ;
    input d_arr_merge2_7__21 ;
    input d_arr_merge2_7__20 ;
    input d_arr_merge2_7__19 ;
    input d_arr_merge2_7__18 ;
    input d_arr_merge2_7__17 ;
    input d_arr_merge2_7__16 ;
    input d_arr_merge2_7__15 ;
    input d_arr_merge2_7__14 ;
    input d_arr_merge2_7__13 ;
    input d_arr_merge2_7__12 ;
    input d_arr_merge2_7__11 ;
    input d_arr_merge2_7__10 ;
    input d_arr_merge2_7__9 ;
    input d_arr_merge2_7__8 ;
    input d_arr_merge2_7__7 ;
    input d_arr_merge2_7__6 ;
    input d_arr_merge2_7__5 ;
    input d_arr_merge2_7__4 ;
    input d_arr_merge2_7__3 ;
    input d_arr_merge2_7__2 ;
    input d_arr_merge2_7__1 ;
    input d_arr_merge2_7__0 ;
    input d_arr_merge2_8__31 ;
    input d_arr_merge2_8__30 ;
    input d_arr_merge2_8__29 ;
    input d_arr_merge2_8__28 ;
    input d_arr_merge2_8__27 ;
    input d_arr_merge2_8__26 ;
    input d_arr_merge2_8__25 ;
    input d_arr_merge2_8__24 ;
    input d_arr_merge2_8__23 ;
    input d_arr_merge2_8__22 ;
    input d_arr_merge2_8__21 ;
    input d_arr_merge2_8__20 ;
    input d_arr_merge2_8__19 ;
    input d_arr_merge2_8__18 ;
    input d_arr_merge2_8__17 ;
    input d_arr_merge2_8__16 ;
    input d_arr_merge2_8__15 ;
    input d_arr_merge2_8__14 ;
    input d_arr_merge2_8__13 ;
    input d_arr_merge2_8__12 ;
    input d_arr_merge2_8__11 ;
    input d_arr_merge2_8__10 ;
    input d_arr_merge2_8__9 ;
    input d_arr_merge2_8__8 ;
    input d_arr_merge2_8__7 ;
    input d_arr_merge2_8__6 ;
    input d_arr_merge2_8__5 ;
    input d_arr_merge2_8__4 ;
    input d_arr_merge2_8__3 ;
    input d_arr_merge2_8__2 ;
    input d_arr_merge2_8__1 ;
    input d_arr_merge2_8__0 ;
    input d_arr_merge2_9__31 ;
    input d_arr_merge2_9__30 ;
    input d_arr_merge2_9__29 ;
    input d_arr_merge2_9__28 ;
    input d_arr_merge2_9__27 ;
    input d_arr_merge2_9__26 ;
    input d_arr_merge2_9__25 ;
    input d_arr_merge2_9__24 ;
    input d_arr_merge2_9__23 ;
    input d_arr_merge2_9__22 ;
    input d_arr_merge2_9__21 ;
    input d_arr_merge2_9__20 ;
    input d_arr_merge2_9__19 ;
    input d_arr_merge2_9__18 ;
    input d_arr_merge2_9__17 ;
    input d_arr_merge2_9__16 ;
    input d_arr_merge2_9__15 ;
    input d_arr_merge2_9__14 ;
    input d_arr_merge2_9__13 ;
    input d_arr_merge2_9__12 ;
    input d_arr_merge2_9__11 ;
    input d_arr_merge2_9__10 ;
    input d_arr_merge2_9__9 ;
    input d_arr_merge2_9__8 ;
    input d_arr_merge2_9__7 ;
    input d_arr_merge2_9__6 ;
    input d_arr_merge2_9__5 ;
    input d_arr_merge2_9__4 ;
    input d_arr_merge2_9__3 ;
    input d_arr_merge2_9__2 ;
    input d_arr_merge2_9__1 ;
    input d_arr_merge2_9__0 ;
    input d_arr_merge2_10__31 ;
    input d_arr_merge2_10__30 ;
    input d_arr_merge2_10__29 ;
    input d_arr_merge2_10__28 ;
    input d_arr_merge2_10__27 ;
    input d_arr_merge2_10__26 ;
    input d_arr_merge2_10__25 ;
    input d_arr_merge2_10__24 ;
    input d_arr_merge2_10__23 ;
    input d_arr_merge2_10__22 ;
    input d_arr_merge2_10__21 ;
    input d_arr_merge2_10__20 ;
    input d_arr_merge2_10__19 ;
    input d_arr_merge2_10__18 ;
    input d_arr_merge2_10__17 ;
    input d_arr_merge2_10__16 ;
    input d_arr_merge2_10__15 ;
    input d_arr_merge2_10__14 ;
    input d_arr_merge2_10__13 ;
    input d_arr_merge2_10__12 ;
    input d_arr_merge2_10__11 ;
    input d_arr_merge2_10__10 ;
    input d_arr_merge2_10__9 ;
    input d_arr_merge2_10__8 ;
    input d_arr_merge2_10__7 ;
    input d_arr_merge2_10__6 ;
    input d_arr_merge2_10__5 ;
    input d_arr_merge2_10__4 ;
    input d_arr_merge2_10__3 ;
    input d_arr_merge2_10__2 ;
    input d_arr_merge2_10__1 ;
    input d_arr_merge2_10__0 ;
    input d_arr_merge2_11__31 ;
    input d_arr_merge2_11__30 ;
    input d_arr_merge2_11__29 ;
    input d_arr_merge2_11__28 ;
    input d_arr_merge2_11__27 ;
    input d_arr_merge2_11__26 ;
    input d_arr_merge2_11__25 ;
    input d_arr_merge2_11__24 ;
    input d_arr_merge2_11__23 ;
    input d_arr_merge2_11__22 ;
    input d_arr_merge2_11__21 ;
    input d_arr_merge2_11__20 ;
    input d_arr_merge2_11__19 ;
    input d_arr_merge2_11__18 ;
    input d_arr_merge2_11__17 ;
    input d_arr_merge2_11__16 ;
    input d_arr_merge2_11__15 ;
    input d_arr_merge2_11__14 ;
    input d_arr_merge2_11__13 ;
    input d_arr_merge2_11__12 ;
    input d_arr_merge2_11__11 ;
    input d_arr_merge2_11__10 ;
    input d_arr_merge2_11__9 ;
    input d_arr_merge2_11__8 ;
    input d_arr_merge2_11__7 ;
    input d_arr_merge2_11__6 ;
    input d_arr_merge2_11__5 ;
    input d_arr_merge2_11__4 ;
    input d_arr_merge2_11__3 ;
    input d_arr_merge2_11__2 ;
    input d_arr_merge2_11__1 ;
    input d_arr_merge2_11__0 ;
    input d_arr_merge2_12__31 ;
    input d_arr_merge2_12__30 ;
    input d_arr_merge2_12__29 ;
    input d_arr_merge2_12__28 ;
    input d_arr_merge2_12__27 ;
    input d_arr_merge2_12__26 ;
    input d_arr_merge2_12__25 ;
    input d_arr_merge2_12__24 ;
    input d_arr_merge2_12__23 ;
    input d_arr_merge2_12__22 ;
    input d_arr_merge2_12__21 ;
    input d_arr_merge2_12__20 ;
    input d_arr_merge2_12__19 ;
    input d_arr_merge2_12__18 ;
    input d_arr_merge2_12__17 ;
    input d_arr_merge2_12__16 ;
    input d_arr_merge2_12__15 ;
    input d_arr_merge2_12__14 ;
    input d_arr_merge2_12__13 ;
    input d_arr_merge2_12__12 ;
    input d_arr_merge2_12__11 ;
    input d_arr_merge2_12__10 ;
    input d_arr_merge2_12__9 ;
    input d_arr_merge2_12__8 ;
    input d_arr_merge2_12__7 ;
    input d_arr_merge2_12__6 ;
    input d_arr_merge2_12__5 ;
    input d_arr_merge2_12__4 ;
    input d_arr_merge2_12__3 ;
    input d_arr_merge2_12__2 ;
    input d_arr_merge2_12__1 ;
    input d_arr_merge2_12__0 ;
    input d_arr_merge2_13__31 ;
    input d_arr_merge2_13__30 ;
    input d_arr_merge2_13__29 ;
    input d_arr_merge2_13__28 ;
    input d_arr_merge2_13__27 ;
    input d_arr_merge2_13__26 ;
    input d_arr_merge2_13__25 ;
    input d_arr_merge2_13__24 ;
    input d_arr_merge2_13__23 ;
    input d_arr_merge2_13__22 ;
    input d_arr_merge2_13__21 ;
    input d_arr_merge2_13__20 ;
    input d_arr_merge2_13__19 ;
    input d_arr_merge2_13__18 ;
    input d_arr_merge2_13__17 ;
    input d_arr_merge2_13__16 ;
    input d_arr_merge2_13__15 ;
    input d_arr_merge2_13__14 ;
    input d_arr_merge2_13__13 ;
    input d_arr_merge2_13__12 ;
    input d_arr_merge2_13__11 ;
    input d_arr_merge2_13__10 ;
    input d_arr_merge2_13__9 ;
    input d_arr_merge2_13__8 ;
    input d_arr_merge2_13__7 ;
    input d_arr_merge2_13__6 ;
    input d_arr_merge2_13__5 ;
    input d_arr_merge2_13__4 ;
    input d_arr_merge2_13__3 ;
    input d_arr_merge2_13__2 ;
    input d_arr_merge2_13__1 ;
    input d_arr_merge2_13__0 ;
    input d_arr_merge2_14__31 ;
    input d_arr_merge2_14__30 ;
    input d_arr_merge2_14__29 ;
    input d_arr_merge2_14__28 ;
    input d_arr_merge2_14__27 ;
    input d_arr_merge2_14__26 ;
    input d_arr_merge2_14__25 ;
    input d_arr_merge2_14__24 ;
    input d_arr_merge2_14__23 ;
    input d_arr_merge2_14__22 ;
    input d_arr_merge2_14__21 ;
    input d_arr_merge2_14__20 ;
    input d_arr_merge2_14__19 ;
    input d_arr_merge2_14__18 ;
    input d_arr_merge2_14__17 ;
    input d_arr_merge2_14__16 ;
    input d_arr_merge2_14__15 ;
    input d_arr_merge2_14__14 ;
    input d_arr_merge2_14__13 ;
    input d_arr_merge2_14__12 ;
    input d_arr_merge2_14__11 ;
    input d_arr_merge2_14__10 ;
    input d_arr_merge2_14__9 ;
    input d_arr_merge2_14__8 ;
    input d_arr_merge2_14__7 ;
    input d_arr_merge2_14__6 ;
    input d_arr_merge2_14__5 ;
    input d_arr_merge2_14__4 ;
    input d_arr_merge2_14__3 ;
    input d_arr_merge2_14__2 ;
    input d_arr_merge2_14__1 ;
    input d_arr_merge2_14__0 ;
    input d_arr_merge2_15__31 ;
    input d_arr_merge2_15__30 ;
    input d_arr_merge2_15__29 ;
    input d_arr_merge2_15__28 ;
    input d_arr_merge2_15__27 ;
    input d_arr_merge2_15__26 ;
    input d_arr_merge2_15__25 ;
    input d_arr_merge2_15__24 ;
    input d_arr_merge2_15__23 ;
    input d_arr_merge2_15__22 ;
    input d_arr_merge2_15__21 ;
    input d_arr_merge2_15__20 ;
    input d_arr_merge2_15__19 ;
    input d_arr_merge2_15__18 ;
    input d_arr_merge2_15__17 ;
    input d_arr_merge2_15__16 ;
    input d_arr_merge2_15__15 ;
    input d_arr_merge2_15__14 ;
    input d_arr_merge2_15__13 ;
    input d_arr_merge2_15__12 ;
    input d_arr_merge2_15__11 ;
    input d_arr_merge2_15__10 ;
    input d_arr_merge2_15__9 ;
    input d_arr_merge2_15__8 ;
    input d_arr_merge2_15__7 ;
    input d_arr_merge2_15__6 ;
    input d_arr_merge2_15__5 ;
    input d_arr_merge2_15__4 ;
    input d_arr_merge2_15__3 ;
    input d_arr_merge2_15__2 ;
    input d_arr_merge2_15__1 ;
    input d_arr_merge2_15__0 ;
    input d_arr_merge2_16__31 ;
    input d_arr_merge2_16__30 ;
    input d_arr_merge2_16__29 ;
    input d_arr_merge2_16__28 ;
    input d_arr_merge2_16__27 ;
    input d_arr_merge2_16__26 ;
    input d_arr_merge2_16__25 ;
    input d_arr_merge2_16__24 ;
    input d_arr_merge2_16__23 ;
    input d_arr_merge2_16__22 ;
    input d_arr_merge2_16__21 ;
    input d_arr_merge2_16__20 ;
    input d_arr_merge2_16__19 ;
    input d_arr_merge2_16__18 ;
    input d_arr_merge2_16__17 ;
    input d_arr_merge2_16__16 ;
    input d_arr_merge2_16__15 ;
    input d_arr_merge2_16__14 ;
    input d_arr_merge2_16__13 ;
    input d_arr_merge2_16__12 ;
    input d_arr_merge2_16__11 ;
    input d_arr_merge2_16__10 ;
    input d_arr_merge2_16__9 ;
    input d_arr_merge2_16__8 ;
    input d_arr_merge2_16__7 ;
    input d_arr_merge2_16__6 ;
    input d_arr_merge2_16__5 ;
    input d_arr_merge2_16__4 ;
    input d_arr_merge2_16__3 ;
    input d_arr_merge2_16__2 ;
    input d_arr_merge2_16__1 ;
    input d_arr_merge2_16__0 ;
    input d_arr_merge2_17__31 ;
    input d_arr_merge2_17__30 ;
    input d_arr_merge2_17__29 ;
    input d_arr_merge2_17__28 ;
    input d_arr_merge2_17__27 ;
    input d_arr_merge2_17__26 ;
    input d_arr_merge2_17__25 ;
    input d_arr_merge2_17__24 ;
    input d_arr_merge2_17__23 ;
    input d_arr_merge2_17__22 ;
    input d_arr_merge2_17__21 ;
    input d_arr_merge2_17__20 ;
    input d_arr_merge2_17__19 ;
    input d_arr_merge2_17__18 ;
    input d_arr_merge2_17__17 ;
    input d_arr_merge2_17__16 ;
    input d_arr_merge2_17__15 ;
    input d_arr_merge2_17__14 ;
    input d_arr_merge2_17__13 ;
    input d_arr_merge2_17__12 ;
    input d_arr_merge2_17__11 ;
    input d_arr_merge2_17__10 ;
    input d_arr_merge2_17__9 ;
    input d_arr_merge2_17__8 ;
    input d_arr_merge2_17__7 ;
    input d_arr_merge2_17__6 ;
    input d_arr_merge2_17__5 ;
    input d_arr_merge2_17__4 ;
    input d_arr_merge2_17__3 ;
    input d_arr_merge2_17__2 ;
    input d_arr_merge2_17__1 ;
    input d_arr_merge2_17__0 ;
    input d_arr_merge2_18__31 ;
    input d_arr_merge2_18__30 ;
    input d_arr_merge2_18__29 ;
    input d_arr_merge2_18__28 ;
    input d_arr_merge2_18__27 ;
    input d_arr_merge2_18__26 ;
    input d_arr_merge2_18__25 ;
    input d_arr_merge2_18__24 ;
    input d_arr_merge2_18__23 ;
    input d_arr_merge2_18__22 ;
    input d_arr_merge2_18__21 ;
    input d_arr_merge2_18__20 ;
    input d_arr_merge2_18__19 ;
    input d_arr_merge2_18__18 ;
    input d_arr_merge2_18__17 ;
    input d_arr_merge2_18__16 ;
    input d_arr_merge2_18__15 ;
    input d_arr_merge2_18__14 ;
    input d_arr_merge2_18__13 ;
    input d_arr_merge2_18__12 ;
    input d_arr_merge2_18__11 ;
    input d_arr_merge2_18__10 ;
    input d_arr_merge2_18__9 ;
    input d_arr_merge2_18__8 ;
    input d_arr_merge2_18__7 ;
    input d_arr_merge2_18__6 ;
    input d_arr_merge2_18__5 ;
    input d_arr_merge2_18__4 ;
    input d_arr_merge2_18__3 ;
    input d_arr_merge2_18__2 ;
    input d_arr_merge2_18__1 ;
    input d_arr_merge2_18__0 ;
    input d_arr_merge2_19__31 ;
    input d_arr_merge2_19__30 ;
    input d_arr_merge2_19__29 ;
    input d_arr_merge2_19__28 ;
    input d_arr_merge2_19__27 ;
    input d_arr_merge2_19__26 ;
    input d_arr_merge2_19__25 ;
    input d_arr_merge2_19__24 ;
    input d_arr_merge2_19__23 ;
    input d_arr_merge2_19__22 ;
    input d_arr_merge2_19__21 ;
    input d_arr_merge2_19__20 ;
    input d_arr_merge2_19__19 ;
    input d_arr_merge2_19__18 ;
    input d_arr_merge2_19__17 ;
    input d_arr_merge2_19__16 ;
    input d_arr_merge2_19__15 ;
    input d_arr_merge2_19__14 ;
    input d_arr_merge2_19__13 ;
    input d_arr_merge2_19__12 ;
    input d_arr_merge2_19__11 ;
    input d_arr_merge2_19__10 ;
    input d_arr_merge2_19__9 ;
    input d_arr_merge2_19__8 ;
    input d_arr_merge2_19__7 ;
    input d_arr_merge2_19__6 ;
    input d_arr_merge2_19__5 ;
    input d_arr_merge2_19__4 ;
    input d_arr_merge2_19__3 ;
    input d_arr_merge2_19__2 ;
    input d_arr_merge2_19__1 ;
    input d_arr_merge2_19__0 ;
    input d_arr_merge2_20__31 ;
    input d_arr_merge2_20__30 ;
    input d_arr_merge2_20__29 ;
    input d_arr_merge2_20__28 ;
    input d_arr_merge2_20__27 ;
    input d_arr_merge2_20__26 ;
    input d_arr_merge2_20__25 ;
    input d_arr_merge2_20__24 ;
    input d_arr_merge2_20__23 ;
    input d_arr_merge2_20__22 ;
    input d_arr_merge2_20__21 ;
    input d_arr_merge2_20__20 ;
    input d_arr_merge2_20__19 ;
    input d_arr_merge2_20__18 ;
    input d_arr_merge2_20__17 ;
    input d_arr_merge2_20__16 ;
    input d_arr_merge2_20__15 ;
    input d_arr_merge2_20__14 ;
    input d_arr_merge2_20__13 ;
    input d_arr_merge2_20__12 ;
    input d_arr_merge2_20__11 ;
    input d_arr_merge2_20__10 ;
    input d_arr_merge2_20__9 ;
    input d_arr_merge2_20__8 ;
    input d_arr_merge2_20__7 ;
    input d_arr_merge2_20__6 ;
    input d_arr_merge2_20__5 ;
    input d_arr_merge2_20__4 ;
    input d_arr_merge2_20__3 ;
    input d_arr_merge2_20__2 ;
    input d_arr_merge2_20__1 ;
    input d_arr_merge2_20__0 ;
    input d_arr_merge2_21__31 ;
    input d_arr_merge2_21__30 ;
    input d_arr_merge2_21__29 ;
    input d_arr_merge2_21__28 ;
    input d_arr_merge2_21__27 ;
    input d_arr_merge2_21__26 ;
    input d_arr_merge2_21__25 ;
    input d_arr_merge2_21__24 ;
    input d_arr_merge2_21__23 ;
    input d_arr_merge2_21__22 ;
    input d_arr_merge2_21__21 ;
    input d_arr_merge2_21__20 ;
    input d_arr_merge2_21__19 ;
    input d_arr_merge2_21__18 ;
    input d_arr_merge2_21__17 ;
    input d_arr_merge2_21__16 ;
    input d_arr_merge2_21__15 ;
    input d_arr_merge2_21__14 ;
    input d_arr_merge2_21__13 ;
    input d_arr_merge2_21__12 ;
    input d_arr_merge2_21__11 ;
    input d_arr_merge2_21__10 ;
    input d_arr_merge2_21__9 ;
    input d_arr_merge2_21__8 ;
    input d_arr_merge2_21__7 ;
    input d_arr_merge2_21__6 ;
    input d_arr_merge2_21__5 ;
    input d_arr_merge2_21__4 ;
    input d_arr_merge2_21__3 ;
    input d_arr_merge2_21__2 ;
    input d_arr_merge2_21__1 ;
    input d_arr_merge2_21__0 ;
    input d_arr_merge2_22__31 ;
    input d_arr_merge2_22__30 ;
    input d_arr_merge2_22__29 ;
    input d_arr_merge2_22__28 ;
    input d_arr_merge2_22__27 ;
    input d_arr_merge2_22__26 ;
    input d_arr_merge2_22__25 ;
    input d_arr_merge2_22__24 ;
    input d_arr_merge2_22__23 ;
    input d_arr_merge2_22__22 ;
    input d_arr_merge2_22__21 ;
    input d_arr_merge2_22__20 ;
    input d_arr_merge2_22__19 ;
    input d_arr_merge2_22__18 ;
    input d_arr_merge2_22__17 ;
    input d_arr_merge2_22__16 ;
    input d_arr_merge2_22__15 ;
    input d_arr_merge2_22__14 ;
    input d_arr_merge2_22__13 ;
    input d_arr_merge2_22__12 ;
    input d_arr_merge2_22__11 ;
    input d_arr_merge2_22__10 ;
    input d_arr_merge2_22__9 ;
    input d_arr_merge2_22__8 ;
    input d_arr_merge2_22__7 ;
    input d_arr_merge2_22__6 ;
    input d_arr_merge2_22__5 ;
    input d_arr_merge2_22__4 ;
    input d_arr_merge2_22__3 ;
    input d_arr_merge2_22__2 ;
    input d_arr_merge2_22__1 ;
    input d_arr_merge2_22__0 ;
    input d_arr_merge2_23__31 ;
    input d_arr_merge2_23__30 ;
    input d_arr_merge2_23__29 ;
    input d_arr_merge2_23__28 ;
    input d_arr_merge2_23__27 ;
    input d_arr_merge2_23__26 ;
    input d_arr_merge2_23__25 ;
    input d_arr_merge2_23__24 ;
    input d_arr_merge2_23__23 ;
    input d_arr_merge2_23__22 ;
    input d_arr_merge2_23__21 ;
    input d_arr_merge2_23__20 ;
    input d_arr_merge2_23__19 ;
    input d_arr_merge2_23__18 ;
    input d_arr_merge2_23__17 ;
    input d_arr_merge2_23__16 ;
    input d_arr_merge2_23__15 ;
    input d_arr_merge2_23__14 ;
    input d_arr_merge2_23__13 ;
    input d_arr_merge2_23__12 ;
    input d_arr_merge2_23__11 ;
    input d_arr_merge2_23__10 ;
    input d_arr_merge2_23__9 ;
    input d_arr_merge2_23__8 ;
    input d_arr_merge2_23__7 ;
    input d_arr_merge2_23__6 ;
    input d_arr_merge2_23__5 ;
    input d_arr_merge2_23__4 ;
    input d_arr_merge2_23__3 ;
    input d_arr_merge2_23__2 ;
    input d_arr_merge2_23__1 ;
    input d_arr_merge2_23__0 ;
    input d_arr_merge2_24__31 ;
    input d_arr_merge2_24__30 ;
    input d_arr_merge2_24__29 ;
    input d_arr_merge2_24__28 ;
    input d_arr_merge2_24__27 ;
    input d_arr_merge2_24__26 ;
    input d_arr_merge2_24__25 ;
    input d_arr_merge2_24__24 ;
    input d_arr_merge2_24__23 ;
    input d_arr_merge2_24__22 ;
    input d_arr_merge2_24__21 ;
    input d_arr_merge2_24__20 ;
    input d_arr_merge2_24__19 ;
    input d_arr_merge2_24__18 ;
    input d_arr_merge2_24__17 ;
    input d_arr_merge2_24__16 ;
    input d_arr_merge2_24__15 ;
    input d_arr_merge2_24__14 ;
    input d_arr_merge2_24__13 ;
    input d_arr_merge2_24__12 ;
    input d_arr_merge2_24__11 ;
    input d_arr_merge2_24__10 ;
    input d_arr_merge2_24__9 ;
    input d_arr_merge2_24__8 ;
    input d_arr_merge2_24__7 ;
    input d_arr_merge2_24__6 ;
    input d_arr_merge2_24__5 ;
    input d_arr_merge2_24__4 ;
    input d_arr_merge2_24__3 ;
    input d_arr_merge2_24__2 ;
    input d_arr_merge2_24__1 ;
    input d_arr_merge2_24__0 ;
    input d_arr_relu_0__31 ;
    input d_arr_relu_0__30 ;
    input d_arr_relu_0__29 ;
    input d_arr_relu_0__28 ;
    input d_arr_relu_0__27 ;
    input d_arr_relu_0__26 ;
    input d_arr_relu_0__25 ;
    input d_arr_relu_0__24 ;
    input d_arr_relu_0__23 ;
    input d_arr_relu_0__22 ;
    input d_arr_relu_0__21 ;
    input d_arr_relu_0__20 ;
    input d_arr_relu_0__19 ;
    input d_arr_relu_0__18 ;
    input d_arr_relu_0__17 ;
    input d_arr_relu_0__16 ;
    input d_arr_relu_0__15 ;
    input d_arr_relu_0__14 ;
    input d_arr_relu_0__13 ;
    input d_arr_relu_0__12 ;
    input d_arr_relu_0__11 ;
    input d_arr_relu_0__10 ;
    input d_arr_relu_0__9 ;
    input d_arr_relu_0__8 ;
    input d_arr_relu_0__7 ;
    input d_arr_relu_0__6 ;
    input d_arr_relu_0__5 ;
    input d_arr_relu_0__4 ;
    input d_arr_relu_0__3 ;
    input d_arr_relu_0__2 ;
    input d_arr_relu_0__1 ;
    input d_arr_relu_0__0 ;
    input d_arr_relu_1__31 ;
    input d_arr_relu_1__30 ;
    input d_arr_relu_1__29 ;
    input d_arr_relu_1__28 ;
    input d_arr_relu_1__27 ;
    input d_arr_relu_1__26 ;
    input d_arr_relu_1__25 ;
    input d_arr_relu_1__24 ;
    input d_arr_relu_1__23 ;
    input d_arr_relu_1__22 ;
    input d_arr_relu_1__21 ;
    input d_arr_relu_1__20 ;
    input d_arr_relu_1__19 ;
    input d_arr_relu_1__18 ;
    input d_arr_relu_1__17 ;
    input d_arr_relu_1__16 ;
    input d_arr_relu_1__15 ;
    input d_arr_relu_1__14 ;
    input d_arr_relu_1__13 ;
    input d_arr_relu_1__12 ;
    input d_arr_relu_1__11 ;
    input d_arr_relu_1__10 ;
    input d_arr_relu_1__9 ;
    input d_arr_relu_1__8 ;
    input d_arr_relu_1__7 ;
    input d_arr_relu_1__6 ;
    input d_arr_relu_1__5 ;
    input d_arr_relu_1__4 ;
    input d_arr_relu_1__3 ;
    input d_arr_relu_1__2 ;
    input d_arr_relu_1__1 ;
    input d_arr_relu_1__0 ;
    input d_arr_relu_2__31 ;
    input d_arr_relu_2__30 ;
    input d_arr_relu_2__29 ;
    input d_arr_relu_2__28 ;
    input d_arr_relu_2__27 ;
    input d_arr_relu_2__26 ;
    input d_arr_relu_2__25 ;
    input d_arr_relu_2__24 ;
    input d_arr_relu_2__23 ;
    input d_arr_relu_2__22 ;
    input d_arr_relu_2__21 ;
    input d_arr_relu_2__20 ;
    input d_arr_relu_2__19 ;
    input d_arr_relu_2__18 ;
    input d_arr_relu_2__17 ;
    input d_arr_relu_2__16 ;
    input d_arr_relu_2__15 ;
    input d_arr_relu_2__14 ;
    input d_arr_relu_2__13 ;
    input d_arr_relu_2__12 ;
    input d_arr_relu_2__11 ;
    input d_arr_relu_2__10 ;
    input d_arr_relu_2__9 ;
    input d_arr_relu_2__8 ;
    input d_arr_relu_2__7 ;
    input d_arr_relu_2__6 ;
    input d_arr_relu_2__5 ;
    input d_arr_relu_2__4 ;
    input d_arr_relu_2__3 ;
    input d_arr_relu_2__2 ;
    input d_arr_relu_2__1 ;
    input d_arr_relu_2__0 ;
    input d_arr_relu_3__31 ;
    input d_arr_relu_3__30 ;
    input d_arr_relu_3__29 ;
    input d_arr_relu_3__28 ;
    input d_arr_relu_3__27 ;
    input d_arr_relu_3__26 ;
    input d_arr_relu_3__25 ;
    input d_arr_relu_3__24 ;
    input d_arr_relu_3__23 ;
    input d_arr_relu_3__22 ;
    input d_arr_relu_3__21 ;
    input d_arr_relu_3__20 ;
    input d_arr_relu_3__19 ;
    input d_arr_relu_3__18 ;
    input d_arr_relu_3__17 ;
    input d_arr_relu_3__16 ;
    input d_arr_relu_3__15 ;
    input d_arr_relu_3__14 ;
    input d_arr_relu_3__13 ;
    input d_arr_relu_3__12 ;
    input d_arr_relu_3__11 ;
    input d_arr_relu_3__10 ;
    input d_arr_relu_3__9 ;
    input d_arr_relu_3__8 ;
    input d_arr_relu_3__7 ;
    input d_arr_relu_3__6 ;
    input d_arr_relu_3__5 ;
    input d_arr_relu_3__4 ;
    input d_arr_relu_3__3 ;
    input d_arr_relu_3__2 ;
    input d_arr_relu_3__1 ;
    input d_arr_relu_3__0 ;
    input d_arr_relu_4__31 ;
    input d_arr_relu_4__30 ;
    input d_arr_relu_4__29 ;
    input d_arr_relu_4__28 ;
    input d_arr_relu_4__27 ;
    input d_arr_relu_4__26 ;
    input d_arr_relu_4__25 ;
    input d_arr_relu_4__24 ;
    input d_arr_relu_4__23 ;
    input d_arr_relu_4__22 ;
    input d_arr_relu_4__21 ;
    input d_arr_relu_4__20 ;
    input d_arr_relu_4__19 ;
    input d_arr_relu_4__18 ;
    input d_arr_relu_4__17 ;
    input d_arr_relu_4__16 ;
    input d_arr_relu_4__15 ;
    input d_arr_relu_4__14 ;
    input d_arr_relu_4__13 ;
    input d_arr_relu_4__12 ;
    input d_arr_relu_4__11 ;
    input d_arr_relu_4__10 ;
    input d_arr_relu_4__9 ;
    input d_arr_relu_4__8 ;
    input d_arr_relu_4__7 ;
    input d_arr_relu_4__6 ;
    input d_arr_relu_4__5 ;
    input d_arr_relu_4__4 ;
    input d_arr_relu_4__3 ;
    input d_arr_relu_4__2 ;
    input d_arr_relu_4__1 ;
    input d_arr_relu_4__0 ;
    input d_arr_relu_5__31 ;
    input d_arr_relu_5__30 ;
    input d_arr_relu_5__29 ;
    input d_arr_relu_5__28 ;
    input d_arr_relu_5__27 ;
    input d_arr_relu_5__26 ;
    input d_arr_relu_5__25 ;
    input d_arr_relu_5__24 ;
    input d_arr_relu_5__23 ;
    input d_arr_relu_5__22 ;
    input d_arr_relu_5__21 ;
    input d_arr_relu_5__20 ;
    input d_arr_relu_5__19 ;
    input d_arr_relu_5__18 ;
    input d_arr_relu_5__17 ;
    input d_arr_relu_5__16 ;
    input d_arr_relu_5__15 ;
    input d_arr_relu_5__14 ;
    input d_arr_relu_5__13 ;
    input d_arr_relu_5__12 ;
    input d_arr_relu_5__11 ;
    input d_arr_relu_5__10 ;
    input d_arr_relu_5__9 ;
    input d_arr_relu_5__8 ;
    input d_arr_relu_5__7 ;
    input d_arr_relu_5__6 ;
    input d_arr_relu_5__5 ;
    input d_arr_relu_5__4 ;
    input d_arr_relu_5__3 ;
    input d_arr_relu_5__2 ;
    input d_arr_relu_5__1 ;
    input d_arr_relu_5__0 ;
    input d_arr_relu_6__31 ;
    input d_arr_relu_6__30 ;
    input d_arr_relu_6__29 ;
    input d_arr_relu_6__28 ;
    input d_arr_relu_6__27 ;
    input d_arr_relu_6__26 ;
    input d_arr_relu_6__25 ;
    input d_arr_relu_6__24 ;
    input d_arr_relu_6__23 ;
    input d_arr_relu_6__22 ;
    input d_arr_relu_6__21 ;
    input d_arr_relu_6__20 ;
    input d_arr_relu_6__19 ;
    input d_arr_relu_6__18 ;
    input d_arr_relu_6__17 ;
    input d_arr_relu_6__16 ;
    input d_arr_relu_6__15 ;
    input d_arr_relu_6__14 ;
    input d_arr_relu_6__13 ;
    input d_arr_relu_6__12 ;
    input d_arr_relu_6__11 ;
    input d_arr_relu_6__10 ;
    input d_arr_relu_6__9 ;
    input d_arr_relu_6__8 ;
    input d_arr_relu_6__7 ;
    input d_arr_relu_6__6 ;
    input d_arr_relu_6__5 ;
    input d_arr_relu_6__4 ;
    input d_arr_relu_6__3 ;
    input d_arr_relu_6__2 ;
    input d_arr_relu_6__1 ;
    input d_arr_relu_6__0 ;
    input d_arr_relu_7__31 ;
    input d_arr_relu_7__30 ;
    input d_arr_relu_7__29 ;
    input d_arr_relu_7__28 ;
    input d_arr_relu_7__27 ;
    input d_arr_relu_7__26 ;
    input d_arr_relu_7__25 ;
    input d_arr_relu_7__24 ;
    input d_arr_relu_7__23 ;
    input d_arr_relu_7__22 ;
    input d_arr_relu_7__21 ;
    input d_arr_relu_7__20 ;
    input d_arr_relu_7__19 ;
    input d_arr_relu_7__18 ;
    input d_arr_relu_7__17 ;
    input d_arr_relu_7__16 ;
    input d_arr_relu_7__15 ;
    input d_arr_relu_7__14 ;
    input d_arr_relu_7__13 ;
    input d_arr_relu_7__12 ;
    input d_arr_relu_7__11 ;
    input d_arr_relu_7__10 ;
    input d_arr_relu_7__9 ;
    input d_arr_relu_7__8 ;
    input d_arr_relu_7__7 ;
    input d_arr_relu_7__6 ;
    input d_arr_relu_7__5 ;
    input d_arr_relu_7__4 ;
    input d_arr_relu_7__3 ;
    input d_arr_relu_7__2 ;
    input d_arr_relu_7__1 ;
    input d_arr_relu_7__0 ;
    input d_arr_relu_8__31 ;
    input d_arr_relu_8__30 ;
    input d_arr_relu_8__29 ;
    input d_arr_relu_8__28 ;
    input d_arr_relu_8__27 ;
    input d_arr_relu_8__26 ;
    input d_arr_relu_8__25 ;
    input d_arr_relu_8__24 ;
    input d_arr_relu_8__23 ;
    input d_arr_relu_8__22 ;
    input d_arr_relu_8__21 ;
    input d_arr_relu_8__20 ;
    input d_arr_relu_8__19 ;
    input d_arr_relu_8__18 ;
    input d_arr_relu_8__17 ;
    input d_arr_relu_8__16 ;
    input d_arr_relu_8__15 ;
    input d_arr_relu_8__14 ;
    input d_arr_relu_8__13 ;
    input d_arr_relu_8__12 ;
    input d_arr_relu_8__11 ;
    input d_arr_relu_8__10 ;
    input d_arr_relu_8__9 ;
    input d_arr_relu_8__8 ;
    input d_arr_relu_8__7 ;
    input d_arr_relu_8__6 ;
    input d_arr_relu_8__5 ;
    input d_arr_relu_8__4 ;
    input d_arr_relu_8__3 ;
    input d_arr_relu_8__2 ;
    input d_arr_relu_8__1 ;
    input d_arr_relu_8__0 ;
    input d_arr_relu_9__31 ;
    input d_arr_relu_9__30 ;
    input d_arr_relu_9__29 ;
    input d_arr_relu_9__28 ;
    input d_arr_relu_9__27 ;
    input d_arr_relu_9__26 ;
    input d_arr_relu_9__25 ;
    input d_arr_relu_9__24 ;
    input d_arr_relu_9__23 ;
    input d_arr_relu_9__22 ;
    input d_arr_relu_9__21 ;
    input d_arr_relu_9__20 ;
    input d_arr_relu_9__19 ;
    input d_arr_relu_9__18 ;
    input d_arr_relu_9__17 ;
    input d_arr_relu_9__16 ;
    input d_arr_relu_9__15 ;
    input d_arr_relu_9__14 ;
    input d_arr_relu_9__13 ;
    input d_arr_relu_9__12 ;
    input d_arr_relu_9__11 ;
    input d_arr_relu_9__10 ;
    input d_arr_relu_9__9 ;
    input d_arr_relu_9__8 ;
    input d_arr_relu_9__7 ;
    input d_arr_relu_9__6 ;
    input d_arr_relu_9__5 ;
    input d_arr_relu_9__4 ;
    input d_arr_relu_9__3 ;
    input d_arr_relu_9__2 ;
    input d_arr_relu_9__1 ;
    input d_arr_relu_9__0 ;
    input d_arr_relu_10__31 ;
    input d_arr_relu_10__30 ;
    input d_arr_relu_10__29 ;
    input d_arr_relu_10__28 ;
    input d_arr_relu_10__27 ;
    input d_arr_relu_10__26 ;
    input d_arr_relu_10__25 ;
    input d_arr_relu_10__24 ;
    input d_arr_relu_10__23 ;
    input d_arr_relu_10__22 ;
    input d_arr_relu_10__21 ;
    input d_arr_relu_10__20 ;
    input d_arr_relu_10__19 ;
    input d_arr_relu_10__18 ;
    input d_arr_relu_10__17 ;
    input d_arr_relu_10__16 ;
    input d_arr_relu_10__15 ;
    input d_arr_relu_10__14 ;
    input d_arr_relu_10__13 ;
    input d_arr_relu_10__12 ;
    input d_arr_relu_10__11 ;
    input d_arr_relu_10__10 ;
    input d_arr_relu_10__9 ;
    input d_arr_relu_10__8 ;
    input d_arr_relu_10__7 ;
    input d_arr_relu_10__6 ;
    input d_arr_relu_10__5 ;
    input d_arr_relu_10__4 ;
    input d_arr_relu_10__3 ;
    input d_arr_relu_10__2 ;
    input d_arr_relu_10__1 ;
    input d_arr_relu_10__0 ;
    input d_arr_relu_11__31 ;
    input d_arr_relu_11__30 ;
    input d_arr_relu_11__29 ;
    input d_arr_relu_11__28 ;
    input d_arr_relu_11__27 ;
    input d_arr_relu_11__26 ;
    input d_arr_relu_11__25 ;
    input d_arr_relu_11__24 ;
    input d_arr_relu_11__23 ;
    input d_arr_relu_11__22 ;
    input d_arr_relu_11__21 ;
    input d_arr_relu_11__20 ;
    input d_arr_relu_11__19 ;
    input d_arr_relu_11__18 ;
    input d_arr_relu_11__17 ;
    input d_arr_relu_11__16 ;
    input d_arr_relu_11__15 ;
    input d_arr_relu_11__14 ;
    input d_arr_relu_11__13 ;
    input d_arr_relu_11__12 ;
    input d_arr_relu_11__11 ;
    input d_arr_relu_11__10 ;
    input d_arr_relu_11__9 ;
    input d_arr_relu_11__8 ;
    input d_arr_relu_11__7 ;
    input d_arr_relu_11__6 ;
    input d_arr_relu_11__5 ;
    input d_arr_relu_11__4 ;
    input d_arr_relu_11__3 ;
    input d_arr_relu_11__2 ;
    input d_arr_relu_11__1 ;
    input d_arr_relu_11__0 ;
    input d_arr_relu_12__31 ;
    input d_arr_relu_12__30 ;
    input d_arr_relu_12__29 ;
    input d_arr_relu_12__28 ;
    input d_arr_relu_12__27 ;
    input d_arr_relu_12__26 ;
    input d_arr_relu_12__25 ;
    input d_arr_relu_12__24 ;
    input d_arr_relu_12__23 ;
    input d_arr_relu_12__22 ;
    input d_arr_relu_12__21 ;
    input d_arr_relu_12__20 ;
    input d_arr_relu_12__19 ;
    input d_arr_relu_12__18 ;
    input d_arr_relu_12__17 ;
    input d_arr_relu_12__16 ;
    input d_arr_relu_12__15 ;
    input d_arr_relu_12__14 ;
    input d_arr_relu_12__13 ;
    input d_arr_relu_12__12 ;
    input d_arr_relu_12__11 ;
    input d_arr_relu_12__10 ;
    input d_arr_relu_12__9 ;
    input d_arr_relu_12__8 ;
    input d_arr_relu_12__7 ;
    input d_arr_relu_12__6 ;
    input d_arr_relu_12__5 ;
    input d_arr_relu_12__4 ;
    input d_arr_relu_12__3 ;
    input d_arr_relu_12__2 ;
    input d_arr_relu_12__1 ;
    input d_arr_relu_12__0 ;
    input d_arr_relu_13__31 ;
    input d_arr_relu_13__30 ;
    input d_arr_relu_13__29 ;
    input d_arr_relu_13__28 ;
    input d_arr_relu_13__27 ;
    input d_arr_relu_13__26 ;
    input d_arr_relu_13__25 ;
    input d_arr_relu_13__24 ;
    input d_arr_relu_13__23 ;
    input d_arr_relu_13__22 ;
    input d_arr_relu_13__21 ;
    input d_arr_relu_13__20 ;
    input d_arr_relu_13__19 ;
    input d_arr_relu_13__18 ;
    input d_arr_relu_13__17 ;
    input d_arr_relu_13__16 ;
    input d_arr_relu_13__15 ;
    input d_arr_relu_13__14 ;
    input d_arr_relu_13__13 ;
    input d_arr_relu_13__12 ;
    input d_arr_relu_13__11 ;
    input d_arr_relu_13__10 ;
    input d_arr_relu_13__9 ;
    input d_arr_relu_13__8 ;
    input d_arr_relu_13__7 ;
    input d_arr_relu_13__6 ;
    input d_arr_relu_13__5 ;
    input d_arr_relu_13__4 ;
    input d_arr_relu_13__3 ;
    input d_arr_relu_13__2 ;
    input d_arr_relu_13__1 ;
    input d_arr_relu_13__0 ;
    input d_arr_relu_14__31 ;
    input d_arr_relu_14__30 ;
    input d_arr_relu_14__29 ;
    input d_arr_relu_14__28 ;
    input d_arr_relu_14__27 ;
    input d_arr_relu_14__26 ;
    input d_arr_relu_14__25 ;
    input d_arr_relu_14__24 ;
    input d_arr_relu_14__23 ;
    input d_arr_relu_14__22 ;
    input d_arr_relu_14__21 ;
    input d_arr_relu_14__20 ;
    input d_arr_relu_14__19 ;
    input d_arr_relu_14__18 ;
    input d_arr_relu_14__17 ;
    input d_arr_relu_14__16 ;
    input d_arr_relu_14__15 ;
    input d_arr_relu_14__14 ;
    input d_arr_relu_14__13 ;
    input d_arr_relu_14__12 ;
    input d_arr_relu_14__11 ;
    input d_arr_relu_14__10 ;
    input d_arr_relu_14__9 ;
    input d_arr_relu_14__8 ;
    input d_arr_relu_14__7 ;
    input d_arr_relu_14__6 ;
    input d_arr_relu_14__5 ;
    input d_arr_relu_14__4 ;
    input d_arr_relu_14__3 ;
    input d_arr_relu_14__2 ;
    input d_arr_relu_14__1 ;
    input d_arr_relu_14__0 ;
    input d_arr_relu_15__31 ;
    input d_arr_relu_15__30 ;
    input d_arr_relu_15__29 ;
    input d_arr_relu_15__28 ;
    input d_arr_relu_15__27 ;
    input d_arr_relu_15__26 ;
    input d_arr_relu_15__25 ;
    input d_arr_relu_15__24 ;
    input d_arr_relu_15__23 ;
    input d_arr_relu_15__22 ;
    input d_arr_relu_15__21 ;
    input d_arr_relu_15__20 ;
    input d_arr_relu_15__19 ;
    input d_arr_relu_15__18 ;
    input d_arr_relu_15__17 ;
    input d_arr_relu_15__16 ;
    input d_arr_relu_15__15 ;
    input d_arr_relu_15__14 ;
    input d_arr_relu_15__13 ;
    input d_arr_relu_15__12 ;
    input d_arr_relu_15__11 ;
    input d_arr_relu_15__10 ;
    input d_arr_relu_15__9 ;
    input d_arr_relu_15__8 ;
    input d_arr_relu_15__7 ;
    input d_arr_relu_15__6 ;
    input d_arr_relu_15__5 ;
    input d_arr_relu_15__4 ;
    input d_arr_relu_15__3 ;
    input d_arr_relu_15__2 ;
    input d_arr_relu_15__1 ;
    input d_arr_relu_15__0 ;
    input d_arr_relu_16__31 ;
    input d_arr_relu_16__30 ;
    input d_arr_relu_16__29 ;
    input d_arr_relu_16__28 ;
    input d_arr_relu_16__27 ;
    input d_arr_relu_16__26 ;
    input d_arr_relu_16__25 ;
    input d_arr_relu_16__24 ;
    input d_arr_relu_16__23 ;
    input d_arr_relu_16__22 ;
    input d_arr_relu_16__21 ;
    input d_arr_relu_16__20 ;
    input d_arr_relu_16__19 ;
    input d_arr_relu_16__18 ;
    input d_arr_relu_16__17 ;
    input d_arr_relu_16__16 ;
    input d_arr_relu_16__15 ;
    input d_arr_relu_16__14 ;
    input d_arr_relu_16__13 ;
    input d_arr_relu_16__12 ;
    input d_arr_relu_16__11 ;
    input d_arr_relu_16__10 ;
    input d_arr_relu_16__9 ;
    input d_arr_relu_16__8 ;
    input d_arr_relu_16__7 ;
    input d_arr_relu_16__6 ;
    input d_arr_relu_16__5 ;
    input d_arr_relu_16__4 ;
    input d_arr_relu_16__3 ;
    input d_arr_relu_16__2 ;
    input d_arr_relu_16__1 ;
    input d_arr_relu_16__0 ;
    input d_arr_relu_17__31 ;
    input d_arr_relu_17__30 ;
    input d_arr_relu_17__29 ;
    input d_arr_relu_17__28 ;
    input d_arr_relu_17__27 ;
    input d_arr_relu_17__26 ;
    input d_arr_relu_17__25 ;
    input d_arr_relu_17__24 ;
    input d_arr_relu_17__23 ;
    input d_arr_relu_17__22 ;
    input d_arr_relu_17__21 ;
    input d_arr_relu_17__20 ;
    input d_arr_relu_17__19 ;
    input d_arr_relu_17__18 ;
    input d_arr_relu_17__17 ;
    input d_arr_relu_17__16 ;
    input d_arr_relu_17__15 ;
    input d_arr_relu_17__14 ;
    input d_arr_relu_17__13 ;
    input d_arr_relu_17__12 ;
    input d_arr_relu_17__11 ;
    input d_arr_relu_17__10 ;
    input d_arr_relu_17__9 ;
    input d_arr_relu_17__8 ;
    input d_arr_relu_17__7 ;
    input d_arr_relu_17__6 ;
    input d_arr_relu_17__5 ;
    input d_arr_relu_17__4 ;
    input d_arr_relu_17__3 ;
    input d_arr_relu_17__2 ;
    input d_arr_relu_17__1 ;
    input d_arr_relu_17__0 ;
    input d_arr_relu_18__31 ;
    input d_arr_relu_18__30 ;
    input d_arr_relu_18__29 ;
    input d_arr_relu_18__28 ;
    input d_arr_relu_18__27 ;
    input d_arr_relu_18__26 ;
    input d_arr_relu_18__25 ;
    input d_arr_relu_18__24 ;
    input d_arr_relu_18__23 ;
    input d_arr_relu_18__22 ;
    input d_arr_relu_18__21 ;
    input d_arr_relu_18__20 ;
    input d_arr_relu_18__19 ;
    input d_arr_relu_18__18 ;
    input d_arr_relu_18__17 ;
    input d_arr_relu_18__16 ;
    input d_arr_relu_18__15 ;
    input d_arr_relu_18__14 ;
    input d_arr_relu_18__13 ;
    input d_arr_relu_18__12 ;
    input d_arr_relu_18__11 ;
    input d_arr_relu_18__10 ;
    input d_arr_relu_18__9 ;
    input d_arr_relu_18__8 ;
    input d_arr_relu_18__7 ;
    input d_arr_relu_18__6 ;
    input d_arr_relu_18__5 ;
    input d_arr_relu_18__4 ;
    input d_arr_relu_18__3 ;
    input d_arr_relu_18__2 ;
    input d_arr_relu_18__1 ;
    input d_arr_relu_18__0 ;
    input d_arr_relu_19__31 ;
    input d_arr_relu_19__30 ;
    input d_arr_relu_19__29 ;
    input d_arr_relu_19__28 ;
    input d_arr_relu_19__27 ;
    input d_arr_relu_19__26 ;
    input d_arr_relu_19__25 ;
    input d_arr_relu_19__24 ;
    input d_arr_relu_19__23 ;
    input d_arr_relu_19__22 ;
    input d_arr_relu_19__21 ;
    input d_arr_relu_19__20 ;
    input d_arr_relu_19__19 ;
    input d_arr_relu_19__18 ;
    input d_arr_relu_19__17 ;
    input d_arr_relu_19__16 ;
    input d_arr_relu_19__15 ;
    input d_arr_relu_19__14 ;
    input d_arr_relu_19__13 ;
    input d_arr_relu_19__12 ;
    input d_arr_relu_19__11 ;
    input d_arr_relu_19__10 ;
    input d_arr_relu_19__9 ;
    input d_arr_relu_19__8 ;
    input d_arr_relu_19__7 ;
    input d_arr_relu_19__6 ;
    input d_arr_relu_19__5 ;
    input d_arr_relu_19__4 ;
    input d_arr_relu_19__3 ;
    input d_arr_relu_19__2 ;
    input d_arr_relu_19__1 ;
    input d_arr_relu_19__0 ;
    input d_arr_relu_20__31 ;
    input d_arr_relu_20__30 ;
    input d_arr_relu_20__29 ;
    input d_arr_relu_20__28 ;
    input d_arr_relu_20__27 ;
    input d_arr_relu_20__26 ;
    input d_arr_relu_20__25 ;
    input d_arr_relu_20__24 ;
    input d_arr_relu_20__23 ;
    input d_arr_relu_20__22 ;
    input d_arr_relu_20__21 ;
    input d_arr_relu_20__20 ;
    input d_arr_relu_20__19 ;
    input d_arr_relu_20__18 ;
    input d_arr_relu_20__17 ;
    input d_arr_relu_20__16 ;
    input d_arr_relu_20__15 ;
    input d_arr_relu_20__14 ;
    input d_arr_relu_20__13 ;
    input d_arr_relu_20__12 ;
    input d_arr_relu_20__11 ;
    input d_arr_relu_20__10 ;
    input d_arr_relu_20__9 ;
    input d_arr_relu_20__8 ;
    input d_arr_relu_20__7 ;
    input d_arr_relu_20__6 ;
    input d_arr_relu_20__5 ;
    input d_arr_relu_20__4 ;
    input d_arr_relu_20__3 ;
    input d_arr_relu_20__2 ;
    input d_arr_relu_20__1 ;
    input d_arr_relu_20__0 ;
    input d_arr_relu_21__31 ;
    input d_arr_relu_21__30 ;
    input d_arr_relu_21__29 ;
    input d_arr_relu_21__28 ;
    input d_arr_relu_21__27 ;
    input d_arr_relu_21__26 ;
    input d_arr_relu_21__25 ;
    input d_arr_relu_21__24 ;
    input d_arr_relu_21__23 ;
    input d_arr_relu_21__22 ;
    input d_arr_relu_21__21 ;
    input d_arr_relu_21__20 ;
    input d_arr_relu_21__19 ;
    input d_arr_relu_21__18 ;
    input d_arr_relu_21__17 ;
    input d_arr_relu_21__16 ;
    input d_arr_relu_21__15 ;
    input d_arr_relu_21__14 ;
    input d_arr_relu_21__13 ;
    input d_arr_relu_21__12 ;
    input d_arr_relu_21__11 ;
    input d_arr_relu_21__10 ;
    input d_arr_relu_21__9 ;
    input d_arr_relu_21__8 ;
    input d_arr_relu_21__7 ;
    input d_arr_relu_21__6 ;
    input d_arr_relu_21__5 ;
    input d_arr_relu_21__4 ;
    input d_arr_relu_21__3 ;
    input d_arr_relu_21__2 ;
    input d_arr_relu_21__1 ;
    input d_arr_relu_21__0 ;
    input d_arr_relu_22__31 ;
    input d_arr_relu_22__30 ;
    input d_arr_relu_22__29 ;
    input d_arr_relu_22__28 ;
    input d_arr_relu_22__27 ;
    input d_arr_relu_22__26 ;
    input d_arr_relu_22__25 ;
    input d_arr_relu_22__24 ;
    input d_arr_relu_22__23 ;
    input d_arr_relu_22__22 ;
    input d_arr_relu_22__21 ;
    input d_arr_relu_22__20 ;
    input d_arr_relu_22__19 ;
    input d_arr_relu_22__18 ;
    input d_arr_relu_22__17 ;
    input d_arr_relu_22__16 ;
    input d_arr_relu_22__15 ;
    input d_arr_relu_22__14 ;
    input d_arr_relu_22__13 ;
    input d_arr_relu_22__12 ;
    input d_arr_relu_22__11 ;
    input d_arr_relu_22__10 ;
    input d_arr_relu_22__9 ;
    input d_arr_relu_22__8 ;
    input d_arr_relu_22__7 ;
    input d_arr_relu_22__6 ;
    input d_arr_relu_22__5 ;
    input d_arr_relu_22__4 ;
    input d_arr_relu_22__3 ;
    input d_arr_relu_22__2 ;
    input d_arr_relu_22__1 ;
    input d_arr_relu_22__0 ;
    input d_arr_relu_23__31 ;
    input d_arr_relu_23__30 ;
    input d_arr_relu_23__29 ;
    input d_arr_relu_23__28 ;
    input d_arr_relu_23__27 ;
    input d_arr_relu_23__26 ;
    input d_arr_relu_23__25 ;
    input d_arr_relu_23__24 ;
    input d_arr_relu_23__23 ;
    input d_arr_relu_23__22 ;
    input d_arr_relu_23__21 ;
    input d_arr_relu_23__20 ;
    input d_arr_relu_23__19 ;
    input d_arr_relu_23__18 ;
    input d_arr_relu_23__17 ;
    input d_arr_relu_23__16 ;
    input d_arr_relu_23__15 ;
    input d_arr_relu_23__14 ;
    input d_arr_relu_23__13 ;
    input d_arr_relu_23__12 ;
    input d_arr_relu_23__11 ;
    input d_arr_relu_23__10 ;
    input d_arr_relu_23__9 ;
    input d_arr_relu_23__8 ;
    input d_arr_relu_23__7 ;
    input d_arr_relu_23__6 ;
    input d_arr_relu_23__5 ;
    input d_arr_relu_23__4 ;
    input d_arr_relu_23__3 ;
    input d_arr_relu_23__2 ;
    input d_arr_relu_23__1 ;
    input d_arr_relu_23__0 ;
    input d_arr_relu_24__31 ;
    input d_arr_relu_24__30 ;
    input d_arr_relu_24__29 ;
    input d_arr_relu_24__28 ;
    input d_arr_relu_24__27 ;
    input d_arr_relu_24__26 ;
    input d_arr_relu_24__25 ;
    input d_arr_relu_24__24 ;
    input d_arr_relu_24__23 ;
    input d_arr_relu_24__22 ;
    input d_arr_relu_24__21 ;
    input d_arr_relu_24__20 ;
    input d_arr_relu_24__19 ;
    input d_arr_relu_24__18 ;
    input d_arr_relu_24__17 ;
    input d_arr_relu_24__16 ;
    input d_arr_relu_24__15 ;
    input d_arr_relu_24__14 ;
    input d_arr_relu_24__13 ;
    input d_arr_relu_24__12 ;
    input d_arr_relu_24__11 ;
    input d_arr_relu_24__10 ;
    input d_arr_relu_24__9 ;
    input d_arr_relu_24__8 ;
    input d_arr_relu_24__7 ;
    input d_arr_relu_24__6 ;
    input d_arr_relu_24__5 ;
    input d_arr_relu_24__4 ;
    input d_arr_relu_24__3 ;
    input d_arr_relu_24__2 ;
    input d_arr_relu_24__1 ;
    input d_arr_relu_24__0 ;
    input sel_mux ;
    input sel_mul ;
    input sel_add ;
    input sel_merge1 ;
    input sel_merge2 ;
    input sel_relu ;
    output d_arr_0__31 ;
    output d_arr_0__30 ;
    output d_arr_0__29 ;
    output d_arr_0__28 ;
    output d_arr_0__27 ;
    output d_arr_0__26 ;
    output d_arr_0__25 ;
    output d_arr_0__24 ;
    output d_arr_0__23 ;
    output d_arr_0__22 ;
    output d_arr_0__21 ;
    output d_arr_0__20 ;
    output d_arr_0__19 ;
    output d_arr_0__18 ;
    output d_arr_0__17 ;
    output d_arr_0__16 ;
    output d_arr_0__15 ;
    output d_arr_0__14 ;
    output d_arr_0__13 ;
    output d_arr_0__12 ;
    output d_arr_0__11 ;
    output d_arr_0__10 ;
    output d_arr_0__9 ;
    output d_arr_0__8 ;
    output d_arr_0__7 ;
    output d_arr_0__6 ;
    output d_arr_0__5 ;
    output d_arr_0__4 ;
    output d_arr_0__3 ;
    output d_arr_0__2 ;
    output d_arr_0__1 ;
    output d_arr_0__0 ;
    output d_arr_1__31 ;
    output d_arr_1__30 ;
    output d_arr_1__29 ;
    output d_arr_1__28 ;
    output d_arr_1__27 ;
    output d_arr_1__26 ;
    output d_arr_1__25 ;
    output d_arr_1__24 ;
    output d_arr_1__23 ;
    output d_arr_1__22 ;
    output d_arr_1__21 ;
    output d_arr_1__20 ;
    output d_arr_1__19 ;
    output d_arr_1__18 ;
    output d_arr_1__17 ;
    output d_arr_1__16 ;
    output d_arr_1__15 ;
    output d_arr_1__14 ;
    output d_arr_1__13 ;
    output d_arr_1__12 ;
    output d_arr_1__11 ;
    output d_arr_1__10 ;
    output d_arr_1__9 ;
    output d_arr_1__8 ;
    output d_arr_1__7 ;
    output d_arr_1__6 ;
    output d_arr_1__5 ;
    output d_arr_1__4 ;
    output d_arr_1__3 ;
    output d_arr_1__2 ;
    output d_arr_1__1 ;
    output d_arr_1__0 ;
    output d_arr_2__31 ;
    output d_arr_2__30 ;
    output d_arr_2__29 ;
    output d_arr_2__28 ;
    output d_arr_2__27 ;
    output d_arr_2__26 ;
    output d_arr_2__25 ;
    output d_arr_2__24 ;
    output d_arr_2__23 ;
    output d_arr_2__22 ;
    output d_arr_2__21 ;
    output d_arr_2__20 ;
    output d_arr_2__19 ;
    output d_arr_2__18 ;
    output d_arr_2__17 ;
    output d_arr_2__16 ;
    output d_arr_2__15 ;
    output d_arr_2__14 ;
    output d_arr_2__13 ;
    output d_arr_2__12 ;
    output d_arr_2__11 ;
    output d_arr_2__10 ;
    output d_arr_2__9 ;
    output d_arr_2__8 ;
    output d_arr_2__7 ;
    output d_arr_2__6 ;
    output d_arr_2__5 ;
    output d_arr_2__4 ;
    output d_arr_2__3 ;
    output d_arr_2__2 ;
    output d_arr_2__1 ;
    output d_arr_2__0 ;
    output d_arr_3__31 ;
    output d_arr_3__30 ;
    output d_arr_3__29 ;
    output d_arr_3__28 ;
    output d_arr_3__27 ;
    output d_arr_3__26 ;
    output d_arr_3__25 ;
    output d_arr_3__24 ;
    output d_arr_3__23 ;
    output d_arr_3__22 ;
    output d_arr_3__21 ;
    output d_arr_3__20 ;
    output d_arr_3__19 ;
    output d_arr_3__18 ;
    output d_arr_3__17 ;
    output d_arr_3__16 ;
    output d_arr_3__15 ;
    output d_arr_3__14 ;
    output d_arr_3__13 ;
    output d_arr_3__12 ;
    output d_arr_3__11 ;
    output d_arr_3__10 ;
    output d_arr_3__9 ;
    output d_arr_3__8 ;
    output d_arr_3__7 ;
    output d_arr_3__6 ;
    output d_arr_3__5 ;
    output d_arr_3__4 ;
    output d_arr_3__3 ;
    output d_arr_3__2 ;
    output d_arr_3__1 ;
    output d_arr_3__0 ;
    output d_arr_4__31 ;
    output d_arr_4__30 ;
    output d_arr_4__29 ;
    output d_arr_4__28 ;
    output d_arr_4__27 ;
    output d_arr_4__26 ;
    output d_arr_4__25 ;
    output d_arr_4__24 ;
    output d_arr_4__23 ;
    output d_arr_4__22 ;
    output d_arr_4__21 ;
    output d_arr_4__20 ;
    output d_arr_4__19 ;
    output d_arr_4__18 ;
    output d_arr_4__17 ;
    output d_arr_4__16 ;
    output d_arr_4__15 ;
    output d_arr_4__14 ;
    output d_arr_4__13 ;
    output d_arr_4__12 ;
    output d_arr_4__11 ;
    output d_arr_4__10 ;
    output d_arr_4__9 ;
    output d_arr_4__8 ;
    output d_arr_4__7 ;
    output d_arr_4__6 ;
    output d_arr_4__5 ;
    output d_arr_4__4 ;
    output d_arr_4__3 ;
    output d_arr_4__2 ;
    output d_arr_4__1 ;
    output d_arr_4__0 ;
    output d_arr_5__31 ;
    output d_arr_5__30 ;
    output d_arr_5__29 ;
    output d_arr_5__28 ;
    output d_arr_5__27 ;
    output d_arr_5__26 ;
    output d_arr_5__25 ;
    output d_arr_5__24 ;
    output d_arr_5__23 ;
    output d_arr_5__22 ;
    output d_arr_5__21 ;
    output d_arr_5__20 ;
    output d_arr_5__19 ;
    output d_arr_5__18 ;
    output d_arr_5__17 ;
    output d_arr_5__16 ;
    output d_arr_5__15 ;
    output d_arr_5__14 ;
    output d_arr_5__13 ;
    output d_arr_5__12 ;
    output d_arr_5__11 ;
    output d_arr_5__10 ;
    output d_arr_5__9 ;
    output d_arr_5__8 ;
    output d_arr_5__7 ;
    output d_arr_5__6 ;
    output d_arr_5__5 ;
    output d_arr_5__4 ;
    output d_arr_5__3 ;
    output d_arr_5__2 ;
    output d_arr_5__1 ;
    output d_arr_5__0 ;
    output d_arr_6__31 ;
    output d_arr_6__30 ;
    output d_arr_6__29 ;
    output d_arr_6__28 ;
    output d_arr_6__27 ;
    output d_arr_6__26 ;
    output d_arr_6__25 ;
    output d_arr_6__24 ;
    output d_arr_6__23 ;
    output d_arr_6__22 ;
    output d_arr_6__21 ;
    output d_arr_6__20 ;
    output d_arr_6__19 ;
    output d_arr_6__18 ;
    output d_arr_6__17 ;
    output d_arr_6__16 ;
    output d_arr_6__15 ;
    output d_arr_6__14 ;
    output d_arr_6__13 ;
    output d_arr_6__12 ;
    output d_arr_6__11 ;
    output d_arr_6__10 ;
    output d_arr_6__9 ;
    output d_arr_6__8 ;
    output d_arr_6__7 ;
    output d_arr_6__6 ;
    output d_arr_6__5 ;
    output d_arr_6__4 ;
    output d_arr_6__3 ;
    output d_arr_6__2 ;
    output d_arr_6__1 ;
    output d_arr_6__0 ;
    output d_arr_7__31 ;
    output d_arr_7__30 ;
    output d_arr_7__29 ;
    output d_arr_7__28 ;
    output d_arr_7__27 ;
    output d_arr_7__26 ;
    output d_arr_7__25 ;
    output d_arr_7__24 ;
    output d_arr_7__23 ;
    output d_arr_7__22 ;
    output d_arr_7__21 ;
    output d_arr_7__20 ;
    output d_arr_7__19 ;
    output d_arr_7__18 ;
    output d_arr_7__17 ;
    output d_arr_7__16 ;
    output d_arr_7__15 ;
    output d_arr_7__14 ;
    output d_arr_7__13 ;
    output d_arr_7__12 ;
    output d_arr_7__11 ;
    output d_arr_7__10 ;
    output d_arr_7__9 ;
    output d_arr_7__8 ;
    output d_arr_7__7 ;
    output d_arr_7__6 ;
    output d_arr_7__5 ;
    output d_arr_7__4 ;
    output d_arr_7__3 ;
    output d_arr_7__2 ;
    output d_arr_7__1 ;
    output d_arr_7__0 ;
    output d_arr_8__31 ;
    output d_arr_8__30 ;
    output d_arr_8__29 ;
    output d_arr_8__28 ;
    output d_arr_8__27 ;
    output d_arr_8__26 ;
    output d_arr_8__25 ;
    output d_arr_8__24 ;
    output d_arr_8__23 ;
    output d_arr_8__22 ;
    output d_arr_8__21 ;
    output d_arr_8__20 ;
    output d_arr_8__19 ;
    output d_arr_8__18 ;
    output d_arr_8__17 ;
    output d_arr_8__16 ;
    output d_arr_8__15 ;
    output d_arr_8__14 ;
    output d_arr_8__13 ;
    output d_arr_8__12 ;
    output d_arr_8__11 ;
    output d_arr_8__10 ;
    output d_arr_8__9 ;
    output d_arr_8__8 ;
    output d_arr_8__7 ;
    output d_arr_8__6 ;
    output d_arr_8__5 ;
    output d_arr_8__4 ;
    output d_arr_8__3 ;
    output d_arr_8__2 ;
    output d_arr_8__1 ;
    output d_arr_8__0 ;
    output d_arr_9__31 ;
    output d_arr_9__30 ;
    output d_arr_9__29 ;
    output d_arr_9__28 ;
    output d_arr_9__27 ;
    output d_arr_9__26 ;
    output d_arr_9__25 ;
    output d_arr_9__24 ;
    output d_arr_9__23 ;
    output d_arr_9__22 ;
    output d_arr_9__21 ;
    output d_arr_9__20 ;
    output d_arr_9__19 ;
    output d_arr_9__18 ;
    output d_arr_9__17 ;
    output d_arr_9__16 ;
    output d_arr_9__15 ;
    output d_arr_9__14 ;
    output d_arr_9__13 ;
    output d_arr_9__12 ;
    output d_arr_9__11 ;
    output d_arr_9__10 ;
    output d_arr_9__9 ;
    output d_arr_9__8 ;
    output d_arr_9__7 ;
    output d_arr_9__6 ;
    output d_arr_9__5 ;
    output d_arr_9__4 ;
    output d_arr_9__3 ;
    output d_arr_9__2 ;
    output d_arr_9__1 ;
    output d_arr_9__0 ;
    output d_arr_10__31 ;
    output d_arr_10__30 ;
    output d_arr_10__29 ;
    output d_arr_10__28 ;
    output d_arr_10__27 ;
    output d_arr_10__26 ;
    output d_arr_10__25 ;
    output d_arr_10__24 ;
    output d_arr_10__23 ;
    output d_arr_10__22 ;
    output d_arr_10__21 ;
    output d_arr_10__20 ;
    output d_arr_10__19 ;
    output d_arr_10__18 ;
    output d_arr_10__17 ;
    output d_arr_10__16 ;
    output d_arr_10__15 ;
    output d_arr_10__14 ;
    output d_arr_10__13 ;
    output d_arr_10__12 ;
    output d_arr_10__11 ;
    output d_arr_10__10 ;
    output d_arr_10__9 ;
    output d_arr_10__8 ;
    output d_arr_10__7 ;
    output d_arr_10__6 ;
    output d_arr_10__5 ;
    output d_arr_10__4 ;
    output d_arr_10__3 ;
    output d_arr_10__2 ;
    output d_arr_10__1 ;
    output d_arr_10__0 ;
    output d_arr_11__31 ;
    output d_arr_11__30 ;
    output d_arr_11__29 ;
    output d_arr_11__28 ;
    output d_arr_11__27 ;
    output d_arr_11__26 ;
    output d_arr_11__25 ;
    output d_arr_11__24 ;
    output d_arr_11__23 ;
    output d_arr_11__22 ;
    output d_arr_11__21 ;
    output d_arr_11__20 ;
    output d_arr_11__19 ;
    output d_arr_11__18 ;
    output d_arr_11__17 ;
    output d_arr_11__16 ;
    output d_arr_11__15 ;
    output d_arr_11__14 ;
    output d_arr_11__13 ;
    output d_arr_11__12 ;
    output d_arr_11__11 ;
    output d_arr_11__10 ;
    output d_arr_11__9 ;
    output d_arr_11__8 ;
    output d_arr_11__7 ;
    output d_arr_11__6 ;
    output d_arr_11__5 ;
    output d_arr_11__4 ;
    output d_arr_11__3 ;
    output d_arr_11__2 ;
    output d_arr_11__1 ;
    output d_arr_11__0 ;
    output d_arr_12__31 ;
    output d_arr_12__30 ;
    output d_arr_12__29 ;
    output d_arr_12__28 ;
    output d_arr_12__27 ;
    output d_arr_12__26 ;
    output d_arr_12__25 ;
    output d_arr_12__24 ;
    output d_arr_12__23 ;
    output d_arr_12__22 ;
    output d_arr_12__21 ;
    output d_arr_12__20 ;
    output d_arr_12__19 ;
    output d_arr_12__18 ;
    output d_arr_12__17 ;
    output d_arr_12__16 ;
    output d_arr_12__15 ;
    output d_arr_12__14 ;
    output d_arr_12__13 ;
    output d_arr_12__12 ;
    output d_arr_12__11 ;
    output d_arr_12__10 ;
    output d_arr_12__9 ;
    output d_arr_12__8 ;
    output d_arr_12__7 ;
    output d_arr_12__6 ;
    output d_arr_12__5 ;
    output d_arr_12__4 ;
    output d_arr_12__3 ;
    output d_arr_12__2 ;
    output d_arr_12__1 ;
    output d_arr_12__0 ;
    output d_arr_13__31 ;
    output d_arr_13__30 ;
    output d_arr_13__29 ;
    output d_arr_13__28 ;
    output d_arr_13__27 ;
    output d_arr_13__26 ;
    output d_arr_13__25 ;
    output d_arr_13__24 ;
    output d_arr_13__23 ;
    output d_arr_13__22 ;
    output d_arr_13__21 ;
    output d_arr_13__20 ;
    output d_arr_13__19 ;
    output d_arr_13__18 ;
    output d_arr_13__17 ;
    output d_arr_13__16 ;
    output d_arr_13__15 ;
    output d_arr_13__14 ;
    output d_arr_13__13 ;
    output d_arr_13__12 ;
    output d_arr_13__11 ;
    output d_arr_13__10 ;
    output d_arr_13__9 ;
    output d_arr_13__8 ;
    output d_arr_13__7 ;
    output d_arr_13__6 ;
    output d_arr_13__5 ;
    output d_arr_13__4 ;
    output d_arr_13__3 ;
    output d_arr_13__2 ;
    output d_arr_13__1 ;
    output d_arr_13__0 ;
    output d_arr_14__31 ;
    output d_arr_14__30 ;
    output d_arr_14__29 ;
    output d_arr_14__28 ;
    output d_arr_14__27 ;
    output d_arr_14__26 ;
    output d_arr_14__25 ;
    output d_arr_14__24 ;
    output d_arr_14__23 ;
    output d_arr_14__22 ;
    output d_arr_14__21 ;
    output d_arr_14__20 ;
    output d_arr_14__19 ;
    output d_arr_14__18 ;
    output d_arr_14__17 ;
    output d_arr_14__16 ;
    output d_arr_14__15 ;
    output d_arr_14__14 ;
    output d_arr_14__13 ;
    output d_arr_14__12 ;
    output d_arr_14__11 ;
    output d_arr_14__10 ;
    output d_arr_14__9 ;
    output d_arr_14__8 ;
    output d_arr_14__7 ;
    output d_arr_14__6 ;
    output d_arr_14__5 ;
    output d_arr_14__4 ;
    output d_arr_14__3 ;
    output d_arr_14__2 ;
    output d_arr_14__1 ;
    output d_arr_14__0 ;
    output d_arr_15__31 ;
    output d_arr_15__30 ;
    output d_arr_15__29 ;
    output d_arr_15__28 ;
    output d_arr_15__27 ;
    output d_arr_15__26 ;
    output d_arr_15__25 ;
    output d_arr_15__24 ;
    output d_arr_15__23 ;
    output d_arr_15__22 ;
    output d_arr_15__21 ;
    output d_arr_15__20 ;
    output d_arr_15__19 ;
    output d_arr_15__18 ;
    output d_arr_15__17 ;
    output d_arr_15__16 ;
    output d_arr_15__15 ;
    output d_arr_15__14 ;
    output d_arr_15__13 ;
    output d_arr_15__12 ;
    output d_arr_15__11 ;
    output d_arr_15__10 ;
    output d_arr_15__9 ;
    output d_arr_15__8 ;
    output d_arr_15__7 ;
    output d_arr_15__6 ;
    output d_arr_15__5 ;
    output d_arr_15__4 ;
    output d_arr_15__3 ;
    output d_arr_15__2 ;
    output d_arr_15__1 ;
    output d_arr_15__0 ;
    output d_arr_16__31 ;
    output d_arr_16__30 ;
    output d_arr_16__29 ;
    output d_arr_16__28 ;
    output d_arr_16__27 ;
    output d_arr_16__26 ;
    output d_arr_16__25 ;
    output d_arr_16__24 ;
    output d_arr_16__23 ;
    output d_arr_16__22 ;
    output d_arr_16__21 ;
    output d_arr_16__20 ;
    output d_arr_16__19 ;
    output d_arr_16__18 ;
    output d_arr_16__17 ;
    output d_arr_16__16 ;
    output d_arr_16__15 ;
    output d_arr_16__14 ;
    output d_arr_16__13 ;
    output d_arr_16__12 ;
    output d_arr_16__11 ;
    output d_arr_16__10 ;
    output d_arr_16__9 ;
    output d_arr_16__8 ;
    output d_arr_16__7 ;
    output d_arr_16__6 ;
    output d_arr_16__5 ;
    output d_arr_16__4 ;
    output d_arr_16__3 ;
    output d_arr_16__2 ;
    output d_arr_16__1 ;
    output d_arr_16__0 ;
    output d_arr_17__31 ;
    output d_arr_17__30 ;
    output d_arr_17__29 ;
    output d_arr_17__28 ;
    output d_arr_17__27 ;
    output d_arr_17__26 ;
    output d_arr_17__25 ;
    output d_arr_17__24 ;
    output d_arr_17__23 ;
    output d_arr_17__22 ;
    output d_arr_17__21 ;
    output d_arr_17__20 ;
    output d_arr_17__19 ;
    output d_arr_17__18 ;
    output d_arr_17__17 ;
    output d_arr_17__16 ;
    output d_arr_17__15 ;
    output d_arr_17__14 ;
    output d_arr_17__13 ;
    output d_arr_17__12 ;
    output d_arr_17__11 ;
    output d_arr_17__10 ;
    output d_arr_17__9 ;
    output d_arr_17__8 ;
    output d_arr_17__7 ;
    output d_arr_17__6 ;
    output d_arr_17__5 ;
    output d_arr_17__4 ;
    output d_arr_17__3 ;
    output d_arr_17__2 ;
    output d_arr_17__1 ;
    output d_arr_17__0 ;
    output d_arr_18__31 ;
    output d_arr_18__30 ;
    output d_arr_18__29 ;
    output d_arr_18__28 ;
    output d_arr_18__27 ;
    output d_arr_18__26 ;
    output d_arr_18__25 ;
    output d_arr_18__24 ;
    output d_arr_18__23 ;
    output d_arr_18__22 ;
    output d_arr_18__21 ;
    output d_arr_18__20 ;
    output d_arr_18__19 ;
    output d_arr_18__18 ;
    output d_arr_18__17 ;
    output d_arr_18__16 ;
    output d_arr_18__15 ;
    output d_arr_18__14 ;
    output d_arr_18__13 ;
    output d_arr_18__12 ;
    output d_arr_18__11 ;
    output d_arr_18__10 ;
    output d_arr_18__9 ;
    output d_arr_18__8 ;
    output d_arr_18__7 ;
    output d_arr_18__6 ;
    output d_arr_18__5 ;
    output d_arr_18__4 ;
    output d_arr_18__3 ;
    output d_arr_18__2 ;
    output d_arr_18__1 ;
    output d_arr_18__0 ;
    output d_arr_19__31 ;
    output d_arr_19__30 ;
    output d_arr_19__29 ;
    output d_arr_19__28 ;
    output d_arr_19__27 ;
    output d_arr_19__26 ;
    output d_arr_19__25 ;
    output d_arr_19__24 ;
    output d_arr_19__23 ;
    output d_arr_19__22 ;
    output d_arr_19__21 ;
    output d_arr_19__20 ;
    output d_arr_19__19 ;
    output d_arr_19__18 ;
    output d_arr_19__17 ;
    output d_arr_19__16 ;
    output d_arr_19__15 ;
    output d_arr_19__14 ;
    output d_arr_19__13 ;
    output d_arr_19__12 ;
    output d_arr_19__11 ;
    output d_arr_19__10 ;
    output d_arr_19__9 ;
    output d_arr_19__8 ;
    output d_arr_19__7 ;
    output d_arr_19__6 ;
    output d_arr_19__5 ;
    output d_arr_19__4 ;
    output d_arr_19__3 ;
    output d_arr_19__2 ;
    output d_arr_19__1 ;
    output d_arr_19__0 ;
    output d_arr_20__31 ;
    output d_arr_20__30 ;
    output d_arr_20__29 ;
    output d_arr_20__28 ;
    output d_arr_20__27 ;
    output d_arr_20__26 ;
    output d_arr_20__25 ;
    output d_arr_20__24 ;
    output d_arr_20__23 ;
    output d_arr_20__22 ;
    output d_arr_20__21 ;
    output d_arr_20__20 ;
    output d_arr_20__19 ;
    output d_arr_20__18 ;
    output d_arr_20__17 ;
    output d_arr_20__16 ;
    output d_arr_20__15 ;
    output d_arr_20__14 ;
    output d_arr_20__13 ;
    output d_arr_20__12 ;
    output d_arr_20__11 ;
    output d_arr_20__10 ;
    output d_arr_20__9 ;
    output d_arr_20__8 ;
    output d_arr_20__7 ;
    output d_arr_20__6 ;
    output d_arr_20__5 ;
    output d_arr_20__4 ;
    output d_arr_20__3 ;
    output d_arr_20__2 ;
    output d_arr_20__1 ;
    output d_arr_20__0 ;
    output d_arr_21__31 ;
    output d_arr_21__30 ;
    output d_arr_21__29 ;
    output d_arr_21__28 ;
    output d_arr_21__27 ;
    output d_arr_21__26 ;
    output d_arr_21__25 ;
    output d_arr_21__24 ;
    output d_arr_21__23 ;
    output d_arr_21__22 ;
    output d_arr_21__21 ;
    output d_arr_21__20 ;
    output d_arr_21__19 ;
    output d_arr_21__18 ;
    output d_arr_21__17 ;
    output d_arr_21__16 ;
    output d_arr_21__15 ;
    output d_arr_21__14 ;
    output d_arr_21__13 ;
    output d_arr_21__12 ;
    output d_arr_21__11 ;
    output d_arr_21__10 ;
    output d_arr_21__9 ;
    output d_arr_21__8 ;
    output d_arr_21__7 ;
    output d_arr_21__6 ;
    output d_arr_21__5 ;
    output d_arr_21__4 ;
    output d_arr_21__3 ;
    output d_arr_21__2 ;
    output d_arr_21__1 ;
    output d_arr_21__0 ;
    output d_arr_22__31 ;
    output d_arr_22__30 ;
    output d_arr_22__29 ;
    output d_arr_22__28 ;
    output d_arr_22__27 ;
    output d_arr_22__26 ;
    output d_arr_22__25 ;
    output d_arr_22__24 ;
    output d_arr_22__23 ;
    output d_arr_22__22 ;
    output d_arr_22__21 ;
    output d_arr_22__20 ;
    output d_arr_22__19 ;
    output d_arr_22__18 ;
    output d_arr_22__17 ;
    output d_arr_22__16 ;
    output d_arr_22__15 ;
    output d_arr_22__14 ;
    output d_arr_22__13 ;
    output d_arr_22__12 ;
    output d_arr_22__11 ;
    output d_arr_22__10 ;
    output d_arr_22__9 ;
    output d_arr_22__8 ;
    output d_arr_22__7 ;
    output d_arr_22__6 ;
    output d_arr_22__5 ;
    output d_arr_22__4 ;
    output d_arr_22__3 ;
    output d_arr_22__2 ;
    output d_arr_22__1 ;
    output d_arr_22__0 ;
    output d_arr_23__31 ;
    output d_arr_23__30 ;
    output d_arr_23__29 ;
    output d_arr_23__28 ;
    output d_arr_23__27 ;
    output d_arr_23__26 ;
    output d_arr_23__25 ;
    output d_arr_23__24 ;
    output d_arr_23__23 ;
    output d_arr_23__22 ;
    output d_arr_23__21 ;
    output d_arr_23__20 ;
    output d_arr_23__19 ;
    output d_arr_23__18 ;
    output d_arr_23__17 ;
    output d_arr_23__16 ;
    output d_arr_23__15 ;
    output d_arr_23__14 ;
    output d_arr_23__13 ;
    output d_arr_23__12 ;
    output d_arr_23__11 ;
    output d_arr_23__10 ;
    output d_arr_23__9 ;
    output d_arr_23__8 ;
    output d_arr_23__7 ;
    output d_arr_23__6 ;
    output d_arr_23__5 ;
    output d_arr_23__4 ;
    output d_arr_23__3 ;
    output d_arr_23__2 ;
    output d_arr_23__1 ;
    output d_arr_23__0 ;
    output d_arr_24__31 ;
    output d_arr_24__30 ;
    output d_arr_24__29 ;
    output d_arr_24__28 ;
    output d_arr_24__27 ;
    output d_arr_24__26 ;
    output d_arr_24__25 ;
    output d_arr_24__24 ;
    output d_arr_24__23 ;
    output d_arr_24__22 ;
    output d_arr_24__21 ;
    output d_arr_24__20 ;
    output d_arr_24__19 ;
    output d_arr_24__18 ;
    output d_arr_24__17 ;
    output d_arr_24__16 ;
    output d_arr_24__15 ;
    output d_arr_24__14 ;
    output d_arr_24__13 ;
    output d_arr_24__12 ;
    output d_arr_24__11 ;
    output d_arr_24__10 ;
    output d_arr_24__9 ;
    output d_arr_24__8 ;
    output d_arr_24__7 ;
    output d_arr_24__6 ;
    output d_arr_24__5 ;
    output d_arr_24__4 ;
    output d_arr_24__3 ;
    output d_arr_24__2 ;
    output d_arr_24__1 ;
    output d_arr_24__0 ;

    wire nx4, nx8, nx12, nx18, nx28, nx36, nx44, nx52, nx60, nx68, nx76, nx84, 
         nx92, nx100, nx108, nx116, nx124, nx132, nx140, nx146, nx152, nx158, 
         nx164, nx170, nx176, nx182, nx188, nx194, nx200, nx206, nx212, nx218, 
         nx224, nx230, nx236, nx244, nx252, nx260, nx268, nx276, nx284, nx292, 
         nx300, nx308, nx316, nx324, nx332, nx340, nx348, nx356, nx364, nx370, 
         nx376, nx382, nx388, nx394, nx400, nx406, nx412, nx418, nx424, nx430, 
         nx436, nx442, nx448, nx454, nx460, nx468, nx476, nx484, nx492, nx500, 
         nx508, nx516, nx524, nx532, nx540, nx548, nx556, nx564, nx572, nx580, 
         nx588, nx594, nx600, nx606, nx612, nx618, nx624, nx630, nx636, nx642, 
         nx648, nx654, nx660, nx666, nx672, nx678, nx684, nx694, nx700, nx712, 
         nx724, nx736, nx748, nx760, nx772, nx784, nx796, nx808, nx820, nx832, 
         nx844, nx856, nx868, nx880, nx890, nx900, nx910, nx920, nx930, nx940, 
         nx950, nx960, nx970, nx980, nx990, nx1000, nx1010, nx1020, nx1030, 
         nx1040, nx1052, nx1064, nx1076, nx1088, nx1100, nx1112, nx1124, nx1136, 
         nx1148, nx1160, nx1172, nx1184, nx1196, nx1208, nx1220, nx1232, nx1242, 
         nx1252, nx1262, nx1272, nx1282, nx1292, nx1302, nx1312, nx1322, nx1332, 
         nx1342, nx1352, nx1362, nx1372, nx1382, nx1392, nx1404, nx1416, nx1428, 
         nx1440, nx1452, nx1464, nx1476, nx1488, nx1500, nx1512, nx1524, nx1536, 
         nx1548, nx1560, nx1572, nx1584, nx1594, nx1604, nx1614, nx1624, nx1634, 
         nx1644, nx1654, nx1664, nx1674, nx1684, nx1694, nx1704, nx1714, nx1724, 
         nx1734, nx1744, nx1756, nx1768, nx1780, nx1792, nx1804, nx1816, nx1828, 
         nx1840, nx1852, nx1864, nx1876, nx1888, nx1900, nx1912, nx1924, nx1936, 
         nx1946, nx1956, nx1966, nx1976, nx1986, nx1996, nx2006, nx2016, nx2026, 
         nx2036, nx2046, nx2056, nx2066, nx2076, nx2086, nx2096, nx2104, nx2112, 
         nx2120, nx2128, nx2136, nx2144, nx2152, nx2160, nx2168, nx2176, nx2184, 
         nx2192, nx2200, nx2208, nx2216, nx2224, nx2232, nx2240, nx2248, nx2256, 
         nx2264, nx2272, nx2280, nx2288, nx2296, nx2304, nx2312, nx2320, nx2328, 
         nx2336, nx2344, nx2352, nx2360, nx2368, nx2376, nx2384, nx2392, nx2400, 
         nx2408, nx2416, nx2424, nx2432, nx2440, nx2448, nx2456, nx2464, nx2472, 
         nx2480, nx2488, nx2496, nx2504, nx2512, nx2520, nx2528, nx2536, nx2544, 
         nx2552, nx2560, nx2568, nx2576, nx2584, nx2592, nx2600, nx2608, nx2616, 
         nx2624, nx2632, nx2640, nx2648, nx2656, nx2664, nx2672, nx2680, nx2688, 
         nx2696, nx2704, nx2712, nx2720, nx2728, nx2736, nx2744, nx2752, nx2760, 
         nx2768, nx2776, nx2784, nx2792, nx2800, nx2808, nx2816, nx2824, nx2832, 
         nx2840, nx2848, nx2856, nx2864, nx2872, nx2880, nx2888, nx2896, nx2904, 
         nx2912, nx2920, nx2928, nx2936, nx2944, nx2952, nx2960, nx2968, nx2976, 
         nx2984, nx2992, nx3000, nx3008, nx3016, nx3024, nx3032, nx3040, nx3048, 
         nx3056, nx3064, nx3072, nx3080, nx3088, nx3096, nx3104, nx3112, nx3120, 
         nx3132, nx3144, nx3156, nx3168, nx3180, nx3192, nx3204, nx3216, nx3228, 
         nx3240, nx3252, nx3264, nx3276, nx3288, nx3300, nx3312, nx3324, nx3336, 
         nx3348, nx3360, nx3372, nx3384, nx3396, nx3408, nx3420, nx3432, nx3444, 
         nx3456, nx3468, nx3480, nx3492, nx3504, nx3516, nx3528, nx3540, nx3552, 
         nx3564, nx3576, nx3588, nx3600, nx3612, nx3624, nx3636, nx3648, nx3660, 
         nx3672, nx3684, nx3696, nx3708, nx3720, nx3732, nx3744, nx3756, nx3768, 
         nx3780, nx3792, nx3804, nx3816, nx3828, nx3840, nx3852, nx3864, nx3876, 
         nx3888, nx3900, nx3912, nx3924, nx3936, nx3948, nx3960, nx3972, nx3984, 
         nx3996, nx4008, nx4020, nx4032, nx4044, nx4056, nx4068, nx4080, nx4092, 
         nx4104, nx4116, nx4128, nx4140, nx4152, nx4164, nx4176, nx4188, nx4200, 
         nx4212, nx4224, nx4236, nx4248, nx4260, nx4272, nx4284, nx4296, nx4308, 
         nx4320, nx4332, nx4344, nx4356, nx4368, nx4380, nx4392, nx4404, nx4416, 
         nx4428, nx4440, nx4452, nx4464, nx4476, nx4488, nx4500, nx4512, nx4524, 
         nx4536, nx4548, nx4560, nx4572, nx4584, nx4596, nx4608, nx4620, nx4632, 
         nx4644, nx4656, nx4668, nx4680, nx4692, nx4704, nx4716, nx4728, nx4740, 
         nx4752, nx4764, nx4776, nx4788, nx4800, nx4812, nx4824, nx4836, nx4848, 
         nx4860, nx4872, nx4884, nx4896, nx4908, nx4920, nx4932, nx4944, nx4956, 
         nx4968, nx4980, nx4992, nx5004, nx5016, nx5028, nx5040, nx5048, nx5056, 
         nx5064, nx5072, nx5080, nx5088, nx5096, nx5104, nx5112, nx5120, nx5128, 
         nx5136, nx5144, nx5152, nx5160, nx5168, nx5174, nx5180, nx5186, nx5192, 
         nx5198, nx5204, nx5210, nx5216, nx5222, nx5228, nx5234, nx5240, nx5246, 
         nx5252, nx5258, nx5264, nx5272, nx5280, nx5288, nx5296, nx5304, nx5312, 
         nx5320, nx5328, nx5336, nx5344, nx5352, nx5360, nx5368, nx5376, nx5384, 
         nx5392, nx5398, nx5404, nx5410, nx5416, nx5422, nx5428, nx5434, nx5440, 
         nx5446, nx5452, nx5458, nx5464, nx5470, nx5476, nx5482, nx5488, nx5496, 
         nx5504, nx5512, nx5520, nx5528, nx5536, nx5544, nx5552, nx5560, nx5568, 
         nx5576, nx5584, nx5592, nx5600, nx5608, nx5616, nx5622, nx5628, nx5634, 
         nx5640, nx5646, nx5652, nx5658, nx5664, nx5670, nx5676, nx5682, nx5688, 
         nx5694, nx5700, nx5706, nx5712, nx5720, nx5728, nx5736, nx5744, nx5752, 
         nx5760, nx5768, nx5776, nx5784, nx5792, nx5800, nx5808, nx5816, nx5824, 
         nx5832, nx5840, nx5846, nx5852, nx5858, nx5864, nx5870, nx5876, nx5882, 
         nx5888, nx5894, nx5900, nx5906, nx5912, nx5918, nx5924, nx5930, nx5936, 
         nx5948, nx5960, nx5972, nx5984, nx5996, nx6008, nx6020, nx6032, nx6044, 
         nx6056, nx6068, nx6080, nx6092, nx6104, nx6116, nx6128, nx6138, nx6148, 
         nx6158, nx6168, nx6178, nx6188, nx6198, nx6208, nx6218, nx6228, nx6238, 
         nx6248, nx6258, nx6268, nx6278, nx6288, nx6300, nx6312, nx6324, nx6336, 
         nx6348, nx6360, nx6372, nx6384, nx6396, nx6408, nx6420, nx6432, nx6444, 
         nx6456, nx6468, nx6480, nx6490, nx6500, nx6510, nx6520, nx6530, nx6540, 
         nx6550, nx6560, nx6570, nx6580, nx6590, nx6600, nx6610, nx6620, nx6630, 
         nx6640, nx6652, nx6664, nx6676, nx6688, nx6700, nx6712, nx6724, nx6736, 
         nx6748, nx6760, nx6772, nx6784, nx6796, nx6808, nx6820, nx6832, nx6842, 
         nx6852, nx6862, nx6872, nx6882, nx6892, nx6902, nx6912, nx6922, nx6932, 
         nx6942, nx6952, nx6962, nx6972, nx6982, nx6992, nx7002, nx7018, nx7028, 
         nx7036, nx7060, nx7084, nx7108, nx7132, nx7156, nx7180, nx7204, nx7228, 
         nx7252, nx7276, nx7300, nx7324, nx7348, nx7372, nx7392, nx7414, nx7436, 
         nx7458, nx7480, nx7502, nx7524, nx7546, nx7568, nx7590, nx7612, nx7634, 
         nx7656, nx7678, nx7700, nx7722, nx7744, nx7768, nx7792, nx7816, nx7840, 
         nx7864, nx7888, nx7912, nx7936, nx7960, nx7984, nx8008, nx8032, nx8056, 
         nx8080, nx8104, nx8124, nx8146, nx8168, nx8190, nx8212, nx8234, nx8256, 
         nx8278, nx8300, nx8322, nx8344, nx8366, nx8388, nx8410, nx8432, nx8454, 
         nx8476, nx7201, nx7205, nx7209, nx7215, nx7221, nx7227, nx7233, nx7239, 
         nx7245, nx7251, nx7257, nx7263, nx7269, nx7275, nx7281, nx7287, nx7293, 
         nx7295, nx7301, nx7305, nx7311, nx7317, nx7323, nx7329, nx7335, nx7341, 
         nx7347, nx7353, nx7359, nx7365, nx7371, nx7377, nx7383, nx7389, nx7395, 
         nx7401, nx7407, nx7413, nx7419, nx7425, nx7431, nx7437, nx7441, nx7447, 
         nx7453, nx7459, nx7463, nx7469, nx7475, nx7481, nx7483, nx7489, nx7495, 
         nx7501, nx7507, nx7513, nx7519, nx7525, nx7529, nx7535, nx7541, nx7547, 
         nx7551, nx7557, nx7563, nx7569, nx7573, nx7579, nx7585, nx7591, nx7595, 
         nx7601, nx7607, nx7613, nx7617, nx7623, nx7629, nx7635, nx7639, nx7645, 
         nx7651, nx7657, nx7661, nx7663, nx7669, nx7675, nx7681, nx7687, nx7693, 
         nx7699, nx7705, nx7711, nx7717, nx7723, nx7727, nx7733, nx7739, nx7745, 
         nx7749, nx7755, nx7761, nx7767, nx7773, nx7779, nx7785, nx7791, nx7797, 
         nx7803, nx7809, nx7815, nx7821, nx7827, nx7833, nx7839, nx7845, nx7851, 
         nx7853, nx7859, nx7865, nx7869, nx7875, nx7881, nx7887, nx7893, nx7899, 
         nx7905, nx7911, nx7917, nx7923, nx7929, nx7935, nx7941, nx7947, nx8423, 
         nx8429, nx8435, nx8441, nx8447, nx8453, nx8459, nx8465, nx8471, nx8477, 
         nx8481, nx8485, nx8489, nx8493, nx8497, nx8501, nx8505, nx8509, nx8513, 
         nx8517, nx8521, nx8525, nx8529, nx8533, nx8537, nx8541, nx8545, nx8549, 
         nx8553, nx8557, nx8561, nx8565, nx8569, nx8573, nx8577, nx8581, nx8585, 
         nx8589, nx8593, nx8597, nx8601, nx8605, nx8609, nx8613, nx8617, nx8621, 
         nx8625, nx8629, nx8633, nx8637, nx8641, nx8645, nx8649, nx8653, nx8657, 
         nx8661, nx8665, nx8669, nx8673, nx8677, nx8681, nx8685, nx8689, nx8693, 
         nx8697, nx8701, nx8705, nx8709, nx8713, nx8717, nx8721, nx8725, nx8729, 
         nx8733, nx8737, nx8741, nx8745, nx8749, nx8753, nx8757, nx8761, nx8765, 
         nx8769, nx8773, nx8777, nx8781, nx8785, nx8789, nx8793, nx8797, nx8801, 
         nx8805, nx8809, nx8813, nx8817, nx8821, nx8825, nx8829, nx8833, nx8837, 
         nx8841, nx8845, nx8849, nx8853, nx8857, nx8861, nx8865, nx8869, nx8873, 
         nx8877, nx8881, nx8885, nx8889, nx8893, nx8897, nx8901, nx8905, nx8909, 
         nx8913, nx8917, nx8921, nx8925, nx8929, nx8933, nx8937, nx8941, nx8945, 
         nx8949, nx8953, nx8957, nx8961, nx8965, nx8969, nx8973, nx8977, nx8981, 
         nx8985, nx8989, nx8993, nx8997, nx9001, nx9005, nx9009, nx9013, nx9017, 
         nx9021, nx9025, nx9029, nx9033, nx9037, nx9041, nx9045, nx9049, nx9053, 
         nx9057, nx9061, nx9065, nx9069, nx9073, nx9077, nx9341, nx9345, nx9349, 
         nx9353, nx9357, nx9361, nx9365, nx9369, nx9373, nx9377, nx9381, nx9385, 
         nx9389, nx9393, nx9397, nx9401, nx9403, nx9407, nx9411, nx9415, nx9419, 
         nx9423, nx9427, nx9431, nx9435, nx9439, nx9443, nx9447, nx9451, nx9455, 
         nx9459, nx9463, nx9467, nx9471, nx9475, nx9479, nx9483, nx9487, nx9491, 
         nx9495, nx9499, nx9503, nx9507, nx9511, nx9515, nx9519, nx9523, nx9527, 
         nx9531, nx9533, nx9537, nx9541, nx9545, nx9549, nx9553, nx9557, nx9561, 
         nx9565, nx9569, nx9573, nx9577, nx9581, nx9585, nx9589, nx9593, nx9597, 
         nx9601, nx9605, nx9609, nx9613, nx9617, nx9621, nx9625, nx9629, nx9633, 
         nx9637, nx9641, nx9645, nx9649, nx9653, nx9657, nx9661, nx9663, nx9667, 
         nx9671, nx9675, nx9679, nx9683, nx9687, nx9691, nx9695, nx9699, nx9703, 
         nx9707, nx9711, nx9715, nx9719, nx9723, nx9727, nx9731, nx9734, nx9737, 
         nx9739, nx9742, nx9746, nx9748, nx9752, nx9754, nx9758, nx9760, nx9764, 
         nx9766, nx9770, nx9772, nx9776, nx9778, nx9782, nx9784, nx9788, nx9790, 
         nx9794, nx9796, nx9800, nx9802, nx9806, nx9808, nx9812, nx9814, nx9818, 
         nx9820, nx9824, nx9826, nx9830, nx9832, nx9834, nx9838, nx9840, nx9844, 
         nx9846, nx9850, nx9852, nx9856, nx9858, nx9862, nx9864, nx9868, nx9870, 
         nx9874, nx9876, nx9880, nx9882, nx9886, nx9888, nx9892, nx9894, nx9898, 
         nx9900, nx9904, nx9906, nx9910, nx9912, nx9916, nx9918, nx9922, nx9924, 
         nx9928, nx9930, nx9934, nx9936, nx9940, nx9942, nx9946, nx9948, nx9952, 
         nx9954, nx9958, nx9960, nx9964, nx9966, nx9970, nx9972, nx9976, nx9978, 
         nx9982, nx9984, nx9988, nx9990, nx9994, nx9996, nx10000, nx10002, 
         nx10006, nx10008, nx10012, nx10014, nx10018, nx10020, nx10024, nx10026, 
         nx10028, nx10032, nx10034, nx10038, nx10040, nx10044, nx10046, nx10050, 
         nx10052, nx10056, nx10058, nx10062, nx10064, nx10068, nx10070, nx10074, 
         nx10076, nx10080, nx10082, nx10086, nx10088, nx10092, nx10094, nx10098, 
         nx10100, nx10104, nx10106, nx10110, nx10112, nx10116, nx10118, nx10122, 
         nx10124, nx10133, nx10135, nx10137, nx10139, nx10141, nx10143, nx10145, 
         nx10147, nx10149, nx10151, nx10153, nx10155, nx10157, nx10159, nx10161, 
         nx10163, nx10165, nx10167, nx10169, nx10171, nx10173, nx10175, nx10177, 
         nx10179, nx10181, nx10183, nx10185, nx10187, nx10189, nx10191, nx10193, 
         nx10195, nx10197, nx10199, nx10201, nx10203, nx10205, nx10207, nx10209, 
         nx10211, nx10213, nx10215, nx10217, nx10219, nx10221, nx10223, nx10225, 
         nx10227, nx10229, nx10231, nx10233, nx10235, nx10237, nx10239, nx10241, 
         nx10243, nx10245, nx10247, nx10249, nx10251, nx10253, nx10255, nx10257, 
         nx10259, nx10261, nx10263, nx10265, nx10267, nx10269, nx10271, nx10273, 
         nx10275, nx10277, nx10279, nx10281, nx10283, nx10285, nx10287, nx10289, 
         nx10291, nx10293, nx10295, nx10297, nx10299, nx10301, nx10303, nx10305, 
         nx10307, nx10309, nx10311, nx10313, nx10315, nx10317, nx10319, nx10321, 
         nx10323, nx10325, nx10327, nx10329, nx10331, nx10333, nx10335, nx10337, 
         nx10339, nx10341, nx10343, nx10345, nx10347, nx10349, nx10351, nx10353, 
         nx10355, nx10357, nx10359, nx10361, nx10365, nx10367, nx10369, nx10373, 
         nx10375, nx10377, nx10383, nx10385, nx10387, nx10391, nx10393, nx10395, 
         nx10397, nx10399, nx10401, nx10403, nx10405, nx10407, nx10409, nx10411, 
         nx10413, nx10415, nx10417, nx10419, nx10421, nx10423, nx10425, nx10427, 
         nx10429, nx10431, nx10433, nx10435, nx10437, nx10439, nx10441, nx10443, 
         nx10445, nx10447, nx10449, nx10451, nx10453, nx10455, nx10457, nx10459, 
         nx10461, nx10463, nx10465, nx10467, nx10469, nx10471, nx10473, nx10475, 
         nx10477, nx10479, nx10481, nx10483, nx10485, nx10487, nx10489, nx10491, 
         nx10493, nx10495, nx10497, nx10499, nx10501, nx10503, nx10505, nx10507, 
         nx10509, nx10511, nx10513, nx10515, nx10519, nx10521, nx10523, nx10529, 
         nx10531, nx10533, nx10537, nx10539, nx10541, nx10547, nx10549, nx10551, 
         nx10553, nx10555, nx10557, nx10559, nx10561, nx10563, nx10565, nx10567, 
         nx10569, nx10571, nx10573, nx10575, nx10577, nx10579, nx10581, nx10583, 
         nx10585, nx10587, nx10589, nx10591, nx10593, nx10595, nx10603, nx10611, 
         nx10621, nx10623, nx10625, nx10627, nx10629, nx10631, nx10633, nx10635, 
         nx10637, nx10639, nx10641, nx10643, nx10645, nx10647, nx10649, nx10651, 
         nx10653, nx10655, nx10657, nx10659, nx10661, nx10663, nx10665, nx10667, 
         nx10669, nx10671, nx10673, nx10675, nx10677, nx10679, nx10681, nx10683, 
         nx10685, nx10687, nx10689, nx10691, nx10693, nx10695, nx10697, nx10699, 
         nx10701, nx10703, nx10705, nx10707, nx10709, nx10711, nx10713, nx10715, 
         nx10717, nx10719, nx10721, nx10723, nx10725, nx10727, nx10729, nx10731, 
         nx10733, nx10735, nx10737, nx10739, nx10741, nx10743, nx10745, nx10747, 
         nx10749, nx10757, nx10765, nx10773, nx10781, nx10783, nx10785, nx10787, 
         nx10789, nx10791, nx10793, nx10795, nx10797, nx10799, nx10801, nx10803, 
         nx10805, nx10807, nx10809, nx10811, nx10813, nx10815, nx10817, nx10819, 
         nx10821, nx10823, nx10825, nx10827, nx10829, nx10831, nx10833, nx10835, 
         nx10837, nx10839, nx10841, nx10843, nx10845, nx10847, nx10849, nx10851, 
         nx10853, nx10855, nx10857, nx10859, nx10861, nx10863, nx10865, nx10867, 
         nx10869, nx10871, nx10873, nx10875, nx10877, nx10879, nx10881, nx10883, 
         nx10885, nx10887, nx10889, nx10891, nx10893, nx10895, nx10897, nx10899, 
         nx10901, nx10903, nx10905, nx10907, nx10909, nx10911, nx10913, nx10915, 
         nx10917, nx10919, nx10921, nx10923, nx10925, nx10927, nx10929, nx10931, 
         nx10933, nx10935, nx10937, nx10939, nx10941, nx10943, nx10945, nx10947, 
         nx10949, nx10951, nx10953, nx10955, nx10957, nx10959, nx10961, nx10963, 
         nx10965, nx10967, nx10969, nx10971, nx10973, nx10979, nx10981, nx10983, 
         nx10985, nx10987, nx10989, nx10991, nx10993, nx10995, nx10997, nx10999, 
         nx11005, nx11007, nx11009, nx11011, nx11013, nx11015, nx11017, nx11019, 
         nx11021, nx11023, nx11025, nx11027, nx11029, nx11031, nx11033, nx11035, 
         nx11037, nx11039, nx11041, nx11043, nx11045, nx11047, nx11049, nx11051, 
         nx11053, nx11055, nx11057, nx11059, nx11061, nx11063, nx11065, nx11067, 
         nx11069, nx11071, nx11073, nx11075, nx11077, nx11079, nx11081, nx11083, 
         nx11085, nx11087, nx11089, nx11091, nx11093, nx11095, nx11097, nx11099, 
         nx11101, nx11103, nx11105, nx11107, nx11109, nx11111, nx11113, nx11115, 
         nx11117, nx11119, nx11121, nx11123, nx11125, nx11127, nx11129, nx11131, 
         nx11133, nx11135, nx11137, nx11139, nx11141, nx11143, nx11145, nx11147, 
         nx11149, nx11151, nx11153, nx11155, nx11157, nx11159, nx11161, nx11163, 
         nx11165, nx11167, nx11169, nx11171, nx11173, nx11175, nx11177, nx11179, 
         nx11181, nx11183, nx11185, nx11187, nx11189, nx11191, nx11193, nx11195, 
         nx11197, nx11199, nx11201, nx11203, nx11205, nx11207, nx11209, nx11211, 
         nx11213, nx11215, nx11217, nx11219, nx11221, nx11223, nx11225, nx11227, 
         nx11229, nx11231, nx11233, nx11235, nx11237, nx11239, nx11241, nx11245, 
         nx11247, nx11249, nx11251, nx11253, nx11255, nx11257, nx11259, nx11261, 
         nx11263, nx11265, nx11267, nx11269, nx11271, nx11273, nx11275, nx11277, 
         nx11279, nx11281, nx11283, nx11285, nx11287, nx11289, nx11291, nx11293, 
         nx11295, nx11297, nx11299, nx11301, nx11303, nx11305, nx11307, nx11309, 
         nx11311, nx11313, nx11315, nx11317, nx11319, nx11321, nx11323, nx11325, 
         nx11327, nx11329, nx11331, nx11333, nx11335, nx11337, nx11339, nx11341, 
         nx11343, nx11345, nx11347, nx11349, nx11351, nx11353, nx11355, nx11357, 
         nx11359, nx11361, nx11363, nx11365, nx11367, nx11369, nx11371, nx11373, 
         nx11375, nx11377, nx11379, nx11381, nx11383, nx11385, nx11387, nx11389, 
         nx11391, nx11393, nx11395, nx11397, nx11399, nx11401, nx11403, nx11405, 
         nx11407, nx11409, nx11411, nx11413, nx11415, nx11417, nx11419, nx11421, 
         nx11423, nx11425, nx11427, nx11429, nx11431, nx11433, nx11435, nx11437, 
         nx11439, nx11441, nx11443, nx11445, nx11447, nx11449, nx11451, nx11453, 
         nx11455, nx11457, nx11459, nx11461, nx11463, nx11465, nx11467, nx11469, 
         nx11471, nx11473, nx11475, nx11477, nx11479, nx11481, nx11483, nx11485, 
         nx11487, nx11489, nx11491, nx11493, nx11495, nx11497, nx11499, nx11501, 
         nx11503, nx11505, nx11511, nx11517, nx11519, nx11524, nx11525;



    latch lat_d_arr_24__0 (.Q (d_arr_24__0), .D (nx18), .CLK (nx10133)) ;
    ao22 ix19 (.Y (nx18), .A0 (d_arr_mux_24__0), .A1 (nx11245), .B0 (
         d_arr_mul_24__0), .B1 (nx10365)) ;
    nor02ii ix13 (.Y (nx12), .A0 (nx11245), .A1 (sel_mul)) ;
    or03 ix9 (.Y (nx8), .A0 (sel_merge2), .A1 (sel_relu), .A2 (nx4)) ;
    latch lat_d_arr_24__1 (.Q (d_arr_24__1), .D (nx28), .CLK (nx10133)) ;
    ao22 ix29 (.Y (nx28), .A0 (d_arr_mux_24__1), .A1 (nx11245), .B0 (
         d_arr_mul_24__1), .B1 (nx10365)) ;
    latch lat_d_arr_24__2 (.Q (d_arr_24__2), .D (nx36), .CLK (nx10133)) ;
    ao22 ix37 (.Y (nx36), .A0 (d_arr_mux_24__2), .A1 (nx11245), .B0 (
         d_arr_mul_24__2), .B1 (nx10365)) ;
    latch lat_d_arr_24__3 (.Q (d_arr_24__3), .D (nx44), .CLK (nx10133)) ;
    ao22 ix45 (.Y (nx44), .A0 (d_arr_mux_24__3), .A1 (nx11245), .B0 (
         d_arr_mul_24__3), .B1 (nx10365)) ;
    latch lat_d_arr_24__4 (.Q (d_arr_24__4), .D (nx52), .CLK (nx10133)) ;
    ao22 ix53 (.Y (nx52), .A0 (d_arr_mux_24__4), .A1 (nx11245), .B0 (
         d_arr_mul_24__4), .B1 (nx10365)) ;
    latch lat_d_arr_24__5 (.Q (d_arr_24__5), .D (nx60), .CLK (nx10133)) ;
    ao22 ix61 (.Y (nx60), .A0 (d_arr_mux_24__5), .A1 (nx11245), .B0 (
         d_arr_mul_24__5), .B1 (nx10365)) ;
    latch lat_d_arr_24__6 (.Q (d_arr_24__6), .D (nx68), .CLK (nx10133)) ;
    ao22 ix69 (.Y (nx68), .A0 (d_arr_mux_24__6), .A1 (nx11247), .B0 (
         d_arr_mul_24__6), .B1 (nx10365)) ;
    latch lat_d_arr_24__7 (.Q (d_arr_24__7), .D (nx76), .CLK (nx10135)) ;
    ao22 ix77 (.Y (nx76), .A0 (d_arr_mux_24__7), .A1 (nx11247), .B0 (
         d_arr_mul_24__7), .B1 (nx10367)) ;
    latch lat_d_arr_24__8 (.Q (d_arr_24__8), .D (nx84), .CLK (nx10135)) ;
    ao22 ix85 (.Y (nx84), .A0 (d_arr_mux_24__8), .A1 (nx11247), .B0 (
         d_arr_mul_24__8), .B1 (nx10367)) ;
    latch lat_d_arr_24__9 (.Q (d_arr_24__9), .D (nx92), .CLK (nx10135)) ;
    ao22 ix93 (.Y (nx92), .A0 (d_arr_mux_24__9), .A1 (nx11247), .B0 (
         d_arr_mul_24__9), .B1 (nx10367)) ;
    latch lat_d_arr_24__10 (.Q (d_arr_24__10), .D (nx100), .CLK (nx10135)) ;
    ao22 ix101 (.Y (nx100), .A0 (d_arr_mux_24__10), .A1 (nx11247), .B0 (
         d_arr_mul_24__10), .B1 (nx10367)) ;
    latch lat_d_arr_24__11 (.Q (d_arr_24__11), .D (nx108), .CLK (nx10135)) ;
    ao22 ix109 (.Y (nx108), .A0 (d_arr_mux_24__11), .A1 (nx11247), .B0 (
         d_arr_mul_24__11), .B1 (nx10367)) ;
    latch lat_d_arr_24__12 (.Q (d_arr_24__12), .D (nx116), .CLK (nx10135)) ;
    ao22 ix117 (.Y (nx116), .A0 (d_arr_mux_24__12), .A1 (nx11247), .B0 (
         d_arr_mul_24__12), .B1 (nx10367)) ;
    latch lat_d_arr_24__13 (.Q (d_arr_24__13), .D (nx124), .CLK (nx10135)) ;
    ao22 ix125 (.Y (nx124), .A0 (d_arr_mux_24__13), .A1 (nx11249), .B0 (
         d_arr_mul_24__13), .B1 (nx10367)) ;
    latch lat_d_arr_24__14 (.Q (d_arr_24__14), .D (nx132), .CLK (nx10137)) ;
    ao22 ix133 (.Y (nx132), .A0 (d_arr_mux_24__14), .A1 (nx11249), .B0 (
         d_arr_mul_24__14), .B1 (nx10369)) ;
    latch lat_d_arr_24__15 (.Q (d_arr_24__15), .D (nx140), .CLK (nx10137)) ;
    latch lat_d_arr_24__16 (.Q (d_arr_24__16), .D (nx146), .CLK (nx10137)) ;
    latch lat_d_arr_24__17 (.Q (d_arr_24__17), .D (nx152), .CLK (nx10137)) ;
    latch lat_d_arr_24__18 (.Q (d_arr_24__18), .D (nx158), .CLK (nx10137)) ;
    latch lat_d_arr_24__19 (.Q (d_arr_24__19), .D (nx164), .CLK (nx10137)) ;
    latch lat_d_arr_24__20 (.Q (d_arr_24__20), .D (nx170), .CLK (nx10137)) ;
    latch lat_d_arr_24__21 (.Q (d_arr_24__21), .D (nx176), .CLK (nx10139)) ;
    latch lat_d_arr_24__22 (.Q (d_arr_24__22), .D (nx182), .CLK (nx10139)) ;
    latch lat_d_arr_24__23 (.Q (d_arr_24__23), .D (nx188), .CLK (nx10139)) ;
    latch lat_d_arr_24__24 (.Q (d_arr_24__24), .D (nx194), .CLK (nx10139)) ;
    latch lat_d_arr_24__25 (.Q (d_arr_24__25), .D (nx200), .CLK (nx10139)) ;
    latch lat_d_arr_24__26 (.Q (d_arr_24__26), .D (nx206), .CLK (nx10139)) ;
    latch lat_d_arr_24__27 (.Q (d_arr_24__27), .D (nx212), .CLK (nx10139)) ;
    latch lat_d_arr_24__28 (.Q (d_arr_24__28), .D (nx218), .CLK (nx10141)) ;
    latch lat_d_arr_24__29 (.Q (d_arr_24__29), .D (nx224), .CLK (nx10141)) ;
    latch lat_d_arr_24__30 (.Q (d_arr_24__30), .D (nx230), .CLK (nx10141)) ;
    latch lat_d_arr_24__31 (.Q (d_arr_24__31), .D (nx236), .CLK (nx10141)) ;
    latch lat_d_arr_23__0 (.Q (d_arr_23__0), .D (nx244), .CLK (nx10141)) ;
    ao22 ix245 (.Y (nx244), .A0 (d_arr_mux_23__0), .A1 (nx11249), .B0 (
         d_arr_mul_23__0), .B1 (nx10373)) ;
    latch lat_d_arr_23__1 (.Q (d_arr_23__1), .D (nx252), .CLK (nx10141)) ;
    ao22 ix253 (.Y (nx252), .A0 (d_arr_mux_23__1), .A1 (nx11249), .B0 (
         d_arr_mul_23__1), .B1 (nx10373)) ;
    latch lat_d_arr_23__2 (.Q (d_arr_23__2), .D (nx260), .CLK (nx10141)) ;
    ao22 ix261 (.Y (nx260), .A0 (d_arr_mux_23__2), .A1 (nx11249), .B0 (
         d_arr_mul_23__2), .B1 (nx10373)) ;
    latch lat_d_arr_23__3 (.Q (d_arr_23__3), .D (nx268), .CLK (nx10143)) ;
    ao22 ix269 (.Y (nx268), .A0 (d_arr_mux_23__3), .A1 (nx11249), .B0 (
         d_arr_mul_23__3), .B1 (nx10375)) ;
    latch lat_d_arr_23__4 (.Q (d_arr_23__4), .D (nx276), .CLK (nx10143)) ;
    ao22 ix277 (.Y (nx276), .A0 (d_arr_mux_23__4), .A1 (nx11249), .B0 (
         d_arr_mul_23__4), .B1 (nx10375)) ;
    latch lat_d_arr_23__5 (.Q (d_arr_23__5), .D (nx284), .CLK (nx10143)) ;
    ao22 ix285 (.Y (nx284), .A0 (d_arr_mux_23__5), .A1 (nx11251), .B0 (
         d_arr_mul_23__5), .B1 (nx10375)) ;
    latch lat_d_arr_23__6 (.Q (d_arr_23__6), .D (nx292), .CLK (nx10143)) ;
    ao22 ix293 (.Y (nx292), .A0 (d_arr_mux_23__6), .A1 (nx11251), .B0 (
         d_arr_mul_23__6), .B1 (nx10375)) ;
    latch lat_d_arr_23__7 (.Q (d_arr_23__7), .D (nx300), .CLK (nx10143)) ;
    ao22 ix301 (.Y (nx300), .A0 (d_arr_mux_23__7), .A1 (nx11251), .B0 (
         d_arr_mul_23__7), .B1 (nx10375)) ;
    latch lat_d_arr_23__8 (.Q (d_arr_23__8), .D (nx308), .CLK (nx10143)) ;
    ao22 ix309 (.Y (nx308), .A0 (d_arr_mux_23__8), .A1 (nx11251), .B0 (
         d_arr_mul_23__8), .B1 (nx10375)) ;
    latch lat_d_arr_23__9 (.Q (d_arr_23__9), .D (nx316), .CLK (nx10143)) ;
    ao22 ix317 (.Y (nx316), .A0 (d_arr_mux_23__9), .A1 (nx11251), .B0 (
         d_arr_mul_23__9), .B1 (nx10375)) ;
    latch lat_d_arr_23__10 (.Q (d_arr_23__10), .D (nx324), .CLK (nx10145)) ;
    ao22 ix325 (.Y (nx324), .A0 (d_arr_mux_23__10), .A1 (nx11251), .B0 (
         d_arr_mul_23__10), .B1 (nx10377)) ;
    latch lat_d_arr_23__11 (.Q (d_arr_23__11), .D (nx332), .CLK (nx10145)) ;
    ao22 ix333 (.Y (nx332), .A0 (d_arr_mux_23__11), .A1 (nx11251), .B0 (
         d_arr_mul_23__11), .B1 (nx10377)) ;
    latch lat_d_arr_23__12 (.Q (d_arr_23__12), .D (nx340), .CLK (nx10145)) ;
    ao22 ix341 (.Y (nx340), .A0 (d_arr_mux_23__12), .A1 (nx11253), .B0 (
         d_arr_mul_23__12), .B1 (nx10377)) ;
    latch lat_d_arr_23__13 (.Q (d_arr_23__13), .D (nx348), .CLK (nx10145)) ;
    ao22 ix349 (.Y (nx348), .A0 (d_arr_mux_23__13), .A1 (nx11253), .B0 (
         d_arr_mul_23__13), .B1 (nx10377)) ;
    latch lat_d_arr_23__14 (.Q (d_arr_23__14), .D (nx356), .CLK (nx10145)) ;
    ao22 ix357 (.Y (nx356), .A0 (d_arr_mux_23__14), .A1 (nx11253), .B0 (
         d_arr_mul_23__14), .B1 (nx10377)) ;
    latch lat_d_arr_23__15 (.Q (d_arr_23__15), .D (nx364), .CLK (nx10145)) ;
    latch lat_d_arr_23__16 (.Q (d_arr_23__16), .D (nx370), .CLK (nx10145)) ;
    latch lat_d_arr_23__17 (.Q (d_arr_23__17), .D (nx376), .CLK (nx10147)) ;
    latch lat_d_arr_23__18 (.Q (d_arr_23__18), .D (nx382), .CLK (nx10147)) ;
    latch lat_d_arr_23__19 (.Q (d_arr_23__19), .D (nx388), .CLK (nx10147)) ;
    latch lat_d_arr_23__20 (.Q (d_arr_23__20), .D (nx394), .CLK (nx10147)) ;
    latch lat_d_arr_23__21 (.Q (d_arr_23__21), .D (nx400), .CLK (nx10147)) ;
    latch lat_d_arr_23__22 (.Q (d_arr_23__22), .D (nx406), .CLK (nx10147)) ;
    latch lat_d_arr_23__23 (.Q (d_arr_23__23), .D (nx412), .CLK (nx10147)) ;
    latch lat_d_arr_23__24 (.Q (d_arr_23__24), .D (nx418), .CLK (nx10149)) ;
    latch lat_d_arr_23__25 (.Q (d_arr_23__25), .D (nx424), .CLK (nx10149)) ;
    latch lat_d_arr_23__26 (.Q (d_arr_23__26), .D (nx430), .CLK (nx10149)) ;
    latch lat_d_arr_23__27 (.Q (d_arr_23__27), .D (nx436), .CLK (nx10149)) ;
    latch lat_d_arr_23__28 (.Q (d_arr_23__28), .D (nx442), .CLK (nx10149)) ;
    latch lat_d_arr_23__29 (.Q (d_arr_23__29), .D (nx448), .CLK (nx10149)) ;
    latch lat_d_arr_23__30 (.Q (d_arr_23__30), .D (nx454), .CLK (nx10149)) ;
    latch lat_d_arr_23__31 (.Q (d_arr_23__31), .D (nx460), .CLK (nx10151)) ;
    latch lat_d_arr_22__0 (.Q (d_arr_22__0), .D (nx468), .CLK (nx10151)) ;
    ao22 ix469 (.Y (nx468), .A0 (d_arr_mux_22__0), .A1 (nx11253), .B0 (
         d_arr_mul_22__0), .B1 (nx10383)) ;
    latch lat_d_arr_22__1 (.Q (d_arr_22__1), .D (nx476), .CLK (nx10151)) ;
    ao22 ix477 (.Y (nx476), .A0 (d_arr_mux_22__1), .A1 (nx11253), .B0 (
         d_arr_mul_22__1), .B1 (nx10383)) ;
    latch lat_d_arr_22__2 (.Q (d_arr_22__2), .D (nx484), .CLK (nx10151)) ;
    ao22 ix485 (.Y (nx484), .A0 (d_arr_mux_22__2), .A1 (nx11253), .B0 (
         d_arr_mul_22__2), .B1 (nx10383)) ;
    latch lat_d_arr_22__3 (.Q (d_arr_22__3), .D (nx492), .CLK (nx10151)) ;
    ao22 ix493 (.Y (nx492), .A0 (d_arr_mux_22__3), .A1 (nx11253), .B0 (
         d_arr_mul_22__3), .B1 (nx10383)) ;
    latch lat_d_arr_22__4 (.Q (d_arr_22__4), .D (nx500), .CLK (nx10151)) ;
    ao22 ix501 (.Y (nx500), .A0 (d_arr_mux_22__4), .A1 (nx11255), .B0 (
         d_arr_mul_22__4), .B1 (nx10383)) ;
    latch lat_d_arr_22__5 (.Q (d_arr_22__5), .D (nx508), .CLK (nx10151)) ;
    ao22 ix509 (.Y (nx508), .A0 (d_arr_mux_22__5), .A1 (nx11255), .B0 (
         d_arr_mul_22__5), .B1 (nx10383)) ;
    latch lat_d_arr_22__6 (.Q (d_arr_22__6), .D (nx516), .CLK (nx10153)) ;
    ao22 ix517 (.Y (nx516), .A0 (d_arr_mux_22__6), .A1 (nx11255), .B0 (
         d_arr_mul_22__6), .B1 (nx10385)) ;
    latch lat_d_arr_22__7 (.Q (d_arr_22__7), .D (nx524), .CLK (nx10153)) ;
    ao22 ix525 (.Y (nx524), .A0 (d_arr_mux_22__7), .A1 (nx11255), .B0 (
         d_arr_mul_22__7), .B1 (nx10385)) ;
    latch lat_d_arr_22__8 (.Q (d_arr_22__8), .D (nx532), .CLK (nx10153)) ;
    ao22 ix533 (.Y (nx532), .A0 (d_arr_mux_22__8), .A1 (nx11255), .B0 (
         d_arr_mul_22__8), .B1 (nx10385)) ;
    latch lat_d_arr_22__9 (.Q (d_arr_22__9), .D (nx540), .CLK (nx10153)) ;
    ao22 ix541 (.Y (nx540), .A0 (d_arr_mux_22__9), .A1 (nx11255), .B0 (
         d_arr_mul_22__9), .B1 (nx10385)) ;
    latch lat_d_arr_22__10 (.Q (d_arr_22__10), .D (nx548), .CLK (nx10153)) ;
    ao22 ix549 (.Y (nx548), .A0 (d_arr_mux_22__10), .A1 (nx11255), .B0 (
         d_arr_mul_22__10), .B1 (nx10385)) ;
    latch lat_d_arr_22__11 (.Q (d_arr_22__11), .D (nx556), .CLK (nx10153)) ;
    ao22 ix557 (.Y (nx556), .A0 (d_arr_mux_22__11), .A1 (nx11257), .B0 (
         d_arr_mul_22__11), .B1 (nx10385)) ;
    latch lat_d_arr_22__12 (.Q (d_arr_22__12), .D (nx564), .CLK (nx10153)) ;
    ao22 ix565 (.Y (nx564), .A0 (d_arr_mux_22__12), .A1 (nx11257), .B0 (
         d_arr_mul_22__12), .B1 (nx10385)) ;
    latch lat_d_arr_22__13 (.Q (d_arr_22__13), .D (nx572), .CLK (nx10155)) ;
    ao22 ix573 (.Y (nx572), .A0 (d_arr_mux_22__13), .A1 (nx11257), .B0 (
         d_arr_mul_22__13), .B1 (nx10387)) ;
    latch lat_d_arr_22__14 (.Q (d_arr_22__14), .D (nx580), .CLK (nx10155)) ;
    ao22 ix581 (.Y (nx580), .A0 (d_arr_mux_22__14), .A1 (nx11257), .B0 (
         d_arr_mul_22__14), .B1 (nx10387)) ;
    latch lat_d_arr_22__15 (.Q (d_arr_22__15), .D (nx588), .CLK (nx10155)) ;
    latch lat_d_arr_22__16 (.Q (d_arr_22__16), .D (nx594), .CLK (nx10155)) ;
    latch lat_d_arr_22__17 (.Q (d_arr_22__17), .D (nx600), .CLK (nx10155)) ;
    latch lat_d_arr_22__18 (.Q (d_arr_22__18), .D (nx606), .CLK (nx10155)) ;
    latch lat_d_arr_22__19 (.Q (d_arr_22__19), .D (nx612), .CLK (nx10155)) ;
    latch lat_d_arr_22__20 (.Q (d_arr_22__20), .D (nx618), .CLK (nx10157)) ;
    latch lat_d_arr_22__21 (.Q (d_arr_22__21), .D (nx624), .CLK (nx10157)) ;
    latch lat_d_arr_22__22 (.Q (d_arr_22__22), .D (nx630), .CLK (nx10157)) ;
    latch lat_d_arr_22__23 (.Q (d_arr_22__23), .D (nx636), .CLK (nx10157)) ;
    latch lat_d_arr_22__24 (.Q (d_arr_22__24), .D (nx642), .CLK (nx10157)) ;
    latch lat_d_arr_22__25 (.Q (d_arr_22__25), .D (nx648), .CLK (nx10157)) ;
    latch lat_d_arr_22__26 (.Q (d_arr_22__26), .D (nx654), .CLK (nx10157)) ;
    latch lat_d_arr_22__27 (.Q (d_arr_22__27), .D (nx660), .CLK (nx10159)) ;
    latch lat_d_arr_22__28 (.Q (d_arr_22__28), .D (nx666), .CLK (nx10159)) ;
    latch lat_d_arr_22__29 (.Q (d_arr_22__29), .D (nx672), .CLK (nx10159)) ;
    latch lat_d_arr_22__30 (.Q (d_arr_22__30), .D (nx678), .CLK (nx10159)) ;
    latch lat_d_arr_22__31 (.Q (d_arr_22__31), .D (nx684), .CLK (nx10159)) ;
    latch lat_d_arr_21__0 (.Q (d_arr_21__0), .D (nx700), .CLK (nx10159)) ;
    inv01 ix701 (.Y (nx700), .A (nx7201)) ;
    aoi222 ix7202 (.Y (nx7201), .A0 (d_arr_mux_21__0), .A1 (nx11257), .B0 (
           d_arr_mul_21__0), .B1 (nx10391), .C0 (d_arr_add_21__0), .C1 (nx10621)
           ) ;
    nor03_2x ix695 (.Y (nx694), .A0 (nx7205), .A1 (nx11257), .A2 (sel_mul)) ;
    inv01 ix7206 (.Y (nx7205), .A (sel_add)) ;
    latch lat_d_arr_21__1 (.Q (d_arr_21__1), .D (nx712), .CLK (nx10159)) ;
    inv01 ix713 (.Y (nx712), .A (nx7209)) ;
    aoi222 ix7210 (.Y (nx7209), .A0 (d_arr_mux_21__1), .A1 (nx11257), .B0 (
           d_arr_mul_21__1), .B1 (nx10391), .C0 (d_arr_add_21__1), .C1 (nx10621)
           ) ;
    latch lat_d_arr_21__2 (.Q (d_arr_21__2), .D (nx724), .CLK (nx10161)) ;
    inv01 ix725 (.Y (nx724), .A (nx7215)) ;
    aoi222 ix7216 (.Y (nx7215), .A0 (d_arr_mux_21__2), .A1 (nx11259), .B0 (
           d_arr_mul_21__2), .B1 (nx10393), .C0 (d_arr_add_21__2), .C1 (nx10621)
           ) ;
    latch lat_d_arr_21__3 (.Q (d_arr_21__3), .D (nx736), .CLK (nx10161)) ;
    inv01 ix737 (.Y (nx736), .A (nx7221)) ;
    aoi222 ix7222 (.Y (nx7221), .A0 (d_arr_mux_21__3), .A1 (nx11259), .B0 (
           d_arr_mul_21__3), .B1 (nx10393), .C0 (d_arr_add_21__3), .C1 (nx10621)
           ) ;
    latch lat_d_arr_21__4 (.Q (d_arr_21__4), .D (nx748), .CLK (nx10161)) ;
    inv01 ix749 (.Y (nx748), .A (nx7227)) ;
    aoi222 ix7228 (.Y (nx7227), .A0 (d_arr_mux_21__4), .A1 (nx11259), .B0 (
           d_arr_mul_21__4), .B1 (nx10393), .C0 (d_arr_add_21__4), .C1 (nx10621)
           ) ;
    latch lat_d_arr_21__5 (.Q (d_arr_21__5), .D (nx760), .CLK (nx10161)) ;
    inv01 ix761 (.Y (nx760), .A (nx7233)) ;
    aoi222 ix7234 (.Y (nx7233), .A0 (d_arr_mux_21__5), .A1 (nx11259), .B0 (
           d_arr_mul_21__5), .B1 (nx10393), .C0 (d_arr_add_21__5), .C1 (nx10621)
           ) ;
    latch lat_d_arr_21__6 (.Q (d_arr_21__6), .D (nx772), .CLK (nx10161)) ;
    inv01 ix773 (.Y (nx772), .A (nx7239)) ;
    aoi222 ix7240 (.Y (nx7239), .A0 (d_arr_mux_21__6), .A1 (nx11259), .B0 (
           d_arr_mul_21__6), .B1 (nx10393), .C0 (d_arr_add_21__6), .C1 (nx10621)
           ) ;
    latch lat_d_arr_21__7 (.Q (d_arr_21__7), .D (nx784), .CLK (nx10161)) ;
    inv01 ix785 (.Y (nx784), .A (nx7245)) ;
    aoi222 ix7246 (.Y (nx7245), .A0 (d_arr_mux_21__7), .A1 (nx11259), .B0 (
           d_arr_mul_21__7), .B1 (nx10393), .C0 (d_arr_add_21__7), .C1 (nx10623)
           ) ;
    latch lat_d_arr_21__8 (.Q (d_arr_21__8), .D (nx796), .CLK (nx10161)) ;
    inv01 ix797 (.Y (nx796), .A (nx7251)) ;
    aoi222 ix7252 (.Y (nx7251), .A0 (d_arr_mux_21__8), .A1 (nx11259), .B0 (
           d_arr_mul_21__8), .B1 (nx10393), .C0 (d_arr_add_21__8), .C1 (nx10623)
           ) ;
    latch lat_d_arr_21__9 (.Q (d_arr_21__9), .D (nx808), .CLK (nx10163)) ;
    inv01 ix809 (.Y (nx808), .A (nx7257)) ;
    aoi222 ix7258 (.Y (nx7257), .A0 (d_arr_mux_21__9), .A1 (nx11261), .B0 (
           d_arr_mul_21__9), .B1 (nx10395), .C0 (d_arr_add_21__9), .C1 (nx10623)
           ) ;
    latch lat_d_arr_21__10 (.Q (d_arr_21__10), .D (nx820), .CLK (nx10163)) ;
    inv01 ix821 (.Y (nx820), .A (nx7263)) ;
    aoi222 ix7264 (.Y (nx7263), .A0 (d_arr_mux_21__10), .A1 (nx11261), .B0 (
           d_arr_mul_21__10), .B1 (nx10395), .C0 (d_arr_add_21__10), .C1 (
           nx10623)) ;
    latch lat_d_arr_21__11 (.Q (d_arr_21__11), .D (nx832), .CLK (nx10163)) ;
    inv01 ix833 (.Y (nx832), .A (nx7269)) ;
    aoi222 ix7270 (.Y (nx7269), .A0 (d_arr_mux_21__11), .A1 (nx11261), .B0 (
           d_arr_mul_21__11), .B1 (nx10395), .C0 (d_arr_add_21__11), .C1 (
           nx10623)) ;
    latch lat_d_arr_21__12 (.Q (d_arr_21__12), .D (nx844), .CLK (nx10163)) ;
    inv01 ix845 (.Y (nx844), .A (nx7275)) ;
    aoi222 ix7276 (.Y (nx7275), .A0 (d_arr_mux_21__12), .A1 (nx11261), .B0 (
           d_arr_mul_21__12), .B1 (nx10395), .C0 (d_arr_add_21__12), .C1 (
           nx10623)) ;
    latch lat_d_arr_21__13 (.Q (d_arr_21__13), .D (nx856), .CLK (nx10163)) ;
    inv01 ix857 (.Y (nx856), .A (nx7281)) ;
    aoi222 ix7282 (.Y (nx7281), .A0 (d_arr_mux_21__13), .A1 (nx11261), .B0 (
           d_arr_mul_21__13), .B1 (nx10395), .C0 (d_arr_add_21__13), .C1 (
           nx10623)) ;
    latch lat_d_arr_21__14 (.Q (d_arr_21__14), .D (nx868), .CLK (nx10163)) ;
    inv01 ix869 (.Y (nx868), .A (nx7287)) ;
    aoi222 ix7288 (.Y (nx7287), .A0 (d_arr_mux_21__14), .A1 (nx11261), .B0 (
           d_arr_mul_21__14), .B1 (nx10395), .C0 (d_arr_add_21__14), .C1 (
           nx10625)) ;
    latch lat_d_arr_21__15 (.Q (d_arr_21__15), .D (nx880), .CLK (nx10163)) ;
    nand02 ix881 (.Y (nx880), .A0 (nx7293), .A1 (nx10845)) ;
    aoi22 ix7294 (.Y (nx7293), .A0 (d_arr_mul_21__15), .A1 (nx10395), .B0 (
          d_arr_add_21__15), .B1 (nx10625)) ;
    nand02 ix7296 (.Y (nx7295), .A0 (d_arr_mux_21__31), .A1 (nx11261)) ;
    latch lat_d_arr_21__16 (.Q (d_arr_21__16), .D (nx890), .CLK (nx10165)) ;
    nand02 ix891 (.Y (nx890), .A0 (nx7301), .A1 (nx10845)) ;
    aoi22 ix7302 (.Y (nx7301), .A0 (d_arr_mul_21__16), .A1 (nx10397), .B0 (
          d_arr_add_21__16), .B1 (nx10625)) ;
    latch lat_d_arr_21__17 (.Q (d_arr_21__17), .D (nx900), .CLK (nx10165)) ;
    nand02 ix901 (.Y (nx900), .A0 (nx7305), .A1 (nx10845)) ;
    aoi22 ix7306 (.Y (nx7305), .A0 (d_arr_mul_21__17), .A1 (nx10397), .B0 (
          d_arr_add_21__17), .B1 (nx10625)) ;
    latch lat_d_arr_21__18 (.Q (d_arr_21__18), .D (nx910), .CLK (nx10165)) ;
    nand02 ix911 (.Y (nx910), .A0 (nx7311), .A1 (nx10845)) ;
    aoi22 ix7312 (.Y (nx7311), .A0 (d_arr_mul_21__18), .A1 (nx10397), .B0 (
          d_arr_add_21__18), .B1 (nx10625)) ;
    latch lat_d_arr_21__19 (.Q (d_arr_21__19), .D (nx920), .CLK (nx10165)) ;
    nand02 ix921 (.Y (nx920), .A0 (nx7317), .A1 (nx10845)) ;
    aoi22 ix7318 (.Y (nx7317), .A0 (d_arr_mul_21__19), .A1 (nx10397), .B0 (
          d_arr_add_21__19), .B1 (nx10625)) ;
    latch lat_d_arr_21__20 (.Q (d_arr_21__20), .D (nx930), .CLK (nx10165)) ;
    nand02 ix931 (.Y (nx930), .A0 (nx7323), .A1 (nx10845)) ;
    aoi22 ix7324 (.Y (nx7323), .A0 (d_arr_mul_21__20), .A1 (nx10397), .B0 (
          d_arr_add_21__20), .B1 (nx10625)) ;
    latch lat_d_arr_21__21 (.Q (d_arr_21__21), .D (nx940), .CLK (nx10165)) ;
    nand02 ix941 (.Y (nx940), .A0 (nx7329), .A1 (nx10845)) ;
    aoi22 ix7330 (.Y (nx7329), .A0 (d_arr_mul_21__21), .A1 (nx10397), .B0 (
          d_arr_add_21__21), .B1 (nx10627)) ;
    latch lat_d_arr_21__22 (.Q (d_arr_21__22), .D (nx950), .CLK (nx10165)) ;
    nand02 ix951 (.Y (nx950), .A0 (nx7335), .A1 (nx10847)) ;
    aoi22 ix7336 (.Y (nx7335), .A0 (d_arr_mul_21__22), .A1 (nx10397), .B0 (
          d_arr_add_21__22), .B1 (nx10627)) ;
    latch lat_d_arr_21__23 (.Q (d_arr_21__23), .D (nx960), .CLK (nx10167)) ;
    nand02 ix961 (.Y (nx960), .A0 (nx7341), .A1 (nx10847)) ;
    aoi22 ix7342 (.Y (nx7341), .A0 (d_arr_mul_21__23), .A1 (nx10399), .B0 (
          d_arr_add_21__23), .B1 (nx10627)) ;
    latch lat_d_arr_21__24 (.Q (d_arr_21__24), .D (nx970), .CLK (nx10167)) ;
    nand02 ix971 (.Y (nx970), .A0 (nx7347), .A1 (nx10847)) ;
    aoi22 ix7348 (.Y (nx7347), .A0 (d_arr_mul_21__24), .A1 (nx10399), .B0 (
          d_arr_add_21__24), .B1 (nx10627)) ;
    latch lat_d_arr_21__25 (.Q (d_arr_21__25), .D (nx980), .CLK (nx10167)) ;
    nand02 ix981 (.Y (nx980), .A0 (nx7353), .A1 (nx10847)) ;
    aoi22 ix7354 (.Y (nx7353), .A0 (d_arr_mul_21__25), .A1 (nx10399), .B0 (
          d_arr_add_21__25), .B1 (nx10627)) ;
    latch lat_d_arr_21__26 (.Q (d_arr_21__26), .D (nx990), .CLK (nx10167)) ;
    nand02 ix991 (.Y (nx990), .A0 (nx7359), .A1 (nx10847)) ;
    aoi22 ix7360 (.Y (nx7359), .A0 (d_arr_mul_21__26), .A1 (nx10399), .B0 (
          d_arr_add_21__26), .B1 (nx10627)) ;
    latch lat_d_arr_21__27 (.Q (d_arr_21__27), .D (nx1000), .CLK (nx10167)) ;
    nand02 ix1001 (.Y (nx1000), .A0 (nx7365), .A1 (nx10847)) ;
    aoi22 ix7366 (.Y (nx7365), .A0 (d_arr_mul_21__27), .A1 (nx10399), .B0 (
          d_arr_add_21__27), .B1 (nx10627)) ;
    latch lat_d_arr_21__28 (.Q (d_arr_21__28), .D (nx1010), .CLK (nx10167)) ;
    nand02 ix1011 (.Y (nx1010), .A0 (nx7371), .A1 (nx10847)) ;
    aoi22 ix7372 (.Y (nx7371), .A0 (d_arr_mul_21__28), .A1 (nx10399), .B0 (
          d_arr_add_21__28), .B1 (nx10629)) ;
    latch lat_d_arr_21__29 (.Q (d_arr_21__29), .D (nx1020), .CLK (nx10167)) ;
    nand02 ix1021 (.Y (nx1020), .A0 (nx7377), .A1 (nx7295)) ;
    aoi22 ix7378 (.Y (nx7377), .A0 (d_arr_mul_21__29), .A1 (nx10399), .B0 (
          d_arr_add_21__29), .B1 (nx10629)) ;
    latch lat_d_arr_21__30 (.Q (d_arr_21__30), .D (nx1030), .CLK (nx10169)) ;
    nand02 ix1031 (.Y (nx1030), .A0 (nx7383), .A1 (nx7295)) ;
    aoi22 ix7384 (.Y (nx7383), .A0 (d_arr_mul_21__30), .A1 (nx10401), .B0 (
          d_arr_add_21__30), .B1 (nx10629)) ;
    latch lat_d_arr_21__31 (.Q (d_arr_21__31), .D (nx1040), .CLK (nx10169)) ;
    nand02 ix1041 (.Y (nx1040), .A0 (nx7389), .A1 (nx7295)) ;
    aoi22 ix7390 (.Y (nx7389), .A0 (d_arr_mul_21__31), .A1 (nx10401), .B0 (
          d_arr_add_21__31), .B1 (nx10629)) ;
    latch lat_d_arr_20__0 (.Q (d_arr_20__0), .D (nx1052), .CLK (nx10169)) ;
    inv01 ix1053 (.Y (nx1052), .A (nx7395)) ;
    aoi222 ix7396 (.Y (nx7395), .A0 (d_arr_mux_20__0), .A1 (nx11263), .B0 (
           d_arr_mul_20__0), .B1 (nx10401), .C0 (d_arr_add_20__0), .C1 (nx10629)
           ) ;
    latch lat_d_arr_20__1 (.Q (d_arr_20__1), .D (nx1064), .CLK (nx10169)) ;
    inv01 ix1065 (.Y (nx1064), .A (nx7401)) ;
    aoi222 ix7402 (.Y (nx7401), .A0 (d_arr_mux_20__1), .A1 (nx11263), .B0 (
           d_arr_mul_20__1), .B1 (nx10401), .C0 (d_arr_add_20__1), .C1 (nx10629)
           ) ;
    latch lat_d_arr_20__2 (.Q (d_arr_20__2), .D (nx1076), .CLK (nx10169)) ;
    inv01 ix1077 (.Y (nx1076), .A (nx7407)) ;
    aoi222 ix7408 (.Y (nx7407), .A0 (d_arr_mux_20__2), .A1 (nx11263), .B0 (
           d_arr_mul_20__2), .B1 (nx10401), .C0 (d_arr_add_20__2), .C1 (nx10629)
           ) ;
    latch lat_d_arr_20__3 (.Q (d_arr_20__3), .D (nx1088), .CLK (nx10169)) ;
    inv01 ix1089 (.Y (nx1088), .A (nx7413)) ;
    aoi222 ix7414 (.Y (nx7413), .A0 (d_arr_mux_20__3), .A1 (nx11263), .B0 (
           d_arr_mul_20__3), .B1 (nx10401), .C0 (d_arr_add_20__3), .C1 (nx10631)
           ) ;
    latch lat_d_arr_20__4 (.Q (d_arr_20__4), .D (nx1100), .CLK (nx10169)) ;
    inv01 ix1101 (.Y (nx1100), .A (nx7419)) ;
    aoi222 ix7420 (.Y (nx7419), .A0 (d_arr_mux_20__4), .A1 (nx11263), .B0 (
           d_arr_mul_20__4), .B1 (nx10401), .C0 (d_arr_add_20__4), .C1 (nx10631)
           ) ;
    latch lat_d_arr_20__5 (.Q (d_arr_20__5), .D (nx1112), .CLK (nx10171)) ;
    inv01 ix1113 (.Y (nx1112), .A (nx7425)) ;
    aoi222 ix7426 (.Y (nx7425), .A0 (d_arr_mux_20__5), .A1 (nx11263), .B0 (
           d_arr_mul_20__5), .B1 (nx10403), .C0 (d_arr_add_20__5), .C1 (nx10631)
           ) ;
    latch lat_d_arr_20__6 (.Q (d_arr_20__6), .D (nx1124), .CLK (nx10171)) ;
    inv01 ix1125 (.Y (nx1124), .A (nx7431)) ;
    aoi222 ix7432 (.Y (nx7431), .A0 (d_arr_mux_20__6), .A1 (nx11263), .B0 (
           d_arr_mul_20__6), .B1 (nx10403), .C0 (d_arr_add_20__6), .C1 (nx10631)
           ) ;
    latch lat_d_arr_20__7 (.Q (d_arr_20__7), .D (nx1136), .CLK (nx10171)) ;
    inv01 ix1137 (.Y (nx1136), .A (nx7437)) ;
    aoi222 ix7438 (.Y (nx7437), .A0 (d_arr_mux_20__7), .A1 (nx11265), .B0 (
           d_arr_mul_20__7), .B1 (nx10403), .C0 (d_arr_add_20__7), .C1 (nx10631)
           ) ;
    latch lat_d_arr_20__8 (.Q (d_arr_20__8), .D (nx1148), .CLK (nx10171)) ;
    inv01 ix1149 (.Y (nx1148), .A (nx7441)) ;
    aoi222 ix7442 (.Y (nx7441), .A0 (d_arr_mux_20__8), .A1 (nx11265), .B0 (
           d_arr_mul_20__8), .B1 (nx10403), .C0 (d_arr_add_20__8), .C1 (nx10631)
           ) ;
    latch lat_d_arr_20__9 (.Q (d_arr_20__9), .D (nx1160), .CLK (nx10171)) ;
    inv01 ix1161 (.Y (nx1160), .A (nx7447)) ;
    aoi222 ix7448 (.Y (nx7447), .A0 (d_arr_mux_20__9), .A1 (nx11265), .B0 (
           d_arr_mul_20__9), .B1 (nx10403), .C0 (d_arr_add_20__9), .C1 (nx10631)
           ) ;
    latch lat_d_arr_20__10 (.Q (d_arr_20__10), .D (nx1172), .CLK (nx10171)) ;
    inv01 ix1173 (.Y (nx1172), .A (nx7453)) ;
    aoi222 ix7454 (.Y (nx7453), .A0 (d_arr_mux_20__10), .A1 (nx11265), .B0 (
           d_arr_mul_20__10), .B1 (nx10403), .C0 (d_arr_add_20__10), .C1 (
           nx10633)) ;
    latch lat_d_arr_20__11 (.Q (d_arr_20__11), .D (nx1184), .CLK (nx10171)) ;
    inv01 ix1185 (.Y (nx1184), .A (nx7459)) ;
    aoi222 ix7460 (.Y (nx7459), .A0 (d_arr_mux_20__11), .A1 (nx11265), .B0 (
           d_arr_mul_20__11), .B1 (nx10403), .C0 (d_arr_add_20__11), .C1 (
           nx10633)) ;
    latch lat_d_arr_20__12 (.Q (d_arr_20__12), .D (nx1196), .CLK (nx10173)) ;
    inv01 ix1197 (.Y (nx1196), .A (nx7463)) ;
    aoi222 ix7464 (.Y (nx7463), .A0 (d_arr_mux_20__12), .A1 (nx11265), .B0 (
           d_arr_mul_20__12), .B1 (nx10405), .C0 (d_arr_add_20__12), .C1 (
           nx10633)) ;
    latch lat_d_arr_20__13 (.Q (d_arr_20__13), .D (nx1208), .CLK (nx10173)) ;
    inv01 ix1209 (.Y (nx1208), .A (nx7469)) ;
    aoi222 ix7470 (.Y (nx7469), .A0 (d_arr_mux_20__13), .A1 (nx11265), .B0 (
           d_arr_mul_20__13), .B1 (nx10405), .C0 (d_arr_add_20__13), .C1 (
           nx10633)) ;
    latch lat_d_arr_20__14 (.Q (d_arr_20__14), .D (nx1220), .CLK (nx10173)) ;
    inv01 ix1221 (.Y (nx1220), .A (nx7475)) ;
    aoi222 ix7476 (.Y (nx7475), .A0 (d_arr_mux_20__14), .A1 (nx11267), .B0 (
           d_arr_mul_20__14), .B1 (nx10405), .C0 (d_arr_add_20__14), .C1 (
           nx10633)) ;
    latch lat_d_arr_20__15 (.Q (d_arr_20__15), .D (nx1232), .CLK (nx10173)) ;
    nand02 ix1233 (.Y (nx1232), .A0 (nx7481), .A1 (nx10849)) ;
    aoi22 ix7482 (.Y (nx7481), .A0 (d_arr_mul_20__15), .A1 (nx10405), .B0 (
          d_arr_add_20__15), .B1 (nx10633)) ;
    nand02 ix7484 (.Y (nx7483), .A0 (d_arr_mux_20__31), .A1 (nx11267)) ;
    latch lat_d_arr_20__16 (.Q (d_arr_20__16), .D (nx1242), .CLK (nx10173)) ;
    nand02 ix1243 (.Y (nx1242), .A0 (nx7489), .A1 (nx10849)) ;
    aoi22 ix7490 (.Y (nx7489), .A0 (d_arr_mul_20__16), .A1 (nx10405), .B0 (
          d_arr_add_20__16), .B1 (nx10633)) ;
    latch lat_d_arr_20__17 (.Q (d_arr_20__17), .D (nx1252), .CLK (nx10173)) ;
    nand02 ix1253 (.Y (nx1252), .A0 (nx7495), .A1 (nx10849)) ;
    aoi22 ix7496 (.Y (nx7495), .A0 (d_arr_mul_20__17), .A1 (nx10405), .B0 (
          d_arr_add_20__17), .B1 (nx10635)) ;
    latch lat_d_arr_20__18 (.Q (d_arr_20__18), .D (nx1262), .CLK (nx10173)) ;
    nand02 ix1263 (.Y (nx1262), .A0 (nx7501), .A1 (nx10849)) ;
    aoi22 ix7502 (.Y (nx7501), .A0 (d_arr_mul_20__18), .A1 (nx10405), .B0 (
          d_arr_add_20__18), .B1 (nx10635)) ;
    latch lat_d_arr_20__19 (.Q (d_arr_20__19), .D (nx1272), .CLK (nx10175)) ;
    nand02 ix1273 (.Y (nx1272), .A0 (nx7507), .A1 (nx10849)) ;
    aoi22 ix7508 (.Y (nx7507), .A0 (d_arr_mul_20__19), .A1 (nx10407), .B0 (
          d_arr_add_20__19), .B1 (nx10635)) ;
    latch lat_d_arr_20__20 (.Q (d_arr_20__20), .D (nx1282), .CLK (nx10175)) ;
    nand02 ix1283 (.Y (nx1282), .A0 (nx7513), .A1 (nx10849)) ;
    aoi22 ix7514 (.Y (nx7513), .A0 (d_arr_mul_20__20), .A1 (nx10407), .B0 (
          d_arr_add_20__20), .B1 (nx10635)) ;
    latch lat_d_arr_20__21 (.Q (d_arr_20__21), .D (nx1292), .CLK (nx10175)) ;
    nand02 ix1293 (.Y (nx1292), .A0 (nx7519), .A1 (nx10849)) ;
    aoi22 ix7520 (.Y (nx7519), .A0 (d_arr_mul_20__21), .A1 (nx10407), .B0 (
          d_arr_add_20__21), .B1 (nx10635)) ;
    latch lat_d_arr_20__22 (.Q (d_arr_20__22), .D (nx1302), .CLK (nx10175)) ;
    nand02 ix1303 (.Y (nx1302), .A0 (nx7525), .A1 (nx10851)) ;
    aoi22 ix7526 (.Y (nx7525), .A0 (d_arr_mul_20__22), .A1 (nx10407), .B0 (
          d_arr_add_20__22), .B1 (nx10635)) ;
    latch lat_d_arr_20__23 (.Q (d_arr_20__23), .D (nx1312), .CLK (nx10175)) ;
    nand02 ix1313 (.Y (nx1312), .A0 (nx7529), .A1 (nx10851)) ;
    aoi22 ix7530 (.Y (nx7529), .A0 (d_arr_mul_20__23), .A1 (nx10407), .B0 (
          d_arr_add_20__23), .B1 (nx10635)) ;
    latch lat_d_arr_20__24 (.Q (d_arr_20__24), .D (nx1322), .CLK (nx10175)) ;
    nand02 ix1323 (.Y (nx1322), .A0 (nx7535), .A1 (nx10851)) ;
    aoi22 ix7536 (.Y (nx7535), .A0 (d_arr_mul_20__24), .A1 (nx10407), .B0 (
          d_arr_add_20__24), .B1 (nx10637)) ;
    latch lat_d_arr_20__25 (.Q (d_arr_20__25), .D (nx1332), .CLK (nx10175)) ;
    nand02 ix1333 (.Y (nx1332), .A0 (nx7541), .A1 (nx10851)) ;
    aoi22 ix7542 (.Y (nx7541), .A0 (d_arr_mul_20__25), .A1 (nx10407), .B0 (
          d_arr_add_20__25), .B1 (nx10637)) ;
    latch lat_d_arr_20__26 (.Q (d_arr_20__26), .D (nx1342), .CLK (nx10177)) ;
    nand02 ix1343 (.Y (nx1342), .A0 (nx7547), .A1 (nx10851)) ;
    aoi22 ix7548 (.Y (nx7547), .A0 (d_arr_mul_20__26), .A1 (nx10409), .B0 (
          d_arr_add_20__26), .B1 (nx10637)) ;
    latch lat_d_arr_20__27 (.Q (d_arr_20__27), .D (nx1352), .CLK (nx10177)) ;
    nand02 ix1353 (.Y (nx1352), .A0 (nx7551), .A1 (nx10851)) ;
    aoi22 ix7552 (.Y (nx7551), .A0 (d_arr_mul_20__27), .A1 (nx10409), .B0 (
          d_arr_add_20__27), .B1 (nx10637)) ;
    latch lat_d_arr_20__28 (.Q (d_arr_20__28), .D (nx1362), .CLK (nx10177)) ;
    nand02 ix1363 (.Y (nx1362), .A0 (nx7557), .A1 (nx10851)) ;
    aoi22 ix7558 (.Y (nx7557), .A0 (d_arr_mul_20__28), .A1 (nx10409), .B0 (
          d_arr_add_20__28), .B1 (nx10637)) ;
    latch lat_d_arr_20__29 (.Q (d_arr_20__29), .D (nx1372), .CLK (nx10177)) ;
    nand02 ix1373 (.Y (nx1372), .A0 (nx7563), .A1 (nx7483)) ;
    aoi22 ix7564 (.Y (nx7563), .A0 (d_arr_mul_20__29), .A1 (nx10409), .B0 (
          d_arr_add_20__29), .B1 (nx10637)) ;
    latch lat_d_arr_20__30 (.Q (d_arr_20__30), .D (nx1382), .CLK (nx10177)) ;
    nand02 ix1383 (.Y (nx1382), .A0 (nx7569), .A1 (nx7483)) ;
    aoi22 ix7570 (.Y (nx7569), .A0 (d_arr_mul_20__30), .A1 (nx10409), .B0 (
          d_arr_add_20__30), .B1 (nx10637)) ;
    latch lat_d_arr_20__31 (.Q (d_arr_20__31), .D (nx1392), .CLK (nx10177)) ;
    nand02 ix1393 (.Y (nx1392), .A0 (nx7573), .A1 (nx7483)) ;
    aoi22 ix7574 (.Y (nx7573), .A0 (d_arr_mul_20__31), .A1 (nx10409), .B0 (
          d_arr_add_20__31), .B1 (nx10639)) ;
    latch lat_d_arr_19__0 (.Q (d_arr_19__0), .D (nx1404), .CLK (nx10177)) ;
    inv01 ix1405 (.Y (nx1404), .A (nx7579)) ;
    aoi222 ix7580 (.Y (nx7579), .A0 (d_arr_mux_19__0), .A1 (nx11267), .B0 (
           d_arr_mul_19__0), .B1 (nx10409), .C0 (d_arr_add_19__0), .C1 (nx10639)
           ) ;
    latch lat_d_arr_19__1 (.Q (d_arr_19__1), .D (nx1416), .CLK (nx10179)) ;
    inv01 ix1417 (.Y (nx1416), .A (nx7585)) ;
    aoi222 ix7586 (.Y (nx7585), .A0 (d_arr_mux_19__1), .A1 (nx11267), .B0 (
           d_arr_mul_19__1), .B1 (nx10411), .C0 (d_arr_add_19__1), .C1 (nx10639)
           ) ;
    latch lat_d_arr_19__2 (.Q (d_arr_19__2), .D (nx1428), .CLK (nx10179)) ;
    inv01 ix1429 (.Y (nx1428), .A (nx7591)) ;
    aoi222 ix7592 (.Y (nx7591), .A0 (d_arr_mux_19__2), .A1 (nx11267), .B0 (
           d_arr_mul_19__2), .B1 (nx10411), .C0 (d_arr_add_19__2), .C1 (nx10639)
           ) ;
    latch lat_d_arr_19__3 (.Q (d_arr_19__3), .D (nx1440), .CLK (nx10179)) ;
    inv01 ix1441 (.Y (nx1440), .A (nx7595)) ;
    aoi222 ix7596 (.Y (nx7595), .A0 (d_arr_mux_19__3), .A1 (nx11267), .B0 (
           d_arr_mul_19__3), .B1 (nx10411), .C0 (d_arr_add_19__3), .C1 (nx10639)
           ) ;
    latch lat_d_arr_19__4 (.Q (d_arr_19__4), .D (nx1452), .CLK (nx10179)) ;
    inv01 ix1453 (.Y (nx1452), .A (nx7601)) ;
    aoi222 ix7602 (.Y (nx7601), .A0 (d_arr_mux_19__4), .A1 (nx11267), .B0 (
           d_arr_mul_19__4), .B1 (nx10411), .C0 (d_arr_add_19__4), .C1 (nx10639)
           ) ;
    latch lat_d_arr_19__5 (.Q (d_arr_19__5), .D (nx1464), .CLK (nx10179)) ;
    inv01 ix1465 (.Y (nx1464), .A (nx7607)) ;
    aoi222 ix7608 (.Y (nx7607), .A0 (d_arr_mux_19__5), .A1 (nx11269), .B0 (
           d_arr_mul_19__5), .B1 (nx10411), .C0 (d_arr_add_19__5), .C1 (nx10639)
           ) ;
    latch lat_d_arr_19__6 (.Q (d_arr_19__6), .D (nx1476), .CLK (nx10179)) ;
    inv01 ix1477 (.Y (nx1476), .A (nx7613)) ;
    aoi222 ix7614 (.Y (nx7613), .A0 (d_arr_mux_19__6), .A1 (nx11269), .B0 (
           d_arr_mul_19__6), .B1 (nx10411), .C0 (d_arr_add_19__6), .C1 (nx10641)
           ) ;
    latch lat_d_arr_19__7 (.Q (d_arr_19__7), .D (nx1488), .CLK (nx10179)) ;
    inv01 ix1489 (.Y (nx1488), .A (nx7617)) ;
    aoi222 ix7618 (.Y (nx7617), .A0 (d_arr_mux_19__7), .A1 (nx11269), .B0 (
           d_arr_mul_19__7), .B1 (nx10411), .C0 (d_arr_add_19__7), .C1 (nx10641)
           ) ;
    latch lat_d_arr_19__8 (.Q (d_arr_19__8), .D (nx1500), .CLK (nx10181)) ;
    inv01 ix1501 (.Y (nx1500), .A (nx7623)) ;
    aoi222 ix7624 (.Y (nx7623), .A0 (d_arr_mux_19__8), .A1 (nx11269), .B0 (
           d_arr_mul_19__8), .B1 (nx10413), .C0 (d_arr_add_19__8), .C1 (nx10641)
           ) ;
    latch lat_d_arr_19__9 (.Q (d_arr_19__9), .D (nx1512), .CLK (nx10181)) ;
    inv01 ix1513 (.Y (nx1512), .A (nx7629)) ;
    aoi222 ix7630 (.Y (nx7629), .A0 (d_arr_mux_19__9), .A1 (nx11269), .B0 (
           d_arr_mul_19__9), .B1 (nx10413), .C0 (d_arr_add_19__9), .C1 (nx10641)
           ) ;
    latch lat_d_arr_19__10 (.Q (d_arr_19__10), .D (nx1524), .CLK (nx10181)) ;
    inv01 ix1525 (.Y (nx1524), .A (nx7635)) ;
    aoi222 ix7636 (.Y (nx7635), .A0 (d_arr_mux_19__10), .A1 (nx11269), .B0 (
           d_arr_mul_19__10), .B1 (nx10413), .C0 (d_arr_add_19__10), .C1 (
           nx10641)) ;
    latch lat_d_arr_19__11 (.Q (d_arr_19__11), .D (nx1536), .CLK (nx10181)) ;
    inv01 ix1537 (.Y (nx1536), .A (nx7639)) ;
    aoi222 ix7640 (.Y (nx7639), .A0 (d_arr_mux_19__11), .A1 (nx11269), .B0 (
           d_arr_mul_19__11), .B1 (nx10413), .C0 (d_arr_add_19__11), .C1 (
           nx10641)) ;
    latch lat_d_arr_19__12 (.Q (d_arr_19__12), .D (nx1548), .CLK (nx10181)) ;
    inv01 ix1549 (.Y (nx1548), .A (nx7645)) ;
    aoi222 ix7646 (.Y (nx7645), .A0 (d_arr_mux_19__12), .A1 (nx11271), .B0 (
           d_arr_mul_19__12), .B1 (nx10413), .C0 (d_arr_add_19__12), .C1 (
           nx10641)) ;
    latch lat_d_arr_19__13 (.Q (d_arr_19__13), .D (nx1560), .CLK (nx10181)) ;
    inv01 ix1561 (.Y (nx1560), .A (nx7651)) ;
    aoi222 ix7652 (.Y (nx7651), .A0 (d_arr_mux_19__13), .A1 (nx11271), .B0 (
           d_arr_mul_19__13), .B1 (nx10413), .C0 (d_arr_add_19__13), .C1 (
           nx10643)) ;
    latch lat_d_arr_19__14 (.Q (d_arr_19__14), .D (nx1572), .CLK (nx10181)) ;
    inv01 ix1573 (.Y (nx1572), .A (nx7657)) ;
    aoi222 ix7658 (.Y (nx7657), .A0 (d_arr_mux_19__14), .A1 (nx11271), .B0 (
           d_arr_mul_19__14), .B1 (nx10413), .C0 (d_arr_add_19__14), .C1 (
           nx10643)) ;
    latch lat_d_arr_19__15 (.Q (d_arr_19__15), .D (nx1584), .CLK (nx10183)) ;
    nand02 ix1585 (.Y (nx1584), .A0 (nx7661), .A1 (nx10853)) ;
    aoi22 ix7662 (.Y (nx7661), .A0 (d_arr_mul_19__15), .A1 (nx10415), .B0 (
          d_arr_add_19__15), .B1 (nx10643)) ;
    nand02 ix7664 (.Y (nx7663), .A0 (d_arr_mux_19__31), .A1 (nx11271)) ;
    latch lat_d_arr_19__16 (.Q (d_arr_19__16), .D (nx1594), .CLK (nx10183)) ;
    nand02 ix1595 (.Y (nx1594), .A0 (nx7669), .A1 (nx10853)) ;
    aoi22 ix7670 (.Y (nx7669), .A0 (d_arr_mul_19__16), .A1 (nx10415), .B0 (
          d_arr_add_19__16), .B1 (nx10643)) ;
    latch lat_d_arr_19__17 (.Q (d_arr_19__17), .D (nx1604), .CLK (nx10183)) ;
    nand02 ix1605 (.Y (nx1604), .A0 (nx7675), .A1 (nx10853)) ;
    aoi22 ix7676 (.Y (nx7675), .A0 (d_arr_mul_19__17), .A1 (nx10415), .B0 (
          d_arr_add_19__17), .B1 (nx10643)) ;
    latch lat_d_arr_19__18 (.Q (d_arr_19__18), .D (nx1614), .CLK (nx10183)) ;
    nand02 ix1615 (.Y (nx1614), .A0 (nx7681), .A1 (nx10853)) ;
    aoi22 ix7682 (.Y (nx7681), .A0 (d_arr_mul_19__18), .A1 (nx10415), .B0 (
          d_arr_add_19__18), .B1 (nx10643)) ;
    latch lat_d_arr_19__19 (.Q (d_arr_19__19), .D (nx1624), .CLK (nx10183)) ;
    nand02 ix1625 (.Y (nx1624), .A0 (nx7687), .A1 (nx10853)) ;
    aoi22 ix7688 (.Y (nx7687), .A0 (d_arr_mul_19__19), .A1 (nx10415), .B0 (
          d_arr_add_19__19), .B1 (nx10643)) ;
    latch lat_d_arr_19__20 (.Q (d_arr_19__20), .D (nx1634), .CLK (nx10183)) ;
    nand02 ix1635 (.Y (nx1634), .A0 (nx7693), .A1 (nx10853)) ;
    aoi22 ix7694 (.Y (nx7693), .A0 (d_arr_mul_19__20), .A1 (nx10415), .B0 (
          d_arr_add_19__20), .B1 (nx10645)) ;
    latch lat_d_arr_19__21 (.Q (d_arr_19__21), .D (nx1644), .CLK (nx10183)) ;
    nand02 ix1645 (.Y (nx1644), .A0 (nx7699), .A1 (nx10853)) ;
    aoi22 ix7700 (.Y (nx7699), .A0 (d_arr_mul_19__21), .A1 (nx10415), .B0 (
          d_arr_add_19__21), .B1 (nx10645)) ;
    latch lat_d_arr_19__22 (.Q (d_arr_19__22), .D (nx1654), .CLK (nx10185)) ;
    nand02 ix1655 (.Y (nx1654), .A0 (nx7705), .A1 (nx10855)) ;
    aoi22 ix7706 (.Y (nx7705), .A0 (d_arr_mul_19__22), .A1 (nx10417), .B0 (
          d_arr_add_19__22), .B1 (nx10645)) ;
    latch lat_d_arr_19__23 (.Q (d_arr_19__23), .D (nx1664), .CLK (nx10185)) ;
    nand02 ix1665 (.Y (nx1664), .A0 (nx7711), .A1 (nx10855)) ;
    aoi22 ix7712 (.Y (nx7711), .A0 (d_arr_mul_19__23), .A1 (nx10417), .B0 (
          d_arr_add_19__23), .B1 (nx10645)) ;
    latch lat_d_arr_19__24 (.Q (d_arr_19__24), .D (nx1674), .CLK (nx10185)) ;
    nand02 ix1675 (.Y (nx1674), .A0 (nx7717), .A1 (nx10855)) ;
    aoi22 ix7718 (.Y (nx7717), .A0 (d_arr_mul_19__24), .A1 (nx10417), .B0 (
          d_arr_add_19__24), .B1 (nx10645)) ;
    latch lat_d_arr_19__25 (.Q (d_arr_19__25), .D (nx1684), .CLK (nx10185)) ;
    nand02 ix1685 (.Y (nx1684), .A0 (nx7723), .A1 (nx10855)) ;
    aoi22 ix7724 (.Y (nx7723), .A0 (d_arr_mul_19__25), .A1 (nx10417), .B0 (
          d_arr_add_19__25), .B1 (nx10645)) ;
    latch lat_d_arr_19__26 (.Q (d_arr_19__26), .D (nx1694), .CLK (nx10185)) ;
    nand02 ix1695 (.Y (nx1694), .A0 (nx7727), .A1 (nx10855)) ;
    aoi22 ix7728 (.Y (nx7727), .A0 (d_arr_mul_19__26), .A1 (nx10417), .B0 (
          d_arr_add_19__26), .B1 (nx10645)) ;
    latch lat_d_arr_19__27 (.Q (d_arr_19__27), .D (nx1704), .CLK (nx10185)) ;
    nand02 ix1705 (.Y (nx1704), .A0 (nx7733), .A1 (nx10855)) ;
    aoi22 ix7734 (.Y (nx7733), .A0 (d_arr_mul_19__27), .A1 (nx10417), .B0 (
          d_arr_add_19__27), .B1 (nx10647)) ;
    latch lat_d_arr_19__28 (.Q (d_arr_19__28), .D (nx1714), .CLK (nx10185)) ;
    nand02 ix1715 (.Y (nx1714), .A0 (nx7739), .A1 (nx10855)) ;
    aoi22 ix7740 (.Y (nx7739), .A0 (d_arr_mul_19__28), .A1 (nx10417), .B0 (
          d_arr_add_19__28), .B1 (nx10647)) ;
    latch lat_d_arr_19__29 (.Q (d_arr_19__29), .D (nx1724), .CLK (nx10187)) ;
    nand02 ix1725 (.Y (nx1724), .A0 (nx7745), .A1 (nx7663)) ;
    aoi22 ix7746 (.Y (nx7745), .A0 (d_arr_mul_19__29), .A1 (nx10419), .B0 (
          d_arr_add_19__29), .B1 (nx10647)) ;
    latch lat_d_arr_19__30 (.Q (d_arr_19__30), .D (nx1734), .CLK (nx10187)) ;
    nand02 ix1735 (.Y (nx1734), .A0 (nx7749), .A1 (nx7663)) ;
    aoi22 ix7750 (.Y (nx7749), .A0 (d_arr_mul_19__30), .A1 (nx10419), .B0 (
          d_arr_add_19__30), .B1 (nx10647)) ;
    latch lat_d_arr_19__31 (.Q (d_arr_19__31), .D (nx1744), .CLK (nx10187)) ;
    nand02 ix1745 (.Y (nx1744), .A0 (nx7755), .A1 (nx7663)) ;
    aoi22 ix7756 (.Y (nx7755), .A0 (d_arr_mul_19__31), .A1 (nx10419), .B0 (
          d_arr_add_19__31), .B1 (nx10647)) ;
    latch lat_d_arr_18__0 (.Q (d_arr_18__0), .D (nx1756), .CLK (nx10187)) ;
    inv01 ix1757 (.Y (nx1756), .A (nx7761)) ;
    aoi222 ix7762 (.Y (nx7761), .A0 (d_arr_mux_18__0), .A1 (nx11271), .B0 (
           d_arr_mul_18__0), .B1 (nx10419), .C0 (d_arr_add_18__0), .C1 (nx10647)
           ) ;
    latch lat_d_arr_18__1 (.Q (d_arr_18__1), .D (nx1768), .CLK (nx10187)) ;
    inv01 ix1769 (.Y (nx1768), .A (nx7767)) ;
    aoi222 ix7768 (.Y (nx7767), .A0 (d_arr_mux_18__1), .A1 (nx11271), .B0 (
           d_arr_mul_18__1), .B1 (nx10419), .C0 (d_arr_add_18__1), .C1 (nx10647)
           ) ;
    latch lat_d_arr_18__2 (.Q (d_arr_18__2), .D (nx1780), .CLK (nx10187)) ;
    inv01 ix1781 (.Y (nx1780), .A (nx7773)) ;
    aoi222 ix7774 (.Y (nx7773), .A0 (d_arr_mux_18__2), .A1 (nx11271), .B0 (
           d_arr_mul_18__2), .B1 (nx10419), .C0 (d_arr_add_18__2), .C1 (nx10649)
           ) ;
    latch lat_d_arr_18__3 (.Q (d_arr_18__3), .D (nx1792), .CLK (nx10187)) ;
    inv01 ix1793 (.Y (nx1792), .A (nx7779)) ;
    aoi222 ix7780 (.Y (nx7779), .A0 (d_arr_mux_18__3), .A1 (nx11273), .B0 (
           d_arr_mul_18__3), .B1 (nx10419), .C0 (d_arr_add_18__3), .C1 (nx10649)
           ) ;
    latch lat_d_arr_18__4 (.Q (d_arr_18__4), .D (nx1804), .CLK (nx10189)) ;
    inv01 ix1805 (.Y (nx1804), .A (nx7785)) ;
    aoi222 ix7786 (.Y (nx7785), .A0 (d_arr_mux_18__4), .A1 (nx11273), .B0 (
           d_arr_mul_18__4), .B1 (nx10421), .C0 (d_arr_add_18__4), .C1 (nx10649)
           ) ;
    latch lat_d_arr_18__5 (.Q (d_arr_18__5), .D (nx1816), .CLK (nx10189)) ;
    inv01 ix1817 (.Y (nx1816), .A (nx7791)) ;
    aoi222 ix7792 (.Y (nx7791), .A0 (d_arr_mux_18__5), .A1 (nx11273), .B0 (
           d_arr_mul_18__5), .B1 (nx10421), .C0 (d_arr_add_18__5), .C1 (nx10649)
           ) ;
    latch lat_d_arr_18__6 (.Q (d_arr_18__6), .D (nx1828), .CLK (nx10189)) ;
    inv01 ix1829 (.Y (nx1828), .A (nx7797)) ;
    aoi222 ix7798 (.Y (nx7797), .A0 (d_arr_mux_18__6), .A1 (nx11273), .B0 (
           d_arr_mul_18__6), .B1 (nx10421), .C0 (d_arr_add_18__6), .C1 (nx10649)
           ) ;
    latch lat_d_arr_18__7 (.Q (d_arr_18__7), .D (nx1840), .CLK (nx10189)) ;
    inv01 ix1841 (.Y (nx1840), .A (nx7803)) ;
    aoi222 ix7804 (.Y (nx7803), .A0 (d_arr_mux_18__7), .A1 (nx11273), .B0 (
           d_arr_mul_18__7), .B1 (nx10421), .C0 (d_arr_add_18__7), .C1 (nx10649)
           ) ;
    latch lat_d_arr_18__8 (.Q (d_arr_18__8), .D (nx1852), .CLK (nx10189)) ;
    inv01 ix1853 (.Y (nx1852), .A (nx7809)) ;
    aoi222 ix7810 (.Y (nx7809), .A0 (d_arr_mux_18__8), .A1 (nx11273), .B0 (
           d_arr_mul_18__8), .B1 (nx10421), .C0 (d_arr_add_18__8), .C1 (nx10649)
           ) ;
    latch lat_d_arr_18__9 (.Q (d_arr_18__9), .D (nx1864), .CLK (nx10189)) ;
    inv01 ix1865 (.Y (nx1864), .A (nx7815)) ;
    aoi222 ix7816 (.Y (nx7815), .A0 (d_arr_mux_18__9), .A1 (nx11273), .B0 (
           d_arr_mul_18__9), .B1 (nx10421), .C0 (d_arr_add_18__9), .C1 (nx10651)
           ) ;
    latch lat_d_arr_18__10 (.Q (d_arr_18__10), .D (nx1876), .CLK (nx10189)) ;
    inv01 ix1877 (.Y (nx1876), .A (nx7821)) ;
    aoi222 ix7822 (.Y (nx7821), .A0 (d_arr_mux_18__10), .A1 (nx11275), .B0 (
           d_arr_mul_18__10), .B1 (nx10421), .C0 (d_arr_add_18__10), .C1 (
           nx10651)) ;
    latch lat_d_arr_18__11 (.Q (d_arr_18__11), .D (nx1888), .CLK (nx10191)) ;
    inv01 ix1889 (.Y (nx1888), .A (nx7827)) ;
    aoi222 ix7828 (.Y (nx7827), .A0 (d_arr_mux_18__11), .A1 (nx11275), .B0 (
           d_arr_mul_18__11), .B1 (nx10423), .C0 (d_arr_add_18__11), .C1 (
           nx10651)) ;
    latch lat_d_arr_18__12 (.Q (d_arr_18__12), .D (nx1900), .CLK (nx10191)) ;
    inv01 ix1901 (.Y (nx1900), .A (nx7833)) ;
    aoi222 ix7834 (.Y (nx7833), .A0 (d_arr_mux_18__12), .A1 (nx11275), .B0 (
           d_arr_mul_18__12), .B1 (nx10423), .C0 (d_arr_add_18__12), .C1 (
           nx10651)) ;
    latch lat_d_arr_18__13 (.Q (d_arr_18__13), .D (nx1912), .CLK (nx10191)) ;
    inv01 ix1913 (.Y (nx1912), .A (nx7839)) ;
    aoi222 ix7840 (.Y (nx7839), .A0 (d_arr_mux_18__13), .A1 (nx11275), .B0 (
           d_arr_mul_18__13), .B1 (nx10423), .C0 (d_arr_add_18__13), .C1 (
           nx10651)) ;
    latch lat_d_arr_18__14 (.Q (d_arr_18__14), .D (nx1924), .CLK (nx10191)) ;
    inv01 ix1925 (.Y (nx1924), .A (nx7845)) ;
    aoi222 ix7846 (.Y (nx7845), .A0 (d_arr_mux_18__14), .A1 (nx11275), .B0 (
           d_arr_mul_18__14), .B1 (nx10423), .C0 (d_arr_add_18__14), .C1 (
           nx10651)) ;
    latch lat_d_arr_18__15 (.Q (d_arr_18__15), .D (nx1936), .CLK (nx10191)) ;
    nand02 ix1937 (.Y (nx1936), .A0 (nx7851), .A1 (nx10857)) ;
    aoi22 ix7852 (.Y (nx7851), .A0 (d_arr_mul_18__15), .A1 (nx10423), .B0 (
          d_arr_add_18__15), .B1 (nx10651)) ;
    nand02 ix7854 (.Y (nx7853), .A0 (d_arr_mux_18__31), .A1 (nx11275)) ;
    latch lat_d_arr_18__16 (.Q (d_arr_18__16), .D (nx1946), .CLK (nx10191)) ;
    nand02 ix1947 (.Y (nx1946), .A0 (nx7859), .A1 (nx10857)) ;
    aoi22 ix7860 (.Y (nx7859), .A0 (d_arr_mul_18__16), .A1 (nx10423), .B0 (
          d_arr_add_18__16), .B1 (nx10653)) ;
    latch lat_d_arr_18__17 (.Q (d_arr_18__17), .D (nx1956), .CLK (nx10191)) ;
    nand02 ix1957 (.Y (nx1956), .A0 (nx7865), .A1 (nx10857)) ;
    aoi22 ix7866 (.Y (nx7865), .A0 (d_arr_mul_18__17), .A1 (nx10423), .B0 (
          d_arr_add_18__17), .B1 (nx10653)) ;
    latch lat_d_arr_18__18 (.Q (d_arr_18__18), .D (nx1966), .CLK (nx10193)) ;
    nand02 ix1967 (.Y (nx1966), .A0 (nx7869), .A1 (nx10857)) ;
    aoi22 ix7870 (.Y (nx7869), .A0 (d_arr_mul_18__18), .A1 (nx10425), .B0 (
          d_arr_add_18__18), .B1 (nx10653)) ;
    latch lat_d_arr_18__19 (.Q (d_arr_18__19), .D (nx1976), .CLK (nx10193)) ;
    nand02 ix1977 (.Y (nx1976), .A0 (nx7875), .A1 (nx10857)) ;
    aoi22 ix7876 (.Y (nx7875), .A0 (d_arr_mul_18__19), .A1 (nx10425), .B0 (
          d_arr_add_18__19), .B1 (nx10653)) ;
    latch lat_d_arr_18__20 (.Q (d_arr_18__20), .D (nx1986), .CLK (nx10193)) ;
    nand02 ix1987 (.Y (nx1986), .A0 (nx7881), .A1 (nx10857)) ;
    aoi22 ix7882 (.Y (nx7881), .A0 (d_arr_mul_18__20), .A1 (nx10425), .B0 (
          d_arr_add_18__20), .B1 (nx10653)) ;
    latch lat_d_arr_18__21 (.Q (d_arr_18__21), .D (nx1996), .CLK (nx10193)) ;
    nand02 ix1997 (.Y (nx1996), .A0 (nx7887), .A1 (nx10857)) ;
    aoi22 ix7888 (.Y (nx7887), .A0 (d_arr_mul_18__21), .A1 (nx10425), .B0 (
          d_arr_add_18__21), .B1 (nx10653)) ;
    latch lat_d_arr_18__22 (.Q (d_arr_18__22), .D (nx2006), .CLK (nx10193)) ;
    nand02 ix2007 (.Y (nx2006), .A0 (nx7893), .A1 (nx10859)) ;
    aoi22 ix7894 (.Y (nx7893), .A0 (d_arr_mul_18__22), .A1 (nx10425), .B0 (
          d_arr_add_18__22), .B1 (nx10653)) ;
    latch lat_d_arr_18__23 (.Q (d_arr_18__23), .D (nx2016), .CLK (nx10193)) ;
    nand02 ix2017 (.Y (nx2016), .A0 (nx7899), .A1 (nx10859)) ;
    aoi22 ix7900 (.Y (nx7899), .A0 (d_arr_mul_18__23), .A1 (nx10425), .B0 (
          d_arr_add_18__23), .B1 (nx10655)) ;
    latch lat_d_arr_18__24 (.Q (d_arr_18__24), .D (nx2026), .CLK (nx10193)) ;
    nand02 ix2027 (.Y (nx2026), .A0 (nx7905), .A1 (nx10859)) ;
    aoi22 ix7906 (.Y (nx7905), .A0 (d_arr_mul_18__24), .A1 (nx10425), .B0 (
          d_arr_add_18__24), .B1 (nx10655)) ;
    latch lat_d_arr_18__25 (.Q (d_arr_18__25), .D (nx2036), .CLK (nx10195)) ;
    nand02 ix2037 (.Y (nx2036), .A0 (nx7911), .A1 (nx10859)) ;
    aoi22 ix7912 (.Y (nx7911), .A0 (d_arr_mul_18__25), .A1 (nx10427), .B0 (
          d_arr_add_18__25), .B1 (nx10655)) ;
    latch lat_d_arr_18__26 (.Q (d_arr_18__26), .D (nx2046), .CLK (nx10195)) ;
    nand02 ix2047 (.Y (nx2046), .A0 (nx7917), .A1 (nx10859)) ;
    aoi22 ix7918 (.Y (nx7917), .A0 (d_arr_mul_18__26), .A1 (nx10427), .B0 (
          d_arr_add_18__26), .B1 (nx10655)) ;
    latch lat_d_arr_18__27 (.Q (d_arr_18__27), .D (nx2056), .CLK (nx10195)) ;
    nand02 ix2057 (.Y (nx2056), .A0 (nx7923), .A1 (nx10859)) ;
    aoi22 ix7924 (.Y (nx7923), .A0 (d_arr_mul_18__27), .A1 (nx10427), .B0 (
          d_arr_add_18__27), .B1 (nx10655)) ;
    latch lat_d_arr_18__28 (.Q (d_arr_18__28), .D (nx2066), .CLK (nx10195)) ;
    nand02 ix2067 (.Y (nx2066), .A0 (nx7929), .A1 (nx10859)) ;
    aoi22 ix7930 (.Y (nx7929), .A0 (d_arr_mul_18__28), .A1 (nx10427), .B0 (
          d_arr_add_18__28), .B1 (nx10655)) ;
    latch lat_d_arr_18__29 (.Q (d_arr_18__29), .D (nx2076), .CLK (nx10195)) ;
    nand02 ix2077 (.Y (nx2076), .A0 (nx7935), .A1 (nx7853)) ;
    aoi22 ix7936 (.Y (nx7935), .A0 (d_arr_mul_18__29), .A1 (nx10427), .B0 (
          d_arr_add_18__29), .B1 (nx10655)) ;
    latch lat_d_arr_18__30 (.Q (d_arr_18__30), .D (nx2086), .CLK (nx10195)) ;
    nand02 ix2087 (.Y (nx2086), .A0 (nx7941), .A1 (nx7853)) ;
    aoi22 ix7942 (.Y (nx7941), .A0 (d_arr_mul_18__30), .A1 (nx10427), .B0 (
          d_arr_add_18__30), .B1 (nx10657)) ;
    latch lat_d_arr_18__31 (.Q (d_arr_18__31), .D (nx2096), .CLK (nx10195)) ;
    nand02 ix2097 (.Y (nx2096), .A0 (nx7947), .A1 (nx7853)) ;
    aoi22 ix7948 (.Y (nx7947), .A0 (d_arr_mul_18__31), .A1 (nx10427), .B0 (
          d_arr_add_18__31), .B1 (nx10657)) ;
    latch lat_d_arr_17__0 (.Q (d_arr_17__0), .D (nx2104), .CLK (nx10197)) ;
    ao22 ix2105 (.Y (nx2104), .A0 (d_arr_mux_17__0), .A1 (nx11275), .B0 (
         d_arr_mul_17__0), .B1 (nx10429)) ;
    latch lat_d_arr_17__1 (.Q (d_arr_17__1), .D (nx2112), .CLK (nx10197)) ;
    ao22 ix2113 (.Y (nx2112), .A0 (d_arr_mux_17__1), .A1 (nx11277), .B0 (
         d_arr_mul_17__1), .B1 (nx10429)) ;
    latch lat_d_arr_17__2 (.Q (d_arr_17__2), .D (nx2120), .CLK (nx10197)) ;
    ao22 ix2121 (.Y (nx2120), .A0 (d_arr_mux_17__2), .A1 (nx11277), .B0 (
         d_arr_mul_17__2), .B1 (nx10429)) ;
    latch lat_d_arr_17__3 (.Q (d_arr_17__3), .D (nx2128), .CLK (nx10197)) ;
    ao22 ix2129 (.Y (nx2128), .A0 (d_arr_mux_17__3), .A1 (nx11277), .B0 (
         d_arr_mul_17__3), .B1 (nx10429)) ;
    latch lat_d_arr_17__4 (.Q (d_arr_17__4), .D (nx2136), .CLK (nx10197)) ;
    ao22 ix2137 (.Y (nx2136), .A0 (d_arr_mux_17__4), .A1 (nx11277), .B0 (
         d_arr_mul_17__4), .B1 (nx10429)) ;
    latch lat_d_arr_17__5 (.Q (d_arr_17__5), .D (nx2144), .CLK (nx10197)) ;
    ao22 ix2145 (.Y (nx2144), .A0 (d_arr_mux_17__5), .A1 (nx11277), .B0 (
         d_arr_mul_17__5), .B1 (nx10429)) ;
    latch lat_d_arr_17__6 (.Q (d_arr_17__6), .D (nx2152), .CLK (nx10197)) ;
    ao22 ix2153 (.Y (nx2152), .A0 (d_arr_mux_17__6), .A1 (nx11277), .B0 (
         d_arr_mul_17__6), .B1 (nx10429)) ;
    latch lat_d_arr_17__7 (.Q (d_arr_17__7), .D (nx2160), .CLK (nx10199)) ;
    ao22 ix2161 (.Y (nx2160), .A0 (d_arr_mux_17__7), .A1 (nx11277), .B0 (
         d_arr_mul_17__7), .B1 (nx10431)) ;
    latch lat_d_arr_17__8 (.Q (d_arr_17__8), .D (nx2168), .CLK (nx10199)) ;
    ao22 ix2169 (.Y (nx2168), .A0 (d_arr_mux_17__8), .A1 (nx11279), .B0 (
         d_arr_mul_17__8), .B1 (nx10431)) ;
    latch lat_d_arr_17__9 (.Q (d_arr_17__9), .D (nx2176), .CLK (nx10199)) ;
    ao22 ix2177 (.Y (nx2176), .A0 (d_arr_mux_17__9), .A1 (nx11279), .B0 (
         d_arr_mul_17__9), .B1 (nx10431)) ;
    latch lat_d_arr_17__10 (.Q (d_arr_17__10), .D (nx2184), .CLK (nx10199)) ;
    ao22 ix2185 (.Y (nx2184), .A0 (d_arr_mux_17__10), .A1 (nx11279), .B0 (
         d_arr_mul_17__10), .B1 (nx10431)) ;
    latch lat_d_arr_17__11 (.Q (d_arr_17__11), .D (nx2192), .CLK (nx10199)) ;
    ao22 ix2193 (.Y (nx2192), .A0 (d_arr_mux_17__11), .A1 (nx11279), .B0 (
         d_arr_mul_17__11), .B1 (nx10431)) ;
    latch lat_d_arr_17__12 (.Q (d_arr_17__12), .D (nx2200), .CLK (nx10199)) ;
    ao22 ix2201 (.Y (nx2200), .A0 (d_arr_mux_17__12), .A1 (nx11279), .B0 (
         d_arr_mul_17__12), .B1 (nx10431)) ;
    latch lat_d_arr_17__13 (.Q (d_arr_17__13), .D (nx2208), .CLK (nx10199)) ;
    ao22 ix2209 (.Y (nx2208), .A0 (d_arr_mux_17__13), .A1 (nx11279), .B0 (
         d_arr_mul_17__13), .B1 (nx10431)) ;
    latch lat_d_arr_17__14 (.Q (d_arr_17__14), .D (nx2216), .CLK (nx10201)) ;
    ao22 ix2217 (.Y (nx2216), .A0 (d_arr_mux_17__14), .A1 (nx11279), .B0 (
         d_arr_mul_17__14), .B1 (nx10433)) ;
    latch lat_d_arr_17__15 (.Q (d_arr_17__15), .D (nx2224), .CLK (nx10201)) ;
    ao22 ix2225 (.Y (nx2224), .A0 (d_arr_mux_17__15), .A1 (nx11281), .B0 (
         d_arr_mul_17__15), .B1 (nx10433)) ;
    latch lat_d_arr_17__16 (.Q (d_arr_17__16), .D (nx2232), .CLK (nx10201)) ;
    ao22 ix2233 (.Y (nx2232), .A0 (d_arr_mux_17__16), .A1 (nx11281), .B0 (
         d_arr_mul_17__16), .B1 (nx10433)) ;
    latch lat_d_arr_17__17 (.Q (d_arr_17__17), .D (nx2240), .CLK (nx10201)) ;
    ao22 ix2241 (.Y (nx2240), .A0 (d_arr_mux_17__17), .A1 (nx11281), .B0 (
         d_arr_mul_17__17), .B1 (nx10433)) ;
    latch lat_d_arr_17__18 (.Q (d_arr_17__18), .D (nx2248), .CLK (nx10201)) ;
    ao22 ix2249 (.Y (nx2248), .A0 (d_arr_mux_17__18), .A1 (nx11281), .B0 (
         d_arr_mul_17__18), .B1 (nx10433)) ;
    latch lat_d_arr_17__19 (.Q (d_arr_17__19), .D (nx2256), .CLK (nx10201)) ;
    ao22 ix2257 (.Y (nx2256), .A0 (d_arr_mux_17__19), .A1 (nx11281), .B0 (
         d_arr_mul_17__19), .B1 (nx10433)) ;
    latch lat_d_arr_17__20 (.Q (d_arr_17__20), .D (nx2264), .CLK (nx10201)) ;
    ao22 ix2265 (.Y (nx2264), .A0 (d_arr_mux_17__20), .A1 (nx11281), .B0 (
         d_arr_mul_17__20), .B1 (nx10433)) ;
    latch lat_d_arr_17__21 (.Q (d_arr_17__21), .D (nx2272), .CLK (nx10203)) ;
    ao22 ix2273 (.Y (nx2272), .A0 (d_arr_mux_17__21), .A1 (nx11281), .B0 (
         d_arr_mul_17__21), .B1 (nx10435)) ;
    latch lat_d_arr_17__22 (.Q (d_arr_17__22), .D (nx2280), .CLK (nx10203)) ;
    ao22 ix2281 (.Y (nx2280), .A0 (d_arr_mux_17__22), .A1 (nx11283), .B0 (
         d_arr_mul_17__22), .B1 (nx10435)) ;
    latch lat_d_arr_17__23 (.Q (d_arr_17__23), .D (nx2288), .CLK (nx10203)) ;
    ao22 ix2289 (.Y (nx2288), .A0 (d_arr_mux_17__23), .A1 (nx11283), .B0 (
         d_arr_mul_17__23), .B1 (nx10435)) ;
    latch lat_d_arr_17__24 (.Q (d_arr_17__24), .D (nx2296), .CLK (nx10203)) ;
    ao22 ix2297 (.Y (nx2296), .A0 (d_arr_mux_17__24), .A1 (nx11283), .B0 (
         d_arr_mul_17__24), .B1 (nx10435)) ;
    latch lat_d_arr_17__25 (.Q (d_arr_17__25), .D (nx2304), .CLK (nx10203)) ;
    ao22 ix2305 (.Y (nx2304), .A0 (d_arr_mux_17__25), .A1 (nx11283), .B0 (
         d_arr_mul_17__25), .B1 (nx10435)) ;
    latch lat_d_arr_17__26 (.Q (d_arr_17__26), .D (nx2312), .CLK (nx10203)) ;
    ao22 ix2313 (.Y (nx2312), .A0 (d_arr_mux_17__26), .A1 (nx11283), .B0 (
         d_arr_mul_17__26), .B1 (nx10435)) ;
    latch lat_d_arr_17__27 (.Q (d_arr_17__27), .D (nx2320), .CLK (nx10203)) ;
    ao22 ix2321 (.Y (nx2320), .A0 (d_arr_mux_17__27), .A1 (nx11283), .B0 (
         d_arr_mul_17__27), .B1 (nx10435)) ;
    latch lat_d_arr_17__28 (.Q (d_arr_17__28), .D (nx2328), .CLK (nx10205)) ;
    ao22 ix2329 (.Y (nx2328), .A0 (d_arr_mux_17__28), .A1 (nx11283), .B0 (
         d_arr_mul_17__28), .B1 (nx10437)) ;
    latch lat_d_arr_17__29 (.Q (d_arr_17__29), .D (nx2336), .CLK (nx10205)) ;
    ao22 ix2337 (.Y (nx2336), .A0 (d_arr_mux_17__29), .A1 (nx11285), .B0 (
         d_arr_mul_17__29), .B1 (nx10437)) ;
    latch lat_d_arr_17__30 (.Q (d_arr_17__30), .D (nx2344), .CLK (nx10205)) ;
    ao22 ix2345 (.Y (nx2344), .A0 (d_arr_mux_17__30), .A1 (nx11285), .B0 (
         d_arr_mul_17__30), .B1 (nx10437)) ;
    latch lat_d_arr_17__31 (.Q (d_arr_17__31), .D (nx2352), .CLK (nx10205)) ;
    ao22 ix2353 (.Y (nx2352), .A0 (d_arr_mux_17__31), .A1 (nx11285), .B0 (
         d_arr_mul_17__31), .B1 (nx10437)) ;
    latch lat_d_arr_16__0 (.Q (d_arr_16__0), .D (nx2360), .CLK (nx10205)) ;
    ao22 ix2361 (.Y (nx2360), .A0 (d_arr_mux_16__0), .A1 (nx11285), .B0 (
         d_arr_mul_16__0), .B1 (nx10437)) ;
    latch lat_d_arr_16__1 (.Q (d_arr_16__1), .D (nx2368), .CLK (nx10205)) ;
    ao22 ix2369 (.Y (nx2368), .A0 (d_arr_mux_16__1), .A1 (nx11285), .B0 (
         d_arr_mul_16__1), .B1 (nx10437)) ;
    latch lat_d_arr_16__2 (.Q (d_arr_16__2), .D (nx2376), .CLK (nx10205)) ;
    ao22 ix2377 (.Y (nx2376), .A0 (d_arr_mux_16__2), .A1 (nx11285), .B0 (
         d_arr_mul_16__2), .B1 (nx10437)) ;
    latch lat_d_arr_16__3 (.Q (d_arr_16__3), .D (nx2384), .CLK (nx10207)) ;
    ao22 ix2385 (.Y (nx2384), .A0 (d_arr_mux_16__3), .A1 (nx11285), .B0 (
         d_arr_mul_16__3), .B1 (nx10439)) ;
    latch lat_d_arr_16__4 (.Q (d_arr_16__4), .D (nx2392), .CLK (nx10207)) ;
    ao22 ix2393 (.Y (nx2392), .A0 (d_arr_mux_16__4), .A1 (nx11287), .B0 (
         d_arr_mul_16__4), .B1 (nx10439)) ;
    latch lat_d_arr_16__5 (.Q (d_arr_16__5), .D (nx2400), .CLK (nx10207)) ;
    ao22 ix2401 (.Y (nx2400), .A0 (d_arr_mux_16__5), .A1 (nx11287), .B0 (
         d_arr_mul_16__5), .B1 (nx10439)) ;
    latch lat_d_arr_16__6 (.Q (d_arr_16__6), .D (nx2408), .CLK (nx10207)) ;
    ao22 ix2409 (.Y (nx2408), .A0 (d_arr_mux_16__6), .A1 (nx11287), .B0 (
         d_arr_mul_16__6), .B1 (nx10439)) ;
    latch lat_d_arr_16__7 (.Q (d_arr_16__7), .D (nx2416), .CLK (nx10207)) ;
    ao22 ix2417 (.Y (nx2416), .A0 (d_arr_mux_16__7), .A1 (nx11287), .B0 (
         d_arr_mul_16__7), .B1 (nx10439)) ;
    latch lat_d_arr_16__8 (.Q (d_arr_16__8), .D (nx2424), .CLK (nx10207)) ;
    ao22 ix2425 (.Y (nx2424), .A0 (d_arr_mux_16__8), .A1 (nx11287), .B0 (
         d_arr_mul_16__8), .B1 (nx10439)) ;
    latch lat_d_arr_16__9 (.Q (d_arr_16__9), .D (nx2432), .CLK (nx10207)) ;
    ao22 ix2433 (.Y (nx2432), .A0 (d_arr_mux_16__9), .A1 (nx11287), .B0 (
         d_arr_mul_16__9), .B1 (nx10439)) ;
    latch lat_d_arr_16__10 (.Q (d_arr_16__10), .D (nx2440), .CLK (nx10209)) ;
    ao22 ix2441 (.Y (nx2440), .A0 (d_arr_mux_16__10), .A1 (nx11287), .B0 (
         d_arr_mul_16__10), .B1 (nx10441)) ;
    latch lat_d_arr_16__11 (.Q (d_arr_16__11), .D (nx2448), .CLK (nx10209)) ;
    ao22 ix2449 (.Y (nx2448), .A0 (d_arr_mux_16__11), .A1 (nx11289), .B0 (
         d_arr_mul_16__11), .B1 (nx10441)) ;
    latch lat_d_arr_16__12 (.Q (d_arr_16__12), .D (nx2456), .CLK (nx10209)) ;
    ao22 ix2457 (.Y (nx2456), .A0 (d_arr_mux_16__12), .A1 (nx11289), .B0 (
         d_arr_mul_16__12), .B1 (nx10441)) ;
    latch lat_d_arr_16__13 (.Q (d_arr_16__13), .D (nx2464), .CLK (nx10209)) ;
    ao22 ix2465 (.Y (nx2464), .A0 (d_arr_mux_16__13), .A1 (nx11289), .B0 (
         d_arr_mul_16__13), .B1 (nx10441)) ;
    latch lat_d_arr_16__14 (.Q (d_arr_16__14), .D (nx2472), .CLK (nx10209)) ;
    ao22 ix2473 (.Y (nx2472), .A0 (d_arr_mux_16__14), .A1 (nx11289), .B0 (
         d_arr_mul_16__14), .B1 (nx10441)) ;
    latch lat_d_arr_16__15 (.Q (d_arr_16__15), .D (nx2480), .CLK (nx10209)) ;
    ao22 ix2481 (.Y (nx2480), .A0 (d_arr_mux_16__15), .A1 (nx11289), .B0 (
         d_arr_mul_16__15), .B1 (nx10441)) ;
    latch lat_d_arr_16__16 (.Q (d_arr_16__16), .D (nx2488), .CLK (nx10209)) ;
    ao22 ix2489 (.Y (nx2488), .A0 (d_arr_mux_16__16), .A1 (nx11289), .B0 (
         d_arr_mul_16__16), .B1 (nx10441)) ;
    latch lat_d_arr_16__17 (.Q (d_arr_16__17), .D (nx2496), .CLK (nx10211)) ;
    ao22 ix2497 (.Y (nx2496), .A0 (d_arr_mux_16__17), .A1 (nx11289), .B0 (
         d_arr_mul_16__17), .B1 (nx10443)) ;
    latch lat_d_arr_16__18 (.Q (d_arr_16__18), .D (nx2504), .CLK (nx10211)) ;
    ao22 ix2505 (.Y (nx2504), .A0 (d_arr_mux_16__18), .A1 (nx11291), .B0 (
         d_arr_mul_16__18), .B1 (nx10443)) ;
    latch lat_d_arr_16__19 (.Q (d_arr_16__19), .D (nx2512), .CLK (nx10211)) ;
    ao22 ix2513 (.Y (nx2512), .A0 (d_arr_mux_16__19), .A1 (nx11291), .B0 (
         d_arr_mul_16__19), .B1 (nx10443)) ;
    latch lat_d_arr_16__20 (.Q (d_arr_16__20), .D (nx2520), .CLK (nx10211)) ;
    ao22 ix2521 (.Y (nx2520), .A0 (d_arr_mux_16__20), .A1 (nx11291), .B0 (
         d_arr_mul_16__20), .B1 (nx10443)) ;
    latch lat_d_arr_16__21 (.Q (d_arr_16__21), .D (nx2528), .CLK (nx10211)) ;
    ao22 ix2529 (.Y (nx2528), .A0 (d_arr_mux_16__21), .A1 (nx11291), .B0 (
         d_arr_mul_16__21), .B1 (nx10443)) ;
    latch lat_d_arr_16__22 (.Q (d_arr_16__22), .D (nx2536), .CLK (nx10211)) ;
    ao22 ix2537 (.Y (nx2536), .A0 (d_arr_mux_16__22), .A1 (nx11291), .B0 (
         d_arr_mul_16__22), .B1 (nx10443)) ;
    latch lat_d_arr_16__23 (.Q (d_arr_16__23), .D (nx2544), .CLK (nx10211)) ;
    ao22 ix2545 (.Y (nx2544), .A0 (d_arr_mux_16__23), .A1 (nx11291), .B0 (
         d_arr_mul_16__23), .B1 (nx10443)) ;
    latch lat_d_arr_16__24 (.Q (d_arr_16__24), .D (nx2552), .CLK (nx10213)) ;
    ao22 ix2553 (.Y (nx2552), .A0 (d_arr_mux_16__24), .A1 (nx11291), .B0 (
         d_arr_mul_16__24), .B1 (nx10445)) ;
    latch lat_d_arr_16__25 (.Q (d_arr_16__25), .D (nx2560), .CLK (nx10213)) ;
    ao22 ix2561 (.Y (nx2560), .A0 (d_arr_mux_16__25), .A1 (nx11293), .B0 (
         d_arr_mul_16__25), .B1 (nx10445)) ;
    latch lat_d_arr_16__26 (.Q (d_arr_16__26), .D (nx2568), .CLK (nx10213)) ;
    ao22 ix2569 (.Y (nx2568), .A0 (d_arr_mux_16__26), .A1 (nx11293), .B0 (
         d_arr_mul_16__26), .B1 (nx10445)) ;
    latch lat_d_arr_16__27 (.Q (d_arr_16__27), .D (nx2576), .CLK (nx10213)) ;
    ao22 ix2577 (.Y (nx2576), .A0 (d_arr_mux_16__27), .A1 (nx11293), .B0 (
         d_arr_mul_16__27), .B1 (nx10445)) ;
    latch lat_d_arr_16__28 (.Q (d_arr_16__28), .D (nx2584), .CLK (nx10213)) ;
    ao22 ix2585 (.Y (nx2584), .A0 (d_arr_mux_16__28), .A1 (nx11293), .B0 (
         d_arr_mul_16__28), .B1 (nx10445)) ;
    latch lat_d_arr_16__29 (.Q (d_arr_16__29), .D (nx2592), .CLK (nx10213)) ;
    ao22 ix2593 (.Y (nx2592), .A0 (d_arr_mux_16__29), .A1 (nx11293), .B0 (
         d_arr_mul_16__29), .B1 (nx10445)) ;
    latch lat_d_arr_16__30 (.Q (d_arr_16__30), .D (nx2600), .CLK (nx10213)) ;
    ao22 ix2601 (.Y (nx2600), .A0 (d_arr_mux_16__30), .A1 (nx11293), .B0 (
         d_arr_mul_16__30), .B1 (nx10445)) ;
    latch lat_d_arr_16__31 (.Q (d_arr_16__31), .D (nx2608), .CLK (nx10215)) ;
    ao22 ix2609 (.Y (nx2608), .A0 (d_arr_mux_16__31), .A1 (nx11293), .B0 (
         d_arr_mul_16__31), .B1 (nx10447)) ;
    latch lat_d_arr_15__0 (.Q (d_arr_15__0), .D (nx2616), .CLK (nx10215)) ;
    ao22 ix2617 (.Y (nx2616), .A0 (d_arr_mux_15__0), .A1 (nx11295), .B0 (
         d_arr_mul_15__0), .B1 (nx10447)) ;
    latch lat_d_arr_15__1 (.Q (d_arr_15__1), .D (nx2624), .CLK (nx10215)) ;
    ao22 ix2625 (.Y (nx2624), .A0 (d_arr_mux_15__1), .A1 (nx11295), .B0 (
         d_arr_mul_15__1), .B1 (nx10447)) ;
    latch lat_d_arr_15__2 (.Q (d_arr_15__2), .D (nx2632), .CLK (nx10215)) ;
    ao22 ix2633 (.Y (nx2632), .A0 (d_arr_mux_15__2), .A1 (nx11295), .B0 (
         d_arr_mul_15__2), .B1 (nx10447)) ;
    latch lat_d_arr_15__3 (.Q (d_arr_15__3), .D (nx2640), .CLK (nx10215)) ;
    ao22 ix2641 (.Y (nx2640), .A0 (d_arr_mux_15__3), .A1 (nx11295), .B0 (
         d_arr_mul_15__3), .B1 (nx10447)) ;
    latch lat_d_arr_15__4 (.Q (d_arr_15__4), .D (nx2648), .CLK (nx10215)) ;
    ao22 ix2649 (.Y (nx2648), .A0 (d_arr_mux_15__4), .A1 (nx11295), .B0 (
         d_arr_mul_15__4), .B1 (nx10447)) ;
    latch lat_d_arr_15__5 (.Q (d_arr_15__5), .D (nx2656), .CLK (nx10215)) ;
    ao22 ix2657 (.Y (nx2656), .A0 (d_arr_mux_15__5), .A1 (nx11295), .B0 (
         d_arr_mul_15__5), .B1 (nx10447)) ;
    latch lat_d_arr_15__6 (.Q (d_arr_15__6), .D (nx2664), .CLK (nx10217)) ;
    ao22 ix2665 (.Y (nx2664), .A0 (d_arr_mux_15__6), .A1 (nx11295), .B0 (
         d_arr_mul_15__6), .B1 (nx10449)) ;
    latch lat_d_arr_15__7 (.Q (d_arr_15__7), .D (nx2672), .CLK (nx10217)) ;
    ao22 ix2673 (.Y (nx2672), .A0 (d_arr_mux_15__7), .A1 (nx11297), .B0 (
         d_arr_mul_15__7), .B1 (nx10449)) ;
    latch lat_d_arr_15__8 (.Q (d_arr_15__8), .D (nx2680), .CLK (nx10217)) ;
    ao22 ix2681 (.Y (nx2680), .A0 (d_arr_mux_15__8), .A1 (nx11297), .B0 (
         d_arr_mul_15__8), .B1 (nx10449)) ;
    latch lat_d_arr_15__9 (.Q (d_arr_15__9), .D (nx2688), .CLK (nx10217)) ;
    ao22 ix2689 (.Y (nx2688), .A0 (d_arr_mux_15__9), .A1 (nx11297), .B0 (
         d_arr_mul_15__9), .B1 (nx10449)) ;
    latch lat_d_arr_15__10 (.Q (d_arr_15__10), .D (nx2696), .CLK (nx10217)) ;
    ao22 ix2697 (.Y (nx2696), .A0 (d_arr_mux_15__10), .A1 (nx11297), .B0 (
         d_arr_mul_15__10), .B1 (nx10449)) ;
    latch lat_d_arr_15__11 (.Q (d_arr_15__11), .D (nx2704), .CLK (nx10217)) ;
    ao22 ix2705 (.Y (nx2704), .A0 (d_arr_mux_15__11), .A1 (nx11297), .B0 (
         d_arr_mul_15__11), .B1 (nx10449)) ;
    latch lat_d_arr_15__12 (.Q (d_arr_15__12), .D (nx2712), .CLK (nx10217)) ;
    ao22 ix2713 (.Y (nx2712), .A0 (d_arr_mux_15__12), .A1 (nx11297), .B0 (
         d_arr_mul_15__12), .B1 (nx10449)) ;
    latch lat_d_arr_15__13 (.Q (d_arr_15__13), .D (nx2720), .CLK (nx10219)) ;
    ao22 ix2721 (.Y (nx2720), .A0 (d_arr_mux_15__13), .A1 (nx11297), .B0 (
         d_arr_mul_15__13), .B1 (nx10451)) ;
    latch lat_d_arr_15__14 (.Q (d_arr_15__14), .D (nx2728), .CLK (nx10219)) ;
    ao22 ix2729 (.Y (nx2728), .A0 (d_arr_mux_15__14), .A1 (nx11299), .B0 (
         d_arr_mul_15__14), .B1 (nx10451)) ;
    latch lat_d_arr_15__15 (.Q (d_arr_15__15), .D (nx2736), .CLK (nx10219)) ;
    ao22 ix2737 (.Y (nx2736), .A0 (d_arr_mux_15__15), .A1 (nx11299), .B0 (
         d_arr_mul_15__15), .B1 (nx10451)) ;
    latch lat_d_arr_15__16 (.Q (d_arr_15__16), .D (nx2744), .CLK (nx10219)) ;
    ao22 ix2745 (.Y (nx2744), .A0 (d_arr_mux_15__16), .A1 (nx11299), .B0 (
         d_arr_mul_15__16), .B1 (nx10451)) ;
    latch lat_d_arr_15__17 (.Q (d_arr_15__17), .D (nx2752), .CLK (nx10219)) ;
    ao22 ix2753 (.Y (nx2752), .A0 (d_arr_mux_15__17), .A1 (nx11299), .B0 (
         d_arr_mul_15__17), .B1 (nx10451)) ;
    latch lat_d_arr_15__18 (.Q (d_arr_15__18), .D (nx2760), .CLK (nx10219)) ;
    ao22 ix2761 (.Y (nx2760), .A0 (d_arr_mux_15__18), .A1 (nx11299), .B0 (
         d_arr_mul_15__18), .B1 (nx10451)) ;
    latch lat_d_arr_15__19 (.Q (d_arr_15__19), .D (nx2768), .CLK (nx10219)) ;
    ao22 ix2769 (.Y (nx2768), .A0 (d_arr_mux_15__19), .A1 (nx11299), .B0 (
         d_arr_mul_15__19), .B1 (nx10451)) ;
    latch lat_d_arr_15__20 (.Q (d_arr_15__20), .D (nx2776), .CLK (nx10221)) ;
    ao22 ix2777 (.Y (nx2776), .A0 (d_arr_mux_15__20), .A1 (nx11299), .B0 (
         d_arr_mul_15__20), .B1 (nx10453)) ;
    latch lat_d_arr_15__21 (.Q (d_arr_15__21), .D (nx2784), .CLK (nx10221)) ;
    ao22 ix2785 (.Y (nx2784), .A0 (d_arr_mux_15__21), .A1 (nx11301), .B0 (
         d_arr_mul_15__21), .B1 (nx10453)) ;
    latch lat_d_arr_15__22 (.Q (d_arr_15__22), .D (nx2792), .CLK (nx10221)) ;
    ao22 ix2793 (.Y (nx2792), .A0 (d_arr_mux_15__22), .A1 (nx11301), .B0 (
         d_arr_mul_15__22), .B1 (nx10453)) ;
    latch lat_d_arr_15__23 (.Q (d_arr_15__23), .D (nx2800), .CLK (nx10221)) ;
    ao22 ix2801 (.Y (nx2800), .A0 (d_arr_mux_15__23), .A1 (nx11301), .B0 (
         d_arr_mul_15__23), .B1 (nx10453)) ;
    latch lat_d_arr_15__24 (.Q (d_arr_15__24), .D (nx2808), .CLK (nx10221)) ;
    ao22 ix2809 (.Y (nx2808), .A0 (d_arr_mux_15__24), .A1 (nx11301), .B0 (
         d_arr_mul_15__24), .B1 (nx10453)) ;
    latch lat_d_arr_15__25 (.Q (d_arr_15__25), .D (nx2816), .CLK (nx10221)) ;
    ao22 ix2817 (.Y (nx2816), .A0 (d_arr_mux_15__25), .A1 (nx11301), .B0 (
         d_arr_mul_15__25), .B1 (nx10453)) ;
    latch lat_d_arr_15__26 (.Q (d_arr_15__26), .D (nx2824), .CLK (nx10221)) ;
    ao22 ix2825 (.Y (nx2824), .A0 (d_arr_mux_15__26), .A1 (nx11301), .B0 (
         d_arr_mul_15__26), .B1 (nx10453)) ;
    latch lat_d_arr_15__27 (.Q (d_arr_15__27), .D (nx2832), .CLK (nx10223)) ;
    ao22 ix2833 (.Y (nx2832), .A0 (d_arr_mux_15__27), .A1 (nx11301), .B0 (
         d_arr_mul_15__27), .B1 (nx10455)) ;
    latch lat_d_arr_15__28 (.Q (d_arr_15__28), .D (nx2840), .CLK (nx10223)) ;
    ao22 ix2841 (.Y (nx2840), .A0 (d_arr_mux_15__28), .A1 (nx11303), .B0 (
         d_arr_mul_15__28), .B1 (nx10455)) ;
    latch lat_d_arr_15__29 (.Q (d_arr_15__29), .D (nx2848), .CLK (nx10223)) ;
    ao22 ix2849 (.Y (nx2848), .A0 (d_arr_mux_15__29), .A1 (nx11303), .B0 (
         d_arr_mul_15__29), .B1 (nx10455)) ;
    latch lat_d_arr_15__30 (.Q (d_arr_15__30), .D (nx2856), .CLK (nx10223)) ;
    ao22 ix2857 (.Y (nx2856), .A0 (d_arr_mux_15__30), .A1 (nx11303), .B0 (
         d_arr_mul_15__30), .B1 (nx10455)) ;
    latch lat_d_arr_15__31 (.Q (d_arr_15__31), .D (nx2864), .CLK (nx10223)) ;
    ao22 ix2865 (.Y (nx2864), .A0 (d_arr_mux_15__31), .A1 (nx11303), .B0 (
         d_arr_mul_15__31), .B1 (nx10455)) ;
    latch lat_d_arr_14__0 (.Q (d_arr_14__0), .D (nx2872), .CLK (nx10223)) ;
    ao22 ix2873 (.Y (nx2872), .A0 (d_arr_mux_14__0), .A1 (nx11303), .B0 (
         d_arr_mul_14__0), .B1 (nx10455)) ;
    latch lat_d_arr_14__1 (.Q (d_arr_14__1), .D (nx2880), .CLK (nx10223)) ;
    ao22 ix2881 (.Y (nx2880), .A0 (d_arr_mux_14__1), .A1 (nx11303), .B0 (
         d_arr_mul_14__1), .B1 (nx10455)) ;
    latch lat_d_arr_14__2 (.Q (d_arr_14__2), .D (nx2888), .CLK (nx10225)) ;
    ao22 ix2889 (.Y (nx2888), .A0 (d_arr_mux_14__2), .A1 (nx11303), .B0 (
         d_arr_mul_14__2), .B1 (nx10457)) ;
    latch lat_d_arr_14__3 (.Q (d_arr_14__3), .D (nx2896), .CLK (nx10225)) ;
    ao22 ix2897 (.Y (nx2896), .A0 (d_arr_mux_14__3), .A1 (nx11305), .B0 (
         d_arr_mul_14__3), .B1 (nx10457)) ;
    latch lat_d_arr_14__4 (.Q (d_arr_14__4), .D (nx2904), .CLK (nx10225)) ;
    ao22 ix2905 (.Y (nx2904), .A0 (d_arr_mux_14__4), .A1 (nx11305), .B0 (
         d_arr_mul_14__4), .B1 (nx10457)) ;
    latch lat_d_arr_14__5 (.Q (d_arr_14__5), .D (nx2912), .CLK (nx10225)) ;
    ao22 ix2913 (.Y (nx2912), .A0 (d_arr_mux_14__5), .A1 (nx11305), .B0 (
         d_arr_mul_14__5), .B1 (nx10457)) ;
    latch lat_d_arr_14__6 (.Q (d_arr_14__6), .D (nx2920), .CLK (nx10225)) ;
    ao22 ix2921 (.Y (nx2920), .A0 (d_arr_mux_14__6), .A1 (nx11305), .B0 (
         d_arr_mul_14__6), .B1 (nx10457)) ;
    latch lat_d_arr_14__7 (.Q (d_arr_14__7), .D (nx2928), .CLK (nx10225)) ;
    ao22 ix2929 (.Y (nx2928), .A0 (d_arr_mux_14__7), .A1 (nx11305), .B0 (
         d_arr_mul_14__7), .B1 (nx10457)) ;
    latch lat_d_arr_14__8 (.Q (d_arr_14__8), .D (nx2936), .CLK (nx10225)) ;
    ao22 ix2937 (.Y (nx2936), .A0 (d_arr_mux_14__8), .A1 (nx11305), .B0 (
         d_arr_mul_14__8), .B1 (nx10457)) ;
    latch lat_d_arr_14__9 (.Q (d_arr_14__9), .D (nx2944), .CLK (nx10227)) ;
    ao22 ix2945 (.Y (nx2944), .A0 (d_arr_mux_14__9), .A1 (nx11305), .B0 (
         d_arr_mul_14__9), .B1 (nx10459)) ;
    latch lat_d_arr_14__10 (.Q (d_arr_14__10), .D (nx2952), .CLK (nx10227)) ;
    ao22 ix2953 (.Y (nx2952), .A0 (d_arr_mux_14__10), .A1 (nx11307), .B0 (
         d_arr_mul_14__10), .B1 (nx10459)) ;
    latch lat_d_arr_14__11 (.Q (d_arr_14__11), .D (nx2960), .CLK (nx10227)) ;
    ao22 ix2961 (.Y (nx2960), .A0 (d_arr_mux_14__11), .A1 (nx11307), .B0 (
         d_arr_mul_14__11), .B1 (nx10459)) ;
    latch lat_d_arr_14__12 (.Q (d_arr_14__12), .D (nx2968), .CLK (nx10227)) ;
    ao22 ix2969 (.Y (nx2968), .A0 (d_arr_mux_14__12), .A1 (nx11307), .B0 (
         d_arr_mul_14__12), .B1 (nx10459)) ;
    latch lat_d_arr_14__13 (.Q (d_arr_14__13), .D (nx2976), .CLK (nx10227)) ;
    ao22 ix2977 (.Y (nx2976), .A0 (d_arr_mux_14__13), .A1 (nx11307), .B0 (
         d_arr_mul_14__13), .B1 (nx10459)) ;
    latch lat_d_arr_14__14 (.Q (d_arr_14__14), .D (nx2984), .CLK (nx10227)) ;
    ao22 ix2985 (.Y (nx2984), .A0 (d_arr_mux_14__14), .A1 (nx11307), .B0 (
         d_arr_mul_14__14), .B1 (nx10459)) ;
    latch lat_d_arr_14__15 (.Q (d_arr_14__15), .D (nx2992), .CLK (nx10227)) ;
    ao22 ix2993 (.Y (nx2992), .A0 (d_arr_mux_14__15), .A1 (nx11307), .B0 (
         d_arr_mul_14__15), .B1 (nx10459)) ;
    latch lat_d_arr_14__16 (.Q (d_arr_14__16), .D (nx3000), .CLK (nx10229)) ;
    ao22 ix3001 (.Y (nx3000), .A0 (d_arr_mux_14__16), .A1 (nx11307), .B0 (
         d_arr_mul_14__16), .B1 (nx10461)) ;
    latch lat_d_arr_14__17 (.Q (d_arr_14__17), .D (nx3008), .CLK (nx10229)) ;
    ao22 ix3009 (.Y (nx3008), .A0 (d_arr_mux_14__17), .A1 (nx11309), .B0 (
         d_arr_mul_14__17), .B1 (nx10461)) ;
    latch lat_d_arr_14__18 (.Q (d_arr_14__18), .D (nx3016), .CLK (nx10229)) ;
    ao22 ix3017 (.Y (nx3016), .A0 (d_arr_mux_14__18), .A1 (nx11309), .B0 (
         d_arr_mul_14__18), .B1 (nx10461)) ;
    latch lat_d_arr_14__19 (.Q (d_arr_14__19), .D (nx3024), .CLK (nx10229)) ;
    ao22 ix3025 (.Y (nx3024), .A0 (d_arr_mux_14__19), .A1 (nx11309), .B0 (
         d_arr_mul_14__19), .B1 (nx10461)) ;
    latch lat_d_arr_14__20 (.Q (d_arr_14__20), .D (nx3032), .CLK (nx10229)) ;
    ao22 ix3033 (.Y (nx3032), .A0 (d_arr_mux_14__20), .A1 (nx11309), .B0 (
         d_arr_mul_14__20), .B1 (nx10461)) ;
    latch lat_d_arr_14__21 (.Q (d_arr_14__21), .D (nx3040), .CLK (nx10229)) ;
    ao22 ix3041 (.Y (nx3040), .A0 (d_arr_mux_14__21), .A1 (nx11309), .B0 (
         d_arr_mul_14__21), .B1 (nx10461)) ;
    latch lat_d_arr_14__22 (.Q (d_arr_14__22), .D (nx3048), .CLK (nx10229)) ;
    ao22 ix3049 (.Y (nx3048), .A0 (d_arr_mux_14__22), .A1 (nx11309), .B0 (
         d_arr_mul_14__22), .B1 (nx10461)) ;
    latch lat_d_arr_14__23 (.Q (d_arr_14__23), .D (nx3056), .CLK (nx10231)) ;
    ao22 ix3057 (.Y (nx3056), .A0 (d_arr_mux_14__23), .A1 (nx11309), .B0 (
         d_arr_mul_14__23), .B1 (nx10463)) ;
    latch lat_d_arr_14__24 (.Q (d_arr_14__24), .D (nx3064), .CLK (nx10231)) ;
    ao22 ix3065 (.Y (nx3064), .A0 (d_arr_mux_14__24), .A1 (nx11311), .B0 (
         d_arr_mul_14__24), .B1 (nx10463)) ;
    latch lat_d_arr_14__25 (.Q (d_arr_14__25), .D (nx3072), .CLK (nx10231)) ;
    ao22 ix3073 (.Y (nx3072), .A0 (d_arr_mux_14__25), .A1 (nx11311), .B0 (
         d_arr_mul_14__25), .B1 (nx10463)) ;
    latch lat_d_arr_14__26 (.Q (d_arr_14__26), .D (nx3080), .CLK (nx10231)) ;
    ao22 ix3081 (.Y (nx3080), .A0 (d_arr_mux_14__26), .A1 (nx11311), .B0 (
         d_arr_mul_14__26), .B1 (nx10463)) ;
    latch lat_d_arr_14__27 (.Q (d_arr_14__27), .D (nx3088), .CLK (nx10231)) ;
    ao22 ix3089 (.Y (nx3088), .A0 (d_arr_mux_14__27), .A1 (nx11311), .B0 (
         d_arr_mul_14__27), .B1 (nx10463)) ;
    latch lat_d_arr_14__28 (.Q (d_arr_14__28), .D (nx3096), .CLK (nx10231)) ;
    ao22 ix3097 (.Y (nx3096), .A0 (d_arr_mux_14__28), .A1 (nx11311), .B0 (
         d_arr_mul_14__28), .B1 (nx10463)) ;
    latch lat_d_arr_14__29 (.Q (d_arr_14__29), .D (nx3104), .CLK (nx10231)) ;
    ao22 ix3105 (.Y (nx3104), .A0 (d_arr_mux_14__29), .A1 (nx11311), .B0 (
         d_arr_mul_14__29), .B1 (nx10463)) ;
    latch lat_d_arr_14__30 (.Q (d_arr_14__30), .D (nx3112), .CLK (nx10233)) ;
    ao22 ix3113 (.Y (nx3112), .A0 (d_arr_mux_14__30), .A1 (nx11311), .B0 (
         d_arr_mul_14__30), .B1 (nx10465)) ;
    latch lat_d_arr_14__31 (.Q (d_arr_14__31), .D (nx3120), .CLK (nx10233)) ;
    ao22 ix3121 (.Y (nx3120), .A0 (d_arr_mux_14__31), .A1 (nx11313), .B0 (
         d_arr_mul_14__31), .B1 (nx10465)) ;
    latch lat_d_arr_13__0 (.Q (d_arr_13__0), .D (nx3132), .CLK (nx10233)) ;
    inv01 ix3133 (.Y (nx3132), .A (nx8423)) ;
    aoi222 ix8424 (.Y (nx8423), .A0 (d_arr_mux_13__0), .A1 (nx11313), .B0 (
           d_arr_mul_13__0), .B1 (nx10465), .C0 (d_arr_add_13__0), .C1 (nx10657)
           ) ;
    latch lat_d_arr_13__1 (.Q (d_arr_13__1), .D (nx3144), .CLK (nx10233)) ;
    inv01 ix3145 (.Y (nx3144), .A (nx8429)) ;
    aoi222 ix8430 (.Y (nx8429), .A0 (d_arr_mux_13__1), .A1 (nx11313), .B0 (
           d_arr_mul_13__1), .B1 (nx10465), .C0 (d_arr_add_13__1), .C1 (nx10657)
           ) ;
    latch lat_d_arr_13__2 (.Q (d_arr_13__2), .D (nx3156), .CLK (nx10233)) ;
    inv01 ix3157 (.Y (nx3156), .A (nx8435)) ;
    aoi222 ix8436 (.Y (nx8435), .A0 (d_arr_mux_13__2), .A1 (nx11313), .B0 (
           d_arr_mul_13__2), .B1 (nx10465), .C0 (d_arr_add_13__2), .C1 (nx10657)
           ) ;
    latch lat_d_arr_13__3 (.Q (d_arr_13__3), .D (nx3168), .CLK (nx10233)) ;
    inv01 ix3169 (.Y (nx3168), .A (nx8441)) ;
    aoi222 ix8442 (.Y (nx8441), .A0 (d_arr_mux_13__3), .A1 (nx11313), .B0 (
           d_arr_mul_13__3), .B1 (nx10465), .C0 (d_arr_add_13__3), .C1 (nx10657)
           ) ;
    latch lat_d_arr_13__4 (.Q (d_arr_13__4), .D (nx3180), .CLK (nx10233)) ;
    inv01 ix3181 (.Y (nx3180), .A (nx8447)) ;
    aoi222 ix8448 (.Y (nx8447), .A0 (d_arr_mux_13__4), .A1 (nx11313), .B0 (
           d_arr_mul_13__4), .B1 (nx10465), .C0 (d_arr_add_13__4), .C1 (nx10657)
           ) ;
    latch lat_d_arr_13__5 (.Q (d_arr_13__5), .D (nx3192), .CLK (nx10235)) ;
    inv01 ix3193 (.Y (nx3192), .A (nx8453)) ;
    aoi222 ix8454 (.Y (nx8453), .A0 (d_arr_mux_13__5), .A1 (nx11313), .B0 (
           d_arr_mul_13__5), .B1 (nx10467), .C0 (d_arr_add_13__5), .C1 (nx10659)
           ) ;
    latch lat_d_arr_13__6 (.Q (d_arr_13__6), .D (nx3204), .CLK (nx10235)) ;
    inv01 ix3205 (.Y (nx3204), .A (nx8459)) ;
    aoi222 ix8460 (.Y (nx8459), .A0 (d_arr_mux_13__6), .A1 (nx11315), .B0 (
           d_arr_mul_13__6), .B1 (nx10467), .C0 (d_arr_add_13__6), .C1 (nx10659)
           ) ;
    latch lat_d_arr_13__7 (.Q (d_arr_13__7), .D (nx3216), .CLK (nx10235)) ;
    inv01 ix3217 (.Y (nx3216), .A (nx8465)) ;
    aoi222 ix8466 (.Y (nx8465), .A0 (d_arr_mux_13__7), .A1 (nx11315), .B0 (
           d_arr_mul_13__7), .B1 (nx10467), .C0 (d_arr_add_13__7), .C1 (nx10659)
           ) ;
    latch lat_d_arr_13__8 (.Q (d_arr_13__8), .D (nx3228), .CLK (nx10235)) ;
    inv01 ix3229 (.Y (nx3228), .A (nx8471)) ;
    aoi222 ix8472 (.Y (nx8471), .A0 (d_arr_mux_13__8), .A1 (nx11315), .B0 (
           d_arr_mul_13__8), .B1 (nx10467), .C0 (d_arr_add_13__8), .C1 (nx10659)
           ) ;
    latch lat_d_arr_13__9 (.Q (d_arr_13__9), .D (nx3240), .CLK (nx10235)) ;
    inv01 ix3241 (.Y (nx3240), .A (nx8477)) ;
    aoi222 ix8478 (.Y (nx8477), .A0 (d_arr_mux_13__9), .A1 (nx11315), .B0 (
           d_arr_mul_13__9), .B1 (nx10467), .C0 (d_arr_add_13__9), .C1 (nx10659)
           ) ;
    latch lat_d_arr_13__10 (.Q (d_arr_13__10), .D (nx3252), .CLK (nx10235)) ;
    inv01 ix3253 (.Y (nx3252), .A (nx8481)) ;
    aoi222 ix8482 (.Y (nx8481), .A0 (d_arr_mux_13__10), .A1 (nx11315), .B0 (
           d_arr_mul_13__10), .B1 (nx10467), .C0 (d_arr_add_13__10), .C1 (
           nx10659)) ;
    latch lat_d_arr_13__11 (.Q (d_arr_13__11), .D (nx3264), .CLK (nx10235)) ;
    inv01 ix3265 (.Y (nx3264), .A (nx8485)) ;
    aoi222 ix8486 (.Y (nx8485), .A0 (d_arr_mux_13__11), .A1 (nx11315), .B0 (
           d_arr_mul_13__11), .B1 (nx10467), .C0 (d_arr_add_13__11), .C1 (
           nx10659)) ;
    latch lat_d_arr_13__12 (.Q (d_arr_13__12), .D (nx3276), .CLK (nx10237)) ;
    inv01 ix3277 (.Y (nx3276), .A (nx8489)) ;
    aoi222 ix8490 (.Y (nx8489), .A0 (d_arr_mux_13__12), .A1 (nx11315), .B0 (
           d_arr_mul_13__12), .B1 (nx10469), .C0 (d_arr_add_13__12), .C1 (
           nx10661)) ;
    latch lat_d_arr_13__13 (.Q (d_arr_13__13), .D (nx3288), .CLK (nx10237)) ;
    inv01 ix3289 (.Y (nx3288), .A (nx8493)) ;
    aoi222 ix8494 (.Y (nx8493), .A0 (d_arr_mux_13__13), .A1 (nx11317), .B0 (
           d_arr_mul_13__13), .B1 (nx10469), .C0 (d_arr_add_13__13), .C1 (
           nx10661)) ;
    latch lat_d_arr_13__14 (.Q (d_arr_13__14), .D (nx3300), .CLK (nx10237)) ;
    inv01 ix3301 (.Y (nx3300), .A (nx8497)) ;
    aoi222 ix8498 (.Y (nx8497), .A0 (d_arr_mux_13__14), .A1 (nx11317), .B0 (
           d_arr_mul_13__14), .B1 (nx10469), .C0 (d_arr_add_13__14), .C1 (
           nx10661)) ;
    latch lat_d_arr_13__15 (.Q (d_arr_13__15), .D (nx3312), .CLK (nx10237)) ;
    inv01 ix3313 (.Y (nx3312), .A (nx8501)) ;
    aoi222 ix8502 (.Y (nx8501), .A0 (d_arr_mux_13__15), .A1 (nx11317), .B0 (
           d_arr_mul_13__15), .B1 (nx10469), .C0 (d_arr_add_13__15), .C1 (
           nx10661)) ;
    latch lat_d_arr_13__16 (.Q (d_arr_13__16), .D (nx3324), .CLK (nx10237)) ;
    inv01 ix3325 (.Y (nx3324), .A (nx8505)) ;
    aoi222 ix8506 (.Y (nx8505), .A0 (d_arr_mux_13__16), .A1 (nx11317), .B0 (
           d_arr_mul_13__16), .B1 (nx10469), .C0 (d_arr_add_13__16), .C1 (
           nx10661)) ;
    latch lat_d_arr_13__17 (.Q (d_arr_13__17), .D (nx3336), .CLK (nx10237)) ;
    inv01 ix3337 (.Y (nx3336), .A (nx8509)) ;
    aoi222 ix8510 (.Y (nx8509), .A0 (d_arr_mux_13__17), .A1 (nx11317), .B0 (
           d_arr_mul_13__17), .B1 (nx10469), .C0 (d_arr_add_13__17), .C1 (
           nx10661)) ;
    latch lat_d_arr_13__18 (.Q (d_arr_13__18), .D (nx3348), .CLK (nx10237)) ;
    inv01 ix3349 (.Y (nx3348), .A (nx8513)) ;
    aoi222 ix8514 (.Y (nx8513), .A0 (d_arr_mux_13__18), .A1 (nx11317), .B0 (
           d_arr_mul_13__18), .B1 (nx10469), .C0 (d_arr_add_13__18), .C1 (
           nx10661)) ;
    latch lat_d_arr_13__19 (.Q (d_arr_13__19), .D (nx3360), .CLK (nx10239)) ;
    inv01 ix3361 (.Y (nx3360), .A (nx8517)) ;
    aoi222 ix8518 (.Y (nx8517), .A0 (d_arr_mux_13__19), .A1 (nx11317), .B0 (
           d_arr_mul_13__19), .B1 (nx10471), .C0 (d_arr_add_13__19), .C1 (
           nx10663)) ;
    latch lat_d_arr_13__20 (.Q (d_arr_13__20), .D (nx3372), .CLK (nx10239)) ;
    inv01 ix3373 (.Y (nx3372), .A (nx8521)) ;
    aoi222 ix8522 (.Y (nx8521), .A0 (d_arr_mux_13__20), .A1 (nx11319), .B0 (
           d_arr_mul_13__20), .B1 (nx10471), .C0 (d_arr_add_13__20), .C1 (
           nx10663)) ;
    latch lat_d_arr_13__21 (.Q (d_arr_13__21), .D (nx3384), .CLK (nx10239)) ;
    inv01 ix3385 (.Y (nx3384), .A (nx8525)) ;
    aoi222 ix8526 (.Y (nx8525), .A0 (d_arr_mux_13__21), .A1 (nx11319), .B0 (
           d_arr_mul_13__21), .B1 (nx10471), .C0 (d_arr_add_13__21), .C1 (
           nx10663)) ;
    latch lat_d_arr_13__22 (.Q (d_arr_13__22), .D (nx3396), .CLK (nx10239)) ;
    inv01 ix3397 (.Y (nx3396), .A (nx8529)) ;
    aoi222 ix8530 (.Y (nx8529), .A0 (d_arr_mux_13__22), .A1 (nx11319), .B0 (
           d_arr_mul_13__22), .B1 (nx10471), .C0 (d_arr_add_13__22), .C1 (
           nx10663)) ;
    latch lat_d_arr_13__23 (.Q (d_arr_13__23), .D (nx3408), .CLK (nx10239)) ;
    inv01 ix3409 (.Y (nx3408), .A (nx8533)) ;
    aoi222 ix8534 (.Y (nx8533), .A0 (d_arr_mux_13__23), .A1 (nx11319), .B0 (
           d_arr_mul_13__23), .B1 (nx10471), .C0 (d_arr_add_13__23), .C1 (
           nx10663)) ;
    latch lat_d_arr_13__24 (.Q (d_arr_13__24), .D (nx3420), .CLK (nx10239)) ;
    inv01 ix3421 (.Y (nx3420), .A (nx8537)) ;
    aoi222 ix8538 (.Y (nx8537), .A0 (d_arr_mux_13__24), .A1 (nx11319), .B0 (
           d_arr_mul_13__24), .B1 (nx10471), .C0 (d_arr_add_13__24), .C1 (
           nx10663)) ;
    latch lat_d_arr_13__25 (.Q (d_arr_13__25), .D (nx3432), .CLK (nx10239)) ;
    inv01 ix3433 (.Y (nx3432), .A (nx8541)) ;
    aoi222 ix8542 (.Y (nx8541), .A0 (d_arr_mux_13__25), .A1 (nx11319), .B0 (
           d_arr_mul_13__25), .B1 (nx10471), .C0 (d_arr_add_13__25), .C1 (
           nx10663)) ;
    latch lat_d_arr_13__26 (.Q (d_arr_13__26), .D (nx3444), .CLK (nx10241)) ;
    inv01 ix3445 (.Y (nx3444), .A (nx8545)) ;
    aoi222 ix8546 (.Y (nx8545), .A0 (d_arr_mux_13__26), .A1 (nx11319), .B0 (
           d_arr_mul_13__26), .B1 (nx10473), .C0 (d_arr_add_13__26), .C1 (
           nx10665)) ;
    latch lat_d_arr_13__27 (.Q (d_arr_13__27), .D (nx3456), .CLK (nx10241)) ;
    inv01 ix3457 (.Y (nx3456), .A (nx8549)) ;
    aoi222 ix8550 (.Y (nx8549), .A0 (d_arr_mux_13__27), .A1 (nx11321), .B0 (
           d_arr_mul_13__27), .B1 (nx10473), .C0 (d_arr_add_13__27), .C1 (
           nx10665)) ;
    latch lat_d_arr_13__28 (.Q (d_arr_13__28), .D (nx3468), .CLK (nx10241)) ;
    inv01 ix3469 (.Y (nx3468), .A (nx8553)) ;
    aoi222 ix8554 (.Y (nx8553), .A0 (d_arr_mux_13__28), .A1 (nx11321), .B0 (
           d_arr_mul_13__28), .B1 (nx10473), .C0 (d_arr_add_13__28), .C1 (
           nx10665)) ;
    latch lat_d_arr_13__29 (.Q (d_arr_13__29), .D (nx3480), .CLK (nx10241)) ;
    inv01 ix3481 (.Y (nx3480), .A (nx8557)) ;
    aoi222 ix8558 (.Y (nx8557), .A0 (d_arr_mux_13__29), .A1 (nx11321), .B0 (
           d_arr_mul_13__29), .B1 (nx10473), .C0 (d_arr_add_13__29), .C1 (
           nx10665)) ;
    latch lat_d_arr_13__30 (.Q (d_arr_13__30), .D (nx3492), .CLK (nx10241)) ;
    inv01 ix3493 (.Y (nx3492), .A (nx8561)) ;
    aoi222 ix8562 (.Y (nx8561), .A0 (d_arr_mux_13__30), .A1 (nx11321), .B0 (
           d_arr_mul_13__30), .B1 (nx10473), .C0 (d_arr_add_13__30), .C1 (
           nx10665)) ;
    latch lat_d_arr_13__31 (.Q (d_arr_13__31), .D (nx3504), .CLK (nx10241)) ;
    inv01 ix3505 (.Y (nx3504), .A (nx8565)) ;
    aoi222 ix8566 (.Y (nx8565), .A0 (d_arr_mux_13__31), .A1 (nx11321), .B0 (
           d_arr_mul_13__31), .B1 (nx10473), .C0 (d_arr_add_13__31), .C1 (
           nx10665)) ;
    latch lat_d_arr_12__0 (.Q (d_arr_12__0), .D (nx3516), .CLK (nx10241)) ;
    inv01 ix3517 (.Y (nx3516), .A (nx8569)) ;
    aoi222 ix8570 (.Y (nx8569), .A0 (d_arr_mux_12__0), .A1 (nx11321), .B0 (
           d_arr_mul_12__0), .B1 (nx10473), .C0 (d_arr_add_12__0), .C1 (nx10665)
           ) ;
    latch lat_d_arr_12__1 (.Q (d_arr_12__1), .D (nx3528), .CLK (nx10243)) ;
    inv01 ix3529 (.Y (nx3528), .A (nx8573)) ;
    aoi222 ix8574 (.Y (nx8573), .A0 (d_arr_mux_12__1), .A1 (nx11321), .B0 (
           d_arr_mul_12__1), .B1 (nx10475), .C0 (d_arr_add_12__1), .C1 (nx10667)
           ) ;
    latch lat_d_arr_12__2 (.Q (d_arr_12__2), .D (nx3540), .CLK (nx10243)) ;
    inv01 ix3541 (.Y (nx3540), .A (nx8577)) ;
    aoi222 ix8578 (.Y (nx8577), .A0 (d_arr_mux_12__2), .A1 (nx11323), .B0 (
           d_arr_mul_12__2), .B1 (nx10475), .C0 (d_arr_add_12__2), .C1 (nx10667)
           ) ;
    latch lat_d_arr_12__3 (.Q (d_arr_12__3), .D (nx3552), .CLK (nx10243)) ;
    inv01 ix3553 (.Y (nx3552), .A (nx8581)) ;
    aoi222 ix8582 (.Y (nx8581), .A0 (d_arr_mux_12__3), .A1 (nx11323), .B0 (
           d_arr_mul_12__3), .B1 (nx10475), .C0 (d_arr_add_12__3), .C1 (nx10667)
           ) ;
    latch lat_d_arr_12__4 (.Q (d_arr_12__4), .D (nx3564), .CLK (nx10243)) ;
    inv01 ix3565 (.Y (nx3564), .A (nx8585)) ;
    aoi222 ix8586 (.Y (nx8585), .A0 (d_arr_mux_12__4), .A1 (nx11323), .B0 (
           d_arr_mul_12__4), .B1 (nx10475), .C0 (d_arr_add_12__4), .C1 (nx10667)
           ) ;
    latch lat_d_arr_12__5 (.Q (d_arr_12__5), .D (nx3576), .CLK (nx10243)) ;
    inv01 ix3577 (.Y (nx3576), .A (nx8589)) ;
    aoi222 ix8590 (.Y (nx8589), .A0 (d_arr_mux_12__5), .A1 (nx11323), .B0 (
           d_arr_mul_12__5), .B1 (nx10475), .C0 (d_arr_add_12__5), .C1 (nx10667)
           ) ;
    latch lat_d_arr_12__6 (.Q (d_arr_12__6), .D (nx3588), .CLK (nx10243)) ;
    inv01 ix3589 (.Y (nx3588), .A (nx8593)) ;
    aoi222 ix8594 (.Y (nx8593), .A0 (d_arr_mux_12__6), .A1 (nx11323), .B0 (
           d_arr_mul_12__6), .B1 (nx10475), .C0 (d_arr_add_12__6), .C1 (nx10667)
           ) ;
    latch lat_d_arr_12__7 (.Q (d_arr_12__7), .D (nx3600), .CLK (nx10243)) ;
    inv01 ix3601 (.Y (nx3600), .A (nx8597)) ;
    aoi222 ix8598 (.Y (nx8597), .A0 (d_arr_mux_12__7), .A1 (nx11323), .B0 (
           d_arr_mul_12__7), .B1 (nx10475), .C0 (d_arr_add_12__7), .C1 (nx10667)
           ) ;
    latch lat_d_arr_12__8 (.Q (d_arr_12__8), .D (nx3612), .CLK (nx10245)) ;
    inv01 ix3613 (.Y (nx3612), .A (nx8601)) ;
    aoi222 ix8602 (.Y (nx8601), .A0 (d_arr_mux_12__8), .A1 (nx11323), .B0 (
           d_arr_mul_12__8), .B1 (nx10477), .C0 (d_arr_add_12__8), .C1 (nx10669)
           ) ;
    latch lat_d_arr_12__9 (.Q (d_arr_12__9), .D (nx3624), .CLK (nx10245)) ;
    inv01 ix3625 (.Y (nx3624), .A (nx8605)) ;
    aoi222 ix8606 (.Y (nx8605), .A0 (d_arr_mux_12__9), .A1 (nx11325), .B0 (
           d_arr_mul_12__9), .B1 (nx10477), .C0 (d_arr_add_12__9), .C1 (nx10669)
           ) ;
    latch lat_d_arr_12__10 (.Q (d_arr_12__10), .D (nx3636), .CLK (nx10245)) ;
    inv01 ix3637 (.Y (nx3636), .A (nx8609)) ;
    aoi222 ix8610 (.Y (nx8609), .A0 (d_arr_mux_12__10), .A1 (nx11325), .B0 (
           d_arr_mul_12__10), .B1 (nx10477), .C0 (d_arr_add_12__10), .C1 (
           nx10669)) ;
    latch lat_d_arr_12__11 (.Q (d_arr_12__11), .D (nx3648), .CLK (nx10245)) ;
    inv01 ix3649 (.Y (nx3648), .A (nx8613)) ;
    aoi222 ix8614 (.Y (nx8613), .A0 (d_arr_mux_12__11), .A1 (nx11325), .B0 (
           d_arr_mul_12__11), .B1 (nx10477), .C0 (d_arr_add_12__11), .C1 (
           nx10669)) ;
    latch lat_d_arr_12__12 (.Q (d_arr_12__12), .D (nx3660), .CLK (nx10245)) ;
    inv01 ix3661 (.Y (nx3660), .A (nx8617)) ;
    aoi222 ix8618 (.Y (nx8617), .A0 (d_arr_mux_12__12), .A1 (nx11325), .B0 (
           d_arr_mul_12__12), .B1 (nx10477), .C0 (d_arr_add_12__12), .C1 (
           nx10669)) ;
    latch lat_d_arr_12__13 (.Q (d_arr_12__13), .D (nx3672), .CLK (nx10245)) ;
    inv01 ix3673 (.Y (nx3672), .A (nx8621)) ;
    aoi222 ix8622 (.Y (nx8621), .A0 (d_arr_mux_12__13), .A1 (nx11325), .B0 (
           d_arr_mul_12__13), .B1 (nx10477), .C0 (d_arr_add_12__13), .C1 (
           nx10669)) ;
    latch lat_d_arr_12__14 (.Q (d_arr_12__14), .D (nx3684), .CLK (nx10245)) ;
    inv01 ix3685 (.Y (nx3684), .A (nx8625)) ;
    aoi222 ix8626 (.Y (nx8625), .A0 (d_arr_mux_12__14), .A1 (nx11325), .B0 (
           d_arr_mul_12__14), .B1 (nx10477), .C0 (d_arr_add_12__14), .C1 (
           nx10669)) ;
    latch lat_d_arr_12__15 (.Q (d_arr_12__15), .D (nx3696), .CLK (nx10247)) ;
    inv01 ix3697 (.Y (nx3696), .A (nx8629)) ;
    aoi222 ix8630 (.Y (nx8629), .A0 (d_arr_mux_12__15), .A1 (nx11325), .B0 (
           d_arr_mul_12__15), .B1 (nx10479), .C0 (d_arr_add_12__15), .C1 (
           nx10671)) ;
    latch lat_d_arr_12__16 (.Q (d_arr_12__16), .D (nx3708), .CLK (nx10247)) ;
    inv01 ix3709 (.Y (nx3708), .A (nx8633)) ;
    aoi222 ix8634 (.Y (nx8633), .A0 (d_arr_mux_12__16), .A1 (nx11327), .B0 (
           d_arr_mul_12__16), .B1 (nx10479), .C0 (d_arr_add_12__16), .C1 (
           nx10671)) ;
    latch lat_d_arr_12__17 (.Q (d_arr_12__17), .D (nx3720), .CLK (nx10247)) ;
    inv01 ix3721 (.Y (nx3720), .A (nx8637)) ;
    aoi222 ix8638 (.Y (nx8637), .A0 (d_arr_mux_12__17), .A1 (nx11327), .B0 (
           d_arr_mul_12__17), .B1 (nx10479), .C0 (d_arr_add_12__17), .C1 (
           nx10671)) ;
    latch lat_d_arr_12__18 (.Q (d_arr_12__18), .D (nx3732), .CLK (nx10247)) ;
    inv01 ix3733 (.Y (nx3732), .A (nx8641)) ;
    aoi222 ix8642 (.Y (nx8641), .A0 (d_arr_mux_12__18), .A1 (nx11327), .B0 (
           d_arr_mul_12__18), .B1 (nx10479), .C0 (d_arr_add_12__18), .C1 (
           nx10671)) ;
    latch lat_d_arr_12__19 (.Q (d_arr_12__19), .D (nx3744), .CLK (nx10247)) ;
    inv01 ix3745 (.Y (nx3744), .A (nx8645)) ;
    aoi222 ix8646 (.Y (nx8645), .A0 (d_arr_mux_12__19), .A1 (nx11327), .B0 (
           d_arr_mul_12__19), .B1 (nx10479), .C0 (d_arr_add_12__19), .C1 (
           nx10671)) ;
    latch lat_d_arr_12__20 (.Q (d_arr_12__20), .D (nx3756), .CLK (nx10247)) ;
    inv01 ix3757 (.Y (nx3756), .A (nx8649)) ;
    aoi222 ix8650 (.Y (nx8649), .A0 (d_arr_mux_12__20), .A1 (nx11327), .B0 (
           d_arr_mul_12__20), .B1 (nx10479), .C0 (d_arr_add_12__20), .C1 (
           nx10671)) ;
    latch lat_d_arr_12__21 (.Q (d_arr_12__21), .D (nx3768), .CLK (nx10247)) ;
    inv01 ix3769 (.Y (nx3768), .A (nx8653)) ;
    aoi222 ix8654 (.Y (nx8653), .A0 (d_arr_mux_12__21), .A1 (nx11327), .B0 (
           d_arr_mul_12__21), .B1 (nx10479), .C0 (d_arr_add_12__21), .C1 (
           nx10671)) ;
    latch lat_d_arr_12__22 (.Q (d_arr_12__22), .D (nx3780), .CLK (nx10249)) ;
    inv01 ix3781 (.Y (nx3780), .A (nx8657)) ;
    aoi222 ix8658 (.Y (nx8657), .A0 (d_arr_mux_12__22), .A1 (nx11327), .B0 (
           d_arr_mul_12__22), .B1 (nx10481), .C0 (d_arr_add_12__22), .C1 (
           nx10673)) ;
    latch lat_d_arr_12__23 (.Q (d_arr_12__23), .D (nx3792), .CLK (nx10249)) ;
    inv01 ix3793 (.Y (nx3792), .A (nx8661)) ;
    aoi222 ix8662 (.Y (nx8661), .A0 (d_arr_mux_12__23), .A1 (nx11329), .B0 (
           d_arr_mul_12__23), .B1 (nx10481), .C0 (d_arr_add_12__23), .C1 (
           nx10673)) ;
    latch lat_d_arr_12__24 (.Q (d_arr_12__24), .D (nx3804), .CLK (nx10249)) ;
    inv01 ix3805 (.Y (nx3804), .A (nx8665)) ;
    aoi222 ix8666 (.Y (nx8665), .A0 (d_arr_mux_12__24), .A1 (nx11329), .B0 (
           d_arr_mul_12__24), .B1 (nx10481), .C0 (d_arr_add_12__24), .C1 (
           nx10673)) ;
    latch lat_d_arr_12__25 (.Q (d_arr_12__25), .D (nx3816), .CLK (nx10249)) ;
    inv01 ix3817 (.Y (nx3816), .A (nx8669)) ;
    aoi222 ix8670 (.Y (nx8669), .A0 (d_arr_mux_12__25), .A1 (nx11329), .B0 (
           d_arr_mul_12__25), .B1 (nx10481), .C0 (d_arr_add_12__25), .C1 (
           nx10673)) ;
    latch lat_d_arr_12__26 (.Q (d_arr_12__26), .D (nx3828), .CLK (nx10249)) ;
    inv01 ix3829 (.Y (nx3828), .A (nx8673)) ;
    aoi222 ix8674 (.Y (nx8673), .A0 (d_arr_mux_12__26), .A1 (nx11329), .B0 (
           d_arr_mul_12__26), .B1 (nx10481), .C0 (d_arr_add_12__26), .C1 (
           nx10673)) ;
    latch lat_d_arr_12__27 (.Q (d_arr_12__27), .D (nx3840), .CLK (nx10249)) ;
    inv01 ix3841 (.Y (nx3840), .A (nx8677)) ;
    aoi222 ix8678 (.Y (nx8677), .A0 (d_arr_mux_12__27), .A1 (nx11329), .B0 (
           d_arr_mul_12__27), .B1 (nx10481), .C0 (d_arr_add_12__27), .C1 (
           nx10673)) ;
    latch lat_d_arr_12__28 (.Q (d_arr_12__28), .D (nx3852), .CLK (nx10249)) ;
    inv01 ix3853 (.Y (nx3852), .A (nx8681)) ;
    aoi222 ix8682 (.Y (nx8681), .A0 (d_arr_mux_12__28), .A1 (nx11329), .B0 (
           d_arr_mul_12__28), .B1 (nx10481), .C0 (d_arr_add_12__28), .C1 (
           nx10673)) ;
    latch lat_d_arr_12__29 (.Q (d_arr_12__29), .D (nx3864), .CLK (nx10251)) ;
    inv01 ix3865 (.Y (nx3864), .A (nx8685)) ;
    aoi222 ix8686 (.Y (nx8685), .A0 (d_arr_mux_12__29), .A1 (nx11329), .B0 (
           d_arr_mul_12__29), .B1 (nx10483), .C0 (d_arr_add_12__29), .C1 (
           nx10675)) ;
    latch lat_d_arr_12__30 (.Q (d_arr_12__30), .D (nx3876), .CLK (nx10251)) ;
    inv01 ix3877 (.Y (nx3876), .A (nx8689)) ;
    aoi222 ix8690 (.Y (nx8689), .A0 (d_arr_mux_12__30), .A1 (nx11331), .B0 (
           d_arr_mul_12__30), .B1 (nx10483), .C0 (d_arr_add_12__30), .C1 (
           nx10675)) ;
    latch lat_d_arr_12__31 (.Q (d_arr_12__31), .D (nx3888), .CLK (nx10251)) ;
    inv01 ix3889 (.Y (nx3888), .A (nx8693)) ;
    aoi222 ix8694 (.Y (nx8693), .A0 (d_arr_mux_12__31), .A1 (nx11331), .B0 (
           d_arr_mul_12__31), .B1 (nx10483), .C0 (d_arr_add_12__31), .C1 (
           nx10675)) ;
    latch lat_d_arr_11__0 (.Q (d_arr_11__0), .D (nx3900), .CLK (nx10251)) ;
    inv01 ix3901 (.Y (nx3900), .A (nx8697)) ;
    aoi222 ix8698 (.Y (nx8697), .A0 (d_arr_mux_11__0), .A1 (nx11331), .B0 (
           d_arr_mul_11__0), .B1 (nx10483), .C0 (d_arr_add_11__0), .C1 (nx10675)
           ) ;
    latch lat_d_arr_11__1 (.Q (d_arr_11__1), .D (nx3912), .CLK (nx10251)) ;
    inv01 ix3913 (.Y (nx3912), .A (nx8701)) ;
    aoi222 ix8702 (.Y (nx8701), .A0 (d_arr_mux_11__1), .A1 (nx11331), .B0 (
           d_arr_mul_11__1), .B1 (nx10483), .C0 (d_arr_add_11__1), .C1 (nx10675)
           ) ;
    latch lat_d_arr_11__2 (.Q (d_arr_11__2), .D (nx3924), .CLK (nx10251)) ;
    inv01 ix3925 (.Y (nx3924), .A (nx8705)) ;
    aoi222 ix8706 (.Y (nx8705), .A0 (d_arr_mux_11__2), .A1 (nx11331), .B0 (
           d_arr_mul_11__2), .B1 (nx10483), .C0 (d_arr_add_11__2), .C1 (nx10675)
           ) ;
    latch lat_d_arr_11__3 (.Q (d_arr_11__3), .D (nx3936), .CLK (nx10251)) ;
    inv01 ix3937 (.Y (nx3936), .A (nx8709)) ;
    aoi222 ix8710 (.Y (nx8709), .A0 (d_arr_mux_11__3), .A1 (nx11331), .B0 (
           d_arr_mul_11__3), .B1 (nx10483), .C0 (d_arr_add_11__3), .C1 (nx10675)
           ) ;
    latch lat_d_arr_11__4 (.Q (d_arr_11__4), .D (nx3948), .CLK (nx10253)) ;
    inv01 ix3949 (.Y (nx3948), .A (nx8713)) ;
    aoi222 ix8714 (.Y (nx8713), .A0 (d_arr_mux_11__4), .A1 (nx11331), .B0 (
           d_arr_mul_11__4), .B1 (nx10485), .C0 (d_arr_add_11__4), .C1 (nx10677)
           ) ;
    latch lat_d_arr_11__5 (.Q (d_arr_11__5), .D (nx3960), .CLK (nx10253)) ;
    inv01 ix3961 (.Y (nx3960), .A (nx8717)) ;
    aoi222 ix8718 (.Y (nx8717), .A0 (d_arr_mux_11__5), .A1 (nx11333), .B0 (
           d_arr_mul_11__5), .B1 (nx10485), .C0 (d_arr_add_11__5), .C1 (nx10677)
           ) ;
    latch lat_d_arr_11__6 (.Q (d_arr_11__6), .D (nx3972), .CLK (nx10253)) ;
    inv01 ix3973 (.Y (nx3972), .A (nx8721)) ;
    aoi222 ix8722 (.Y (nx8721), .A0 (d_arr_mux_11__6), .A1 (nx11333), .B0 (
           d_arr_mul_11__6), .B1 (nx10485), .C0 (d_arr_add_11__6), .C1 (nx10677)
           ) ;
    latch lat_d_arr_11__7 (.Q (d_arr_11__7), .D (nx3984), .CLK (nx10253)) ;
    inv01 ix3985 (.Y (nx3984), .A (nx8725)) ;
    aoi222 ix8726 (.Y (nx8725), .A0 (d_arr_mux_11__7), .A1 (nx11333), .B0 (
           d_arr_mul_11__7), .B1 (nx10485), .C0 (d_arr_add_11__7), .C1 (nx10677)
           ) ;
    latch lat_d_arr_11__8 (.Q (d_arr_11__8), .D (nx3996), .CLK (nx10253)) ;
    inv01 ix3997 (.Y (nx3996), .A (nx8729)) ;
    aoi222 ix8730 (.Y (nx8729), .A0 (d_arr_mux_11__8), .A1 (nx11333), .B0 (
           d_arr_mul_11__8), .B1 (nx10485), .C0 (d_arr_add_11__8), .C1 (nx10677)
           ) ;
    latch lat_d_arr_11__9 (.Q (d_arr_11__9), .D (nx4008), .CLK (nx10253)) ;
    inv01 ix4009 (.Y (nx4008), .A (nx8733)) ;
    aoi222 ix8734 (.Y (nx8733), .A0 (d_arr_mux_11__9), .A1 (nx11333), .B0 (
           d_arr_mul_11__9), .B1 (nx10485), .C0 (d_arr_add_11__9), .C1 (nx10677)
           ) ;
    latch lat_d_arr_11__10 (.Q (d_arr_11__10), .D (nx4020), .CLK (nx10253)) ;
    inv01 ix4021 (.Y (nx4020), .A (nx8737)) ;
    aoi222 ix8738 (.Y (nx8737), .A0 (d_arr_mux_11__10), .A1 (nx11333), .B0 (
           d_arr_mul_11__10), .B1 (nx10485), .C0 (d_arr_add_11__10), .C1 (
           nx10677)) ;
    latch lat_d_arr_11__11 (.Q (d_arr_11__11), .D (nx4032), .CLK (nx10255)) ;
    inv01 ix4033 (.Y (nx4032), .A (nx8741)) ;
    aoi222 ix8742 (.Y (nx8741), .A0 (d_arr_mux_11__11), .A1 (nx11333), .B0 (
           d_arr_mul_11__11), .B1 (nx10487), .C0 (d_arr_add_11__11), .C1 (
           nx10679)) ;
    latch lat_d_arr_11__12 (.Q (d_arr_11__12), .D (nx4044), .CLK (nx10255)) ;
    inv01 ix4045 (.Y (nx4044), .A (nx8745)) ;
    aoi222 ix8746 (.Y (nx8745), .A0 (d_arr_mux_11__12), .A1 (nx11335), .B0 (
           d_arr_mul_11__12), .B1 (nx10487), .C0 (d_arr_add_11__12), .C1 (
           nx10679)) ;
    latch lat_d_arr_11__13 (.Q (d_arr_11__13), .D (nx4056), .CLK (nx10255)) ;
    inv01 ix4057 (.Y (nx4056), .A (nx8749)) ;
    aoi222 ix8750 (.Y (nx8749), .A0 (d_arr_mux_11__13), .A1 (nx11335), .B0 (
           d_arr_mul_11__13), .B1 (nx10487), .C0 (d_arr_add_11__13), .C1 (
           nx10679)) ;
    latch lat_d_arr_11__14 (.Q (d_arr_11__14), .D (nx4068), .CLK (nx10255)) ;
    inv01 ix4069 (.Y (nx4068), .A (nx8753)) ;
    aoi222 ix8754 (.Y (nx8753), .A0 (d_arr_mux_11__14), .A1 (nx11335), .B0 (
           d_arr_mul_11__14), .B1 (nx10487), .C0 (d_arr_add_11__14), .C1 (
           nx10679)) ;
    latch lat_d_arr_11__15 (.Q (d_arr_11__15), .D (nx4080), .CLK (nx10255)) ;
    inv01 ix4081 (.Y (nx4080), .A (nx8757)) ;
    aoi222 ix8758 (.Y (nx8757), .A0 (d_arr_mux_11__15), .A1 (nx11335), .B0 (
           d_arr_mul_11__15), .B1 (nx10487), .C0 (d_arr_add_11__15), .C1 (
           nx10679)) ;
    latch lat_d_arr_11__16 (.Q (d_arr_11__16), .D (nx4092), .CLK (nx10255)) ;
    inv01 ix4093 (.Y (nx4092), .A (nx8761)) ;
    aoi222 ix8762 (.Y (nx8761), .A0 (d_arr_mux_11__16), .A1 (nx11335), .B0 (
           d_arr_mul_11__16), .B1 (nx10487), .C0 (d_arr_add_11__16), .C1 (
           nx10679)) ;
    latch lat_d_arr_11__17 (.Q (d_arr_11__17), .D (nx4104), .CLK (nx10255)) ;
    inv01 ix4105 (.Y (nx4104), .A (nx8765)) ;
    aoi222 ix8766 (.Y (nx8765), .A0 (d_arr_mux_11__17), .A1 (nx11335), .B0 (
           d_arr_mul_11__17), .B1 (nx10487), .C0 (d_arr_add_11__17), .C1 (
           nx10679)) ;
    latch lat_d_arr_11__18 (.Q (d_arr_11__18), .D (nx4116), .CLK (nx10257)) ;
    inv01 ix4117 (.Y (nx4116), .A (nx8769)) ;
    aoi222 ix8770 (.Y (nx8769), .A0 (d_arr_mux_11__18), .A1 (nx11335), .B0 (
           d_arr_mul_11__18), .B1 (nx10489), .C0 (d_arr_add_11__18), .C1 (
           nx10681)) ;
    latch lat_d_arr_11__19 (.Q (d_arr_11__19), .D (nx4128), .CLK (nx10257)) ;
    inv01 ix4129 (.Y (nx4128), .A (nx8773)) ;
    aoi222 ix8774 (.Y (nx8773), .A0 (d_arr_mux_11__19), .A1 (nx11337), .B0 (
           d_arr_mul_11__19), .B1 (nx10489), .C0 (d_arr_add_11__19), .C1 (
           nx10681)) ;
    latch lat_d_arr_11__20 (.Q (d_arr_11__20), .D (nx4140), .CLK (nx10257)) ;
    inv01 ix4141 (.Y (nx4140), .A (nx8777)) ;
    aoi222 ix8778 (.Y (nx8777), .A0 (d_arr_mux_11__20), .A1 (nx11337), .B0 (
           d_arr_mul_11__20), .B1 (nx10489), .C0 (d_arr_add_11__20), .C1 (
           nx10681)) ;
    latch lat_d_arr_11__21 (.Q (d_arr_11__21), .D (nx4152), .CLK (nx10257)) ;
    inv01 ix4153 (.Y (nx4152), .A (nx8781)) ;
    aoi222 ix8782 (.Y (nx8781), .A0 (d_arr_mux_11__21), .A1 (nx11337), .B0 (
           d_arr_mul_11__21), .B1 (nx10489), .C0 (d_arr_add_11__21), .C1 (
           nx10681)) ;
    latch lat_d_arr_11__22 (.Q (d_arr_11__22), .D (nx4164), .CLK (nx10257)) ;
    inv01 ix4165 (.Y (nx4164), .A (nx8785)) ;
    aoi222 ix8786 (.Y (nx8785), .A0 (d_arr_mux_11__22), .A1 (nx11337), .B0 (
           d_arr_mul_11__22), .B1 (nx10489), .C0 (d_arr_add_11__22), .C1 (
           nx10681)) ;
    latch lat_d_arr_11__23 (.Q (d_arr_11__23), .D (nx4176), .CLK (nx10257)) ;
    inv01 ix4177 (.Y (nx4176), .A (nx8789)) ;
    aoi222 ix8790 (.Y (nx8789), .A0 (d_arr_mux_11__23), .A1 (nx11337), .B0 (
           d_arr_mul_11__23), .B1 (nx10489), .C0 (d_arr_add_11__23), .C1 (
           nx10681)) ;
    latch lat_d_arr_11__24 (.Q (d_arr_11__24), .D (nx4188), .CLK (nx10257)) ;
    inv01 ix4189 (.Y (nx4188), .A (nx8793)) ;
    aoi222 ix8794 (.Y (nx8793), .A0 (d_arr_mux_11__24), .A1 (nx11337), .B0 (
           d_arr_mul_11__24), .B1 (nx10489), .C0 (d_arr_add_11__24), .C1 (
           nx10681)) ;
    latch lat_d_arr_11__25 (.Q (d_arr_11__25), .D (nx4200), .CLK (nx10259)) ;
    inv01 ix4201 (.Y (nx4200), .A (nx8797)) ;
    aoi222 ix8798 (.Y (nx8797), .A0 (d_arr_mux_11__25), .A1 (nx11337), .B0 (
           d_arr_mul_11__25), .B1 (nx10491), .C0 (d_arr_add_11__25), .C1 (
           nx10683)) ;
    latch lat_d_arr_11__26 (.Q (d_arr_11__26), .D (nx4212), .CLK (nx10259)) ;
    inv01 ix4213 (.Y (nx4212), .A (nx8801)) ;
    aoi222 ix8802 (.Y (nx8801), .A0 (d_arr_mux_11__26), .A1 (nx11339), .B0 (
           d_arr_mul_11__26), .B1 (nx10491), .C0 (d_arr_add_11__26), .C1 (
           nx10683)) ;
    latch lat_d_arr_11__27 (.Q (d_arr_11__27), .D (nx4224), .CLK (nx10259)) ;
    inv01 ix4225 (.Y (nx4224), .A (nx8805)) ;
    aoi222 ix8806 (.Y (nx8805), .A0 (d_arr_mux_11__27), .A1 (nx11339), .B0 (
           d_arr_mul_11__27), .B1 (nx10491), .C0 (d_arr_add_11__27), .C1 (
           nx10683)) ;
    latch lat_d_arr_11__28 (.Q (d_arr_11__28), .D (nx4236), .CLK (nx10259)) ;
    inv01 ix4237 (.Y (nx4236), .A (nx8809)) ;
    aoi222 ix8810 (.Y (nx8809), .A0 (d_arr_mux_11__28), .A1 (nx11339), .B0 (
           d_arr_mul_11__28), .B1 (nx10491), .C0 (d_arr_add_11__28), .C1 (
           nx10683)) ;
    latch lat_d_arr_11__29 (.Q (d_arr_11__29), .D (nx4248), .CLK (nx10259)) ;
    inv01 ix4249 (.Y (nx4248), .A (nx8813)) ;
    aoi222 ix8814 (.Y (nx8813), .A0 (d_arr_mux_11__29), .A1 (nx11339), .B0 (
           d_arr_mul_11__29), .B1 (nx10491), .C0 (d_arr_add_11__29), .C1 (
           nx10683)) ;
    latch lat_d_arr_11__30 (.Q (d_arr_11__30), .D (nx4260), .CLK (nx10259)) ;
    inv01 ix4261 (.Y (nx4260), .A (nx8817)) ;
    aoi222 ix8818 (.Y (nx8817), .A0 (d_arr_mux_11__30), .A1 (nx11339), .B0 (
           d_arr_mul_11__30), .B1 (nx10491), .C0 (d_arr_add_11__30), .C1 (
           nx10683)) ;
    latch lat_d_arr_11__31 (.Q (d_arr_11__31), .D (nx4272), .CLK (nx10259)) ;
    inv01 ix4273 (.Y (nx4272), .A (nx8821)) ;
    aoi222 ix8822 (.Y (nx8821), .A0 (d_arr_mux_11__31), .A1 (nx11339), .B0 (
           d_arr_mul_11__31), .B1 (nx10491), .C0 (d_arr_add_11__31), .C1 (
           nx10683)) ;
    latch lat_d_arr_10__0 (.Q (d_arr_10__0), .D (nx4284), .CLK (nx10261)) ;
    inv01 ix4285 (.Y (nx4284), .A (nx8825)) ;
    aoi222 ix8826 (.Y (nx8825), .A0 (d_arr_mux_10__0), .A1 (nx11339), .B0 (
           d_arr_mul_10__0), .B1 (nx10493), .C0 (d_arr_add_10__0), .C1 (nx10685)
           ) ;
    latch lat_d_arr_10__1 (.Q (d_arr_10__1), .D (nx4296), .CLK (nx10261)) ;
    inv01 ix4297 (.Y (nx4296), .A (nx8829)) ;
    aoi222 ix8830 (.Y (nx8829), .A0 (d_arr_mux_10__1), .A1 (nx11341), .B0 (
           d_arr_mul_10__1), .B1 (nx10493), .C0 (d_arr_add_10__1), .C1 (nx10685)
           ) ;
    latch lat_d_arr_10__2 (.Q (d_arr_10__2), .D (nx4308), .CLK (nx10261)) ;
    inv01 ix4309 (.Y (nx4308), .A (nx8833)) ;
    aoi222 ix8834 (.Y (nx8833), .A0 (d_arr_mux_10__2), .A1 (nx11341), .B0 (
           d_arr_mul_10__2), .B1 (nx10493), .C0 (d_arr_add_10__2), .C1 (nx10685)
           ) ;
    latch lat_d_arr_10__3 (.Q (d_arr_10__3), .D (nx4320), .CLK (nx10261)) ;
    inv01 ix4321 (.Y (nx4320), .A (nx8837)) ;
    aoi222 ix8838 (.Y (nx8837), .A0 (d_arr_mux_10__3), .A1 (nx11341), .B0 (
           d_arr_mul_10__3), .B1 (nx10493), .C0 (d_arr_add_10__3), .C1 (nx10685)
           ) ;
    latch lat_d_arr_10__4 (.Q (d_arr_10__4), .D (nx4332), .CLK (nx10261)) ;
    inv01 ix4333 (.Y (nx4332), .A (nx8841)) ;
    aoi222 ix8842 (.Y (nx8841), .A0 (d_arr_mux_10__4), .A1 (nx11341), .B0 (
           d_arr_mul_10__4), .B1 (nx10493), .C0 (d_arr_add_10__4), .C1 (nx10685)
           ) ;
    latch lat_d_arr_10__5 (.Q (d_arr_10__5), .D (nx4344), .CLK (nx10261)) ;
    inv01 ix4345 (.Y (nx4344), .A (nx8845)) ;
    aoi222 ix8846 (.Y (nx8845), .A0 (d_arr_mux_10__5), .A1 (nx11341), .B0 (
           d_arr_mul_10__5), .B1 (nx10493), .C0 (d_arr_add_10__5), .C1 (nx10685)
           ) ;
    latch lat_d_arr_10__6 (.Q (d_arr_10__6), .D (nx4356), .CLK (nx10261)) ;
    inv01 ix4357 (.Y (nx4356), .A (nx8849)) ;
    aoi222 ix8850 (.Y (nx8849), .A0 (d_arr_mux_10__6), .A1 (nx11341), .B0 (
           d_arr_mul_10__6), .B1 (nx10493), .C0 (d_arr_add_10__6), .C1 (nx10685)
           ) ;
    latch lat_d_arr_10__7 (.Q (d_arr_10__7), .D (nx4368), .CLK (nx10263)) ;
    inv01 ix4369 (.Y (nx4368), .A (nx8853)) ;
    aoi222 ix8854 (.Y (nx8853), .A0 (d_arr_mux_10__7), .A1 (nx11341), .B0 (
           d_arr_mul_10__7), .B1 (nx10495), .C0 (d_arr_add_10__7), .C1 (nx10687)
           ) ;
    latch lat_d_arr_10__8 (.Q (d_arr_10__8), .D (nx4380), .CLK (nx10263)) ;
    inv01 ix4381 (.Y (nx4380), .A (nx8857)) ;
    aoi222 ix8858 (.Y (nx8857), .A0 (d_arr_mux_10__8), .A1 (nx11343), .B0 (
           d_arr_mul_10__8), .B1 (nx10495), .C0 (d_arr_add_10__8), .C1 (nx10687)
           ) ;
    latch lat_d_arr_10__9 (.Q (d_arr_10__9), .D (nx4392), .CLK (nx10263)) ;
    inv01 ix4393 (.Y (nx4392), .A (nx8861)) ;
    aoi222 ix8862 (.Y (nx8861), .A0 (d_arr_mux_10__9), .A1 (nx11343), .B0 (
           d_arr_mul_10__9), .B1 (nx10495), .C0 (d_arr_add_10__9), .C1 (nx10687)
           ) ;
    latch lat_d_arr_10__10 (.Q (d_arr_10__10), .D (nx4404), .CLK (nx10263)) ;
    inv01 ix4405 (.Y (nx4404), .A (nx8865)) ;
    aoi222 ix8866 (.Y (nx8865), .A0 (d_arr_mux_10__10), .A1 (nx11343), .B0 (
           d_arr_mul_10__10), .B1 (nx10495), .C0 (d_arr_add_10__10), .C1 (
           nx10687)) ;
    latch lat_d_arr_10__11 (.Q (d_arr_10__11), .D (nx4416), .CLK (nx10263)) ;
    inv01 ix4417 (.Y (nx4416), .A (nx8869)) ;
    aoi222 ix8870 (.Y (nx8869), .A0 (d_arr_mux_10__11), .A1 (nx11343), .B0 (
           d_arr_mul_10__11), .B1 (nx10495), .C0 (d_arr_add_10__11), .C1 (
           nx10687)) ;
    latch lat_d_arr_10__12 (.Q (d_arr_10__12), .D (nx4428), .CLK (nx10263)) ;
    inv01 ix4429 (.Y (nx4428), .A (nx8873)) ;
    aoi222 ix8874 (.Y (nx8873), .A0 (d_arr_mux_10__12), .A1 (nx11343), .B0 (
           d_arr_mul_10__12), .B1 (nx10495), .C0 (d_arr_add_10__12), .C1 (
           nx10687)) ;
    latch lat_d_arr_10__13 (.Q (d_arr_10__13), .D (nx4440), .CLK (nx10263)) ;
    inv01 ix4441 (.Y (nx4440), .A (nx8877)) ;
    aoi222 ix8878 (.Y (nx8877), .A0 (d_arr_mux_10__13), .A1 (nx11343), .B0 (
           d_arr_mul_10__13), .B1 (nx10495), .C0 (d_arr_add_10__13), .C1 (
           nx10687)) ;
    latch lat_d_arr_10__14 (.Q (d_arr_10__14), .D (nx4452), .CLK (nx10265)) ;
    inv01 ix4453 (.Y (nx4452), .A (nx8881)) ;
    aoi222 ix8882 (.Y (nx8881), .A0 (d_arr_mux_10__14), .A1 (nx11343), .B0 (
           d_arr_mul_10__14), .B1 (nx10497), .C0 (d_arr_add_10__14), .C1 (
           nx10689)) ;
    latch lat_d_arr_10__15 (.Q (d_arr_10__15), .D (nx4464), .CLK (nx10265)) ;
    inv01 ix4465 (.Y (nx4464), .A (nx8885)) ;
    aoi222 ix8886 (.Y (nx8885), .A0 (d_arr_mux_10__15), .A1 (nx11345), .B0 (
           d_arr_mul_10__15), .B1 (nx10497), .C0 (d_arr_add_10__15), .C1 (
           nx10689)) ;
    latch lat_d_arr_10__16 (.Q (d_arr_10__16), .D (nx4476), .CLK (nx10265)) ;
    inv01 ix4477 (.Y (nx4476), .A (nx8889)) ;
    aoi222 ix8890 (.Y (nx8889), .A0 (d_arr_mux_10__16), .A1 (nx11345), .B0 (
           d_arr_mul_10__16), .B1 (nx10497), .C0 (d_arr_add_10__16), .C1 (
           nx10689)) ;
    latch lat_d_arr_10__17 (.Q (d_arr_10__17), .D (nx4488), .CLK (nx10265)) ;
    inv01 ix4489 (.Y (nx4488), .A (nx8893)) ;
    aoi222 ix8894 (.Y (nx8893), .A0 (d_arr_mux_10__17), .A1 (nx11345), .B0 (
           d_arr_mul_10__17), .B1 (nx10497), .C0 (d_arr_add_10__17), .C1 (
           nx10689)) ;
    latch lat_d_arr_10__18 (.Q (d_arr_10__18), .D (nx4500), .CLK (nx10265)) ;
    inv01 ix4501 (.Y (nx4500), .A (nx8897)) ;
    aoi222 ix8898 (.Y (nx8897), .A0 (d_arr_mux_10__18), .A1 (nx11345), .B0 (
           d_arr_mul_10__18), .B1 (nx10497), .C0 (d_arr_add_10__18), .C1 (
           nx10689)) ;
    latch lat_d_arr_10__19 (.Q (d_arr_10__19), .D (nx4512), .CLK (nx10265)) ;
    inv01 ix4513 (.Y (nx4512), .A (nx8901)) ;
    aoi222 ix8902 (.Y (nx8901), .A0 (d_arr_mux_10__19), .A1 (nx11345), .B0 (
           d_arr_mul_10__19), .B1 (nx10497), .C0 (d_arr_add_10__19), .C1 (
           nx10689)) ;
    latch lat_d_arr_10__20 (.Q (d_arr_10__20), .D (nx4524), .CLK (nx10265)) ;
    inv01 ix4525 (.Y (nx4524), .A (nx8905)) ;
    aoi222 ix8906 (.Y (nx8905), .A0 (d_arr_mux_10__20), .A1 (nx11345), .B0 (
           d_arr_mul_10__20), .B1 (nx10497), .C0 (d_arr_add_10__20), .C1 (
           nx10689)) ;
    latch lat_d_arr_10__21 (.Q (d_arr_10__21), .D (nx4536), .CLK (nx10267)) ;
    inv01 ix4537 (.Y (nx4536), .A (nx8909)) ;
    aoi222 ix8910 (.Y (nx8909), .A0 (d_arr_mux_10__21), .A1 (nx11345), .B0 (
           d_arr_mul_10__21), .B1 (nx10499), .C0 (d_arr_add_10__21), .C1 (
           nx10691)) ;
    latch lat_d_arr_10__22 (.Q (d_arr_10__22), .D (nx4548), .CLK (nx10267)) ;
    inv01 ix4549 (.Y (nx4548), .A (nx8913)) ;
    aoi222 ix8914 (.Y (nx8913), .A0 (d_arr_mux_10__22), .A1 (nx11347), .B0 (
           d_arr_mul_10__22), .B1 (nx10499), .C0 (d_arr_add_10__22), .C1 (
           nx10691)) ;
    latch lat_d_arr_10__23 (.Q (d_arr_10__23), .D (nx4560), .CLK (nx10267)) ;
    inv01 ix4561 (.Y (nx4560), .A (nx8917)) ;
    aoi222 ix8918 (.Y (nx8917), .A0 (d_arr_mux_10__23), .A1 (nx11347), .B0 (
           d_arr_mul_10__23), .B1 (nx10499), .C0 (d_arr_add_10__23), .C1 (
           nx10691)) ;
    latch lat_d_arr_10__24 (.Q (d_arr_10__24), .D (nx4572), .CLK (nx10267)) ;
    inv01 ix4573 (.Y (nx4572), .A (nx8921)) ;
    aoi222 ix8922 (.Y (nx8921), .A0 (d_arr_mux_10__24), .A1 (nx11347), .B0 (
           d_arr_mul_10__24), .B1 (nx10499), .C0 (d_arr_add_10__24), .C1 (
           nx10691)) ;
    latch lat_d_arr_10__25 (.Q (d_arr_10__25), .D (nx4584), .CLK (nx10267)) ;
    inv01 ix4585 (.Y (nx4584), .A (nx8925)) ;
    aoi222 ix8926 (.Y (nx8925), .A0 (d_arr_mux_10__25), .A1 (nx11347), .B0 (
           d_arr_mul_10__25), .B1 (nx10499), .C0 (d_arr_add_10__25), .C1 (
           nx10691)) ;
    latch lat_d_arr_10__26 (.Q (d_arr_10__26), .D (nx4596), .CLK (nx10267)) ;
    inv01 ix4597 (.Y (nx4596), .A (nx8929)) ;
    aoi222 ix8930 (.Y (nx8929), .A0 (d_arr_mux_10__26), .A1 (nx11347), .B0 (
           d_arr_mul_10__26), .B1 (nx10499), .C0 (d_arr_add_10__26), .C1 (
           nx10691)) ;
    latch lat_d_arr_10__27 (.Q (d_arr_10__27), .D (nx4608), .CLK (nx10267)) ;
    inv01 ix4609 (.Y (nx4608), .A (nx8933)) ;
    aoi222 ix8934 (.Y (nx8933), .A0 (d_arr_mux_10__27), .A1 (nx11347), .B0 (
           d_arr_mul_10__27), .B1 (nx10499), .C0 (d_arr_add_10__27), .C1 (
           nx10691)) ;
    latch lat_d_arr_10__28 (.Q (d_arr_10__28), .D (nx4620), .CLK (nx10269)) ;
    inv01 ix4621 (.Y (nx4620), .A (nx8937)) ;
    aoi222 ix8938 (.Y (nx8937), .A0 (d_arr_mux_10__28), .A1 (nx11347), .B0 (
           d_arr_mul_10__28), .B1 (nx10501), .C0 (d_arr_add_10__28), .C1 (
           nx10693)) ;
    latch lat_d_arr_10__29 (.Q (d_arr_10__29), .D (nx4632), .CLK (nx10269)) ;
    inv01 ix4633 (.Y (nx4632), .A (nx8941)) ;
    aoi222 ix8942 (.Y (nx8941), .A0 (d_arr_mux_10__29), .A1 (nx11349), .B0 (
           d_arr_mul_10__29), .B1 (nx10501), .C0 (d_arr_add_10__29), .C1 (
           nx10693)) ;
    latch lat_d_arr_10__30 (.Q (d_arr_10__30), .D (nx4644), .CLK (nx10269)) ;
    inv01 ix4645 (.Y (nx4644), .A (nx8945)) ;
    aoi222 ix8946 (.Y (nx8945), .A0 (d_arr_mux_10__30), .A1 (nx11349), .B0 (
           d_arr_mul_10__30), .B1 (nx10501), .C0 (d_arr_add_10__30), .C1 (
           nx10693)) ;
    latch lat_d_arr_10__31 (.Q (d_arr_10__31), .D (nx4656), .CLK (nx10269)) ;
    inv01 ix4657 (.Y (nx4656), .A (nx8949)) ;
    aoi222 ix8950 (.Y (nx8949), .A0 (d_arr_mux_10__31), .A1 (nx11349), .B0 (
           d_arr_mul_10__31), .B1 (nx10501), .C0 (d_arr_add_10__31), .C1 (
           nx10693)) ;
    latch lat_d_arr_9__0 (.Q (d_arr_9__0), .D (nx4668), .CLK (nx10269)) ;
    inv01 ix4669 (.Y (nx4668), .A (nx8953)) ;
    aoi222 ix8954 (.Y (nx8953), .A0 (d_arr_mux_9__0), .A1 (nx11349), .B0 (
           d_arr_mul_9__0), .B1 (nx10501), .C0 (d_arr_add_9__0), .C1 (nx10693)
           ) ;
    latch lat_d_arr_9__1 (.Q (d_arr_9__1), .D (nx4680), .CLK (nx10269)) ;
    inv01 ix4681 (.Y (nx4680), .A (nx8957)) ;
    aoi222 ix8958 (.Y (nx8957), .A0 (d_arr_mux_9__1), .A1 (nx11349), .B0 (
           d_arr_mul_9__1), .B1 (nx10501), .C0 (d_arr_add_9__1), .C1 (nx10693)
           ) ;
    latch lat_d_arr_9__2 (.Q (d_arr_9__2), .D (nx4692), .CLK (nx10269)) ;
    inv01 ix4693 (.Y (nx4692), .A (nx8961)) ;
    aoi222 ix8962 (.Y (nx8961), .A0 (d_arr_mux_9__2), .A1 (nx11349), .B0 (
           d_arr_mul_9__2), .B1 (nx10501), .C0 (d_arr_add_9__2), .C1 (nx10693)
           ) ;
    latch lat_d_arr_9__3 (.Q (d_arr_9__3), .D (nx4704), .CLK (nx10271)) ;
    inv01 ix4705 (.Y (nx4704), .A (nx8965)) ;
    aoi222 ix8966 (.Y (nx8965), .A0 (d_arr_mux_9__3), .A1 (nx11349), .B0 (
           d_arr_mul_9__3), .B1 (nx10503), .C0 (d_arr_add_9__3), .C1 (nx10695)
           ) ;
    latch lat_d_arr_9__4 (.Q (d_arr_9__4), .D (nx4716), .CLK (nx10271)) ;
    inv01 ix4717 (.Y (nx4716), .A (nx8969)) ;
    aoi222 ix8970 (.Y (nx8969), .A0 (d_arr_mux_9__4), .A1 (nx11351), .B0 (
           d_arr_mul_9__4), .B1 (nx10503), .C0 (d_arr_add_9__4), .C1 (nx10695)
           ) ;
    latch lat_d_arr_9__5 (.Q (d_arr_9__5), .D (nx4728), .CLK (nx10271)) ;
    inv01 ix4729 (.Y (nx4728), .A (nx8973)) ;
    aoi222 ix8974 (.Y (nx8973), .A0 (d_arr_mux_9__5), .A1 (nx11351), .B0 (
           d_arr_mul_9__5), .B1 (nx10503), .C0 (d_arr_add_9__5), .C1 (nx10695)
           ) ;
    latch lat_d_arr_9__6 (.Q (d_arr_9__6), .D (nx4740), .CLK (nx10271)) ;
    inv01 ix4741 (.Y (nx4740), .A (nx8977)) ;
    aoi222 ix8978 (.Y (nx8977), .A0 (d_arr_mux_9__6), .A1 (nx11351), .B0 (
           d_arr_mul_9__6), .B1 (nx10503), .C0 (d_arr_add_9__6), .C1 (nx10695)
           ) ;
    latch lat_d_arr_9__7 (.Q (d_arr_9__7), .D (nx4752), .CLK (nx10271)) ;
    inv01 ix4753 (.Y (nx4752), .A (nx8981)) ;
    aoi222 ix8982 (.Y (nx8981), .A0 (d_arr_mux_9__7), .A1 (nx11351), .B0 (
           d_arr_mul_9__7), .B1 (nx10503), .C0 (d_arr_add_9__7), .C1 (nx10695)
           ) ;
    latch lat_d_arr_9__8 (.Q (d_arr_9__8), .D (nx4764), .CLK (nx10271)) ;
    inv01 ix4765 (.Y (nx4764), .A (nx8985)) ;
    aoi222 ix8986 (.Y (nx8985), .A0 (d_arr_mux_9__8), .A1 (nx11351), .B0 (
           d_arr_mul_9__8), .B1 (nx10503), .C0 (d_arr_add_9__8), .C1 (nx10695)
           ) ;
    latch lat_d_arr_9__9 (.Q (d_arr_9__9), .D (nx4776), .CLK (nx10271)) ;
    inv01 ix4777 (.Y (nx4776), .A (nx8989)) ;
    aoi222 ix8990 (.Y (nx8989), .A0 (d_arr_mux_9__9), .A1 (nx11351), .B0 (
           d_arr_mul_9__9), .B1 (nx10503), .C0 (d_arr_add_9__9), .C1 (nx10695)
           ) ;
    latch lat_d_arr_9__10 (.Q (d_arr_9__10), .D (nx4788), .CLK (nx10273)) ;
    inv01 ix4789 (.Y (nx4788), .A (nx8993)) ;
    aoi222 ix8994 (.Y (nx8993), .A0 (d_arr_mux_9__10), .A1 (nx11351), .B0 (
           d_arr_mul_9__10), .B1 (nx10505), .C0 (d_arr_add_9__10), .C1 (nx10697)
           ) ;
    latch lat_d_arr_9__11 (.Q (d_arr_9__11), .D (nx4800), .CLK (nx10273)) ;
    inv01 ix4801 (.Y (nx4800), .A (nx8997)) ;
    aoi222 ix8998 (.Y (nx8997), .A0 (d_arr_mux_9__11), .A1 (nx11353), .B0 (
           d_arr_mul_9__11), .B1 (nx10505), .C0 (d_arr_add_9__11), .C1 (nx10697)
           ) ;
    latch lat_d_arr_9__12 (.Q (d_arr_9__12), .D (nx4812), .CLK (nx10273)) ;
    inv01 ix4813 (.Y (nx4812), .A (nx9001)) ;
    aoi222 ix9002 (.Y (nx9001), .A0 (d_arr_mux_9__12), .A1 (nx11353), .B0 (
           d_arr_mul_9__12), .B1 (nx10505), .C0 (d_arr_add_9__12), .C1 (nx10697)
           ) ;
    latch lat_d_arr_9__13 (.Q (d_arr_9__13), .D (nx4824), .CLK (nx10273)) ;
    inv01 ix4825 (.Y (nx4824), .A (nx9005)) ;
    aoi222 ix9006 (.Y (nx9005), .A0 (d_arr_mux_9__13), .A1 (nx11353), .B0 (
           d_arr_mul_9__13), .B1 (nx10505), .C0 (d_arr_add_9__13), .C1 (nx10697)
           ) ;
    latch lat_d_arr_9__14 (.Q (d_arr_9__14), .D (nx4836), .CLK (nx10273)) ;
    inv01 ix4837 (.Y (nx4836), .A (nx9009)) ;
    aoi222 ix9010 (.Y (nx9009), .A0 (d_arr_mux_9__14), .A1 (nx11353), .B0 (
           d_arr_mul_9__14), .B1 (nx10505), .C0 (d_arr_add_9__14), .C1 (nx10697)
           ) ;
    latch lat_d_arr_9__15 (.Q (d_arr_9__15), .D (nx4848), .CLK (nx10273)) ;
    inv01 ix4849 (.Y (nx4848), .A (nx9013)) ;
    aoi222 ix9014 (.Y (nx9013), .A0 (d_arr_mux_9__15), .A1 (nx11353), .B0 (
           d_arr_mul_9__15), .B1 (nx10505), .C0 (d_arr_add_9__15), .C1 (nx10697)
           ) ;
    latch lat_d_arr_9__16 (.Q (d_arr_9__16), .D (nx4860), .CLK (nx10273)) ;
    inv01 ix4861 (.Y (nx4860), .A (nx9017)) ;
    aoi222 ix9018 (.Y (nx9017), .A0 (d_arr_mux_9__16), .A1 (nx11353), .B0 (
           d_arr_mul_9__16), .B1 (nx10505), .C0 (d_arr_add_9__16), .C1 (nx10697)
           ) ;
    latch lat_d_arr_9__17 (.Q (d_arr_9__17), .D (nx4872), .CLK (nx10275)) ;
    inv01 ix4873 (.Y (nx4872), .A (nx9021)) ;
    aoi222 ix9022 (.Y (nx9021), .A0 (d_arr_mux_9__17), .A1 (nx11353), .B0 (
           d_arr_mul_9__17), .B1 (nx10507), .C0 (d_arr_add_9__17), .C1 (nx10699)
           ) ;
    latch lat_d_arr_9__18 (.Q (d_arr_9__18), .D (nx4884), .CLK (nx10275)) ;
    inv01 ix4885 (.Y (nx4884), .A (nx9025)) ;
    aoi222 ix9026 (.Y (nx9025), .A0 (d_arr_mux_9__18), .A1 (nx11355), .B0 (
           d_arr_mul_9__18), .B1 (nx10507), .C0 (d_arr_add_9__18), .C1 (nx10699)
           ) ;
    latch lat_d_arr_9__19 (.Q (d_arr_9__19), .D (nx4896), .CLK (nx10275)) ;
    inv01 ix4897 (.Y (nx4896), .A (nx9029)) ;
    aoi222 ix9030 (.Y (nx9029), .A0 (d_arr_mux_9__19), .A1 (nx11355), .B0 (
           d_arr_mul_9__19), .B1 (nx10507), .C0 (d_arr_add_9__19), .C1 (nx10699)
           ) ;
    latch lat_d_arr_9__20 (.Q (d_arr_9__20), .D (nx4908), .CLK (nx10275)) ;
    inv01 ix4909 (.Y (nx4908), .A (nx9033)) ;
    aoi222 ix9034 (.Y (nx9033), .A0 (d_arr_mux_9__20), .A1 (nx11355), .B0 (
           d_arr_mul_9__20), .B1 (nx10507), .C0 (d_arr_add_9__20), .C1 (nx10699)
           ) ;
    latch lat_d_arr_9__21 (.Q (d_arr_9__21), .D (nx4920), .CLK (nx10275)) ;
    inv01 ix4921 (.Y (nx4920), .A (nx9037)) ;
    aoi222 ix9038 (.Y (nx9037), .A0 (d_arr_mux_9__21), .A1 (nx11355), .B0 (
           d_arr_mul_9__21), .B1 (nx10507), .C0 (d_arr_add_9__21), .C1 (nx10699)
           ) ;
    latch lat_d_arr_9__22 (.Q (d_arr_9__22), .D (nx4932), .CLK (nx10275)) ;
    inv01 ix4933 (.Y (nx4932), .A (nx9041)) ;
    aoi222 ix9042 (.Y (nx9041), .A0 (d_arr_mux_9__22), .A1 (nx11355), .B0 (
           d_arr_mul_9__22), .B1 (nx10507), .C0 (d_arr_add_9__22), .C1 (nx10699)
           ) ;
    latch lat_d_arr_9__23 (.Q (d_arr_9__23), .D (nx4944), .CLK (nx10275)) ;
    inv01 ix4945 (.Y (nx4944), .A (nx9045)) ;
    aoi222 ix9046 (.Y (nx9045), .A0 (d_arr_mux_9__23), .A1 (nx11355), .B0 (
           d_arr_mul_9__23), .B1 (nx10507), .C0 (d_arr_add_9__23), .C1 (nx10699)
           ) ;
    latch lat_d_arr_9__24 (.Q (d_arr_9__24), .D (nx4956), .CLK (nx10277)) ;
    inv01 ix4957 (.Y (nx4956), .A (nx9049)) ;
    aoi222 ix9050 (.Y (nx9049), .A0 (d_arr_mux_9__24), .A1 (nx11355), .B0 (
           d_arr_mul_9__24), .B1 (nx10509), .C0 (d_arr_add_9__24), .C1 (nx10701)
           ) ;
    latch lat_d_arr_9__25 (.Q (d_arr_9__25), .D (nx4968), .CLK (nx10277)) ;
    inv01 ix4969 (.Y (nx4968), .A (nx9053)) ;
    aoi222 ix9054 (.Y (nx9053), .A0 (d_arr_mux_9__25), .A1 (nx11357), .B0 (
           d_arr_mul_9__25), .B1 (nx10509), .C0 (d_arr_add_9__25), .C1 (nx10701)
           ) ;
    latch lat_d_arr_9__26 (.Q (d_arr_9__26), .D (nx4980), .CLK (nx10277)) ;
    inv01 ix4981 (.Y (nx4980), .A (nx9057)) ;
    aoi222 ix9058 (.Y (nx9057), .A0 (d_arr_mux_9__26), .A1 (nx11357), .B0 (
           d_arr_mul_9__26), .B1 (nx10509), .C0 (d_arr_add_9__26), .C1 (nx10701)
           ) ;
    latch lat_d_arr_9__27 (.Q (d_arr_9__27), .D (nx4992), .CLK (nx10277)) ;
    inv01 ix4993 (.Y (nx4992), .A (nx9061)) ;
    aoi222 ix9062 (.Y (nx9061), .A0 (d_arr_mux_9__27), .A1 (nx11357), .B0 (
           d_arr_mul_9__27), .B1 (nx10509), .C0 (d_arr_add_9__27), .C1 (nx10701)
           ) ;
    latch lat_d_arr_9__28 (.Q (d_arr_9__28), .D (nx5004), .CLK (nx10277)) ;
    inv01 ix5005 (.Y (nx5004), .A (nx9065)) ;
    aoi222 ix9066 (.Y (nx9065), .A0 (d_arr_mux_9__28), .A1 (nx11357), .B0 (
           d_arr_mul_9__28), .B1 (nx10509), .C0 (d_arr_add_9__28), .C1 (nx10701)
           ) ;
    latch lat_d_arr_9__29 (.Q (d_arr_9__29), .D (nx5016), .CLK (nx10277)) ;
    inv01 ix5017 (.Y (nx5016), .A (nx9069)) ;
    aoi222 ix9070 (.Y (nx9069), .A0 (d_arr_mux_9__29), .A1 (nx11357), .B0 (
           d_arr_mul_9__29), .B1 (nx10509), .C0 (d_arr_add_9__29), .C1 (nx10701)
           ) ;
    latch lat_d_arr_9__30 (.Q (d_arr_9__30), .D (nx5028), .CLK (nx10277)) ;
    inv01 ix5029 (.Y (nx5028), .A (nx9073)) ;
    aoi222 ix9074 (.Y (nx9073), .A0 (d_arr_mux_9__30), .A1 (nx11357), .B0 (
           d_arr_mul_9__30), .B1 (nx10509), .C0 (d_arr_add_9__30), .C1 (nx10701)
           ) ;
    latch lat_d_arr_9__31 (.Q (d_arr_9__31), .D (nx5040), .CLK (nx10279)) ;
    inv01 ix5041 (.Y (nx5040), .A (nx9077)) ;
    aoi222 ix9078 (.Y (nx9077), .A0 (d_arr_mux_9__31), .A1 (nx11357), .B0 (
           d_arr_mul_9__31), .B1 (nx10511), .C0 (d_arr_add_9__31), .C1 (nx10703)
           ) ;
    latch lat_d_arr_8__0 (.Q (d_arr_8__0), .D (nx5048), .CLK (nx10279)) ;
    ao22 ix5049 (.Y (nx5048), .A0 (d_arr_mux_8__0), .A1 (nx11359), .B0 (
         d_arr_mul_8__0), .B1 (nx10511)) ;
    latch lat_d_arr_8__1 (.Q (d_arr_8__1), .D (nx5056), .CLK (nx10279)) ;
    ao22 ix5057 (.Y (nx5056), .A0 (d_arr_mux_8__1), .A1 (nx11359), .B0 (
         d_arr_mul_8__1), .B1 (nx10511)) ;
    latch lat_d_arr_8__2 (.Q (d_arr_8__2), .D (nx5064), .CLK (nx10279)) ;
    ao22 ix5065 (.Y (nx5064), .A0 (d_arr_mux_8__2), .A1 (nx11359), .B0 (
         d_arr_mul_8__2), .B1 (nx10511)) ;
    latch lat_d_arr_8__3 (.Q (d_arr_8__3), .D (nx5072), .CLK (nx10279)) ;
    ao22 ix5073 (.Y (nx5072), .A0 (d_arr_mux_8__3), .A1 (nx11359), .B0 (
         d_arr_mul_8__3), .B1 (nx10511)) ;
    latch lat_d_arr_8__4 (.Q (d_arr_8__4), .D (nx5080), .CLK (nx10279)) ;
    ao22 ix5081 (.Y (nx5080), .A0 (d_arr_mux_8__4), .A1 (nx11359), .B0 (
         d_arr_mul_8__4), .B1 (nx10511)) ;
    latch lat_d_arr_8__5 (.Q (d_arr_8__5), .D (nx5088), .CLK (nx10279)) ;
    ao22 ix5089 (.Y (nx5088), .A0 (d_arr_mux_8__5), .A1 (nx11359), .B0 (
         d_arr_mul_8__5), .B1 (nx10511)) ;
    latch lat_d_arr_8__6 (.Q (d_arr_8__6), .D (nx5096), .CLK (nx10281)) ;
    ao22 ix5097 (.Y (nx5096), .A0 (d_arr_mux_8__6), .A1 (nx11359), .B0 (
         d_arr_mul_8__6), .B1 (nx10513)) ;
    latch lat_d_arr_8__7 (.Q (d_arr_8__7), .D (nx5104), .CLK (nx10281)) ;
    ao22 ix5105 (.Y (nx5104), .A0 (d_arr_mux_8__7), .A1 (nx11361), .B0 (
         d_arr_mul_8__7), .B1 (nx10513)) ;
    latch lat_d_arr_8__8 (.Q (d_arr_8__8), .D (nx5112), .CLK (nx10281)) ;
    ao22 ix5113 (.Y (nx5112), .A0 (d_arr_mux_8__8), .A1 (nx11361), .B0 (
         d_arr_mul_8__8), .B1 (nx10513)) ;
    latch lat_d_arr_8__9 (.Q (d_arr_8__9), .D (nx5120), .CLK (nx10281)) ;
    ao22 ix5121 (.Y (nx5120), .A0 (d_arr_mux_8__9), .A1 (nx11361), .B0 (
         d_arr_mul_8__9), .B1 (nx10513)) ;
    latch lat_d_arr_8__10 (.Q (d_arr_8__10), .D (nx5128), .CLK (nx10281)) ;
    ao22 ix5129 (.Y (nx5128), .A0 (d_arr_mux_8__10), .A1 (nx11361), .B0 (
         d_arr_mul_8__10), .B1 (nx10513)) ;
    latch lat_d_arr_8__11 (.Q (d_arr_8__11), .D (nx5136), .CLK (nx10281)) ;
    ao22 ix5137 (.Y (nx5136), .A0 (d_arr_mux_8__11), .A1 (nx11361), .B0 (
         d_arr_mul_8__11), .B1 (nx10513)) ;
    latch lat_d_arr_8__12 (.Q (d_arr_8__12), .D (nx5144), .CLK (nx10281)) ;
    ao22 ix5145 (.Y (nx5144), .A0 (d_arr_mux_8__12), .A1 (nx11361), .B0 (
         d_arr_mul_8__12), .B1 (nx10513)) ;
    latch lat_d_arr_8__13 (.Q (d_arr_8__13), .D (nx5152), .CLK (nx10283)) ;
    ao22 ix5153 (.Y (nx5152), .A0 (d_arr_mux_8__13), .A1 (nx11361), .B0 (
         d_arr_mul_8__13), .B1 (nx10515)) ;
    latch lat_d_arr_8__14 (.Q (d_arr_8__14), .D (nx5160), .CLK (nx10283)) ;
    ao22 ix5161 (.Y (nx5160), .A0 (d_arr_mux_8__14), .A1 (nx11363), .B0 (
         d_arr_mul_8__14), .B1 (nx10515)) ;
    latch lat_d_arr_8__15 (.Q (d_arr_8__15), .D (nx5168), .CLK (nx10283)) ;
    latch lat_d_arr_8__16 (.Q (d_arr_8__16), .D (nx5174), .CLK (nx10283)) ;
    latch lat_d_arr_8__17 (.Q (d_arr_8__17), .D (nx5180), .CLK (nx10283)) ;
    latch lat_d_arr_8__18 (.Q (d_arr_8__18), .D (nx5186), .CLK (nx10283)) ;
    latch lat_d_arr_8__19 (.Q (d_arr_8__19), .D (nx5192), .CLK (nx10283)) ;
    latch lat_d_arr_8__20 (.Q (d_arr_8__20), .D (nx5198), .CLK (nx10285)) ;
    latch lat_d_arr_8__21 (.Q (d_arr_8__21), .D (nx5204), .CLK (nx10285)) ;
    latch lat_d_arr_8__22 (.Q (d_arr_8__22), .D (nx5210), .CLK (nx10285)) ;
    latch lat_d_arr_8__23 (.Q (d_arr_8__23), .D (nx5216), .CLK (nx10285)) ;
    latch lat_d_arr_8__24 (.Q (d_arr_8__24), .D (nx5222), .CLK (nx10285)) ;
    latch lat_d_arr_8__25 (.Q (d_arr_8__25), .D (nx5228), .CLK (nx10285)) ;
    latch lat_d_arr_8__26 (.Q (d_arr_8__26), .D (nx5234), .CLK (nx10285)) ;
    latch lat_d_arr_8__27 (.Q (d_arr_8__27), .D (nx5240), .CLK (nx10287)) ;
    latch lat_d_arr_8__28 (.Q (d_arr_8__28), .D (nx5246), .CLK (nx10287)) ;
    latch lat_d_arr_8__29 (.Q (d_arr_8__29), .D (nx5252), .CLK (nx10287)) ;
    latch lat_d_arr_8__30 (.Q (d_arr_8__30), .D (nx5258), .CLK (nx10287)) ;
    latch lat_d_arr_8__31 (.Q (d_arr_8__31), .D (nx5264), .CLK (nx10287)) ;
    latch lat_d_arr_7__0 (.Q (d_arr_7__0), .D (nx5272), .CLK (nx10287)) ;
    ao22 ix5273 (.Y (nx5272), .A0 (d_arr_mux_7__0), .A1 (nx11363), .B0 (
         d_arr_mul_7__0), .B1 (nx10519)) ;
    latch lat_d_arr_7__1 (.Q (d_arr_7__1), .D (nx5280), .CLK (nx10287)) ;
    ao22 ix5281 (.Y (nx5280), .A0 (d_arr_mux_7__1), .A1 (nx11363), .B0 (
         d_arr_mul_7__1), .B1 (nx10519)) ;
    latch lat_d_arr_7__2 (.Q (d_arr_7__2), .D (nx5288), .CLK (nx10289)) ;
    ao22 ix5289 (.Y (nx5288), .A0 (d_arr_mux_7__2), .A1 (nx11363), .B0 (
         d_arr_mul_7__2), .B1 (nx10521)) ;
    latch lat_d_arr_7__3 (.Q (d_arr_7__3), .D (nx5296), .CLK (nx10289)) ;
    ao22 ix5297 (.Y (nx5296), .A0 (d_arr_mux_7__3), .A1 (nx11363), .B0 (
         d_arr_mul_7__3), .B1 (nx10521)) ;
    latch lat_d_arr_7__4 (.Q (d_arr_7__4), .D (nx5304), .CLK (nx10289)) ;
    ao22 ix5305 (.Y (nx5304), .A0 (d_arr_mux_7__4), .A1 (nx11363), .B0 (
         d_arr_mul_7__4), .B1 (nx10521)) ;
    latch lat_d_arr_7__5 (.Q (d_arr_7__5), .D (nx5312), .CLK (nx10289)) ;
    ao22 ix5313 (.Y (nx5312), .A0 (d_arr_mux_7__5), .A1 (nx11363), .B0 (
         d_arr_mul_7__5), .B1 (nx10521)) ;
    latch lat_d_arr_7__6 (.Q (d_arr_7__6), .D (nx5320), .CLK (nx10289)) ;
    ao22 ix5321 (.Y (nx5320), .A0 (d_arr_mux_7__6), .A1 (nx11365), .B0 (
         d_arr_mul_7__6), .B1 (nx10521)) ;
    latch lat_d_arr_7__7 (.Q (d_arr_7__7), .D (nx5328), .CLK (nx10289)) ;
    ao22 ix5329 (.Y (nx5328), .A0 (d_arr_mux_7__7), .A1 (nx11365), .B0 (
         d_arr_mul_7__7), .B1 (nx10521)) ;
    latch lat_d_arr_7__8 (.Q (d_arr_7__8), .D (nx5336), .CLK (nx10289)) ;
    ao22 ix5337 (.Y (nx5336), .A0 (d_arr_mux_7__8), .A1 (nx11365), .B0 (
         d_arr_mul_7__8), .B1 (nx10521)) ;
    latch lat_d_arr_7__9 (.Q (d_arr_7__9), .D (nx5344), .CLK (nx10291)) ;
    ao22 ix5345 (.Y (nx5344), .A0 (d_arr_mux_7__9), .A1 (nx11365), .B0 (
         d_arr_mul_7__9), .B1 (nx10523)) ;
    latch lat_d_arr_7__10 (.Q (d_arr_7__10), .D (nx5352), .CLK (nx10291)) ;
    ao22 ix5353 (.Y (nx5352), .A0 (d_arr_mux_7__10), .A1 (nx11365), .B0 (
         d_arr_mul_7__10), .B1 (nx10523)) ;
    latch lat_d_arr_7__11 (.Q (d_arr_7__11), .D (nx5360), .CLK (nx10291)) ;
    ao22 ix5361 (.Y (nx5360), .A0 (d_arr_mux_7__11), .A1 (nx11365), .B0 (
         d_arr_mul_7__11), .B1 (nx10523)) ;
    latch lat_d_arr_7__12 (.Q (d_arr_7__12), .D (nx5368), .CLK (nx10291)) ;
    ao22 ix5369 (.Y (nx5368), .A0 (d_arr_mux_7__12), .A1 (nx11365), .B0 (
         d_arr_mul_7__12), .B1 (nx10523)) ;
    latch lat_d_arr_7__13 (.Q (d_arr_7__13), .D (nx5376), .CLK (nx10291)) ;
    ao22 ix5377 (.Y (nx5376), .A0 (d_arr_mux_7__13), .A1 (nx11367), .B0 (
         d_arr_mul_7__13), .B1 (nx10523)) ;
    latch lat_d_arr_7__14 (.Q (d_arr_7__14), .D (nx5384), .CLK (nx10291)) ;
    ao22 ix5385 (.Y (nx5384), .A0 (d_arr_mux_7__14), .A1 (nx11367), .B0 (
         d_arr_mul_7__14), .B1 (nx10523)) ;
    latch lat_d_arr_7__15 (.Q (d_arr_7__15), .D (nx5392), .CLK (nx10291)) ;
    latch lat_d_arr_7__16 (.Q (d_arr_7__16), .D (nx5398), .CLK (nx10293)) ;
    latch lat_d_arr_7__17 (.Q (d_arr_7__17), .D (nx5404), .CLK (nx10293)) ;
    latch lat_d_arr_7__18 (.Q (d_arr_7__18), .D (nx5410), .CLK (nx10293)) ;
    latch lat_d_arr_7__19 (.Q (d_arr_7__19), .D (nx5416), .CLK (nx10293)) ;
    latch lat_d_arr_7__20 (.Q (d_arr_7__20), .D (nx5422), .CLK (nx10293)) ;
    latch lat_d_arr_7__21 (.Q (d_arr_7__21), .D (nx5428), .CLK (nx10293)) ;
    latch lat_d_arr_7__22 (.Q (d_arr_7__22), .D (nx5434), .CLK (nx10293)) ;
    latch lat_d_arr_7__23 (.Q (d_arr_7__23), .D (nx5440), .CLK (nx10295)) ;
    latch lat_d_arr_7__24 (.Q (d_arr_7__24), .D (nx5446), .CLK (nx10295)) ;
    latch lat_d_arr_7__25 (.Q (d_arr_7__25), .D (nx5452), .CLK (nx10295)) ;
    latch lat_d_arr_7__26 (.Q (d_arr_7__26), .D (nx5458), .CLK (nx10295)) ;
    latch lat_d_arr_7__27 (.Q (d_arr_7__27), .D (nx5464), .CLK (nx10295)) ;
    latch lat_d_arr_7__28 (.Q (d_arr_7__28), .D (nx5470), .CLK (nx10295)) ;
    latch lat_d_arr_7__29 (.Q (d_arr_7__29), .D (nx5476), .CLK (nx10295)) ;
    latch lat_d_arr_7__30 (.Q (d_arr_7__30), .D (nx5482), .CLK (nx10297)) ;
    latch lat_d_arr_7__31 (.Q (d_arr_7__31), .D (nx5488), .CLK (nx10297)) ;
    latch lat_d_arr_6__0 (.Q (d_arr_6__0), .D (nx5496), .CLK (nx10297)) ;
    ao22 ix5497 (.Y (nx5496), .A0 (d_arr_mux_6__0), .A1 (nx11367), .B0 (
         d_arr_mul_6__0), .B1 (nx10529)) ;
    latch lat_d_arr_6__1 (.Q (d_arr_6__1), .D (nx5504), .CLK (nx10297)) ;
    ao22 ix5505 (.Y (nx5504), .A0 (d_arr_mux_6__1), .A1 (nx11367), .B0 (
         d_arr_mul_6__1), .B1 (nx10529)) ;
    latch lat_d_arr_6__2 (.Q (d_arr_6__2), .D (nx5512), .CLK (nx10297)) ;
    ao22 ix5513 (.Y (nx5512), .A0 (d_arr_mux_6__2), .A1 (nx11367), .B0 (
         d_arr_mul_6__2), .B1 (nx10529)) ;
    latch lat_d_arr_6__3 (.Q (d_arr_6__3), .D (nx5520), .CLK (nx10297)) ;
    ao22 ix5521 (.Y (nx5520), .A0 (d_arr_mux_6__3), .A1 (nx11367), .B0 (
         d_arr_mul_6__3), .B1 (nx10529)) ;
    latch lat_d_arr_6__4 (.Q (d_arr_6__4), .D (nx5528), .CLK (nx10297)) ;
    ao22 ix5529 (.Y (nx5528), .A0 (d_arr_mux_6__4), .A1 (nx11367), .B0 (
         d_arr_mul_6__4), .B1 (nx10529)) ;
    latch lat_d_arr_6__5 (.Q (d_arr_6__5), .D (nx5536), .CLK (nx10299)) ;
    ao22 ix5537 (.Y (nx5536), .A0 (d_arr_mux_6__5), .A1 (nx11369), .B0 (
         d_arr_mul_6__5), .B1 (nx10531)) ;
    latch lat_d_arr_6__6 (.Q (d_arr_6__6), .D (nx5544), .CLK (nx10299)) ;
    ao22 ix5545 (.Y (nx5544), .A0 (d_arr_mux_6__6), .A1 (nx11369), .B0 (
         d_arr_mul_6__6), .B1 (nx10531)) ;
    latch lat_d_arr_6__7 (.Q (d_arr_6__7), .D (nx5552), .CLK (nx10299)) ;
    ao22 ix5553 (.Y (nx5552), .A0 (d_arr_mux_6__7), .A1 (nx11369), .B0 (
         d_arr_mul_6__7), .B1 (nx10531)) ;
    latch lat_d_arr_6__8 (.Q (d_arr_6__8), .D (nx5560), .CLK (nx10299)) ;
    ao22 ix5561 (.Y (nx5560), .A0 (d_arr_mux_6__8), .A1 (nx11369), .B0 (
         d_arr_mul_6__8), .B1 (nx10531)) ;
    latch lat_d_arr_6__9 (.Q (d_arr_6__9), .D (nx5568), .CLK (nx10299)) ;
    ao22 ix5569 (.Y (nx5568), .A0 (d_arr_mux_6__9), .A1 (nx11369), .B0 (
         d_arr_mul_6__9), .B1 (nx10531)) ;
    latch lat_d_arr_6__10 (.Q (d_arr_6__10), .D (nx5576), .CLK (nx10299)) ;
    ao22 ix5577 (.Y (nx5576), .A0 (d_arr_mux_6__10), .A1 (nx11369), .B0 (
         d_arr_mul_6__10), .B1 (nx10531)) ;
    latch lat_d_arr_6__11 (.Q (d_arr_6__11), .D (nx5584), .CLK (nx10299)) ;
    ao22 ix5585 (.Y (nx5584), .A0 (d_arr_mux_6__11), .A1 (nx11369), .B0 (
         d_arr_mul_6__11), .B1 (nx10531)) ;
    latch lat_d_arr_6__12 (.Q (d_arr_6__12), .D (nx5592), .CLK (nx10301)) ;
    ao22 ix5593 (.Y (nx5592), .A0 (d_arr_mux_6__12), .A1 (nx11371), .B0 (
         d_arr_mul_6__12), .B1 (nx10533)) ;
    latch lat_d_arr_6__13 (.Q (d_arr_6__13), .D (nx5600), .CLK (nx10301)) ;
    ao22 ix5601 (.Y (nx5600), .A0 (d_arr_mux_6__13), .A1 (nx11371), .B0 (
         d_arr_mul_6__13), .B1 (nx10533)) ;
    latch lat_d_arr_6__14 (.Q (d_arr_6__14), .D (nx5608), .CLK (nx10301)) ;
    ao22 ix5609 (.Y (nx5608), .A0 (d_arr_mux_6__14), .A1 (nx11371), .B0 (
         d_arr_mul_6__14), .B1 (nx10533)) ;
    latch lat_d_arr_6__15 (.Q (d_arr_6__15), .D (nx5616), .CLK (nx10301)) ;
    latch lat_d_arr_6__16 (.Q (d_arr_6__16), .D (nx5622), .CLK (nx10301)) ;
    latch lat_d_arr_6__17 (.Q (d_arr_6__17), .D (nx5628), .CLK (nx10301)) ;
    latch lat_d_arr_6__18 (.Q (d_arr_6__18), .D (nx5634), .CLK (nx10301)) ;
    latch lat_d_arr_6__19 (.Q (d_arr_6__19), .D (nx5640), .CLK (nx10303)) ;
    latch lat_d_arr_6__20 (.Q (d_arr_6__20), .D (nx5646), .CLK (nx10303)) ;
    latch lat_d_arr_6__21 (.Q (d_arr_6__21), .D (nx5652), .CLK (nx10303)) ;
    latch lat_d_arr_6__22 (.Q (d_arr_6__22), .D (nx5658), .CLK (nx10303)) ;
    latch lat_d_arr_6__23 (.Q (d_arr_6__23), .D (nx5664), .CLK (nx10303)) ;
    latch lat_d_arr_6__24 (.Q (d_arr_6__24), .D (nx5670), .CLK (nx10303)) ;
    latch lat_d_arr_6__25 (.Q (d_arr_6__25), .D (nx5676), .CLK (nx10303)) ;
    latch lat_d_arr_6__26 (.Q (d_arr_6__26), .D (nx5682), .CLK (nx10305)) ;
    latch lat_d_arr_6__27 (.Q (d_arr_6__27), .D (nx5688), .CLK (nx10305)) ;
    latch lat_d_arr_6__28 (.Q (d_arr_6__28), .D (nx5694), .CLK (nx10305)) ;
    latch lat_d_arr_6__29 (.Q (d_arr_6__29), .D (nx5700), .CLK (nx10305)) ;
    latch lat_d_arr_6__30 (.Q (d_arr_6__30), .D (nx5706), .CLK (nx10305)) ;
    latch lat_d_arr_6__31 (.Q (d_arr_6__31), .D (nx5712), .CLK (nx10305)) ;
    latch lat_d_arr_5__0 (.Q (d_arr_5__0), .D (nx5720), .CLK (nx10305)) ;
    ao22 ix5721 (.Y (nx5720), .A0 (d_arr_mux_5__0), .A1 (nx11371), .B0 (
         d_arr_mul_5__0), .B1 (nx10537)) ;
    latch lat_d_arr_5__1 (.Q (d_arr_5__1), .D (nx5728), .CLK (nx10307)) ;
    ao22 ix5729 (.Y (nx5728), .A0 (d_arr_mux_5__1), .A1 (nx11371), .B0 (
         d_arr_mul_5__1), .B1 (nx10539)) ;
    latch lat_d_arr_5__2 (.Q (d_arr_5__2), .D (nx5736), .CLK (nx10307)) ;
    ao22 ix5737 (.Y (nx5736), .A0 (d_arr_mux_5__2), .A1 (nx11371), .B0 (
         d_arr_mul_5__2), .B1 (nx10539)) ;
    latch lat_d_arr_5__3 (.Q (d_arr_5__3), .D (nx5744), .CLK (nx10307)) ;
    ao22 ix5745 (.Y (nx5744), .A0 (d_arr_mux_5__3), .A1 (nx11371), .B0 (
         d_arr_mul_5__3), .B1 (nx10539)) ;
    latch lat_d_arr_5__4 (.Q (d_arr_5__4), .D (nx5752), .CLK (nx10307)) ;
    ao22 ix5753 (.Y (nx5752), .A0 (d_arr_mux_5__4), .A1 (nx11373), .B0 (
         d_arr_mul_5__4), .B1 (nx10539)) ;
    latch lat_d_arr_5__5 (.Q (d_arr_5__5), .D (nx5760), .CLK (nx10307)) ;
    ao22 ix5761 (.Y (nx5760), .A0 (d_arr_mux_5__5), .A1 (nx11373), .B0 (
         d_arr_mul_5__5), .B1 (nx10539)) ;
    latch lat_d_arr_5__6 (.Q (d_arr_5__6), .D (nx5768), .CLK (nx10307)) ;
    ao22 ix5769 (.Y (nx5768), .A0 (d_arr_mux_5__6), .A1 (nx11373), .B0 (
         d_arr_mul_5__6), .B1 (nx10539)) ;
    latch lat_d_arr_5__7 (.Q (d_arr_5__7), .D (nx5776), .CLK (nx10307)) ;
    ao22 ix5777 (.Y (nx5776), .A0 (d_arr_mux_5__7), .A1 (nx11373), .B0 (
         d_arr_mul_5__7), .B1 (nx10539)) ;
    latch lat_d_arr_5__8 (.Q (d_arr_5__8), .D (nx5784), .CLK (nx10309)) ;
    ao22 ix5785 (.Y (nx5784), .A0 (d_arr_mux_5__8), .A1 (nx11373), .B0 (
         d_arr_mul_5__8), .B1 (nx10541)) ;
    latch lat_d_arr_5__9 (.Q (d_arr_5__9), .D (nx5792), .CLK (nx10309)) ;
    ao22 ix5793 (.Y (nx5792), .A0 (d_arr_mux_5__9), .A1 (nx11373), .B0 (
         d_arr_mul_5__9), .B1 (nx10541)) ;
    latch lat_d_arr_5__10 (.Q (d_arr_5__10), .D (nx5800), .CLK (nx10309)) ;
    ao22 ix5801 (.Y (nx5800), .A0 (d_arr_mux_5__10), .A1 (nx11373), .B0 (
         d_arr_mul_5__10), .B1 (nx10541)) ;
    latch lat_d_arr_5__11 (.Q (d_arr_5__11), .D (nx5808), .CLK (nx10309)) ;
    ao22 ix5809 (.Y (nx5808), .A0 (d_arr_mux_5__11), .A1 (nx11375), .B0 (
         d_arr_mul_5__11), .B1 (nx10541)) ;
    latch lat_d_arr_5__12 (.Q (d_arr_5__12), .D (nx5816), .CLK (nx10309)) ;
    ao22 ix5817 (.Y (nx5816), .A0 (d_arr_mux_5__12), .A1 (nx11375), .B0 (
         d_arr_mul_5__12), .B1 (nx10541)) ;
    latch lat_d_arr_5__13 (.Q (d_arr_5__13), .D (nx5824), .CLK (nx10309)) ;
    ao22 ix5825 (.Y (nx5824), .A0 (d_arr_mux_5__13), .A1 (nx11375), .B0 (
         d_arr_mul_5__13), .B1 (nx10541)) ;
    latch lat_d_arr_5__14 (.Q (d_arr_5__14), .D (nx5832), .CLK (nx10309)) ;
    ao22 ix5833 (.Y (nx5832), .A0 (d_arr_mux_5__14), .A1 (nx11375), .B0 (
         d_arr_mul_5__14), .B1 (nx10541)) ;
    latch lat_d_arr_5__15 (.Q (d_arr_5__15), .D (nx5840), .CLK (nx10311)) ;
    latch lat_d_arr_5__16 (.Q (d_arr_5__16), .D (nx5846), .CLK (nx10311)) ;
    latch lat_d_arr_5__17 (.Q (d_arr_5__17), .D (nx5852), .CLK (nx10311)) ;
    latch lat_d_arr_5__18 (.Q (d_arr_5__18), .D (nx5858), .CLK (nx10311)) ;
    latch lat_d_arr_5__19 (.Q (d_arr_5__19), .D (nx5864), .CLK (nx10311)) ;
    latch lat_d_arr_5__20 (.Q (d_arr_5__20), .D (nx5870), .CLK (nx10311)) ;
    latch lat_d_arr_5__21 (.Q (d_arr_5__21), .D (nx5876), .CLK (nx10311)) ;
    latch lat_d_arr_5__22 (.Q (d_arr_5__22), .D (nx5882), .CLK (nx10313)) ;
    latch lat_d_arr_5__23 (.Q (d_arr_5__23), .D (nx5888), .CLK (nx10313)) ;
    latch lat_d_arr_5__24 (.Q (d_arr_5__24), .D (nx5894), .CLK (nx10313)) ;
    latch lat_d_arr_5__25 (.Q (d_arr_5__25), .D (nx5900), .CLK (nx10313)) ;
    latch lat_d_arr_5__26 (.Q (d_arr_5__26), .D (nx5906), .CLK (nx10313)) ;
    latch lat_d_arr_5__27 (.Q (d_arr_5__27), .D (nx5912), .CLK (nx10313)) ;
    latch lat_d_arr_5__28 (.Q (d_arr_5__28), .D (nx5918), .CLK (nx10313)) ;
    latch lat_d_arr_5__29 (.Q (d_arr_5__29), .D (nx5924), .CLK (nx10315)) ;
    latch lat_d_arr_5__30 (.Q (d_arr_5__30), .D (nx5930), .CLK (nx10315)) ;
    latch lat_d_arr_5__31 (.Q (d_arr_5__31), .D (nx5936), .CLK (nx10315)) ;
    latch lat_d_arr_4__0 (.Q (d_arr_4__0), .D (nx5948), .CLK (nx10315)) ;
    inv01 ix5949 (.Y (nx5948), .A (nx9341)) ;
    aoi222 ix9342 (.Y (nx9341), .A0 (d_arr_mux_4__0), .A1 (nx11375), .B0 (
           d_arr_mul_4__0), .B1 (nx10547), .C0 (d_arr_add_4__0), .C1 (nx10703)
           ) ;
    latch lat_d_arr_4__1 (.Q (d_arr_4__1), .D (nx5960), .CLK (nx10315)) ;
    inv01 ix5961 (.Y (nx5960), .A (nx9345)) ;
    aoi222 ix9346 (.Y (nx9345), .A0 (d_arr_mux_4__1), .A1 (nx11375), .B0 (
           d_arr_mul_4__1), .B1 (nx10547), .C0 (d_arr_add_4__1), .C1 (nx10703)
           ) ;
    latch lat_d_arr_4__2 (.Q (d_arr_4__2), .D (nx5972), .CLK (nx10315)) ;
    inv01 ix5973 (.Y (nx5972), .A (nx9349)) ;
    aoi222 ix9350 (.Y (nx9349), .A0 (d_arr_mux_4__2), .A1 (nx11375), .B0 (
           d_arr_mul_4__2), .B1 (nx10547), .C0 (d_arr_add_4__2), .C1 (nx10703)
           ) ;
    latch lat_d_arr_4__3 (.Q (d_arr_4__3), .D (nx5984), .CLK (nx10315)) ;
    inv01 ix5985 (.Y (nx5984), .A (nx9353)) ;
    aoi222 ix9354 (.Y (nx9353), .A0 (d_arr_mux_4__3), .A1 (nx11377), .B0 (
           d_arr_mul_4__3), .B1 (nx10547), .C0 (d_arr_add_4__3), .C1 (nx10703)
           ) ;
    latch lat_d_arr_4__4 (.Q (d_arr_4__4), .D (nx5996), .CLK (nx10317)) ;
    inv01 ix5997 (.Y (nx5996), .A (nx9357)) ;
    aoi222 ix9358 (.Y (nx9357), .A0 (d_arr_mux_4__4), .A1 (nx11377), .B0 (
           d_arr_mul_4__4), .B1 (nx10549), .C0 (d_arr_add_4__4), .C1 (nx10703)
           ) ;
    latch lat_d_arr_4__5 (.Q (d_arr_4__5), .D (nx6008), .CLK (nx10317)) ;
    inv01 ix6009 (.Y (nx6008), .A (nx9361)) ;
    aoi222 ix9362 (.Y (nx9361), .A0 (d_arr_mux_4__5), .A1 (nx11377), .B0 (
           d_arr_mul_4__5), .B1 (nx10549), .C0 (d_arr_add_4__5), .C1 (nx10703)
           ) ;
    latch lat_d_arr_4__6 (.Q (d_arr_4__6), .D (nx6020), .CLK (nx10317)) ;
    inv01 ix6021 (.Y (nx6020), .A (nx9365)) ;
    aoi222 ix9366 (.Y (nx9365), .A0 (d_arr_mux_4__6), .A1 (nx11377), .B0 (
           d_arr_mul_4__6), .B1 (nx10549), .C0 (d_arr_add_4__6), .C1 (nx10705)
           ) ;
    latch lat_d_arr_4__7 (.Q (d_arr_4__7), .D (nx6032), .CLK (nx10317)) ;
    inv01 ix6033 (.Y (nx6032), .A (nx9369)) ;
    aoi222 ix9370 (.Y (nx9369), .A0 (d_arr_mux_4__7), .A1 (nx11377), .B0 (
           d_arr_mul_4__7), .B1 (nx10549), .C0 (d_arr_add_4__7), .C1 (nx10705)
           ) ;
    latch lat_d_arr_4__8 (.Q (d_arr_4__8), .D (nx6044), .CLK (nx10317)) ;
    inv01 ix6045 (.Y (nx6044), .A (nx9373)) ;
    aoi222 ix9374 (.Y (nx9373), .A0 (d_arr_mux_4__8), .A1 (nx11377), .B0 (
           d_arr_mul_4__8), .B1 (nx10549), .C0 (d_arr_add_4__8), .C1 (nx10705)
           ) ;
    latch lat_d_arr_4__9 (.Q (d_arr_4__9), .D (nx6056), .CLK (nx10317)) ;
    inv01 ix6057 (.Y (nx6056), .A (nx9377)) ;
    aoi222 ix9378 (.Y (nx9377), .A0 (d_arr_mux_4__9), .A1 (nx11377), .B0 (
           d_arr_mul_4__9), .B1 (nx10549), .C0 (d_arr_add_4__9), .C1 (nx10705)
           ) ;
    latch lat_d_arr_4__10 (.Q (d_arr_4__10), .D (nx6068), .CLK (nx10317)) ;
    inv01 ix6069 (.Y (nx6068), .A (nx9381)) ;
    aoi222 ix9382 (.Y (nx9381), .A0 (d_arr_mux_4__10), .A1 (nx11379), .B0 (
           d_arr_mul_4__10), .B1 (nx10549), .C0 (d_arr_add_4__10), .C1 (nx10705)
           ) ;
    latch lat_d_arr_4__11 (.Q (d_arr_4__11), .D (nx6080), .CLK (nx10319)) ;
    inv01 ix6081 (.Y (nx6080), .A (nx9385)) ;
    aoi222 ix9386 (.Y (nx9385), .A0 (d_arr_mux_4__11), .A1 (nx11379), .B0 (
           d_arr_mul_4__11), .B1 (nx10551), .C0 (d_arr_add_4__11), .C1 (nx10705)
           ) ;
    latch lat_d_arr_4__12 (.Q (d_arr_4__12), .D (nx6092), .CLK (nx10319)) ;
    inv01 ix6093 (.Y (nx6092), .A (nx9389)) ;
    aoi222 ix9390 (.Y (nx9389), .A0 (d_arr_mux_4__12), .A1 (nx11379), .B0 (
           d_arr_mul_4__12), .B1 (nx10551), .C0 (d_arr_add_4__12), .C1 (nx10705)
           ) ;
    latch lat_d_arr_4__13 (.Q (d_arr_4__13), .D (nx6104), .CLK (nx10319)) ;
    inv01 ix6105 (.Y (nx6104), .A (nx9393)) ;
    aoi222 ix9394 (.Y (nx9393), .A0 (d_arr_mux_4__13), .A1 (nx11379), .B0 (
           d_arr_mul_4__13), .B1 (nx10551), .C0 (d_arr_add_4__13), .C1 (nx10707)
           ) ;
    latch lat_d_arr_4__14 (.Q (d_arr_4__14), .D (nx6116), .CLK (nx10319)) ;
    inv01 ix6117 (.Y (nx6116), .A (nx9397)) ;
    aoi222 ix9398 (.Y (nx9397), .A0 (d_arr_mux_4__14), .A1 (nx11379), .B0 (
           d_arr_mul_4__14), .B1 (nx10551), .C0 (d_arr_add_4__14), .C1 (nx10707)
           ) ;
    latch lat_d_arr_4__15 (.Q (d_arr_4__15), .D (nx6128), .CLK (nx10319)) ;
    nand02 ix6129 (.Y (nx6128), .A0 (nx9401), .A1 (nx10861)) ;
    aoi22 ix9402 (.Y (nx9401), .A0 (d_arr_mul_4__15), .A1 (nx10551), .B0 (
          d_arr_add_4__15), .B1 (nx10707)) ;
    nand02 ix9404 (.Y (nx9403), .A0 (d_arr_mux_4__31), .A1 (nx11379)) ;
    latch lat_d_arr_4__16 (.Q (d_arr_4__16), .D (nx6138), .CLK (nx10319)) ;
    nand02 ix6139 (.Y (nx6138), .A0 (nx9407), .A1 (nx10861)) ;
    aoi22 ix9408 (.Y (nx9407), .A0 (d_arr_mul_4__16), .A1 (nx10551), .B0 (
          d_arr_add_4__16), .B1 (nx10707)) ;
    latch lat_d_arr_4__17 (.Q (d_arr_4__17), .D (nx6148), .CLK (nx10319)) ;
    nand02 ix6149 (.Y (nx6148), .A0 (nx9411), .A1 (nx10861)) ;
    aoi22 ix9412 (.Y (nx9411), .A0 (d_arr_mul_4__17), .A1 (nx10551), .B0 (
          d_arr_add_4__17), .B1 (nx10707)) ;
    latch lat_d_arr_4__18 (.Q (d_arr_4__18), .D (nx6158), .CLK (nx10321)) ;
    nand02 ix6159 (.Y (nx6158), .A0 (nx9415), .A1 (nx10861)) ;
    aoi22 ix9416 (.Y (nx9415), .A0 (d_arr_mul_4__18), .A1 (nx10553), .B0 (
          d_arr_add_4__18), .B1 (nx10707)) ;
    latch lat_d_arr_4__19 (.Q (d_arr_4__19), .D (nx6168), .CLK (nx10321)) ;
    nand02 ix6169 (.Y (nx6168), .A0 (nx9419), .A1 (nx10861)) ;
    aoi22 ix9420 (.Y (nx9419), .A0 (d_arr_mul_4__19), .A1 (nx10553), .B0 (
          d_arr_add_4__19), .B1 (nx10707)) ;
    latch lat_d_arr_4__20 (.Q (d_arr_4__20), .D (nx6178), .CLK (nx10321)) ;
    nand02 ix6179 (.Y (nx6178), .A0 (nx9423), .A1 (nx10861)) ;
    aoi22 ix9424 (.Y (nx9423), .A0 (d_arr_mul_4__20), .A1 (nx10553), .B0 (
          d_arr_add_4__20), .B1 (nx10709)) ;
    latch lat_d_arr_4__21 (.Q (d_arr_4__21), .D (nx6188), .CLK (nx10321)) ;
    nand02 ix6189 (.Y (nx6188), .A0 (nx9427), .A1 (nx10861)) ;
    aoi22 ix9428 (.Y (nx9427), .A0 (d_arr_mul_4__21), .A1 (nx10553), .B0 (
          d_arr_add_4__21), .B1 (nx10709)) ;
    latch lat_d_arr_4__22 (.Q (d_arr_4__22), .D (nx6198), .CLK (nx10321)) ;
    nand02 ix6199 (.Y (nx6198), .A0 (nx9431), .A1 (nx10863)) ;
    aoi22 ix9432 (.Y (nx9431), .A0 (d_arr_mul_4__22), .A1 (nx10553), .B0 (
          d_arr_add_4__22), .B1 (nx10709)) ;
    latch lat_d_arr_4__23 (.Q (d_arr_4__23), .D (nx6208), .CLK (nx10321)) ;
    nand02 ix6209 (.Y (nx6208), .A0 (nx9435), .A1 (nx10863)) ;
    aoi22 ix9436 (.Y (nx9435), .A0 (d_arr_mul_4__23), .A1 (nx10553), .B0 (
          d_arr_add_4__23), .B1 (nx10709)) ;
    latch lat_d_arr_4__24 (.Q (d_arr_4__24), .D (nx6218), .CLK (nx10321)) ;
    nand02 ix6219 (.Y (nx6218), .A0 (nx9439), .A1 (nx10863)) ;
    aoi22 ix9440 (.Y (nx9439), .A0 (d_arr_mul_4__24), .A1 (nx10553), .B0 (
          d_arr_add_4__24), .B1 (nx10709)) ;
    latch lat_d_arr_4__25 (.Q (d_arr_4__25), .D (nx6228), .CLK (nx10323)) ;
    nand02 ix6229 (.Y (nx6228), .A0 (nx9443), .A1 (nx10863)) ;
    aoi22 ix9444 (.Y (nx9443), .A0 (d_arr_mul_4__25), .A1 (nx10555), .B0 (
          d_arr_add_4__25), .B1 (nx10709)) ;
    latch lat_d_arr_4__26 (.Q (d_arr_4__26), .D (nx6238), .CLK (nx10323)) ;
    nand02 ix6239 (.Y (nx6238), .A0 (nx9447), .A1 (nx10863)) ;
    aoi22 ix9448 (.Y (nx9447), .A0 (d_arr_mul_4__26), .A1 (nx10555), .B0 (
          d_arr_add_4__26), .B1 (nx10709)) ;
    latch lat_d_arr_4__27 (.Q (d_arr_4__27), .D (nx6248), .CLK (nx10323)) ;
    nand02 ix6249 (.Y (nx6248), .A0 (nx9451), .A1 (nx10863)) ;
    aoi22 ix9452 (.Y (nx9451), .A0 (d_arr_mul_4__27), .A1 (nx10555), .B0 (
          d_arr_add_4__27), .B1 (nx10711)) ;
    latch lat_d_arr_4__28 (.Q (d_arr_4__28), .D (nx6258), .CLK (nx10323)) ;
    nand02 ix6259 (.Y (nx6258), .A0 (nx9455), .A1 (nx10863)) ;
    aoi22 ix9456 (.Y (nx9455), .A0 (d_arr_mul_4__28), .A1 (nx10555), .B0 (
          d_arr_add_4__28), .B1 (nx10711)) ;
    latch lat_d_arr_4__29 (.Q (d_arr_4__29), .D (nx6268), .CLK (nx10323)) ;
    nand02 ix6269 (.Y (nx6268), .A0 (nx9459), .A1 (nx9403)) ;
    aoi22 ix9460 (.Y (nx9459), .A0 (d_arr_mul_4__29), .A1 (nx10555), .B0 (
          d_arr_add_4__29), .B1 (nx10711)) ;
    latch lat_d_arr_4__30 (.Q (d_arr_4__30), .D (nx6278), .CLK (nx10323)) ;
    nand02 ix6279 (.Y (nx6278), .A0 (nx9463), .A1 (nx9403)) ;
    aoi22 ix9464 (.Y (nx9463), .A0 (d_arr_mul_4__30), .A1 (nx10555), .B0 (
          d_arr_add_4__30), .B1 (nx10711)) ;
    latch lat_d_arr_4__31 (.Q (d_arr_4__31), .D (nx6288), .CLK (nx10323)) ;
    nand02 ix6289 (.Y (nx6288), .A0 (nx9467), .A1 (nx9403)) ;
    aoi22 ix9468 (.Y (nx9467), .A0 (d_arr_mul_4__31), .A1 (nx10555), .B0 (
          d_arr_add_4__31), .B1 (nx10711)) ;
    latch lat_d_arr_3__0 (.Q (d_arr_3__0), .D (nx6300), .CLK (nx10325)) ;
    inv01 ix6301 (.Y (nx6300), .A (nx9471)) ;
    aoi222 ix9472 (.Y (nx9471), .A0 (d_arr_mux_3__0), .A1 (nx11379), .B0 (
           d_arr_mul_3__0), .B1 (nx10557), .C0 (d_arr_add_3__0), .C1 (nx10711)
           ) ;
    latch lat_d_arr_3__1 (.Q (d_arr_3__1), .D (nx6312), .CLK (nx10325)) ;
    inv01 ix6313 (.Y (nx6312), .A (nx9475)) ;
    aoi222 ix9476 (.Y (nx9475), .A0 (d_arr_mux_3__1), .A1 (nx11381), .B0 (
           d_arr_mul_3__1), .B1 (nx10557), .C0 (d_arr_add_3__1), .C1 (nx10711)
           ) ;
    latch lat_d_arr_3__2 (.Q (d_arr_3__2), .D (nx6324), .CLK (nx10325)) ;
    inv01 ix6325 (.Y (nx6324), .A (nx9479)) ;
    aoi222 ix9480 (.Y (nx9479), .A0 (d_arr_mux_3__2), .A1 (nx11381), .B0 (
           d_arr_mul_3__2), .B1 (nx10557), .C0 (d_arr_add_3__2), .C1 (nx10713)
           ) ;
    latch lat_d_arr_3__3 (.Q (d_arr_3__3), .D (nx6336), .CLK (nx10325)) ;
    inv01 ix6337 (.Y (nx6336), .A (nx9483)) ;
    aoi222 ix9484 (.Y (nx9483), .A0 (d_arr_mux_3__3), .A1 (nx11381), .B0 (
           d_arr_mul_3__3), .B1 (nx10557), .C0 (d_arr_add_3__3), .C1 (nx10713)
           ) ;
    latch lat_d_arr_3__4 (.Q (d_arr_3__4), .D (nx6348), .CLK (nx10325)) ;
    inv01 ix6349 (.Y (nx6348), .A (nx9487)) ;
    aoi222 ix9488 (.Y (nx9487), .A0 (d_arr_mux_3__4), .A1 (nx11381), .B0 (
           d_arr_mul_3__4), .B1 (nx10557), .C0 (d_arr_add_3__4), .C1 (nx10713)
           ) ;
    latch lat_d_arr_3__5 (.Q (d_arr_3__5), .D (nx6360), .CLK (nx10325)) ;
    inv01 ix6361 (.Y (nx6360), .A (nx9491)) ;
    aoi222 ix9492 (.Y (nx9491), .A0 (d_arr_mux_3__5), .A1 (nx11381), .B0 (
           d_arr_mul_3__5), .B1 (nx10557), .C0 (d_arr_add_3__5), .C1 (nx10713)
           ) ;
    latch lat_d_arr_3__6 (.Q (d_arr_3__6), .D (nx6372), .CLK (nx10325)) ;
    inv01 ix6373 (.Y (nx6372), .A (nx9495)) ;
    aoi222 ix9496 (.Y (nx9495), .A0 (d_arr_mux_3__6), .A1 (nx11381), .B0 (
           d_arr_mul_3__6), .B1 (nx10557), .C0 (d_arr_add_3__6), .C1 (nx10713)
           ) ;
    latch lat_d_arr_3__7 (.Q (d_arr_3__7), .D (nx6384), .CLK (nx10327)) ;
    inv01 ix6385 (.Y (nx6384), .A (nx9499)) ;
    aoi222 ix9500 (.Y (nx9499), .A0 (d_arr_mux_3__7), .A1 (nx11381), .B0 (
           d_arr_mul_3__7), .B1 (nx10559), .C0 (d_arr_add_3__7), .C1 (nx10713)
           ) ;
    latch lat_d_arr_3__8 (.Q (d_arr_3__8), .D (nx6396), .CLK (nx10327)) ;
    inv01 ix6397 (.Y (nx6396), .A (nx9503)) ;
    aoi222 ix9504 (.Y (nx9503), .A0 (d_arr_mux_3__8), .A1 (nx11383), .B0 (
           d_arr_mul_3__8), .B1 (nx10559), .C0 (d_arr_add_3__8), .C1 (nx10713)
           ) ;
    latch lat_d_arr_3__9 (.Q (d_arr_3__9), .D (nx6408), .CLK (nx10327)) ;
    inv01 ix6409 (.Y (nx6408), .A (nx9507)) ;
    aoi222 ix9508 (.Y (nx9507), .A0 (d_arr_mux_3__9), .A1 (nx11383), .B0 (
           d_arr_mul_3__9), .B1 (nx10559), .C0 (d_arr_add_3__9), .C1 (nx10715)
           ) ;
    latch lat_d_arr_3__10 (.Q (d_arr_3__10), .D (nx6420), .CLK (nx10327)) ;
    inv01 ix6421 (.Y (nx6420), .A (nx9511)) ;
    aoi222 ix9512 (.Y (nx9511), .A0 (d_arr_mux_3__10), .A1 (nx11383), .B0 (
           d_arr_mul_3__10), .B1 (nx10559), .C0 (d_arr_add_3__10), .C1 (nx10715)
           ) ;
    latch lat_d_arr_3__11 (.Q (d_arr_3__11), .D (nx6432), .CLK (nx10327)) ;
    inv01 ix6433 (.Y (nx6432), .A (nx9515)) ;
    aoi222 ix9516 (.Y (nx9515), .A0 (d_arr_mux_3__11), .A1 (nx11383), .B0 (
           d_arr_mul_3__11), .B1 (nx10559), .C0 (d_arr_add_3__11), .C1 (nx10715)
           ) ;
    latch lat_d_arr_3__12 (.Q (d_arr_3__12), .D (nx6444), .CLK (nx10327)) ;
    inv01 ix6445 (.Y (nx6444), .A (nx9519)) ;
    aoi222 ix9520 (.Y (nx9519), .A0 (d_arr_mux_3__12), .A1 (nx11383), .B0 (
           d_arr_mul_3__12), .B1 (nx10559), .C0 (d_arr_add_3__12), .C1 (nx10715)
           ) ;
    latch lat_d_arr_3__13 (.Q (d_arr_3__13), .D (nx6456), .CLK (nx10327)) ;
    inv01 ix6457 (.Y (nx6456), .A (nx9523)) ;
    aoi222 ix9524 (.Y (nx9523), .A0 (d_arr_mux_3__13), .A1 (nx11383), .B0 (
           d_arr_mul_3__13), .B1 (nx10559), .C0 (d_arr_add_3__13), .C1 (nx10715)
           ) ;
    latch lat_d_arr_3__14 (.Q (d_arr_3__14), .D (nx6468), .CLK (nx10329)) ;
    inv01 ix6469 (.Y (nx6468), .A (nx9527)) ;
    aoi222 ix9528 (.Y (nx9527), .A0 (d_arr_mux_3__14), .A1 (nx11383), .B0 (
           d_arr_mul_3__14), .B1 (nx10561), .C0 (d_arr_add_3__14), .C1 (nx10715)
           ) ;
    latch lat_d_arr_3__15 (.Q (d_arr_3__15), .D (nx6480), .CLK (nx10329)) ;
    nand02 ix6481 (.Y (nx6480), .A0 (nx9531), .A1 (nx10865)) ;
    aoi22 ix9532 (.Y (nx9531), .A0 (d_arr_mul_3__15), .A1 (nx10561), .B0 (
          d_arr_add_3__15), .B1 (nx10715)) ;
    nand02 ix9534 (.Y (nx9533), .A0 (d_arr_mux_3__31), .A1 (nx11385)) ;
    latch lat_d_arr_3__16 (.Q (d_arr_3__16), .D (nx6490), .CLK (nx10329)) ;
    nand02 ix6491 (.Y (nx6490), .A0 (nx9537), .A1 (nx10865)) ;
    aoi22 ix9538 (.Y (nx9537), .A0 (d_arr_mul_3__16), .A1 (nx10561), .B0 (
          d_arr_add_3__16), .B1 (nx10717)) ;
    latch lat_d_arr_3__17 (.Q (d_arr_3__17), .D (nx6500), .CLK (nx10329)) ;
    nand02 ix6501 (.Y (nx6500), .A0 (nx9541), .A1 (nx10865)) ;
    aoi22 ix9542 (.Y (nx9541), .A0 (d_arr_mul_3__17), .A1 (nx10561), .B0 (
          d_arr_add_3__17), .B1 (nx10717)) ;
    latch lat_d_arr_3__18 (.Q (d_arr_3__18), .D (nx6510), .CLK (nx10329)) ;
    nand02 ix6511 (.Y (nx6510), .A0 (nx9545), .A1 (nx10865)) ;
    aoi22 ix9546 (.Y (nx9545), .A0 (d_arr_mul_3__18), .A1 (nx10561), .B0 (
          d_arr_add_3__18), .B1 (nx10717)) ;
    latch lat_d_arr_3__19 (.Q (d_arr_3__19), .D (nx6520), .CLK (nx10329)) ;
    nand02 ix6521 (.Y (nx6520), .A0 (nx9549), .A1 (nx10865)) ;
    aoi22 ix9550 (.Y (nx9549), .A0 (d_arr_mul_3__19), .A1 (nx10561), .B0 (
          d_arr_add_3__19), .B1 (nx10717)) ;
    latch lat_d_arr_3__20 (.Q (d_arr_3__20), .D (nx6530), .CLK (nx10329)) ;
    nand02 ix6531 (.Y (nx6530), .A0 (nx9553), .A1 (nx10865)) ;
    aoi22 ix9554 (.Y (nx9553), .A0 (d_arr_mul_3__20), .A1 (nx10561), .B0 (
          d_arr_add_3__20), .B1 (nx10717)) ;
    latch lat_d_arr_3__21 (.Q (d_arr_3__21), .D (nx6540), .CLK (nx10331)) ;
    nand02 ix6541 (.Y (nx6540), .A0 (nx9557), .A1 (nx10865)) ;
    aoi22 ix9558 (.Y (nx9557), .A0 (d_arr_mul_3__21), .A1 (nx10563), .B0 (
          d_arr_add_3__21), .B1 (nx10717)) ;
    latch lat_d_arr_3__22 (.Q (d_arr_3__22), .D (nx6550), .CLK (nx10331)) ;
    nand02 ix6551 (.Y (nx6550), .A0 (nx9561), .A1 (nx10867)) ;
    aoi22 ix9562 (.Y (nx9561), .A0 (d_arr_mul_3__22), .A1 (nx10563), .B0 (
          d_arr_add_3__22), .B1 (nx10717)) ;
    latch lat_d_arr_3__23 (.Q (d_arr_3__23), .D (nx6560), .CLK (nx10331)) ;
    nand02 ix6561 (.Y (nx6560), .A0 (nx9565), .A1 (nx10867)) ;
    aoi22 ix9566 (.Y (nx9565), .A0 (d_arr_mul_3__23), .A1 (nx10563), .B0 (
          d_arr_add_3__23), .B1 (nx10719)) ;
    latch lat_d_arr_3__24 (.Q (d_arr_3__24), .D (nx6570), .CLK (nx10331)) ;
    nand02 ix6571 (.Y (nx6570), .A0 (nx9569), .A1 (nx10867)) ;
    aoi22 ix9570 (.Y (nx9569), .A0 (d_arr_mul_3__24), .A1 (nx10563), .B0 (
          d_arr_add_3__24), .B1 (nx10719)) ;
    latch lat_d_arr_3__25 (.Q (d_arr_3__25), .D (nx6580), .CLK (nx10331)) ;
    nand02 ix6581 (.Y (nx6580), .A0 (nx9573), .A1 (nx10867)) ;
    aoi22 ix9574 (.Y (nx9573), .A0 (d_arr_mul_3__25), .A1 (nx10563), .B0 (
          d_arr_add_3__25), .B1 (nx10719)) ;
    latch lat_d_arr_3__26 (.Q (d_arr_3__26), .D (nx6590), .CLK (nx10331)) ;
    nand02 ix6591 (.Y (nx6590), .A0 (nx9577), .A1 (nx10867)) ;
    aoi22 ix9578 (.Y (nx9577), .A0 (d_arr_mul_3__26), .A1 (nx10563), .B0 (
          d_arr_add_3__26), .B1 (nx10719)) ;
    latch lat_d_arr_3__27 (.Q (d_arr_3__27), .D (nx6600), .CLK (nx10331)) ;
    nand02 ix6601 (.Y (nx6600), .A0 (nx9581), .A1 (nx10867)) ;
    aoi22 ix9582 (.Y (nx9581), .A0 (d_arr_mul_3__27), .A1 (nx10563), .B0 (
          d_arr_add_3__27), .B1 (nx10719)) ;
    latch lat_d_arr_3__28 (.Q (d_arr_3__28), .D (nx6610), .CLK (nx10333)) ;
    nand02 ix6611 (.Y (nx6610), .A0 (nx9585), .A1 (nx10867)) ;
    aoi22 ix9586 (.Y (nx9585), .A0 (d_arr_mul_3__28), .A1 (nx10565), .B0 (
          d_arr_add_3__28), .B1 (nx10719)) ;
    latch lat_d_arr_3__29 (.Q (d_arr_3__29), .D (nx6620), .CLK (nx10333)) ;
    nand02 ix6621 (.Y (nx6620), .A0 (nx9589), .A1 (nx9533)) ;
    aoi22 ix9590 (.Y (nx9589), .A0 (d_arr_mul_3__29), .A1 (nx10565), .B0 (
          d_arr_add_3__29), .B1 (nx10719)) ;
    latch lat_d_arr_3__30 (.Q (d_arr_3__30), .D (nx6630), .CLK (nx10333)) ;
    nand02 ix6631 (.Y (nx6630), .A0 (nx9593), .A1 (nx9533)) ;
    aoi22 ix9594 (.Y (nx9593), .A0 (d_arr_mul_3__30), .A1 (nx10565), .B0 (
          d_arr_add_3__30), .B1 (nx10721)) ;
    latch lat_d_arr_3__31 (.Q (d_arr_3__31), .D (nx6640), .CLK (nx10333)) ;
    nand02 ix6641 (.Y (nx6640), .A0 (nx9597), .A1 (nx9533)) ;
    aoi22 ix9598 (.Y (nx9597), .A0 (d_arr_mul_3__31), .A1 (nx10565), .B0 (
          d_arr_add_3__31), .B1 (nx10721)) ;
    latch lat_d_arr_2__0 (.Q (d_arr_2__0), .D (nx6652), .CLK (nx10333)) ;
    inv01 ix6653 (.Y (nx6652), .A (nx9601)) ;
    aoi222 ix9602 (.Y (nx9601), .A0 (d_arr_mux_2__0), .A1 (nx11385), .B0 (
           d_arr_mul_2__0), .B1 (nx10565), .C0 (d_arr_add_2__0), .C1 (nx10721)
           ) ;
    latch lat_d_arr_2__1 (.Q (d_arr_2__1), .D (nx6664), .CLK (nx10333)) ;
    inv01 ix6665 (.Y (nx6664), .A (nx9605)) ;
    aoi222 ix9606 (.Y (nx9605), .A0 (d_arr_mux_2__1), .A1 (nx11385), .B0 (
           d_arr_mul_2__1), .B1 (nx10565), .C0 (d_arr_add_2__1), .C1 (nx10721)
           ) ;
    latch lat_d_arr_2__2 (.Q (d_arr_2__2), .D (nx6676), .CLK (nx10333)) ;
    inv01 ix6677 (.Y (nx6676), .A (nx9609)) ;
    aoi222 ix9610 (.Y (nx9609), .A0 (d_arr_mux_2__2), .A1 (nx11385), .B0 (
           d_arr_mul_2__2), .B1 (nx10565), .C0 (d_arr_add_2__2), .C1 (nx10721)
           ) ;
    latch lat_d_arr_2__3 (.Q (d_arr_2__3), .D (nx6688), .CLK (nx10335)) ;
    inv01 ix6689 (.Y (nx6688), .A (nx9613)) ;
    aoi222 ix9614 (.Y (nx9613), .A0 (d_arr_mux_2__3), .A1 (nx11385), .B0 (
           d_arr_mul_2__3), .B1 (nx10567), .C0 (d_arr_add_2__3), .C1 (nx10721)
           ) ;
    latch lat_d_arr_2__4 (.Q (d_arr_2__4), .D (nx6700), .CLK (nx10335)) ;
    inv01 ix6701 (.Y (nx6700), .A (nx9617)) ;
    aoi222 ix9618 (.Y (nx9617), .A0 (d_arr_mux_2__4), .A1 (nx11385), .B0 (
           d_arr_mul_2__4), .B1 (nx10567), .C0 (d_arr_add_2__4), .C1 (nx10721)
           ) ;
    latch lat_d_arr_2__5 (.Q (d_arr_2__5), .D (nx6712), .CLK (nx10335)) ;
    inv01 ix6713 (.Y (nx6712), .A (nx9621)) ;
    aoi222 ix9622 (.Y (nx9621), .A0 (d_arr_mux_2__5), .A1 (nx11385), .B0 (
           d_arr_mul_2__5), .B1 (nx10567), .C0 (d_arr_add_2__5), .C1 (nx10723)
           ) ;
    latch lat_d_arr_2__6 (.Q (d_arr_2__6), .D (nx6724), .CLK (nx10335)) ;
    inv01 ix6725 (.Y (nx6724), .A (nx9625)) ;
    aoi222 ix9626 (.Y (nx9625), .A0 (d_arr_mux_2__6), .A1 (nx11387), .B0 (
           d_arr_mul_2__6), .B1 (nx10567), .C0 (d_arr_add_2__6), .C1 (nx10723)
           ) ;
    latch lat_d_arr_2__7 (.Q (d_arr_2__7), .D (nx6736), .CLK (nx10335)) ;
    inv01 ix6737 (.Y (nx6736), .A (nx9629)) ;
    aoi222 ix9630 (.Y (nx9629), .A0 (d_arr_mux_2__7), .A1 (nx11387), .B0 (
           d_arr_mul_2__7), .B1 (nx10567), .C0 (d_arr_add_2__7), .C1 (nx10723)
           ) ;
    latch lat_d_arr_2__8 (.Q (d_arr_2__8), .D (nx6748), .CLK (nx10335)) ;
    inv01 ix6749 (.Y (nx6748), .A (nx9633)) ;
    aoi222 ix9634 (.Y (nx9633), .A0 (d_arr_mux_2__8), .A1 (nx11387), .B0 (
           d_arr_mul_2__8), .B1 (nx10567), .C0 (d_arr_add_2__8), .C1 (nx10723)
           ) ;
    latch lat_d_arr_2__9 (.Q (d_arr_2__9), .D (nx6760), .CLK (nx10335)) ;
    inv01 ix6761 (.Y (nx6760), .A (nx9637)) ;
    aoi222 ix9638 (.Y (nx9637), .A0 (d_arr_mux_2__9), .A1 (nx11387), .B0 (
           d_arr_mul_2__9), .B1 (nx10567), .C0 (d_arr_add_2__9), .C1 (nx10723)
           ) ;
    latch lat_d_arr_2__10 (.Q (d_arr_2__10), .D (nx6772), .CLK (nx10337)) ;
    inv01 ix6773 (.Y (nx6772), .A (nx9641)) ;
    aoi222 ix9642 (.Y (nx9641), .A0 (d_arr_mux_2__10), .A1 (nx11387), .B0 (
           d_arr_mul_2__10), .B1 (nx10569), .C0 (d_arr_add_2__10), .C1 (nx10723)
           ) ;
    latch lat_d_arr_2__11 (.Q (d_arr_2__11), .D (nx6784), .CLK (nx10337)) ;
    inv01 ix6785 (.Y (nx6784), .A (nx9645)) ;
    aoi222 ix9646 (.Y (nx9645), .A0 (d_arr_mux_2__11), .A1 (nx11387), .B0 (
           d_arr_mul_2__11), .B1 (nx10569), .C0 (d_arr_add_2__11), .C1 (nx10723)
           ) ;
    latch lat_d_arr_2__12 (.Q (d_arr_2__12), .D (nx6796), .CLK (nx10337)) ;
    inv01 ix6797 (.Y (nx6796), .A (nx9649)) ;
    aoi222 ix9650 (.Y (nx9649), .A0 (d_arr_mux_2__12), .A1 (nx11387), .B0 (
           d_arr_mul_2__12), .B1 (nx10569), .C0 (d_arr_add_2__12), .C1 (nx10725)
           ) ;
    latch lat_d_arr_2__13 (.Q (d_arr_2__13), .D (nx6808), .CLK (nx10337)) ;
    inv01 ix6809 (.Y (nx6808), .A (nx9653)) ;
    aoi222 ix9654 (.Y (nx9653), .A0 (d_arr_mux_2__13), .A1 (nx11389), .B0 (
           d_arr_mul_2__13), .B1 (nx10569), .C0 (d_arr_add_2__13), .C1 (nx10725)
           ) ;
    latch lat_d_arr_2__14 (.Q (d_arr_2__14), .D (nx6820), .CLK (nx10337)) ;
    inv01 ix6821 (.Y (nx6820), .A (nx9657)) ;
    aoi222 ix9658 (.Y (nx9657), .A0 (d_arr_mux_2__14), .A1 (nx11389), .B0 (
           d_arr_mul_2__14), .B1 (nx10569), .C0 (d_arr_add_2__14), .C1 (nx10725)
           ) ;
    latch lat_d_arr_2__15 (.Q (d_arr_2__15), .D (nx6832), .CLK (nx10337)) ;
    nand02 ix6833 (.Y (nx6832), .A0 (nx9661), .A1 (nx10869)) ;
    aoi22 ix9662 (.Y (nx9661), .A0 (d_arr_mul_2__15), .A1 (nx10569), .B0 (
          d_arr_add_2__15), .B1 (nx10725)) ;
    nand02 ix9664 (.Y (nx9663), .A0 (d_arr_mux_2__31), .A1 (nx11389)) ;
    latch lat_d_arr_2__16 (.Q (d_arr_2__16), .D (nx6842), .CLK (nx10337)) ;
    nand02 ix6843 (.Y (nx6842), .A0 (nx9667), .A1 (nx10869)) ;
    aoi22 ix9668 (.Y (nx9667), .A0 (d_arr_mul_2__16), .A1 (nx10569), .B0 (
          d_arr_add_2__16), .B1 (nx10725)) ;
    latch lat_d_arr_2__17 (.Q (d_arr_2__17), .D (nx6852), .CLK (nx10339)) ;
    nand02 ix6853 (.Y (nx6852), .A0 (nx9671), .A1 (nx10869)) ;
    aoi22 ix9672 (.Y (nx9671), .A0 (d_arr_mul_2__17), .A1 (nx10571), .B0 (
          d_arr_add_2__17), .B1 (nx10725)) ;
    latch lat_d_arr_2__18 (.Q (d_arr_2__18), .D (nx6862), .CLK (nx10339)) ;
    nand02 ix6863 (.Y (nx6862), .A0 (nx9675), .A1 (nx10869)) ;
    aoi22 ix9676 (.Y (nx9675), .A0 (d_arr_mul_2__18), .A1 (nx10571), .B0 (
          d_arr_add_2__18), .B1 (nx10725)) ;
    latch lat_d_arr_2__19 (.Q (d_arr_2__19), .D (nx6872), .CLK (nx10339)) ;
    nand02 ix6873 (.Y (nx6872), .A0 (nx9679), .A1 (nx10869)) ;
    aoi22 ix9680 (.Y (nx9679), .A0 (d_arr_mul_2__19), .A1 (nx10571), .B0 (
          d_arr_add_2__19), .B1 (nx10727)) ;
    latch lat_d_arr_2__20 (.Q (d_arr_2__20), .D (nx6882), .CLK (nx10339)) ;
    nand02 ix6883 (.Y (nx6882), .A0 (nx9683), .A1 (nx10869)) ;
    aoi22 ix9684 (.Y (nx9683), .A0 (d_arr_mul_2__20), .A1 (nx10571), .B0 (
          d_arr_add_2__20), .B1 (nx10727)) ;
    latch lat_d_arr_2__21 (.Q (d_arr_2__21), .D (nx6892), .CLK (nx10339)) ;
    nand02 ix6893 (.Y (nx6892), .A0 (nx9687), .A1 (nx10869)) ;
    aoi22 ix9688 (.Y (nx9687), .A0 (d_arr_mul_2__21), .A1 (nx10571), .B0 (
          d_arr_add_2__21), .B1 (nx10727)) ;
    latch lat_d_arr_2__22 (.Q (d_arr_2__22), .D (nx6902), .CLK (nx10339)) ;
    nand02 ix6903 (.Y (nx6902), .A0 (nx9691), .A1 (nx10871)) ;
    aoi22 ix9692 (.Y (nx9691), .A0 (d_arr_mul_2__22), .A1 (nx10571), .B0 (
          d_arr_add_2__22), .B1 (nx10727)) ;
    latch lat_d_arr_2__23 (.Q (d_arr_2__23), .D (nx6912), .CLK (nx10339)) ;
    nand02 ix6913 (.Y (nx6912), .A0 (nx9695), .A1 (nx10871)) ;
    aoi22 ix9696 (.Y (nx9695), .A0 (d_arr_mul_2__23), .A1 (nx10571), .B0 (
          d_arr_add_2__23), .B1 (nx10727)) ;
    latch lat_d_arr_2__24 (.Q (d_arr_2__24), .D (nx6922), .CLK (nx10341)) ;
    nand02 ix6923 (.Y (nx6922), .A0 (nx9699), .A1 (nx10871)) ;
    aoi22 ix9700 (.Y (nx9699), .A0 (d_arr_mul_2__24), .A1 (nx10573), .B0 (
          d_arr_add_2__24), .B1 (nx10727)) ;
    latch lat_d_arr_2__25 (.Q (d_arr_2__25), .D (nx6932), .CLK (nx10341)) ;
    nand02 ix6933 (.Y (nx6932), .A0 (nx9703), .A1 (nx10871)) ;
    aoi22 ix9704 (.Y (nx9703), .A0 (d_arr_mul_2__25), .A1 (nx10573), .B0 (
          d_arr_add_2__25), .B1 (nx10727)) ;
    latch lat_d_arr_2__26 (.Q (d_arr_2__26), .D (nx6942), .CLK (nx10341)) ;
    nand02 ix6943 (.Y (nx6942), .A0 (nx9707), .A1 (nx10871)) ;
    aoi22 ix9708 (.Y (nx9707), .A0 (d_arr_mul_2__26), .A1 (nx10573), .B0 (
          d_arr_add_2__26), .B1 (nx10729)) ;
    latch lat_d_arr_2__27 (.Q (d_arr_2__27), .D (nx6952), .CLK (nx10341)) ;
    nand02 ix6953 (.Y (nx6952), .A0 (nx9711), .A1 (nx10871)) ;
    aoi22 ix9712 (.Y (nx9711), .A0 (d_arr_mul_2__27), .A1 (nx10573), .B0 (
          d_arr_add_2__27), .B1 (nx10729)) ;
    latch lat_d_arr_2__28 (.Q (d_arr_2__28), .D (nx6962), .CLK (nx10341)) ;
    nand02 ix6963 (.Y (nx6962), .A0 (nx9715), .A1 (nx10871)) ;
    aoi22 ix9716 (.Y (nx9715), .A0 (d_arr_mul_2__28), .A1 (nx10573), .B0 (
          d_arr_add_2__28), .B1 (nx10729)) ;
    latch lat_d_arr_2__29 (.Q (d_arr_2__29), .D (nx6972), .CLK (nx10341)) ;
    nand02 ix6973 (.Y (nx6972), .A0 (nx9719), .A1 (nx9663)) ;
    aoi22 ix9720 (.Y (nx9719), .A0 (d_arr_mul_2__29), .A1 (nx10573), .B0 (
          d_arr_add_2__29), .B1 (nx10729)) ;
    latch lat_d_arr_2__30 (.Q (d_arr_2__30), .D (nx6982), .CLK (nx10341)) ;
    nand02 ix6983 (.Y (nx6982), .A0 (nx9723), .A1 (nx9663)) ;
    aoi22 ix9724 (.Y (nx9723), .A0 (d_arr_mul_2__30), .A1 (nx10573), .B0 (
          d_arr_add_2__30), .B1 (nx10729)) ;
    latch lat_d_arr_2__31 (.Q (d_arr_2__31), .D (nx6992), .CLK (nx10343)) ;
    nand02 ix6993 (.Y (nx6992), .A0 (nx9727), .A1 (nx9663)) ;
    aoi22 ix9728 (.Y (nx9727), .A0 (d_arr_mul_2__31), .A1 (nx10575), .B0 (
          d_arr_add_2__31), .B1 (nx10729)) ;
    latch lat_d_arr_1__0 (.Q (d_arr_1__0), .D (nx7036), .CLK (nx10343)) ;
    nand02 ix7037 (.Y (nx7036), .A0 (nx9731), .A1 (nx9739)) ;
    aoi222 ix9732 (.Y (nx9731), .A0 (d_arr_mux_1__0), .A1 (nx11389), .B0 (
           d_arr_merge2_1__0), .B1 (nx10805), .C0 (d_arr_relu_1__0), .C1 (
           nx10827)) ;
    and02 ix7019 (.Y (nx7018), .A0 (sel_merge2), .A1 (nx9734)) ;
    nor04 ix9735 (.Y (nx9734), .A0 (sel_add), .A1 (sel_merge1), .A2 (nx11389), .A3 (
          sel_mul)) ;
    and03 ix7029 (.Y (nx7028), .A0 (nx9734), .A1 (sel_relu), .A2 (nx9737)) ;
    inv01 ix9738 (.Y (nx9737), .A (sel_merge2)) ;
    aoi222 ix9740 (.Y (nx9739), .A0 (d_arr_mul_1__0), .A1 (nx10575), .B0 (
           d_arr_add_1__0), .B1 (nx10729), .C0 (d_arr_merge1_1__0), .C1 (nx10783
           )) ;
    nor04 ix7003 (.Y (nx7002), .A0 (nx11389), .A1 (sel_mul), .A2 (nx9742), .A3 (
          sel_add)) ;
    inv01 ix9743 (.Y (nx9742), .A (sel_merge1)) ;
    latch lat_d_arr_1__1 (.Q (d_arr_1__1), .D (nx7060), .CLK (nx10343)) ;
    nand02 ix7061 (.Y (nx7060), .A0 (nx9746), .A1 (nx9748)) ;
    aoi222 ix9747 (.Y (nx9746), .A0 (d_arr_mux_1__1), .A1 (nx11389), .B0 (
           d_arr_merge2_1__1), .B1 (nx10805), .C0 (d_arr_relu_1__1), .C1 (
           nx10827)) ;
    aoi222 ix9749 (.Y (nx9748), .A0 (d_arr_mul_1__1), .A1 (nx10575), .B0 (
           d_arr_add_1__1), .B1 (nx10731), .C0 (d_arr_merge1_1__1), .C1 (nx10783
           )) ;
    latch lat_d_arr_1__2 (.Q (d_arr_1__2), .D (nx7084), .CLK (nx10343)) ;
    nand02 ix7085 (.Y (nx7084), .A0 (nx9752), .A1 (nx9754)) ;
    aoi222 ix9753 (.Y (nx9752), .A0 (d_arr_mux_1__2), .A1 (nx11391), .B0 (
           d_arr_merge2_1__2), .B1 (nx10805), .C0 (d_arr_relu_1__2), .C1 (
           nx10827)) ;
    aoi222 ix9755 (.Y (nx9754), .A0 (d_arr_mul_1__2), .A1 (nx10575), .B0 (
           d_arr_add_1__2), .B1 (nx10731), .C0 (d_arr_merge1_1__2), .C1 (nx10783
           )) ;
    latch lat_d_arr_1__3 (.Q (d_arr_1__3), .D (nx7108), .CLK (nx10343)) ;
    nand02 ix7109 (.Y (nx7108), .A0 (nx9758), .A1 (nx9760)) ;
    aoi222 ix9759 (.Y (nx9758), .A0 (d_arr_mux_1__3), .A1 (nx11391), .B0 (
           d_arr_merge2_1__3), .B1 (nx10805), .C0 (d_arr_relu_1__3), .C1 (
           nx10827)) ;
    aoi222 ix9761 (.Y (nx9760), .A0 (d_arr_mul_1__3), .A1 (nx10575), .B0 (
           d_arr_add_1__3), .B1 (nx10731), .C0 (d_arr_merge1_1__3), .C1 (nx10783
           )) ;
    latch lat_d_arr_1__4 (.Q (d_arr_1__4), .D (nx7132), .CLK (nx10343)) ;
    nand02 ix7133 (.Y (nx7132), .A0 (nx9764), .A1 (nx9766)) ;
    aoi222 ix9765 (.Y (nx9764), .A0 (d_arr_mux_1__4), .A1 (nx11391), .B0 (
           d_arr_merge2_1__4), .B1 (nx10805), .C0 (d_arr_relu_1__4), .C1 (
           nx10827)) ;
    aoi222 ix9767 (.Y (nx9766), .A0 (d_arr_mul_1__4), .A1 (nx10575), .B0 (
           d_arr_add_1__4), .B1 (nx10731), .C0 (d_arr_merge1_1__4), .C1 (nx10783
           )) ;
    latch lat_d_arr_1__5 (.Q (d_arr_1__5), .D (nx7156), .CLK (nx10343)) ;
    nand02 ix7157 (.Y (nx7156), .A0 (nx9770), .A1 (nx9772)) ;
    aoi222 ix9771 (.Y (nx9770), .A0 (d_arr_mux_1__5), .A1 (nx11391), .B0 (
           d_arr_merge2_1__5), .B1 (nx10805), .C0 (d_arr_relu_1__5), .C1 (
           nx10827)) ;
    aoi222 ix9773 (.Y (nx9772), .A0 (d_arr_mul_1__5), .A1 (nx10575), .B0 (
           d_arr_add_1__5), .B1 (nx10731), .C0 (d_arr_merge1_1__5), .C1 (nx10783
           )) ;
    latch lat_d_arr_1__6 (.Q (d_arr_1__6), .D (nx7180), .CLK (nx10345)) ;
    nand02 ix7181 (.Y (nx7180), .A0 (nx9776), .A1 (nx9778)) ;
    aoi222 ix9777 (.Y (nx9776), .A0 (d_arr_mux_1__6), .A1 (nx11391), .B0 (
           d_arr_merge2_1__6), .B1 (nx10805), .C0 (d_arr_relu_1__6), .C1 (
           nx10827)) ;
    aoi222 ix9779 (.Y (nx9778), .A0 (d_arr_mul_1__6), .A1 (nx10577), .B0 (
           d_arr_add_1__6), .B1 (nx10731), .C0 (d_arr_merge1_1__6), .C1 (nx10783
           )) ;
    latch lat_d_arr_1__7 (.Q (d_arr_1__7), .D (nx7204), .CLK (nx10345)) ;
    nand02 ix7205 (.Y (nx7204), .A0 (nx9782), .A1 (nx9784)) ;
    aoi222 ix9783 (.Y (nx9782), .A0 (d_arr_mux_1__7), .A1 (nx11391), .B0 (
           d_arr_merge2_1__7), .B1 (nx10807), .C0 (d_arr_relu_1__7), .C1 (
           nx10829)) ;
    aoi222 ix9785 (.Y (nx9784), .A0 (d_arr_mul_1__7), .A1 (nx10577), .B0 (
           d_arr_add_1__7), .B1 (nx10731), .C0 (d_arr_merge1_1__7), .C1 (nx10785
           )) ;
    latch lat_d_arr_1__8 (.Q (d_arr_1__8), .D (nx7228), .CLK (nx10345)) ;
    nand02 ix7229 (.Y (nx7228), .A0 (nx9788), .A1 (nx9790)) ;
    aoi222 ix9789 (.Y (nx9788), .A0 (d_arr_mux_1__8), .A1 (nx11391), .B0 (
           d_arr_merge2_1__8), .B1 (nx10807), .C0 (d_arr_relu_1__8), .C1 (
           nx10829)) ;
    aoi222 ix9791 (.Y (nx9790), .A0 (d_arr_mul_1__8), .A1 (nx10577), .B0 (
           d_arr_add_1__8), .B1 (nx10733), .C0 (d_arr_merge1_1__8), .C1 (nx10785
           )) ;
    latch lat_d_arr_1__9 (.Q (d_arr_1__9), .D (nx7252), .CLK (nx10345)) ;
    nand02 ix7253 (.Y (nx7252), .A0 (nx9794), .A1 (nx9796)) ;
    aoi222 ix9795 (.Y (nx9794), .A0 (d_arr_mux_1__9), .A1 (nx11393), .B0 (
           d_arr_merge2_1__9), .B1 (nx10807), .C0 (d_arr_relu_1__9), .C1 (
           nx10829)) ;
    aoi222 ix9797 (.Y (nx9796), .A0 (d_arr_mul_1__9), .A1 (nx10577), .B0 (
           d_arr_add_1__9), .B1 (nx10733), .C0 (d_arr_merge1_1__9), .C1 (nx10785
           )) ;
    latch lat_d_arr_1__10 (.Q (d_arr_1__10), .D (nx7276), .CLK (nx10345)) ;
    nand02 ix7277 (.Y (nx7276), .A0 (nx9800), .A1 (nx9802)) ;
    aoi222 ix9801 (.Y (nx9800), .A0 (d_arr_mux_1__10), .A1 (nx11393), .B0 (
           d_arr_merge2_1__10), .B1 (nx10807), .C0 (d_arr_relu_1__10), .C1 (
           nx10829)) ;
    aoi222 ix9803 (.Y (nx9802), .A0 (d_arr_mul_1__10), .A1 (nx10577), .B0 (
           d_arr_add_1__10), .B1 (nx10733), .C0 (d_arr_merge1_1__10), .C1 (
           nx10785)) ;
    latch lat_d_arr_1__11 (.Q (d_arr_1__11), .D (nx7300), .CLK (nx10345)) ;
    nand02 ix7301 (.Y (nx7300), .A0 (nx9806), .A1 (nx9808)) ;
    aoi222 ix9807 (.Y (nx9806), .A0 (d_arr_mux_1__11), .A1 (nx11393), .B0 (
           d_arr_merge2_1__11), .B1 (nx10807), .C0 (d_arr_relu_1__11), .C1 (
           nx10829)) ;
    aoi222 ix9809 (.Y (nx9808), .A0 (d_arr_mul_1__11), .A1 (nx10577), .B0 (
           d_arr_add_1__11), .B1 (nx10733), .C0 (d_arr_merge1_1__11), .C1 (
           nx10785)) ;
    latch lat_d_arr_1__12 (.Q (d_arr_1__12), .D (nx7324), .CLK (nx10345)) ;
    nand02 ix7325 (.Y (nx7324), .A0 (nx9812), .A1 (nx9814)) ;
    aoi222 ix9813 (.Y (nx9812), .A0 (d_arr_mux_1__12), .A1 (nx11393), .B0 (
           d_arr_merge2_1__12), .B1 (nx10807), .C0 (d_arr_relu_1__12), .C1 (
           nx10829)) ;
    aoi222 ix9815 (.Y (nx9814), .A0 (d_arr_mul_1__12), .A1 (nx10577), .B0 (
           d_arr_add_1__12), .B1 (nx10733), .C0 (d_arr_merge1_1__12), .C1 (
           nx10785)) ;
    latch lat_d_arr_1__13 (.Q (d_arr_1__13), .D (nx7348), .CLK (nx10347)) ;
    nand02 ix7349 (.Y (nx7348), .A0 (nx9818), .A1 (nx9820)) ;
    aoi222 ix9819 (.Y (nx9818), .A0 (d_arr_mux_1__13), .A1 (nx11393), .B0 (
           d_arr_merge2_1__13), .B1 (nx10807), .C0 (d_arr_relu_1__13), .C1 (
           nx10829)) ;
    aoi222 ix9821 (.Y (nx9820), .A0 (d_arr_mul_1__13), .A1 (nx10579), .B0 (
           d_arr_add_1__13), .B1 (nx10733), .C0 (d_arr_merge1_1__13), .C1 (
           nx10785)) ;
    latch lat_d_arr_1__14 (.Q (d_arr_1__14), .D (nx7372), .CLK (nx10347)) ;
    nand02 ix7373 (.Y (nx7372), .A0 (nx9824), .A1 (nx9826)) ;
    aoi222 ix9825 (.Y (nx9824), .A0 (d_arr_mux_1__14), .A1 (nx11393), .B0 (
           d_arr_merge2_1__14), .B1 (nx10809), .C0 (d_arr_relu_1__14), .C1 (
           nx10831)) ;
    aoi222 ix9827 (.Y (nx9826), .A0 (d_arr_mul_1__14), .A1 (nx10579), .B0 (
           d_arr_add_1__14), .B1 (nx10733), .C0 (d_arr_merge1_1__14), .C1 (
           nx10787)) ;
    latch lat_d_arr_1__15 (.Q (d_arr_1__15), .D (nx7392), .CLK (nx10347)) ;
    nand03 ix7393 (.Y (nx7392), .A0 (nx9830), .A1 (nx10873), .A2 (nx9834)) ;
    nand02 ix9831 (.Y (nx9830), .A0 (d_arr_merge2_1__15), .A1 (nx10809)) ;
    nand02 ix9833 (.Y (nx9832), .A0 (d_arr_mux_1__31), .A1 (nx11393)) ;
    aoi222 ix9835 (.Y (nx9834), .A0 (d_arr_mul_1__15), .A1 (nx10579), .B0 (
           d_arr_add_1__15), .B1 (nx10735), .C0 (d_arr_merge1_1__15), .C1 (
           nx10787)) ;
    latch lat_d_arr_1__16 (.Q (d_arr_1__16), .D (nx7414), .CLK (nx10347)) ;
    nand03 ix7415 (.Y (nx7414), .A0 (nx9838), .A1 (nx10873), .A2 (nx9840)) ;
    aoi22 ix9839 (.Y (nx9838), .A0 (d_arr_merge2_1__16), .A1 (nx10809), .B0 (
          d_arr_relu_1__16), .B1 (nx10831)) ;
    aoi222 ix9841 (.Y (nx9840), .A0 (d_arr_mul_1__16), .A1 (nx10579), .B0 (
           d_arr_add_1__16), .B1 (nx10735), .C0 (d_arr_merge1_1__16), .C1 (
           nx10787)) ;
    latch lat_d_arr_1__17 (.Q (d_arr_1__17), .D (nx7436), .CLK (nx10347)) ;
    nand03 ix7437 (.Y (nx7436), .A0 (nx9844), .A1 (nx10873), .A2 (nx9846)) ;
    aoi22 ix9845 (.Y (nx9844), .A0 (d_arr_merge2_1__17), .A1 (nx10809), .B0 (
          d_arr_relu_1__17), .B1 (nx10831)) ;
    aoi222 ix9847 (.Y (nx9846), .A0 (d_arr_mul_1__17), .A1 (nx10579), .B0 (
           d_arr_add_1__17), .B1 (nx10735), .C0 (d_arr_merge1_1__17), .C1 (
           nx10787)) ;
    latch lat_d_arr_1__18 (.Q (d_arr_1__18), .D (nx7458), .CLK (nx10347)) ;
    nand03 ix7459 (.Y (nx7458), .A0 (nx9850), .A1 (nx10873), .A2 (nx9852)) ;
    aoi22 ix9851 (.Y (nx9850), .A0 (d_arr_merge2_1__18), .A1 (nx10809), .B0 (
          d_arr_relu_1__18), .B1 (nx10831)) ;
    aoi222 ix9853 (.Y (nx9852), .A0 (d_arr_mul_1__18), .A1 (nx10579), .B0 (
           d_arr_add_1__18), .B1 (nx10735), .C0 (d_arr_merge1_1__18), .C1 (
           nx10787)) ;
    latch lat_d_arr_1__19 (.Q (d_arr_1__19), .D (nx7480), .CLK (nx10347)) ;
    nand03 ix7481 (.Y (nx7480), .A0 (nx9856), .A1 (nx10873), .A2 (nx9858)) ;
    aoi22 ix9857 (.Y (nx9856), .A0 (d_arr_merge2_1__19), .A1 (nx10809), .B0 (
          d_arr_relu_1__19), .B1 (nx10831)) ;
    aoi222 ix9859 (.Y (nx9858), .A0 (d_arr_mul_1__19), .A1 (nx10579), .B0 (
           d_arr_add_1__19), .B1 (nx10735), .C0 (d_arr_merge1_1__19), .C1 (
           nx10787)) ;
    latch lat_d_arr_1__20 (.Q (d_arr_1__20), .D (nx7502), .CLK (nx10349)) ;
    nand03 ix7503 (.Y (nx7502), .A0 (nx9862), .A1 (nx10873), .A2 (nx9864)) ;
    aoi22 ix9863 (.Y (nx9862), .A0 (d_arr_merge2_1__20), .A1 (nx10809), .B0 (
          d_arr_relu_1__20), .B1 (nx10831)) ;
    aoi222 ix9865 (.Y (nx9864), .A0 (d_arr_mul_1__20), .A1 (nx10581), .B0 (
           d_arr_add_1__20), .B1 (nx10735), .C0 (d_arr_merge1_1__20), .C1 (
           nx10787)) ;
    latch lat_d_arr_1__21 (.Q (d_arr_1__21), .D (nx7524), .CLK (nx10349)) ;
    nand03 ix7525 (.Y (nx7524), .A0 (nx9868), .A1 (nx10873), .A2 (nx9870)) ;
    aoi22 ix9869 (.Y (nx9868), .A0 (d_arr_merge2_1__21), .A1 (nx10811), .B0 (
          d_arr_relu_1__21), .B1 (nx10831)) ;
    aoi222 ix9871 (.Y (nx9870), .A0 (d_arr_mul_1__21), .A1 (nx10581), .B0 (
           d_arr_add_1__21), .B1 (nx10735), .C0 (d_arr_merge1_1__21), .C1 (
           nx10789)) ;
    latch lat_d_arr_1__22 (.Q (d_arr_1__22), .D (nx7546), .CLK (nx10349)) ;
    nand03 ix7547 (.Y (nx7546), .A0 (nx9874), .A1 (nx10875), .A2 (nx9876)) ;
    aoi22 ix9875 (.Y (nx9874), .A0 (d_arr_merge2_1__22), .A1 (nx10811), .B0 (
          d_arr_relu_1__22), .B1 (nx10833)) ;
    aoi222 ix9877 (.Y (nx9876), .A0 (d_arr_mul_1__22), .A1 (nx10581), .B0 (
           d_arr_add_1__22), .B1 (nx10737), .C0 (d_arr_merge1_1__22), .C1 (
           nx10789)) ;
    latch lat_d_arr_1__23 (.Q (d_arr_1__23), .D (nx7568), .CLK (nx10349)) ;
    nand03 ix7569 (.Y (nx7568), .A0 (nx9880), .A1 (nx10875), .A2 (nx9882)) ;
    aoi22 ix9881 (.Y (nx9880), .A0 (d_arr_merge2_1__23), .A1 (nx10811), .B0 (
          d_arr_relu_1__23), .B1 (nx10833)) ;
    aoi222 ix9883 (.Y (nx9882), .A0 (d_arr_mul_1__23), .A1 (nx10581), .B0 (
           d_arr_add_1__23), .B1 (nx10737), .C0 (d_arr_merge1_1__23), .C1 (
           nx10789)) ;
    latch lat_d_arr_1__24 (.Q (d_arr_1__24), .D (nx7590), .CLK (nx10349)) ;
    nand03 ix7591 (.Y (nx7590), .A0 (nx9886), .A1 (nx10875), .A2 (nx9888)) ;
    aoi22 ix9887 (.Y (nx9886), .A0 (d_arr_merge2_1__24), .A1 (nx10811), .B0 (
          d_arr_relu_1__24), .B1 (nx10833)) ;
    aoi222 ix9889 (.Y (nx9888), .A0 (d_arr_mul_1__24), .A1 (nx10581), .B0 (
           d_arr_add_1__24), .B1 (nx10737), .C0 (d_arr_merge1_1__24), .C1 (
           nx10789)) ;
    latch lat_d_arr_1__25 (.Q (d_arr_1__25), .D (nx7612), .CLK (nx10349)) ;
    nand03 ix7613 (.Y (nx7612), .A0 (nx9892), .A1 (nx10875), .A2 (nx9894)) ;
    aoi22 ix9893 (.Y (nx9892), .A0 (d_arr_merge2_1__25), .A1 (nx10811), .B0 (
          d_arr_relu_1__25), .B1 (nx10833)) ;
    aoi222 ix9895 (.Y (nx9894), .A0 (d_arr_mul_1__25), .A1 (nx10581), .B0 (
           d_arr_add_1__25), .B1 (nx10737), .C0 (d_arr_merge1_1__25), .C1 (
           nx10789)) ;
    latch lat_d_arr_1__26 (.Q (d_arr_1__26), .D (nx7634), .CLK (nx10349)) ;
    nand03 ix7635 (.Y (nx7634), .A0 (nx9898), .A1 (nx10875), .A2 (nx9900)) ;
    aoi22 ix9899 (.Y (nx9898), .A0 (d_arr_merge2_1__26), .A1 (nx10811), .B0 (
          d_arr_relu_1__26), .B1 (nx10833)) ;
    aoi222 ix9901 (.Y (nx9900), .A0 (d_arr_mul_1__26), .A1 (nx10581), .B0 (
           d_arr_add_1__26), .B1 (nx10737), .C0 (d_arr_merge1_1__26), .C1 (
           nx10789)) ;
    latch lat_d_arr_1__27 (.Q (d_arr_1__27), .D (nx7656), .CLK (nx10351)) ;
    nand03 ix7657 (.Y (nx7656), .A0 (nx9904), .A1 (nx10875), .A2 (nx9906)) ;
    aoi22 ix9905 (.Y (nx9904), .A0 (d_arr_merge2_1__27), .A1 (nx10811), .B0 (
          d_arr_relu_1__27), .B1 (nx10833)) ;
    aoi222 ix9907 (.Y (nx9906), .A0 (d_arr_mul_1__27), .A1 (nx10583), .B0 (
           d_arr_add_1__27), .B1 (nx10737), .C0 (d_arr_merge1_1__27), .C1 (
           nx10789)) ;
    latch lat_d_arr_1__28 (.Q (d_arr_1__28), .D (nx7678), .CLK (nx10351)) ;
    nand03 ix7679 (.Y (nx7678), .A0 (nx9910), .A1 (nx10875), .A2 (nx9912)) ;
    aoi22 ix9911 (.Y (nx9910), .A0 (d_arr_merge2_1__28), .A1 (nx10813), .B0 (
          d_arr_relu_1__28), .B1 (nx10833)) ;
    aoi222 ix9913 (.Y (nx9912), .A0 (d_arr_mul_1__28), .A1 (nx10583), .B0 (
           d_arr_add_1__28), .B1 (nx10737), .C0 (d_arr_merge1_1__28), .C1 (
           nx10791)) ;
    latch lat_d_arr_1__29 (.Q (d_arr_1__29), .D (nx7700), .CLK (nx10351)) ;
    nand03 ix7701 (.Y (nx7700), .A0 (nx9916), .A1 (nx9832), .A2 (nx9918)) ;
    aoi22 ix9917 (.Y (nx9916), .A0 (d_arr_merge2_1__29), .A1 (nx10813), .B0 (
          d_arr_relu_1__29), .B1 (nx10835)) ;
    aoi222 ix9919 (.Y (nx9918), .A0 (d_arr_mul_1__29), .A1 (nx10583), .B0 (
           d_arr_add_1__29), .B1 (nx10739), .C0 (d_arr_merge1_1__29), .C1 (
           nx10791)) ;
    latch lat_d_arr_1__30 (.Q (d_arr_1__30), .D (nx7722), .CLK (nx10351)) ;
    nand03 ix7723 (.Y (nx7722), .A0 (nx9922), .A1 (nx9832), .A2 (nx9924)) ;
    aoi22 ix9923 (.Y (nx9922), .A0 (d_arr_merge2_1__30), .A1 (nx10813), .B0 (
          d_arr_relu_1__30), .B1 (nx10835)) ;
    aoi222 ix9925 (.Y (nx9924), .A0 (d_arr_mul_1__30), .A1 (nx10583), .B0 (
           d_arr_add_1__30), .B1 (nx10739), .C0 (d_arr_merge1_1__30), .C1 (
           nx10791)) ;
    latch lat_d_arr_1__31 (.Q (d_arr_1__31), .D (nx7744), .CLK (nx10351)) ;
    nand03 ix7745 (.Y (nx7744), .A0 (nx9928), .A1 (nx9832), .A2 (nx9930)) ;
    aoi22 ix9929 (.Y (nx9928), .A0 (d_arr_merge2_1__31), .A1 (nx10813), .B0 (
          d_arr_relu_1__31), .B1 (nx10835)) ;
    aoi222 ix9931 (.Y (nx9930), .A0 (d_arr_mul_1__31), .A1 (nx10583), .B0 (
           d_arr_add_1__31), .B1 (nx10739), .C0 (d_arr_merge1_1__31), .C1 (
           nx10791)) ;
    latch lat_d_arr_0__0 (.Q (d_arr_0__0), .D (nx7768), .CLK (nx10351)) ;
    nand02 ix7769 (.Y (nx7768), .A0 (nx9934), .A1 (nx9936)) ;
    aoi222 ix9935 (.Y (nx9934), .A0 (d_arr_mux_0__0), .A1 (nx11395), .B0 (
           d_arr_merge2_0__0), .B1 (nx10813), .C0 (d_arr_relu_0__0), .C1 (
           nx10835)) ;
    aoi222 ix9937 (.Y (nx9936), .A0 (d_arr_mul_0__0), .A1 (nx10583), .B0 (
           d_arr_add_0__0), .B1 (nx10739), .C0 (d_arr_merge1_0__0), .C1 (nx10791
           )) ;
    latch lat_d_arr_0__1 (.Q (d_arr_0__1), .D (nx7792), .CLK (nx10351)) ;
    nand02 ix7793 (.Y (nx7792), .A0 (nx9940), .A1 (nx9942)) ;
    aoi222 ix9941 (.Y (nx9940), .A0 (d_arr_mux_0__1), .A1 (nx11395), .B0 (
           d_arr_merge2_0__1), .B1 (nx10813), .C0 (d_arr_relu_0__1), .C1 (
           nx10835)) ;
    aoi222 ix9943 (.Y (nx9942), .A0 (d_arr_mul_0__1), .A1 (nx10583), .B0 (
           d_arr_add_0__1), .B1 (nx10739), .C0 (d_arr_merge1_0__1), .C1 (nx10791
           )) ;
    latch lat_d_arr_0__2 (.Q (d_arr_0__2), .D (nx7816), .CLK (nx10353)) ;
    nand02 ix7817 (.Y (nx7816), .A0 (nx9946), .A1 (nx9948)) ;
    aoi222 ix9947 (.Y (nx9946), .A0 (d_arr_mux_0__2), .A1 (nx11395), .B0 (
           d_arr_merge2_0__2), .B1 (nx10813), .C0 (d_arr_relu_0__2), .C1 (
           nx10835)) ;
    aoi222 ix9949 (.Y (nx9948), .A0 (d_arr_mul_0__2), .A1 (nx10585), .B0 (
           d_arr_add_0__2), .B1 (nx10739), .C0 (d_arr_merge1_0__2), .C1 (nx10791
           )) ;
    latch lat_d_arr_0__3 (.Q (d_arr_0__3), .D (nx7840), .CLK (nx10353)) ;
    nand02 ix7841 (.Y (nx7840), .A0 (nx9952), .A1 (nx9954)) ;
    aoi222 ix9953 (.Y (nx9952), .A0 (d_arr_mux_0__3), .A1 (nx11395), .B0 (
           d_arr_merge2_0__3), .B1 (nx10815), .C0 (d_arr_relu_0__3), .C1 (
           nx10835)) ;
    aoi222 ix9955 (.Y (nx9954), .A0 (d_arr_mul_0__3), .A1 (nx10585), .B0 (
           d_arr_add_0__3), .B1 (nx10739), .C0 (d_arr_merge1_0__3), .C1 (nx10793
           )) ;
    latch lat_d_arr_0__4 (.Q (d_arr_0__4), .D (nx7864), .CLK (nx10353)) ;
    nand02 ix7865 (.Y (nx7864), .A0 (nx9958), .A1 (nx9960)) ;
    aoi222 ix9959 (.Y (nx9958), .A0 (d_arr_mux_0__4), .A1 (nx11395), .B0 (
           d_arr_merge2_0__4), .B1 (nx10815), .C0 (d_arr_relu_0__4), .C1 (
           nx10837)) ;
    aoi222 ix9961 (.Y (nx9960), .A0 (d_arr_mul_0__4), .A1 (nx10585), .B0 (
           d_arr_add_0__4), .B1 (nx10741), .C0 (d_arr_merge1_0__4), .C1 (nx10793
           )) ;
    latch lat_d_arr_0__5 (.Q (d_arr_0__5), .D (nx7888), .CLK (nx10353)) ;
    nand02 ix7889 (.Y (nx7888), .A0 (nx9964), .A1 (nx9966)) ;
    aoi222 ix9965 (.Y (nx9964), .A0 (d_arr_mux_0__5), .A1 (nx11395), .B0 (
           d_arr_merge2_0__5), .B1 (nx10815), .C0 (d_arr_relu_0__5), .C1 (
           nx10837)) ;
    aoi222 ix9967 (.Y (nx9966), .A0 (d_arr_mul_0__5), .A1 (nx10585), .B0 (
           d_arr_add_0__5), .B1 (nx10741), .C0 (d_arr_merge1_0__5), .C1 (nx10793
           )) ;
    latch lat_d_arr_0__6 (.Q (d_arr_0__6), .D (nx7912), .CLK (nx10353)) ;
    nand02 ix7913 (.Y (nx7912), .A0 (nx9970), .A1 (nx9972)) ;
    aoi222 ix9971 (.Y (nx9970), .A0 (d_arr_mux_0__6), .A1 (nx11395), .B0 (
           d_arr_merge2_0__6), .B1 (nx10815), .C0 (d_arr_relu_0__6), .C1 (
           nx10837)) ;
    aoi222 ix9973 (.Y (nx9972), .A0 (d_arr_mul_0__6), .A1 (nx10585), .B0 (
           d_arr_add_0__6), .B1 (nx10741), .C0 (d_arr_merge1_0__6), .C1 (nx10793
           )) ;
    latch lat_d_arr_0__7 (.Q (d_arr_0__7), .D (nx7936), .CLK (nx10353)) ;
    nand02 ix7937 (.Y (nx7936), .A0 (nx9976), .A1 (nx9978)) ;
    aoi222 ix9977 (.Y (nx9976), .A0 (d_arr_mux_0__7), .A1 (nx11397), .B0 (
           d_arr_merge2_0__7), .B1 (nx10815), .C0 (d_arr_relu_0__7), .C1 (
           nx10837)) ;
    aoi222 ix9979 (.Y (nx9978), .A0 (d_arr_mul_0__7), .A1 (nx10585), .B0 (
           d_arr_add_0__7), .B1 (nx10741), .C0 (d_arr_merge1_0__7), .C1 (nx10793
           )) ;
    latch lat_d_arr_0__8 (.Q (d_arr_0__8), .D (nx7960), .CLK (nx10353)) ;
    nand02 ix7961 (.Y (nx7960), .A0 (nx9982), .A1 (nx9984)) ;
    aoi222 ix9983 (.Y (nx9982), .A0 (d_arr_mux_0__8), .A1 (nx11397), .B0 (
           d_arr_merge2_0__8), .B1 (nx10815), .C0 (d_arr_relu_0__8), .C1 (
           nx10837)) ;
    aoi222 ix9985 (.Y (nx9984), .A0 (d_arr_mul_0__8), .A1 (nx10585), .B0 (
           d_arr_add_0__8), .B1 (nx10741), .C0 (d_arr_merge1_0__8), .C1 (nx10793
           )) ;
    latch lat_d_arr_0__9 (.Q (d_arr_0__9), .D (nx7984), .CLK (nx10355)) ;
    nand02 ix7985 (.Y (nx7984), .A0 (nx9988), .A1 (nx9990)) ;
    aoi222 ix9989 (.Y (nx9988), .A0 (d_arr_mux_0__9), .A1 (nx11397), .B0 (
           d_arr_merge2_0__9), .B1 (nx10815), .C0 (d_arr_relu_0__9), .C1 (
           nx10837)) ;
    aoi222 ix9991 (.Y (nx9990), .A0 (d_arr_mul_0__9), .A1 (nx10587), .B0 (
           d_arr_add_0__9), .B1 (nx10741), .C0 (d_arr_merge1_0__9), .C1 (nx10793
           )) ;
    latch lat_d_arr_0__10 (.Q (d_arr_0__10), .D (nx8008), .CLK (nx10355)) ;
    nand02 ix8009 (.Y (nx8008), .A0 (nx9994), .A1 (nx9996)) ;
    aoi222 ix9995 (.Y (nx9994), .A0 (d_arr_mux_0__10), .A1 (nx11397), .B0 (
           d_arr_merge2_0__10), .B1 (nx10817), .C0 (d_arr_relu_0__10), .C1 (
           nx10837)) ;
    aoi222 ix9997 (.Y (nx9996), .A0 (d_arr_mul_0__10), .A1 (nx10587), .B0 (
           d_arr_add_0__10), .B1 (nx10741), .C0 (d_arr_merge1_0__10), .C1 (
           nx10795)) ;
    latch lat_d_arr_0__11 (.Q (d_arr_0__11), .D (nx8032), .CLK (nx10355)) ;
    nand02 ix8033 (.Y (nx8032), .A0 (nx10000), .A1 (nx10002)) ;
    aoi222 ix10001 (.Y (nx10000), .A0 (d_arr_mux_0__11), .A1 (nx11397), .B0 (
           d_arr_merge2_0__11), .B1 (nx10817), .C0 (d_arr_relu_0__11), .C1 (
           nx10839)) ;
    aoi222 ix10003 (.Y (nx10002), .A0 (d_arr_mul_0__11), .A1 (nx10587), .B0 (
           d_arr_add_0__11), .B1 (nx10743), .C0 (d_arr_merge1_0__11), .C1 (
           nx10795)) ;
    latch lat_d_arr_0__12 (.Q (d_arr_0__12), .D (nx8056), .CLK (nx10355)) ;
    nand02 ix8057 (.Y (nx8056), .A0 (nx10006), .A1 (nx10008)) ;
    aoi222 ix10007 (.Y (nx10006), .A0 (d_arr_mux_0__12), .A1 (nx11397), .B0 (
           d_arr_merge2_0__12), .B1 (nx10817), .C0 (d_arr_relu_0__12), .C1 (
           nx10839)) ;
    aoi222 ix10009 (.Y (nx10008), .A0 (d_arr_mul_0__12), .A1 (nx10587), .B0 (
           d_arr_add_0__12), .B1 (nx10743), .C0 (d_arr_merge1_0__12), .C1 (
           nx10795)) ;
    latch lat_d_arr_0__13 (.Q (d_arr_0__13), .D (nx8080), .CLK (nx10355)) ;
    nand02 ix8081 (.Y (nx8080), .A0 (nx10012), .A1 (nx10014)) ;
    aoi222 ix10013 (.Y (nx10012), .A0 (d_arr_mux_0__13), .A1 (nx11397), .B0 (
           d_arr_merge2_0__13), .B1 (nx10817), .C0 (d_arr_relu_0__13), .C1 (
           nx10839)) ;
    aoi222 ix10015 (.Y (nx10014), .A0 (d_arr_mul_0__13), .A1 (nx10587), .B0 (
           d_arr_add_0__13), .B1 (nx10743), .C0 (d_arr_merge1_0__13), .C1 (
           nx10795)) ;
    latch lat_d_arr_0__14 (.Q (d_arr_0__14), .D (nx8104), .CLK (nx10355)) ;
    nand02 ix8105 (.Y (nx8104), .A0 (nx10018), .A1 (nx10020)) ;
    aoi222 ix10019 (.Y (nx10018), .A0 (d_arr_mux_0__14), .A1 (nx11399), .B0 (
           d_arr_merge2_0__14), .B1 (nx10817), .C0 (d_arr_relu_0__14), .C1 (
           nx10839)) ;
    aoi222 ix10021 (.Y (nx10020), .A0 (d_arr_mul_0__14), .A1 (nx10587), .B0 (
           d_arr_add_0__14), .B1 (nx10743), .C0 (d_arr_merge1_0__14), .C1 (
           nx10795)) ;
    latch lat_d_arr_0__15 (.Q (d_arr_0__15), .D (nx8124), .CLK (nx10355)) ;
    nand03 ix8125 (.Y (nx8124), .A0 (nx10024), .A1 (nx10877), .A2 (nx10028)) ;
    nand02 ix10025 (.Y (nx10024), .A0 (d_arr_merge2_0__15), .A1 (nx10817)) ;
    nand02 ix10027 (.Y (nx10026), .A0 (d_arr_mux_0__31), .A1 (nx11399)) ;
    aoi222 ix10029 (.Y (nx10028), .A0 (d_arr_mul_0__15), .A1 (nx10587), .B0 (
           d_arr_add_0__15), .B1 (nx10743), .C0 (d_arr_merge1_0__15), .C1 (
           nx10795)) ;
    latch lat_d_arr_0__16 (.Q (d_arr_0__16), .D (nx8146), .CLK (nx10357)) ;
    nand03 ix8147 (.Y (nx8146), .A0 (nx10032), .A1 (nx10877), .A2 (nx10034)) ;
    aoi22 ix10033 (.Y (nx10032), .A0 (d_arr_merge2_0__16), .A1 (nx10817), .B0 (
          d_arr_relu_0__16), .B1 (nx10839)) ;
    aoi222 ix10035 (.Y (nx10034), .A0 (d_arr_mul_0__16), .A1 (nx10589), .B0 (
           d_arr_add_0__16), .B1 (nx10743), .C0 (d_arr_merge1_0__16), .C1 (
           nx10795)) ;
    latch lat_d_arr_0__17 (.Q (d_arr_0__17), .D (nx8168), .CLK (nx10357)) ;
    nand03 ix8169 (.Y (nx8168), .A0 (nx10038), .A1 (nx10877), .A2 (nx10040)) ;
    aoi22 ix10039 (.Y (nx10038), .A0 (d_arr_merge2_0__17), .A1 (nx10819), .B0 (
          d_arr_relu_0__17), .B1 (nx10839)) ;
    aoi222 ix10041 (.Y (nx10040), .A0 (d_arr_mul_0__17), .A1 (nx10589), .B0 (
           d_arr_add_0__17), .B1 (nx10743), .C0 (d_arr_merge1_0__17), .C1 (
           nx10797)) ;
    latch lat_d_arr_0__18 (.Q (d_arr_0__18), .D (nx8190), .CLK (nx10357)) ;
    nand03 ix8191 (.Y (nx8190), .A0 (nx10044), .A1 (nx10877), .A2 (nx10046)) ;
    aoi22 ix10045 (.Y (nx10044), .A0 (d_arr_merge2_0__18), .A1 (nx10819), .B0 (
          d_arr_relu_0__18), .B1 (nx10839)) ;
    aoi222 ix10047 (.Y (nx10046), .A0 (d_arr_mul_0__18), .A1 (nx10589), .B0 (
           d_arr_add_0__18), .B1 (nx10745), .C0 (d_arr_merge1_0__18), .C1 (
           nx10797)) ;
    latch lat_d_arr_0__19 (.Q (d_arr_0__19), .D (nx8212), .CLK (nx10357)) ;
    nand03 ix8213 (.Y (nx8212), .A0 (nx10050), .A1 (nx10877), .A2 (nx10052)) ;
    aoi22 ix10051 (.Y (nx10050), .A0 (d_arr_merge2_0__19), .A1 (nx10819), .B0 (
          d_arr_relu_0__19), .B1 (nx10841)) ;
    aoi222 ix10053 (.Y (nx10052), .A0 (d_arr_mul_0__19), .A1 (nx10589), .B0 (
           d_arr_add_0__19), .B1 (nx10745), .C0 (d_arr_merge1_0__19), .C1 (
           nx10797)) ;
    latch lat_d_arr_0__20 (.Q (d_arr_0__20), .D (nx8234), .CLK (nx10357)) ;
    nand03 ix8235 (.Y (nx8234), .A0 (nx10056), .A1 (nx10877), .A2 (nx10058)) ;
    aoi22 ix10057 (.Y (nx10056), .A0 (d_arr_merge2_0__20), .A1 (nx10819), .B0 (
          d_arr_relu_0__20), .B1 (nx10841)) ;
    aoi222 ix10059 (.Y (nx10058), .A0 (d_arr_mul_0__20), .A1 (nx10589), .B0 (
           d_arr_add_0__20), .B1 (nx10745), .C0 (d_arr_merge1_0__20), .C1 (
           nx10797)) ;
    latch lat_d_arr_0__21 (.Q (d_arr_0__21), .D (nx8256), .CLK (nx10357)) ;
    nand03 ix8257 (.Y (nx8256), .A0 (nx10062), .A1 (nx10877), .A2 (nx10064)) ;
    aoi22 ix10063 (.Y (nx10062), .A0 (d_arr_merge2_0__21), .A1 (nx10819), .B0 (
          d_arr_relu_0__21), .B1 (nx10841)) ;
    aoi222 ix10065 (.Y (nx10064), .A0 (d_arr_mul_0__21), .A1 (nx10589), .B0 (
           d_arr_add_0__21), .B1 (nx10745), .C0 (d_arr_merge1_0__21), .C1 (
           nx10797)) ;
    latch lat_d_arr_0__22 (.Q (d_arr_0__22), .D (nx8278), .CLK (nx10357)) ;
    nand03 ix8279 (.Y (nx8278), .A0 (nx10068), .A1 (nx10879), .A2 (nx10070)) ;
    aoi22 ix10069 (.Y (nx10068), .A0 (d_arr_merge2_0__22), .A1 (nx10819), .B0 (
          d_arr_relu_0__22), .B1 (nx10841)) ;
    aoi222 ix10071 (.Y (nx10070), .A0 (d_arr_mul_0__22), .A1 (nx10589), .B0 (
           d_arr_add_0__22), .B1 (nx10745), .C0 (d_arr_merge1_0__22), .C1 (
           nx10797)) ;
    latch lat_d_arr_0__23 (.Q (d_arr_0__23), .D (nx8300), .CLK (nx10359)) ;
    nand03 ix8301 (.Y (nx8300), .A0 (nx10074), .A1 (nx10879), .A2 (nx10076)) ;
    aoi22 ix10075 (.Y (nx10074), .A0 (d_arr_merge2_0__23), .A1 (nx10819), .B0 (
          d_arr_relu_0__23), .B1 (nx10841)) ;
    aoi222 ix10077 (.Y (nx10076), .A0 (d_arr_mul_0__23), .A1 (nx10591), .B0 (
           d_arr_add_0__23), .B1 (nx10745), .C0 (d_arr_merge1_0__23), .C1 (
           nx10797)) ;
    latch lat_d_arr_0__24 (.Q (d_arr_0__24), .D (nx8322), .CLK (nx10359)) ;
    nand03 ix8323 (.Y (nx8322), .A0 (nx10080), .A1 (nx10879), .A2 (nx10082)) ;
    aoi22 ix10081 (.Y (nx10080), .A0 (d_arr_merge2_0__24), .A1 (nx10821), .B0 (
          d_arr_relu_0__24), .B1 (nx10841)) ;
    aoi222 ix10083 (.Y (nx10082), .A0 (d_arr_mul_0__24), .A1 (nx10591), .B0 (
           d_arr_add_0__24), .B1 (nx10745), .C0 (d_arr_merge1_0__24), .C1 (
           nx10799)) ;
    latch lat_d_arr_0__25 (.Q (d_arr_0__25), .D (nx8344), .CLK (nx10359)) ;
    nand03 ix8345 (.Y (nx8344), .A0 (nx10086), .A1 (nx10879), .A2 (nx10088)) ;
    aoi22 ix10087 (.Y (nx10086), .A0 (d_arr_merge2_0__25), .A1 (nx10821), .B0 (
          d_arr_relu_0__25), .B1 (nx10841)) ;
    aoi222 ix10089 (.Y (nx10088), .A0 (d_arr_mul_0__25), .A1 (nx10591), .B0 (
           d_arr_add_0__25), .B1 (nx10747), .C0 (d_arr_merge1_0__25), .C1 (
           nx10799)) ;
    latch lat_d_arr_0__26 (.Q (d_arr_0__26), .D (nx8366), .CLK (nx10359)) ;
    nand03 ix8367 (.Y (nx8366), .A0 (nx10092), .A1 (nx10879), .A2 (nx10094)) ;
    aoi22 ix10093 (.Y (nx10092), .A0 (d_arr_merge2_0__26), .A1 (nx10821), .B0 (
          d_arr_relu_0__26), .B1 (nx10843)) ;
    aoi222 ix10095 (.Y (nx10094), .A0 (d_arr_mul_0__26), .A1 (nx10591), .B0 (
           d_arr_add_0__26), .B1 (nx10747), .C0 (d_arr_merge1_0__26), .C1 (
           nx10799)) ;
    latch lat_d_arr_0__27 (.Q (d_arr_0__27), .D (nx8388), .CLK (nx10359)) ;
    nand03 ix8389 (.Y (nx8388), .A0 (nx10098), .A1 (nx10879), .A2 (nx10100)) ;
    aoi22 ix10099 (.Y (nx10098), .A0 (d_arr_merge2_0__27), .A1 (nx10821), .B0 (
          d_arr_relu_0__27), .B1 (nx10843)) ;
    aoi222 ix10101 (.Y (nx10100), .A0 (d_arr_mul_0__27), .A1 (nx10591), .B0 (
           d_arr_add_0__27), .B1 (nx10747), .C0 (d_arr_merge1_0__27), .C1 (
           nx10799)) ;
    latch lat_d_arr_0__28 (.Q (d_arr_0__28), .D (nx8410), .CLK (nx10359)) ;
    nand03 ix8411 (.Y (nx8410), .A0 (nx10104), .A1 (nx10879), .A2 (nx10106)) ;
    aoi22 ix10105 (.Y (nx10104), .A0 (d_arr_merge2_0__28), .A1 (nx10821), .B0 (
          d_arr_relu_0__28), .B1 (nx10843)) ;
    aoi222 ix10107 (.Y (nx10106), .A0 (d_arr_mul_0__28), .A1 (nx10591), .B0 (
           d_arr_add_0__28), .B1 (nx10747), .C0 (d_arr_merge1_0__28), .C1 (
           nx10799)) ;
    latch lat_d_arr_0__29 (.Q (d_arr_0__29), .D (nx8432), .CLK (nx10359)) ;
    nand03 ix8433 (.Y (nx8432), .A0 (nx10110), .A1 (nx10026), .A2 (nx10112)) ;
    aoi22 ix10111 (.Y (nx10110), .A0 (d_arr_merge2_0__29), .A1 (nx10821), .B0 (
          d_arr_relu_0__29), .B1 (nx10843)) ;
    aoi222 ix10113 (.Y (nx10112), .A0 (d_arr_mul_0__29), .A1 (nx10591), .B0 (
           d_arr_add_0__29), .B1 (nx10747), .C0 (d_arr_merge1_0__29), .C1 (
           nx10799)) ;
    latch lat_d_arr_0__30 (.Q (d_arr_0__30), .D (nx8454), .CLK (nx10361)) ;
    nand03 ix8455 (.Y (nx8454), .A0 (nx10116), .A1 (nx10026), .A2 (nx10118)) ;
    aoi22 ix10117 (.Y (nx10116), .A0 (d_arr_merge2_0__30), .A1 (nx10821), .B0 (
          d_arr_relu_0__30), .B1 (nx10843)) ;
    aoi222 ix10119 (.Y (nx10118), .A0 (d_arr_mul_0__30), .A1 (nx10593), .B0 (
           d_arr_add_0__30), .B1 (nx10747), .C0 (d_arr_merge1_0__30), .C1 (
           nx10799)) ;
    latch lat_d_arr_0__31 (.Q (d_arr_0__31), .D (nx8476), .CLK (nx10361)) ;
    nand03 ix8477 (.Y (nx8476), .A0 (nx10122), .A1 (nx10026), .A2 (nx10124)) ;
    aoi22 ix10123 (.Y (nx10122), .A0 (d_arr_merge2_0__31), .A1 (nx10823), .B0 (
          d_arr_relu_0__31), .B1 (nx10843)) ;
    aoi222 ix10125 (.Y (nx10124), .A0 (d_arr_mul_0__31), .A1 (nx10593), .B0 (
           d_arr_add_0__31), .B1 (nx10747), .C0 (d_arr_merge1_0__31), .C1 (
           nx10801)) ;
    inv01 ix5 (.Y (nx4), .A (nx9734)) ;
    inv02 ix10132 (.Y (nx10133), .A (nx10995)) ;
    inv02 ix10134 (.Y (nx10135), .A (nx10995)) ;
    inv02 ix10136 (.Y (nx10137), .A (nx10995)) ;
    inv02 ix10138 (.Y (nx10139), .A (nx10995)) ;
    inv02 ix10140 (.Y (nx10141), .A (nx10995)) ;
    inv02 ix10142 (.Y (nx10143), .A (nx10995)) ;
    inv02 ix10144 (.Y (nx10145), .A (nx10995)) ;
    inv02 ix10146 (.Y (nx10147), .A (nx10883)) ;
    inv02 ix10148 (.Y (nx10149), .A (nx10883)) ;
    inv02 ix10150 (.Y (nx10151), .A (nx10883)) ;
    inv02 ix10152 (.Y (nx10153), .A (nx10883)) ;
    inv02 ix10154 (.Y (nx10155), .A (nx10883)) ;
    inv02 ix10156 (.Y (nx10157), .A (nx10883)) ;
    inv02 ix10158 (.Y (nx10159), .A (nx10883)) ;
    inv02 ix10160 (.Y (nx10161), .A (nx10885)) ;
    inv02 ix10162 (.Y (nx10163), .A (nx10885)) ;
    inv02 ix10164 (.Y (nx10165), .A (nx10885)) ;
    inv02 ix10166 (.Y (nx10167), .A (nx10885)) ;
    inv02 ix10168 (.Y (nx10169), .A (nx10885)) ;
    inv02 ix10170 (.Y (nx10171), .A (nx10885)) ;
    inv02 ix10172 (.Y (nx10173), .A (nx10885)) ;
    inv02 ix10174 (.Y (nx10175), .A (nx10887)) ;
    inv02 ix10176 (.Y (nx10177), .A (nx10887)) ;
    inv02 ix10178 (.Y (nx10179), .A (nx10887)) ;
    inv02 ix10180 (.Y (nx10181), .A (nx10887)) ;
    inv02 ix10182 (.Y (nx10183), .A (nx10887)) ;
    inv02 ix10184 (.Y (nx10185), .A (nx10887)) ;
    inv02 ix10186 (.Y (nx10187), .A (nx10887)) ;
    inv02 ix10188 (.Y (nx10189), .A (nx10889)) ;
    inv02 ix10190 (.Y (nx10191), .A (nx10889)) ;
    inv02 ix10192 (.Y (nx10193), .A (nx10889)) ;
    inv02 ix10194 (.Y (nx10195), .A (nx10889)) ;
    inv02 ix10196 (.Y (nx10197), .A (nx10889)) ;
    inv02 ix10198 (.Y (nx10199), .A (nx10889)) ;
    inv02 ix10200 (.Y (nx10201), .A (nx10889)) ;
    inv02 ix10202 (.Y (nx10203), .A (nx10891)) ;
    inv02 ix10204 (.Y (nx10205), .A (nx10891)) ;
    inv02 ix10206 (.Y (nx10207), .A (nx10891)) ;
    inv02 ix10208 (.Y (nx10209), .A (nx10891)) ;
    inv02 ix10210 (.Y (nx10211), .A (nx10891)) ;
    inv02 ix10212 (.Y (nx10213), .A (nx10891)) ;
    inv02 ix10214 (.Y (nx10215), .A (nx10891)) ;
    inv02 ix10216 (.Y (nx10217), .A (nx10893)) ;
    inv02 ix10218 (.Y (nx10219), .A (nx10893)) ;
    inv02 ix10220 (.Y (nx10221), .A (nx10893)) ;
    inv02 ix10222 (.Y (nx10223), .A (nx10893)) ;
    inv02 ix10224 (.Y (nx10225), .A (nx10893)) ;
    inv02 ix10226 (.Y (nx10227), .A (nx10893)) ;
    inv02 ix10228 (.Y (nx10229), .A (nx10893)) ;
    inv02 ix10230 (.Y (nx10231), .A (nx10895)) ;
    inv02 ix10232 (.Y (nx10233), .A (nx10895)) ;
    inv02 ix10234 (.Y (nx10235), .A (nx10895)) ;
    inv02 ix10236 (.Y (nx10237), .A (nx10895)) ;
    inv02 ix10238 (.Y (nx10239), .A (nx10895)) ;
    inv02 ix10240 (.Y (nx10241), .A (nx10895)) ;
    inv02 ix10242 (.Y (nx10243), .A (nx10895)) ;
    inv02 ix10244 (.Y (nx10245), .A (nx10897)) ;
    inv02 ix10246 (.Y (nx10247), .A (nx10897)) ;
    inv02 ix10248 (.Y (nx10249), .A (nx10897)) ;
    inv02 ix10250 (.Y (nx10251), .A (nx10897)) ;
    inv02 ix10252 (.Y (nx10253), .A (nx10897)) ;
    inv02 ix10254 (.Y (nx10255), .A (nx10897)) ;
    inv02 ix10256 (.Y (nx10257), .A (nx10897)) ;
    inv02 ix10258 (.Y (nx10259), .A (nx10899)) ;
    inv02 ix10260 (.Y (nx10261), .A (nx10899)) ;
    inv02 ix10262 (.Y (nx10263), .A (nx10899)) ;
    inv02 ix10264 (.Y (nx10265), .A (nx10899)) ;
    inv02 ix10266 (.Y (nx10267), .A (nx10899)) ;
    inv02 ix10268 (.Y (nx10269), .A (nx10899)) ;
    inv02 ix10270 (.Y (nx10271), .A (nx10899)) ;
    inv02 ix10272 (.Y (nx10273), .A (nx10901)) ;
    inv02 ix10274 (.Y (nx10275), .A (nx10901)) ;
    inv02 ix10276 (.Y (nx10277), .A (nx10901)) ;
    inv02 ix10278 (.Y (nx10279), .A (nx10901)) ;
    inv02 ix10280 (.Y (nx10281), .A (nx10901)) ;
    inv02 ix10282 (.Y (nx10283), .A (nx10901)) ;
    inv02 ix10284 (.Y (nx10285), .A (nx10901)) ;
    inv02 ix10286 (.Y (nx10287), .A (nx10903)) ;
    inv02 ix10288 (.Y (nx10289), .A (nx10903)) ;
    inv02 ix10290 (.Y (nx10291), .A (nx10903)) ;
    inv02 ix10292 (.Y (nx10293), .A (nx10903)) ;
    inv02 ix10294 (.Y (nx10295), .A (nx10903)) ;
    inv02 ix10296 (.Y (nx10297), .A (nx10903)) ;
    inv02 ix10298 (.Y (nx10299), .A (nx10903)) ;
    inv02 ix10300 (.Y (nx10301), .A (nx10905)) ;
    inv02 ix10302 (.Y (nx10303), .A (nx10905)) ;
    inv02 ix10304 (.Y (nx10305), .A (nx10905)) ;
    inv02 ix10306 (.Y (nx10307), .A (nx10905)) ;
    inv02 ix10308 (.Y (nx10309), .A (nx10905)) ;
    inv02 ix10310 (.Y (nx10311), .A (nx10905)) ;
    inv02 ix10312 (.Y (nx10313), .A (nx10905)) ;
    inv02 ix10314 (.Y (nx10315), .A (nx10907)) ;
    inv02 ix10316 (.Y (nx10317), .A (nx10907)) ;
    inv02 ix10318 (.Y (nx10319), .A (nx10907)) ;
    inv02 ix10320 (.Y (nx10321), .A (nx10907)) ;
    inv02 ix10322 (.Y (nx10323), .A (nx10907)) ;
    inv02 ix10324 (.Y (nx10325), .A (nx10907)) ;
    inv02 ix10326 (.Y (nx10327), .A (nx10907)) ;
    inv02 ix10328 (.Y (nx10329), .A (nx10909)) ;
    inv02 ix10330 (.Y (nx10331), .A (nx10909)) ;
    inv02 ix10332 (.Y (nx10333), .A (nx10909)) ;
    inv02 ix10334 (.Y (nx10335), .A (nx10909)) ;
    inv02 ix10336 (.Y (nx10337), .A (nx10909)) ;
    inv02 ix10338 (.Y (nx10339), .A (nx10909)) ;
    inv02 ix10340 (.Y (nx10341), .A (nx10909)) ;
    inv02 ix10342 (.Y (nx10343), .A (nx10911)) ;
    inv02 ix10344 (.Y (nx10345), .A (nx10911)) ;
    inv02 ix10346 (.Y (nx10347), .A (nx10911)) ;
    inv02 ix10348 (.Y (nx10349), .A (nx10911)) ;
    inv02 ix10350 (.Y (nx10351), .A (nx10911)) ;
    inv02 ix10352 (.Y (nx10353), .A (nx10911)) ;
    inv02 ix10354 (.Y (nx10355), .A (nx10911)) ;
    inv02 ix10356 (.Y (nx10357), .A (nx10913)) ;
    inv02 ix10358 (.Y (nx10359), .A (nx10913)) ;
    inv02 ix10360 (.Y (nx10361), .A (nx10913)) ;
    inv02 ix10364 (.Y (nx10365), .A (nx11471)) ;
    inv02 ix10366 (.Y (nx10367), .A (nx11471)) ;
    inv02 ix10368 (.Y (nx10369), .A (nx11471)) ;
    inv02 ix10372 (.Y (nx10373), .A (nx11471)) ;
    inv02 ix10374 (.Y (nx10375), .A (nx11471)) ;
    inv02 ix10376 (.Y (nx10377), .A (nx11471)) ;
    inv02 ix10382 (.Y (nx10383), .A (nx11435)) ;
    inv02 ix10384 (.Y (nx10385), .A (nx11435)) ;
    inv02 ix10386 (.Y (nx10387), .A (nx11435)) ;
    inv02 ix10390 (.Y (nx10391), .A (nx11435)) ;
    inv02 ix10392 (.Y (nx10393), .A (nx10919)) ;
    inv02 ix10394 (.Y (nx10395), .A (nx10919)) ;
    inv02 ix10396 (.Y (nx10397), .A (nx10919)) ;
    inv02 ix10398 (.Y (nx10399), .A (nx10919)) ;
    inv02 ix10400 (.Y (nx10401), .A (nx10919)) ;
    inv02 ix10402 (.Y (nx10403), .A (nx10919)) ;
    inv02 ix10404 (.Y (nx10405), .A (nx10919)) ;
    inv02 ix10406 (.Y (nx10407), .A (nx10921)) ;
    inv02 ix10408 (.Y (nx10409), .A (nx10921)) ;
    inv02 ix10410 (.Y (nx10411), .A (nx10921)) ;
    inv02 ix10412 (.Y (nx10413), .A (nx10921)) ;
    inv02 ix10414 (.Y (nx10415), .A (nx10921)) ;
    inv02 ix10416 (.Y (nx10417), .A (nx10921)) ;
    inv02 ix10418 (.Y (nx10419), .A (nx10921)) ;
    inv02 ix10420 (.Y (nx10421), .A (nx10923)) ;
    inv02 ix10422 (.Y (nx10423), .A (nx10923)) ;
    inv02 ix10424 (.Y (nx10425), .A (nx10923)) ;
    inv02 ix10426 (.Y (nx10427), .A (nx10923)) ;
    inv02 ix10428 (.Y (nx10429), .A (nx10923)) ;
    inv02 ix10430 (.Y (nx10431), .A (nx10923)) ;
    inv02 ix10432 (.Y (nx10433), .A (nx10923)) ;
    inv02 ix10434 (.Y (nx10435), .A (nx10925)) ;
    inv02 ix10436 (.Y (nx10437), .A (nx10925)) ;
    inv02 ix10438 (.Y (nx10439), .A (nx10925)) ;
    inv02 ix10440 (.Y (nx10441), .A (nx10925)) ;
    inv02 ix10442 (.Y (nx10443), .A (nx10925)) ;
    inv02 ix10444 (.Y (nx10445), .A (nx10925)) ;
    inv02 ix10446 (.Y (nx10447), .A (nx10925)) ;
    inv02 ix10448 (.Y (nx10449), .A (nx10927)) ;
    inv02 ix10450 (.Y (nx10451), .A (nx10927)) ;
    inv02 ix10452 (.Y (nx10453), .A (nx10927)) ;
    inv02 ix10454 (.Y (nx10455), .A (nx10927)) ;
    inv02 ix10456 (.Y (nx10457), .A (nx10927)) ;
    inv02 ix10458 (.Y (nx10459), .A (nx10927)) ;
    inv02 ix10460 (.Y (nx10461), .A (nx10927)) ;
    inv02 ix10462 (.Y (nx10463), .A (nx10929)) ;
    inv02 ix10464 (.Y (nx10465), .A (nx10929)) ;
    inv02 ix10466 (.Y (nx10467), .A (nx10929)) ;
    inv02 ix10468 (.Y (nx10469), .A (nx10929)) ;
    inv02 ix10470 (.Y (nx10471), .A (nx10929)) ;
    inv02 ix10472 (.Y (nx10473), .A (nx10929)) ;
    inv02 ix10474 (.Y (nx10475), .A (nx10929)) ;
    inv02 ix10476 (.Y (nx10477), .A (nx10931)) ;
    inv02 ix10478 (.Y (nx10479), .A (nx10931)) ;
    inv02 ix10480 (.Y (nx10481), .A (nx10931)) ;
    inv02 ix10482 (.Y (nx10483), .A (nx10931)) ;
    inv02 ix10484 (.Y (nx10485), .A (nx10931)) ;
    inv02 ix10486 (.Y (nx10487), .A (nx10931)) ;
    inv02 ix10488 (.Y (nx10489), .A (nx10931)) ;
    inv02 ix10490 (.Y (nx10491), .A (nx10933)) ;
    inv02 ix10492 (.Y (nx10493), .A (nx10933)) ;
    inv02 ix10494 (.Y (nx10495), .A (nx10933)) ;
    inv02 ix10496 (.Y (nx10497), .A (nx10933)) ;
    inv02 ix10498 (.Y (nx10499), .A (nx10933)) ;
    inv02 ix10500 (.Y (nx10501), .A (nx10933)) ;
    inv02 ix10502 (.Y (nx10503), .A (nx10933)) ;
    inv02 ix10504 (.Y (nx10505), .A (nx11445)) ;
    inv02 ix10506 (.Y (nx10507), .A (nx11445)) ;
    inv02 ix10508 (.Y (nx10509), .A (nx11445)) ;
    inv02 ix10510 (.Y (nx10511), .A (nx11445)) ;
    inv02 ix10512 (.Y (nx10513), .A (nx11445)) ;
    inv02 ix10514 (.Y (nx10515), .A (nx11445)) ;
    inv02 ix10518 (.Y (nx10519), .A (nx11449)) ;
    inv02 ix10520 (.Y (nx10521), .A (nx11449)) ;
    inv02 ix10522 (.Y (nx10523), .A (nx11449)) ;
    inv02 ix10528 (.Y (nx10529), .A (nx11449)) ;
    inv02 ix10530 (.Y (nx10531), .A (nx11449)) ;
    inv02 ix10532 (.Y (nx10533), .A (nx11455)) ;
    inv02 ix10536 (.Y (nx10537), .A (nx11455)) ;
    inv02 ix10538 (.Y (nx10539), .A (nx11455)) ;
    inv02 ix10540 (.Y (nx10541), .A (nx11455)) ;
    inv02 ix10546 (.Y (nx10547), .A (nx11463)) ;
    inv02 ix10548 (.Y (nx10549), .A (nx11463)) ;
    inv02 ix10550 (.Y (nx10551), .A (nx11463)) ;
    inv02 ix10552 (.Y (nx10553), .A (nx11463)) ;
    inv02 ix10554 (.Y (nx10555), .A (nx11463)) ;
    inv02 ix10556 (.Y (nx10557), .A (nx11463)) ;
    inv02 ix10558 (.Y (nx10559), .A (nx11463)) ;
    inv02 ix10560 (.Y (nx10561), .A (nx10943)) ;
    inv02 ix10562 (.Y (nx10563), .A (nx10943)) ;
    inv02 ix10564 (.Y (nx10565), .A (nx10943)) ;
    inv02 ix10566 (.Y (nx10567), .A (nx10943)) ;
    inv02 ix10568 (.Y (nx10569), .A (nx10943)) ;
    inv02 ix10570 (.Y (nx10571), .A (nx10943)) ;
    inv02 ix10572 (.Y (nx10573), .A (nx10943)) ;
    inv02 ix10574 (.Y (nx10575), .A (nx10945)) ;
    inv02 ix10576 (.Y (nx10577), .A (nx10945)) ;
    inv02 ix10578 (.Y (nx10579), .A (nx10945)) ;
    inv02 ix10580 (.Y (nx10581), .A (nx10945)) ;
    inv02 ix10582 (.Y (nx10583), .A (nx10945)) ;
    inv02 ix10584 (.Y (nx10585), .A (nx10945)) ;
    inv02 ix10586 (.Y (nx10587), .A (nx10945)) ;
    inv02 ix10588 (.Y (nx10589), .A (nx10947)) ;
    inv02 ix10590 (.Y (nx10591), .A (nx10947)) ;
    inv02 ix10592 (.Y (nx10593), .A (nx10947)) ;
    inv02 ix10620 (.Y (nx10621), .A (nx10999)) ;
    inv02 ix10622 (.Y (nx10623), .A (nx10999)) ;
    inv02 ix10624 (.Y (nx10625), .A (nx10999)) ;
    inv02 ix10626 (.Y (nx10627), .A (nx10999)) ;
    inv02 ix10628 (.Y (nx10629), .A (nx10999)) ;
    inv02 ix10630 (.Y (nx10631), .A (nx10999)) ;
    inv02 ix10632 (.Y (nx10633), .A (nx10949)) ;
    inv02 ix10634 (.Y (nx10635), .A (nx10951)) ;
    inv02 ix10636 (.Y (nx10637), .A (nx10951)) ;
    inv02 ix10638 (.Y (nx10639), .A (nx10951)) ;
    inv02 ix10640 (.Y (nx10641), .A (nx10951)) ;
    inv02 ix10642 (.Y (nx10643), .A (nx10951)) ;
    inv02 ix10644 (.Y (nx10645), .A (nx10951)) ;
    inv02 ix10646 (.Y (nx10647), .A (nx10951)) ;
    inv02 ix10648 (.Y (nx10649), .A (nx10953)) ;
    inv02 ix10650 (.Y (nx10651), .A (nx10953)) ;
    inv02 ix10652 (.Y (nx10653), .A (nx10953)) ;
    inv02 ix10654 (.Y (nx10655), .A (nx10953)) ;
    inv02 ix10656 (.Y (nx10657), .A (nx10953)) ;
    inv02 ix10658 (.Y (nx10659), .A (nx10953)) ;
    inv02 ix10660 (.Y (nx10661), .A (nx10953)) ;
    inv02 ix10662 (.Y (nx10663), .A (nx10955)) ;
    inv02 ix10664 (.Y (nx10665), .A (nx10955)) ;
    inv02 ix10666 (.Y (nx10667), .A (nx10955)) ;
    inv02 ix10668 (.Y (nx10669), .A (nx10955)) ;
    inv02 ix10670 (.Y (nx10671), .A (nx10955)) ;
    inv02 ix10672 (.Y (nx10673), .A (nx10955)) ;
    inv02 ix10674 (.Y (nx10675), .A (nx10955)) ;
    inv02 ix10676 (.Y (nx10677), .A (nx10957)) ;
    inv02 ix10678 (.Y (nx10679), .A (nx10957)) ;
    inv02 ix10680 (.Y (nx10681), .A (nx10957)) ;
    inv02 ix10682 (.Y (nx10683), .A (nx10957)) ;
    inv02 ix10684 (.Y (nx10685), .A (nx10957)) ;
    inv02 ix10686 (.Y (nx10687), .A (nx10957)) ;
    inv02 ix10688 (.Y (nx10689), .A (nx10957)) ;
    inv02 ix10690 (.Y (nx10691), .A (nx10959)) ;
    inv02 ix10692 (.Y (nx10693), .A (nx10959)) ;
    inv02 ix10694 (.Y (nx10695), .A (nx10959)) ;
    inv02 ix10696 (.Y (nx10697), .A (nx10959)) ;
    inv02 ix10698 (.Y (nx10699), .A (nx10959)) ;
    inv02 ix10700 (.Y (nx10701), .A (nx10959)) ;
    inv02 ix10702 (.Y (nx10703), .A (nx10959)) ;
    inv02 ix10704 (.Y (nx10705), .A (nx10961)) ;
    inv02 ix10706 (.Y (nx10707), .A (nx10961)) ;
    inv02 ix10708 (.Y (nx10709), .A (nx10961)) ;
    inv02 ix10710 (.Y (nx10711), .A (nx10961)) ;
    inv02 ix10712 (.Y (nx10713), .A (nx10961)) ;
    inv02 ix10714 (.Y (nx10715), .A (nx10961)) ;
    inv02 ix10716 (.Y (nx10717), .A (nx10961)) ;
    inv02 ix10718 (.Y (nx10719), .A (nx10963)) ;
    inv02 ix10720 (.Y (nx10721), .A (nx10963)) ;
    inv02 ix10722 (.Y (nx10723), .A (nx10963)) ;
    inv02 ix10724 (.Y (nx10725), .A (nx10963)) ;
    inv02 ix10726 (.Y (nx10727), .A (nx10963)) ;
    inv02 ix10728 (.Y (nx10729), .A (nx10963)) ;
    inv02 ix10730 (.Y (nx10731), .A (nx10963)) ;
    inv02 ix10732 (.Y (nx10733), .A (nx10965)) ;
    inv02 ix10734 (.Y (nx10735), .A (nx10965)) ;
    inv02 ix10736 (.Y (nx10737), .A (nx10965)) ;
    inv02 ix10738 (.Y (nx10739), .A (nx10965)) ;
    inv02 ix10740 (.Y (nx10741), .A (nx10965)) ;
    inv02 ix10742 (.Y (nx10743), .A (nx10965)) ;
    inv02 ix10744 (.Y (nx10745), .A (nx10965)) ;
    inv02 ix10746 (.Y (nx10747), .A (nx10967)) ;
    inv01 ix10780 (.Y (nx10781), .A (nx7002)) ;
    inv02 ix10782 (.Y (nx10783), .A (nx10969)) ;
    inv02 ix10784 (.Y (nx10785), .A (nx10969)) ;
    inv02 ix10786 (.Y (nx10787), .A (nx10969)) ;
    inv02 ix10788 (.Y (nx10789), .A (nx10969)) ;
    inv02 ix10790 (.Y (nx10791), .A (nx10969)) ;
    inv02 ix10792 (.Y (nx10793), .A (nx10781)) ;
    inv02 ix10794 (.Y (nx10795), .A (nx10781)) ;
    inv02 ix10796 (.Y (nx10797), .A (nx10781)) ;
    inv02 ix10798 (.Y (nx10799), .A (nx10781)) ;
    inv02 ix10800 (.Y (nx10801), .A (nx10781)) ;
    inv01 ix10802 (.Y (nx10803), .A (nx7018)) ;
    inv02 ix10804 (.Y (nx10805), .A (nx10971)) ;
    inv02 ix10806 (.Y (nx10807), .A (nx10971)) ;
    inv02 ix10808 (.Y (nx10809), .A (nx10971)) ;
    inv02 ix10810 (.Y (nx10811), .A (nx10971)) ;
    inv02 ix10812 (.Y (nx10813), .A (nx10971)) ;
    inv02 ix10814 (.Y (nx10815), .A (nx10803)) ;
    inv02 ix10816 (.Y (nx10817), .A (nx10803)) ;
    inv02 ix10818 (.Y (nx10819), .A (nx10803)) ;
    inv02 ix10820 (.Y (nx10821), .A (nx10803)) ;
    inv02 ix10822 (.Y (nx10823), .A (nx10803)) ;
    inv01 ix10824 (.Y (nx10825), .A (nx7028)) ;
    inv02 ix10826 (.Y (nx10827), .A (nx10973)) ;
    inv02 ix10828 (.Y (nx10829), .A (nx10973)) ;
    inv02 ix10830 (.Y (nx10831), .A (nx10973)) ;
    inv02 ix10832 (.Y (nx10833), .A (nx10973)) ;
    inv02 ix10834 (.Y (nx10835), .A (nx10973)) ;
    inv02 ix10836 (.Y (nx10837), .A (nx10825)) ;
    inv02 ix10838 (.Y (nx10839), .A (nx10825)) ;
    inv02 ix10840 (.Y (nx10841), .A (nx10825)) ;
    inv02 ix10842 (.Y (nx10843), .A (nx10825)) ;
    nand02 ix10844 (.Y (nx10845), .A0 (d_arr_mux_21__31), .A1 (nx11399)) ;
    nand02 ix10846 (.Y (nx10847), .A0 (d_arr_mux_21__31), .A1 (nx11399)) ;
    nand02 ix10848 (.Y (nx10849), .A0 (d_arr_mux_20__31), .A1 (nx11399)) ;
    nand02 ix10850 (.Y (nx10851), .A0 (d_arr_mux_20__31), .A1 (nx11399)) ;
    nand02 ix10852 (.Y (nx10853), .A0 (d_arr_mux_19__31), .A1 (nx11399)) ;
    nand02 ix10854 (.Y (nx10855), .A0 (d_arr_mux_19__31), .A1 (nx11401)) ;
    nand02 ix10856 (.Y (nx10857), .A0 (d_arr_mux_18__31), .A1 (nx11401)) ;
    nand02 ix10858 (.Y (nx10859), .A0 (d_arr_mux_18__31), .A1 (nx11401)) ;
    nand02 ix10860 (.Y (nx10861), .A0 (d_arr_mux_4__31), .A1 (nx11401)) ;
    nand02 ix10862 (.Y (nx10863), .A0 (d_arr_mux_4__31), .A1 (nx11401)) ;
    nand02 ix10864 (.Y (nx10865), .A0 (d_arr_mux_3__31), .A1 (nx11401)) ;
    nand02 ix10866 (.Y (nx10867), .A0 (d_arr_mux_3__31), .A1 (nx11401)) ;
    nand02 ix10868 (.Y (nx10869), .A0 (d_arr_mux_2__31), .A1 (nx11501)) ;
    nand02 ix10870 (.Y (nx10871), .A0 (d_arr_mux_2__31), .A1 (nx11501)) ;
    nand02 ix10872 (.Y (nx10873), .A0 (d_arr_mux_1__31), .A1 (nx11501)) ;
    nand02 ix10874 (.Y (nx10875), .A0 (d_arr_mux_1__31), .A1 (nx11501)) ;
    nand02 ix10876 (.Y (nx10877), .A0 (d_arr_mux_0__31), .A1 (nx11501)) ;
    nand02 ix10878 (.Y (nx10879), .A0 (d_arr_mux_0__31), .A1 (nx11501)) ;
    inv02 ix10880 (.Y (nx10881), .A (nx8)) ;
    inv02 ix10882 (.Y (nx10883), .A (nx10979)) ;
    inv02 ix10884 (.Y (nx10885), .A (nx10979)) ;
    inv02 ix10886 (.Y (nx10887), .A (nx10979)) ;
    inv02 ix10888 (.Y (nx10889), .A (nx10979)) ;
    inv02 ix10890 (.Y (nx10891), .A (nx10979)) ;
    inv02 ix10892 (.Y (nx10893), .A (nx10979)) ;
    inv02 ix10894 (.Y (nx10895), .A (nx10979)) ;
    inv02 ix10896 (.Y (nx10897), .A (nx10981)) ;
    inv02 ix10898 (.Y (nx10899), .A (nx10981)) ;
    inv02 ix10900 (.Y (nx10901), .A (nx10981)) ;
    inv02 ix10902 (.Y (nx10903), .A (nx10981)) ;
    inv02 ix10904 (.Y (nx10905), .A (nx10981)) ;
    inv02 ix10906 (.Y (nx10907), .A (nx10981)) ;
    inv02 ix10908 (.Y (nx10909), .A (nx10981)) ;
    inv02 ix10910 (.Y (nx10911), .A (nx10983)) ;
    inv02 ix10912 (.Y (nx10913), .A (nx10983)) ;
    inv02 ix10914 (.Y (nx10915), .A (nx12)) ;
    inv02 ix10916 (.Y (nx10917), .A (nx11465)) ;
    inv02 ix10918 (.Y (nx10919), .A (nx11465)) ;
    inv02 ix10920 (.Y (nx10921), .A (nx11465)) ;
    inv02 ix10922 (.Y (nx10923), .A (nx11465)) ;
    inv02 ix10924 (.Y (nx10925), .A (nx11465)) ;
    inv02 ix10926 (.Y (nx10927), .A (nx11465)) ;
    inv02 ix10928 (.Y (nx10929), .A (nx11465)) ;
    inv02 ix10930 (.Y (nx10931), .A (nx11467)) ;
    inv02 ix10932 (.Y (nx10933), .A (nx11467)) ;
    inv02 ix10934 (.Y (nx10935), .A (nx11467)) ;
    inv02 ix10936 (.Y (nx10937), .A (nx11467)) ;
    inv02 ix10938 (.Y (nx10939), .A (nx11467)) ;
    inv02 ix10940 (.Y (nx10941), .A (nx11467)) ;
    inv02 ix10942 (.Y (nx10943), .A (nx11467)) ;
    inv02 ix10944 (.Y (nx10945), .A (nx10989)) ;
    inv02 ix10946 (.Y (nx10947), .A (nx10989)) ;
    inv02 ix10948 (.Y (nx10949), .A (nx694)) ;
    inv02 ix10950 (.Y (nx10951), .A (nx10991)) ;
    inv02 ix10952 (.Y (nx10953), .A (nx10991)) ;
    inv02 ix10954 (.Y (nx10955), .A (nx10991)) ;
    inv02 ix10956 (.Y (nx10957), .A (nx10991)) ;
    inv02 ix10958 (.Y (nx10959), .A (nx10991)) ;
    inv02 ix10960 (.Y (nx10961), .A (nx10993)) ;
    inv02 ix10962 (.Y (nx10963), .A (nx10993)) ;
    inv02 ix10964 (.Y (nx10965), .A (nx10993)) ;
    inv02 ix10966 (.Y (nx10967), .A (nx10993)) ;
    inv01 ix10968 (.Y (nx10969), .A (nx7002)) ;
    inv01 ix10970 (.Y (nx10971), .A (nx7018)) ;
    inv01 ix10972 (.Y (nx10973), .A (nx7028)) ;
    inv02 ix10978 (.Y (nx10979), .A (nx10881)) ;
    inv02 ix10980 (.Y (nx10981), .A (nx10881)) ;
    inv02 ix10982 (.Y (nx10983), .A (nx10881)) ;
    inv02 ix10984 (.Y (nx10985), .A (nx10915)) ;
    inv02 ix10986 (.Y (nx10987), .A (nx10915)) ;
    inv02 ix10988 (.Y (nx10989), .A (nx10915)) ;
    inv01 ix10990 (.Y (nx10991), .A (nx10999)) ;
    inv01 ix10992 (.Y (nx10993), .A (nx10949)) ;
    inv02 ix10994 (.Y (nx10995), .A (nx8)) ;
    inv02 ix10996 (.Y (nx10997), .A (nx11511)) ;
    inv02 ix10998 (.Y (nx10999), .A (nx694)) ;
    oai21 ix141 (.Y (nx140), .A0 (nx11005), .A1 (nx11471), .B0 (nx11407)) ;
    inv01 ix11004 (.Y (nx11005), .A (d_arr_mul_24__15)) ;
    nand02 ix137 (.Y (nx10595), .A0 (nx11501), .A1 (d_arr_mux_24__31)) ;
    oai21 ix147 (.Y (nx146), .A0 (nx11007), .A1 (nx11473), .B0 (nx11407)) ;
    inv01 ix11006 (.Y (nx11007), .A (d_arr_mul_24__16)) ;
    oai21 ix153 (.Y (nx152), .A0 (nx11009), .A1 (nx11473), .B0 (nx11407)) ;
    inv01 ix11008 (.Y (nx11009), .A (d_arr_mul_24__17)) ;
    oai21 ix159 (.Y (nx158), .A0 (nx11011), .A1 (nx11473), .B0 (nx11407)) ;
    inv01 ix11010 (.Y (nx11011), .A (d_arr_mul_24__18)) ;
    oai21 ix165 (.Y (nx164), .A0 (nx11013), .A1 (nx11473), .B0 (nx11407)) ;
    inv01 ix11012 (.Y (nx11013), .A (d_arr_mul_24__19)) ;
    oai21 ix171 (.Y (nx170), .A0 (nx11015), .A1 (nx11473), .B0 (nx11407)) ;
    inv01 ix11014 (.Y (nx11015), .A (d_arr_mul_24__20)) ;
    oai21 ix177 (.Y (nx176), .A0 (nx11017), .A1 (nx11473), .B0 (nx11407)) ;
    inv01 ix11016 (.Y (nx11017), .A (d_arr_mul_24__21)) ;
    oai21 ix183 (.Y (nx182), .A0 (nx11019), .A1 (nx11473), .B0 (nx11409)) ;
    inv01 ix11018 (.Y (nx11019), .A (d_arr_mul_24__22)) ;
    oai21 ix189 (.Y (nx188), .A0 (nx11021), .A1 (nx11475), .B0 (nx11409)) ;
    inv01 ix11020 (.Y (nx11021), .A (d_arr_mul_24__23)) ;
    oai21 ix195 (.Y (nx194), .A0 (nx11023), .A1 (nx11475), .B0 (nx11409)) ;
    inv01 ix11022 (.Y (nx11023), .A (d_arr_mul_24__24)) ;
    oai21 ix201 (.Y (nx200), .A0 (nx11025), .A1 (nx11475), .B0 (nx11409)) ;
    inv01 ix11024 (.Y (nx11025), .A (d_arr_mul_24__25)) ;
    oai21 ix207 (.Y (nx206), .A0 (nx11027), .A1 (nx11475), .B0 (nx11409)) ;
    inv01 ix11026 (.Y (nx11027), .A (d_arr_mul_24__26)) ;
    oai21 ix213 (.Y (nx212), .A0 (nx11029), .A1 (nx11475), .B0 (nx11409)) ;
    inv01 ix11028 (.Y (nx11029), .A (d_arr_mul_24__27)) ;
    oai21 ix219 (.Y (nx218), .A0 (nx11031), .A1 (nx11475), .B0 (nx11409)) ;
    inv01 ix11030 (.Y (nx11031), .A (d_arr_mul_24__28)) ;
    oai21 ix225 (.Y (nx224), .A0 (nx11033), .A1 (nx11475), .B0 (nx10595)) ;
    inv01 ix11032 (.Y (nx11033), .A (d_arr_mul_24__29)) ;
    oai21 ix231 (.Y (nx230), .A0 (nx11035), .A1 (nx10997), .B0 (nx10595)) ;
    inv01 ix11034 (.Y (nx11035), .A (d_arr_mul_24__30)) ;
    oai21 ix237 (.Y (nx236), .A0 (nx11037), .A1 (nx10997), .B0 (nx10595)) ;
    inv01 ix11036 (.Y (nx11037), .A (d_arr_mul_24__31)) ;
    oai21 ix365 (.Y (nx364), .A0 (nx11039), .A1 (nx10997), .B0 (nx11411)) ;
    inv01 ix11038 (.Y (nx11039), .A (d_arr_mul_23__15)) ;
    nand02 ix361 (.Y (nx10603), .A0 (nx11503), .A1 (d_arr_mux_23__31)) ;
    oai21 ix371 (.Y (nx370), .A0 (nx11041), .A1 (nx10997), .B0 (nx11411)) ;
    inv01 ix11040 (.Y (nx11041), .A (d_arr_mul_23__16)) ;
    oai21 ix377 (.Y (nx376), .A0 (nx11043), .A1 (nx11435), .B0 (nx11411)) ;
    inv01 ix11042 (.Y (nx11043), .A (d_arr_mul_23__17)) ;
    oai21 ix383 (.Y (nx382), .A0 (nx11045), .A1 (nx11435), .B0 (nx11411)) ;
    inv01 ix11044 (.Y (nx11045), .A (d_arr_mul_23__18)) ;
    oai21 ix389 (.Y (nx388), .A0 (nx11047), .A1 (nx11435), .B0 (nx11411)) ;
    inv01 ix11046 (.Y (nx11047), .A (d_arr_mul_23__19)) ;
    oai21 ix395 (.Y (nx394), .A0 (nx11049), .A1 (nx11437), .B0 (nx11411)) ;
    inv01 ix11048 (.Y (nx11049), .A (d_arr_mul_23__20)) ;
    oai21 ix401 (.Y (nx400), .A0 (nx11051), .A1 (nx11437), .B0 (nx11411)) ;
    inv01 ix11050 (.Y (nx11051), .A (d_arr_mul_23__21)) ;
    oai21 ix407 (.Y (nx406), .A0 (nx11053), .A1 (nx11437), .B0 (nx11413)) ;
    inv01 ix11052 (.Y (nx11053), .A (d_arr_mul_23__22)) ;
    oai21 ix413 (.Y (nx412), .A0 (nx11055), .A1 (nx11437), .B0 (nx11413)) ;
    inv01 ix11054 (.Y (nx11055), .A (d_arr_mul_23__23)) ;
    oai21 ix419 (.Y (nx418), .A0 (nx11057), .A1 (nx11437), .B0 (nx11413)) ;
    inv01 ix11056 (.Y (nx11057), .A (d_arr_mul_23__24)) ;
    oai21 ix425 (.Y (nx424), .A0 (nx11059), .A1 (nx11437), .B0 (nx11413)) ;
    inv01 ix11058 (.Y (nx11059), .A (d_arr_mul_23__25)) ;
    oai21 ix431 (.Y (nx430), .A0 (nx11061), .A1 (nx11437), .B0 (nx11413)) ;
    inv01 ix11060 (.Y (nx11061), .A (d_arr_mul_23__26)) ;
    oai21 ix437 (.Y (nx436), .A0 (nx11063), .A1 (nx11439), .B0 (nx11413)) ;
    inv01 ix11062 (.Y (nx11063), .A (d_arr_mul_23__27)) ;
    oai21 ix443 (.Y (nx442), .A0 (nx11065), .A1 (nx11439), .B0 (nx11413)) ;
    inv01 ix11064 (.Y (nx11065), .A (d_arr_mul_23__28)) ;
    oai21 ix449 (.Y (nx448), .A0 (nx11067), .A1 (nx11439), .B0 (nx10603)) ;
    inv01 ix11066 (.Y (nx11067), .A (d_arr_mul_23__29)) ;
    oai21 ix455 (.Y (nx454), .A0 (nx11069), .A1 (nx11439), .B0 (nx10603)) ;
    inv01 ix11068 (.Y (nx11069), .A (d_arr_mul_23__30)) ;
    oai21 ix461 (.Y (nx460), .A0 (nx11071), .A1 (nx11439), .B0 (nx10603)) ;
    inv01 ix11070 (.Y (nx11071), .A (d_arr_mul_23__31)) ;
    oai21 ix589 (.Y (nx588), .A0 (nx11073), .A1 (nx11439), .B0 (nx11415)) ;
    inv01 ix11072 (.Y (nx11073), .A (d_arr_mul_22__15)) ;
    nand02 ix585 (.Y (nx10611), .A0 (nx11503), .A1 (d_arr_mux_22__31)) ;
    oai21 ix595 (.Y (nx594), .A0 (nx11075), .A1 (nx11439), .B0 (nx11415)) ;
    inv01 ix11074 (.Y (nx11075), .A (d_arr_mul_22__16)) ;
    oai21 ix601 (.Y (nx600), .A0 (nx11077), .A1 (nx11441), .B0 (nx11415)) ;
    inv01 ix11076 (.Y (nx11077), .A (d_arr_mul_22__17)) ;
    oai21 ix607 (.Y (nx606), .A0 (nx11079), .A1 (nx11441), .B0 (nx11415)) ;
    inv01 ix11078 (.Y (nx11079), .A (d_arr_mul_22__18)) ;
    oai21 ix613 (.Y (nx612), .A0 (nx11081), .A1 (nx11441), .B0 (nx11415)) ;
    inv01 ix11080 (.Y (nx11081), .A (d_arr_mul_22__19)) ;
    oai21 ix619 (.Y (nx618), .A0 (nx11083), .A1 (nx11441), .B0 (nx11415)) ;
    inv01 ix11082 (.Y (nx11083), .A (d_arr_mul_22__20)) ;
    oai21 ix625 (.Y (nx624), .A0 (nx11085), .A1 (nx11441), .B0 (nx11415)) ;
    inv01 ix11084 (.Y (nx11085), .A (d_arr_mul_22__21)) ;
    oai21 ix631 (.Y (nx630), .A0 (nx11087), .A1 (nx11441), .B0 (nx11417)) ;
    inv01 ix11086 (.Y (nx11087), .A (d_arr_mul_22__22)) ;
    oai21 ix637 (.Y (nx636), .A0 (nx11089), .A1 (nx11441), .B0 (nx11417)) ;
    inv01 ix11088 (.Y (nx11089), .A (d_arr_mul_22__23)) ;
    oai21 ix643 (.Y (nx642), .A0 (nx11091), .A1 (nx11443), .B0 (nx11417)) ;
    inv01 ix11090 (.Y (nx11091), .A (d_arr_mul_22__24)) ;
    oai21 ix649 (.Y (nx648), .A0 (nx11093), .A1 (nx11443), .B0 (nx11417)) ;
    inv01 ix11092 (.Y (nx11093), .A (d_arr_mul_22__25)) ;
    oai21 ix655 (.Y (nx654), .A0 (nx11095), .A1 (nx11443), .B0 (nx11417)) ;
    inv01 ix11094 (.Y (nx11095), .A (d_arr_mul_22__26)) ;
    oai21 ix661 (.Y (nx660), .A0 (nx11097), .A1 (nx11443), .B0 (nx11417)) ;
    inv01 ix11096 (.Y (nx11097), .A (d_arr_mul_22__27)) ;
    oai21 ix667 (.Y (nx666), .A0 (nx11099), .A1 (nx11443), .B0 (nx11417)) ;
    inv01 ix11098 (.Y (nx11099), .A (d_arr_mul_22__28)) ;
    oai21 ix673 (.Y (nx672), .A0 (nx11101), .A1 (nx11443), .B0 (nx10611)) ;
    inv01 ix11100 (.Y (nx11101), .A (d_arr_mul_22__29)) ;
    oai21 ix679 (.Y (nx678), .A0 (nx11103), .A1 (nx11443), .B0 (nx10611)) ;
    inv01 ix11102 (.Y (nx11103), .A (d_arr_mul_22__30)) ;
    oai21 ix685 (.Y (nx684), .A0 (nx11105), .A1 (nx10917), .B0 (nx10611)) ;
    inv01 ix11104 (.Y (nx11105), .A (d_arr_mul_22__31)) ;
    oai21 ix5169 (.Y (nx5168), .A0 (nx11107), .A1 (nx11445), .B0 (nx11419)) ;
    inv01 ix11106 (.Y (nx11107), .A (d_arr_mul_8__15)) ;
    nand02 ix5165 (.Y (nx10749), .A0 (nx11503), .A1 (d_arr_mux_8__31)) ;
    oai21 ix5175 (.Y (nx5174), .A0 (nx11109), .A1 (nx11447), .B0 (nx11419)) ;
    inv01 ix11108 (.Y (nx11109), .A (d_arr_mul_8__16)) ;
    oai21 ix5181 (.Y (nx5180), .A0 (nx11111), .A1 (nx11447), .B0 (nx11419)) ;
    inv01 ix11110 (.Y (nx11111), .A (d_arr_mul_8__17)) ;
    oai21 ix5187 (.Y (nx5186), .A0 (nx11113), .A1 (nx11447), .B0 (nx11419)) ;
    inv01 ix11112 (.Y (nx11113), .A (d_arr_mul_8__18)) ;
    oai21 ix5193 (.Y (nx5192), .A0 (nx11115), .A1 (nx11447), .B0 (nx11419)) ;
    inv01 ix11114 (.Y (nx11115), .A (d_arr_mul_8__19)) ;
    oai21 ix5199 (.Y (nx5198), .A0 (nx11117), .A1 (nx11447), .B0 (nx11419)) ;
    inv01 ix11116 (.Y (nx11117), .A (d_arr_mul_8__20)) ;
    oai21 ix5205 (.Y (nx5204), .A0 (nx11119), .A1 (nx11447), .B0 (nx11419)) ;
    inv01 ix11118 (.Y (nx11119), .A (d_arr_mul_8__21)) ;
    oai21 ix5211 (.Y (nx5210), .A0 (nx11121), .A1 (nx11447), .B0 (nx11421)) ;
    inv01 ix11120 (.Y (nx11121), .A (d_arr_mul_8__22)) ;
    oai21 ix5217 (.Y (nx5216), .A0 (nx11123), .A1 (nx10935), .B0 (nx11421)) ;
    inv01 ix11122 (.Y (nx11123), .A (d_arr_mul_8__23)) ;
    oai21 ix5223 (.Y (nx5222), .A0 (nx11125), .A1 (nx10935), .B0 (nx11421)) ;
    inv01 ix11124 (.Y (nx11125), .A (d_arr_mul_8__24)) ;
    oai21 ix5229 (.Y (nx5228), .A0 (nx11127), .A1 (nx10935), .B0 (nx11421)) ;
    inv01 ix11126 (.Y (nx11127), .A (d_arr_mul_8__25)) ;
    oai21 ix5235 (.Y (nx5234), .A0 (nx11129), .A1 (nx10935), .B0 (nx11421)) ;
    inv01 ix11128 (.Y (nx11129), .A (d_arr_mul_8__26)) ;
    oai21 ix5241 (.Y (nx5240), .A0 (nx11131), .A1 (nx11449), .B0 (nx11421)) ;
    inv01 ix11130 (.Y (nx11131), .A (d_arr_mul_8__27)) ;
    oai21 ix5247 (.Y (nx5246), .A0 (nx11133), .A1 (nx11449), .B0 (nx11421)) ;
    inv01 ix11132 (.Y (nx11133), .A (d_arr_mul_8__28)) ;
    oai21 ix5253 (.Y (nx5252), .A0 (nx11135), .A1 (nx11451), .B0 (nx10749)) ;
    inv01 ix11134 (.Y (nx11135), .A (d_arr_mul_8__29)) ;
    oai21 ix5259 (.Y (nx5258), .A0 (nx11137), .A1 (nx11451), .B0 (nx10749)) ;
    inv01 ix11136 (.Y (nx11137), .A (d_arr_mul_8__30)) ;
    oai21 ix5265 (.Y (nx5264), .A0 (nx11139), .A1 (nx11451), .B0 (nx10749)) ;
    inv01 ix11138 (.Y (nx11139), .A (d_arr_mul_8__31)) ;
    oai21 ix5393 (.Y (nx5392), .A0 (nx11141), .A1 (nx11451), .B0 (nx11423)) ;
    inv01 ix11140 (.Y (nx11141), .A (d_arr_mul_7__15)) ;
    nand02 ix5389 (.Y (nx10757), .A0 (nx11503), .A1 (d_arr_mux_7__31)) ;
    oai21 ix5399 (.Y (nx5398), .A0 (nx11143), .A1 (nx11451), .B0 (nx11423)) ;
    inv01 ix11142 (.Y (nx11143), .A (d_arr_mul_7__16)) ;
    oai21 ix5405 (.Y (nx5404), .A0 (nx11145), .A1 (nx11451), .B0 (nx11423)) ;
    inv01 ix11144 (.Y (nx11145), .A (d_arr_mul_7__17)) ;
    oai21 ix5411 (.Y (nx5410), .A0 (nx11147), .A1 (nx11451), .B0 (nx11423)) ;
    inv01 ix11146 (.Y (nx11147), .A (d_arr_mul_7__18)) ;
    oai21 ix5417 (.Y (nx5416), .A0 (nx11149), .A1 (nx11453), .B0 (nx11423)) ;
    inv01 ix11148 (.Y (nx11149), .A (d_arr_mul_7__19)) ;
    oai21 ix5423 (.Y (nx5422), .A0 (nx11151), .A1 (nx11453), .B0 (nx11423)) ;
    inv01 ix11150 (.Y (nx11151), .A (d_arr_mul_7__20)) ;
    oai21 ix5429 (.Y (nx5428), .A0 (nx11153), .A1 (nx11453), .B0 (nx11423)) ;
    inv01 ix11152 (.Y (nx11153), .A (d_arr_mul_7__21)) ;
    oai21 ix5435 (.Y (nx5434), .A0 (nx11155), .A1 (nx11453), .B0 (nx11425)) ;
    inv01 ix11154 (.Y (nx11155), .A (d_arr_mul_7__22)) ;
    oai21 ix5441 (.Y (nx5440), .A0 (nx11157), .A1 (nx11453), .B0 (nx11425)) ;
    inv01 ix11156 (.Y (nx11157), .A (d_arr_mul_7__23)) ;
    oai21 ix5447 (.Y (nx5446), .A0 (nx11159), .A1 (nx11453), .B0 (nx11425)) ;
    inv01 ix11158 (.Y (nx11159), .A (d_arr_mul_7__24)) ;
    oai21 ix5453 (.Y (nx5452), .A0 (nx11161), .A1 (nx11453), .B0 (nx11425)) ;
    inv01 ix11160 (.Y (nx11161), .A (d_arr_mul_7__25)) ;
    oai21 ix5459 (.Y (nx5458), .A0 (nx11163), .A1 (nx10937), .B0 (nx11425)) ;
    inv01 ix11162 (.Y (nx11163), .A (d_arr_mul_7__26)) ;
    oai21 ix5465 (.Y (nx5464), .A0 (nx11165), .A1 (nx10937), .B0 (nx11425)) ;
    inv01 ix11164 (.Y (nx11165), .A (d_arr_mul_7__27)) ;
    oai21 ix5471 (.Y (nx5470), .A0 (nx11167), .A1 (nx10937), .B0 (nx11425)) ;
    inv01 ix11166 (.Y (nx11167), .A (d_arr_mul_7__28)) ;
    oai21 ix5477 (.Y (nx5476), .A0 (nx11169), .A1 (nx10937), .B0 (nx10757)) ;
    inv01 ix11168 (.Y (nx11169), .A (d_arr_mul_7__29)) ;
    oai21 ix5483 (.Y (nx5482), .A0 (nx11171), .A1 (nx10937), .B0 (nx10757)) ;
    inv01 ix11170 (.Y (nx11171), .A (d_arr_mul_7__30)) ;
    oai21 ix5489 (.Y (nx5488), .A0 (nx11173), .A1 (nx10937), .B0 (nx10757)) ;
    inv01 ix11172 (.Y (nx11173), .A (d_arr_mul_7__31)) ;
    oai21 ix5617 (.Y (nx5616), .A0 (nx11175), .A1 (nx11455), .B0 (nx11427)) ;
    inv01 ix11174 (.Y (nx11175), .A (d_arr_mul_6__15)) ;
    nand02 ix5613 (.Y (nx10765), .A0 (nx11503), .A1 (d_arr_mux_6__31)) ;
    oai21 ix5623 (.Y (nx5622), .A0 (nx11177), .A1 (nx11455), .B0 (nx11427)) ;
    inv01 ix11176 (.Y (nx11177), .A (d_arr_mul_6__16)) ;
    oai21 ix5629 (.Y (nx5628), .A0 (nx11179), .A1 (nx11455), .B0 (nx11427)) ;
    inv01 ix11178 (.Y (nx11179), .A (d_arr_mul_6__17)) ;
    oai21 ix5635 (.Y (nx5634), .A0 (nx11181), .A1 (nx11457), .B0 (nx11427)) ;
    inv01 ix11180 (.Y (nx11181), .A (d_arr_mul_6__18)) ;
    oai21 ix5641 (.Y (nx5640), .A0 (nx11183), .A1 (nx11457), .B0 (nx11427)) ;
    inv01 ix11182 (.Y (nx11183), .A (d_arr_mul_6__19)) ;
    oai21 ix5647 (.Y (nx5646), .A0 (nx11185), .A1 (nx11457), .B0 (nx11427)) ;
    inv01 ix11184 (.Y (nx11185), .A (d_arr_mul_6__20)) ;
    oai21 ix5653 (.Y (nx5652), .A0 (nx11187), .A1 (nx11457), .B0 (nx11427)) ;
    inv01 ix11186 (.Y (nx11187), .A (d_arr_mul_6__21)) ;
    oai21 ix5659 (.Y (nx5658), .A0 (nx11189), .A1 (nx11457), .B0 (nx11429)) ;
    inv01 ix11188 (.Y (nx11189), .A (d_arr_mul_6__22)) ;
    oai21 ix5665 (.Y (nx5664), .A0 (nx11191), .A1 (nx11457), .B0 (nx11429)) ;
    inv01 ix11190 (.Y (nx11191), .A (d_arr_mul_6__23)) ;
    oai21 ix5671 (.Y (nx5670), .A0 (nx11193), .A1 (nx11457), .B0 (nx11429)) ;
    inv01 ix11192 (.Y (nx11193), .A (d_arr_mul_6__24)) ;
    oai21 ix5677 (.Y (nx5676), .A0 (nx11195), .A1 (nx11459), .B0 (nx11429)) ;
    inv01 ix11194 (.Y (nx11195), .A (d_arr_mul_6__25)) ;
    oai21 ix5683 (.Y (nx5682), .A0 (nx11197), .A1 (nx11459), .B0 (nx11429)) ;
    inv01 ix11196 (.Y (nx11197), .A (d_arr_mul_6__26)) ;
    oai21 ix5689 (.Y (nx5688), .A0 (nx11199), .A1 (nx11459), .B0 (nx11429)) ;
    inv01 ix11198 (.Y (nx11199), .A (d_arr_mul_6__27)) ;
    oai21 ix5695 (.Y (nx5694), .A0 (nx11201), .A1 (nx11459), .B0 (nx11429)) ;
    inv01 ix11200 (.Y (nx11201), .A (d_arr_mul_6__28)) ;
    oai21 ix5701 (.Y (nx5700), .A0 (nx11203), .A1 (nx11459), .B0 (nx10765)) ;
    inv01 ix11202 (.Y (nx11203), .A (d_arr_mul_6__29)) ;
    oai21 ix5707 (.Y (nx5706), .A0 (nx11205), .A1 (nx11459), .B0 (nx10765)) ;
    inv01 ix11204 (.Y (nx11205), .A (d_arr_mul_6__30)) ;
    oai21 ix5713 (.Y (nx5712), .A0 (nx11207), .A1 (nx11459), .B0 (nx10765)) ;
    inv01 ix11206 (.Y (nx11207), .A (d_arr_mul_6__31)) ;
    oai21 ix5841 (.Y (nx5840), .A0 (nx11209), .A1 (nx11461), .B0 (nx11431)) ;
    inv01 ix11208 (.Y (nx11209), .A (d_arr_mul_5__15)) ;
    nand02 ix5837 (.Y (nx10773), .A0 (nx11503), .A1 (d_arr_mux_5__31)) ;
    oai21 ix5847 (.Y (nx5846), .A0 (nx11211), .A1 (nx11461), .B0 (nx11431)) ;
    inv01 ix11210 (.Y (nx11211), .A (d_arr_mul_5__16)) ;
    oai21 ix5853 (.Y (nx5852), .A0 (nx11213), .A1 (nx11461), .B0 (nx11431)) ;
    inv01 ix11212 (.Y (nx11213), .A (d_arr_mul_5__17)) ;
    oai21 ix5859 (.Y (nx5858), .A0 (nx11215), .A1 (nx11461), .B0 (nx11431)) ;
    inv01 ix11214 (.Y (nx11215), .A (d_arr_mul_5__18)) ;
    oai21 ix5865 (.Y (nx5864), .A0 (nx11217), .A1 (nx11461), .B0 (nx11431)) ;
    inv01 ix11216 (.Y (nx11217), .A (d_arr_mul_5__19)) ;
    oai21 ix5871 (.Y (nx5870), .A0 (nx11219), .A1 (nx11461), .B0 (nx11431)) ;
    inv01 ix11218 (.Y (nx11219), .A (d_arr_mul_5__20)) ;
    oai21 ix5877 (.Y (nx5876), .A0 (nx11221), .A1 (nx11461), .B0 (nx11431)) ;
    inv01 ix11220 (.Y (nx11221), .A (d_arr_mul_5__21)) ;
    oai21 ix5883 (.Y (nx5882), .A0 (nx11223), .A1 (nx10939), .B0 (nx11433)) ;
    inv01 ix11222 (.Y (nx11223), .A (d_arr_mul_5__22)) ;
    oai21 ix5889 (.Y (nx5888), .A0 (nx11225), .A1 (nx10939), .B0 (nx11433)) ;
    inv01 ix11224 (.Y (nx11225), .A (d_arr_mul_5__23)) ;
    oai21 ix5895 (.Y (nx5894), .A0 (nx11227), .A1 (nx10939), .B0 (nx11433)) ;
    inv01 ix11226 (.Y (nx11227), .A (d_arr_mul_5__24)) ;
    oai21 ix5901 (.Y (nx5900), .A0 (nx11229), .A1 (nx10939), .B0 (nx11433)) ;
    inv01 ix11228 (.Y (nx11229), .A (d_arr_mul_5__25)) ;
    oai21 ix5907 (.Y (nx5906), .A0 (nx11231), .A1 (nx10939), .B0 (nx11433)) ;
    inv01 ix11230 (.Y (nx11231), .A (d_arr_mul_5__26)) ;
    oai21 ix5913 (.Y (nx5912), .A0 (nx11233), .A1 (nx10939), .B0 (nx11433)) ;
    inv01 ix11232 (.Y (nx11233), .A (d_arr_mul_5__27)) ;
    oai21 ix5919 (.Y (nx5918), .A0 (nx11235), .A1 (nx10939), .B0 (nx11433)) ;
    inv01 ix11234 (.Y (nx11235), .A (d_arr_mul_5__28)) ;
    oai21 ix5925 (.Y (nx5924), .A0 (nx11237), .A1 (nx10941), .B0 (nx10773)) ;
    inv01 ix11236 (.Y (nx11237), .A (d_arr_mul_5__29)) ;
    oai21 ix5931 (.Y (nx5930), .A0 (nx11239), .A1 (nx10941), .B0 (nx10773)) ;
    inv01 ix11238 (.Y (nx11239), .A (d_arr_mul_5__30)) ;
    oai21 ix5937 (.Y (nx5936), .A0 (nx11241), .A1 (nx10941), .B0 (nx10773)) ;
    inv01 ix11240 (.Y (nx11241), .A (d_arr_mul_5__31)) ;
    inv02 ix11244 (.Y (nx11245), .A (nx11524)) ;
    inv02 ix11246 (.Y (nx11247), .A (nx11524)) ;
    inv02 ix11248 (.Y (nx11249), .A (nx11524)) ;
    inv02 ix11250 (.Y (nx11251), .A (nx11524)) ;
    inv02 ix11252 (.Y (nx11253), .A (nx11525)) ;
    inv02 ix11254 (.Y (nx11255), .A (nx11525)) ;
    inv02 ix11256 (.Y (nx11257), .A (nx11525)) ;
    inv02 ix11258 (.Y (nx11259), .A (nx11479)) ;
    inv02 ix11260 (.Y (nx11261), .A (nx11479)) ;
    inv02 ix11262 (.Y (nx11263), .A (nx11479)) ;
    inv02 ix11264 (.Y (nx11265), .A (nx11479)) ;
    inv02 ix11266 (.Y (nx11267), .A (nx11479)) ;
    inv02 ix11268 (.Y (nx11269), .A (nx11479)) ;
    inv02 ix11270 (.Y (nx11271), .A (nx11479)) ;
    inv02 ix11272 (.Y (nx11273), .A (nx11481)) ;
    inv02 ix11274 (.Y (nx11275), .A (nx11481)) ;
    inv02 ix11276 (.Y (nx11277), .A (nx11481)) ;
    inv02 ix11278 (.Y (nx11279), .A (nx11481)) ;
    inv02 ix11280 (.Y (nx11281), .A (nx11481)) ;
    inv02 ix11282 (.Y (nx11283), .A (nx11481)) ;
    inv02 ix11284 (.Y (nx11285), .A (nx11481)) ;
    inv02 ix11286 (.Y (nx11287), .A (nx11483)) ;
    inv02 ix11288 (.Y (nx11289), .A (nx11483)) ;
    inv02 ix11290 (.Y (nx11291), .A (nx11483)) ;
    inv02 ix11292 (.Y (nx11293), .A (nx11483)) ;
    inv02 ix11294 (.Y (nx11295), .A (nx11483)) ;
    inv02 ix11296 (.Y (nx11297), .A (nx11483)) ;
    inv02 ix11298 (.Y (nx11299), .A (nx11483)) ;
    inv02 ix11300 (.Y (nx11301), .A (nx11485)) ;
    inv02 ix11302 (.Y (nx11303), .A (nx11485)) ;
    inv02 ix11304 (.Y (nx11305), .A (nx11485)) ;
    inv02 ix11306 (.Y (nx11307), .A (nx11485)) ;
    inv02 ix11308 (.Y (nx11309), .A (nx11485)) ;
    inv02 ix11310 (.Y (nx11311), .A (nx11485)) ;
    inv02 ix11312 (.Y (nx11313), .A (nx11485)) ;
    inv02 ix11314 (.Y (nx11315), .A (nx11487)) ;
    inv02 ix11316 (.Y (nx11317), .A (nx11487)) ;
    inv02 ix11318 (.Y (nx11319), .A (nx11487)) ;
    inv02 ix11320 (.Y (nx11321), .A (nx11487)) ;
    inv02 ix11322 (.Y (nx11323), .A (nx11487)) ;
    inv02 ix11324 (.Y (nx11325), .A (nx11487)) ;
    inv02 ix11326 (.Y (nx11327), .A (nx11487)) ;
    inv02 ix11328 (.Y (nx11329), .A (nx11489)) ;
    inv02 ix11330 (.Y (nx11331), .A (nx11489)) ;
    inv02 ix11332 (.Y (nx11333), .A (nx11489)) ;
    inv02 ix11334 (.Y (nx11335), .A (nx11489)) ;
    inv02 ix11336 (.Y (nx11337), .A (nx11489)) ;
    inv02 ix11338 (.Y (nx11339), .A (nx11489)) ;
    inv02 ix11340 (.Y (nx11341), .A (nx11489)) ;
    inv02 ix11342 (.Y (nx11343), .A (nx11491)) ;
    inv02 ix11344 (.Y (nx11345), .A (nx11491)) ;
    inv02 ix11346 (.Y (nx11347), .A (nx11491)) ;
    inv02 ix11348 (.Y (nx11349), .A (nx11491)) ;
    inv02 ix11350 (.Y (nx11351), .A (nx11491)) ;
    inv02 ix11352 (.Y (nx11353), .A (nx11491)) ;
    inv02 ix11354 (.Y (nx11355), .A (nx11491)) ;
    inv02 ix11356 (.Y (nx11357), .A (nx11493)) ;
    inv02 ix11358 (.Y (nx11359), .A (nx11493)) ;
    inv02 ix11360 (.Y (nx11361), .A (nx11493)) ;
    inv02 ix11362 (.Y (nx11363), .A (nx11493)) ;
    inv02 ix11364 (.Y (nx11365), .A (nx11493)) ;
    inv02 ix11366 (.Y (nx11367), .A (nx11493)) ;
    inv02 ix11368 (.Y (nx11369), .A (nx11493)) ;
    inv02 ix11370 (.Y (nx11371), .A (nx11495)) ;
    inv02 ix11372 (.Y (nx11373), .A (nx11495)) ;
    inv02 ix11374 (.Y (nx11375), .A (nx11495)) ;
    inv02 ix11376 (.Y (nx11377), .A (nx11495)) ;
    inv02 ix11378 (.Y (nx11379), .A (nx11495)) ;
    inv02 ix11380 (.Y (nx11381), .A (nx11495)) ;
    inv02 ix11382 (.Y (nx11383), .A (nx11495)) ;
    inv02 ix11384 (.Y (nx11385), .A (nx11497)) ;
    inv02 ix11386 (.Y (nx11387), .A (nx11497)) ;
    inv02 ix11388 (.Y (nx11389), .A (nx11497)) ;
    inv02 ix11390 (.Y (nx11391), .A (nx11497)) ;
    inv02 ix11392 (.Y (nx11393), .A (nx11497)) ;
    inv02 ix11394 (.Y (nx11395), .A (nx11497)) ;
    inv02 ix11396 (.Y (nx11397), .A (nx11497)) ;
    inv02 ix11398 (.Y (nx11399), .A (nx11499)) ;
    inv02 ix11400 (.Y (nx11401), .A (nx11499)) ;
    inv02 ix11402 (.Y (nx11403), .A (nx11499)) ;
    inv02 ix11404 (.Y (nx11405), .A (nx11499)) ;
    nand02 ix11406 (.Y (nx11407), .A0 (nx11403), .A1 (d_arr_mux_24__31)) ;
    nand02 ix11408 (.Y (nx11409), .A0 (nx11403), .A1 (d_arr_mux_24__31)) ;
    nand02 ix11410 (.Y (nx11411), .A0 (nx11503), .A1 (d_arr_mux_23__31)) ;
    nand02 ix11412 (.Y (nx11413), .A0 (nx11505), .A1 (d_arr_mux_23__31)) ;
    nand02 ix11414 (.Y (nx11415), .A0 (nx11505), .A1 (d_arr_mux_22__31)) ;
    nand02 ix11416 (.Y (nx11417), .A0 (nx11505), .A1 (d_arr_mux_22__31)) ;
    nand02 ix11418 (.Y (nx11419), .A0 (nx11505), .A1 (d_arr_mux_8__31)) ;
    nand02 ix11420 (.Y (nx11421), .A0 (nx11505), .A1 (d_arr_mux_8__31)) ;
    nand02 ix11422 (.Y (nx11423), .A0 (nx11505), .A1 (d_arr_mux_7__31)) ;
    nand02 ix11424 (.Y (nx11425), .A0 (nx11505), .A1 (d_arr_mux_7__31)) ;
    nand02 ix11426 (.Y (nx11427), .A0 (nx11405), .A1 (d_arr_mux_6__31)) ;
    nand02 ix11428 (.Y (nx11429), .A0 (nx11405), .A1 (d_arr_mux_6__31)) ;
    nand02 ix11430 (.Y (nx11431), .A0 (nx11405), .A1 (d_arr_mux_5__31)) ;
    nand02 ix11432 (.Y (nx11433), .A0 (nx11405), .A1 (d_arr_mux_5__31)) ;
    inv02 ix11434 (.Y (nx11435), .A (nx10985)) ;
    inv02 ix11436 (.Y (nx11437), .A (nx10985)) ;
    inv02 ix11438 (.Y (nx11439), .A (nx10985)) ;
    inv02 ix11440 (.Y (nx11441), .A (nx10985)) ;
    inv02 ix11442 (.Y (nx11443), .A (nx10985)) ;
    inv02 ix11444 (.Y (nx11445), .A (nx11469)) ;
    inv02 ix11446 (.Y (nx11447), .A (nx11469)) ;
    inv02 ix11448 (.Y (nx11449), .A (nx11469)) ;
    inv02 ix11450 (.Y (nx11451), .A (nx11469)) ;
    inv02 ix11452 (.Y (nx11453), .A (nx11469)) ;
    inv02 ix11454 (.Y (nx11455), .A (nx11469)) ;
    inv02 ix11456 (.Y (nx11457), .A (nx11469)) ;
    inv02 ix11458 (.Y (nx11459), .A (nx10987)) ;
    inv02 ix11460 (.Y (nx11461), .A (nx10987)) ;
    inv02 ix11462 (.Y (nx11463), .A (nx10987)) ;
    inv02 ix11464 (.Y (nx11465), .A (nx10915)) ;
    inv02 ix11466 (.Y (nx11467), .A (nx10915)) ;
    inv02 ix11468 (.Y (nx11469), .A (nx10915)) ;
    inv02 ix11470 (.Y (nx11471), .A (nx11511)) ;
    inv02 ix11472 (.Y (nx11473), .A (nx11511)) ;
    inv02 ix11474 (.Y (nx11475), .A (nx11511)) ;
    inv02 ix11476 (.Y (nx11477), .A (sel_mux)) ;
    inv02 ix11478 (.Y (nx11479), .A (nx11517)) ;
    inv02 ix11480 (.Y (nx11481), .A (nx11517)) ;
    inv02 ix11482 (.Y (nx11483), .A (nx11517)) ;
    inv02 ix11484 (.Y (nx11485), .A (nx11517)) ;
    inv02 ix11486 (.Y (nx11487), .A (nx11517)) ;
    inv02 ix11488 (.Y (nx11489), .A (nx11517)) ;
    inv02 ix11490 (.Y (nx11491), .A (nx11517)) ;
    inv02 ix11492 (.Y (nx11493), .A (nx11519)) ;
    inv02 ix11494 (.Y (nx11495), .A (nx11519)) ;
    inv02 ix11496 (.Y (nx11497), .A (nx11519)) ;
    inv02 ix11498 (.Y (nx11499), .A (nx11519)) ;
    inv02 ix11500 (.Y (nx11501), .A (nx11499)) ;
    inv02 ix11502 (.Y (nx11503), .A (nx11499)) ;
    inv02 ix11504 (.Y (nx11505), .A (nx11499)) ;
    inv01 ix11510 (.Y (nx11511), .A (nx10915)) ;
    inv02 ix11516 (.Y (nx11517), .A (nx11525)) ;
    inv02 ix11518 (.Y (nx11519), .A (nx11525)) ;
    buf16 ix11526 (.Y (nx11524), .A (nx11477)) ;
    buf16 ix11527 (.Y (nx11525), .A (nx11477)) ;
endmodule


module Controller_16_16_5_16 ( clk, reset, io_ready_in, io_done_out, mem_data_in, 
                               mem_data_out, mem_addr_out, mem_write_out, 
                               mem_read_out, wind_en, wind_rst, 
                               wind_col_in_4__15, wind_col_in_4__14, 
                               wind_col_in_4__13, wind_col_in_4__12, 
                               wind_col_in_4__11, wind_col_in_4__10, 
                               wind_col_in_4__9, wind_col_in_4__8, 
                               wind_col_in_4__7, wind_col_in_4__6, 
                               wind_col_in_4__5, wind_col_in_4__4, 
                               wind_col_in_4__3, wind_col_in_4__2, 
                               wind_col_in_4__1, wind_col_in_4__0, 
                               wind_col_in_3__15, wind_col_in_3__14, 
                               wind_col_in_3__13, wind_col_in_3__12, 
                               wind_col_in_3__11, wind_col_in_3__10, 
                               wind_col_in_3__9, wind_col_in_3__8, 
                               wind_col_in_3__7, wind_col_in_3__6, 
                               wind_col_in_3__5, wind_col_in_3__4, 
                               wind_col_in_3__3, wind_col_in_3__2, 
                               wind_col_in_3__1, wind_col_in_3__0, 
                               wind_col_in_2__15, wind_col_in_2__14, 
                               wind_col_in_2__13, wind_col_in_2__12, 
                               wind_col_in_2__11, wind_col_in_2__10, 
                               wind_col_in_2__9, wind_col_in_2__8, 
                               wind_col_in_2__7, wind_col_in_2__6, 
                               wind_col_in_2__5, wind_col_in_2__4, 
                               wind_col_in_2__3, wind_col_in_2__2, 
                               wind_col_in_2__1, wind_col_in_2__0, 
                               wind_col_in_1__15, wind_col_in_1__14, 
                               wind_col_in_1__13, wind_col_in_1__12, 
                               wind_col_in_1__11, wind_col_in_1__10, 
                               wind_col_in_1__9, wind_col_in_1__8, 
                               wind_col_in_1__7, wind_col_in_1__6, 
                               wind_col_in_1__5, wind_col_in_1__4, 
                               wind_col_in_1__3, wind_col_in_1__2, 
                               wind_col_in_1__1, wind_col_in_1__0, 
                               wind_col_in_0__15, wind_col_in_0__14, 
                               wind_col_in_0__13, wind_col_in_0__12, 
                               wind_col_in_0__11, wind_col_in_0__10, 
                               wind_col_in_0__9, wind_col_in_0__8, 
                               wind_col_in_0__7, wind_col_in_0__6, 
                               wind_col_in_0__5, wind_col_in_0__4, 
                               wind_col_in_0__3, wind_col_in_0__2, 
                               wind_col_in_0__1, wind_col_in_0__0, 
                               filter_data_out, filter_ready_out, filter_reset, 
                               comp_unit_ready, comp_unit_operation, 
                               comp_unit_flt_size, comp_unit_relu, 
                               comp_unit_data1_out, comp_unit_data2_out, 
                               comp_unit_buffer_finished, comp_unit_finished, 
                               comp_unit_data1_in, comp_unit_data2_in, 
                               argmax_ready, argmax_data_out, argmax_data_in ) ;

    input clk ;
    input reset ;
    input io_ready_in ;
    output io_done_out ;
    input [15:0]mem_data_in ;
    output [15:0]mem_data_out ;
    output [15:0]mem_addr_out ;
    output mem_write_out ;
    output mem_read_out ;
    output wind_en ;
    output wind_rst ;
    output wind_col_in_4__15 ;
    output wind_col_in_4__14 ;
    output wind_col_in_4__13 ;
    output wind_col_in_4__12 ;
    output wind_col_in_4__11 ;
    output wind_col_in_4__10 ;
    output wind_col_in_4__9 ;
    output wind_col_in_4__8 ;
    output wind_col_in_4__7 ;
    output wind_col_in_4__6 ;
    output wind_col_in_4__5 ;
    output wind_col_in_4__4 ;
    output wind_col_in_4__3 ;
    output wind_col_in_4__2 ;
    output wind_col_in_4__1 ;
    output wind_col_in_4__0 ;
    output wind_col_in_3__15 ;
    output wind_col_in_3__14 ;
    output wind_col_in_3__13 ;
    output wind_col_in_3__12 ;
    output wind_col_in_3__11 ;
    output wind_col_in_3__10 ;
    output wind_col_in_3__9 ;
    output wind_col_in_3__8 ;
    output wind_col_in_3__7 ;
    output wind_col_in_3__6 ;
    output wind_col_in_3__5 ;
    output wind_col_in_3__4 ;
    output wind_col_in_3__3 ;
    output wind_col_in_3__2 ;
    output wind_col_in_3__1 ;
    output wind_col_in_3__0 ;
    output wind_col_in_2__15 ;
    output wind_col_in_2__14 ;
    output wind_col_in_2__13 ;
    output wind_col_in_2__12 ;
    output wind_col_in_2__11 ;
    output wind_col_in_2__10 ;
    output wind_col_in_2__9 ;
    output wind_col_in_2__8 ;
    output wind_col_in_2__7 ;
    output wind_col_in_2__6 ;
    output wind_col_in_2__5 ;
    output wind_col_in_2__4 ;
    output wind_col_in_2__3 ;
    output wind_col_in_2__2 ;
    output wind_col_in_2__1 ;
    output wind_col_in_2__0 ;
    output wind_col_in_1__15 ;
    output wind_col_in_1__14 ;
    output wind_col_in_1__13 ;
    output wind_col_in_1__12 ;
    output wind_col_in_1__11 ;
    output wind_col_in_1__10 ;
    output wind_col_in_1__9 ;
    output wind_col_in_1__8 ;
    output wind_col_in_1__7 ;
    output wind_col_in_1__6 ;
    output wind_col_in_1__5 ;
    output wind_col_in_1__4 ;
    output wind_col_in_1__3 ;
    output wind_col_in_1__2 ;
    output wind_col_in_1__1 ;
    output wind_col_in_1__0 ;
    output wind_col_in_0__15 ;
    output wind_col_in_0__14 ;
    output wind_col_in_0__13 ;
    output wind_col_in_0__12 ;
    output wind_col_in_0__11 ;
    output wind_col_in_0__10 ;
    output wind_col_in_0__9 ;
    output wind_col_in_0__8 ;
    output wind_col_in_0__7 ;
    output wind_col_in_0__6 ;
    output wind_col_in_0__5 ;
    output wind_col_in_0__4 ;
    output wind_col_in_0__3 ;
    output wind_col_in_0__2 ;
    output wind_col_in_0__1 ;
    output wind_col_in_0__0 ;
    output [15:0]filter_data_out ;
    output filter_ready_out ;
    output filter_reset ;
    output comp_unit_ready ;
    output comp_unit_operation ;
    output comp_unit_flt_size ;
    output comp_unit_relu ;
    output [15:0]comp_unit_data1_out ;
    output [15:0]comp_unit_data2_out ;
    input comp_unit_buffer_finished ;
    input comp_unit_finished ;
    input [15:0]comp_unit_data1_in ;
    input [15:0]comp_unit_data2_in ;
    output argmax_ready ;
    output [15:0]argmax_data_out ;
    input [15:0]argmax_data_in ;

    wire current_state_13, wind_width_count_4, wind_width_count_3, 
         wind_width_count_2, wind_width_count_1, wind_width_count_0, 
         cache_height_count_en, cache_height_ended, max_height_2, max_height_0, 
         cache_width_count_4, cache_width_count_3, cache_width_count_2, 
         cache_width_count_1, cache_width_count_0, cache_data_in_15, 
         cache_data_in_14, cache_data_in_13, cache_data_in_12, cache_data_in_11, 
         cache_data_in_10, cache_data_in_9, cache_data_in_8, cache_data_in_7, 
         cache_data_in_6, cache_data_in_5, cache_data_in_4, cache_data_in_3, 
         cache_data_in_2, cache_data_in_1, cache_data_in_0, cache_data_out_4__15, 
         cache_data_out_4__14, cache_data_out_4__13, cache_data_out_4__12, 
         cache_data_out_4__11, cache_data_out_4__10, cache_data_out_4__9, 
         cache_data_out_4__8, cache_data_out_4__7, cache_data_out_4__6, 
         cache_data_out_4__5, cache_data_out_4__4, cache_data_out_4__3, 
         cache_data_out_4__2, cache_data_out_4__1, cache_data_out_4__0, 
         cache_data_out_3__15, cache_data_out_3__14, cache_data_out_3__13, 
         cache_data_out_3__12, cache_data_out_3__11, cache_data_out_3__10, 
         cache_data_out_3__9, cache_data_out_3__8, cache_data_out_3__7, 
         cache_data_out_3__6, cache_data_out_3__5, cache_data_out_3__4, 
         cache_data_out_3__3, cache_data_out_3__2, cache_data_out_3__1, 
         cache_data_out_3__0, cache_data_out_2__15, cache_data_out_2__14, 
         cache_data_out_2__13, cache_data_out_2__12, cache_data_out_2__11, 
         cache_data_out_2__10, cache_data_out_2__9, cache_data_out_2__8, 
         cache_data_out_2__7, cache_data_out_2__6, cache_data_out_2__5, 
         cache_data_out_2__4, cache_data_out_2__3, cache_data_out_2__2, 
         cache_data_out_2__1, cache_data_out_2__0, cache_data_out_1__15, 
         cache_data_out_1__14, cache_data_out_1__13, cache_data_out_1__12, 
         cache_data_out_1__11, cache_data_out_1__10, cache_data_out_1__9, 
         cache_data_out_1__8, cache_data_out_1__7, cache_data_out_1__6, 
         cache_data_out_1__5, cache_data_out_1__4, cache_data_out_1__3, 
         cache_data_out_1__2, cache_data_out_1__1, cache_data_out_1__0, 
         cache_data_out_0__15, cache_data_out_0__14, cache_data_out_0__13, 
         cache_data_out_0__12, cache_data_out_0__11, cache_data_out_0__10, 
         cache_data_out_0__9, cache_data_out_0__8, cache_data_out_0__7, 
         cache_data_out_0__6, cache_data_out_0__5, cache_data_out_0__4, 
         cache_data_out_0__3, cache_data_out_0__2, cache_data_out_0__1, 
         cache_data_out_0__0, cache_load, cache_rst_actual, max_height_4, 
         max_height_3, max_height_1, current_state_21, current_state_20, 
         layer_type_out_1, current_state_3, nx1409, current_state_24, 
         ftc_cntrl_reg_out_12, current_state_16, ftc_cntrl_reg_out_8, nx1411, 
         nx4, nx14, ftc_cntrl_reg_out_14, current_state_12, current_state_25, 
         nflt_layer_out_3, current_state_4, nflt_layer_out_1, nflt_layer_out_0, 
         nx98, nx1419, nx112, current_state_9, current_state_8, current_state_7, 
         current_state_6, current_state_5, nx136, nx146, nx1421, nx152, 
         cntr1_inst_counter_out_1, cntr1_inst_counter_out_0, nx176, 
         cntr1_inst_counter_out_3, cntr1_inst_counter_out_2, nx200, nx214, 
         cntr1_inst_counter_out_4, nx1425, nx232, nx246, nx248, flt_size_out_0, 
         flt_size_out_2, flt_size_out_1, nx278, nx280, nx286, nx300, nx1427, 
         nx306, ftc_cntrl_reg_out_13, nx320, nx332, ftc_cntrl_reg_out_11, nx1429, 
         window_width_cntr_counter_out_14, nx1430, 
         window_width_cntr_counter_out_13, window_width_cntr_counter_out_12, 
         nx1432, window_width_cntr_counter_out_11, 
         window_width_cntr_counter_out_10, nx1434, 
         window_width_cntr_counter_out_9, window_width_cntr_counter_out_8, 
         nx1436, window_width_cntr_counter_out_7, 
         window_width_cntr_counter_out_6, nx1439, 
         window_width_cntr_counter_out_5, nx348, nx354, nx362, nx370, nx378, 
         nx398, nx422, nx446, nx470, nx494, nx520, nx534, nx546, img_width_out_0, 
         new_width_out_0, nx572, nx574, nx582, img_width_out_1, new_width_out_1, 
         nx600, nx606, nx610, img_width_out_2, new_width_out_2, nx644, 
         img_width_out_3, new_width_out_3, nx674, img_width_out_4, 
         new_width_out_4, nx692, nx702, current_state_15, 
         write_offset_data_out_0, nx730, new_size_squared_out_0, 
         write_offset_data_out_1, nx750, new_size_squared_out_1, 
         write_offset_data_out_2, new_size_squared_out_2, 
         write_offset_data_out_3, nx802, new_size_squared_out_3, nx820, 
         write_offset_data_out_4, nx822, nx828, new_size_squared_out_4, 
         write_offset_data_out_5, new_size_squared_out_5, 
         write_offset_data_out_6, nx868, nx874, new_size_squared_out_6, 
         write_offset_data_out_7, new_size_squared_out_7, nx914, 
         write_offset_data_out_8, nx918, nx924, new_size_squared_out_8, 
         write_offset_data_out_9, new_size_squared_out_9, 
         write_offset_data_out_10, nx964, nx970, new_size_squared_out_10, 
         write_offset_data_out_11, new_size_squared_out_11, nx1010, 
         write_offset_data_out_12, nx1012, nx1018, new_size_squared_out_12, 
         write_offset_data_out_13, new_size_squared_out_13, 
         write_offset_data_out_14, nx1058, nx1064, new_size_squared_out_14, 
         write_offset_data_out_15, new_size_squared_out_15, nx1098, nx1108, 
         ftc_cntrl_reg_out_9, nx1116, nx1124, nx1138, ftc_cntrl_reg_out_10, 
         nx1152, nx1166, cache_width_cntr_counter_out_14, nx1447, 
         cache_width_cntr_counter_out_13, cache_width_cntr_counter_out_12, 
         nx1449, cache_width_cntr_counter_out_11, 
         cache_width_cntr_counter_out_10, nx1451, cache_width_cntr_counter_out_9, 
         cache_width_cntr_counter_out_8, nx1454, cache_width_cntr_counter_out_7, 
         cache_width_cntr_counter_out_6, nx1456, nx1192, nx1198, nx1206, nx1214, 
         nx1222, cache_width_cntr_counter_out_5, nx1228, nx1248, nx1272, nx1296, 
         nx1320, nx1344, nx1370, nx1384, nx1402, nx1404, nx1406, nx1414, nx1416, 
         nx1424, nx1428, current_state_19, current_state_18, nx1446, nx1452, 
         nx1468, nx1459, nx1486, nx1492, nx1502, nx1461, nx1516, 
         num_channels_out_3, nflt_layer_temp_3, nx1528, nx1463, 
         num_channels_out_2, nflt_layer_temp_2, nx1464, num_channels_out_1, 
         nflt_layer_temp_1, num_channels_out_0, current_state_2, nx1572, nx1578, 
         nflt_layer_temp_0, max_num_channels_data_out_0, nx1594, nx1602, nx1610, 
         nx1620, nx1630, max_num_channels_data_out_1, nx1646, nx1652, nx1664, 
         max_num_channels_data_out_2, nx1678, nx1690, 
         max_num_channels_data_out_3, nx1704, nx1716, 
         max_num_channels_data_out_4, nlayers_counter_out_0, 
         nlayers_counter_out_2, nlayers_counter_out_1, nx1768, nx1784, nx1800, 
         nx1469, nx1842, nx1880, current_state_28, current_state_27, 
         class_cntr_counter_out_3, class_cntr_counter_out_2, 
         class_cntr_counter_out_1, class_cntr_counter_out_0, nx1908, nx1916, 
         nx1942, nx1950, flt_bias_out_0, nx2084, nx2096, nx2098, flt_bias_out_1, 
         nx2124, flt_bias_out_2, nx2150, flt_bias_out_3, nx2176, flt_bias_out_4, 
         nx2202, flt_bias_out_5, nx2228, flt_bias_out_6, nx2254, flt_bias_out_7, 
         nx2280, flt_bias_out_8, nx2306, flt_bias_out_9, nx2332, flt_bias_out_10, 
         nx2358, flt_bias_out_11, nx2384, flt_bias_out_12, nx2410, 
         flt_bias_out_13, nx2436, flt_bias_out_14, nx2462, flt_bias_out_15, 
         nx2488, nx2502, ftc_cntrl_reg_out_15, nx2522, nx2536, nx2580, nx2582, 
         bias_offset_data_out_0, nx2620, nx2626, img_base_addr_0, 
         write_base_prev_data_out_0, nx2636, nx2640, img_addr_offset_0, nx2680, 
         addr1_data_0, nx2706, write_base_data_out_1, nx2752, nx2760, nx2766, 
         addr1_data_1, bias_offset_data_out_1, nx2794, nx2796, img_base_addr_1, 
         write_base_prev_data_out_1, img_addr_offset_1, nx2832, nx2834, 
         write_base_data_out_2, nx2872, nx2882, nx2884, nx2886, nx2894, 
         addr1_data_2, nx2904, bias_offset_data_out_2, nx2932, img_base_addr_2, 
         write_base_prev_data_out_2, nx2950, nx2956, img_addr_offset_2, nx2970, 
         nx2978, write_base_data_out_3, nx3004, nx3006, nx3016, nx3032, nx3034, 
         addr1_data_3, nx3048, nx3066, bias_offset_data_out_3, nx3074, nx3076, 
         nx3086, img_base_addr_3, write_base_prev_data_out_3, nx3100, 
         img_addr_offset_3, nx3114, nx3120, nx3122, nx3138, 
         write_base_data_out_4, nx3158, nx3160, nx3170, nx3186, addr1_data_4, 
         nx3190, nx3196, bias_offset_data_out_4, nx3224, img_base_addr_4, nx3242, 
         nx3248, img_addr_offset_4, nx3256, nx3262, nx3270, 
         write_base_data_out_5, nx3294, nx3296, nx3298, nx3308, nx3312, nx3318, 
         nx3326, addr1_data_5, nx3354, bias_offset_data_out_5, nx3362, nx3364, 
         nx3374, img_base_addr_5, write_base_prev_data_out_5, nx3388, 
         img_addr_offset_5, nx3408, nx3410, nx3426, write_base_data_out_6, 
         nx3446, nx3448, nx3460, nx3466, addr1_data_6, nx3470, nx3476, 
         bias_offset_data_out_6, nx3504, img_base_addr_6, nx3522, nx3528, 
         img_addr_offset_6, nx3536, nx3542, nx3550, write_base_data_out_7, 
         nx3574, nx3576, nx3578, nx3588, nx3592, nx3598, nx3606, addr1_data_7, 
         nx3634, bias_offset_data_out_7, nx3642, nx3644, nx3654, img_base_addr_7, 
         write_base_prev_data_out_7, nx3668, img_addr_offset_7, nx3688, nx3690, 
         nx3706, write_base_data_out_8, nx3726, nx3728, nx3740, nx3746, 
         addr1_data_8, nx3750, nx3756, bias_offset_data_out_8, nx3784, 
         img_base_addr_8, nx3802, nx3808, img_addr_offset_8, nx3816, nx3822, 
         nx3830, write_base_data_out_9, nx3854, nx3856, nx3858, nx3868, nx3872, 
         nx3878, nx3886, addr1_data_9, nx3914, bias_offset_data_out_9, nx3922, 
         nx3924, nx3934, img_base_addr_9, write_base_prev_data_out_9, nx3948, 
         img_addr_offset_9, nx3968, nx3970, nx3986, write_base_data_out_10, 
         nx4006, nx4008, nx4020, nx4026, addr1_data_10, nx4030, nx4036, 
         bias_offset_data_out_10, nx4064, img_base_addr_10, nx4082, nx4088, 
         img_addr_offset_10, nx4096, nx4102, nx4110, write_base_data_out_11, 
         nx4134, nx4136, nx4138, nx4148, nx4152, nx4158, nx4166, addr1_data_11, 
         nx4194, bias_offset_data_out_11, nx4202, nx4204, nx4214, 
         img_base_addr_11, write_base_prev_data_out_11, nx4228, 
         img_addr_offset_11, nx4248, nx4250, nx4266, write_base_data_out_12, 
         nx4286, nx4288, nx4300, nx4306, addr1_data_12, nx4310, nx4316, 
         bias_offset_data_out_12, nx4344, img_base_addr_12, nx4362, nx4368, 
         img_addr_offset_12, nx4376, nx4382, nx4390, write_base_data_out_13, 
         nx4418, nx4428, nx4432, nx4438, nx4446, addr1_data_13, nx4474, 
         bias_offset_data_out_13, nx4482, nx4484, nx4494, img_base_addr_13, 
         write_base_prev_data_out_13, nx4508, img_addr_offset_13, nx4528, nx4530, 
         nx4546, write_base_data_out_14, nx4566, nx4568, nx4580, nx4586, 
         addr1_data_14, nx4590, nx4596, bias_offset_data_out_14, nx4624, 
         img_base_addr_14, nx4642, nx4648, img_addr_offset_14, nx4656, nx4662, 
         nx4670, nx4686, bias_offset_data_out_15, write_base_data_out_15, nx4714, 
         addr1_data_15, nx4734, nx4736, nx4744, nx4746, nx4756, img_base_addr_15, 
         write_base_prev_data_out_15, nx4764, nx4780, nx1479, nx1489, nx1499, 
         nx1509, nx1519, nx1529, nx1539, nx1549, nx1559, nx1569, nx1579, nx1589, 
         nx1599, nx1609, nx1619, nx1629, nx1639, nx1649, nx1659, nx1669, nx1679, 
         nx1689, nx1699, nx1709, nx1719, nx1729, nx1739, nx1749, nx1759, nx1769, 
         nx1779, nx1789, nx1799, nx1809, nx1819, nx1829, nx1839, nx1849, nx1859, 
         nx1869, nx1879, nx1889, nx1899, nx1909, nx1919, nx1929, nx1939, nx1949, 
         nx1959, nx1969, nx1979, nx1989, nx1999, nx2009, nx2019, nx2029, nx2039, 
         nx2049, nx2059, nx2069, nx2079, nx2089, nx2099, nx2109, nx2119, nx2129, 
         nx2139, nx2149, nx2159, nx2169, nx2179, nx2189, nx2199, nx2209, nx2219, 
         nx2229, nx2239, nx2249, nx2259, nx2269, nx2279, nx2289, nx2299, nx2309, 
         nx2319, nx2329, nx2339, nx2349, nx2359, nx2369, nx2379, nx2389, nx2399, 
         nx2409, nx2419, nx2429, nx2439, nx2449, nx2459, nx2469, nx2479, nx2489, 
         nx2499, nx2509, nx2519, nx2529, nx2539, nx2549, nx2559, nx2569, nx2579, 
         nx2589, nx2599, nx2609, nx2619, nx2629, nx2639, nx2649, nx2659, nx2669, 
         nx2679, nx2689, nx2699, nx2709, nx2719, nx2729, nx2739, nx2749, nx2759, 
         nx2769, nx2779, nx2789, nx2799, nx2809, nx2819, nx2829, nx2839, nx2849, 
         nx2859, nx2869, nx2879, nx2889, nx2899, nx2909, nx2919, nx2929, nx2939, 
         nx2949, nx2959, nx2969, nx2979, nx2989, nx2999, nx3009, nx3019, nx3029, 
         nx3039, nx3049, nx3059, nx3069, nx3079, nx3089, nx3099, nx3109, nx3119, 
         nx3129, nx3139, nx3149, nx3159, nx3169, nx3179, nx3189, nx3199, nx3209, 
         nx3219, nx3229, nx3239, nx3249, nx3259, nx3269, nx3279, nx3289, nx3299, 
         nx3309, nx3319, nx3329, nx3339, nx3349, nx3359, nx3369, nx3379, nx3389, 
         nx3399, nx3409, nx3419, nx3429, nx3439, nx3449, nx3459, nx3469, nx3479, 
         nx3489, nx3499, nx3509, nx3519, nx3529, nx3539, nx3549, nx3559, nx3569, 
         nx3579, nx3589, nx3599, nx3609, nx3619, nx3629, nx3639, nx3649, nx3659, 
         nx3669, nx3679, nx3689, nx3699, nx3709, nx3719, nx3729, nx3739, nx3749, 
         nx3759, nx3769, nx3779, nx3789, nx3799, nx3809, nx3819, nx3829, nx3839, 
         nx3849, nx3859, nx3869, nx3879, nx3889, nx3909, nx3919, nx3929, nx3939, 
         nx3957, nx3959, nx3967, nx3975, nx3979, nx3981, nx3989, nx3999, nx4004, 
         nx4009, nx4017, nx4019, nx4027, nx4031, nx4033, nx4039, nx4041, nx4043, 
         nx4045, nx4047, nx4053, nx4055, nx4057, nx4059, nx4065, nx4067, nx4069, 
         nx4073, nx4077, nx4080, nx4087, nx4099, nx4105, nx4109, nx4111, nx4115, 
         nx4119, nx4123, nx4129, nx4143, nx4149, nx4151, nx4153, nx4157, nx4163, 
         nx4167, nx4175, nx4180, nx4183, nx4191, nx4197, nx4200, nx4207, nx4213, 
         nx4217, nx4223, nx4229, nx4235, nx4239, nx4246, nx4251, nx4253, nx4257, 
         nx4265, nx4271, nx4277, nx4281, nx4284, nx4287, nx4293, nx4295, nx4299, 
         nx4301, nx4303, nx4305, nx4307, nx4314, nx4320, nx4321, nx4328, nx4335, 
         nx4337, nx4343, nx4349, nx4351, nx4358, nx4363, nx4365, nx4372, nx4377, 
         nx4379, nx4386, nx4391, nx4393, nx4400, nx4407, nx4408, nx4417, nx4423, 
         nx4427, nx4433, nx4435, nx4441, nx4447, nx4453, nx4459, nx4460, nx4465, 
         nx4469, nx4471, nx4480, nx4485, nx4487, nx4493, nx4497, nx4499, nx4503, 
         nx4507, nx4513, nx4515, nx4519, nx4526, nx4531, nx4533, nx4535, nx4543, 
         nx4553, nx4561, nx4563, nx4565, nx4571, nx4575, nx4579, nx4581, nx4583, 
         nx4589, nx4601, nx4609, nx4617, nx4621, nx4633, nx4635, nx4637, nx4638, 
         nx4647, nx4655, nx4657, nx4663, nx4669, nx4673, nx4681, nx4689, nx4692, 
         nx4701, nx4703, nx4705, nx4711, nx4717, nx4723, nx4725, nx4731, nx4735, 
         nx4743, nx4747, nx4751, nx4759, nx4761, nx4765, nx4767, nx4770, nx4776, 
         nx4781, nx4783, nx4787, nx4795, nx4801, nx4803, nx4807, nx4813, nx4819, 
         nx4821, nx4825, nx4833, nx4839, nx4841, nx4845, nx4853, nx4861, nx4879, 
         nx4881, nx4883, nx4895, nx4903, nx4911, nx4913, nx4927, nx4941, nx4957, 
         nx4961, nx4975, nx4977, nx4981, nx4993, nx4997, nx5009, nx5011, nx5013, 
         nx5019, nx5023, nx5031, nx5037, nx5041, nx5049, nx5055, nx5059, nx5067, 
         nx5072, nx5077, nx5083, nx5089, nx5099, nx5107, nx5113, nx5115, nx5122, 
         nx5128, nx5134, nx5137, nx5140, nx5142, nx5144, nx5146, nx5148, nx5155, 
         nx5157, nx5162, nx5164, nx5168, nx5188, nx5194, nx5197, nx5202, nx5204, 
         nx5206, nx5208, nx5216, nx5218, nx5243, nx5330, nx5334, nx5379, nx5383, 
         nx5386, nx5390, nx5393, nx5396, nx5399, nx5402, nx5405, nx5408, nx5411, 
         nx5414, nx5417, nx5420, nx5423, nx5426, nx5429, nx5432, nx5435, nx5438, 
         nx5441, nx5444, nx5447, nx5450, nx5453, nx5456, nx5459, nx5462, nx5465, 
         nx5468, nx5471, nx5474, nx5477, nx5480, nx5482, nx5501, nx5587, nx5593, 
         nx5596, nx5598, nx5605, nx5607, nx5611, nx5614, nx5616, nx5619, nx5621, 
         nx5629, nx5632, nx5636, nx5647, nx5651, nx5653, nx5657, nx5659, nx5662, 
         nx5664, nx5670, nx5673, nx5677, nx5679, nx5685, nx5687, nx5692, nx5696, 
         nx5698, nx5700, nx5703, nx5707, nx5709, nx5712, nx5714, nx5718, nx5720, 
         nx5722, nx5728, nx5731, nx5734, nx5737, nx5742, nx5747, nx5749, nx5758, 
         nx5762, nx5764, nx5767, nx5771, nx5773, nx5777, nx5783, nx5790, nx5794, 
         nx5805, nx5807, nx5809, nx5815, nx5820, nx5826, nx5829, nx5831, nx5834, 
         nx5836, nx5838, nx5843, nx5850, nx5853, nx5856, nx5859, nx5864, nx5869, 
         nx5871, nx5873, nx5876, nx5879, nx5882, nx5886, nx5888, nx5892, nx5895, 
         nx5900, nx5901, nx5906, nx5908, nx5913, nx5917, nx5921, nx5925, nx5936, 
         nx5938, nx5943, nx5945, nx5947, nx5951, nx5955, nx5957, nx5961, nx5963, 
         nx5965, nx5968, nx5971, nx5974, nx5977, nx5980, nx5983, nx5986, nx5991, 
         nx5996, nx5998, nx6000, nx6003, nx6006, nx6009, nx6013, nx6017, nx6020, 
         nx6025, nx6026, nx6031, nx6034, nx6037, nx6039, nx6042, nx6045, nx6049, 
         nx6060, nx6062, nx6067, nx6069, nx6071, nx6075, nx6079, nx6081, nx6085, 
         nx6088, nx6090, nx6097, nx6100, nx6103, nx6106, nx6109, nx6114, nx6119, 
         nx6121, nx6123, nx6126, nx6129, nx6132, nx6136, nx6140, nx6143, nx6148, 
         nx6149, nx6154, nx6157, nx6160, nx6162, nx6164, nx6167, nx6171, nx6182, 
         nx6184, nx6189, nx6191, nx6193, nx6197, nx6201, nx6203, nx6207, nx6210, 
         nx6212, nx6219, nx6222, nx6225, nx6228, nx6231, nx6236, nx6241, nx6243, 
         nx6245, nx6248, nx6251, nx6254, nx6258, nx6262, nx6265, nx6270, nx6271, 
         nx6276, nx6279, nx6282, nx6284, nx6286, nx6289, nx6293, nx6304, nx6306, 
         nx6311, nx6313, nx6315, nx6319, nx6323, nx6325, nx6329, nx6332, nx6334, 
         nx6341, nx6344, nx6347, nx6350, nx6353, nx6358, nx6363, nx6365, nx6367, 
         nx6373, nx6376, nx6380, nx6384, nx6387, nx6392, nx6393, nx6398, nx6400, 
         nx6402, nx6404, nx6408, nx6411, nx6415, nx6426, nx6428, nx6433, nx6435, 
         nx6437, nx6441, nx6445, nx6447, nx6451, nx6454, nx6456, nx6463, nx6466, 
         nx6469, nx6472, nx6475, nx6484, nx6486, nx6493, nx6494, nx6496, nx6500, 
         nx6502, nx6505, nx6510, nx6511, nx6516, nx6518, nx6520, nx6524, nx6527, 
         nx6532, nx6543, nx6555, nx6558, nx6560, nx6563, nx6569, nx6572, nx6576, 
         nx6580, nx6583, nx6586, nx6589, nx6592, nx6599, nx6601, nx6603, nx6605, 
         nx6607, nx6609, nx6611, nx6613, nx6615, nx6617, nx6619, nx6621, nx6623, 
         nx6625, nx6627, nx6629, nx6631, nx6633, nx6635, nx6637, nx6639, nx6641, 
         nx6643, nx6651, nx6653, nx6655, nx6657, nx6659, nx6663, nx6665, nx6667, 
         nx6673, nx6675, nx6677, nx6679, nx6681, nx6683, nx6685, nx6687, nx6689, 
         nx6691, nx6693, nx6695, nx6699, nx6705, nx6713, nx6721, nx6723, nx6725, 
         nx6727, nx6729, nx6731, nx6733, nx6735, nx6737, nx6739, nx6741, nx6743, 
         nx6749, nx6759, nx6761, nx6763, nx6765, nx6767, nx6769, nx6771, nx6773, 
         nx6781, nx6787, nx6793, nx6795, nx6797, nx6799, nx6801, nx6803, nx6805, 
         nx6807, nx6809, nx6811, nx6813, nx6815, nx6817, nx6819, nx6821, nx6823, 
         nx6825, nx6827, nx6829, nx6831, nx6833, nx6835, nx6837, nx6839, nx6851, 
         nx6855, nx6857, nx6859, nx6871, nx6897, nx6899, nx6901, nx6903, nx6905, 
         nx6927, nx6929, nx6931, nx6933, nx6939, nx6941, nx6943, nx6945, nx6947, 
         nx6949, nx6951, nx6953, nx6955, nx6957, nx6959, nx6961, nx6963, nx6965, 
         nx6967, nx6969, nx6971, nx6973, nx6975, nx6977, nx6979, nx6981, nx6983, 
         nx6985, nx6987, nx6989, nx6991, nx6993, nx6995, nx6997, nx6999, nx7001, 
         nx7003, nx7005, nx7007, nx7009, nx7011, nx7013, nx7015, nx7017, nx7019, 
         nx7021, nx7023, nx7025, nx7027, nx7033, nx7035, nx7037, nx7039, nx7041, 
         nx7043, nx7049, nx7051, nx7053, nx7055, nx7057, nx7059, nx7061, nx7065, 
         nx7071, nx7073, nx7075, nx7077, nx7079, nx7081, nx7083, nx7085, nx7087, 
         nx7089, nx7091, nx7093, nx7095, nx7097, nx7099, nx7101, nx7103, nx7105, 
         nx7107, nx7109, nx7111, nx7113, nx7115, nx7117, nx7119, nx7121, nx7123, 
         nx7125, nx7127, nx7129, nx7131, nx7133, nx7135, nx7137, nx7139, nx7145, 
         nx7029, nx4593, nx4665, nx7063, nx7031, nx6711, nx7293, nx7294, nx7295, 
         nx7296, nx7297, nx7298, nx7299, nx7300, nx7301, nx7302, nx7303, nx7304, 
         nx7305, nx3899, nx7306, nx7307, nx6488, nx7308, nx7309, nx6491, nx4414, 
         nx7310, nx7311, nx6370, nx7312, nx7313, nx7314, nx7315, nx7316, nx7317, 
         nx7318, nx7319, nx7320, nx7321, nx7322, nx3002, nx7323, nx5751, nx5754, 
         nx5689, nx7324, nx5191, argmax_ready_dup0, nx7325, nx7326, nx7327, 
         nx7328, nx1930, nx7329, nx7330, nx7331, nx7332, nx7333, nx7334, nx7335, 
         nx5847, nx7336, nx7337, nx2850, nx5667, nx5725, nx6775, nx7047, nx7338, 
         nx7339, nx7340, argmax_ready_XX0_XREP5, nx7341, nx7342, nx7343, nx7344, 
         nx7345, nx7346, nx7347, nx7348, nx7349, nx7350, nx7351, nx7352, nx7353, 
         NOT_nx4700, nx7354, nx7355, nx7356, nx7357, nx7358, nx7359, nx7360, 
         nx7361, nx7362, nx7363, nx7364, nx7365, nx7366, nx7367, nx7445;
    wire [138:0] \$dummy ;




    assign wind_rst = io_done_out ;
    assign filter_reset = io_done_out ;
    Cache_5_16_28_5 img_cache (.in_word ({cache_data_in_15,cache_data_in_14,
                    cache_data_in_13,cache_data_in_12,cache_data_in_11,
                    cache_data_in_10,cache_data_in_9,cache_data_in_8,
                    cache_data_in_7,cache_data_in_6,cache_data_in_5,
                    cache_data_in_4,cache_data_in_3,cache_data_in_2,
                    cache_data_in_1,cache_data_in_0}), .cache_in_sel ({nx6611,
                    cache_width_count_3,nx6615,cache_width_count_1,
                    cache_width_count_0}), .cache_out_sel ({wind_width_count_4,
                    wind_width_count_3,wind_width_count_2,wind_width_count_1,
                    nx6607}), .decoder_enable (cache_load), .out_column_0__15 (
                    cache_data_out_4__15), .out_column_0__14 (
                    cache_data_out_4__14), .out_column_0__13 (
                    cache_data_out_4__13), .out_column_0__12 (
                    cache_data_out_4__12), .out_column_0__11 (
                    cache_data_out_4__11), .out_column_0__10 (
                    cache_data_out_4__10), .out_column_0__9 (cache_data_out_4__9
                    ), .out_column_0__8 (cache_data_out_4__8), .out_column_0__7 (
                    cache_data_out_4__7), .out_column_0__6 (cache_data_out_4__6)
                    , .out_column_0__5 (cache_data_out_4__5), .out_column_0__4 (
                    cache_data_out_4__4), .out_column_0__3 (cache_data_out_4__3)
                    , .out_column_0__2 (cache_data_out_4__2), .out_column_0__1 (
                    cache_data_out_4__1), .out_column_0__0 (cache_data_out_4__0)
                    , .out_column_1__15 (cache_data_out_3__15), .out_column_1__14 (
                    cache_data_out_3__14), .out_column_1__13 (
                    cache_data_out_3__13), .out_column_1__12 (
                    cache_data_out_3__12), .out_column_1__11 (
                    cache_data_out_3__11), .out_column_1__10 (
                    cache_data_out_3__10), .out_column_1__9 (cache_data_out_3__9
                    ), .out_column_1__8 (cache_data_out_3__8), .out_column_1__7 (
                    cache_data_out_3__7), .out_column_1__6 (cache_data_out_3__6)
                    , .out_column_1__5 (cache_data_out_3__5), .out_column_1__4 (
                    cache_data_out_3__4), .out_column_1__3 (cache_data_out_3__3)
                    , .out_column_1__2 (cache_data_out_3__2), .out_column_1__1 (
                    cache_data_out_3__1), .out_column_1__0 (cache_data_out_3__0)
                    , .out_column_2__15 (cache_data_out_2__15), .out_column_2__14 (
                    cache_data_out_2__14), .out_column_2__13 (
                    cache_data_out_2__13), .out_column_2__12 (
                    cache_data_out_2__12), .out_column_2__11 (
                    cache_data_out_2__11), .out_column_2__10 (
                    cache_data_out_2__10), .out_column_2__9 (cache_data_out_2__9
                    ), .out_column_2__8 (cache_data_out_2__8), .out_column_2__7 (
                    cache_data_out_2__7), .out_column_2__6 (cache_data_out_2__6)
                    , .out_column_2__5 (cache_data_out_2__5), .out_column_2__4 (
                    cache_data_out_2__4), .out_column_2__3 (cache_data_out_2__3)
                    , .out_column_2__2 (cache_data_out_2__2), .out_column_2__1 (
                    cache_data_out_2__1), .out_column_2__0 (cache_data_out_2__0)
                    , .out_column_3__15 (cache_data_out_1__15), .out_column_3__14 (
                    cache_data_out_1__14), .out_column_3__13 (
                    cache_data_out_1__13), .out_column_3__12 (
                    cache_data_out_1__12), .out_column_3__11 (
                    cache_data_out_1__11), .out_column_3__10 (
                    cache_data_out_1__10), .out_column_3__9 (cache_data_out_1__9
                    ), .out_column_3__8 (cache_data_out_1__8), .out_column_3__7 (
                    cache_data_out_1__7), .out_column_3__6 (cache_data_out_1__6)
                    , .out_column_3__5 (cache_data_out_1__5), .out_column_3__4 (
                    cache_data_out_1__4), .out_column_3__3 (cache_data_out_1__3)
                    , .out_column_3__2 (cache_data_out_1__2), .out_column_3__1 (
                    cache_data_out_1__1), .out_column_3__0 (cache_data_out_1__0)
                    , .out_column_4__15 (cache_data_out_0__15), .out_column_4__14 (
                    cache_data_out_0__14), .out_column_4__13 (
                    cache_data_out_0__13), .out_column_4__12 (
                    cache_data_out_0__12), .out_column_4__11 (
                    cache_data_out_0__11), .out_column_4__10 (
                    cache_data_out_0__10), .out_column_4__9 (cache_data_out_0__9
                    ), .out_column_4__8 (cache_data_out_0__8), .out_column_4__7 (
                    cache_data_out_0__7), .out_column_4__6 (cache_data_out_0__6)
                    , .out_column_4__5 (cache_data_out_0__5), .out_column_4__4 (
                    cache_data_out_0__4), .out_column_4__3 (cache_data_out_0__3)
                    , .out_column_4__2 (cache_data_out_0__2), .out_column_4__1 (
                    cache_data_out_0__1), .out_column_4__0 (cache_data_out_0__0)
                    , .clk (nx6619), .reset (cache_rst_actual)) ;
    AdvancedCounter_16 cache_height_cntr (.clk (clk), .reset (nx6601), .enable (
                       cache_height_count_en), .mode_in ({io_done_out,
                       io_done_out}), .max_val_in ({io_done_out,io_done_out,
                       io_done_out,io_done_out,io_done_out,io_done_out,
                       io_done_out,io_done_out,io_done_out,io_done_out,
                       io_done_out,max_height_4,max_height_3,max_height_2,
                       max_height_1,max_height_0}), .max_reached_out (
                       cache_height_ended), .counter_out ({\$dummy [0],
                       \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],
                       \$dummy [5],\$dummy [6],\$dummy [7],\$dummy [8],
                       \$dummy [9],\$dummy [10],\$dummy [11],\$dummy [12],
                       \$dummy [13],\$dummy [14],\$dummy [15]})) ;
    fake_gnd ix1260 (.Y (io_done_out)) ;
    ao22 ix2001 (.Y (mem_data_out[4]), .A0 (comp_unit_data2_in[4]), .A1 (nx6673)
         , .B0 (comp_unit_data1_in[4]), .B1 (nx6679)) ;
    nand02 ix1487 (.Y (nx1486), .A0 (nx3957), .A1 (nx5011)) ;
    aoi32 ix3958 (.Y (nx3957), .A0 (nx3959), .A1 (comp_unit_finished), .A2 (
          current_state_19), .B0 (nx4563), .B1 (nx1459)) ;
    dffr layer_type_reg_q_0 (.Q (comp_unit_operation), .QB (\$dummy [16]), .D (
         nx1519), .CLK (clk), .R (reset)) ;
    mux21_ni ix1520 (.Y (nx1519), .A0 (nx6927), .A1 (mem_data_in[0]), .S0 (
             current_state_3)) ;
    dffr reg_current_state_3 (.Q (current_state_3), .QB (\$dummy [17]), .D (
         nx1461), .CLK (nx6627), .R (reset)) ;
    dffr reg_current_state_2 (.Q (current_state_2), .QB (nx3967), .D (nx1578), .CLK (
         nx6619), .R (reset)) ;
    oai21 ix1573 (.Y (nx1572), .A0 (io_ready_in), .A1 (nx3975), .B0 (nx3979)) ;
    dffr reg_current_state_1 (.Q (\$dummy [18]), .QB (nx3975), .D (nx1572), .CLK (
         nx6619), .R (reset)) ;
    dffs_ni reg_current_state_0 (.Q (\$dummy [19]), .QB (nx3979), .D (
            io_done_out), .CLK (nx6619), .S (reset)) ;
    nand02 ix1737 (.Y (nx1409), .A0 (nx3989), .A1 (nx4503)) ;
    mux21_ni ix2470 (.Y (nx2469), .A0 (nx1620), .A1 (num_channels_out_0), .S0 (
             nx4115)) ;
    nand03 ix1611 (.Y (nx1610), .A0 (nx3999), .A1 (nx4105), .A2 (nx3967)) ;
    oai21 ix4000 (.Y (nx3999), .A0 (nx1602), .A1 (current_state_25), .B0 (
          max_num_channels_data_out_0)) ;
    mux21_ni ix2590 (.Y (nx2589), .A0 (layer_type_out_1), .A1 (mem_data_in[1]), 
             .S0 (current_state_3)) ;
    dffr layer_type_reg_q_1 (.Q (layer_type_out_1), .QB (nx4004), .D (nx2589), .CLK (
         clk), .R (reset)) ;
    dffr reg_current_state_26 (.Q (\$dummy [20]), .QB (nx3981), .D (nx1800), .CLK (
         nx6619), .R (reset)) ;
    dffr reg_current_state_25 (.Q (current_state_25), .QB (nx4073), .D (nx112), 
         .CLK (nx6619), .R (reset)) ;
    oai32 ix1480 (.Y (nx1479), .A0 (nx4019), .A1 (nx6689), .A2 (current_state_25
          ), .B0 (nx4027), .B1 (nx7017)) ;
    dffr reg_current_state_4 (.Q (current_state_4), .QB (\$dummy [21]), .D (
         current_state_3), .CLK (nx6619), .R (reset)) ;
    dffr reg_nflt_layer_out_0 (.Q (nflt_layer_out_0), .QB (nx4019), .D (nx1479)
         , .CLK (clk), .R (reset)) ;
    inv01 ix4032 (.Y (nx4031), .A (mem_data_in[0])) ;
    oai32 ix1490 (.Y (nx1489), .A0 (nx4039), .A1 (nx6689), .A2 (current_state_25
          ), .B0 (nx4041), .B1 (nx7017)) ;
    dffr reg_nflt_layer_out_1 (.Q (nflt_layer_out_1), .QB (nx4039), .D (nx1489)
         , .CLK (clk), .R (reset)) ;
    mux21_ni ix4042 (.Y (nx4041), .A0 (nx4043), .A1 (nx4047), .S0 (nx6689)) ;
    aoi21 ix4044 (.Y (nx4043), .A0 (nflt_layer_out_1), .A1 (nflt_layer_out_0), .B0 (
          nx4045)) ;
    inv01 ix4048 (.Y (nx4047), .A (mem_data_in[1])) ;
    oai32 ix1500 (.Y (nx1499), .A0 (nx4053), .A1 (nx6689), .A2 (current_state_25
          ), .B0 (nx4055), .B1 (nx7017)) ;
    dffr nflt_layer_out_2 (.Q (\$dummy [22]), .QB (nx4053), .D (nx1499), .CLK (
         clk), .R (reset)) ;
    mux21_ni ix4056 (.Y (nx4055), .A0 (nx4057), .A1 (nx4059), .S0 (nx6689)) ;
    inv01 ix4060 (.Y (nx4059), .A (mem_data_in[2])) ;
    dffr reg_nflt_layer_out_3 (.Q (nflt_layer_out_3), .QB (\$dummy [23]), .D (
         nx1509), .CLK (clk), .R (reset)) ;
    mux21_ni ix1510 (.Y (nx1509), .A0 (nx98), .A1 (nflt_layer_out_3), .S0 (
             nx7017)) ;
    mux21 ix99 (.Y (nx98), .A0 (nx4065), .A1 (nx4069), .S0 (nx6691)) ;
    xnor2 ix4066 (.Y (nx4065), .A0 (nflt_layer_out_3), .A1 (nx4067)) ;
    inv01 ix4070 (.Y (nx4069), .A (mem_data_in[3])) ;
    oai222 ix2460 (.Y (nx2459), .A0 (nx4077), .A1 (nx1594), .B0 (nx4099), .B1 (
           nx7019), .C0 (nx4031), .C1 (nx6821)) ;
    dffs_ni max_num_channels_inst_reg_q_0 (.Q (max_num_channels_data_out_0), .QB (
            nx4077), .D (nx2459), .CLK (clk), .S (reset)) ;
    nand02 ix1595 (.Y (nx1594), .A0 (nx7019), .A1 (nx6821)) ;
    dffr reg_current_state_9 (.Q (current_state_9), .QB (\$dummy [24]), .D (
         nx136), .CLK (nx6621), .R (reset)) ;
    nor03_2x ix137 (.Y (nx136), .A0 (nx4087), .A1 (nx6927), .A2 (nx4004)) ;
    dffr reg_current_state_8 (.Q (current_state_8), .QB (nx4087), .D (nx6699), .CLK (
         nx6621), .R (reset)) ;
    dffr reg_current_state_7 (.Q (current_state_7), .QB (\$dummy [25]), .D (
         current_state_6), .CLK (nx6621), .R (reset)) ;
    dffr reg_current_state_6 (.Q (current_state_6), .QB (\$dummy [26]), .D (
         current_state_5), .CLK (nx6621), .R (reset)) ;
    dffr reg_current_state_5 (.Q (current_state_5), .QB (\$dummy [27]), .D (
         nx6691), .CLK (nx6621), .R (reset)) ;
    mux21_ni ix2450 (.Y (nx2449), .A0 (nflt_layer_temp_0), .A1 (mem_data_in[0])
             , .S0 (nx6691)) ;
    dffr nflt_layer_total_reg_q_0 (.Q (nflt_layer_temp_0), .QB (nx4099), .D (
         nx2449), .CLK (clk), .R (reset)) ;
    aoi22 ix4106 (.Y (nx4105), .A0 (mem_data_in[0]), .A1 (nx6693), .B0 (
          nflt_layer_temp_0), .B1 (nx1528)) ;
    dffr reg_num_channels_out_0 (.Q (num_channels_out_0), .QB (nx4111), .D (
         nx2469), .CLK (clk), .R (reset)) ;
    nor02_2x ix4116 (.Y (nx4115), .A0 (nx1516), .A1 (nx1421)) ;
    nor02ii ix1513 (.Y (nx1421), .A0 (nx4123), .A1 (nx1409)) ;
    nand02 ix4124 (.Y (nx4123), .A0 (current_state_24), .A1 (nx4153)) ;
    dffr reg_current_state_24 (.Q (current_state_24), .QB (nx4151), .D (nx1502)
         , .CLK (nx6623), .R (reset)) ;
    oai21 ix1503 (.Y (nx1502), .A0 (nx4129), .A1 (nx6641), .B0 (nx4149)) ;
    dffr reg_current_state_22 (.Q (\$dummy [28]), .QB (nx4129), .D (nx1486), .CLK (
         nx6621), .R (reset)) ;
    mux21_ni ix1590 (.Y (nx1589), .A0 (flt_size_out_0), .A1 (mem_data_in[0]), .S0 (
             current_state_5)) ;
    dffr flt_size_reg_q_0 (.Q (flt_size_out_0), .QB (\$dummy [29]), .D (nx1589)
         , .CLK (clk), .R (reset)) ;
    dffr flt_size_reg_q_2 (.Q (flt_size_out_2), .QB (nx4143), .D (nx1599), .CLK (
         clk), .R (reset)) ;
    mux21_ni ix1600 (.Y (nx1599), .A0 (flt_size_out_2), .A1 (mem_data_in[2]), .S0 (
             current_state_5)) ;
    mux21_ni ix1610 (.Y (nx1609), .A0 (flt_size_out_1), .A1 (mem_data_in[1]), .S0 (
             current_state_5)) ;
    dffr flt_size_reg_q_1 (.Q (flt_size_out_1), .QB (\$dummy [30]), .D (nx1609)
         , .CLK (clk), .R (reset)) ;
    dffr reg_current_state_23 (.Q (\$dummy [31]), .QB (nx4149), .D (nx1492), .CLK (
         nx6621), .R (reset)) ;
    nor04 ix4154 (.Y (nx4153), .A0 (nx1098), .A1 (nx1010), .A2 (nx914), .A3 (
          nx820)) ;
    nand04 ix1099 (.Y (nx1098), .A0 (nx4157), .A1 (nx4314), .A2 (nx4321), .A3 (
           nx4328)) ;
    oai22 ix2210 (.Y (nx2209), .A0 (nx4163), .A1 (nx6833), .B0 (nx4307), .B1 (
          nx6735)) ;
    dffr reg_write_offset_reg_q_14 (.Q (write_offset_data_out_14), .QB (nx4167)
         , .D (nx2189), .CLK (nx6623), .R (reset)) ;
    nand02 ix4176 (.Y (nx4175), .A0 (write_offset_data_out_13), .A1 (nx1012)) ;
    oai22 ix2170 (.Y (nx2169), .A0 (nx4180), .A1 (nx6833), .B0 (nx4305), .B1 (
          nx6733)) ;
    oai21 ix4181 (.Y (nx4180), .A0 (nx1012), .A1 (write_offset_data_out_13), .B0 (
          nx4175)) ;
    dffr reg_write_offset_reg_q_12 (.Q (write_offset_data_out_12), .QB (nx4183)
         , .D (nx2149), .CLK (nx6623), .R (reset)) ;
    nand02 ix4192 (.Y (nx4191), .A0 (write_offset_data_out_11), .A1 (nx964)) ;
    oai22 ix2130 (.Y (nx2129), .A0 (nx4197), .A1 (nx6831), .B0 (nx4303), .B1 (
          nx6733)) ;
    oai21 ix4198 (.Y (nx4197), .A0 (nx964), .A1 (write_offset_data_out_11), .B0 (
          nx4191)) ;
    dffr reg_write_offset_reg_q_10 (.Q (write_offset_data_out_10), .QB (nx4200)
         , .D (nx2109), .CLK (nx6623), .R (reset)) ;
    nand02 ix4208 (.Y (nx4207), .A0 (write_offset_data_out_9), .A1 (nx918)) ;
    oai22 ix2090 (.Y (nx2089), .A0 (nx4213), .A1 (nx6831), .B0 (nx4301), .B1 (
          nx6733)) ;
    oai21 ix4214 (.Y (nx4213), .A0 (nx918), .A1 (write_offset_data_out_9), .B0 (
          nx4207)) ;
    dffr reg_write_offset_reg_q_8 (.Q (write_offset_data_out_8), .QB (nx4217), .D (
         nx2069), .CLK (nx6623), .R (reset)) ;
    nand02 ix4224 (.Y (nx4223), .A0 (write_offset_data_out_7), .A1 (nx868)) ;
    oai22 ix2050 (.Y (nx2049), .A0 (nx4229), .A1 (nx6731), .B0 (nx4235), .B1 (
          nx6831)) ;
    dffr reg_write_offset_reg_q_7 (.Q (write_offset_data_out_7), .QB (nx4229), .D (
         nx2049), .CLK (nx6623), .R (reset)) ;
    oai21 ix4236 (.Y (nx4235), .A0 (nx868), .A1 (write_offset_data_out_7), .B0 (
          nx4223)) ;
    dffr reg_write_offset_reg_q_6 (.Q (write_offset_data_out_6), .QB (nx4239), .D (
         nx2029), .CLK (nx6623), .R (reset)) ;
    nand02 ix4247 (.Y (nx4246), .A0 (write_offset_data_out_5), .A1 (nx822)) ;
    oai22 ix2010 (.Y (nx2009), .A0 (nx4251), .A1 (nx6731), .B0 (nx4253), .B1 (
          nx6829)) ;
    dffr reg_write_offset_reg_q_5 (.Q (write_offset_data_out_5), .QB (nx4251), .D (
         nx2009), .CLK (nx6625), .R (reset)) ;
    oai21 ix4254 (.Y (nx4253), .A0 (nx822), .A1 (write_offset_data_out_5), .B0 (
          nx4246)) ;
    dffr reg_write_offset_reg_q_4 (.Q (write_offset_data_out_4), .QB (nx4257), .D (
         nx1989), .CLK (nx6625), .R (reset)) ;
    dffr reg_write_offset_reg_q_3 (.Q (write_offset_data_out_3), .QB (nx4271), .D (
         nx1969), .CLK (nx6625), .R (reset)) ;
    oai22 ix1950 (.Y (nx1949), .A0 (nx4277), .A1 (nx6731), .B0 (nx4281), .B1 (
          nx6829)) ;
    oai21 ix4282 (.Y (nx4281), .A0 (nx750), .A1 (write_offset_data_out_2), .B0 (
          nx4299)) ;
    oai22 ix1930 (.Y (nx1929), .A0 (nx7355), .A1 (nx6731), .B0 (nx4287), .B1 (
          nx6829)) ;
    oai21 ix4288 (.Y (nx4287), .A0 (write_offset_data_out_0), .A1 (
          write_offset_data_out_1), .B0 (nx4295)) ;
    dffr reg_write_offset_reg_q_0 (.Q (write_offset_data_out_0), .QB (nx4293), .D (
         nx1909), .CLK (nx6625), .R (reset)) ;
    dffr reg_write_offset_reg_q_1 (.Q (write_offset_data_out_1), .QB (nx4284), .D (
         nx1929), .CLK (nx6625), .R (reset)) ;
    dffr reg_write_offset_reg_q_2 (.Q (write_offset_data_out_2), .QB (nx4277), .D (
         nx1949), .CLK (nx6625), .R (reset)) ;
    dffr reg_write_offset_reg_q_9 (.Q (write_offset_data_out_9), .QB (nx4301), .D (
         nx2089), .CLK (nx6625), .R (reset)) ;
    dffr reg_write_offset_reg_q_11 (.Q (write_offset_data_out_11), .QB (nx4303)
         , .D (nx2129), .CLK (nx6627), .R (reset)) ;
    dffr reg_write_offset_reg_q_13 (.Q (write_offset_data_out_13), .QB (nx4305)
         , .D (nx2169), .CLK (nx6627), .R (reset)) ;
    dffr reg_write_offset_reg_q_15 (.Q (write_offset_data_out_15), .QB (nx4307)
         , .D (nx2209), .CLK (nx6627), .R (reset)) ;
    dffr new_size_squared_reg_q_15 (.Q (new_size_squared_out_15), .QB (
         \$dummy [32]), .D (nx2219), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_14 (.Q (new_size_squared_out_14), .QB (nx4320), 
         .D (nx2199), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_13 (.Q (new_size_squared_out_13), .QB (
         \$dummy [33]), .D (nx2179), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_12 (.Q (new_size_squared_out_12), .QB (nx4335), 
         .D (nx2159), .CLK (clk), .R (reset)) ;
    nand04 ix1011 (.Y (nx1010), .A0 (nx4337), .A1 (nx4343), .A2 (nx4351), .A3 (
           nx4358)) ;
    dffr new_size_squared_reg_q_11 (.Q (new_size_squared_out_11), .QB (
         \$dummy [34]), .D (nx2139), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_10 (.Q (new_size_squared_out_10), .QB (nx4349), 
         .D (nx2119), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_9 (.Q (new_size_squared_out_9), .QB (
         \$dummy [35]), .D (nx2099), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_8 (.Q (new_size_squared_out_8), .QB (nx4363), .D (
         nx2079), .CLK (clk), .R (reset)) ;
    nand04 ix915 (.Y (nx914), .A0 (nx4365), .A1 (nx4372), .A2 (nx4379), .A3 (
           nx4386)) ;
    dffr new_size_squared_reg_q_7 (.Q (new_size_squared_out_7), .QB (
         \$dummy [36]), .D (nx2059), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_6 (.Q (new_size_squared_out_6), .QB (nx4377), .D (
         nx2039), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_5 (.Q (new_size_squared_out_5), .QB (
         \$dummy [37]), .D (nx2019), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_4 (.Q (new_size_squared_out_4), .QB (nx4391), .D (
         nx1999), .CLK (clk), .R (reset)) ;
    nand04 ix821 (.Y (nx820), .A0 (nx4393), .A1 (nx4400), .A2 (nx4408), .A3 (
           nx4417)) ;
    dffr new_size_squared_reg_q_3 (.Q (new_size_squared_out_3), .QB (
         \$dummy [38]), .D (nx1979), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_2 (.Q (new_size_squared_out_2), .QB (nx4407), .D (
         nx1959), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_1 (.Q (new_size_squared_out_1), .QB (
         \$dummy [39]), .D (nx1939), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_0 (.Q (new_size_squared_out_0), .QB (nx4423), .D (
         nx1919), .CLK (clk), .R (reset)) ;
    dffr reg_num_channels_out_1 (.Q (num_channels_out_1), .QB (nx4447), .D (
         nx2489), .CLK (clk), .R (reset)) ;
    mux21_ni ix2490 (.Y (nx2489), .A0 (nx1652), .A1 (num_channels_out_1), .S0 (
             nx4115)) ;
    oai21 ix1653 (.Y (nx1652), .A0 (nx4427), .A1 (nx6825), .B0 (nx4435)) ;
    aoi22 ix4428 (.Y (nx4427), .A0 (mem_data_in[1]), .A1 (nx6693), .B0 (
          nflt_layer_temp_1), .B1 (nx1528)) ;
    dffr nflt_layer_total_reg_q_1 (.Q (nflt_layer_temp_1), .QB (nx4433), .D (
         nx2439), .CLK (clk), .R (reset)) ;
    mux21_ni ix2440 (.Y (nx2439), .A0 (nflt_layer_temp_1), .A1 (mem_data_in[1])
             , .S0 (nx6691)) ;
    aoi22 ix4436 (.Y (nx4435), .A0 (max_num_channels_data_out_1), .A1 (nx1646), 
          .B0 (nx6825), .B1 (nx1630)) ;
    oai222 ix2480 (.Y (nx2479), .A0 (nx4441), .A1 (nx1594), .B0 (nx4433), .B1 (
           nx7019), .C0 (nx4047), .C1 (nx6821)) ;
    dffr max_num_channels_inst_reg_q_1 (.Q (max_num_channels_data_out_1), .QB (
         nx4441), .D (nx2479), .CLK (clk), .R (reset)) ;
    oai21 ix1647 (.Y (nx1646), .A0 (nx7009), .A1 (nx6705), .B0 (nx4073)) ;
    mux21_ni ix2510 (.Y (nx2509), .A0 (nx1678), .A1 (num_channels_out_2), .S0 (
             nx4115)) ;
    oai21 ix1679 (.Y (nx1678), .A0 (nx4453), .A1 (nx6825), .B0 (nx4460)) ;
    aoi22 ix4454 (.Y (nx4453), .A0 (mem_data_in[2]), .A1 (nx6693), .B0 (
          nflt_layer_temp_2), .B1 (nx1528)) ;
    dffr nflt_layer_total_reg_q_2 (.Q (nflt_layer_temp_2), .QB (nx4459), .D (
         nx2429), .CLK (clk), .R (reset)) ;
    mux21_ni ix2430 (.Y (nx2429), .A0 (nflt_layer_temp_2), .A1 (mem_data_in[2])
             , .S0 (nx6691)) ;
    aoi22 ix4461 (.Y (nx4460), .A0 (max_num_channels_data_out_2), .A1 (nx1646), 
          .B0 (nx6825), .B1 (nx1664)) ;
    oai222 ix2500 (.Y (nx2499), .A0 (nx4465), .A1 (nx1594), .B0 (nx4459), .B1 (
           nx7019), .C0 (nx4059), .C1 (nx6821)) ;
    dffr max_num_channels_inst_reg_q_2 (.Q (max_num_channels_data_out_2), .QB (
         nx4465), .D (nx2499), .CLK (clk), .R (reset)) ;
    oai21 ix1665 (.Y (nx1664), .A0 (nx4469), .A1 (nx4471), .B0 (nx1464)) ;
    dffr reg_num_channels_out_2 (.Q (num_channels_out_2), .QB (nx4469), .D (
         nx2509), .CLK (clk), .R (reset)) ;
    mux21_ni ix2530 (.Y (nx2529), .A0 (nx1704), .A1 (num_channels_out_3), .S0 (
             nx4115)) ;
    oai21 ix1705 (.Y (nx1704), .A0 (nx4480), .A1 (nx6825), .B0 (nx4487)) ;
    aoi22 ix4481 (.Y (nx4480), .A0 (mem_data_in[3]), .A1 (nx6693), .B0 (
          nflt_layer_temp_3), .B1 (nx1528)) ;
    dffr nflt_layer_total_reg_q_3 (.Q (nflt_layer_temp_3), .QB (nx4485), .D (
         nx2419), .CLK (clk), .R (reset)) ;
    mux21_ni ix2420 (.Y (nx2419), .A0 (nflt_layer_temp_3), .A1 (mem_data_in[3])
             , .S0 (nx6691)) ;
    aoi22 ix4488 (.Y (nx4487), .A0 (max_num_channels_data_out_3), .A1 (nx1646), 
          .B0 (nx6825), .B1 (nx1690)) ;
    oai222 ix2520 (.Y (nx2519), .A0 (nx4493), .A1 (nx1594), .B0 (nx4485), .B1 (
           nx7019), .C0 (nx4069), .C1 (nx6821)) ;
    dffr max_num_channels_inst_reg_q_3 (.Q (max_num_channels_data_out_3), .QB (
         nx4493), .D (nx2519), .CLK (clk), .R (reset)) ;
    oai21 ix1691 (.Y (nx1690), .A0 (nx4497), .A1 (nx4499), .B0 (nx1463)) ;
    dffr reg_num_channels_out_3 (.Q (num_channels_out_3), .QB (nx4497), .D (
         nx2529), .CLK (clk), .R (reset)) ;
    dffr num_channels_out_4 (.Q (\$dummy [40]), .QB (nx4503), .D (nx2549), .CLK (
         clk), .R (reset)) ;
    mux21 ix2550 (.Y (nx2549), .A0 (nx4507), .A1 (nx4503), .S0 (nx4115)) ;
    aoi222 ix4508 (.Y (nx4507), .A0 (max_num_channels_data_out_4), .A1 (nx1646)
           , .B0 (mem_data_in[4]), .B1 (nx6693), .C0 (nx6827), .C1 (nx1716)) ;
    oai22 ix2540 (.Y (nx2539), .A0 (nx4513), .A1 (nx1594), .B0 (nx4515), .B1 (
          nx6821)) ;
    dffr max_num_channels_inst_reg_q_4 (.Q (max_num_channels_data_out_4), .QB (
         nx4513), .D (nx2539), .CLK (clk), .R (reset)) ;
    inv01 ix4516 (.Y (nx4515), .A (mem_data_in[4])) ;
    oai21 ix1717 (.Y (nx1716), .A0 (nx4503), .A1 (nx3989), .B0 (nx1409)) ;
    nor03_2x ix4520 (.Y (nx4519), .A0 (nlayers_counter_out_1), .A1 (
             nlayers_counter_out_2), .A2 (nx4531)) ;
    dffr reg_nlayers_counter_out_1 (.Q (nlayers_counter_out_1), .QB (
         \$dummy [41]), .D (nx2569), .CLK (clk), .R (reset)) ;
    mux21_ni ix2570 (.Y (nx2569), .A0 (nx1768), .A1 (nlayers_counter_out_1), .S0 (
             nx4009)) ;
    aoi21 ix4527 (.Y (nx4526), .A0 (nlayers_counter_out_1), .A1 (
          nlayers_counter_out_0), .B0 (nx4535)) ;
    oai32 ix2560 (.Y (nx2559), .A0 (nx4531), .A1 (current_state_2), .A2 (nx6665)
          , .B0 (nx4533), .B1 (nx4009)) ;
    dffr reg_nlayers_counter_out_0 (.Q (nlayers_counter_out_0), .QB (nx4531), .D (
         nx2559), .CLK (clk), .R (reset)) ;
    dffr reg_nlayers_counter_out_2 (.Q (nlayers_counter_out_2), .QB (
         \$dummy [42]), .D (nx2579), .CLK (clk), .R (reset)) ;
    mux21_ni ix2580 (.Y (nx2579), .A0 (nx1784), .A1 (nlayers_counter_out_2), .S0 (
             nx4009)) ;
    xnor2 ix4544 (.Y (nx4543), .A0 (nlayers_counter_out_2), .A1 (nx4535)) ;
    oai221 ix1469 (.Y (nx1468), .A0 (nx7023), .A1 (nx6643), .B0 (
           comp_unit_finished), .B1 (nx4581), .C0 (nx6851)) ;
    dffr reg_current_state_17 (.Q (\$dummy [43]), .QB (nx4553), .D (nx1446), .CLK (
         nx6633), .R (reset)) ;
    mux21 ix1900 (.Y (nx1899), .A0 (nx4561), .A1 (nx4583), .S0 (nx6835)) ;
    aoi32 ix4562 (.Y (nx4561), .A0 (nx4563), .A1 (ftc_cntrl_reg_out_11), .A2 (
          current_state_21), .B0 (ftc_cntrl_reg_out_8), .B1 (nx14)) ;
    mux21_ni ix1630 (.Y (nx1629), .A0 (nx332), .A1 (ftc_cntrl_reg_out_14), .S0 (
             nx6835)) ;
    oai22 ix333 (.Y (nx332), .A0 (nx4563), .A1 (nx4571), .B0 (nx4565), .B1 (
          nx5164)) ;
    oai321 ix1843 (.Y (nx1842), .A0 (nx3959), .A1 (nx4579), .A2 (nx4581), .B0 (
           nx4583), .B1 (nx4673), .C0 (nx5162)) ;
    inv01 ix4580 (.Y (nx4579), .A (comp_unit_finished)) ;
    dffr reg_current_state_19 (.Q (current_state_19), .QB (nx4581), .D (nx1468)
         , .CLK (nx6627), .R (reset)) ;
    dffr ftc_cntrl_reg_reg_q_8 (.Q (ftc_cntrl_reg_out_8), .QB (nx4583), .D (
         nx1899), .CLK (nx6627), .R (nx6601)) ;
    dffr reg_current_state_13 (.Q (current_state_13), .QB (\$dummy [44]), .D (
         nx300), .CLK (nx6629), .R (reset)) ;
    oai22 ix301 (.Y (nx300), .A0 (nx7029), .A1 (nx286), .B0 (nx4637), .B1 (
          nx6705)) ;
    dffr reg_cntr1_inst_counter_out_4 (.Q (cntr1_inst_counter_out_4), .QB (
         nx4647), .D (nx1569), .CLK (clk), .R (nx6713)) ;
    nand04 ix4602 (.Y (nx4601), .A0 (cntr1_inst_counter_out_3), .A1 (
           cntr1_inst_counter_out_2), .A2 (cntr1_inst_counter_out_1), .A3 (
           cntr1_inst_counter_out_0)) ;
    dffr reg_cntr1_inst_counter_out_3 (.Q (cntr1_inst_counter_out_3), .QB (
         \$dummy [45]), .D (nx1559), .CLK (clk), .R (nx6713)) ;
    xnor2 ix215 (.Y (nx214), .A0 (cntr1_inst_counter_out_3), .A1 (nx4609)) ;
    nand03 ix4610 (.Y (nx4609), .A0 (cntr1_inst_counter_out_2), .A1 (
           cntr1_inst_counter_out_1), .A2 (cntr1_inst_counter_out_0)) ;
    dffr reg_cntr1_inst_counter_out_2 (.Q (cntr1_inst_counter_out_2), .QB (
         \$dummy [46]), .D (nx1549), .CLK (clk), .R (nx6713)) ;
    xnor2 ix201 (.Y (nx200), .A0 (cntr1_inst_counter_out_2), .A1 (nx4617)) ;
    nand02 ix4618 (.Y (nx4617), .A0 (cntr1_inst_counter_out_1), .A1 (
           cntr1_inst_counter_out_0)) ;
    dffr reg_cntr1_inst_counter_out_1 (.Q (cntr1_inst_counter_out_1), .QB (
         nx4621), .D (nx1539), .CLK (clk), .R (nx6713)) ;
    dffr reg_current_state_10 (.Q (\$dummy [47]), .QB (nx4637), .D (nx152), .CLK (
         nx6629), .R (reset)) ;
    or02 ix153 (.Y (nx152), .A0 (nx1421), .A1 (current_state_12)) ;
    dffr reg_current_state_12 (.Q (current_state_12), .QB (nx4635), .D (nx146), 
         .CLK (nx6627), .R (reset)) ;
    nand03 ix147 (.Y (nx146), .A0 (nx4633), .A1 (nx6821), .A2 (nx4073)) ;
    oai21 ix4634 (.Y (nx4633), .A0 (nx6927), .A1 (nx4004), .B0 (current_state_8)
          ) ;
    oai21 ix4639 (.Y (nx4638), .A0 (cntr1_inst_counter_out_0), .A1 (
          cntr1_inst_counter_out_1), .B0 (nx4617)) ;
    dffr reg_cntr1_inst_counter_out_0 (.Q (cntr1_inst_counter_out_0), .QB (
         \$dummy [48]), .D (nx1529), .CLK (clk), .R (nx6713)) ;
    xnor2 ix1530 (.Y (nx1529), .A0 (cntr1_inst_counter_out_0), .A1 (nx7029)) ;
    dffr reg_current_state_11 (.Q (\$dummy [49]), .QB (nx4589), .D (nx6659), .CLK (
         nx6629), .R (reset)) ;
    dffr cntr1_inst_counter_out_5 (.Q (\$dummy [50]), .QB (nx4655), .D (nx1579)
         , .CLK (clk), .R (nx6713)) ;
    nand04 ix287 (.Y (nx286), .A0 (nx4669), .A1 (cntr1_inst_counter_out_0), .A2 (
           cntr1_inst_counter_out_3), .A3 (nx4663)) ;
    nor03_2x ix4670 (.Y (nx4669), .A0 (nx280), .A1 (nx248), .A2 (nx246)) ;
    mux21 ix2410 (.Y (nx2409), .A0 (nx4681), .A1 (nx4705), .S0 (nx6835)) ;
    nand04 ix4682 (.Y (nx4681), .A0 (nx1370), .A1 (nx1384), .A2 (nx1402), .A3 (
           nx1424)) ;
    dffr reg_cache_width_cntr_counter_out_14 (.Q (
         cache_width_cntr_counter_out_14), .QB (nx4692), .D (nx2389), .CLK (clk)
         , .R (nx6739)) ;
    nand02 ix1193 (.Y (nx1192), .A0 (nx4701), .A1 (nx5011)) ;
    aoi21 ix4702 (.Y (nx4701), .A0 (nx4703), .A1 (nx6685), .B0 (nx6603)) ;
    dffr ftc_cntrl_reg_reg_q_12 (.Q (ftc_cntrl_reg_out_12), .QB (nx4705), .D (
         nx2409), .CLK (nx6629), .R (nx6601)) ;
    or02 ix307 (.Y (nx306), .A0 (nx1427), .A1 (nx6603)) ;
    dffr reg_current_state_14 (.Q (\$dummy [51]), .QB (nx4711), .D (nx306), .CLK (
         nx6629), .R (reset)) ;
    mux21_ni ix1620 (.Y (nx1619), .A0 (cache_height_ended), .A1 (
             ftc_cntrl_reg_out_13), .S0 (nx6835)) ;
    dffr reg_current_state_15 (.Q (current_state_15), .QB (nx4725), .D (nx1108)
         , .CLK (nx6629), .R (reset)) ;
    oai22 ix1109 (.Y (nx1108), .A0 (nx4151), .A1 (nx4153), .B0 (nx7033), .B1 (
          nx4723)) ;
    dffr ftc_cntrl_reg_reg_q_13 (.Q (ftc_cntrl_reg_out_13), .QB (nx4723), .D (
         nx1619), .CLK (nx6629), .R (nx6601)) ;
    nand02 ix1139 (.Y (nx1138), .A0 (nx6977), .A1 (nx4751)) ;
    mux21 ix1890 (.Y (nx1889), .A0 (nx4735), .A1 (nx4731), .S0 (nx6835)) ;
    nand04 ix4736 (.Y (nx4735), .A0 (nx520), .A1 (nx534), .A2 (nx582), .A3 (
           nx702)) ;
    dffr window_width_cntr_counter_out_15 (.Q (\$dummy [52]), .QB (nx4743), .D (
         nx1779), .CLK (clk), .R (nx6723)) ;
    nand02 ix349 (.Y (nx348), .A0 (nx4747), .A1 (nx4751)) ;
    aoi22 ix4748 (.Y (nx4747), .A0 (nx6685), .A1 (ftc_cntrl_reg_out_13), .B0 (
          current_state_20), .B1 (ftc_cntrl_reg_out_12)) ;
    dffr reg_current_state_20 (.Q (current_state_20), .QB (nx4575), .D (nx1842)
         , .CLK (nx6631), .R (reset)) ;
    mux21_ni ix2230 (.Y (nx2229), .A0 (nx1124), .A1 (ftc_cntrl_reg_out_9), .S0 (
             nx6835)) ;
    oai21 ix1125 (.Y (nx1124), .A0 (nx4759), .A1 (nx4761), .B0 (nx4747)) ;
    dffr ftc_cntrl_reg_reg_q_9 (.Q (ftc_cntrl_reg_out_9), .QB (nx4759), .D (
         nx2229), .CLK (nx6631), .R (nx6601)) ;
    aoi21 ix4762 (.Y (nx4761), .A0 (nx6977), .A1 (nx1116), .B0 (nx6685)) ;
    dffr reg_current_state_16 (.Q (current_state_16), .QB (nx4765), .D (nx1138)
         , .CLK (nx6631), .R (reset)) ;
    dffr reg_window_width_cntr_counter_out_14 (.Q (
         window_width_cntr_counter_out_14), .QB (nx4770), .D (nx1769), .CLK (clk
         ), .R (nx6723)) ;
    nand02 ix4777 (.Y (nx4776), .A0 (window_width_cntr_counter_out_13), .A1 (
           nx1432)) ;
    dffr reg_window_width_cntr_counter_out_13 (.Q (
         window_width_cntr_counter_out_13), .QB (nx4781), .D (nx1759), .CLK (clk
         ), .R (nx6723)) ;
    oai21 ix4784 (.Y (nx4783), .A0 (nx1432), .A1 (
          window_width_cntr_counter_out_13), .B0 (nx4776)) ;
    dffr reg_window_width_cntr_counter_out_12 (.Q (
         window_width_cntr_counter_out_12), .QB (nx4787), .D (nx1749), .CLK (clk
         ), .R (nx6723)) ;
    nand02 ix4796 (.Y (nx4795), .A0 (window_width_cntr_counter_out_11), .A1 (
           nx1434)) ;
    dffr reg_window_width_cntr_counter_out_11 (.Q (
         window_width_cntr_counter_out_11), .QB (nx4801), .D (nx1739), .CLK (clk
         ), .R (nx6723)) ;
    oai21 ix4804 (.Y (nx4803), .A0 (nx1434), .A1 (
          window_width_cntr_counter_out_11), .B0 (nx4795)) ;
    dffr reg_window_width_cntr_counter_out_10 (.Q (
         window_width_cntr_counter_out_10), .QB (nx4807), .D (nx1729), .CLK (clk
         ), .R (nx6723)) ;
    nand02 ix4814 (.Y (nx4813), .A0 (window_width_cntr_counter_out_9), .A1 (
           nx1436)) ;
    dffr reg_window_width_cntr_counter_out_9 (.Q (
         window_width_cntr_counter_out_9), .QB (nx4819), .D (nx1719), .CLK (clk)
         , .R (nx6723)) ;
    oai21 ix4822 (.Y (nx4821), .A0 (nx1436), .A1 (
          window_width_cntr_counter_out_9), .B0 (nx4813)) ;
    dffr reg_window_width_cntr_counter_out_8 (.Q (
         window_width_cntr_counter_out_8), .QB (nx4825), .D (nx1709), .CLK (clk)
         , .R (nx6725)) ;
    nand02 ix4834 (.Y (nx4833), .A0 (window_width_cntr_counter_out_7), .A1 (
           nx1439)) ;
    dffr reg_window_width_cntr_counter_out_7 (.Q (
         window_width_cntr_counter_out_7), .QB (nx4839), .D (nx1699), .CLK (clk)
         , .R (nx6725)) ;
    oai21 ix4842 (.Y (nx4841), .A0 (nx1439), .A1 (
          window_width_cntr_counter_out_7), .B0 (nx4833)) ;
    dffr reg_window_width_cntr_counter_out_6 (.Q (
         window_width_cntr_counter_out_6), .QB (nx4845), .D (nx1689), .CLK (clk)
         , .R (nx6725)) ;
    dffr reg_wind_width_count_4 (.Q (wind_width_count_4), .QB (\$dummy [53]), .D (
         nx2599), .CLK (clk), .R (nx6727)) ;
    xnor2 ix1881 (.Y (nx1880), .A0 (wind_width_count_4), .A1 (nx4861)) ;
    nand04 ix4862 (.Y (nx4861), .A0 (wind_width_count_1), .A1 (nx6607), .A2 (
           wind_width_count_2), .A3 (wind_width_count_3)) ;
    dffr reg_wind_width_count_1 (.Q (wind_width_count_1), .QB (\$dummy [54]), .D (
         nx1649), .CLK (clk), .R (nx6725)) ;
    xor2 ix355 (.Y (nx354), .A0 (wind_width_count_1), .A1 (nx6607)) ;
    dffr reg_wind_width_count_0 (.Q (wind_width_count_0), .QB (\$dummy [55]), .D (
         nx1639), .CLK (clk), .R (nx6725)) ;
    oai21 ix1863 (.Y (nx1411), .A0 (nx4879), .A1 (nx4563), .B0 (nx4881)) ;
    dffr reg_current_state_21 (.Q (current_state_21), .QB (nx4879), .D (nx1411)
         , .CLK (nx6631), .R (reset)) ;
    nand03 ix4882 (.Y (nx4881), .A0 (nx1469), .A1 (nx4583), .A2 (nx4563)) ;
    dffr ftc_cntrl_reg_reg_q_11 (.Q (ftc_cntrl_reg_out_11), .QB (nx4731), .D (
         nx1889), .CLK (nx6631), .R (nx6601)) ;
    oai22 ix1879 (.Y (nx1429), .A0 (ftc_cntrl_reg_out_9), .A1 (nx6977), .B0 (
          nx4879), .B1 (ftc_cntrl_reg_out_11)) ;
    dffr reg_wind_width_count_2 (.Q (wind_width_count_2), .QB (\$dummy [56]), .D (
         nx1659), .CLK (clk), .R (nx6725)) ;
    xnor2 ix363 (.Y (nx362), .A0 (wind_width_count_2), .A1 (nx4895)) ;
    nand02 ix4896 (.Y (nx4895), .A0 (wind_width_count_1), .A1 (nx6609)) ;
    dffr reg_wind_width_count_3 (.Q (wind_width_count_3), .QB (\$dummy [57]), .D (
         nx1669), .CLK (clk), .R (nx6725)) ;
    xnor2 ix371 (.Y (nx370), .A0 (wind_width_count_3), .A1 (nx4903)) ;
    nand03 ix4904 (.Y (nx4903), .A0 (wind_width_count_1), .A1 (nx6609), .A2 (
           wind_width_count_2)) ;
    dffr reg_window_width_cntr_counter_out_5 (.Q (
         window_width_cntr_counter_out_5), .QB (nx4911), .D (nx1679), .CLK (clk)
         , .R (nx6727)) ;
    oai21 ix4914 (.Y (nx4913), .A0 (nx378), .A1 (window_width_cntr_counter_out_5
          ), .B0 (nx4853)) ;
    nor02ii ix379 (.Y (nx378), .A0 (nx4861), .A1 (wind_width_count_4)) ;
    xor2 ix575 (.Y (nx574), .A0 (nx572), .A1 (nx6609)) ;
    dffr img_width_reg_q_0 (.Q (img_width_out_0), .QB (nx4927), .D (nx1799), .CLK (
         clk), .R (reset)) ;
    mux21_ni ix1790 (.Y (nx1789), .A0 (new_width_out_0), .A1 (mem_data_in[0]), .S0 (
             current_state_6)) ;
    dffr new_width_reg_q_0 (.Q (new_width_out_0), .QB (\$dummy [58]), .D (nx1789
         ), .CLK (clk), .R (reset)) ;
    and04 ix703 (.Y (nx702), .A0 (nx4941), .A1 (nx4957), .A2 (nx4977), .A3 (
          nx4993)) ;
    xnor2 ix4942 (.Y (nx4941), .A0 (wind_width_count_1), .A1 (nx610)) ;
    dffr img_width_reg_q_1 (.Q (img_width_out_1), .QB (\$dummy [59]), .D (nx1819
         ), .CLK (clk), .R (reset)) ;
    ao22 ix1820 (.Y (nx1819), .A0 (nx6665), .A1 (new_width_out_1), .B0 (
         img_width_out_1), .B1 (nx4119)) ;
    dffr new_width_reg_q_1 (.Q (new_width_out_1), .QB (\$dummy [60]), .D (nx1809
         ), .CLK (clk), .R (reset)) ;
    mux21_ni ix1810 (.Y (nx1809), .A0 (new_width_out_1), .A1 (mem_data_in[1]), .S0 (
             current_state_6)) ;
    xnor2 ix4958 (.Y (nx4957), .A0 (wind_width_count_2), .A1 (nx644)) ;
    mux21 ix645 (.Y (nx644), .A0 (nx6641), .A1 (nx6839), .S0 (nx6977)) ;
    aoi21 ix4962 (.Y (nx4961), .A0 (img_width_out_2), .A1 (nx600), .B0 (nx4975)
          ) ;
    dffs_ni img_width_reg_q_2 (.Q (img_width_out_2), .QB (\$dummy [61]), .D (
            nx1839), .CLK (clk), .S (reset)) ;
    ao221 ix1840 (.Y (nx1839), .A0 (nx6665), .A1 (new_width_out_2), .B0 (
          img_width_out_2), .B1 (nx4119), .C0 (nx6695)) ;
    dffr new_width_reg_q_2 (.Q (new_width_out_2), .QB (\$dummy [62]), .D (nx1829
         ), .CLK (clk), .R (reset)) ;
    mux21_ni ix1830 (.Y (nx1829), .A0 (new_width_out_2), .A1 (mem_data_in[2]), .S0 (
             current_state_6)) ;
    nor03_2x ix4976 (.Y (nx4975), .A0 (img_width_out_0), .A1 (img_width_out_1), 
             .A2 (img_width_out_2)) ;
    xnor2 ix4978 (.Y (nx4977), .A0 (wind_width_count_3), .A1 (nx674)) ;
    xnor2 ix4982 (.Y (nx4981), .A0 (img_width_out_3), .A1 (nx4975)) ;
    dffs_ni img_width_reg_q_3 (.Q (img_width_out_3), .QB (\$dummy [63]), .D (
            nx1859), .CLK (clk), .S (reset)) ;
    ao22 ix1860 (.Y (nx1859), .A0 (nx6667), .A1 (new_width_out_3), .B0 (
         img_width_out_3), .B1 (nx4119)) ;
    dffr new_width_reg_q_3 (.Q (new_width_out_3), .QB (\$dummy [64]), .D (nx1849
         ), .CLK (clk), .R (reset)) ;
    mux21_ni ix1850 (.Y (nx1849), .A0 (new_width_out_3), .A1 (mem_data_in[3]), .S0 (
             current_state_6)) ;
    xnor2 ix4994 (.Y (nx4993), .A0 (wind_width_count_4), .A1 (nx692)) ;
    xnor2 ix4998 (.Y (nx4997), .A0 (img_width_out_4), .A1 (nx5009)) ;
    dffs_ni img_width_reg_q_4 (.Q (img_width_out_4), .QB (\$dummy [65]), .D (
            nx1879), .CLK (clk), .S (reset)) ;
    ao22 ix1880 (.Y (nx1879), .A0 (nx6667), .A1 (new_width_out_4), .B0 (
         img_width_out_4), .B1 (nx4119)) ;
    dffr new_width_reg_q_4 (.Q (new_width_out_4), .QB (\$dummy [66]), .D (nx1869
         ), .CLK (clk), .R (reset)) ;
    mux21_ni ix1870 (.Y (nx1869), .A0 (new_width_out_4), .A1 (mem_data_in[4]), .S0 (
             current_state_6)) ;
    nor04 ix5010 (.Y (nx5009), .A0 (img_width_out_0), .A1 (img_width_out_1), .A2 (
          img_width_out_2), .A3 (img_width_out_3)) ;
    nand02 ix5014 (.Y (nx5013), .A0 (cache_width_cntr_counter_out_13), .A1 (
           nx1449)) ;
    oai21 ix5020 (.Y (nx5019), .A0 (nx1449), .A1 (
          cache_width_cntr_counter_out_13), .B0 (nx5013)) ;
    dffr reg_cache_width_cntr_counter_out_12 (.Q (
         cache_width_cntr_counter_out_12), .QB (nx5023), .D (nx2369), .CLK (clk)
         , .R (nx6739)) ;
    nand02 ix5032 (.Y (nx5031), .A0 (cache_width_cntr_counter_out_11), .A1 (
           nx1451)) ;
    oai21 ix5038 (.Y (nx5037), .A0 (nx1451), .A1 (
          cache_width_cntr_counter_out_11), .B0 (nx5031)) ;
    dffr reg_cache_width_cntr_counter_out_10 (.Q (
         cache_width_cntr_counter_out_10), .QB (nx5041), .D (nx2349), .CLK (clk)
         , .R (nx6739)) ;
    nand02 ix5050 (.Y (nx5049), .A0 (cache_width_cntr_counter_out_9), .A1 (
           nx1454)) ;
    oai21 ix5056 (.Y (nx5055), .A0 (nx1454), .A1 (cache_width_cntr_counter_out_9
          ), .B0 (nx5049)) ;
    dffr reg_cache_width_cntr_counter_out_8 (.Q (cache_width_cntr_counter_out_8)
         , .QB (nx5059), .D (nx2329), .CLK (clk), .R (nx6739)) ;
    nand02 ix5068 (.Y (nx5067), .A0 (cache_width_cntr_counter_out_7), .A1 (
           nx1456)) ;
    oai21 ix5074 (.Y (nx5072), .A0 (nx1456), .A1 (cache_width_cntr_counter_out_7
          ), .B0 (nx5067)) ;
    dffr reg_cache_width_cntr_counter_out_6 (.Q (cache_width_cntr_counter_out_6)
         , .QB (nx5077), .D (nx2309), .CLK (clk), .R (nx6739)) ;
    dffr reg_cache_width_count_4 (.Q (cache_width_count_4), .QB (\$dummy [67]), 
         .D (nx2289), .CLK (clk), .R (nx6741)) ;
    xnor2 ix1223 (.Y (nx1222), .A0 (nx6611), .A1 (nx5089)) ;
    nand04 ix5090 (.Y (nx5089), .A0 (cache_width_count_1), .A1 (
           cache_width_count_0), .A2 (nx6615), .A3 (cache_width_count_3)) ;
    dffr reg_cache_width_count_1 (.Q (cache_width_count_1), .QB (\$dummy [68]), 
         .D (nx2259), .CLK (clk), .R (nx6739)) ;
    xor2 ix1199 (.Y (nx1198), .A0 (cache_width_count_1), .A1 (
         cache_width_count_0)) ;
    dffr reg_cache_width_count_0 (.Q (cache_width_count_0), .QB (\$dummy [69]), 
         .D (nx2249), .CLK (clk), .R (nx6739)) ;
    oai21 ix5100 (.Y (nx5099), .A0 (nx4), .A1 (nx1152), .B0 (
          ftc_cntrl_reg_out_10)) ;
    nor03_2x ix1153 (.Y (nx1152), .A0 (ftc_cntrl_reg_out_12), .A1 (nx7033), .A2 (
             ftc_cntrl_reg_out_13)) ;
    mux21 ix2240 (.Y (nx2239), .A0 (nx5107), .A1 (nx5115), .S0 (nx6835)) ;
    aoi221 ix5108 (.Y (nx5107), .A0 (current_state_20), .A1 (nx4705), .B0 (
           ftc_cntrl_reg_out_10), .B1 (nx1166), .C0 (nx1152)) ;
    oai21 ix1167 (.Y (nx1166), .A0 (nx7033), .A1 (cache_height_count_en), .B0 (
          nx320)) ;
    nor03_2x ix1159 (.Y (cache_height_count_en), .A0 (nx5113), .A1 (
             ftc_cntrl_reg_out_13), .A2 (nx4705)) ;
    dffr ftc_cntrl_reg_reg_q_10 (.Q (ftc_cntrl_reg_out_10), .QB (nx5115), .D (
         nx2239), .CLK (nx6631), .R (nx6603)) ;
    dffr reg_cache_width_count_2 (.Q (cache_width_count_2), .QB (\$dummy [70]), 
         .D (nx2269), .CLK (clk), .R (nx6741)) ;
    xnor2 ix1207 (.Y (nx1206), .A0 (nx6615), .A1 (nx5122)) ;
    nand02 ix5123 (.Y (nx5122), .A0 (cache_width_count_1), .A1 (
           cache_width_count_0)) ;
    dffr reg_cache_width_count_3 (.Q (cache_width_count_3), .QB (\$dummy [71]), 
         .D (nx2279), .CLK (clk), .R (nx6741)) ;
    xnor2 ix1215 (.Y (nx1214), .A0 (cache_width_count_3), .A1 (nx5128)) ;
    nand03 ix5129 (.Y (nx5128), .A0 (cache_width_count_1), .A1 (
           cache_width_count_0), .A2 (nx6617)) ;
    oai21 ix5135 (.Y (nx5134), .A0 (nx1228), .A1 (cache_width_cntr_counter_out_5
          ), .B0 (nx5083)) ;
    nor02ii ix1229 (.Y (nx1228), .A0 (nx5089), .A1 (nx6613)) ;
    dffr reg_cache_width_cntr_counter_out_5 (.Q (cache_width_cntr_counter_out_5)
         , .QB (nx5137), .D (nx2299), .CLK (clk), .R (nx6741)) ;
    dffr reg_cache_width_cntr_counter_out_7 (.Q (cache_width_cntr_counter_out_7)
         , .QB (nx5140), .D (nx2319), .CLK (clk), .R (nx6741)) ;
    dffr reg_cache_width_cntr_counter_out_9 (.Q (cache_width_cntr_counter_out_9)
         , .QB (nx5142), .D (nx2339), .CLK (clk), .R (nx6741)) ;
    dffr reg_cache_width_cntr_counter_out_11 (.Q (
         cache_width_cntr_counter_out_11), .QB (nx5144), .D (nx2359), .CLK (clk)
         , .R (nx6741)) ;
    dffr reg_cache_width_cntr_counter_out_13 (.Q (
         cache_width_cntr_counter_out_13), .QB (nx5146), .D (nx2379), .CLK (clk)
         , .R (nx6743)) ;
    dffr cache_width_cntr_counter_out_15 (.Q (\$dummy [72]), .QB (nx5148), .D (
         nx2399), .CLK (clk), .R (nx6743)) ;
    nor04 ix1425 (.Y (nx1424), .A0 (nx1404), .A1 (nx1406), .A2 (nx1414), .A3 (
          nx1416)) ;
    aoi21 ix5156 (.Y (nx5155), .A0 (img_width_out_1), .A1 (img_width_out_0), .B0 (
          nx5157)) ;
    xnor2 ix1407 (.Y (nx1406), .A0 (nx6617), .A1 (nx6839)) ;
    xnor2 ix1415 (.Y (nx1414), .A0 (cache_width_count_3), .A1 (nx4981)) ;
    xnor2 ix1417 (.Y (nx1416), .A0 (nx6613), .A1 (nx4997)) ;
    aoi43 ix5163 (.Y (nx5162), .A0 (nx4565), .A1 (nx6641), .A2 (current_state_20
          ), .A3 (nx4705), .B0 (nx4563), .B1 (ftc_cntrl_reg_out_11), .B2 (
          current_state_21)) ;
    aoi22 ix5165 (.Y (nx5164), .A0 (nx6685), .A1 (nx4723), .B0 (nx4879), .B1 (
          nx5113)) ;
    dffr ftc_cntrl_reg_reg_q_14 (.Q (ftc_cntrl_reg_out_14), .QB (nx4565), .D (
         nx1629), .CLK (nx6631), .R (nx6603)) ;
    oai221 ix15 (.Y (nx14), .A0 (nx4575), .A1 (ftc_cntrl_reg_out_12), .B0 (
           nx4879), .B1 (nx4563), .C0 (nx5168)) ;
    nand02 ix5169 (.Y (nx5168), .A0 (nx4879), .A1 (nx5011)) ;
    dffr reg_current_state_18 (.Q (current_state_18), .QB (\$dummy [73]), .D (
         nx1452), .CLK (nx6633), .R (reset)) ;
    ao22 ix2007 (.Y (mem_data_out[5]), .A0 (comp_unit_data2_in[5]), .A1 (nx6673)
         , .B0 (comp_unit_data1_in[5]), .B1 (nx6679)) ;
    ao22 ix2013 (.Y (mem_data_out[6]), .A0 (comp_unit_data2_in[6]), .A1 (nx6673)
         , .B0 (comp_unit_data1_in[6]), .B1 (nx6679)) ;
    ao22 ix2019 (.Y (mem_data_out[7]), .A0 (comp_unit_data2_in[7]), .A1 (nx6673)
         , .B0 (comp_unit_data1_in[7]), .B1 (nx6679)) ;
    ao22 ix2025 (.Y (mem_data_out[8]), .A0 (comp_unit_data2_in[8]), .A1 (nx6673)
         , .B0 (comp_unit_data1_in[8]), .B1 (nx6679)) ;
    ao22 ix2031 (.Y (mem_data_out[9]), .A0 (comp_unit_data2_in[9]), .A1 (nx6673)
         , .B0 (comp_unit_data1_in[9]), .B1 (nx6681)) ;
    ao22 ix2037 (.Y (mem_data_out[10]), .A0 (comp_unit_data2_in[10]), .A1 (
         nx6675), .B0 (comp_unit_data1_in[10]), .B1 (nx6681)) ;
    ao22 ix2043 (.Y (mem_data_out[11]), .A0 (comp_unit_data2_in[11]), .A1 (
         nx6675), .B0 (comp_unit_data1_in[11]), .B1 (nx6681)) ;
    ao22 ix2049 (.Y (mem_data_out[12]), .A0 (comp_unit_data2_in[12]), .A1 (
         nx6675), .B0 (comp_unit_data1_in[12]), .B1 (nx6681)) ;
    ao22 ix2055 (.Y (mem_data_out[13]), .A0 (comp_unit_data2_in[13]), .A1 (
         nx6675), .B0 (comp_unit_data1_in[13]), .B1 (nx6681)) ;
    ao22 ix2061 (.Y (mem_data_out[14]), .A0 (comp_unit_data2_in[14]), .A1 (
         nx6675), .B0 (comp_unit_data1_in[14]), .B1 (nx6681)) ;
    ao22 ix2067 (.Y (mem_data_out[15]), .A0 (comp_unit_data2_in[15]), .A1 (
         nx6675), .B0 (comp_unit_data1_in[15]), .B1 (nx6681)) ;
    nand02 ix1943 (.Y (nx1942), .A0 (nx5188), .A1 (nx7043)) ;
    nand03 ix5189 (.Y (nx5188), .A0 (nx1419), .A1 (nx4519), .A2 (nx4017)) ;
    nor02_2x ix1741 (.Y (nx1419), .A0 (nx1409), .A1 (nx4123)) ;
    dffr reg_current_state_27 (.Q (current_state_27), .QB (nx5197), .D (nx1942)
         , .CLK (nx6633), .R (reset)) ;
    dffr reg_class_cntr_counter_out_0 (.Q (class_cntr_counter_out_0), .QB (
         nx5194), .D (nx2609), .CLK (nx6633), .R (reset)) ;
    dffr reg_class_cntr_counter_out_1 (.Q (class_cntr_counter_out_1), .QB (
         nx5202), .D (nx2619), .CLK (nx6633), .R (reset)) ;
    oai21 ix5205 (.Y (nx5204), .A0 (class_cntr_counter_out_0), .A1 (
          class_cntr_counter_out_1), .B0 (nx5206)) ;
    dffr reg_class_cntr_counter_out_2 (.Q (class_cntr_counter_out_2), .QB (
         nx5208), .D (nx2629), .CLK (nx6633), .R (reset)) ;
    dffr reg_class_cntr_counter_out_3 (.Q (class_cntr_counter_out_3), .QB (
         nx5218), .D (nx2639), .CLK (nx6633), .R (reset)) ;
    dff reg_flt_bias1_reg_q_0 (.Q (flt_bias_out_0), .QB (\$dummy [74]), .D (
        nx2659), .CLK (clk)) ;
    mux21_ni ix2660 (.Y (nx2659), .A0 (flt_bias_out_0), .A1 (mem_data_in[0]), .S0 (
             nx7091)) ;
    oai21 ix2650 (.Y (nx2649), .A0 (nx7053), .A1 (nx152), .B0 (nx4635)) ;
    dffr channel_zero_reg_q_0 (.Q (\$dummy [75]), .QB (nx5243), .D (nx2649), .CLK (
         clk), .R (reset)) ;
    dff reg_flt_bias1_reg_q_1 (.Q (flt_bias_out_1), .QB (\$dummy [76]), .D (
        nx2679), .CLK (clk)) ;
    mux21_ni ix2680 (.Y (nx2679), .A0 (flt_bias_out_1), .A1 (mem_data_in[1]), .S0 (
             nx7091)) ;
    dff reg_flt_bias1_reg_q_2 (.Q (flt_bias_out_2), .QB (\$dummy [77]), .D (
        nx2699), .CLK (clk)) ;
    mux21_ni ix2700 (.Y (nx2699), .A0 (flt_bias_out_2), .A1 (mem_data_in[2]), .S0 (
             nx7091)) ;
    dff reg_flt_bias1_reg_q_3 (.Q (flt_bias_out_3), .QB (\$dummy [78]), .D (
        nx2719), .CLK (clk)) ;
    mux21_ni ix2720 (.Y (nx2719), .A0 (flt_bias_out_3), .A1 (mem_data_in[3]), .S0 (
             nx7091)) ;
    dff reg_flt_bias1_reg_q_4 (.Q (flt_bias_out_4), .QB (\$dummy [79]), .D (
        nx2739), .CLK (clk)) ;
    mux21_ni ix2740 (.Y (nx2739), .A0 (flt_bias_out_4), .A1 (mem_data_in[4]), .S0 (
             nx7091)) ;
    dff reg_flt_bias1_reg_q_5 (.Q (flt_bias_out_5), .QB (\$dummy [80]), .D (
        nx2759), .CLK (clk)) ;
    mux21_ni ix2760 (.Y (nx2759), .A0 (flt_bias_out_5), .A1 (mem_data_in[5]), .S0 (
             nx7091)) ;
    dff reg_flt_bias1_reg_q_6 (.Q (flt_bias_out_6), .QB (\$dummy [81]), .D (
        nx2779), .CLK (clk)) ;
    mux21_ni ix2780 (.Y (nx2779), .A0 (flt_bias_out_6), .A1 (mem_data_in[6]), .S0 (
             nx7093)) ;
    dff reg_flt_bias1_reg_q_7 (.Q (flt_bias_out_7), .QB (\$dummy [82]), .D (
        nx2799), .CLK (clk)) ;
    mux21_ni ix2800 (.Y (nx2799), .A0 (flt_bias_out_7), .A1 (mem_data_in[7]), .S0 (
             nx7093)) ;
    dff reg_flt_bias1_reg_q_8 (.Q (flt_bias_out_8), .QB (\$dummy [83]), .D (
        nx2819), .CLK (clk)) ;
    mux21_ni ix2820 (.Y (nx2819), .A0 (flt_bias_out_8), .A1 (mem_data_in[8]), .S0 (
             nx7093)) ;
    dff reg_flt_bias1_reg_q_9 (.Q (flt_bias_out_9), .QB (\$dummy [84]), .D (
        nx2839), .CLK (clk)) ;
    mux21_ni ix2840 (.Y (nx2839), .A0 (flt_bias_out_9), .A1 (mem_data_in[9]), .S0 (
             nx7093)) ;
    dff reg_flt_bias1_reg_q_10 (.Q (flt_bias_out_10), .QB (\$dummy [85]), .D (
        nx2859), .CLK (clk)) ;
    mux21_ni ix2860 (.Y (nx2859), .A0 (flt_bias_out_10), .A1 (mem_data_in[10]), 
             .S0 (nx7093)) ;
    dff reg_flt_bias1_reg_q_11 (.Q (flt_bias_out_11), .QB (\$dummy [86]), .D (
        nx2879), .CLK (clk)) ;
    mux21_ni ix2880 (.Y (nx2879), .A0 (flt_bias_out_11), .A1 (mem_data_in[11]), 
             .S0 (nx7093)) ;
    dff reg_flt_bias1_reg_q_12 (.Q (flt_bias_out_12), .QB (\$dummy [87]), .D (
        nx2899), .CLK (clk)) ;
    mux21_ni ix2900 (.Y (nx2899), .A0 (flt_bias_out_12), .A1 (mem_data_in[12]), 
             .S0 (nx6993)) ;
    dff reg_flt_bias1_reg_q_13 (.Q (flt_bias_out_13), .QB (\$dummy [88]), .D (
        nx2919), .CLK (clk)) ;
    mux21_ni ix2920 (.Y (nx2919), .A0 (flt_bias_out_13), .A1 (mem_data_in[13]), 
             .S0 (nx6993)) ;
    dff reg_flt_bias1_reg_q_14 (.Q (flt_bias_out_14), .QB (\$dummy [89]), .D (
        nx2939), .CLK (clk)) ;
    mux21_ni ix2940 (.Y (nx2939), .A0 (flt_bias_out_14), .A1 (mem_data_in[14]), 
             .S0 (nx6993)) ;
    dff reg_flt_bias1_reg_q_15 (.Q (flt_bias_out_15), .QB (\$dummy [90]), .D (
        nx2959), .CLK (clk)) ;
    mux21_ni ix2960 (.Y (nx2959), .A0 (flt_bias_out_15), .A1 (mem_data_in[15]), 
             .S0 (nx6993)) ;
    nor03_2x ix5083 (.Y (max_height_3), .A0 (nx4981), .A1 (nx6603), .A2 (nx6687)
             ) ;
    nor03_2x ix5087 (.Y (max_height_4), .A0 (nx4997), .A1 (nx6603), .A2 (nx6687)
             ) ;
    or02 ix4791 (.Y (cache_rst_actual), .A0 (nx6605), .A1 (reset)) ;
    mux21 ix2980 (.Y (nx2979), .A0 (nx5330), .A1 (nx5334), .S0 (nx6837)) ;
    aoi32 ix5331 (.Y (nx5330), .A0 (nx1428), .A1 (cache_height_ended), .A2 (
          current_state_20), .B0 (ftc_cntrl_reg_out_15), .B1 (nx2522)) ;
    dffr ftc_cntrl_reg_reg_q_15 (.Q (ftc_cntrl_reg_out_15), .QB (nx5334), .D (
         nx2979), .CLK (nx6635), .R (nx6605)) ;
    nand02 ix5073 (.Y (max_height_0), .A0 (nx5379), .A1 (img_width_out_0)) ;
    nand02 ix5079 (.Y (max_height_2), .A0 (nx5379), .A1 (nx6839)) ;
    oai21 ix2109 (.Y (comp_unit_data1_out[0]), .A0 (nx6855), .A1 (nx5383), .B0 (
          nx5386)) ;
    dffr bias1_reg_reg_q_0 (.Q (\$dummy [91]), .QB (nx5383), .D (nx2669), .CLK (
         clk), .R (reset)) ;
    nand02 ix5387 (.Y (nx5386), .A0 (nx2096), .A1 (nx6763)) ;
    oai21 ix2135 (.Y (comp_unit_data1_out[1]), .A0 (nx6855), .A1 (nx5390), .B0 (
          nx5393)) ;
    dffr bias1_reg_reg_q_1 (.Q (\$dummy [92]), .QB (nx5390), .D (nx2689), .CLK (
         clk), .R (reset)) ;
    nand02 ix5394 (.Y (nx5393), .A0 (nx2124), .A1 (nx6763)) ;
    oai21 ix2161 (.Y (comp_unit_data1_out[2]), .A0 (nx6855), .A1 (nx5396), .B0 (
          nx5399)) ;
    dffr bias1_reg_reg_q_2 (.Q (\$dummy [93]), .QB (nx5396), .D (nx2709), .CLK (
         clk), .R (reset)) ;
    nand02 ix5400 (.Y (nx5399), .A0 (nx2150), .A1 (nx6763)) ;
    oai21 ix2187 (.Y (comp_unit_data1_out[3]), .A0 (nx6855), .A1 (nx5402), .B0 (
          nx5405)) ;
    dffr bias1_reg_reg_q_3 (.Q (\$dummy [94]), .QB (nx5402), .D (nx2729), .CLK (
         clk), .R (reset)) ;
    nand02 ix5406 (.Y (nx5405), .A0 (nx2176), .A1 (nx6763)) ;
    oai21 ix2213 (.Y (comp_unit_data1_out[4]), .A0 (nx6857), .A1 (nx5408), .B0 (
          nx5411)) ;
    dffr bias1_reg_reg_q_4 (.Q (\$dummy [95]), .QB (nx5408), .D (nx2749), .CLK (
         clk), .R (reset)) ;
    nand02 ix5412 (.Y (nx5411), .A0 (nx2202), .A1 (nx6763)) ;
    oai21 ix2239 (.Y (comp_unit_data1_out[5]), .A0 (nx6857), .A1 (nx5414), .B0 (
          nx5417)) ;
    dffr bias1_reg_reg_q_5 (.Q (\$dummy [96]), .QB (nx5414), .D (nx2769), .CLK (
         clk), .R (reset)) ;
    nand02 ix5418 (.Y (nx5417), .A0 (nx2228), .A1 (nx6763)) ;
    oai21 ix2265 (.Y (comp_unit_data1_out[6]), .A0 (nx6857), .A1 (nx5420), .B0 (
          nx5423)) ;
    dffr bias1_reg_reg_q_6 (.Q (\$dummy [97]), .QB (nx5420), .D (nx2789), .CLK (
         clk), .R (reset)) ;
    nand02 ix5424 (.Y (nx5423), .A0 (nx2254), .A1 (nx6763)) ;
    oai21 ix2291 (.Y (comp_unit_data1_out[7]), .A0 (nx6857), .A1 (nx5426), .B0 (
          nx5429)) ;
    dffr bias1_reg_reg_q_7 (.Q (\$dummy [98]), .QB (nx5426), .D (nx2809), .CLK (
         clk), .R (reset)) ;
    nand02 ix5430 (.Y (nx5429), .A0 (nx2280), .A1 (nx6765)) ;
    oai21 ix2317 (.Y (comp_unit_data1_out[8]), .A0 (nx6857), .A1 (nx5432), .B0 (
          nx5435)) ;
    dffr bias1_reg_reg_q_8 (.Q (\$dummy [99]), .QB (nx5432), .D (nx2829), .CLK (
         clk), .R (reset)) ;
    nand02 ix5436 (.Y (nx5435), .A0 (nx2306), .A1 (nx6765)) ;
    oai21 ix2343 (.Y (comp_unit_data1_out[9]), .A0 (nx6857), .A1 (nx5438), .B0 (
          nx5441)) ;
    dffr bias1_reg_reg_q_9 (.Q (\$dummy [100]), .QB (nx5438), .D (nx2849), .CLK (
         clk), .R (reset)) ;
    nand02 ix5442 (.Y (nx5441), .A0 (nx2332), .A1 (nx6765)) ;
    oai21 ix2369 (.Y (comp_unit_data1_out[10]), .A0 (nx6857), .A1 (nx5444), .B0 (
          nx5447)) ;
    dffr bias1_reg_reg_q_10 (.Q (\$dummy [101]), .QB (nx5444), .D (nx2869), .CLK (
         clk), .R (reset)) ;
    nand02 ix5448 (.Y (nx5447), .A0 (nx2358), .A1 (nx6765)) ;
    oai21 ix2395 (.Y (comp_unit_data1_out[11]), .A0 (nx6859), .A1 (nx5450), .B0 (
          nx5453)) ;
    dffr bias1_reg_reg_q_11 (.Q (\$dummy [102]), .QB (nx5450), .D (nx2889), .CLK (
         clk), .R (reset)) ;
    nand02 ix5454 (.Y (nx5453), .A0 (nx2384), .A1 (nx6765)) ;
    oai21 ix2421 (.Y (comp_unit_data1_out[12]), .A0 (nx6859), .A1 (nx5456), .B0 (
          nx5459)) ;
    dffr bias1_reg_reg_q_12 (.Q (\$dummy [103]), .QB (nx5456), .D (nx2909), .CLK (
         clk), .R (reset)) ;
    nand02 ix5460 (.Y (nx5459), .A0 (nx2410), .A1 (nx6765)) ;
    oai21 ix2447 (.Y (comp_unit_data1_out[13]), .A0 (nx6859), .A1 (nx5462), .B0 (
          nx5465)) ;
    dffr bias1_reg_reg_q_13 (.Q (\$dummy [104]), .QB (nx5462), .D (nx2929), .CLK (
         clk), .R (reset)) ;
    nand02 ix5466 (.Y (nx5465), .A0 (nx2436), .A1 (nx6765)) ;
    oai21 ix2473 (.Y (comp_unit_data1_out[14]), .A0 (nx6859), .A1 (nx5468), .B0 (
          nx5471)) ;
    dffr bias1_reg_reg_q_14 (.Q (\$dummy [105]), .QB (nx5468), .D (nx2949), .CLK (
         clk), .R (reset)) ;
    nand02 ix5472 (.Y (nx5471), .A0 (nx2462), .A1 (nx6767)) ;
    oai21 ix2499 (.Y (comp_unit_data1_out[15]), .A0 (nx6859), .A1 (nx5474), .B0 (
          nx5477)) ;
    dffr bias1_reg_reg_q_15 (.Q (\$dummy [106]), .QB (nx5474), .D (nx2969), .CLK (
         clk), .R (reset)) ;
    nand02 ix5478 (.Y (nx5477), .A0 (nx2488), .A1 (nx6767)) ;
    oai21 ix2073 (.Y (comp_unit_ready), .A0 (nx7023), .A1 (nx6705), .B0 (nx5480)
          ) ;
    aoi21 ix5481 (.Y (nx5480), .A0 (nx6749), .A1 (nx7063), .B0 (nx6985)) ;
    nand03 ix5483 (.Y (nx5482), .A0 (flt_size_out_0), .A1 (nx4143), .A2 (
           flt_size_out_1)) ;
    aoi21 ix4813 (.Y (mem_read_out), .A0 (nx5587), .A1 (nx5593), .B0 (reset)) ;
    nor04 ix5594 (.Y (nx5593), .A0 (nx6769), .A1 (nx6663), .A2 (nx2706), .A3 (
          nx6993)) ;
    nand02 ix2707 (.Y (nx2706), .A0 (nx5596), .A1 (nx5598)) ;
    nor04 ix5597 (.Y (nx5596), .A0 (current_state_2), .A1 (current_state_3), .A2 (
          nx6691), .A3 (current_state_5)) ;
    aoi21 ix4797 (.Y (mem_write_out), .A0 (nx6833), .A1 (nx6899), .B0 (reset)) ;
    dffr reg_current_state_28 (.Q (current_state_28), .QB (\$dummy [107]), .D (
         nx1950), .CLK (nx6635), .R (reset)) ;
    nand04 ix2739 (.Y (mem_addr_out[0]), .A0 (nx5605), .A1 (nx6899), .A2 (nx5629
           ), .A3 (nx5664)) ;
    aoi22 ix5606 (.Y (nx5605), .A0 (nx5607), .A1 (nx6651), .B0 (addr1_data_0), .B1 (
          nx6815)) ;
    oai21 ix5608 (.Y (nx5607), .A0 (class_cntr_counter_out_0), .A1 (nx6775), .B0 (
          nx5621)) ;
    oai21 ix2990 (.Y (nx2989), .A0 (nx7357), .A1 (nx6781), .B0 (nx5616)) ;
    dffr reg_write_base_reg_q_0 (.Q (\$dummy [108]), .QB (nx5611), .D (nx2989), 
         .CLK (nx6635), .R (reset)) ;
    nand02 ix2581 (.Y (nx2580), .A0 (nx5614), .A1 (nx7009)) ;
    aoi21 ix5615 (.Y (nx5614), .A0 (nx7021), .A1 (nx1421), .B0 (current_state_25
          )) ;
    nand03 ix5617 (.Y (nx5616), .A0 (nx2582), .A1 (nx5619), .A2 (nx6781)) ;
    nand02 ix2583 (.Y (nx2582), .A0 (nx7357), .A1 (nx4423)) ;
    dffr reg_addr1_data_0 (.Q (addr1_data_0), .QB (\$dummy [109]), .D (nx3039), 
         .CLK (clk), .R (reset)) ;
    aoi43 ix5630 (.Y (nx5629), .A0 (nx2620), .A1 (nx5636), .A2 (nx6985), .A3 (
          nx7053), .B0 (nx2680), .B1 (nx5662), .B2 (nx6769)) ;
    nand02 ix2621 (.Y (nx2620), .A0 (nx7357), .A1 (nx5632)) ;
    dffr reg_bias_offset_reg_q_0 (.Q (bias_offset_data_out_0), .QB (nx5632), .D (
         nx2999), .CLK (clk), .R (reset)) ;
    or02 ix2681 (.Y (nx2680), .A0 (img_addr_offset_0), .A1 (img_base_addr_0)) ;
    dffr reg_img_addr_offset_0 (.Q (img_addr_offset_0), .QB (\$dummy [110]), .D (
         nx3029), .CLK (clk), .R (nx6807)) ;
    dffs_ni img_base_addr_inst_reg_q_0 (.Q (img_base_addr_0), .QB (\$dummy [111]
            ), .D (nx3019), .CLK (clk), .S (reset)) ;
    dffr reg_write_base_prev_reg_q_0 (.Q (write_base_prev_data_out_0), .QB (
         nx5647), .D (nx3009), .CLK (clk), .R (reset)) ;
    nand04 ix5652 (.Y (nx5651), .A0 (nx5653), .A1 (nx2640), .A2 (nx5657), .A3 (
           nx5659)) ;
    nand02 ix5663 (.Y (nx5662), .A0 (img_base_addr_0), .A1 (img_addr_offset_0)
           ) ;
    oai221 ix5665 (.Y (nx5664), .A0 (nx6787), .A1 (nx6981), .B0 (
           write_offset_data_out_0), .B1 (nx6775), .C0 (nx5667)) ;
    nand03 ix2843 (.Y (mem_addr_out[1]), .A0 (nx5670), .A1 (nx6899), .A2 (nx5709
           )) ;
    aoi22 ix5671 (.Y (nx5670), .A0 (nx2834), .A1 (nx6769), .B0 (nx2796), .B1 (
          nx6801)) ;
    xor2 ix2835 (.Y (nx2834), .A0 (nx5662), .A1 (nx5673)) ;
    dffs_ni img_base_addr_inst_reg_q_1 (.Q (img_base_addr_1), .QB (nx5677), .D (
            nx3089), .CLK (clk), .S (reset)) ;
    aoi21 ix5680 (.Y (nx5679), .A0 (write_base_prev_data_out_1), .A1 (
          write_base_prev_data_out_0), .B0 (nx5692)) ;
    dffr reg_write_base_prev_reg_q_1 (.Q (write_base_prev_data_out_1), .QB (
         \$dummy [112]), .D (nx3079), .CLK (clk), .R (reset)) ;
    dffr reg_write_base_reg_q_1 (.Q (write_base_data_out_1), .QB (nx5685), .D (
         nx3049), .CLK (nx6635), .R (reset)) ;
    xnor2 ix5688 (.Y (nx5687), .A0 (nx5619), .A1 (nx5689)) ;
    oai21 ix5697 (.Y (nx5696), .A0 (img_addr_offset_0), .A1 (img_addr_offset_1)
          , .B0 (nx5698)) ;
    nand02 ix5699 (.Y (nx5698), .A0 (img_addr_offset_1), .A1 (img_addr_offset_0)
           ) ;
    dffr reg_img_addr_offset_1 (.Q (img_addr_offset_1), .QB (nx5700), .D (nx3099
         ), .CLK (clk), .R (nx6807)) ;
    xor2 ix2797 (.Y (nx2796), .A0 (nx5636), .A1 (nx5703)) ;
    dffr reg_bias_offset_reg_q_1 (.Q (bias_offset_data_out_1), .QB (nx5707), .D (
         nx3069), .CLK (clk), .R (reset)) ;
    aoi222 ix5710 (.Y (nx5709), .A0 (nx6651), .A1 (nx2766), .B0 (addr1_data_1), 
           .B1 (nx6815), .C0 (nx2752), .C1 (nx6795)) ;
    xnor2 ix2767 (.Y (nx2766), .A0 (nx5607), .A1 (nx5712)) ;
    xnor2 ix5713 (.Y (nx5712), .A0 (nx5621), .A1 (nx5714)) ;
    oai21 ix5719 (.Y (nx5718), .A0 (addr1_data_0), .A1 (addr1_data_1), .B0 (
          nx5720)) ;
    nand02 ix5721 (.Y (nx5720), .A0 (addr1_data_1), .A1 (addr1_data_0)) ;
    dffr reg_addr1_data_1 (.Q (addr1_data_1), .QB (nx5722), .D (nx3059), .CLK (
         clk), .R (reset)) ;
    xor2 ix2753 (.Y (nx2752), .A0 (nx5667), .A1 (nx5725)) ;
    nand03 ix2987 (.Y (mem_addr_out[2]), .A0 (nx5731), .A1 (nx6899), .A2 (nx5773
           )) ;
    aoi22 ix5732 (.Y (nx5731), .A0 (nx2978), .A1 (nx6769), .B0 (nx2932), .B1 (
          nx6801)) ;
    xor2 ix2979 (.Y (nx2978), .A0 (nx5734), .A1 (nx5737)) ;
    aoi32 ix5735 (.Y (nx5734), .A0 (img_base_addr_0), .A1 (img_addr_offset_0), .A2 (
          nx2832), .B0 (img_addr_offset_1), .B1 (img_base_addr_1)) ;
    dffs_ni img_base_addr_inst_reg_q_2 (.Q (img_base_addr_2), .QB (nx5758), .D (
            nx3149), .CLK (clk), .S (reset)) ;
    oai21 ix2957 (.Y (nx2956), .A0 (nx5742), .A1 (nx5692), .B0 (nx2950)) ;
    dffr reg_write_base_reg_q_2 (.Q (write_base_data_out_2), .QB (nx5747), .D (
         nx3109), .CLK (nx6635), .R (reset)) ;
    xnor2 ix5750 (.Y (nx5749), .A0 (nx5751), .A1 (nx5754)) ;
    dffr reg_write_base_prev_reg_q_2 (.Q (write_base_prev_data_out_2), .QB (
         nx5742), .D (nx3139), .CLK (clk), .R (reset)) ;
    dffr reg_img_addr_offset_2 (.Q (img_addr_offset_2), .QB (nx5762), .D (nx3159
         ), .CLK (clk), .R (nx6807)) ;
    xor2 ix2933 (.Y (nx2932), .A0 (nx5764), .A1 (nx5767)) ;
    aoi32 ix5765 (.Y (nx5764), .A0 (bias_offset_data_out_0), .A1 (nx6775), .A2 (
          nx2794), .B0 (write_base_data_out_1), .B1 (bias_offset_data_out_1)) ;
    dffr reg_bias_offset_reg_q_2 (.Q (bias_offset_data_out_2), .QB (nx5771), .D (
         nx3129), .CLK (clk), .R (reset)) ;
    aoi222 ix5774 (.Y (nx5773), .A0 (nx2872), .A1 (nx6795), .B0 (nx6651), .B1 (
           nx2894), .C0 (addr1_data_2), .C1 (nx6815)) ;
    xnor2 ix2873 (.Y (nx2872), .A0 (nx2850), .A1 (nx5777)) ;
    xnor2 ix2895 (.Y (nx2894), .A0 (nx2760), .A1 (nx2886)) ;
    nand02 ix2761 (.Y (nx2760), .A0 (nx5712), .A1 (nx5607)) ;
    xnor2 ix2887 (.Y (nx2886), .A0 (nx2882), .A1 (nx5783)) ;
    oai22 ix2883 (.Y (nx2882), .A0 (nx5621), .A1 (nx5714), .B0 (nx5202), .B1 (
          nx7359)) ;
    dffr reg_addr1_data_2 (.Q (addr1_data_2), .QB (\$dummy [113]), .D (nx3119), 
         .CLK (clk), .R (reset)) ;
    xnor2 ix2905 (.Y (nx2904), .A0 (addr1_data_2), .A1 (nx5720)) ;
    nand03 ix3131 (.Y (mem_addr_out[3]), .A0 (nx5790), .A1 (nx6899), .A2 (nx5826
           )) ;
    aoi22 ix5791 (.Y (nx5790), .A0 (nx3122), .A1 (nx6769), .B0 (nx3076), .B1 (
          nx6801)) ;
    xnor2 ix3123 (.Y (nx3122), .A0 (nx3086), .A1 (nx5794)) ;
    oai22 ix3087 (.Y (nx3086), .A0 (nx5734), .A1 (nx5737), .B0 (nx5762), .B1 (
          nx5758)) ;
    xnor2 ix5795 (.Y (nx5794), .A0 (img_base_addr_3), .A1 (img_addr_offset_3)) ;
    dffr img_base_addr_inst_reg_q_3 (.Q (img_base_addr_3), .QB (\$dummy [114]), 
         .D (nx3209), .CLK (clk), .R (reset)) ;
    xor2 ix3101 (.Y (nx3100), .A0 (write_base_prev_data_out_3), .A1 (nx5809)) ;
    dffr reg_write_base_prev_reg_q_3 (.Q (write_base_prev_data_out_3), .QB (
         \$dummy [115]), .D (nx3199), .CLK (clk), .R (reset)) ;
    dffs_ni reg_write_base_reg_q_3 (.Q (write_base_data_out_3), .QB (nx5807), .D (
            nx3169), .CLK (nx6635), .S (reset)) ;
    xnor2 ix3007 (.Y (nx3006), .A0 (nx3002), .A1 (nx5805)) ;
    nor03_2x ix5810 (.Y (nx5809), .A0 (write_base_prev_data_out_0), .A1 (
             write_base_prev_data_out_1), .A2 (write_base_prev_data_out_2)) ;
    dffr reg_img_addr_offset_3 (.Q (img_addr_offset_3), .QB (\$dummy [116]), .D (
         nx3219), .CLK (clk), .R (nx6807)) ;
    xnor2 ix3115 (.Y (nx3114), .A0 (img_addr_offset_3), .A1 (nx5815)) ;
    nand03 ix5816 (.Y (nx5815), .A0 (img_addr_offset_2), .A1 (img_addr_offset_1)
           , .A2 (img_addr_offset_0)) ;
    xnor2 ix3077 (.Y (nx3076), .A0 (nx3066), .A1 (nx5820)) ;
    oai22 ix3067 (.Y (nx3066), .A0 (nx5764), .A1 (nx5767), .B0 (nx7361), .B1 (
          nx5771)) ;
    dffr reg_bias_offset_reg_q_3 (.Q (bias_offset_data_out_3), .QB (
         \$dummy [117]), .D (nx3189), .CLK (clk), .R (reset)) ;
    aoi322 ix5827 (.Y (nx5826), .A0 (nx3032), .A1 (nx5838), .A2 (nx6651), .B0 (
           addr1_data_3), .B1 (nx6815), .C0 (nx3016), .C1 (nx6795)) ;
    nand02 ix3033 (.Y (nx3032), .A0 (nx5829), .A1 (nx5836)) ;
    xnor2 ix5830 (.Y (nx5829), .A0 (nx5831), .A1 (nx5834)) ;
    aoi22 ix5832 (.Y (nx5831), .A0 (class_cntr_counter_out_2), .A1 (
          write_base_data_out_2), .B0 (nx2882), .B1 (nx2884)) ;
    nor02_2x ix5837 (.Y (nx5836), .A0 (nx2886), .A1 (nx2760)) ;
    dffr reg_addr1_data_3 (.Q (addr1_data_3), .QB (\$dummy [118]), .D (nx3179), 
         .CLK (clk), .R (reset)) ;
    xnor2 ix3049 (.Y (nx3048), .A0 (addr1_data_3), .A1 (nx5843)) ;
    nand03 ix5844 (.Y (nx5843), .A0 (addr1_data_2), .A1 (addr1_data_1), .A2 (
           addr1_data_0)) ;
    xor2 ix3017 (.Y (nx3016), .A0 (nx5847), .A1 (nx5850)) ;
    nand03 ix3279 (.Y (mem_addr_out[4]), .A0 (nx5853), .A1 (nx6899), .A2 (nx5901
           )) ;
    aoi22 ix5854 (.Y (nx5853), .A0 (nx3270), .A1 (nx6769), .B0 (nx3224), .B1 (
          nx6801)) ;
    xor2 ix3271 (.Y (nx3270), .A0 (nx5856), .A1 (nx5859)) ;
    aoi22 ix5857 (.Y (nx5856), .A0 (img_addr_offset_3), .A1 (img_base_addr_3), .B0 (
          nx3086), .B1 (nx3120)) ;
    dffs_ni img_base_addr_inst_reg_q_4 (.Q (img_base_addr_4), .QB (nx5882), .D (
            nx3269), .CLK (clk), .S (reset)) ;
    oai21 ix3249 (.Y (nx3248), .A0 (nx5864), .A1 (nx5879), .B0 (nx3242)) ;
    dffr reg_write_base_reg_q_4 (.Q (write_base_data_out_4), .QB (nx5869), .D (
         nx3229), .CLK (nx6635), .R (reset)) ;
    xnor2 ix5872 (.Y (nx5871), .A0 (nx5873), .A1 (nx5876)) ;
    aoi22 ix5874 (.Y (nx5873), .A0 (write_base_data_out_3), .A1 (
          new_size_squared_out_3), .B0 (nx7323), .B1 (nx3004)) ;
    dffr reg_write_base_prev_reg_q_4 (.Q (\$dummy [119]), .QB (nx5864), .D (
         nx3259), .CLK (clk), .R (reset)) ;
    nor04 ix5880 (.Y (nx5879), .A0 (write_base_prev_data_out_0), .A1 (
          write_base_prev_data_out_1), .A2 (write_base_prev_data_out_2), .A3 (
          write_base_prev_data_out_3)) ;
    nand02 ix3243 (.Y (nx3242), .A0 (nx5879), .A1 (nx5864)) ;
    aoi21 ix3263 (.Y (nx3262), .A0 (nx5886), .A1 (nx5888), .B0 (nx3256)) ;
    nand04 ix5887 (.Y (nx5886), .A0 (img_addr_offset_3), .A1 (img_addr_offset_2)
           , .A2 (img_addr_offset_1), .A3 (img_addr_offset_0)) ;
    dffr reg_img_addr_offset_4 (.Q (img_addr_offset_4), .QB (nx5888), .D (nx3279
         ), .CLK (clk), .R (nx6807)) ;
    xor2 ix3225 (.Y (nx3224), .A0 (nx5892), .A1 (nx5895)) ;
    aoi22 ix5893 (.Y (nx5892), .A0 (write_base_data_out_3), .A1 (
          bias_offset_data_out_3), .B0 (nx3066), .B1 (nx3074)) ;
    dffr reg_bias_offset_reg_q_4 (.Q (bias_offset_data_out_4), .QB (nx5900), .D (
         nx3249), .CLK (clk), .R (reset)) ;
    aoi21 ix829 (.Y (nx828), .A0 (nx4265), .A1 (nx4257), .B0 (nx822)) ;
    aoi222 ix5902 (.Y (nx5901), .A0 (addr1_data_4), .A1 (nx6815), .B0 (nx3160), 
           .B1 (nx6795), .C0 (nx6651), .C1 (nx3186)) ;
    aoi21 ix3197 (.Y (nx3196), .A0 (nx5906), .A1 (nx5908), .B0 (nx3190)) ;
    nand04 ix5907 (.Y (nx5906), .A0 (addr1_data_3), .A1 (addr1_data_2), .A2 (
           addr1_data_1), .A3 (addr1_data_0)) ;
    dffr reg_addr1_data_4 (.Q (addr1_data_4), .QB (nx5908), .D (nx3239), .CLK (
         clk), .R (reset)) ;
    xnor2 ix3161 (.Y (nx3160), .A0 (nx3138), .A1 (nx5913)) ;
    oai22 ix3139 (.Y (nx3138), .A0 (nx7336), .A1 (nx5850), .B0 (nx4271), .B1 (
          nx5807)) ;
    xor2 ix3187 (.Y (nx3186), .A0 (nx3034), .A1 (nx5917)) ;
    nor02_2x ix3035 (.Y (nx3034), .A0 (nx5836), .A1 (nx5829)) ;
    oai22 ix3171 (.Y (nx3170), .A0 (nx5831), .A1 (nx5834), .B0 (nx5218), .B1 (
          nx5807)) ;
    nand03 ix3419 (.Y (mem_addr_out[5]), .A0 (nx5921), .A1 (nx6899), .A2 (nx5957
           )) ;
    aoi22 ix5922 (.Y (nx5921), .A0 (nx3410), .A1 (nx6771), .B0 (nx3364), .B1 (
          nx6801)) ;
    xnor2 ix3411 (.Y (nx3410), .A0 (nx3374), .A1 (nx5925)) ;
    oai22 ix3375 (.Y (nx3374), .A0 (nx5856), .A1 (nx5859), .B0 (nx5888), .B1 (
          nx5882)) ;
    dffr img_base_addr_inst_reg_q_5 (.Q (img_base_addr_5), .QB (\$dummy [120]), 
         .D (nx3329), .CLK (clk), .R (reset)) ;
    xnor2 ix3389 (.Y (nx3388), .A0 (write_base_prev_data_out_5), .A1 (nx3242)) ;
    dffr reg_write_base_prev_reg_q_5 (.Q (write_base_prev_data_out_5), .QB (
         \$dummy [121]), .D (nx3319), .CLK (clk), .R (reset)) ;
    dffs_ni reg_write_base_reg_q_5 (.Q (write_base_data_out_5), .QB (nx5938), .D (
            nx3289), .CLK (nx6637), .S (reset)) ;
    xnor2 ix3299 (.Y (nx3298), .A0 (nx3294), .A1 (nx5936)) ;
    oai22 ix3295 (.Y (nx3294), .A0 (nx5873), .A1 (nx5876), .B0 (nx5869), .B1 (
          nx4391)) ;
    oai21 ix5944 (.Y (nx5943), .A0 (nx3256), .A1 (img_addr_offset_5), .B0 (
          nx5945)) ;
    nand02 ix5946 (.Y (nx5945), .A0 (img_addr_offset_5), .A1 (nx3256)) ;
    dffr reg_img_addr_offset_5 (.Q (img_addr_offset_5), .QB (nx5947), .D (nx3339
         ), .CLK (clk), .R (nx6807)) ;
    xnor2 ix3365 (.Y (nx3364), .A0 (nx3354), .A1 (nx5951)) ;
    oai22 ix3355 (.Y (nx3354), .A0 (nx5892), .A1 (nx5895), .B0 (nx5869), .B1 (
          nx5900)) ;
    dffr reg_bias_offset_reg_q_5 (.Q (bias_offset_data_out_5), .QB (nx5955), .D (
         nx3309), .CLK (clk), .R (reset)) ;
    aoi222 ix5958 (.Y (nx5957), .A0 (addr1_data_5), .A1 (nx6815), .B0 (nx3308), 
           .B1 (nx6795), .C0 (nx6651), .C1 (nx3326)) ;
    oai21 ix5962 (.Y (nx5961), .A0 (nx3190), .A1 (addr1_data_5), .B0 (nx5963)) ;
    nand02 ix5964 (.Y (nx5963), .A0 (addr1_data_5), .A1 (nx3190)) ;
    dffr reg_addr1_data_5 (.Q (addr1_data_5), .QB (nx5965), .D (nx3299), .CLK (
         clk), .R (reset)) ;
    xor2 ix3309 (.Y (nx3308), .A0 (nx5968), .A1 (nx5971)) ;
    aoi22 ix5969 (.Y (nx5968), .A0 (write_offset_data_out_4), .A1 (
          write_base_data_out_4), .B0 (nx3138), .B1 (nx3158)) ;
    xor2 ix3327 (.Y (nx3326), .A0 (nx5974), .A1 (nx3318)) ;
    nor02ii ix5975 (.Y (nx5974), .A0 (nx3034), .A1 (nx5917)) ;
    nand02 ix5978 (.Y (nx5977), .A0 (write_base_data_out_4), .A1 (nx3170)) ;
    nand03 ix3559 (.Y (mem_addr_out[6]), .A0 (nx5980), .A1 (nx6901), .A2 (nx6026
           )) ;
    aoi22 ix5981 (.Y (nx5980), .A0 (nx3550), .A1 (nx6771), .B0 (nx3504), .B1 (
          nx6801)) ;
    xor2 ix3551 (.Y (nx3550), .A0 (nx5983), .A1 (nx5986)) ;
    aoi22 ix5984 (.Y (nx5983), .A0 (img_addr_offset_5), .A1 (img_base_addr_5), .B0 (
          nx3374), .B1 (nx3408)) ;
    dffs_ni img_base_addr_inst_reg_q_6 (.Q (img_base_addr_6), .QB (nx6009), .D (
            nx3389), .CLK (clk), .S (reset)) ;
    oai21 ix3529 (.Y (nx3528), .A0 (nx5991), .A1 (nx6006), .B0 (nx3522)) ;
    dffs_ni reg_write_base_reg_q_6 (.Q (write_base_data_out_6), .QB (nx5996), .D (
            nx3349), .CLK (nx6637), .S (reset)) ;
    xnor2 ix5999 (.Y (nx5998), .A0 (nx6000), .A1 (nx6003)) ;
    aoi22 ix6001 (.Y (nx6000), .A0 (write_base_data_out_5), .A1 (
          new_size_squared_out_5), .B0 (nx3294), .B1 (nx3296)) ;
    dffr reg_write_base_prev_reg_q_6 (.Q (\$dummy [122]), .QB (nx5991), .D (
         nx3379), .CLK (clk), .R (reset)) ;
    nor02_2x ix6007 (.Y (nx6006), .A0 (nx3242), .A1 (write_base_prev_data_out_5)
             ) ;
    nand02 ix3523 (.Y (nx3522), .A0 (nx6006), .A1 (nx5991)) ;
    aoi21 ix3543 (.Y (nx3542), .A0 (nx5945), .A1 (nx6013), .B0 (nx3536)) ;
    dffr reg_img_addr_offset_6 (.Q (img_addr_offset_6), .QB (nx6013), .D (nx3399
         ), .CLK (clk), .R (nx6807)) ;
    xor2 ix3505 (.Y (nx3504), .A0 (nx6017), .A1 (nx6020)) ;
    aoi22 ix6018 (.Y (nx6017), .A0 (write_base_data_out_5), .A1 (
          bias_offset_data_out_5), .B0 (nx3354), .B1 (nx3362)) ;
    dffr reg_bias_offset_reg_q_6 (.Q (bias_offset_data_out_6), .QB (nx6025), .D (
         nx3369), .CLK (clk), .R (reset)) ;
    aoi21 ix875 (.Y (nx874), .A0 (nx4246), .A1 (nx4239), .B0 (nx868)) ;
    aoi222 ix6027 (.Y (nx6026), .A0 (addr1_data_6), .A1 (nx6815), .B0 (nx3448), 
           .B1 (nx6795), .C0 (nx6651), .C1 (nx3466)) ;
    dffr reg_addr1_data_6 (.Q (addr1_data_6), .QB (nx6031), .D (nx3359), .CLK (
         clk), .R (reset)) ;
    xnor2 ix3449 (.Y (nx3448), .A0 (nx3426), .A1 (nx6034)) ;
    oai22 ix3427 (.Y (nx3426), .A0 (nx5968), .A1 (nx5971), .B0 (nx4251), .B1 (
          nx5938)) ;
    xnor2 ix3467 (.Y (nx3466), .A0 (nx6037), .A1 (nx6039)) ;
    nor02ii ix6038 (.Y (nx6037), .A0 (nx3318), .A1 (nx5974)) ;
    oai21 ix6040 (.Y (nx6039), .A0 (nx3312), .A1 (write_base_data_out_6), .B0 (
          nx6042)) ;
    nand02 ix6043 (.Y (nx6042), .A0 (write_base_data_out_6), .A1 (nx3312)) ;
    nand03 ix3699 (.Y (mem_addr_out[7]), .A0 (nx6045), .A1 (nx6901), .A2 (nx6081
           )) ;
    aoi22 ix6046 (.Y (nx6045), .A0 (nx3690), .A1 (nx6771), .B0 (nx3644), .B1 (
          nx6803)) ;
    xnor2 ix3691 (.Y (nx3690), .A0 (nx3654), .A1 (nx6049)) ;
    oai22 ix3655 (.Y (nx3654), .A0 (nx5983), .A1 (nx5986), .B0 (nx6013), .B1 (
          nx6009)) ;
    dffr img_base_addr_inst_reg_q_7 (.Q (img_base_addr_7), .QB (\$dummy [123]), 
         .D (nx3449), .CLK (clk), .R (reset)) ;
    xnor2 ix3669 (.Y (nx3668), .A0 (write_base_prev_data_out_7), .A1 (nx3522)) ;
    dffr reg_write_base_prev_reg_q_7 (.Q (write_base_prev_data_out_7), .QB (
         \$dummy [124]), .D (nx3439), .CLK (clk), .R (reset)) ;
    dffr reg_write_base_reg_q_7 (.Q (write_base_data_out_7), .QB (nx6062), .D (
         nx3409), .CLK (nx6637), .R (reset)) ;
    xnor2 ix3579 (.Y (nx3578), .A0 (nx3574), .A1 (nx6060)) ;
    oai22 ix3575 (.Y (nx3574), .A0 (nx6000), .A1 (nx6003), .B0 (nx5996), .B1 (
          nx4377)) ;
    oai21 ix6068 (.Y (nx6067), .A0 (nx3536), .A1 (img_addr_offset_7), .B0 (
          nx6069)) ;
    nand02 ix6070 (.Y (nx6069), .A0 (img_addr_offset_7), .A1 (nx3536)) ;
    dffr reg_img_addr_offset_7 (.Q (img_addr_offset_7), .QB (nx6071), .D (nx3459
         ), .CLK (clk), .R (nx6809)) ;
    xnor2 ix3645 (.Y (nx3644), .A0 (nx3634), .A1 (nx6075)) ;
    oai22 ix3635 (.Y (nx3634), .A0 (nx6017), .A1 (nx6020), .B0 (nx5996), .B1 (
          nx6025)) ;
    dffr reg_bias_offset_reg_q_7 (.Q (bias_offset_data_out_7), .QB (nx6079), .D (
         nx3429), .CLK (clk), .R (reset)) ;
    aoi222 ix6082 (.Y (nx6081), .A0 (addr1_data_7), .A1 (nx6817), .B0 (nx6653), 
           .B1 (nx3606), .C0 (nx3588), .C1 (nx6795)) ;
    oai21 ix6086 (.Y (nx6085), .A0 (nx3470), .A1 (addr1_data_7), .B0 (nx6088)) ;
    nand02 ix6089 (.Y (nx6088), .A0 (addr1_data_7), .A1 (nx3470)) ;
    dffr reg_addr1_data_7 (.Q (addr1_data_7), .QB (nx6090), .D (nx3419), .CLK (
         clk), .R (reset)) ;
    xnor2 ix3607 (.Y (nx3606), .A0 (nx3460), .A1 (nx3598)) ;
    nand02 ix3461 (.Y (nx3460), .A0 (nx6039), .A1 (nx6037)) ;
    aoi21 ix3599 (.Y (nx3598), .A0 (nx6042), .A1 (nx6062), .B0 (nx3592)) ;
    xor2 ix3589 (.Y (nx3588), .A0 (nx6097), .A1 (nx6100)) ;
    aoi22 ix6098 (.Y (nx6097), .A0 (write_offset_data_out_6), .A1 (
          write_base_data_out_6), .B0 (nx3426), .B1 (nx3446)) ;
    nand03 ix3839 (.Y (mem_addr_out[8]), .A0 (nx6103), .A1 (nx6901), .A2 (nx6149
           )) ;
    aoi22 ix6104 (.Y (nx6103), .A0 (nx3830), .A1 (nx6771), .B0 (nx3784), .B1 (
          nx6803)) ;
    xor2 ix3831 (.Y (nx3830), .A0 (nx6106), .A1 (nx6109)) ;
    aoi22 ix6107 (.Y (nx6106), .A0 (img_addr_offset_7), .A1 (img_base_addr_7), .B0 (
          nx3654), .B1 (nx3688)) ;
    dffr img_base_addr_inst_reg_q_8 (.Q (img_base_addr_8), .QB (nx6132), .D (
         nx3509), .CLK (clk), .R (reset)) ;
    oai21 ix3809 (.Y (nx3808), .A0 (nx6114), .A1 (nx6129), .B0 (nx3802)) ;
    dffs_ni reg_write_base_reg_q_8 (.Q (write_base_data_out_8), .QB (nx6119), .D (
            nx3469), .CLK (nx6637), .S (reset)) ;
    xnor2 ix6122 (.Y (nx6121), .A0 (nx6123), .A1 (nx6126)) ;
    aoi22 ix6124 (.Y (nx6123), .A0 (write_base_data_out_7), .A1 (
          new_size_squared_out_7), .B0 (nx3574), .B1 (nx3576)) ;
    dffr reg_write_base_prev_reg_q_8 (.Q (\$dummy [125]), .QB (nx6114), .D (
         nx3499), .CLK (clk), .R (reset)) ;
    nor02_2x ix6130 (.Y (nx6129), .A0 (nx3522), .A1 (write_base_prev_data_out_7)
             ) ;
    nand02 ix3803 (.Y (nx3802), .A0 (nx6129), .A1 (nx6114)) ;
    aoi21 ix3823 (.Y (nx3822), .A0 (nx6069), .A1 (nx6136), .B0 (nx3816)) ;
    dffr reg_img_addr_offset_8 (.Q (img_addr_offset_8), .QB (nx6136), .D (nx3519
         ), .CLK (clk), .R (nx6809)) ;
    xor2 ix3785 (.Y (nx3784), .A0 (nx6140), .A1 (nx6143)) ;
    aoi22 ix6141 (.Y (nx6140), .A0 (write_base_data_out_7), .A1 (
          bias_offset_data_out_7), .B0 (nx3634), .B1 (nx3642)) ;
    dffr reg_bias_offset_reg_q_8 (.Q (bias_offset_data_out_8), .QB (nx6148), .D (
         nx3489), .CLK (clk), .R (reset)) ;
    aoi21 ix925 (.Y (nx924), .A0 (nx4223), .A1 (nx4217), .B0 (nx918)) ;
    aoi222 ix6150 (.Y (nx6149), .A0 (addr1_data_8), .A1 (nx6817), .B0 (nx3728), 
           .B1 (nx6797), .C0 (nx6653), .C1 (nx3746)) ;
    dffr reg_addr1_data_8 (.Q (addr1_data_8), .QB (nx6154), .D (nx3479), .CLK (
         clk), .R (reset)) ;
    xnor2 ix3729 (.Y (nx3728), .A0 (nx3706), .A1 (nx6157)) ;
    oai22 ix3707 (.Y (nx3706), .A0 (nx6097), .A1 (nx6100), .B0 (nx4229), .B1 (
          nx6062)) ;
    xnor2 ix3747 (.Y (nx3746), .A0 (nx6160), .A1 (nx6162)) ;
    nor02_2x ix6161 (.Y (nx6160), .A0 (nx3598), .A1 (nx3460)) ;
    oai21 ix6163 (.Y (nx6162), .A0 (nx3592), .A1 (write_base_data_out_8), .B0 (
          nx6164)) ;
    nand02 ix6165 (.Y (nx6164), .A0 (write_base_data_out_8), .A1 (nx3592)) ;
    nand03 ix3979 (.Y (mem_addr_out[9]), .A0 (nx6167), .A1 (nx6901), .A2 (nx6203
           )) ;
    aoi22 ix6168 (.Y (nx6167), .A0 (nx3970), .A1 (nx6771), .B0 (nx3924), .B1 (
          nx6803)) ;
    xnor2 ix3971 (.Y (nx3970), .A0 (nx3934), .A1 (nx6171)) ;
    oai22 ix3935 (.Y (nx3934), .A0 (nx6106), .A1 (nx6109), .B0 (nx6136), .B1 (
          nx6132)) ;
    dffr img_base_addr_inst_reg_q_9 (.Q (img_base_addr_9), .QB (\$dummy [126]), 
         .D (nx3569), .CLK (clk), .R (reset)) ;
    xnor2 ix3949 (.Y (nx3948), .A0 (write_base_prev_data_out_9), .A1 (nx3802)) ;
    dffr reg_write_base_prev_reg_q_9 (.Q (write_base_prev_data_out_9), .QB (
         \$dummy [127]), .D (nx3559), .CLK (clk), .R (reset)) ;
    dffs_ni reg_write_base_reg_q_9 (.Q (write_base_data_out_9), .QB (nx6184), .D (
            nx3529), .CLK (nx6637), .S (reset)) ;
    xnor2 ix3859 (.Y (nx3858), .A0 (nx3854), .A1 (nx6182)) ;
    oai22 ix3855 (.Y (nx3854), .A0 (nx6123), .A1 (nx6126), .B0 (nx6119), .B1 (
          nx4363)) ;
    oai21 ix6190 (.Y (nx6189), .A0 (nx3816), .A1 (img_addr_offset_9), .B0 (
          nx6191)) ;
    nand02 ix6192 (.Y (nx6191), .A0 (img_addr_offset_9), .A1 (nx3816)) ;
    dffr reg_img_addr_offset_9 (.Q (img_addr_offset_9), .QB (nx6193), .D (nx3579
         ), .CLK (clk), .R (nx6809)) ;
    xnor2 ix3925 (.Y (nx3924), .A0 (nx3914), .A1 (nx6197)) ;
    oai22 ix3915 (.Y (nx3914), .A0 (nx6140), .A1 (nx6143), .B0 (nx6119), .B1 (
          nx6148)) ;
    dffr reg_bias_offset_reg_q_9 (.Q (bias_offset_data_out_9), .QB (nx6201), .D (
         nx3549), .CLK (clk), .R (reset)) ;
    aoi222 ix6204 (.Y (nx6203), .A0 (addr1_data_9), .A1 (nx6817), .B0 (nx6653), 
           .B1 (nx3886), .C0 (nx3868), .C1 (nx6797)) ;
    oai21 ix6208 (.Y (nx6207), .A0 (nx3750), .A1 (addr1_data_9), .B0 (nx6210)) ;
    nand02 ix6211 (.Y (nx6210), .A0 (addr1_data_9), .A1 (nx3750)) ;
    dffr reg_addr1_data_9 (.Q (addr1_data_9), .QB (nx6212), .D (nx3539), .CLK (
         clk), .R (reset)) ;
    xnor2 ix3887 (.Y (nx3886), .A0 (nx3740), .A1 (nx3878)) ;
    nand02 ix3741 (.Y (nx3740), .A0 (nx6162), .A1 (nx6160)) ;
    aoi21 ix3879 (.Y (nx3878), .A0 (nx6164), .A1 (nx6184), .B0 (nx3872)) ;
    xor2 ix3869 (.Y (nx3868), .A0 (nx6219), .A1 (nx6222)) ;
    aoi22 ix6220 (.Y (nx6219), .A0 (write_offset_data_out_8), .A1 (
          write_base_data_out_8), .B0 (nx3706), .B1 (nx3726)) ;
    nand03 ix4119 (.Y (mem_addr_out[10]), .A0 (nx6225), .A1 (nx6901), .A2 (
           nx6271)) ;
    aoi22 ix6226 (.Y (nx6225), .A0 (nx4110), .A1 (nx6771), .B0 (nx4064), .B1 (
          nx6803)) ;
    xor2 ix4111 (.Y (nx4110), .A0 (nx6228), .A1 (nx6231)) ;
    aoi22 ix6229 (.Y (nx6228), .A0 (img_addr_offset_9), .A1 (img_base_addr_9), .B0 (
          nx3934), .B1 (nx3968)) ;
    dffr img_base_addr_inst_reg_q_10 (.Q (img_base_addr_10), .QB (nx6254), .D (
         nx3629), .CLK (clk), .R (reset)) ;
    oai21 ix4089 (.Y (nx4088), .A0 (nx6236), .A1 (nx6251), .B0 (nx4082)) ;
    dffr reg_write_base_reg_q_10 (.Q (write_base_data_out_10), .QB (nx6241), .D (
         nx3589), .CLK (nx6637), .R (reset)) ;
    xnor2 ix6244 (.Y (nx6243), .A0 (nx6245), .A1 (nx6248)) ;
    aoi22 ix6246 (.Y (nx6245), .A0 (write_base_data_out_9), .A1 (
          new_size_squared_out_9), .B0 (nx3854), .B1 (nx3856)) ;
    dffr reg_write_base_prev_reg_q_10 (.Q (\$dummy [128]), .QB (nx6236), .D (
         nx3619), .CLK (clk), .R (reset)) ;
    nor02_2x ix6252 (.Y (nx6251), .A0 (nx3802), .A1 (write_base_prev_data_out_9)
             ) ;
    nand02 ix4083 (.Y (nx4082), .A0 (nx6251), .A1 (nx6236)) ;
    aoi21 ix4103 (.Y (nx4102), .A0 (nx6191), .A1 (nx6258), .B0 (nx4096)) ;
    dffr reg_img_addr_offset_10 (.Q (img_addr_offset_10), .QB (nx6258), .D (
         nx3639), .CLK (clk), .R (nx6809)) ;
    xor2 ix4065 (.Y (nx4064), .A0 (nx6262), .A1 (nx6265)) ;
    aoi22 ix6263 (.Y (nx6262), .A0 (write_base_data_out_9), .A1 (
          bias_offset_data_out_9), .B0 (nx3914), .B1 (nx3922)) ;
    dffr reg_bias_offset_reg_q_10 (.Q (bias_offset_data_out_10), .QB (nx6270), .D (
         nx3609), .CLK (clk), .R (reset)) ;
    aoi21 ix971 (.Y (nx970), .A0 (nx4207), .A1 (nx4200), .B0 (nx964)) ;
    aoi222 ix6272 (.Y (nx6271), .A0 (addr1_data_10), .A1 (nx6817), .B0 (nx4008)
           , .B1 (nx6797), .C0 (nx6653), .C1 (nx4026)) ;
    dffr reg_addr1_data_10 (.Q (addr1_data_10), .QB (nx6276), .D (nx3599), .CLK (
         clk), .R (reset)) ;
    xnor2 ix4009 (.Y (nx4008), .A0 (nx3986), .A1 (nx6279)) ;
    oai22 ix3987 (.Y (nx3986), .A0 (nx6219), .A1 (nx6222), .B0 (nx4301), .B1 (
          nx6184)) ;
    xnor2 ix4027 (.Y (nx4026), .A0 (nx6282), .A1 (nx6284)) ;
    nor02_2x ix6283 (.Y (nx6282), .A0 (nx3878), .A1 (nx3740)) ;
    oai21 ix6285 (.Y (nx6284), .A0 (nx3872), .A1 (write_base_data_out_10), .B0 (
          nx6286)) ;
    nand02 ix6287 (.Y (nx6286), .A0 (write_base_data_out_10), .A1 (nx3872)) ;
    nand03 ix4259 (.Y (mem_addr_out[11]), .A0 (nx6289), .A1 (nx6901), .A2 (
           nx6325)) ;
    aoi22 ix6290 (.Y (nx6289), .A0 (nx4250), .A1 (nx6771), .B0 (nx4204), .B1 (
          nx6803)) ;
    xnor2 ix4251 (.Y (nx4250), .A0 (nx4214), .A1 (nx6293)) ;
    oai22 ix4215 (.Y (nx4214), .A0 (nx6228), .A1 (nx6231), .B0 (nx6258), .B1 (
          nx6254)) ;
    dffs_ni img_base_addr_inst_reg_q_11 (.Q (img_base_addr_11), .QB (
            \$dummy [129]), .D (nx3689), .CLK (clk), .S (reset)) ;
    xnor2 ix4229 (.Y (nx4228), .A0 (write_base_prev_data_out_11), .A1 (nx4082)
          ) ;
    dffr reg_write_base_prev_reg_q_11 (.Q (write_base_prev_data_out_11), .QB (
         \$dummy [130]), .D (nx3679), .CLK (clk), .R (reset)) ;
    dffs_ni reg_write_base_reg_q_11 (.Q (write_base_data_out_11), .QB (nx6306), 
            .D (nx3649), .CLK (nx6637), .S (reset)) ;
    xnor2 ix4139 (.Y (nx4138), .A0 (nx4134), .A1 (nx6304)) ;
    oai22 ix4135 (.Y (nx4134), .A0 (nx6245), .A1 (nx6248), .B0 (nx6241), .B1 (
          nx4349)) ;
    oai21 ix6312 (.Y (nx6311), .A0 (nx4096), .A1 (img_addr_offset_11), .B0 (
          nx6313)) ;
    nand02 ix6314 (.Y (nx6313), .A0 (img_addr_offset_11), .A1 (nx4096)) ;
    dffr reg_img_addr_offset_11 (.Q (img_addr_offset_11), .QB (nx6315), .D (
         nx3699), .CLK (clk), .R (nx6809)) ;
    xnor2 ix4205 (.Y (nx4204), .A0 (nx4194), .A1 (nx6319)) ;
    oai22 ix4195 (.Y (nx4194), .A0 (nx6262), .A1 (nx6265), .B0 (nx6241), .B1 (
          nx6270)) ;
    dffr reg_bias_offset_reg_q_11 (.Q (bias_offset_data_out_11), .QB (nx6323), .D (
         nx3669), .CLK (clk), .R (reset)) ;
    aoi222 ix6326 (.Y (nx6325), .A0 (addr1_data_11), .A1 (nx6817), .B0 (nx6653)
           , .B1 (nx4166), .C0 (nx4148), .C1 (nx6797)) ;
    oai21 ix6330 (.Y (nx6329), .A0 (nx4030), .A1 (addr1_data_11), .B0 (nx6332)
          ) ;
    nand02 ix6333 (.Y (nx6332), .A0 (addr1_data_11), .A1 (nx4030)) ;
    dffr reg_addr1_data_11 (.Q (addr1_data_11), .QB (nx6334), .D (nx3659), .CLK (
         clk), .R (reset)) ;
    xnor2 ix4167 (.Y (nx4166), .A0 (nx4020), .A1 (nx4158)) ;
    nand02 ix4021 (.Y (nx4020), .A0 (nx6284), .A1 (nx6282)) ;
    aoi21 ix4159 (.Y (nx4158), .A0 (nx6286), .A1 (nx6306), .B0 (nx4152)) ;
    xor2 ix4149 (.Y (nx4148), .A0 (nx6341), .A1 (nx6344)) ;
    aoi22 ix6342 (.Y (nx6341), .A0 (write_offset_data_out_10), .A1 (
          write_base_data_out_10), .B0 (nx3986), .B1 (nx4006)) ;
    nand03 ix4399 (.Y (mem_addr_out[12]), .A0 (nx6347), .A1 (nx6901), .A2 (
           nx6393)) ;
    aoi22 ix6348 (.Y (nx6347), .A0 (nx4390), .A1 (nx6773), .B0 (nx4344), .B1 (
          nx6803)) ;
    xor2 ix4391 (.Y (nx4390), .A0 (nx6350), .A1 (nx6353)) ;
    aoi22 ix6351 (.Y (nx6350), .A0 (img_addr_offset_11), .A1 (img_base_addr_11)
          , .B0 (nx4214), .B1 (nx4248)) ;
    dffs_ni img_base_addr_inst_reg_q_12 (.Q (img_base_addr_12), .QB (nx6376), .D (
            nx3749), .CLK (clk), .S (reset)) ;
    oai21 ix4369 (.Y (nx4368), .A0 (nx6358), .A1 (nx6373), .B0 (nx4362)) ;
    dffs_ni reg_write_base_reg_q_12 (.Q (write_base_data_out_12), .QB (nx6363), 
            .D (nx3709), .CLK (nx6639), .S (reset)) ;
    xnor2 ix6366 (.Y (nx6365), .A0 (nx7445), .A1 (nx6370)) ;
    aoi22 ix6368 (.Y (nx6367), .A0 (write_base_data_out_11), .A1 (
          new_size_squared_out_11), .B0 (nx4134), .B1 (nx4136)) ;
    dffr reg_write_base_prev_reg_q_12 (.Q (\$dummy [131]), .QB (nx6358), .D (
         nx3739), .CLK (clk), .R (reset)) ;
    nor02_2x ix6374 (.Y (nx6373), .A0 (nx4082), .A1 (write_base_prev_data_out_11
             )) ;
    nand02 ix4363 (.Y (nx4362), .A0 (nx6373), .A1 (nx6358)) ;
    aoi21 ix4383 (.Y (nx4382), .A0 (nx6313), .A1 (nx6380), .B0 (nx4376)) ;
    dffr reg_img_addr_offset_12 (.Q (img_addr_offset_12), .QB (nx6380), .D (
         nx3759), .CLK (clk), .R (nx6809)) ;
    xor2 ix4345 (.Y (nx4344), .A0 (nx6384), .A1 (nx6387)) ;
    aoi22 ix6385 (.Y (nx6384), .A0 (write_base_data_out_11), .A1 (
          bias_offset_data_out_11), .B0 (nx4194), .B1 (nx4202)) ;
    dffr reg_bias_offset_reg_q_12 (.Q (bias_offset_data_out_12), .QB (nx6392), .D (
         nx3729), .CLK (clk), .R (reset)) ;
    aoi21 ix1019 (.Y (nx1018), .A0 (nx4191), .A1 (nx4183), .B0 (nx1012)) ;
    aoi222 ix6394 (.Y (nx6393), .A0 (addr1_data_12), .A1 (nx6817), .B0 (nx6653)
           , .B1 (nx4306), .C0 (nx4288), .C1 (nx6797)) ;
    dffr reg_addr1_data_12 (.Q (addr1_data_12), .QB (nx6398), .D (nx3719), .CLK (
         clk), .R (reset)) ;
    xnor2 ix4307 (.Y (nx4306), .A0 (nx6400), .A1 (nx6402)) ;
    nor02_2x ix6401 (.Y (nx6400), .A0 (nx4158), .A1 (nx4020)) ;
    oai21 ix6403 (.Y (nx6402), .A0 (nx4152), .A1 (write_base_data_out_12), .B0 (
          nx6404)) ;
    nand02 ix6405 (.Y (nx6404), .A0 (write_base_data_out_12), .A1 (nx4152)) ;
    xnor2 ix4289 (.Y (nx4288), .A0 (nx4266), .A1 (nx6408)) ;
    oai22 ix4267 (.Y (nx4266), .A0 (nx6341), .A1 (nx6344), .B0 (nx4303), .B1 (
          nx6306)) ;
    nand03 ix4539 (.Y (mem_addr_out[13]), .A0 (nx6411), .A1 (nx6903), .A2 (
           nx6447)) ;
    aoi22 ix6412 (.Y (nx6411), .A0 (nx4530), .A1 (nx6773), .B0 (nx4484), .B1 (
          nx6803)) ;
    xnor2 ix4531 (.Y (nx4530), .A0 (nx4494), .A1 (nx6415)) ;
    oai22 ix4495 (.Y (nx4494), .A0 (nx6350), .A1 (nx6353), .B0 (nx6380), .B1 (
          nx6376)) ;
    dffr img_base_addr_inst_reg_q_13 (.Q (img_base_addr_13), .QB (\$dummy [132])
         , .D (nx3809), .CLK (clk), .R (reset)) ;
    xnor2 ix4509 (.Y (nx4508), .A0 (write_base_prev_data_out_13), .A1 (nx4362)
          ) ;
    dffr reg_write_base_prev_reg_q_13 (.Q (write_base_prev_data_out_13), .QB (
         \$dummy [133]), .D (nx3799), .CLK (clk), .R (reset)) ;
    dffr reg_write_base_reg_q_13 (.Q (write_base_data_out_13), .QB (nx6428), .D (
         nx3769), .CLK (nx6639), .R (reset)) ;
    xnor2 ix4419 (.Y (nx4418), .A0 (nx4414), .A1 (nx6426)) ;
    oai21 ix6434 (.Y (nx6433), .A0 (nx4376), .A1 (img_addr_offset_13), .B0 (
          nx6435)) ;
    nand02 ix6436 (.Y (nx6435), .A0 (img_addr_offset_13), .A1 (nx4376)) ;
    dffr reg_img_addr_offset_13 (.Q (img_addr_offset_13), .QB (nx6437), .D (
         nx3819), .CLK (clk), .R (nx6809)) ;
    xnor2 ix4485 (.Y (nx4484), .A0 (nx4474), .A1 (nx6441)) ;
    oai22 ix4475 (.Y (nx4474), .A0 (nx6384), .A1 (nx6387), .B0 (nx7363), .B1 (
          nx6392)) ;
    dffr reg_bias_offset_reg_q_13 (.Q (bias_offset_data_out_13), .QB (nx6445), .D (
         nx3789), .CLK (clk), .R (reset)) ;
    aoi222 ix6448 (.Y (nx6447), .A0 (addr1_data_13), .A1 (nx6817), .B0 (nx6653)
           , .B1 (nx4446), .C0 (nx4428), .C1 (nx6797)) ;
    oai21 ix6452 (.Y (nx6451), .A0 (nx4310), .A1 (addr1_data_13), .B0 (nx6454)
          ) ;
    nand02 ix6455 (.Y (nx6454), .A0 (addr1_data_13), .A1 (nx4310)) ;
    dffr reg_addr1_data_13 (.Q (addr1_data_13), .QB (nx6456), .D (nx3779), .CLK (
         clk), .R (reset)) ;
    xnor2 ix4447 (.Y (nx4446), .A0 (nx4300), .A1 (nx4438)) ;
    nand02 ix4301 (.Y (nx4300), .A0 (nx6402), .A1 (nx6400)) ;
    aoi21 ix4439 (.Y (nx4438), .A0 (nx6404), .A1 (nx6428), .B0 (nx4432)) ;
    xor2 ix4429 (.Y (nx4428), .A0 (nx6463), .A1 (nx6466)) ;
    aoi22 ix6464 (.Y (nx6463), .A0 (write_offset_data_out_12), .A1 (
          write_base_data_out_12), .B0 (nx4266), .B1 (nx4286)) ;
    nand03 ix4679 (.Y (mem_addr_out[14]), .A0 (nx6469), .A1 (nx6903), .A2 (
           nx6511)) ;
    aoi22 ix6470 (.Y (nx6469), .A0 (nx4670), .A1 (nx6773), .B0 (nx4624), .B1 (
          nx2626)) ;
    xor2 ix4671 (.Y (nx4670), .A0 (nx6472), .A1 (nx6475)) ;
    aoi22 ix6473 (.Y (nx6472), .A0 (img_addr_offset_13), .A1 (img_base_addr_13)
          , .B0 (nx4494), .B1 (nx4528)) ;
    dffr img_base_addr_inst_reg_q_14 (.Q (img_base_addr_14), .QB (nx6496), .D (
         nx3869), .CLK (clk), .R (reset)) ;
    dffr reg_write_base_prev_reg_q_14 (.Q (\$dummy [134]), .QB (nx6493), .D (
         nx3859), .CLK (clk), .R (reset)) ;
    dffr reg_write_base_reg_q_14 (.Q (write_base_data_out_14), .QB (nx6484), .D (
         nx3829), .CLK (nx6639), .R (reset)) ;
    xnor2 ix6487 (.Y (nx6486), .A0 (nx6488), .A1 (nx6491)) ;
    nor02_2x ix6495 (.Y (nx6494), .A0 (nx4362), .A1 (write_base_prev_data_out_13
             )) ;
    dffr reg_img_addr_offset_14 (.Q (img_addr_offset_14), .QB (nx6500), .D (
         nx3879), .CLK (clk), .R (nx6811)) ;
    xor2 ix4625 (.Y (nx4624), .A0 (nx6502), .A1 (nx6505)) ;
    aoi22 ix6503 (.Y (nx6502), .A0 (write_base_data_out_13), .A1 (
          bias_offset_data_out_13), .B0 (nx4474), .B1 (nx4482)) ;
    dffr reg_bias_offset_reg_q_14 (.Q (bias_offset_data_out_14), .QB (nx6510), .D (
         nx3849), .CLK (clk), .R (reset)) ;
    aoi222 ix6512 (.Y (nx6511), .A0 (addr1_data_14), .A1 (nx6819), .B0 (nx6655)
           , .B1 (nx4586), .C0 (nx4568), .C1 (nx6797)) ;
    dffr reg_addr1_data_14 (.Q (addr1_data_14), .QB (nx6516), .D (nx3839), .CLK (
         clk), .R (reset)) ;
    xnor2 ix4587 (.Y (nx4586), .A0 (nx6518), .A1 (nx6520)) ;
    nor02_2x ix6519 (.Y (nx6518), .A0 (nx4438), .A1 (nx4300)) ;
    xnor2 ix4569 (.Y (nx4568), .A0 (nx4546), .A1 (nx6524)) ;
    oai22 ix4547 (.Y (nx4546), .A0 (nx6463), .A1 (nx6466), .B0 (nx4305), .B1 (
          nx6428)) ;
    nand03 ix4789 (.Y (mem_addr_out[15]), .A0 (nx6527), .A1 (nx6903), .A2 (
           nx6560)) ;
    aoi22 ix6528 (.Y (nx6527), .A0 (nx4746), .A1 (nx6655), .B0 (nx4780), .B1 (
          nx6773)) ;
    xnor2 ix4747 (.Y (nx4746), .A0 (nx4580), .A1 (nx4744)) ;
    nand02 ix4581 (.Y (nx4580), .A0 (nx6520), .A1 (nx6518)) ;
    xnor2 ix4745 (.Y (nx4744), .A0 (nx6532), .A1 (write_base_data_out_15)) ;
    nand02 ix6533 (.Y (nx6532), .A0 (write_base_data_out_14), .A1 (nx4432)) ;
    dffs_ni reg_write_base_reg_q_15 (.Q (write_base_data_out_15), .QB (
            \$dummy [135]), .D (nx3899), .CLK (nx6639), .S (reset)) ;
    xnor2 ix4781 (.Y (nx4780), .A0 (nx4756), .A1 (nx6543)) ;
    oai22 ix4757 (.Y (nx4756), .A0 (nx6472), .A1 (nx6475), .B0 (nx6500), .B1 (
          nx6496)) ;
    dffs_ni img_base_addr_inst_reg_q_15 (.Q (img_base_addr_15), .QB (
            \$dummy [136]), .D (nx3929), .CLK (clk), .S (reset)) ;
    xnor2 ix4765 (.Y (nx4764), .A0 (write_base_prev_data_out_15), .A1 (nx4642)
          ) ;
    dffr reg_write_base_prev_reg_q_15 (.Q (write_base_prev_data_out_15), .QB (
         \$dummy [137]), .D (nx3919), .CLK (clk), .R (reset)) ;
    nand02 ix4643 (.Y (nx4642), .A0 (nx6494), .A1 (nx6493)) ;
    dffr img_addr_offset_15 (.Q (\$dummy [138]), .QB (nx6558), .D (nx3939), .CLK (
         clk), .R (nx6811)) ;
    aoi222 ix6561 (.Y (nx6560), .A0 (nx4736), .A1 (nx6799), .B0 (addr1_data_15)
           , .B1 (nx6819), .C0 (nx4714), .C1 (nx2626)) ;
    xnor2 ix4737 (.Y (nx4736), .A0 (nx6563), .A1 (nx4734)) ;
    aoi22 ix6564 (.Y (nx6563), .A0 (write_offset_data_out_14), .A1 (
          write_base_data_out_14), .B0 (nx4546), .B1 (nx4566)) ;
    dffr reg_addr1_data_15 (.Q (addr1_data_15), .QB (nx6572), .D (nx3909), .CLK (
         clk), .R (reset)) ;
    xnor2 ix4715 (.Y (nx4714), .A0 (nx4686), .A1 (nx6576)) ;
    oai22 ix4687 (.Y (nx4686), .A0 (nx6502), .A1 (nx6505), .B0 (nx7365), .B1 (
          nx6510)) ;
    dffr reg_bias_offset_reg_q_15 (.Q (bias_offset_data_out_15), .QB (nx6580), .D (
         nx3889), .CLK (clk), .R (reset)) ;
    inv01 ix1965 (.Y (mem_data_out[0]), .A (nx6583)) ;
    aoi222 ix6584 (.Y (nx6583), .A0 (comp_unit_data2_in[0]), .A1 (nx6675), .B0 (
           comp_unit_data1_in[0]), .B1 (nx6683), .C0 (argmax_data_in[0]), .C1 (
           current_state_28)) ;
    inv01 ix1975 (.Y (mem_data_out[1]), .A (nx6586)) ;
    aoi222 ix6587 (.Y (nx6586), .A0 (comp_unit_data2_in[1]), .A1 (nx6677), .B0 (
           comp_unit_data1_in[1]), .B1 (nx6683), .C0 (argmax_data_in[1]), .C1 (
           current_state_28)) ;
    inv01 ix1985 (.Y (mem_data_out[2]), .A (nx6589)) ;
    aoi222 ix6590 (.Y (nx6589), .A0 (comp_unit_data2_in[2]), .A1 (nx6677), .B0 (
           comp_unit_data1_in[2]), .B1 (nx6683), .C0 (argmax_data_in[2]), .C1 (
           current_state_28)) ;
    inv01 ix1995 (.Y (mem_data_out[3]), .A (nx6592)) ;
    aoi222 ix6593 (.Y (nx6592), .A0 (comp_unit_data2_in[3]), .A1 (nx6677), .B0 (
           comp_unit_data1_in[3]), .B1 (nx6683), .C0 (argmax_data_in[3]), .C1 (
           current_state_28)) ;
    inv01 ix4567 (.Y (nx4566), .A (nx6524)) ;
    inv01 ix4529 (.Y (nx4528), .A (nx6415)) ;
    inv01 ix4483 (.Y (nx4482), .A (nx6441)) ;
    inv01 ix4287 (.Y (nx4286), .A (nx6408)) ;
    inv01 ix4249 (.Y (nx4248), .A (nx6293)) ;
    inv01 ix4203 (.Y (nx4202), .A (nx6319)) ;
    inv01 ix4137 (.Y (nx4136), .A (nx6304)) ;
    inv01 ix4007 (.Y (nx4006), .A (nx6279)) ;
    inv01 ix3969 (.Y (nx3968), .A (nx6171)) ;
    inv01 ix3923 (.Y (nx3922), .A (nx6197)) ;
    inv01 ix3857 (.Y (nx3856), .A (nx6182)) ;
    inv01 ix3727 (.Y (nx3726), .A (nx6157)) ;
    inv01 ix3689 (.Y (nx3688), .A (nx6049)) ;
    inv01 ix3643 (.Y (nx3642), .A (nx6075)) ;
    inv01 ix3577 (.Y (nx3576), .A (nx6060)) ;
    inv01 ix3447 (.Y (nx3446), .A (nx6034)) ;
    inv01 ix3409 (.Y (nx3408), .A (nx5925)) ;
    inv01 ix3363 (.Y (nx3362), .A (nx5951)) ;
    inv01 ix3297 (.Y (nx3296), .A (nx5936)) ;
    inv01 ix3159 (.Y (nx3158), .A (nx5913)) ;
    inv01 ix3121 (.Y (nx3120), .A (nx5794)) ;
    inv01 ix3075 (.Y (nx3074), .A (nx5820)) ;
    inv01 ix5839 (.Y (nx5838), .A (nx3034)) ;
    inv01 ix3005 (.Y (nx3004), .A (nx5805)) ;
    inv01 ix2951 (.Y (nx2950), .A (nx5809)) ;
    inv01 ix2885 (.Y (nx2884), .A (nx5783)) ;
    inv01 ix2833 (.Y (nx2832), .A (nx5673)) ;
    inv01 ix2795 (.Y (nx2794), .A (nx5703)) ;
    inv01 ix5502 (.Y (nx5501), .A (nx2502)) ;
    inv01 ix1685 (.Y (nx1464), .A (nx4499)) ;
    inv01 ix1711 (.Y (nx1463), .A (nx3989)) ;
    inv01 ix1529 (.Y (nx1528), .A (nx4080)) ;
    inv01 ix1807 (.Y (nx1461), .A (nx4009)) ;
    inv01 ix1429 (.Y (nx1428), .A (nx4681)) ;
    inv01 ix4704 (.Y (nx4703), .A (nx1152)) ;
    inv01 ix751 (.Y (nx750), .A (nx4295)) ;
    inv01 ix607 (.Y (nx606), .A (nx5155)) ;
    inv01 ix601 (.Y (nx600), .A (nx5157)) ;
    inv01 ix4884 (.Y (nx4883), .A (nx546)) ;
    inv01 ix321 (.Y (nx320), .A (nx5113)) ;
    inv01 ix6598 (.Y (nx6599), .A (current_state_13)) ;
    inv02 ix6600 (.Y (nx6601), .A (nx6599)) ;
    inv02 ix6602 (.Y (nx6603), .A (nx6599)) ;
    inv02 ix6604 (.Y (nx6605), .A (nx6599)) ;
    buf02 ix6606 (.Y (nx6607), .A (wind_width_count_0)) ;
    buf02 ix6608 (.Y (nx6609), .A (wind_width_count_0)) ;
    buf02 ix6610 (.Y (nx6611), .A (cache_width_count_4)) ;
    buf02 ix6612 (.Y (nx6613), .A (cache_width_count_4)) ;
    buf02 ix6614 (.Y (nx6615), .A (cache_width_count_2)) ;
    buf02 ix6616 (.Y (nx6617), .A (cache_width_count_2)) ;
    inv02 ix6618 (.Y (nx6619), .A (clk)) ;
    inv02 ix6620 (.Y (nx6621), .A (clk)) ;
    inv02 ix6622 (.Y (nx6623), .A (clk)) ;
    inv02 ix6624 (.Y (nx6625), .A (clk)) ;
    inv02 ix6626 (.Y (nx6627), .A (clk)) ;
    inv02 ix6628 (.Y (nx6629), .A (clk)) ;
    inv02 ix6630 (.Y (nx6631), .A (clk)) ;
    inv02 ix6632 (.Y (nx6633), .A (clk)) ;
    inv02 ix6634 (.Y (nx6635), .A (clk)) ;
    inv02 ix6636 (.Y (nx6637), .A (clk)) ;
    inv02 ix6638 (.Y (nx6639), .A (clk)) ;
    inv02 ix6640 (.Y (nx6641), .A (nx7294)) ;
    inv02 ix6642 (.Y (nx6643), .A (nx7294)) ;
    inv02 ix6650 (.Y (nx6651), .A (nx7043)) ;
    inv02 ix6652 (.Y (nx6653), .A (nx7043)) ;
    inv02 ix6654 (.Y (nx6655), .A (nx7043)) ;
    inv01 ix6656 (.Y (nx6657), .A (nx7293)) ;
    inv02 ix6658 (.Y (nx6659), .A (nx7077)) ;
    inv02 ix6662 (.Y (nx6663), .A (nx7077)) ;
    inv02 ix6664 (.Y (nx6665), .A (nx3981)) ;
    inv02 ix6666 (.Y (nx6667), .A (nx7009)) ;
    inv02 ix6672 (.Y (nx6673), .A (nx4149)) ;
    inv02 ix6674 (.Y (nx6675), .A (nx4149)) ;
    inv02 ix6676 (.Y (nx6677), .A (nx4149)) ;
    inv02 ix6678 (.Y (nx6679), .A (nx4129)) ;
    inv02 ix6680 (.Y (nx6681), .A (nx4129)) ;
    inv02 ix6682 (.Y (nx6683), .A (nx4129)) ;
    inv02 ix6684 (.Y (nx6685), .A (nx4711)) ;
    inv02 ix6686 (.Y (nx6687), .A (nx7033)) ;
    buf02 ix6688 (.Y (nx6689), .A (current_state_4)) ;
    buf02 ix6690 (.Y (nx6691), .A (current_state_4)) ;
    inv02 ix6692 (.Y (nx6693), .A (nx6823)) ;
    inv02 ix6694 (.Y (nx6695), .A (nx6823)) ;
    inv02 ix6698 (.Y (nx6699), .A (nx7081)) ;
    inv02 ix6704 (.Y (nx6705), .A (nx4109)) ;
    buf02 ix6712 (.Y (nx6713), .A (nx176)) ;
    inv01 ix6720 (.Y (nx6721), .A (nx348)) ;
    inv02 ix6722 (.Y (nx6723), .A (nx6721)) ;
    inv02 ix6724 (.Y (nx6725), .A (nx6721)) ;
    inv02 ix6726 (.Y (nx6727), .A (nx6721)) ;
    inv02 ix6730 (.Y (nx6731), .A (nx6729)) ;
    inv02 ix6732 (.Y (nx6733), .A (nx7087)) ;
    inv02 ix6734 (.Y (nx6735), .A (nx7087)) ;
    inv01 ix6736 (.Y (nx6737), .A (nx1192)) ;
    inv02 ix6738 (.Y (nx6739), .A (nx6737)) ;
    inv02 ix6740 (.Y (nx6741), .A (nx6737)) ;
    inv02 ix6742 (.Y (nx6743), .A (nx6737)) ;
    inv02 ix6748 (.Y (nx6749), .A (nx4553)) ;
    inv02 ix6762 (.Y (nx6763), .A (nx6897)) ;
    inv02 ix6764 (.Y (nx6765), .A (nx6897)) ;
    inv02 ix6766 (.Y (nx6767), .A (nx6897)) ;
    inv02 ix6768 (.Y (nx6769), .A (nx7107)) ;
    inv02 ix6770 (.Y (nx6771), .A (nx7107)) ;
    inv02 ix6772 (.Y (nx6773), .A (nx7107)) ;
    inv02 ix6780 (.Y (nx6781), .A (nx7095)) ;
    inv02 ix6786 (.Y (nx6787), .A (nx5728)) ;
    inv02 ix6794 (.Y (nx6795), .A (nx6793)) ;
    inv02 ix6796 (.Y (nx6797), .A (nx6793)) ;
    inv02 ix6798 (.Y (nx6799), .A (nx6793)) ;
    inv02 ix6806 (.Y (nx6807), .A (nx6805)) ;
    inv02 ix6808 (.Y (nx6809), .A (nx6805)) ;
    inv02 ix6810 (.Y (nx6811), .A (nx6805)) ;
    inv02 ix6814 (.Y (nx6815), .A (nx6813)) ;
    inv02 ix6816 (.Y (nx6817), .A (nx6813)) ;
    inv02 ix6818 (.Y (nx6819), .A (nx6813)) ;
    inv02 ix6820 (.Y (nx6821), .A (current_state_9)) ;
    inv02 ix6822 (.Y (nx6823), .A (current_state_9)) ;
    inv02 ix6824 (.Y (nx6825), .A (nx1516)) ;
    inv02 ix6826 (.Y (nx6827), .A (nx1516)) ;
    inv02 ix6828 (.Y (nx6829), .A (nx730)) ;
    inv02 ix6830 (.Y (nx6831), .A (nx6981)) ;
    inv02 ix6832 (.Y (nx6833), .A (nx6981)) ;
    buf02 ix6834 (.Y (nx6835), .A (nx4717)) ;
    buf02 ix6836 (.Y (nx6837), .A (nx4717)) ;
    buf02 ix6838 (.Y (nx6839), .A (nx4961)) ;
    inv02 ix6850 (.Y (nx6851), .A (current_state_18)) ;
    inv02 ix6854 (.Y (nx6855), .A (nx6985)) ;
    inv02 ix6856 (.Y (nx6857), .A (nx6985)) ;
    inv02 ix6858 (.Y (nx6859), .A (nx6985)) ;
    inv02 ix6870 (.Y (nx6871), .A (nx2536)) ;
    inv02 ix6896 (.Y (nx6897), .A (nx2098)) ;
    inv02 ix6898 (.Y (nx6899), .A (current_state_28)) ;
    inv02 ix6900 (.Y (nx6901), .A (current_state_28)) ;
    inv02 ix6902 (.Y (nx6903), .A (current_state_28)) ;
    buf02 ix6926 (.Y (nx6927), .A (comp_unit_operation)) ;
    buf02 ix6928 (.Y (nx6929), .A (comp_unit_operation)) ;
    inv01 ix6930 (.Y (nx6931), .A (nx7145)) ;
    inv01 ix6932 (.Y (nx6933), .A (nx7145)) ;
    nor02_2x ix1493 (.Y (nx1492), .A0 (nx4129), .A1 (nx7294)) ;
    nor02ii ix3960 (.Y (nx3959), .A0 (nx6927), .A1 (layer_type_out_1)) ;
    nor02ii ix1579 (.Y (nx1578), .A0 (nx3975), .A1 (io_ready_in)) ;
    and03 ix1801 (.Y (nx1800), .A0 (nx1419), .A1 (nx6939), .A2 (nx4017)) ;
    inv01 ix6938 (.Y (nx6939), .A (nx4519)) ;
    and04 ix3990 (.Y (nx3989), .A0 (nx4111), .A1 (nx4447), .A2 (nx4469), .A3 (
          nx4497)) ;
    mux21_ni ix1621 (.Y (nx1620), .A0 (nx4111), .A1 (nx1610), .S0 (nx1516)) ;
    nor02ii ix1603 (.Y (nx1602), .A0 (nx4009), .A1 (nx7021)) ;
    nor02ii ix167 (.Y (nx4109), .A0 (layer_type_out_1), .A1 (nx6927)) ;
    and02 ix4010 (.Y (nx4009), .A0 (nx3967), .A1 (nx7009)) ;
    nor02ii ix113 (.Y (nx112), .A0 (nx4017), .A1 (nx1419)) ;
    and04 ix4018 (.Y (nx4017), .A0 (nflt_layer_out_0), .A1 (nx4039), .A2 (nx4053
          ), .A3 (nx6941)) ;
    inv01 ix6940 (.Y (nx6941), .A (nflt_layer_out_3)) ;
    mux21 ix4028 (.Y (nx4027), .A0 (nx4019), .A1 (mem_data_in[0]), .S0 (nx6689)
          ) ;
    nor02ii ix4034 (.Y (nx4033), .A0 (nx6689), .A1 (nx4073)) ;
    and02 ix4046 (.Y (nx4045), .A0 (nx4019), .A1 (nx4039)) ;
    xor2 ix4058 (.Y (nx4057), .A0 (nx4053), .A1 (nx4045)) ;
    and03 ix4068 (.Y (nx4067), .A0 (nx4019), .A1 (nx4039), .A2 (nx4053)) ;
    or02 ix4081 (.Y (nx4080), .A0 (nx7009), .A1 (nx7021)) ;
    nand04 ix4114 (.Y (nx1516), .A0 (nx3967), .A1 (nx7009), .A2 (nx4073), .A3 (
           nx6823)) ;
    and02 ix4120 (.Y (nx4119), .A0 (nx6823), .A1 (nx7009)) ;
    xor2 ix4158 (.Y (nx4157), .A0 (nx4307), .A1 (new_size_squared_out_15)) ;
    xor2 ix4164 (.Y (nx4163), .A0 (nx4307), .A1 (nx1058)) ;
    nor02ii ix1059 (.Y (nx1058), .A0 (nx4175), .A1 (write_offset_data_out_14)) ;
    ao22 ix2190 (.Y (nx2189), .A0 (nx1064), .A1 (nx6981), .B0 (
         write_offset_data_out_14), .B1 (nx7087)) ;
    nor02ii ix1013 (.Y (nx1012), .A0 (nx4191), .A1 (write_offset_data_out_12)) ;
    ao22 ix2150 (.Y (nx2149), .A0 (nx1018), .A1 (nx6981), .B0 (
         write_offset_data_out_12), .B1 (nx7087)) ;
    nor02ii ix965 (.Y (nx964), .A0 (nx4207), .A1 (write_offset_data_out_10)) ;
    ao22 ix2110 (.Y (nx2109), .A0 (nx970), .A1 (nx6981), .B0 (
         write_offset_data_out_10), .B1 (nx7087)) ;
    nor02ii ix919 (.Y (nx918), .A0 (nx4223), .A1 (write_offset_data_out_8)) ;
    ao22 ix2070 (.Y (nx2069), .A0 (nx924), .A1 (nx6983), .B0 (
         write_offset_data_out_8), .B1 (nx7087)) ;
    nor02ii ix733 (.Y (nx6729), .A0 (nx6983), .A1 (nx4123)) ;
    nand02 ix4234 (.Y (nx730), .A0 (nx4129), .A1 (nx4149)) ;
    nor02ii ix869 (.Y (nx868), .A0 (nx4246), .A1 (write_offset_data_out_6)) ;
    ao22 ix2030 (.Y (nx2029), .A0 (nx874), .A1 (nx6983), .B0 (
         write_offset_data_out_6), .B1 (nx7087)) ;
    nor02ii ix823 (.Y (nx822), .A0 (nx4265), .A1 (write_offset_data_out_4)) ;
    ao22 ix1990 (.Y (nx1989), .A0 (write_offset_data_out_4), .A1 (nx7089), .B0 (
         nx828), .B1 (nx6983)) ;
    or04 ix4266 (.Y (nx4265), .A0 (nx4271), .A1 (nx4277), .A2 (nx7355), .A3 (
         nx4293)) ;
    ao22 ix1970 (.Y (nx1969), .A0 (write_offset_data_out_3), .A1 (nx7089), .B0 (
         nx802), .B1 (nx6983)) ;
    mux21_ni ix1910 (.Y (nx1909), .A0 (nx7089), .A1 (nx6983), .S0 (nx4293)) ;
    or02 ix4296 (.Y (nx4295), .A0 (nx7355), .A1 (nx4293)) ;
    or03 ix4300 (.Y (nx4299), .A0 (nx4277), .A1 (nx7355), .A2 (nx4293)) ;
    mux21_ni ix2220 (.Y (nx2219), .A0 (mem_data_in[15]), .A1 (
             new_size_squared_out_15), .S0 (nx7081)) ;
    xnor2 ix4316 (.Y (nx4314), .A0 (nx4167), .A1 (nx4320)) ;
    mux21_ni ix2200 (.Y (nx2199), .A0 (mem_data_in[14]), .A1 (
             new_size_squared_out_14), .S0 (nx7081)) ;
    xor2 ix4322 (.Y (nx4321), .A0 (nx4305), .A1 (new_size_squared_out_13)) ;
    mux21_ni ix2180 (.Y (nx2179), .A0 (mem_data_in[13]), .A1 (
             new_size_squared_out_13), .S0 (nx7081)) ;
    xnor2 ix4330 (.Y (nx4328), .A0 (nx4183), .A1 (nx4335)) ;
    mux21_ni ix2160 (.Y (nx2159), .A0 (mem_data_in[12]), .A1 (
             new_size_squared_out_12), .S0 (nx7081)) ;
    xor2 ix4338 (.Y (nx4337), .A0 (nx4303), .A1 (new_size_squared_out_11)) ;
    mux21_ni ix2140 (.Y (nx2139), .A0 (mem_data_in[11]), .A1 (
             new_size_squared_out_11), .S0 (nx7081)) ;
    xnor2 ix4344 (.Y (nx4343), .A0 (nx4200), .A1 (nx4349)) ;
    mux21_ni ix2120 (.Y (nx2119), .A0 (mem_data_in[10]), .A1 (
             new_size_squared_out_10), .S0 (nx7081)) ;
    xor2 ix4352 (.Y (nx4351), .A0 (nx4301), .A1 (new_size_squared_out_9)) ;
    mux21_ni ix2100 (.Y (nx2099), .A0 (mem_data_in[9]), .A1 (
             new_size_squared_out_9), .S0 (nx7083)) ;
    xnor2 ix4359 (.Y (nx4358), .A0 (nx4217), .A1 (nx4363)) ;
    mux21_ni ix2080 (.Y (nx2079), .A0 (mem_data_in[8]), .A1 (
             new_size_squared_out_8), .S0 (nx7083)) ;
    xor2 ix4366 (.Y (nx4365), .A0 (nx4229), .A1 (new_size_squared_out_7)) ;
    mux21_ni ix2060 (.Y (nx2059), .A0 (mem_data_in[7]), .A1 (
             new_size_squared_out_7), .S0 (nx7083)) ;
    xnor2 ix4373 (.Y (nx4372), .A0 (nx4239), .A1 (nx4377)) ;
    mux21_ni ix2040 (.Y (nx2039), .A0 (mem_data_in[6]), .A1 (
             new_size_squared_out_6), .S0 (nx7083)) ;
    xor2 ix4380 (.Y (nx4379), .A0 (nx4251), .A1 (new_size_squared_out_5)) ;
    mux21_ni ix2020 (.Y (nx2019), .A0 (mem_data_in[5]), .A1 (
             new_size_squared_out_5), .S0 (nx7083)) ;
    xnor2 ix4387 (.Y (nx4386), .A0 (nx4257), .A1 (nx4391)) ;
    mux21_ni ix2000 (.Y (nx1999), .A0 (mem_data_in[4]), .A1 (
             new_size_squared_out_4), .S0 (nx7083)) ;
    xor2 ix4394 (.Y (nx4393), .A0 (nx4271), .A1 (new_size_squared_out_3)) ;
    mux21_ni ix1980 (.Y (nx1979), .A0 (mem_data_in[3]), .A1 (
             new_size_squared_out_3), .S0 (nx7083)) ;
    xnor2 ix4402 (.Y (nx4400), .A0 (nx4277), .A1 (nx4407)) ;
    mux21_ni ix1960 (.Y (nx1959), .A0 (mem_data_in[2]), .A1 (
             new_size_squared_out_2), .S0 (nx7085)) ;
    xor2 ix4410 (.Y (nx4408), .A0 (nx7355), .A1 (new_size_squared_out_1)) ;
    mux21_ni ix1940 (.Y (nx1939), .A0 (mem_data_in[1]), .A1 (
             new_size_squared_out_1), .S0 (nx7085)) ;
    xnor2 ix4418 (.Y (nx4417), .A0 (nx4293), .A1 (nx4423)) ;
    mux21_ni ix1920 (.Y (nx1919), .A0 (mem_data_in[0]), .A1 (
             new_size_squared_out_0), .S0 (nx7085)) ;
    xnor2 ix1631 (.Y (nx1630), .A0 (nx4447), .A1 (nx4111)) ;
    and02 ix4472 (.Y (nx4471), .A0 (nx4111), .A1 (nx4447)) ;
    and03 ix4500 (.Y (nx4499), .A0 (nx4111), .A1 (nx4447), .A2 (nx4469)) ;
    mux21 ix1769 (.Y (nx1768), .A0 (nx4047), .A1 (nx4526), .S0 (nx3967)) ;
    mux21 ix4534 (.Y (nx4533), .A0 (mem_data_in[0]), .A1 (nx4531), .S0 (nx3967)
          ) ;
    nor02ii ix4536 (.Y (nx4535), .A0 (nlayers_counter_out_1), .A1 (nx4531)) ;
    mux21 ix1785 (.Y (nx1784), .A0 (nx4059), .A1 (nx4543), .S0 (nx3967)) ;
    ao32 ix1447 (.Y (nx1446), .A0 (nx4583), .A1 (current_state_15), .A2 (nx4759)
         , .B0 (current_state_16), .B1 (ftc_cntrl_reg_out_11)) ;
    or02 ix4564 (.Y (nx4563), .A0 (ftc_cntrl_reg_out_14), .A1 (nx7294)) ;
    nor02ii ix4572 (.Y (nx4571), .A0 (nx4), .A1 (nx4879)) ;
    and02 ix5 (.Y (nx4), .A0 (current_state_20), .A1 (nx4705)) ;
    xnor2 ix281 (.Y (nx280), .A0 (nx4647), .A1 (nx278)) ;
    mux21_ni ix1570 (.Y (nx1569), .A0 (nx232), .A1 (cntr1_inst_counter_out_4), .S0 (
             nx7029)) ;
    xor2 ix233 (.Y (nx232), .A0 (nx4647), .A1 (nx4601)) ;
    mux21_ni ix1560 (.Y (nx1559), .A0 (nx214), .A1 (cntr1_inst_counter_out_3), .S0 (
             nx7029)) ;
    mux21_ni ix1550 (.Y (nx1549), .A0 (nx200), .A1 (cntr1_inst_counter_out_2), .S0 (
             nx7029)) ;
    mux21 ix1540 (.Y (nx1539), .A0 (nx4638), .A1 (nx4621), .S0 (nx7029)) ;
    oai21 ix177 (.Y (nx176), .A0 (nx4637), .A1 (nx7021), .B0 (nx6599)) ;
    or02 ix279 (.Y (nx278), .A0 (nx7063), .A1 (nx7031)) ;
    xor2 ix249 (.Y (nx248), .A0 (nx7295), .A1 (cntr1_inst_counter_out_2)) ;
    xnor2 ix247 (.Y (nx246), .A0 (nx7295), .A1 (nx4655)) ;
    mux21 ix1580 (.Y (nx1579), .A0 (nx4657), .A1 (nx4655), .S0 (nx7295)) ;
    xor2 ix4658 (.Y (nx4657), .A0 (nx4655), .A1 (nx1425)) ;
    nor02ii ix239 (.Y (nx1425), .A0 (nx4601), .A1 (cntr1_inst_counter_out_4)) ;
    xnor2 ix4664 (.Y (nx4663), .A0 (nx7295), .A1 (cntr1_inst_counter_out_1)) ;
    nor02ii ix4674 (.Y (nx4673), .A0 (nx1469), .A1 (nx4725)) ;
    and02 ix1851 (.Y (nx1469), .A0 (current_state_20), .A1 (nx4705)) ;
    and04 ix1371 (.Y (nx1370), .A0 (nx5148), .A1 (nx4692), .A2 (nx5146), .A3 (
          nx5023)) ;
    mux21 ix2400 (.Y (nx2399), .A0 (nx5148), .A1 (nx4689), .S0 (nx7101)) ;
    xor2 ix4690 (.Y (nx4689), .A0 (nx5148), .A1 (nx1447)) ;
    nor02ii ix1351 (.Y (nx1447), .A0 (nx5013), .A1 (
            cache_width_cntr_counter_out_14)) ;
    mux21_ni ix2390 (.Y (nx2389), .A0 (cache_width_cntr_counter_out_14), .A1 (
             nx1344), .S0 (nx7101)) ;
    xor2 ix1345 (.Y (nx1344), .A0 (nx4692), .A1 (nx5013)) ;
    nor02ii ix319 (.Y (nx1427), .A0 (nx7033), .A1 (nx4723)) ;
    and04 ix4718 (.Y (nx4717), .A0 (nx5113), .A1 (nx4725), .A2 (nx4765), .A3 (
          nx4879)) ;
    or02 ix547 (.Y (nx546), .A0 (ftc_cntrl_reg_out_11), .A1 (nx4765)) ;
    and04 ix521 (.Y (nx520), .A0 (nx4743), .A1 (nx4770), .A2 (nx4781), .A3 (
          nx4787)) ;
    mux21 ix1780 (.Y (nx1779), .A0 (nx4767), .A1 (nx4743), .S0 (nx7037)) ;
    or03 ix4752 (.Y (nx4751), .A0 (ftc_cntrl_reg_out_8), .A1 (nx4725), .A2 (
         nx4759)) ;
    ao21 ix1117 (.Y (nx1116), .A0 (nx7033), .A1 (nx4575), .B0 (current_state_16)
         ) ;
    xor2 ix4768 (.Y (nx4767), .A0 (nx4743), .A1 (nx1430)) ;
    nor02ii ix501 (.Y (nx1430), .A0 (nx4776), .A1 (
            window_width_cntr_counter_out_14)) ;
    mux21_ni ix1770 (.Y (nx1769), .A0 (nx494), .A1 (
             window_width_cntr_counter_out_14), .S0 (nx7037)) ;
    xor2 ix495 (.Y (nx494), .A0 (nx4770), .A1 (nx4776)) ;
    mux21 ix1760 (.Y (nx1759), .A0 (nx4783), .A1 (nx4781), .S0 (nx7037)) ;
    nor02ii ix477 (.Y (nx1432), .A0 (nx4795), .A1 (
            window_width_cntr_counter_out_12)) ;
    mux21_ni ix1750 (.Y (nx1749), .A0 (nx470), .A1 (
             window_width_cntr_counter_out_12), .S0 (nx7037)) ;
    xor2 ix471 (.Y (nx470), .A0 (nx4787), .A1 (nx4795)) ;
    mux21 ix1740 (.Y (nx1739), .A0 (nx4803), .A1 (nx4801), .S0 (nx7037)) ;
    nor02ii ix453 (.Y (nx1434), .A0 (nx4813), .A1 (
            window_width_cntr_counter_out_10)) ;
    mux21_ni ix1730 (.Y (nx1729), .A0 (nx446), .A1 (
             window_width_cntr_counter_out_10), .S0 (nx7037)) ;
    xor2 ix447 (.Y (nx446), .A0 (nx4807), .A1 (nx4813)) ;
    mux21 ix1720 (.Y (nx1719), .A0 (nx4821), .A1 (nx4819), .S0 (nx7037)) ;
    nor02ii ix429 (.Y (nx1436), .A0 (nx4833), .A1 (
            window_width_cntr_counter_out_8)) ;
    mux21_ni ix1710 (.Y (nx1709), .A0 (nx422), .A1 (
             window_width_cntr_counter_out_8), .S0 (nx7039)) ;
    xor2 ix423 (.Y (nx422), .A0 (nx4825), .A1 (nx4833)) ;
    mux21 ix1700 (.Y (nx1699), .A0 (nx4841), .A1 (nx4839), .S0 (nx7039)) ;
    nor02ii ix405 (.Y (nx1439), .A0 (nx4853), .A1 (
            window_width_cntr_counter_out_6)) ;
    mux21_ni ix1690 (.Y (nx1689), .A0 (nx398), .A1 (
             window_width_cntr_counter_out_6), .S0 (nx7039)) ;
    xor2 ix399 (.Y (nx398), .A0 (nx4845), .A1 (nx4853)) ;
    or03 ix4854 (.Y (nx4853), .A0 (nx6943), .A1 (nx4911), .A2 (nx4861)) ;
    inv01 ix6942 (.Y (nx6943), .A (wind_width_count_4)) ;
    mux21_ni ix2600 (.Y (nx2599), .A0 (nx1880), .A1 (wind_width_count_4), .S0 (
             nx7039)) ;
    mux21_ni ix1650 (.Y (nx1649), .A0 (nx354), .A1 (wind_width_count_1), .S0 (
             nx7039)) ;
    xor2 ix1640 (.Y (nx1639), .A0 (nx6607), .A1 (nx1429)) ;
    mux21_ni ix1660 (.Y (nx1659), .A0 (nx362), .A1 (wind_width_count_2), .S0 (
             nx7039)) ;
    mux21_ni ix1670 (.Y (nx1669), .A0 (nx370), .A1 (wind_width_count_3), .S0 (
             nx7039)) ;
    mux21 ix1680 (.Y (nx1679), .A0 (nx4913), .A1 (nx4911), .S0 (nx7041)) ;
    and04 ix535 (.Y (nx534), .A0 (nx4801), .A1 (nx4807), .A2 (nx4819), .A3 (
          nx4825)) ;
    and04 ix583 (.Y (nx582), .A0 (nx4839), .A1 (nx4845), .A2 (nx4911), .A3 (
          nx6945)) ;
    inv01 ix6944 (.Y (nx6945), .A (nx574)) ;
    mux21 ix573 (.Y (nx572), .A0 (nx7063), .A1 (img_width_out_0), .S0 (nx6977)
          ) ;
    ao221 ix1800 (.Y (nx1799), .A0 (img_width_out_0), .A1 (nx4119), .B0 (nx6665)
          , .B1 (new_width_out_0), .C0 (current_state_9)) ;
    mux21 ix611 (.Y (nx610), .A0 (nx7065), .A1 (nx5155), .S0 (nx6977)) ;
    nor02ii ix675 (.Y (nx674), .A0 (nx4981), .A1 (nx6977)) ;
    nor02ii ix693 (.Y (nx692), .A0 (nx4997), .A1 (nx6979)) ;
    or02 ix5012 (.Y (nx5011), .A0 (nx4575), .A1 (nx4705)) ;
    mux21 ix2380 (.Y (nx2379), .A0 (nx5146), .A1 (nx5019), .S0 (nx7101)) ;
    nor02ii ix1327 (.Y (nx1449), .A0 (nx5031), .A1 (
            cache_width_cntr_counter_out_12)) ;
    mux21_ni ix2370 (.Y (nx2369), .A0 (cache_width_cntr_counter_out_12), .A1 (
             nx1320), .S0 (nx7101)) ;
    xor2 ix1321 (.Y (nx1320), .A0 (nx5023), .A1 (nx5031)) ;
    mux21 ix2360 (.Y (nx2359), .A0 (nx5144), .A1 (nx5037), .S0 (nx7101)) ;
    nor02ii ix1303 (.Y (nx1451), .A0 (nx5049), .A1 (
            cache_width_cntr_counter_out_10)) ;
    mux21_ni ix2350 (.Y (nx2349), .A0 (cache_width_cntr_counter_out_10), .A1 (
             nx1296), .S0 (nx7101)) ;
    xor2 ix1297 (.Y (nx1296), .A0 (nx5041), .A1 (nx5049)) ;
    mux21 ix2340 (.Y (nx2339), .A0 (nx5142), .A1 (nx5055), .S0 (nx7101)) ;
    nor02ii ix1279 (.Y (nx1454), .A0 (nx5067), .A1 (
            cache_width_cntr_counter_out_8)) ;
    mux21_ni ix2330 (.Y (nx2329), .A0 (cache_width_cntr_counter_out_8), .A1 (
             nx1272), .S0 (nx7103)) ;
    xor2 ix1273 (.Y (nx1272), .A0 (nx5059), .A1 (nx5067)) ;
    mux21 ix2320 (.Y (nx2319), .A0 (nx5140), .A1 (nx5072), .S0 (nx7103)) ;
    nor02ii ix1255 (.Y (nx1456), .A0 (nx5083), .A1 (
            cache_width_cntr_counter_out_6)) ;
    mux21_ni ix2310 (.Y (nx2309), .A0 (cache_width_cntr_counter_out_6), .A1 (
             nx1248), .S0 (nx7103)) ;
    xor2 ix1249 (.Y (nx1248), .A0 (nx5077), .A1 (nx5083)) ;
    or03 ix5084 (.Y (nx5083), .A0 (nx6947), .A1 (nx5137), .A2 (nx5089)) ;
    inv01 ix6946 (.Y (nx6947), .A (nx6613)) ;
    mux21_ni ix2290 (.Y (nx2289), .A0 (nx6611), .A1 (nx1222), .S0 (nx7103)) ;
    mux21_ni ix2260 (.Y (nx2259), .A0 (cache_width_count_1), .A1 (nx1198), .S0 (
             nx7103)) ;
    xor2 ix2250 (.Y (nx2249), .A0 (cache_width_count_0), .A1 (nx7103)) ;
    and02 ix5114 (.Y (nx5113), .A0 (nx7033), .A1 (nx4575)) ;
    mux21_ni ix2270 (.Y (nx2269), .A0 (nx6615), .A1 (nx1206), .S0 (nx7103)) ;
    mux21_ni ix2280 (.Y (nx2279), .A0 (cache_width_count_3), .A1 (nx1214), .S0 (
             nx7105)) ;
    mux21 ix2300 (.Y (nx2299), .A0 (nx5137), .A1 (nx5134), .S0 (nx7105)) ;
    and04 ix1385 (.Y (nx1384), .A0 (nx5144), .A1 (nx5041), .A2 (nx5142), .A3 (
          nx5059)) ;
    and04 ix1403 (.Y (nx1402), .A0 (nx5140), .A1 (nx5077), .A2 (nx5137), .A3 (
          nx6949)) ;
    xnor2 ix1395 (.Y (nx6949), .A0 (nx4927), .A1 (cache_width_count_0)) ;
    xor2 ix1405 (.Y (nx1404), .A0 (cache_width_count_1), .A1 (nx606)) ;
    nor02ii ix5158 (.Y (nx5157), .A0 (img_width_out_1), .A1 (nx4927)) ;
    nor02_2x ix1453 (.Y (nx1452), .A0 (nx7023), .A1 (nx7065)) ;
    and02 ix1871 (.Y (nx1459), .A0 (current_state_21), .A1 (nx4731)) ;
    mux21 ix2610 (.Y (nx2609), .A0 (current_state_27), .A1 (nx7043), .S0 (nx5194
          )) ;
    mux21 ix2620 (.Y (nx2619), .A0 (nx5204), .A1 (nx5202), .S0 (nx7043)) ;
    or02 ix5207 (.Y (nx5206), .A0 (nx5202), .A1 (nx5194)) ;
    mux21_ni ix2630 (.Y (nx2629), .A0 (nx1908), .A1 (class_cntr_counter_out_2), 
             .S0 (nx7043)) ;
    xor2 ix1909 (.Y (nx1908), .A0 (nx5208), .A1 (nx5206)) ;
    mux21_ni ix2640 (.Y (nx2639), .A0 (nx1916), .A1 (class_cntr_counter_out_3), 
             .S0 (nx5191)) ;
    xor2 ix1917 (.Y (nx1916), .A0 (nx5218), .A1 (nx5216)) ;
    or03 ix5217 (.Y (nx5216), .A0 (nx5208), .A1 (nx5202), .A2 (nx5194)) ;
    nor02ii ix4847 (.Y (argmax_data_out[0]), .A0 (argmax_ready_dup0), .A1 (
            mem_data_in[0])) ;
    nor02ii ix4849 (.Y (argmax_data_out[1]), .A0 (nx7325), .A1 (mem_data_in[1])
            ) ;
    nor02ii ix4851 (.Y (argmax_data_out[2]), .A0 (nx7326), .A1 (mem_data_in[2])
            ) ;
    nor02ii ix4855 (.Y (argmax_data_out[4]), .A0 (nx7327), .A1 (mem_data_in[4])
            ) ;
    nor02ii ix4857 (.Y (argmax_data_out[5]), .A0 (nx7328), .A1 (mem_data_in[5])
            ) ;
    nor02ii ix4861 (.Y (argmax_data_out[7]), .A0 (nx7047), .A1 (mem_data_in[7])
            ) ;
    nor02ii ix4863 (.Y (argmax_data_out[8]), .A0 (nx7047), .A1 (mem_data_in[8])
            ) ;
    nor02ii ix4865 (.Y (argmax_data_out[9]), .A0 (nx7047), .A1 (mem_data_in[9])
            ) ;
    nor02ii ix4867 (.Y (argmax_data_out[10]), .A0 (nx7047), .A1 (mem_data_in[10]
            )) ;
    nor02ii ix4869 (.Y (argmax_data_out[11]), .A0 (nx7047), .A1 (mem_data_in[11]
            )) ;
    nor02ii ix4871 (.Y (argmax_data_out[12]), .A0 (nx7047), .A1 (mem_data_in[12]
            )) ;
    nor02ii ix4873 (.Y (argmax_data_out[13]), .A0 (nx7049), .A1 (mem_data_in[13]
            )) ;
    nor02ii ix4875 (.Y (argmax_data_out[14]), .A0 (nx7049), .A1 (mem_data_in[14]
            )) ;
    nor02ii ix4877 (.Y (argmax_data_out[15]), .A0 (nx7049), .A1 (mem_data_in[15]
            )) ;
    and02 ix4879 (.Y (comp_unit_data2_out[0]), .A0 (nx6985), .A1 (nx2096)) ;
    mux21_ni ix2097 (.Y (nx2096), .A0 (flt_bias_out_0), .A1 (mem_data_in[0]), .S0 (
             nx7053)) ;
    nor02ii ix2085 (.Y (nx2084), .A0 (nx6927), .A1 (current_state_12)) ;
    and02 ix4881 (.Y (comp_unit_data2_out[1]), .A0 (nx6987), .A1 (nx2124)) ;
    mux21_ni ix2125 (.Y (nx2124), .A0 (flt_bias_out_1), .A1 (mem_data_in[1]), .S0 (
             nx7053)) ;
    and02 ix4883 (.Y (comp_unit_data2_out[2]), .A0 (nx6987), .A1 (nx2150)) ;
    mux21_ni ix2151 (.Y (nx2150), .A0 (flt_bias_out_2), .A1 (mem_data_in[2]), .S0 (
             nx7053)) ;
    and02 ix4885 (.Y (comp_unit_data2_out[3]), .A0 (nx6987), .A1 (nx2176)) ;
    mux21_ni ix2177 (.Y (nx2176), .A0 (flt_bias_out_3), .A1 (mem_data_in[3]), .S0 (
             nx7053)) ;
    and02 ix4887 (.Y (comp_unit_data2_out[4]), .A0 (nx6987), .A1 (nx2202)) ;
    mux21_ni ix2203 (.Y (nx2202), .A0 (flt_bias_out_4), .A1 (mem_data_in[4]), .S0 (
             nx7053)) ;
    and02 ix4889 (.Y (comp_unit_data2_out[5]), .A0 (nx6987), .A1 (nx2228)) ;
    mux21_ni ix2229 (.Y (nx2228), .A0 (flt_bias_out_5), .A1 (mem_data_in[5]), .S0 (
             nx7055)) ;
    and02 ix4891 (.Y (comp_unit_data2_out[6]), .A0 (nx6987), .A1 (nx2254)) ;
    mux21_ni ix2255 (.Y (nx2254), .A0 (flt_bias_out_6), .A1 (mem_data_in[6]), .S0 (
             nx7055)) ;
    and02 ix4893 (.Y (comp_unit_data2_out[7]), .A0 (nx6987), .A1 (nx2280)) ;
    mux21_ni ix2281 (.Y (nx2280), .A0 (flt_bias_out_7), .A1 (mem_data_in[7]), .S0 (
             nx7055)) ;
    and02 ix4895 (.Y (comp_unit_data2_out[8]), .A0 (nx6989), .A1 (nx2306)) ;
    mux21_ni ix2307 (.Y (nx2306), .A0 (flt_bias_out_8), .A1 (mem_data_in[8]), .S0 (
             nx7055)) ;
    and02 ix4897 (.Y (comp_unit_data2_out[9]), .A0 (nx6989), .A1 (nx2332)) ;
    mux21_ni ix2333 (.Y (nx2332), .A0 (flt_bias_out_9), .A1 (mem_data_in[9]), .S0 (
             nx7055)) ;
    and02 ix4899 (.Y (comp_unit_data2_out[10]), .A0 (nx6989), .A1 (nx2358)) ;
    mux21_ni ix2359 (.Y (nx2358), .A0 (flt_bias_out_10), .A1 (mem_data_in[10]), 
             .S0 (nx7055)) ;
    and02 ix4901 (.Y (comp_unit_data2_out[11]), .A0 (nx6989), .A1 (nx2384)) ;
    mux21_ni ix2385 (.Y (nx2384), .A0 (flt_bias_out_11), .A1 (mem_data_in[11]), 
             .S0 (nx7055)) ;
    and02 ix4903 (.Y (comp_unit_data2_out[12]), .A0 (nx6989), .A1 (nx2410)) ;
    mux21_ni ix2411 (.Y (nx2410), .A0 (flt_bias_out_12), .A1 (mem_data_in[12]), 
             .S0 (nx7057)) ;
    and02 ix4905 (.Y (comp_unit_data2_out[13]), .A0 (nx6989), .A1 (nx2436)) ;
    mux21_ni ix2437 (.Y (nx2436), .A0 (flt_bias_out_13), .A1 (mem_data_in[13]), 
             .S0 (nx7057)) ;
    and02 ix4907 (.Y (comp_unit_data2_out[14]), .A0 (nx6989), .A1 (nx2462)) ;
    mux21_ni ix2463 (.Y (nx2462), .A0 (flt_bias_out_14), .A1 (mem_data_in[14]), 
             .S0 (nx7057)) ;
    and02 ix4909 (.Y (comp_unit_data2_out[15]), .A0 (nx6991), .A1 (nx2488)) ;
    mux21_ni ix2489 (.Y (nx2488), .A0 (flt_bias_out_15), .A1 (mem_data_in[15]), 
             .S0 (nx7057)) ;
    and03 ix5077 (.Y (max_height_1), .A0 (nx606), .A1 (nx6599), .A2 (nx7035)) ;
    nor04 ix5111 (.Y (comp_unit_relu), .A0 (nx6951), .A1 (nx4111), .A2 (
          num_channels_out_2), .A3 (num_channels_out_1)) ;
    nand04 ix5101 (.Y (nx6951), .A0 (nx4004), .A1 (nx6953), .A2 (nx4503), .A3 (
           nx4497)) ;
    inv01 ix6952 (.Y (nx6953), .A (nx6927)) ;
    oai21 ix2573 (.Y (cache_load), .A0 (nx7065), .A1 (nx6955), .B0 (nx7107)) ;
    inv01 ix6954 (.Y (nx6955), .A (nx4)) ;
    or03 ix2523 (.Y (nx2522), .A0 (nx4723), .A1 (current_state_20), .A2 (nx7035)
         ) ;
    and02 ix2539 (.Y (cache_data_in_0), .A0 (mem_data_in[0]), .A1 (nx6999)) ;
    ao21 ix5340 (.Y (nx2536), .A0 (nx5334), .A1 (nx1469), .B0 (nx1152)) ;
    and02 ix2541 (.Y (cache_data_in_1), .A0 (mem_data_in[1]), .A1 (nx6999)) ;
    and02 ix2543 (.Y (cache_data_in_2), .A0 (mem_data_in[2]), .A1 (nx6999)) ;
    and02 ix2545 (.Y (cache_data_in_3), .A0 (mem_data_in[3]), .A1 (nx6999)) ;
    and02 ix2547 (.Y (cache_data_in_4), .A0 (mem_data_in[4]), .A1 (nx6999)) ;
    and02 ix2549 (.Y (cache_data_in_5), .A0 (mem_data_in[5]), .A1 (nx6999)) ;
    and02 ix2551 (.Y (cache_data_in_6), .A0 (mem_data_in[6]), .A1 (nx6999)) ;
    and02 ix2553 (.Y (cache_data_in_7), .A0 (mem_data_in[7]), .A1 (nx7001)) ;
    and02 ix2555 (.Y (cache_data_in_8), .A0 (mem_data_in[8]), .A1 (nx7001)) ;
    and02 ix2557 (.Y (cache_data_in_9), .A0 (mem_data_in[9]), .A1 (nx7001)) ;
    and02 ix2559 (.Y (cache_data_in_10), .A0 (mem_data_in[10]), .A1 (nx7001)) ;
    and02 ix2561 (.Y (cache_data_in_11), .A0 (mem_data_in[11]), .A1 (nx7001)) ;
    and02 ix2563 (.Y (cache_data_in_12), .A0 (mem_data_in[12]), .A1 (nx7001)) ;
    and02 ix2565 (.Y (cache_data_in_13), .A0 (mem_data_in[13]), .A1 (nx7001)) ;
    and02 ix2567 (.Y (cache_data_in_14), .A0 (mem_data_in[14]), .A1 (nx7003)) ;
    and02 ix2569 (.Y (cache_data_in_15), .A0 (mem_data_in[15]), .A1 (nx7003)) ;
    and02 ix5380 (.Y (nx5379), .A0 (nx6599), .A1 (nx7035)) ;
    mux21 ix2670 (.Y (nx2669), .A0 (nx5386), .A1 (nx5383), .S0 (nx7023)) ;
    mux21 ix2690 (.Y (nx2689), .A0 (nx5393), .A1 (nx5390), .S0 (nx7023)) ;
    mux21 ix2710 (.Y (nx2709), .A0 (nx5399), .A1 (nx5396), .S0 (nx7023)) ;
    mux21 ix2730 (.Y (nx2729), .A0 (nx5405), .A1 (nx5402), .S0 (nx7023)) ;
    mux21 ix2750 (.Y (nx2749), .A0 (nx5411), .A1 (nx5408), .S0 (nx7025)) ;
    mux21 ix2770 (.Y (nx2769), .A0 (nx5417), .A1 (nx5414), .S0 (nx7025)) ;
    mux21 ix2790 (.Y (nx2789), .A0 (nx5423), .A1 (nx5420), .S0 (nx7025)) ;
    mux21 ix2810 (.Y (nx2809), .A0 (nx5429), .A1 (nx5426), .S0 (nx7025)) ;
    mux21 ix2830 (.Y (nx2829), .A0 (nx5435), .A1 (nx5432), .S0 (nx7025)) ;
    mux21 ix2850 (.Y (nx2849), .A0 (nx5441), .A1 (nx5438), .S0 (nx7025)) ;
    mux21 ix2870 (.Y (nx2869), .A0 (nx5447), .A1 (nx5444), .S0 (nx7025)) ;
    mux21 ix2890 (.Y (nx2889), .A0 (nx5453), .A1 (nx5450), .S0 (nx7027)) ;
    mux21 ix2910 (.Y (nx2909), .A0 (nx5459), .A1 (nx5456), .S0 (nx7027)) ;
    mux21 ix2930 (.Y (nx2929), .A0 (nx5465), .A1 (nx5462), .S0 (nx7027)) ;
    mux21 ix2950 (.Y (nx2949), .A0 (nx5471), .A1 (nx5468), .S0 (nx7027)) ;
    mux21 ix2970 (.Y (nx2969), .A0 (nx5477), .A1 (nx5474), .S0 (nx7027)) ;
    nor02ii ix4815 (.Y (filter_data_out[0]), .A0 (nx7077), .A1 (mem_data_in[0])
            ) ;
    nor02ii ix4817 (.Y (filter_data_out[1]), .A0 (nx7077), .A1 (mem_data_in[1])
            ) ;
    nor02ii ix4819 (.Y (filter_data_out[2]), .A0 (nx7077), .A1 (mem_data_in[2])
            ) ;
    nor02ii ix4821 (.Y (filter_data_out[3]), .A0 (nx7077), .A1 (mem_data_in[3])
            ) ;
    nor02ii ix4823 (.Y (filter_data_out[4]), .A0 (nx7077), .A1 (mem_data_in[4])
            ) ;
    nor02ii ix4825 (.Y (filter_data_out[5]), .A0 (nx7079), .A1 (mem_data_in[5])
            ) ;
    nor02ii ix4827 (.Y (filter_data_out[6]), .A0 (nx7079), .A1 (mem_data_in[6])
            ) ;
    nor02ii ix4829 (.Y (filter_data_out[7]), .A0 (nx7079), .A1 (mem_data_in[7])
            ) ;
    nor02ii ix4831 (.Y (filter_data_out[8]), .A0 (nx7079), .A1 (mem_data_in[8])
            ) ;
    nor02ii ix4833 (.Y (filter_data_out[9]), .A0 (nx7079), .A1 (mem_data_in[9])
            ) ;
    nor02ii ix4835 (.Y (filter_data_out[10]), .A0 (nx7079), .A1 (mem_data_in[10]
            )) ;
    nor02ii ix4837 (.Y (filter_data_out[11]), .A0 (nx7079), .A1 (mem_data_in[11]
            )) ;
    nor02ii ix4839 (.Y (filter_data_out[12]), .A0 (nx6657), .A1 (mem_data_in[12]
            )) ;
    nor02ii ix4841 (.Y (filter_data_out[13]), .A0 (nx6657), .A1 (mem_data_in[13]
            )) ;
    nor02ii ix4843 (.Y (filter_data_out[14]), .A0 (nx6657), .A1 (mem_data_in[14]
            )) ;
    nor02ii ix4845 (.Y (filter_data_out[15]), .A0 (nx6657), .A1 (mem_data_in[15]
            )) ;
    and02 ix4911 (.Y (wind_col_in_0__0), .A0 (nx7123), .A1 (cache_data_out_0__0)
          ) ;
    and02 ix4913 (.Y (wind_col_in_0__1), .A0 (nx7123), .A1 (cache_data_out_0__1)
          ) ;
    and02 ix4915 (.Y (wind_col_in_0__2), .A0 (nx7123), .A1 (cache_data_out_0__2)
          ) ;
    and02 ix4917 (.Y (wind_col_in_0__3), .A0 (nx7123), .A1 (cache_data_out_0__3)
          ) ;
    and02 ix4919 (.Y (wind_col_in_0__4), .A0 (nx7123), .A1 (cache_data_out_0__4)
          ) ;
    and02 ix4921 (.Y (wind_col_in_0__5), .A0 (nx7123), .A1 (cache_data_out_0__5)
          ) ;
    and02 ix4923 (.Y (wind_col_in_0__6), .A0 (nx7123), .A1 (cache_data_out_0__6)
          ) ;
    and02 ix4925 (.Y (wind_col_in_0__7), .A0 (nx7125), .A1 (cache_data_out_0__7)
          ) ;
    and02 ix4927 (.Y (wind_col_in_0__8), .A0 (nx7125), .A1 (cache_data_out_0__8)
          ) ;
    and02 ix4929 (.Y (wind_col_in_0__9), .A0 (nx7125), .A1 (cache_data_out_0__9)
          ) ;
    and02 ix4931 (.Y (wind_col_in_0__10), .A0 (nx7125), .A1 (
          cache_data_out_0__10)) ;
    and02 ix4933 (.Y (wind_col_in_0__11), .A0 (nx7125), .A1 (
          cache_data_out_0__11)) ;
    and02 ix4935 (.Y (wind_col_in_0__12), .A0 (nx7125), .A1 (
          cache_data_out_0__12)) ;
    and02 ix4937 (.Y (wind_col_in_0__13), .A0 (nx7125), .A1 (
          cache_data_out_0__13)) ;
    and02 ix4939 (.Y (wind_col_in_0__14), .A0 (nx7127), .A1 (
          cache_data_out_0__14)) ;
    and02 ix4941 (.Y (wind_col_in_0__15), .A0 (nx7127), .A1 (
          cache_data_out_0__15)) ;
    and02 ix4943 (.Y (wind_col_in_1__0), .A0 (nx7127), .A1 (cache_data_out_1__0)
          ) ;
    and02 ix4945 (.Y (wind_col_in_1__1), .A0 (nx7127), .A1 (cache_data_out_1__1)
          ) ;
    and02 ix4947 (.Y (wind_col_in_1__2), .A0 (nx7127), .A1 (cache_data_out_1__2)
          ) ;
    and02 ix4949 (.Y (wind_col_in_1__3), .A0 (nx7127), .A1 (cache_data_out_1__3)
          ) ;
    and02 ix4951 (.Y (wind_col_in_1__4), .A0 (nx7127), .A1 (cache_data_out_1__4)
          ) ;
    and02 ix4953 (.Y (wind_col_in_1__5), .A0 (nx7129), .A1 (cache_data_out_1__5)
          ) ;
    and02 ix4955 (.Y (wind_col_in_1__6), .A0 (nx7129), .A1 (cache_data_out_1__6)
          ) ;
    and02 ix4957 (.Y (wind_col_in_1__7), .A0 (nx7129), .A1 (cache_data_out_1__7)
          ) ;
    and02 ix4959 (.Y (wind_col_in_1__8), .A0 (nx7129), .A1 (cache_data_out_1__8)
          ) ;
    and02 ix4961 (.Y (wind_col_in_1__9), .A0 (nx7129), .A1 (cache_data_out_1__9)
          ) ;
    and02 ix4963 (.Y (wind_col_in_1__10), .A0 (nx7129), .A1 (
          cache_data_out_1__10)) ;
    and02 ix4965 (.Y (wind_col_in_1__11), .A0 (nx7129), .A1 (
          cache_data_out_1__11)) ;
    and02 ix4967 (.Y (wind_col_in_1__12), .A0 (nx7131), .A1 (
          cache_data_out_1__12)) ;
    and02 ix4969 (.Y (wind_col_in_1__13), .A0 (nx7131), .A1 (
          cache_data_out_1__13)) ;
    and02 ix4971 (.Y (wind_col_in_1__14), .A0 (nx7131), .A1 (
          cache_data_out_1__14)) ;
    and02 ix4973 (.Y (wind_col_in_1__15), .A0 (nx7131), .A1 (
          cache_data_out_1__15)) ;
    and02 ix4975 (.Y (wind_col_in_2__0), .A0 (nx7131), .A1 (cache_data_out_2__0)
          ) ;
    and02 ix4977 (.Y (wind_col_in_2__1), .A0 (nx7131), .A1 (cache_data_out_2__1)
          ) ;
    and02 ix4979 (.Y (wind_col_in_2__2), .A0 (nx7131), .A1 (cache_data_out_2__2)
          ) ;
    and02 ix4981 (.Y (wind_col_in_2__3), .A0 (nx6931), .A1 (cache_data_out_2__3)
          ) ;
    and02 ix4983 (.Y (wind_col_in_2__4), .A0 (nx6931), .A1 (cache_data_out_2__4)
          ) ;
    and02 ix4985 (.Y (wind_col_in_2__5), .A0 (nx6931), .A1 (cache_data_out_2__5)
          ) ;
    and02 ix4987 (.Y (wind_col_in_2__6), .A0 (nx6931), .A1 (cache_data_out_2__6)
          ) ;
    and02 ix4989 (.Y (wind_col_in_2__7), .A0 (nx6931), .A1 (cache_data_out_2__7)
          ) ;
    and02 ix4991 (.Y (wind_col_in_2__8), .A0 (nx6931), .A1 (cache_data_out_2__8)
          ) ;
    and02 ix4993 (.Y (wind_col_in_2__9), .A0 (nx6931), .A1 (cache_data_out_2__9)
          ) ;
    and02 ix4995 (.Y (wind_col_in_2__10), .A0 (nx7133), .A1 (
          cache_data_out_2__10)) ;
    and02 ix4997 (.Y (wind_col_in_2__11), .A0 (nx7133), .A1 (
          cache_data_out_2__11)) ;
    and02 ix4999 (.Y (wind_col_in_2__12), .A0 (nx7133), .A1 (
          cache_data_out_2__12)) ;
    and02 ix5001 (.Y (wind_col_in_2__13), .A0 (nx7133), .A1 (
          cache_data_out_2__13)) ;
    and02 ix5003 (.Y (wind_col_in_2__14), .A0 (nx7133), .A1 (
          cache_data_out_2__14)) ;
    and02 ix5005 (.Y (wind_col_in_2__15), .A0 (nx7133), .A1 (
          cache_data_out_2__15)) ;
    and02 ix5007 (.Y (wind_col_in_3__0), .A0 (nx7133), .A1 (cache_data_out_3__0)
          ) ;
    and02 ix5009 (.Y (wind_col_in_3__1), .A0 (nx7135), .A1 (cache_data_out_3__1)
          ) ;
    and02 ix5011 (.Y (wind_col_in_3__2), .A0 (nx7135), .A1 (cache_data_out_3__2)
          ) ;
    and02 ix5013 (.Y (wind_col_in_3__3), .A0 (nx7135), .A1 (cache_data_out_3__3)
          ) ;
    and02 ix5015 (.Y (wind_col_in_3__4), .A0 (nx7135), .A1 (cache_data_out_3__4)
          ) ;
    and02 ix5017 (.Y (wind_col_in_3__5), .A0 (nx7135), .A1 (cache_data_out_3__5)
          ) ;
    and02 ix5019 (.Y (wind_col_in_3__6), .A0 (nx7135), .A1 (cache_data_out_3__6)
          ) ;
    and02 ix5021 (.Y (wind_col_in_3__7), .A0 (nx7135), .A1 (cache_data_out_3__7)
          ) ;
    and02 ix5023 (.Y (wind_col_in_3__8), .A0 (nx7137), .A1 (cache_data_out_3__8)
          ) ;
    and02 ix5025 (.Y (wind_col_in_3__9), .A0 (nx7137), .A1 (cache_data_out_3__9)
          ) ;
    and02 ix5027 (.Y (wind_col_in_3__10), .A0 (nx7137), .A1 (
          cache_data_out_3__10)) ;
    and02 ix5029 (.Y (wind_col_in_3__11), .A0 (nx7137), .A1 (
          cache_data_out_3__11)) ;
    and02 ix5031 (.Y (wind_col_in_3__12), .A0 (nx7137), .A1 (
          cache_data_out_3__12)) ;
    and02 ix5033 (.Y (wind_col_in_3__13), .A0 (nx7137), .A1 (
          cache_data_out_3__13)) ;
    and02 ix5035 (.Y (wind_col_in_3__14), .A0 (nx7137), .A1 (
          cache_data_out_3__14)) ;
    and02 ix5037 (.Y (wind_col_in_3__15), .A0 (nx7139), .A1 (
          cache_data_out_3__15)) ;
    and02 ix5039 (.Y (wind_col_in_4__0), .A0 (nx7139), .A1 (cache_data_out_4__0)
          ) ;
    and02 ix5041 (.Y (wind_col_in_4__1), .A0 (nx7139), .A1 (cache_data_out_4__1)
          ) ;
    and02 ix5043 (.Y (wind_col_in_4__2), .A0 (nx7139), .A1 (cache_data_out_4__2)
          ) ;
    and02 ix5045 (.Y (wind_col_in_4__3), .A0 (nx7139), .A1 (cache_data_out_4__3)
          ) ;
    and02 ix5047 (.Y (wind_col_in_4__4), .A0 (nx7139), .A1 (cache_data_out_4__4)
          ) ;
    and02 ix5049 (.Y (wind_col_in_4__5), .A0 (nx7139), .A1 (cache_data_out_4__5)
          ) ;
    and02 ix5051 (.Y (wind_col_in_4__6), .A0 (nx6933), .A1 (cache_data_out_4__6)
          ) ;
    and02 ix5053 (.Y (wind_col_in_4__7), .A0 (nx6933), .A1 (cache_data_out_4__7)
          ) ;
    and02 ix5055 (.Y (wind_col_in_4__8), .A0 (nx6933), .A1 (cache_data_out_4__8)
          ) ;
    and02 ix5057 (.Y (wind_col_in_4__9), .A0 (nx6933), .A1 (cache_data_out_4__9)
          ) ;
    and02 ix5059 (.Y (wind_col_in_4__10), .A0 (nx6933), .A1 (
          cache_data_out_4__10)) ;
    and02 ix5061 (.Y (wind_col_in_4__11), .A0 (nx6933), .A1 (
          cache_data_out_4__11)) ;
    and02 ix5063 (.Y (wind_col_in_4__12), .A0 (nx6933), .A1 (
          cache_data_out_4__12)) ;
    and02 ix5065 (.Y (wind_col_in_4__13), .A0 (nx2502), .A1 (
          cache_data_out_4__13)) ;
    and02 ix5067 (.Y (wind_col_in_4__14), .A0 (nx2502), .A1 (
          cache_data_out_4__14)) ;
    and02 ix5069 (.Y (wind_col_in_4__15), .A0 (nx2502), .A1 (
          cache_data_out_4__15)) ;
    or03 ix2511 (.Y (wind_en), .A0 (nx4883), .A1 (nx7145), .A2 (nx1459)) ;
    or03 ix2503 (.Y (nx2502), .A0 (nx4731), .A1 (nx4879), .A2 (nx7065)) ;
    and03 ix5588 (.Y (nx5587), .A0 (nx6957), .A1 (nx7049), .A2 (nx7071)) ;
    inv01 ix6956 (.Y (nx6957), .A (nx6801)) ;
    and02 ix2627 (.Y (nx2626), .A0 (nx6991), .A1 (nx7057)) ;
    nand02 ix2603 (.Y (nx5728), .A0 (nx7057), .A1 (nx6995)) ;
    nor02_2x ix5592 (.Y (nx2098), .A0 (nx7027), .A1 (nx7021)) ;
    and04 ix5599 (.Y (nx5598), .A0 (nx6959), .A1 (nx7085), .A2 (nx4087), .A3 (
          nx6823)) ;
    inv01 ix6958 (.Y (nx6959), .A (current_state_6)) ;
    nor02_2x ix1951 (.Y (nx1950), .A0 (nx1930), .A1 (nx5197)) ;
    or02 ix5620 (.Y (nx5619), .A0 (nx4423), .A1 (nx7357)) ;
    or02 ix5622 (.Y (nx5621), .A0 (nx7357), .A1 (nx5194)) ;
    xor2 ix3040 (.Y (nx3039), .A0 (addr1_data_0), .A1 (nx7111)) ;
    or03 ix5626 (.Y (nx6905), .A0 (nx6993), .A1 (nx6711), .A2 (nx2706)) ;
    nor02ii ix2719 (.Y (nx6813), .A0 (nx7111), .A1 (nx4665)) ;
    mux21 ix3000 (.Y (nx2999), .A0 (write_offset_data_out_0), .A1 (nx5632), .S0 (
          nx7071)) ;
    or02 ix5637 (.Y (nx5636), .A0 (nx5632), .A1 (nx7358)) ;
    xor2 ix3030 (.Y (nx3029), .A0 (img_addr_offset_0), .A1 (nx7003)) ;
    nor02_2x ix2675 (.Y (nx6805), .A0 (nx1419), .A1 (reset)) ;
    mux21_ni ix3020 (.Y (nx3019), .A0 (nx5647), .A1 (img_base_addr_0), .S0 (
             nx7011)) ;
    mux21 ix3010 (.Y (nx3009), .A0 (nx5647), .A1 (nx7358), .S0 (nx7117)) ;
    xnor2 ix5654 (.Y (nx5653), .A0 (nx4433), .A1 (nx4039)) ;
    nor02ii ix2641 (.Y (nx2640), .A0 (nx2636), .A1 (current_state_12)) ;
    xnor2 ix2637 (.Y (nx2636), .A0 (nx4099), .A1 (nflt_layer_out_0)) ;
    xnor2 ix5658 (.Y (nx5657), .A0 (nx4459), .A1 (nx4053)) ;
    xor2 ix5660 (.Y (nx5659), .A0 (nx4485), .A1 (nflt_layer_out_3)) ;
    xnor2 ix5674 (.Y (nx5673), .A0 (nx5677), .A1 (nx5700)) ;
    mux21 ix3090 (.Y (nx3089), .A0 (nx5679), .A1 (nx5677), .S0 (nx7011)) ;
    mux21_ni ix3080 (.Y (nx3079), .A0 (write_base_prev_data_out_1), .A1 (
             write_base_data_out_1), .S0 (nx7117)) ;
    mux21 ix3050 (.Y (nx3049), .A0 (nx5687), .A1 (nx7359), .S0 (nx7095)) ;
    nor02ii ix5693 (.Y (nx5692), .A0 (write_base_prev_data_out_1), .A1 (nx5647)
            ) ;
    mux21 ix3100 (.Y (nx3099), .A0 (nx5700), .A1 (nx5696), .S0 (nx7003)) ;
    xnor2 ix5704 (.Y (nx5703), .A0 (nx5707), .A1 (nx7359)) ;
    ao32 ix3070 (.Y (nx3069), .A0 (nx6961), .A1 (nx7057), .A2 (nx6995), .B0 (
         bias_offset_data_out_1), .B1 (nx7071)) ;
    inv01 ix6960 (.Y (nx6961), .A (nx4287)) ;
    xnor2 ix5715 (.Y (nx5714), .A0 (nx7359), .A1 (nx5202)) ;
    mux21 ix3060 (.Y (nx3059), .A0 (nx5722), .A1 (nx5718), .S0 (nx7111)) ;
    nor02ii ix2605 (.Y (nx6793), .A0 (nx6983), .A1 (nx7071)) ;
    xnor2 ix5738 (.Y (nx5737), .A0 (nx5758), .A1 (nx5762)) ;
    mux21_ni ix3150 (.Y (nx3149), .A0 (nx2956), .A1 (img_base_addr_2), .S0 (
             nx7011)) ;
    mux21 ix3140 (.Y (nx3139), .A0 (nx5742), .A1 (nx7361), .S0 (nx7117)) ;
    mux21 ix3110 (.Y (nx3109), .A0 (nx5749), .A1 (nx7361), .S0 (nx7095)) ;
    mux21_ni ix3160 (.Y (nx3159), .A0 (img_addr_offset_2), .A1 (nx2970), .S0 (
             nx7003)) ;
    xor2 ix2971 (.Y (nx2970), .A0 (nx5762), .A1 (nx5698)) ;
    xnor2 ix5768 (.Y (nx5767), .A0 (nx5771), .A1 (nx7361)) ;
    ao32 ix3130 (.Y (nx3129), .A0 (nx6963), .A1 (nx7059), .A2 (nx6995), .B0 (
         bias_offset_data_out_2), .B1 (nx7071)) ;
    inv01 ix6962 (.Y (nx6963), .A (nx4281)) ;
    xnor2 ix5778 (.Y (nx5777), .A0 (nx7362), .A1 (nx4277)) ;
    xnor2 ix5784 (.Y (nx5783), .A0 (nx7362), .A1 (nx5208)) ;
    mux21_ni ix3120 (.Y (nx3119), .A0 (addr1_data_2), .A1 (nx2904), .S0 (nx7111)
             ) ;
    mux21_ni ix3210 (.Y (nx3209), .A0 (nx3100), .A1 (img_base_addr_3), .S0 (
             nx7011)) ;
    mux21_ni ix3200 (.Y (nx3199), .A0 (write_base_prev_data_out_3), .A1 (
             write_base_data_out_3), .S0 (nx7117)) ;
    mux21_ni ix3170 (.Y (nx3169), .A0 (nx3006), .A1 (write_base_data_out_3), .S0 (
             nx7095)) ;
    xor2 ix5806 (.Y (nx5805), .A0 (new_size_squared_out_3), .A1 (nx5807)) ;
    mux21_ni ix3220 (.Y (nx3219), .A0 (img_addr_offset_3), .A1 (nx3114), .S0 (
             nx7003)) ;
    xor2 ix5821 (.Y (nx5820), .A0 (bias_offset_data_out_3), .A1 (nx5807)) ;
    mux21_ni ix3190 (.Y (nx3189), .A0 (nx802), .A1 (bias_offset_data_out_3), .S0 (
             nx7071)) ;
    xor2 ix803 (.Y (nx802), .A0 (nx4271), .A1 (nx4299)) ;
    xnor2 ix5835 (.Y (nx5834), .A0 (nx5807), .A1 (nx5218)) ;
    mux21_ni ix3180 (.Y (nx3179), .A0 (addr1_data_3), .A1 (nx3048), .S0 (nx7111)
             ) ;
    xnor2 ix5851 (.Y (nx5850), .A0 (nx5807), .A1 (nx4271)) ;
    xnor2 ix5860 (.Y (nx5859), .A0 (nx5882), .A1 (nx5888)) ;
    mux21_ni ix3270 (.Y (nx3269), .A0 (nx3248), .A1 (img_base_addr_4), .S0 (
             nx7011)) ;
    mux21 ix3260 (.Y (nx3259), .A0 (nx5864), .A1 (nx5869), .S0 (nx7117)) ;
    mux21 ix3230 (.Y (nx3229), .A0 (nx5871), .A1 (nx5869), .S0 (nx7095)) ;
    xnor2 ix5877 (.Y (nx5876), .A0 (nx4391), .A1 (nx5869)) ;
    mux21_ni ix3280 (.Y (nx3279), .A0 (img_addr_offset_4), .A1 (nx3262), .S0 (
             nx7003)) ;
    nor02ii ix3257 (.Y (nx3256), .A0 (nx5886), .A1 (img_addr_offset_4)) ;
    xnor2 ix5896 (.Y (nx5895), .A0 (nx5900), .A1 (nx5869)) ;
    mux21_ni ix3250 (.Y (nx3249), .A0 (nx828), .A1 (bias_offset_data_out_4), .S0 (
             nx7071)) ;
    mux21_ni ix3240 (.Y (nx3239), .A0 (addr1_data_4), .A1 (nx3196), .S0 (nx7111)
             ) ;
    nor02ii ix3191 (.Y (nx3190), .A0 (nx5906), .A1 (addr1_data_4)) ;
    xnor2 ix5914 (.Y (nx5913), .A0 (nx5869), .A1 (nx4257)) ;
    xor2 ix5918 (.Y (nx5917), .A0 (nx5869), .A1 (nx3170)) ;
    xor2 ix5926 (.Y (nx5925), .A0 (img_base_addr_5), .A1 (nx5947)) ;
    mux21_ni ix3330 (.Y (nx3329), .A0 (nx3388), .A1 (img_base_addr_5), .S0 (
             nx7011)) ;
    mux21_ni ix3320 (.Y (nx3319), .A0 (write_base_prev_data_out_5), .A1 (
             write_base_data_out_5), .S0 (nx7117)) ;
    mux21_ni ix3290 (.Y (nx3289), .A0 (nx3298), .A1 (write_base_data_out_5), .S0 (
             nx7095)) ;
    xor2 ix5937 (.Y (nx5936), .A0 (new_size_squared_out_5), .A1 (nx5938)) ;
    mux21 ix3340 (.Y (nx3339), .A0 (nx5947), .A1 (nx5943), .S0 (nx7005)) ;
    xnor2 ix5952 (.Y (nx5951), .A0 (nx5955), .A1 (nx5938)) ;
    ao32 ix3310 (.Y (nx3309), .A0 (nx6965), .A1 (nx7059), .A2 (nx6995), .B0 (
         bias_offset_data_out_5), .B1 (nx7073)) ;
    inv01 ix6964 (.Y (nx6965), .A (nx4253)) ;
    mux21 ix3300 (.Y (nx3299), .A0 (nx5965), .A1 (nx5961), .S0 (nx7111)) ;
    xnor2 ix5972 (.Y (nx5971), .A0 (nx5938), .A1 (nx4251)) ;
    xor2 ix3319 (.Y (nx3318), .A0 (nx5938), .A1 (nx5977)) ;
    xnor2 ix5987 (.Y (nx5986), .A0 (nx6009), .A1 (nx6013)) ;
    mux21_ni ix3390 (.Y (nx3389), .A0 (nx3528), .A1 (img_base_addr_6), .S0 (
             nx7011)) ;
    mux21 ix3380 (.Y (nx3379), .A0 (nx5991), .A1 (nx5996), .S0 (nx7117)) ;
    mux21 ix3350 (.Y (nx3349), .A0 (nx5998), .A1 (nx5996), .S0 (nx7095)) ;
    xnor2 ix6004 (.Y (nx6003), .A0 (nx4377), .A1 (nx5996)) ;
    mux21_ni ix3400 (.Y (nx3399), .A0 (img_addr_offset_6), .A1 (nx3542), .S0 (
             nx7005)) ;
    nor02ii ix3537 (.Y (nx3536), .A0 (nx5945), .A1 (img_addr_offset_6)) ;
    xnor2 ix6021 (.Y (nx6020), .A0 (nx6025), .A1 (nx5996)) ;
    mux21_ni ix3370 (.Y (nx3369), .A0 (nx874), .A1 (bias_offset_data_out_6), .S0 (
             nx7073)) ;
    mux21_ni ix3360 (.Y (nx3359), .A0 (addr1_data_6), .A1 (nx3476), .S0 (nx7113)
             ) ;
    xor2 ix3477 (.Y (nx3476), .A0 (nx6031), .A1 (nx5963)) ;
    xnor2 ix6035 (.Y (nx6034), .A0 (nx5996), .A1 (nx4239)) ;
    nor02ii ix3313 (.Y (nx3312), .A0 (nx5977), .A1 (write_base_data_out_5)) ;
    xor2 ix6050 (.Y (nx6049), .A0 (img_base_addr_7), .A1 (nx6071)) ;
    mux21_ni ix3450 (.Y (nx3449), .A0 (nx3668), .A1 (img_base_addr_7), .S0 (
             nx7013)) ;
    mux21_ni ix3440 (.Y (nx3439), .A0 (write_base_prev_data_out_7), .A1 (
             write_base_data_out_7), .S0 (nx7119)) ;
    mux21_ni ix3410 (.Y (nx3409), .A0 (nx3578), .A1 (write_base_data_out_7), .S0 (
             nx7097)) ;
    xor2 ix6061 (.Y (nx6060), .A0 (new_size_squared_out_7), .A1 (nx6062)) ;
    mux21 ix3460 (.Y (nx3459), .A0 (nx6071), .A1 (nx6067), .S0 (nx7005)) ;
    xnor2 ix6076 (.Y (nx6075), .A0 (nx6079), .A1 (nx6062)) ;
    ao32 ix3430 (.Y (nx3429), .A0 (nx6967), .A1 (nx7059), .A2 (nx6995), .B0 (
         bias_offset_data_out_7), .B1 (nx7073)) ;
    inv01 ix6966 (.Y (nx6967), .A (nx4235)) ;
    mux21 ix3420 (.Y (nx3419), .A0 (nx6090), .A1 (nx6085), .S0 (nx7113)) ;
    nor02ii ix3471 (.Y (nx3470), .A0 (nx5963), .A1 (addr1_data_6)) ;
    nor02ii ix3593 (.Y (nx3592), .A0 (nx6042), .A1 (write_base_data_out_7)) ;
    xnor2 ix6101 (.Y (nx6100), .A0 (nx6062), .A1 (nx4229)) ;
    xnor2 ix6110 (.Y (nx6109), .A0 (nx6132), .A1 (nx6136)) ;
    mux21_ni ix3510 (.Y (nx3509), .A0 (nx3808), .A1 (img_base_addr_8), .S0 (
             nx7013)) ;
    mux21 ix3500 (.Y (nx3499), .A0 (nx6114), .A1 (nx6119), .S0 (nx7119)) ;
    mux21 ix3470 (.Y (nx3469), .A0 (nx6121), .A1 (nx6119), .S0 (nx7097)) ;
    xnor2 ix6127 (.Y (nx6126), .A0 (nx4363), .A1 (nx6119)) ;
    mux21_ni ix3520 (.Y (nx3519), .A0 (img_addr_offset_8), .A1 (nx3822), .S0 (
             nx7005)) ;
    nor02ii ix3817 (.Y (nx3816), .A0 (nx6069), .A1 (img_addr_offset_8)) ;
    xnor2 ix6144 (.Y (nx6143), .A0 (nx6148), .A1 (nx6119)) ;
    mux21_ni ix3490 (.Y (nx3489), .A0 (nx924), .A1 (bias_offset_data_out_8), .S0 (
             nx7073)) ;
    mux21_ni ix3480 (.Y (nx3479), .A0 (addr1_data_8), .A1 (nx3756), .S0 (nx7113)
             ) ;
    xor2 ix3757 (.Y (nx3756), .A0 (nx6154), .A1 (nx6088)) ;
    xnor2 ix6158 (.Y (nx6157), .A0 (nx6119), .A1 (nx4217)) ;
    xor2 ix6172 (.Y (nx6171), .A0 (img_base_addr_9), .A1 (nx6193)) ;
    mux21_ni ix3570 (.Y (nx3569), .A0 (nx3948), .A1 (img_base_addr_9), .S0 (
             nx7013)) ;
    mux21_ni ix3560 (.Y (nx3559), .A0 (write_base_prev_data_out_9), .A1 (
             write_base_data_out_9), .S0 (nx7119)) ;
    mux21_ni ix3530 (.Y (nx3529), .A0 (nx3858), .A1 (write_base_data_out_9), .S0 (
             nx7097)) ;
    xor2 ix6183 (.Y (nx6182), .A0 (new_size_squared_out_9), .A1 (nx6184)) ;
    mux21 ix3580 (.Y (nx3579), .A0 (nx6193), .A1 (nx6189), .S0 (nx7005)) ;
    xnor2 ix6198 (.Y (nx6197), .A0 (nx6201), .A1 (nx6184)) ;
    ao32 ix3550 (.Y (nx3549), .A0 (nx6969), .A1 (nx7059), .A2 (nx6995), .B0 (
         bias_offset_data_out_9), .B1 (nx7073)) ;
    inv01 ix6968 (.Y (nx6969), .A (nx4213)) ;
    mux21 ix3540 (.Y (nx3539), .A0 (nx6212), .A1 (nx6207), .S0 (nx7113)) ;
    nor02ii ix3751 (.Y (nx3750), .A0 (nx6088), .A1 (addr1_data_8)) ;
    nor02ii ix3873 (.Y (nx3872), .A0 (nx6164), .A1 (write_base_data_out_9)) ;
    xnor2 ix6223 (.Y (nx6222), .A0 (nx6184), .A1 (nx4301)) ;
    xnor2 ix6232 (.Y (nx6231), .A0 (nx6254), .A1 (nx6258)) ;
    mux21_ni ix3630 (.Y (nx3629), .A0 (nx4088), .A1 (img_base_addr_10), .S0 (
             nx7013)) ;
    mux21 ix3620 (.Y (nx3619), .A0 (nx6236), .A1 (nx6241), .S0 (nx7119)) ;
    mux21 ix3590 (.Y (nx3589), .A0 (nx6243), .A1 (nx6241), .S0 (nx7097)) ;
    xnor2 ix6249 (.Y (nx6248), .A0 (nx4349), .A1 (nx6241)) ;
    mux21_ni ix3640 (.Y (nx3639), .A0 (img_addr_offset_10), .A1 (nx4102), .S0 (
             nx7005)) ;
    nor02ii ix4097 (.Y (nx4096), .A0 (nx6191), .A1 (img_addr_offset_10)) ;
    xnor2 ix6266 (.Y (nx6265), .A0 (nx6270), .A1 (nx6241)) ;
    mux21_ni ix3610 (.Y (nx3609), .A0 (nx970), .A1 (bias_offset_data_out_10), .S0 (
             nx7073)) ;
    mux21_ni ix3600 (.Y (nx3599), .A0 (addr1_data_10), .A1 (nx4036), .S0 (nx7113
             )) ;
    xor2 ix4037 (.Y (nx4036), .A0 (nx6276), .A1 (nx6210)) ;
    xnor2 ix6280 (.Y (nx6279), .A0 (nx6241), .A1 (nx4200)) ;
    xor2 ix6294 (.Y (nx6293), .A0 (img_base_addr_11), .A1 (nx6315)) ;
    mux21_ni ix3690 (.Y (nx3689), .A0 (nx4228), .A1 (img_base_addr_11), .S0 (
             nx7013)) ;
    mux21_ni ix3680 (.Y (nx3679), .A0 (write_base_prev_data_out_11), .A1 (
             write_base_data_out_11), .S0 (nx7119)) ;
    mux21_ni ix3650 (.Y (nx3649), .A0 (nx4138), .A1 (write_base_data_out_11), .S0 (
             nx7097)) ;
    xor2 ix6305 (.Y (nx6304), .A0 (new_size_squared_out_11), .A1 (nx6306)) ;
    mux21 ix3700 (.Y (nx3699), .A0 (nx6315), .A1 (nx6311), .S0 (nx7005)) ;
    xnor2 ix6320 (.Y (nx6319), .A0 (nx6323), .A1 (nx6306)) ;
    ao32 ix3670 (.Y (nx3669), .A0 (nx6971), .A1 (nx7059), .A2 (nx6995), .B0 (
         bias_offset_data_out_11), .B1 (nx7073)) ;
    inv01 ix6970 (.Y (nx6971), .A (nx4197)) ;
    mux21 ix3660 (.Y (nx3659), .A0 (nx6334), .A1 (nx6329), .S0 (nx7113)) ;
    nor02ii ix4031 (.Y (nx4030), .A0 (nx6210), .A1 (addr1_data_10)) ;
    nor02ii ix4153 (.Y (nx4152), .A0 (nx6286), .A1 (write_base_data_out_11)) ;
    xnor2 ix6345 (.Y (nx6344), .A0 (nx6306), .A1 (nx4303)) ;
    xnor2 ix6354 (.Y (nx6353), .A0 (nx6376), .A1 (nx6380)) ;
    mux21_ni ix3750 (.Y (nx3749), .A0 (nx4368), .A1 (img_base_addr_12), .S0 (
             nx7013)) ;
    mux21 ix3740 (.Y (nx3739), .A0 (nx6358), .A1 (nx7363), .S0 (nx7119)) ;
    mux21 ix3710 (.Y (nx3709), .A0 (nx6365), .A1 (nx7363), .S0 (nx7097)) ;
    mux21_ni ix3760 (.Y (nx3759), .A0 (img_addr_offset_12), .A1 (nx4382), .S0 (
             nx7007)) ;
    nor02ii ix4377 (.Y (nx4376), .A0 (nx6313), .A1 (img_addr_offset_12)) ;
    xnor2 ix6388 (.Y (nx6387), .A0 (nx6392), .A1 (nx7363)) ;
    mux21_ni ix3730 (.Y (nx3729), .A0 (nx1018), .A1 (bias_offset_data_out_12), .S0 (
             nx7075)) ;
    mux21_ni ix3720 (.Y (nx3719), .A0 (addr1_data_12), .A1 (nx4316), .S0 (nx7113
             )) ;
    xor2 ix4317 (.Y (nx4316), .A0 (nx6398), .A1 (nx6332)) ;
    xnor2 ix6409 (.Y (nx6408), .A0 (nx7363), .A1 (nx4183)) ;
    xor2 ix6416 (.Y (nx6415), .A0 (img_base_addr_13), .A1 (nx6437)) ;
    mux21_ni ix3810 (.Y (nx3809), .A0 (nx4508), .A1 (img_base_addr_13), .S0 (
             nx7013)) ;
    mux21_ni ix3800 (.Y (nx3799), .A0 (write_base_prev_data_out_13), .A1 (
             write_base_data_out_13), .S0 (nx7119)) ;
    mux21_ni ix3770 (.Y (nx3769), .A0 (nx4418), .A1 (write_base_data_out_13), .S0 (
             nx7097)) ;
    xor2_2x ix6427 (.Y (nx6426), .A0 (new_size_squared_out_13), .A1 (nx6428)) ;
    mux21 ix3820 (.Y (nx3819), .A0 (nx6437), .A1 (nx6433), .S0 (nx7007)) ;
    xnor2 ix6442 (.Y (nx6441), .A0 (nx6445), .A1 (nx6428)) ;
    ao32 ix3790 (.Y (nx3789), .A0 (nx6973), .A1 (nx7059), .A2 (nx6997), .B0 (
         bias_offset_data_out_13), .B1 (nx7075)) ;
    inv01 ix6972 (.Y (nx6973), .A (nx4180)) ;
    mux21 ix3780 (.Y (nx3779), .A0 (nx6456), .A1 (nx6451), .S0 (nx7115)) ;
    nor02ii ix4311 (.Y (nx4310), .A0 (nx6332), .A1 (addr1_data_12)) ;
    nor02ii ix4433 (.Y (nx4432), .A0 (nx6404), .A1 (write_base_data_out_13)) ;
    xnor2 ix6467 (.Y (nx6466), .A0 (nx6428), .A1 (nx4305)) ;
    xnor2 ix6476 (.Y (nx6475), .A0 (nx6496), .A1 (nx6500)) ;
    mux21_ni ix3870 (.Y (nx3869), .A0 (nx4648), .A1 (img_base_addr_14), .S0 (
             nx7015)) ;
    xnor2 ix4649 (.Y (nx4648), .A0 (nx6493), .A1 (nx6494)) ;
    mux21 ix3860 (.Y (nx3859), .A0 (nx6493), .A1 (nx7365), .S0 (nx7121)) ;
    mux21 ix3830 (.Y (nx3829), .A0 (nx6486), .A1 (nx7365), .S0 (nx7099)) ;
    mux21_ni ix3880 (.Y (nx3879), .A0 (img_addr_offset_14), .A1 (nx4662), .S0 (
             nx7007)) ;
    xor2 ix4663 (.Y (nx4662), .A0 (nx6500), .A1 (nx6435)) ;
    xnor2 ix6506 (.Y (nx6505), .A0 (nx6510), .A1 (nx7365)) ;
    mux21_ni ix3850 (.Y (nx3849), .A0 (nx1064), .A1 (bias_offset_data_out_14), .S0 (
             nx7075)) ;
    xor2 ix1065 (.Y (nx1064), .A0 (nx4167), .A1 (nx4175)) ;
    mux21_ni ix3840 (.Y (nx3839), .A0 (addr1_data_14), .A1 (nx4596), .S0 (nx7115
             )) ;
    xor2 ix4597 (.Y (nx4596), .A0 (nx6516), .A1 (nx6454)) ;
    xor2 ix6521 (.Y (nx6520), .A0 (nx7365), .A1 (nx4432)) ;
    xnor2 ix6525 (.Y (nx6524), .A0 (nx7366), .A1 (nx4167)) ;
    xor2 ix6544 (.Y (nx6543), .A0 (img_base_addr_15), .A1 (nx6558)) ;
    mux21_ni ix3930 (.Y (nx3929), .A0 (nx4764), .A1 (img_base_addr_15), .S0 (
             nx7015)) ;
    mux21_ni ix3920 (.Y (nx3919), .A0 (write_base_prev_data_out_15), .A1 (
             write_base_data_out_15), .S0 (nx7121)) ;
    mux21 ix3940 (.Y (nx3939), .A0 (nx6558), .A1 (nx6555), .S0 (nx7007)) ;
    xor2 ix6556 (.Y (nx6555), .A0 (nx6558), .A1 (nx4656)) ;
    nor02ii ix4657 (.Y (nx4656), .A0 (nx6435), .A1 (img_addr_offset_14)) ;
    xor2 ix4735 (.Y (nx4734), .A0 (write_base_data_out_15), .A1 (
         write_offset_data_out_15)) ;
    mux21 ix3910 (.Y (nx3909), .A0 (nx6572), .A1 (nx6569), .S0 (nx7115)) ;
    xor2 ix6570 (.Y (nx6569), .A0 (nx6572), .A1 (nx4590)) ;
    nor02ii ix4591 (.Y (nx4590), .A0 (nx6454), .A1 (addr1_data_14)) ;
    xor2 ix6577 (.Y (nx6576), .A0 (nx6580), .A1 (write_base_data_out_15)) ;
    ao32 ix3890 (.Y (nx3889), .A0 (nx6975), .A1 (nx7059), .A2 (nx6997), .B0 (
         bias_offset_data_out_15), .B1 (nx7075)) ;
    inv01 ix6974 (.Y (nx6975), .A (nx4163)) ;
    nor02ii ix6758 (.Y (nx6759), .A0 (nx6929), .A1 (current_state_12)) ;
    nor02ii ix6760 (.Y (nx6761), .A0 (nx6929), .A1 (current_state_12)) ;
    and02 ix6800 (.Y (nx6801), .A0 (nx6991), .A1 (nx7061)) ;
    and02 ix6802 (.Y (nx6803), .A0 (nx6991), .A1 (nx7061)) ;
    inv02 ix6976 (.Y (nx6977), .A (nx4883)) ;
    inv02 ix6978 (.Y (nx6979), .A (nx4883)) ;
    inv01 ix6980 (.Y (nx6981), .A (nx6829)) ;
    inv01 ix6982 (.Y (nx6983), .A (nx6829)) ;
    inv01 ix6984 (.Y (nx6985), .A (nx6851)) ;
    inv01 ix6986 (.Y (nx6987), .A (nx6851)) ;
    inv01 ix6988 (.Y (nx6989), .A (nx6851)) ;
    inv01 ix6990 (.Y (nx6991), .A (nx6851)) ;
    buf02 ix6992 (.Y (nx6993), .A (nx2084)) ;
    inv02 ix6994 (.Y (nx6995), .A (nx6897)) ;
    inv02 ix6996 (.Y (nx6997), .A (nx6897)) ;
    inv02 ix6998 (.Y (nx6999), .A (nx7107)) ;
    inv02 ix7000 (.Y (nx7001), .A (nx7107)) ;
    inv02 ix7002 (.Y (nx7003), .A (nx7107)) ;
    inv02 ix7004 (.Y (nx7005), .A (nx6871)) ;
    inv02 ix7006 (.Y (nx7007), .A (nx6871)) ;
    inv02 ix7008 (.Y (nx7009), .A (nx6665)) ;
    inv02 ix7010 (.Y (nx7011), .A (nx6665)) ;
    inv02 ix7012 (.Y (nx7013), .A (nx6665)) ;
    inv02 ix7014 (.Y (nx7015), .A (nx6665)) ;
    buf02 ix7016 (.Y (nx7017), .A (nx4033)) ;
    inv02 ix7018 (.Y (nx7019), .A (nx1528)) ;
    inv01 ix7020 (.Y (nx7021), .A (nx6705)) ;
    inv02 ix7022 (.Y (nx7023), .A (nx6749)) ;
    inv02 ix7024 (.Y (nx7025), .A (nx6749)) ;
    inv02 ix7026 (.Y (nx7027), .A (nx6749)) ;
    inv02 ix7032 (.Y (nx7033), .A (nx6685)) ;
    inv02 ix7034 (.Y (nx7035), .A (nx6685)) ;
    inv02 ix7036 (.Y (nx7037), .A (nx1429)) ;
    inv02 ix7038 (.Y (nx7039), .A (nx1429)) ;
    inv02 ix7040 (.Y (nx7041), .A (nx1429)) ;
    inv02 ix7042 (.Y (nx7043), .A (argmax_ready)) ;
    inv02 ix7048 (.Y (nx7049), .A (argmax_ready)) ;
    inv01 ix7050 (.Y (nx7051), .A (nx5243)) ;
    inv02 ix7052 (.Y (nx7053), .A (nx7051)) ;
    inv02 ix7054 (.Y (nx7055), .A (nx7051)) ;
    inv02 ix7056 (.Y (nx7057), .A (nx7051)) ;
    inv02 ix7058 (.Y (nx7059), .A (nx7051)) ;
    inv02 ix7060 (.Y (nx7061), .A (nx7051)) ;
    inv02 ix7064 (.Y (nx7065), .A (comp_unit_flt_size)) ;
    inv02 ix7070 (.Y (nx7071), .A (nx6787)) ;
    inv02 ix7072 (.Y (nx7073), .A (nx6787)) ;
    inv02 ix7074 (.Y (nx7075), .A (nx6787)) ;
    inv01 ix7076 (.Y (nx7077), .A (nx7293)) ;
    inv01 ix7078 (.Y (nx7079), .A (nx7293)) ;
    inv02 ix7080 (.Y (nx7081), .A (current_state_7)) ;
    inv02 ix7082 (.Y (nx7083), .A (current_state_7)) ;
    inv02 ix7084 (.Y (nx7085), .A (current_state_7)) ;
    inv02 ix7086 (.Y (nx7087), .A (nx6731)) ;
    inv02 ix7088 (.Y (nx7089), .A (nx6731)) ;
    buf02 ix7090 (.Y (nx7091), .A (nx6759)) ;
    buf02 ix7092 (.Y (nx7093), .A (nx6761)) ;
    inv02 ix7094 (.Y (nx7095), .A (nx2580)) ;
    inv02 ix7096 (.Y (nx7097), .A (nx2580)) ;
    inv02 ix7098 (.Y (nx7099), .A (nx2580)) ;
    inv02 ix7100 (.Y (nx7101), .A (nx5099)) ;
    inv02 ix7102 (.Y (nx7103), .A (nx5099)) ;
    inv02 ix7104 (.Y (nx7105), .A (nx5099)) ;
    inv02 ix7106 (.Y (nx7107), .A (nx2536)) ;
    inv01 ix7108 (.Y (nx7109), .A (nx6905)) ;
    inv02 ix7110 (.Y (nx7111), .A (nx7109)) ;
    inv02 ix7112 (.Y (nx7113), .A (nx7109)) ;
    inv02 ix7114 (.Y (nx7115), .A (nx7109)) ;
    inv02 ix7116 (.Y (nx7117), .A (nx5651)) ;
    inv02 ix7118 (.Y (nx7119), .A (nx5651)) ;
    inv02 ix7120 (.Y (nx7121), .A (nx5651)) ;
    inv01 ix7122 (.Y (nx7123), .A (nx7145)) ;
    inv01 ix7124 (.Y (nx7125), .A (nx7145)) ;
    inv01 ix7126 (.Y (nx7127), .A (nx7145)) ;
    inv01 ix7128 (.Y (nx7129), .A (nx7145)) ;
    inv01 ix7130 (.Y (nx7131), .A (nx5501)) ;
    inv01 ix7132 (.Y (nx7133), .A (nx5501)) ;
    inv01 ix7134 (.Y (nx7135), .A (nx5501)) ;
    inv01 ix7136 (.Y (nx7137), .A (nx5501)) ;
    inv01 ix7138 (.Y (nx7139), .A (nx5501)) ;
    inv01 ix7144 (.Y (nx7145), .A (nx2502)) ;
    oai21 ix291 (.Y (filter_ready_out), .A0 (nx7029), .A1 (nx4593), .B0 (nx4665)
          ) ;
    inv02 ix7028 (.Y (nx7029), .A (nx6711)) ;
    inv01 ix4594 (.Y (nx4593), .A (nx286)) ;
    or02 ix4666 (.Y (nx4665), .A0 (nx4637), .A1 (nx7021)) ;
    inv02 ix7062 (.Y (nx7063), .A (comp_unit_flt_size)) ;
    inv01 ix273 (.Y (comp_unit_flt_size), .A (nx5482)) ;
    inv02 ix7030 (.Y (nx7031), .A (nx6711)) ;
    inv02 ix6710 (.Y (nx6711), .A (nx4589)) ;
    buf04 ix7368 (.Y (nx7293), .A (filter_ready_out)) ;
    buf04 ix7369 (.Y (nx7294), .A (nx7063)) ;
    buf04 ix7370 (.Y (nx7295), .A (nx7031)) ;
    inv02 ix7371 (.Y (nx7296), .A (new_size_squared_out_15)) ;
    inv02 ix7372 (.Y (nx7297), .A (write_base_data_out_15)) ;
    oai32 ix7373 (.Y (nx7298), .A0 (nx7099), .A1 (nx7296), .A2 (
          write_base_data_out_15), .B0 (nx7297), .B1 (new_size_squared_out_15)
          ) ;
    and02 ix7374 (.Y (nx7299), .A0 (nx7364), .A1 (nx4335)) ;
    nor02_2x ix7375 (.Y (nx7300), .A0 (nx7364), .A1 (nx4335)) ;
    and02 ix7376 (.Y (nx7301), .A0 (nx7366), .A1 (nx4320)) ;
    inv02 ix7377 (.Y (nx7302), .A (write_base_data_out_13)) ;
    inv02 ix7378 (.Y (nx7303), .A (new_size_squared_out_13)) ;
    inv02 ix7379 (.Y (nx7304), .A (nx7099)) ;
    aoi32 ix7380 (.Y (nx7305), .A0 (nx7304), .A1 (nx7297), .A2 (nx7296), .B0 (
          write_base_data_out_15), .B1 (new_size_squared_out_15)) ;
    ao221 reg_nx3899 (.Y (nx3899), .A0 (nx7298), .A1 (NOT_nx4700), .B0 (
          write_base_data_out_15), .B1 (nx7099), .C0 (nx7350)) ;
    and02 ix7381 (.Y (nx7306), .A0 (write_base_data_out_13), .A1 (
          new_size_squared_out_13)) ;
    inv02 ix7382 (.Y (nx7307), .A (nx6426)) ;
    oai32 reg_nx6488 (.Y (nx6488), .A0 (nx7306), .A1 (nx7354), .A2 (nx7300), .B0 (
          nx7307), .B1 (nx7306)) ;
    inv01 ix7383 (.Y (nx7308), .A (nx7366)) ;
    inv02 ix7384 (.Y (nx7309), .A (nx4320)) ;
    oai22 reg_nx6491 (.Y (nx6491), .A0 (nx7308), .A1 (nx7309), .B0 (nx7366), .B1 (
          nx4320)) ;
    oai22 reg_nx4414 (.Y (nx4414), .A0 (nx7364), .A1 (nx4335), .B0 (nx7299), .B1 (
          nx7445)) ;
    inv02 ix7385 (.Y (nx7310), .A (nx7364)) ;
    inv02 ix7386 (.Y (nx7311), .A (nx4335)) ;
    oai22 reg_nx6370 (.Y (nx6370), .A0 (nx7310), .A1 (nx7311), .B0 (nx7364), .B1 (
          nx4335)) ;
    inv01 ix7387 (.Y (nx7312), .A (nx7362)) ;
    inv01 ix7388 (.Y (nx7313), .A (nx4407)) ;
    nand02_2x ix7389 (.Y (nx7314), .A0 (nx7362), .A1 (nx4407)) ;
    inv01 ix7390 (.Y (nx7315), .A (nx7359)) ;
    nand03_2x ix7391 (.Y (nx7316), .A0 (new_size_squared_out_0), .A1 (nx6775), .A2 (
              nx7315)) ;
    inv01 ix7392 (.Y (nx7317), .A (new_size_squared_out_1)) ;
    nand02_2x ix7393 (.Y (nx7318), .A0 (new_size_squared_out_1), .A1 (nx7315)) ;
    nand03_2x ix7394 (.Y (nx7319), .A0 (nx7318), .A1 (new_size_squared_out_0), .A2 (
              nx6775)) ;
    inv01 ix7395 (.Y (nx7320), .A (write_base_data_out_1)) ;
    aoi22 ix7396 (.Y (nx7321), .A0 (nx7316), .A1 (nx7317), .B0 (nx7319), .B1 (
          nx7320)) ;
    aoi22 ix7397 (.Y (nx7322), .A0 (nx7312), .A1 (nx7313), .B0 (nx7314), .B1 (
          nx7321)) ;
    inv01 reg_nx3002 (.Y (nx3002), .A (nx7322)) ;
    inv01 ix7398 (.Y (nx7323), .A (nx7322)) ;
    inv01 reg_nx5751 (.Y (nx5751), .A (nx7321)) ;
    oai22 reg_nx5754 (.Y (nx5754), .A0 (nx7312), .A1 (nx7313), .B0 (nx7362), .B1 (
          nx4407)) ;
    oai22 reg_nx5689 (.Y (nx5689), .A0 (nx7315), .A1 (new_size_squared_out_1), .B0 (
          nx7317), .B1 (nx7360)) ;
    inv01 ix7399 (.Y (nx7324), .A (mem_data_in[3])) ;
    nor03_2x reg_argmax_data_out_3 (.Y (argmax_data_out[3]), .A0 (nx7338), .A1 (
             nx7324), .A2 (nx7340)) ;
    inv02 reg_nx5191 (.Y (nx5191), .A (argmax_ready)) ;
    inv01 reg_argmax_ready (.Y (argmax_ready_dup0), .A (argmax_ready)) ;
    inv01 ix7400 (.Y (nx7325), .A (nx7367)) ;
    inv01 ix7401 (.Y (nx7326), .A (nx7367)) ;
    inv01 ix7402 (.Y (nx7327), .A (nx7367)) ;
    inv01 ix7403 (.Y (nx7328), .A (nx7367)) ;
    inv01 reg_nx1930 (.Y (nx1930), .A (nx7338)) ;
    nand02_2x ix7404 (.Y (nx7329), .A0 (write_offset_data_out_2), .A1 (
              write_base_data_out_2)) ;
    inv01 ix7405 (.Y (nx7330), .A (nx7356)) ;
    inv01 ix7406 (.Y (nx7331), .A (nx7360)) ;
    nand02_2x ix7407 (.Y (nx7332), .A0 (nx7356), .A1 (nx7360)) ;
    nor02_2x ix7408 (.Y (nx7333), .A0 (nx7358), .A1 (nx4293)) ;
    aoi22 ix7409 (.Y (nx7334), .A0 (nx7330), .A1 (nx7331), .B0 (nx7332), .B1 (
          nx7333)) ;
    aoi22 ix7410 (.Y (nx7335), .A0 (nx7329), .A1 (nx7334), .B0 (nx5777), .B1 (
          nx7329)) ;
    inv02 reg_nx5847 (.Y (nx5847), .A (nx7335)) ;
    inv01 ix7411 (.Y (nx7336), .A (nx7335)) ;
    and02 ix7412 (.Y (nx7337), .A0 (nx7356), .A1 (nx7360)) ;
    oai32 reg_nx2850 (.Y (nx2850), .A0 (nx7337), .A1 (nx7358), .A2 (nx4293), .B0 (
          nx7356), .B1 (nx7360)) ;
    or02 reg_nx5667 (.Y (nx5667), .A0 (nx7358), .A1 (nx4293)) ;
    oai22 reg_nx5725 (.Y (nx5725), .A0 (nx7330), .A1 (nx7331), .B0 (nx7356), .B1 (
          nx7360)) ;
    inv01 reg_nx6775 (.Y (nx6775), .A (nx7358)) ;
    inv01 reg_nx7047 (.Y (nx7047), .A (nx7367)) ;
    nor04_2x ix7413 (.Y (nx7338), .A0 (class_cntr_counter_out_0), .A1 (
             class_cntr_counter_out_2), .A2 (nx5202), .A3 (nx5218)) ;
    inv01 ix7414 (.Y (nx7339), .A (mem_data_in[6])) ;
    inv01 ix7415 (.Y (nx7340), .A (current_state_27)) ;
    nor03_2x reg_argmax_data_out_6 (.Y (argmax_data_out[6]), .A0 (nx7338), .A1 (
             nx7339), .A2 (nx7340)) ;
    nor02_2x reg_argmax_ready_XX0_XREP5 (.Y (argmax_ready_XX0_XREP5), .A0 (
             nx7340), .A1 (nx7338)) ;
    inv02 ix7416 (.Y (nx7341), .A (nx6426)) ;
    inv01 ix7417 (.Y (nx7342), .A (nx7301)) ;
    inv01 ix7418 (.Y (nx7343), .A (nx7299)) ;
    nand03_2x ix7419 (.Y (nx7344), .A0 (nx7341), .A1 (nx7342), .A2 (nx7343)) ;
    inv01 ix7420 (.Y (nx7345), .A (nx7366)) ;
    inv02 ix7421 (.Y (nx7346), .A (nx4320)) ;
    nor02_2x ix7422 (.Y (nx7347), .A0 (nx7302), .A1 (nx7303)) ;
    nor02ii ix7423 (.Y (nx7348), .A0 (nx6426), .A1 (nx7300)) ;
    aoi222 ix7424 (.Y (nx7349), .A0 (nx7345), .A1 (nx7346), .B0 (nx7342), .B1 (
           nx7347), .C0 (nx7342), .C1 (nx7348)) ;
    oai32 ix7425 (.Y (nx7350), .A0 (nx7305), .A1 (nx7445), .A2 (nx7344), .B0 (
          nx7349), .B1 (nx7305)) ;
    inv02 ix7426 (.Y (nx7351), .A (nx7300)) ;
    oai22 ix7427 (.Y (nx7352), .A0 (nx7351), .A1 (nx6426), .B0 (nx7302), .B1 (
          nx7303)) ;
    nor04_2x ix7428 (.Y (nx7353), .A0 (nx7445), .A1 (nx6426), .A2 (nx7301), .A3 (
             nx7299)) ;
    aoi221 reg_NOT_nx4700 (.Y (NOT_nx4700), .A0 (nx7345), .A1 (nx7346), .B0 (
           nx7352), .B1 (nx7342), .C0 (nx7353)) ;
    nor02_2x ix7429 (.Y (nx7354), .A0 (nx7445), .A1 (nx7299)) ;
    buf16 ix7430 (.Y (nx7355), .A (nx4284)) ;
    buf16 ix7431 (.Y (nx7356), .A (nx4284)) ;
    buf16 ix7432 (.Y (nx7357), .A (nx5611)) ;
    buf16 ix7433 (.Y (nx7358), .A (nx5611)) ;
    buf16 ix7434 (.Y (nx7359), .A (nx5685)) ;
    buf16 ix7435 (.Y (nx7360), .A (nx5685)) ;
    buf16 ix7436 (.Y (nx7361), .A (nx5747)) ;
    buf16 ix7437 (.Y (nx7362), .A (nx5747)) ;
    buf16 ix7438 (.Y (nx7363), .A (nx6363)) ;
    buf16 ix7439 (.Y (nx7364), .A (nx6363)) ;
    buf16 ix7440 (.Y (nx7365), .A (nx6484)) ;
    buf16 ix7441 (.Y (nx7366), .A (nx6484)) ;
    buf16 ix7442 (.Y (argmax_ready), .A (argmax_ready_XX0_XREP5)) ;
    buf16 ix7443 (.Y (nx7367), .A (argmax_ready_XX0_XREP5)) ;
    buf02 ix7444 (.Y (nx7445), .A (nx6367)) ;
endmodule


module AdvancedCounter_16 ( clk, reset, enable, mode_in, max_val_in, 
                            max_reached_out, counter_out ) ;

    input clk ;
    input reset ;
    input enable ;
    input [1:0]mode_in ;
    input [15:0]max_val_in ;
    output max_reached_out ;
    output [15:0]counter_out ;

    wire counter_out_15_rename, counter_out_14_rename, nx149, 
         counter_out_13_rename, counter_out_12_rename, nx152, 
         counter_out_11_rename, counter_out_10_rename, nx155, 
         counter_out_9_rename, counter_out_8_rename, nx157, counter_out_7_rename, 
         counter_out_6_rename, nx159, counter_out_5_rename, counter_out_4_rename, 
         nx161, counter_out_3_rename, counter_out_2_rename, counter_out_1_rename, 
         counter_out_dup0_0, nx22, nx34, nx46, nx70, nx94, nx118, nx142, nx166, 
         nx174, nx192, nx206, nx224, nx246, nx173, nx183, nx193, nx203, nx213, 
         nx223, nx233, nx243, nx253, nx263, nx273, nx283, nx293, nx303, nx313, 
         nx323, nx339, nx344, nx348, nx350, nx353, nx358, nx362, nx364, nx367, 
         nx372, nx376, nx378, nx381, nx386, nx390, nx392, nx395, nx400, nx404, 
         nx406, nx409, nx414, nx419, nx424, nx428, nx430, nx436, nx439, nx445, 
         nx447, nx449, nx451, nx458, nx460, nx462, nx464, nx466, nx468, nx470, 
         nx472, nx474;
    wire [1:0] \$dummy ;




    assign counter_out[14] = counter_out[15] ;
    assign counter_out[13] = counter_out[15] ;
    assign counter_out[12] = counter_out[15] ;
    assign counter_out[11] = counter_out[15] ;
    assign counter_out[10] = counter_out[15] ;
    assign counter_out[9] = counter_out[15] ;
    assign counter_out[8] = counter_out[15] ;
    assign counter_out[7] = counter_out[15] ;
    assign counter_out[6] = counter_out[15] ;
    assign counter_out[5] = counter_out[15] ;
    assign counter_out[4] = counter_out[15] ;
    assign counter_out[3] = counter_out[15] ;
    assign counter_out[2] = counter_out[15] ;
    assign counter_out[1] = counter_out[15] ;
    assign counter_out[0] = counter_out[15] ;
    fake_gnd ix140 (.Y (counter_out[15])) ;
    and04 ix251 (.Y (max_reached_out), .A0 (nx192), .A1 (nx206), .A2 (nx224), .A3 (
          nx246)) ;
    mux21_ni ix324 (.Y (nx323), .A0 (counter_out_15_rename), .A1 (nx174), .S0 (
             nx474)) ;
    mux21_ni ix314 (.Y (nx313), .A0 (counter_out_14_rename), .A1 (nx166), .S0 (
             nx472)) ;
    dffr reg_counter_data_14 (.Q (counter_out_14_rename), .QB (nx339), .D (nx313
         ), .CLK (clk), .R (nx462)) ;
    nand02 ix345 (.Y (nx344), .A0 (counter_out_13_rename), .A1 (nx152)) ;
    mux21 ix304 (.Y (nx303), .A0 (nx348), .A1 (nx350), .S0 (nx472)) ;
    dffr reg_counter_data_13 (.Q (counter_out_13_rename), .QB (nx348), .D (nx303
         ), .CLK (clk), .R (nx462)) ;
    oai21 ix351 (.Y (nx350), .A0 (nx152), .A1 (counter_out_13_rename), .B0 (
          nx344)) ;
    mux21_ni ix294 (.Y (nx293), .A0 (counter_out_12_rename), .A1 (nx142), .S0 (
             nx472)) ;
    dffr reg_counter_data_12 (.Q (counter_out_12_rename), .QB (nx353), .D (nx293
         ), .CLK (clk), .R (nx462)) ;
    nand02 ix359 (.Y (nx358), .A0 (counter_out_11_rename), .A1 (nx155)) ;
    mux21 ix284 (.Y (nx283), .A0 (nx362), .A1 (nx364), .S0 (nx472)) ;
    dffr reg_counter_data_11 (.Q (counter_out_11_rename), .QB (nx362), .D (nx283
         ), .CLK (clk), .R (nx462)) ;
    oai21 ix365 (.Y (nx364), .A0 (nx155), .A1 (counter_out_11_rename), .B0 (
          nx358)) ;
    mux21_ni ix274 (.Y (nx273), .A0 (counter_out_10_rename), .A1 (nx118), .S0 (
             nx472)) ;
    dffr reg_counter_data_10 (.Q (counter_out_10_rename), .QB (nx367), .D (nx273
         ), .CLK (clk), .R (nx462)) ;
    nand02 ix373 (.Y (nx372), .A0 (counter_out_9_rename), .A1 (nx157)) ;
    mux21 ix264 (.Y (nx263), .A0 (nx376), .A1 (nx378), .S0 (nx472)) ;
    dffr reg_counter_data_9 (.Q (counter_out_9_rename), .QB (nx376), .D (nx263)
         , .CLK (clk), .R (nx462)) ;
    oai21 ix379 (.Y (nx378), .A0 (nx157), .A1 (counter_out_9_rename), .B0 (nx372
          )) ;
    mux21_ni ix254 (.Y (nx253), .A0 (counter_out_8_rename), .A1 (nx94), .S0 (
             nx472)) ;
    dffr reg_counter_data_8 (.Q (counter_out_8_rename), .QB (nx381), .D (nx253)
         , .CLK (clk), .R (nx462)) ;
    nand02 ix387 (.Y (nx386), .A0 (counter_out_7_rename), .A1 (nx159)) ;
    mux21 ix244 (.Y (nx243), .A0 (nx390), .A1 (nx392), .S0 (nx470)) ;
    dffr reg_counter_data_7 (.Q (counter_out_7_rename), .QB (nx390), .D (nx243)
         , .CLK (clk), .R (nx464)) ;
    oai21 ix393 (.Y (nx392), .A0 (nx159), .A1 (counter_out_7_rename), .B0 (nx386
          )) ;
    mux21_ni ix234 (.Y (nx233), .A0 (counter_out_6_rename), .A1 (nx70), .S0 (
             nx470)) ;
    dffr reg_counter_data_6 (.Q (counter_out_6_rename), .QB (nx395), .D (nx233)
         , .CLK (clk), .R (nx464)) ;
    nand02 ix401 (.Y (nx400), .A0 (counter_out_5_rename), .A1 (nx161)) ;
    mux21 ix224 (.Y (nx223), .A0 (nx404), .A1 (nx406), .S0 (nx470)) ;
    dffr reg_counter_data_5 (.Q (counter_out_5_rename), .QB (nx404), .D (nx223)
         , .CLK (clk), .R (nx464)) ;
    oai21 ix407 (.Y (nx406), .A0 (nx161), .A1 (counter_out_5_rename), .B0 (nx400
          )) ;
    mux21_ni ix214 (.Y (nx213), .A0 (counter_out_4_rename), .A1 (nx46), .S0 (
             nx470)) ;
    dffr reg_counter_data_4 (.Q (counter_out_4_rename), .QB (nx409), .D (nx213)
         , .CLK (clk), .R (nx464)) ;
    aoi21 ix47 (.Y (nx46), .A0 (nx414), .A1 (nx409), .B0 (nx161)) ;
    nand04 ix415 (.Y (nx414), .A0 (counter_out_3_rename), .A1 (
           counter_out_2_rename), .A2 (counter_out_1_rename), .A3 (
           counter_out_dup0_0)) ;
    dffr reg_counter_data_3 (.Q (counter_out_3_rename), .QB (\$dummy [0]), .D (
         nx203), .CLK (clk), .R (nx466)) ;
    mux21_ni ix204 (.Y (nx203), .A0 (counter_out_3_rename), .A1 (nx34), .S0 (
             nx470)) ;
    xnor2 ix35 (.Y (nx34), .A0 (counter_out_3_rename), .A1 (nx419)) ;
    nand03 ix420 (.Y (nx419), .A0 (counter_out_2_rename), .A1 (
           counter_out_1_rename), .A2 (counter_out_dup0_0)) ;
    dffr reg_counter_data_2 (.Q (counter_out_2_rename), .QB (\$dummy [1]), .D (
         nx193), .CLK (clk), .R (nx464)) ;
    mux21_ni ix194 (.Y (nx193), .A0 (counter_out_2_rename), .A1 (nx22), .S0 (
             nx470)) ;
    xnor2 ix23 (.Y (nx22), .A0 (counter_out_2_rename), .A1 (nx424)) ;
    mux21 ix184 (.Y (nx183), .A0 (nx428), .A1 (nx430), .S0 (nx470)) ;
    dffr reg_counter_data_1 (.Q (counter_out_1_rename), .QB (nx428), .D (nx183)
         , .CLK (clk), .R (nx464)) ;
    oai21 ix431 (.Y (nx430), .A0 (counter_out_dup0_0), .A1 (counter_out_1_rename
          ), .B0 (nx424)) ;
    dffr reg_counter_data_0 (.Q (counter_out_dup0_0), .QB (nx436), .D (nx173), .CLK (
         clk), .R (nx464)) ;
    dffr reg_counter_data_15 (.Q (counter_out_15_rename), .QB (nx439), .D (nx323
         ), .CLK (clk), .R (nx466)) ;
    and04 ix247 (.Y (nx246), .A0 (nx445), .A1 (nx447), .A2 (nx449), .A3 (nx451)
          ) ;
    xnor2 ix448 (.Y (nx447), .A0 (counter_out_2_rename), .A1 (max_val_in[2])) ;
    xnor2 ix450 (.Y (nx449), .A0 (counter_out_3_rename), .A1 (max_val_in[3])) ;
    and04 ix193 (.Y (nx192), .A0 (nx439), .A1 (nx339), .A2 (nx348), .A3 (nx353)
          ) ;
    xor2 ix175 (.Y (nx174), .A0 (nx149), .A1 (counter_out_15_rename)) ;
    nor02ii ix173 (.Y (nx149), .A0 (nx344), .A1 (counter_out_14_rename)) ;
    xor2 ix167 (.Y (nx166), .A0 (nx339), .A1 (nx344)) ;
    nor02ii ix149 (.Y (nx152), .A0 (nx358), .A1 (counter_out_12_rename)) ;
    xor2 ix143 (.Y (nx142), .A0 (nx353), .A1 (nx358)) ;
    nor02ii ix125 (.Y (nx155), .A0 (nx372), .A1 (counter_out_10_rename)) ;
    xor2 ix119 (.Y (nx118), .A0 (nx367), .A1 (nx372)) ;
    nor02ii ix101 (.Y (nx157), .A0 (nx386), .A1 (counter_out_8_rename)) ;
    xor2 ix95 (.Y (nx94), .A0 (nx381), .A1 (nx386)) ;
    nor02ii ix77 (.Y (nx159), .A0 (nx400), .A1 (counter_out_6_rename)) ;
    xor2 ix71 (.Y (nx70), .A0 (nx395), .A1 (nx400)) ;
    nor02ii ix53 (.Y (nx161), .A0 (nx414), .A1 (counter_out_4_rename)) ;
    or02 ix425 (.Y (nx424), .A0 (nx428), .A1 (nx436)) ;
    xnor2 ix174 (.Y (nx173), .A0 (nx436), .A1 (nx474)) ;
    and04 ix207 (.Y (nx206), .A0 (nx362), .A1 (nx367), .A2 (nx376), .A3 (nx381)
          ) ;
    and04 ix225 (.Y (nx224), .A0 (nx390), .A1 (nx395), .A2 (nx404), .A3 (nx458)
          ) ;
    xnor2 ix217 (.Y (nx458), .A0 (max_val_in[0]), .A1 (counter_out_dup0_0)) ;
    xor2 ix446 (.Y (nx445), .A0 (nx428), .A1 (max_val_in[1])) ;
    xor2 ix452 (.Y (nx451), .A0 (nx409), .A1 (max_val_in[4])) ;
    inv01 ix459 (.Y (nx460), .A (reset)) ;
    inv02 ix461 (.Y (nx462), .A (nx460)) ;
    inv02 ix463 (.Y (nx464), .A (nx460)) ;
    inv02 ix465 (.Y (nx466), .A (nx460)) ;
    inv01 ix467 (.Y (nx468), .A (enable)) ;
    inv02 ix469 (.Y (nx470), .A (nx468)) ;
    inv02 ix471 (.Y (nx472), .A (nx468)) ;
    inv02 ix473 (.Y (nx474), .A (nx468)) ;
endmodule


module Cache_5_16_28_5 ( in_word, cache_in_sel, cache_out_sel, decoder_enable, 
                         out_column_0__15, out_column_0__14, out_column_0__13, 
                         out_column_0__12, out_column_0__11, out_column_0__10, 
                         out_column_0__9, out_column_0__8, out_column_0__7, 
                         out_column_0__6, out_column_0__5, out_column_0__4, 
                         out_column_0__3, out_column_0__2, out_column_0__1, 
                         out_column_0__0, out_column_1__15, out_column_1__14, 
                         out_column_1__13, out_column_1__12, out_column_1__11, 
                         out_column_1__10, out_column_1__9, out_column_1__8, 
                         out_column_1__7, out_column_1__6, out_column_1__5, 
                         out_column_1__4, out_column_1__3, out_column_1__2, 
                         out_column_1__1, out_column_1__0, out_column_2__15, 
                         out_column_2__14, out_column_2__13, out_column_2__12, 
                         out_column_2__11, out_column_2__10, out_column_2__9, 
                         out_column_2__8, out_column_2__7, out_column_2__6, 
                         out_column_2__5, out_column_2__4, out_column_2__3, 
                         out_column_2__2, out_column_2__1, out_column_2__0, 
                         out_column_3__15, out_column_3__14, out_column_3__13, 
                         out_column_3__12, out_column_3__11, out_column_3__10, 
                         out_column_3__9, out_column_3__8, out_column_3__7, 
                         out_column_3__6, out_column_3__5, out_column_3__4, 
                         out_column_3__3, out_column_3__2, out_column_3__1, 
                         out_column_3__0, out_column_4__15, out_column_4__14, 
                         out_column_4__13, out_column_4__12, out_column_4__11, 
                         out_column_4__10, out_column_4__9, out_column_4__8, 
                         out_column_4__7, out_column_4__6, out_column_4__5, 
                         out_column_4__4, out_column_4__3, out_column_4__2, 
                         out_column_4__1, out_column_4__0, clk, reset ) ;

    input [15:0]in_word ;
    input [4:0]cache_in_sel ;
    input [4:0]cache_out_sel ;
    input decoder_enable ;
    output out_column_0__15 ;
    output out_column_0__14 ;
    output out_column_0__13 ;
    output out_column_0__12 ;
    output out_column_0__11 ;
    output out_column_0__10 ;
    output out_column_0__9 ;
    output out_column_0__8 ;
    output out_column_0__7 ;
    output out_column_0__6 ;
    output out_column_0__5 ;
    output out_column_0__4 ;
    output out_column_0__3 ;
    output out_column_0__2 ;
    output out_column_0__1 ;
    output out_column_0__0 ;
    output out_column_1__15 ;
    output out_column_1__14 ;
    output out_column_1__13 ;
    output out_column_1__12 ;
    output out_column_1__11 ;
    output out_column_1__10 ;
    output out_column_1__9 ;
    output out_column_1__8 ;
    output out_column_1__7 ;
    output out_column_1__6 ;
    output out_column_1__5 ;
    output out_column_1__4 ;
    output out_column_1__3 ;
    output out_column_1__2 ;
    output out_column_1__1 ;
    output out_column_1__0 ;
    output out_column_2__15 ;
    output out_column_2__14 ;
    output out_column_2__13 ;
    output out_column_2__12 ;
    output out_column_2__11 ;
    output out_column_2__10 ;
    output out_column_2__9 ;
    output out_column_2__8 ;
    output out_column_2__7 ;
    output out_column_2__6 ;
    output out_column_2__5 ;
    output out_column_2__4 ;
    output out_column_2__3 ;
    output out_column_2__2 ;
    output out_column_2__1 ;
    output out_column_2__0 ;
    output out_column_3__15 ;
    output out_column_3__14 ;
    output out_column_3__13 ;
    output out_column_3__12 ;
    output out_column_3__11 ;
    output out_column_3__10 ;
    output out_column_3__9 ;
    output out_column_3__8 ;
    output out_column_3__7 ;
    output out_column_3__6 ;
    output out_column_3__5 ;
    output out_column_3__4 ;
    output out_column_3__3 ;
    output out_column_3__2 ;
    output out_column_3__1 ;
    output out_column_3__0 ;
    output out_column_4__15 ;
    output out_column_4__14 ;
    output out_column_4__13 ;
    output out_column_4__12 ;
    output out_column_4__11 ;
    output out_column_4__10 ;
    output out_column_4__9 ;
    output out_column_4__8 ;
    output out_column_4__7 ;
    output out_column_4__6 ;
    output out_column_4__5 ;
    output out_column_4__4 ;
    output out_column_4__3 ;
    output out_column_4__2 ;
    output out_column_4__1 ;
    output out_column_4__0 ;
    input clk ;
    input reset ;

    wire que_out_0__0__15, que_out_0__0__14, que_out_0__0__13, que_out_0__0__12, 
         que_out_0__0__11, que_out_0__0__10, que_out_0__0__9, que_out_0__0__8, 
         que_out_0__0__7, que_out_0__0__6, que_out_0__0__5, que_out_0__0__4, 
         que_out_0__0__3, que_out_0__0__2, que_out_0__0__1, que_out_0__0__0, 
         que_out_0__1__15, que_out_0__1__14, que_out_0__1__13, que_out_0__1__12, 
         que_out_0__1__11, que_out_0__1__10, que_out_0__1__9, que_out_0__1__8, 
         que_out_0__1__7, que_out_0__1__6, que_out_0__1__5, que_out_0__1__4, 
         que_out_0__1__3, que_out_0__1__2, que_out_0__1__1, que_out_0__1__0, 
         que_out_0__2__15, que_out_0__2__14, que_out_0__2__13, que_out_0__2__12, 
         que_out_0__2__11, que_out_0__2__10, que_out_0__2__9, que_out_0__2__8, 
         que_out_0__2__7, que_out_0__2__6, que_out_0__2__5, que_out_0__2__4, 
         que_out_0__2__3, que_out_0__2__2, que_out_0__2__1, que_out_0__2__0, 
         que_out_0__3__15, que_out_0__3__14, que_out_0__3__13, que_out_0__3__12, 
         que_out_0__3__11, que_out_0__3__10, que_out_0__3__9, que_out_0__3__8, 
         que_out_0__3__7, que_out_0__3__6, que_out_0__3__5, que_out_0__3__4, 
         que_out_0__3__3, que_out_0__3__2, que_out_0__3__1, que_out_0__3__0, 
         que_out_0__4__15, que_out_0__4__14, que_out_0__4__13, que_out_0__4__12, 
         que_out_0__4__11, que_out_0__4__10, que_out_0__4__9, que_out_0__4__8, 
         que_out_0__4__7, que_out_0__4__6, que_out_0__4__5, que_out_0__4__4, 
         que_out_0__4__3, que_out_0__4__2, que_out_0__4__1, que_out_0__4__0, 
         que_out_1__0__15, que_out_1__0__14, que_out_1__0__13, que_out_1__0__12, 
         que_out_1__0__11, que_out_1__0__10, que_out_1__0__9, que_out_1__0__8, 
         que_out_1__0__7, que_out_1__0__6, que_out_1__0__5, que_out_1__0__4, 
         que_out_1__0__3, que_out_1__0__2, que_out_1__0__1, que_out_1__0__0, 
         que_out_1__1__15, que_out_1__1__14, que_out_1__1__13, que_out_1__1__12, 
         que_out_1__1__11, que_out_1__1__10, que_out_1__1__9, que_out_1__1__8, 
         que_out_1__1__7, que_out_1__1__6, que_out_1__1__5, que_out_1__1__4, 
         que_out_1__1__3, que_out_1__1__2, que_out_1__1__1, que_out_1__1__0, 
         que_out_1__2__15, que_out_1__2__14, que_out_1__2__13, que_out_1__2__12, 
         que_out_1__2__11, que_out_1__2__10, que_out_1__2__9, que_out_1__2__8, 
         que_out_1__2__7, que_out_1__2__6, que_out_1__2__5, que_out_1__2__4, 
         que_out_1__2__3, que_out_1__2__2, que_out_1__2__1, que_out_1__2__0, 
         que_out_1__3__15, que_out_1__3__14, que_out_1__3__13, que_out_1__3__12, 
         que_out_1__3__11, que_out_1__3__10, que_out_1__3__9, que_out_1__3__8, 
         que_out_1__3__7, que_out_1__3__6, que_out_1__3__5, que_out_1__3__4, 
         que_out_1__3__3, que_out_1__3__2, que_out_1__3__1, que_out_1__3__0, 
         que_out_1__4__15, que_out_1__4__14, que_out_1__4__13, que_out_1__4__12, 
         que_out_1__4__11, que_out_1__4__10, que_out_1__4__9, que_out_1__4__8, 
         que_out_1__4__7, que_out_1__4__6, que_out_1__4__5, que_out_1__4__4, 
         que_out_1__4__3, que_out_1__4__2, que_out_1__4__1, que_out_1__4__0, 
         que_out_2__0__15, que_out_2__0__14, que_out_2__0__13, que_out_2__0__12, 
         que_out_2__0__11, que_out_2__0__10, que_out_2__0__9, que_out_2__0__8, 
         que_out_2__0__7, que_out_2__0__6, que_out_2__0__5, que_out_2__0__4, 
         que_out_2__0__3, que_out_2__0__2, que_out_2__0__1, que_out_2__0__0, 
         que_out_2__1__15, que_out_2__1__14, que_out_2__1__13, que_out_2__1__12, 
         que_out_2__1__11, que_out_2__1__10, que_out_2__1__9, que_out_2__1__8, 
         que_out_2__1__7, que_out_2__1__6, que_out_2__1__5, que_out_2__1__4, 
         que_out_2__1__3, que_out_2__1__2, que_out_2__1__1, que_out_2__1__0, 
         que_out_2__2__15, que_out_2__2__14, que_out_2__2__13, que_out_2__2__12, 
         que_out_2__2__11, que_out_2__2__10, que_out_2__2__9, que_out_2__2__8, 
         que_out_2__2__7, que_out_2__2__6, que_out_2__2__5, que_out_2__2__4, 
         que_out_2__2__3, que_out_2__2__2, que_out_2__2__1, que_out_2__2__0, 
         que_out_2__3__15, que_out_2__3__14, que_out_2__3__13, que_out_2__3__12, 
         que_out_2__3__11, que_out_2__3__10, que_out_2__3__9, que_out_2__3__8, 
         que_out_2__3__7, que_out_2__3__6, que_out_2__3__5, que_out_2__3__4, 
         que_out_2__3__3, que_out_2__3__2, que_out_2__3__1, que_out_2__3__0, 
         que_out_2__4__15, que_out_2__4__14, que_out_2__4__13, que_out_2__4__12, 
         que_out_2__4__11, que_out_2__4__10, que_out_2__4__9, que_out_2__4__8, 
         que_out_2__4__7, que_out_2__4__6, que_out_2__4__5, que_out_2__4__4, 
         que_out_2__4__3, que_out_2__4__2, que_out_2__4__1, que_out_2__4__0, 
         que_out_3__0__15, que_out_3__0__14, que_out_3__0__13, que_out_3__0__12, 
         que_out_3__0__11, que_out_3__0__10, que_out_3__0__9, que_out_3__0__8, 
         que_out_3__0__7, que_out_3__0__6, que_out_3__0__5, que_out_3__0__4, 
         que_out_3__0__3, que_out_3__0__2, que_out_3__0__1, que_out_3__0__0, 
         que_out_3__1__15, que_out_3__1__14, que_out_3__1__13, que_out_3__1__12, 
         que_out_3__1__11, que_out_3__1__10, que_out_3__1__9, que_out_3__1__8, 
         que_out_3__1__7, que_out_3__1__6, que_out_3__1__5, que_out_3__1__4, 
         que_out_3__1__3, que_out_3__1__2, que_out_3__1__1, que_out_3__1__0, 
         que_out_3__2__15, que_out_3__2__14, que_out_3__2__13, que_out_3__2__12, 
         que_out_3__2__11, que_out_3__2__10, que_out_3__2__9, que_out_3__2__8, 
         que_out_3__2__7, que_out_3__2__6, que_out_3__2__5, que_out_3__2__4, 
         que_out_3__2__3, que_out_3__2__2, que_out_3__2__1, que_out_3__2__0, 
         que_out_3__3__15, que_out_3__3__14, que_out_3__3__13, que_out_3__3__12, 
         que_out_3__3__11, que_out_3__3__10, que_out_3__3__9, que_out_3__3__8, 
         que_out_3__3__7, que_out_3__3__6, que_out_3__3__5, que_out_3__3__4, 
         que_out_3__3__3, que_out_3__3__2, que_out_3__3__1, que_out_3__3__0, 
         que_out_3__4__15, que_out_3__4__14, que_out_3__4__13, que_out_3__4__12, 
         que_out_3__4__11, que_out_3__4__10, que_out_3__4__9, que_out_3__4__8, 
         que_out_3__4__7, que_out_3__4__6, que_out_3__4__5, que_out_3__4__4, 
         que_out_3__4__3, que_out_3__4__2, que_out_3__4__1, que_out_3__4__0, 
         que_out_4__0__15, que_out_4__0__14, que_out_4__0__13, que_out_4__0__12, 
         que_out_4__0__11, que_out_4__0__10, que_out_4__0__9, que_out_4__0__8, 
         que_out_4__0__7, que_out_4__0__6, que_out_4__0__5, que_out_4__0__4, 
         que_out_4__0__3, que_out_4__0__2, que_out_4__0__1, que_out_4__0__0, 
         que_out_4__1__15, que_out_4__1__14, que_out_4__1__13, que_out_4__1__12, 
         que_out_4__1__11, que_out_4__1__10, que_out_4__1__9, que_out_4__1__8, 
         que_out_4__1__7, que_out_4__1__6, que_out_4__1__5, que_out_4__1__4, 
         que_out_4__1__3, que_out_4__1__2, que_out_4__1__1, que_out_4__1__0, 
         que_out_4__2__15, que_out_4__2__14, que_out_4__2__13, que_out_4__2__12, 
         que_out_4__2__11, que_out_4__2__10, que_out_4__2__9, que_out_4__2__8, 
         que_out_4__2__7, que_out_4__2__6, que_out_4__2__5, que_out_4__2__4, 
         que_out_4__2__3, que_out_4__2__2, que_out_4__2__1, que_out_4__2__0, 
         que_out_4__3__15, que_out_4__3__14, que_out_4__3__13, que_out_4__3__12, 
         que_out_4__3__11, que_out_4__3__10, que_out_4__3__9, que_out_4__3__8, 
         que_out_4__3__7, que_out_4__3__6, que_out_4__3__5, que_out_4__3__4, 
         que_out_4__3__3, que_out_4__3__2, que_out_4__3__1, que_out_4__3__0, 
         que_out_4__4__15, que_out_4__4__14, que_out_4__4__13, que_out_4__4__12, 
         que_out_4__4__11, que_out_4__4__10, que_out_4__4__9, que_out_4__4__8, 
         que_out_4__4__7, que_out_4__4__6, que_out_4__4__5, que_out_4__4__4, 
         que_out_4__4__3, que_out_4__4__2, que_out_4__4__1, que_out_4__4__0, 
         que_out_5__0__15, que_out_5__0__14, que_out_5__0__13, que_out_5__0__12, 
         que_out_5__0__11, que_out_5__0__10, que_out_5__0__9, que_out_5__0__8, 
         que_out_5__0__7, que_out_5__0__6, que_out_5__0__5, que_out_5__0__4, 
         que_out_5__0__3, que_out_5__0__2, que_out_5__0__1, que_out_5__0__0, 
         que_out_5__1__15, que_out_5__1__14, que_out_5__1__13, que_out_5__1__12, 
         que_out_5__1__11, que_out_5__1__10, que_out_5__1__9, que_out_5__1__8, 
         que_out_5__1__7, que_out_5__1__6, que_out_5__1__5, que_out_5__1__4, 
         que_out_5__1__3, que_out_5__1__2, que_out_5__1__1, que_out_5__1__0, 
         que_out_5__2__15, que_out_5__2__14, que_out_5__2__13, que_out_5__2__12, 
         que_out_5__2__11, que_out_5__2__10, que_out_5__2__9, que_out_5__2__8, 
         que_out_5__2__7, que_out_5__2__6, que_out_5__2__5, que_out_5__2__4, 
         que_out_5__2__3, que_out_5__2__2, que_out_5__2__1, que_out_5__2__0, 
         que_out_5__3__15, que_out_5__3__14, que_out_5__3__13, que_out_5__3__12, 
         que_out_5__3__11, que_out_5__3__10, que_out_5__3__9, que_out_5__3__8, 
         que_out_5__3__7, que_out_5__3__6, que_out_5__3__5, que_out_5__3__4, 
         que_out_5__3__3, que_out_5__3__2, que_out_5__3__1, que_out_5__3__0, 
         que_out_5__4__15, que_out_5__4__14, que_out_5__4__13, que_out_5__4__12, 
         que_out_5__4__11, que_out_5__4__10, que_out_5__4__9, que_out_5__4__8, 
         que_out_5__4__7, que_out_5__4__6, que_out_5__4__5, que_out_5__4__4, 
         que_out_5__4__3, que_out_5__4__2, que_out_5__4__1, que_out_5__4__0, 
         que_out_6__0__15, que_out_6__0__14, que_out_6__0__13, que_out_6__0__12, 
         que_out_6__0__11, que_out_6__0__10, que_out_6__0__9, que_out_6__0__8, 
         que_out_6__0__7, que_out_6__0__6, que_out_6__0__5, que_out_6__0__4, 
         que_out_6__0__3, que_out_6__0__2, que_out_6__0__1, que_out_6__0__0, 
         que_out_6__1__15, que_out_6__1__14, que_out_6__1__13, que_out_6__1__12, 
         que_out_6__1__11, que_out_6__1__10, que_out_6__1__9, que_out_6__1__8, 
         que_out_6__1__7, que_out_6__1__6, que_out_6__1__5, que_out_6__1__4, 
         que_out_6__1__3, que_out_6__1__2, que_out_6__1__1, que_out_6__1__0, 
         que_out_6__2__15, que_out_6__2__14, que_out_6__2__13, que_out_6__2__12, 
         que_out_6__2__11, que_out_6__2__10, que_out_6__2__9, que_out_6__2__8, 
         que_out_6__2__7, que_out_6__2__6, que_out_6__2__5, que_out_6__2__4, 
         que_out_6__2__3, que_out_6__2__2, que_out_6__2__1, que_out_6__2__0, 
         que_out_6__3__15, que_out_6__3__14, que_out_6__3__13, que_out_6__3__12, 
         que_out_6__3__11, que_out_6__3__10, que_out_6__3__9, que_out_6__3__8, 
         que_out_6__3__7, que_out_6__3__6, que_out_6__3__5, que_out_6__3__4, 
         que_out_6__3__3, que_out_6__3__2, que_out_6__3__1, que_out_6__3__0, 
         que_out_6__4__15, que_out_6__4__14, que_out_6__4__13, que_out_6__4__12, 
         que_out_6__4__11, que_out_6__4__10, que_out_6__4__9, que_out_6__4__8, 
         que_out_6__4__7, que_out_6__4__6, que_out_6__4__5, que_out_6__4__4, 
         que_out_6__4__3, que_out_6__4__2, que_out_6__4__1, que_out_6__4__0, 
         que_out_7__0__15, que_out_7__0__14, que_out_7__0__13, que_out_7__0__12, 
         que_out_7__0__11, que_out_7__0__10, que_out_7__0__9, que_out_7__0__8, 
         que_out_7__0__7, que_out_7__0__6, que_out_7__0__5, que_out_7__0__4, 
         que_out_7__0__3, que_out_7__0__2, que_out_7__0__1, que_out_7__0__0, 
         que_out_7__1__15, que_out_7__1__14, que_out_7__1__13, que_out_7__1__12, 
         que_out_7__1__11, que_out_7__1__10, que_out_7__1__9, que_out_7__1__8, 
         que_out_7__1__7, que_out_7__1__6, que_out_7__1__5, que_out_7__1__4, 
         que_out_7__1__3, que_out_7__1__2, que_out_7__1__1, que_out_7__1__0, 
         que_out_7__2__15, que_out_7__2__14, que_out_7__2__13, que_out_7__2__12, 
         que_out_7__2__11, que_out_7__2__10, que_out_7__2__9, que_out_7__2__8, 
         que_out_7__2__7, que_out_7__2__6, que_out_7__2__5, que_out_7__2__4, 
         que_out_7__2__3, que_out_7__2__2, que_out_7__2__1, que_out_7__2__0, 
         que_out_7__3__15, que_out_7__3__14, que_out_7__3__13, que_out_7__3__12, 
         que_out_7__3__11, que_out_7__3__10, que_out_7__3__9, que_out_7__3__8, 
         que_out_7__3__7, que_out_7__3__6, que_out_7__3__5, que_out_7__3__4, 
         que_out_7__3__3, que_out_7__3__2, que_out_7__3__1, que_out_7__3__0, 
         que_out_7__4__15, que_out_7__4__14, que_out_7__4__13, que_out_7__4__12, 
         que_out_7__4__11, que_out_7__4__10, que_out_7__4__9, que_out_7__4__8, 
         que_out_7__4__7, que_out_7__4__6, que_out_7__4__5, que_out_7__4__4, 
         que_out_7__4__3, que_out_7__4__2, que_out_7__4__1, que_out_7__4__0, 
         que_out_8__0__15, que_out_8__0__14, que_out_8__0__13, que_out_8__0__12, 
         que_out_8__0__11, que_out_8__0__10, que_out_8__0__9, que_out_8__0__8, 
         que_out_8__0__7, que_out_8__0__6, que_out_8__0__5, que_out_8__0__4, 
         que_out_8__0__3, que_out_8__0__2, que_out_8__0__1, que_out_8__0__0, 
         que_out_8__1__15, que_out_8__1__14, que_out_8__1__13, que_out_8__1__12, 
         que_out_8__1__11, que_out_8__1__10, que_out_8__1__9, que_out_8__1__8, 
         que_out_8__1__7, que_out_8__1__6, que_out_8__1__5, que_out_8__1__4, 
         que_out_8__1__3, que_out_8__1__2, que_out_8__1__1, que_out_8__1__0, 
         que_out_8__2__15, que_out_8__2__14, que_out_8__2__13, que_out_8__2__12, 
         que_out_8__2__11, que_out_8__2__10, que_out_8__2__9, que_out_8__2__8, 
         que_out_8__2__7, que_out_8__2__6, que_out_8__2__5, que_out_8__2__4, 
         que_out_8__2__3, que_out_8__2__2, que_out_8__2__1, que_out_8__2__0, 
         que_out_8__3__15, que_out_8__3__14, que_out_8__3__13, que_out_8__3__12, 
         que_out_8__3__11, que_out_8__3__10, que_out_8__3__9, que_out_8__3__8, 
         que_out_8__3__7, que_out_8__3__6, que_out_8__3__5, que_out_8__3__4, 
         que_out_8__3__3, que_out_8__3__2, que_out_8__3__1, que_out_8__3__0, 
         que_out_8__4__15, que_out_8__4__14, que_out_8__4__13, que_out_8__4__12, 
         que_out_8__4__11, que_out_8__4__10, que_out_8__4__9, que_out_8__4__8, 
         que_out_8__4__7, que_out_8__4__6, que_out_8__4__5, que_out_8__4__4, 
         que_out_8__4__3, que_out_8__4__2, que_out_8__4__1, que_out_8__4__0, 
         que_out_9__0__15, que_out_9__0__14, que_out_9__0__13, que_out_9__0__12, 
         que_out_9__0__11, que_out_9__0__10, que_out_9__0__9, que_out_9__0__8, 
         que_out_9__0__7, que_out_9__0__6, que_out_9__0__5, que_out_9__0__4, 
         que_out_9__0__3, que_out_9__0__2, que_out_9__0__1, que_out_9__0__0, 
         que_out_9__1__15, que_out_9__1__14, que_out_9__1__13, que_out_9__1__12, 
         que_out_9__1__11, que_out_9__1__10, que_out_9__1__9, que_out_9__1__8, 
         que_out_9__1__7, que_out_9__1__6, que_out_9__1__5, que_out_9__1__4, 
         que_out_9__1__3, que_out_9__1__2, que_out_9__1__1, que_out_9__1__0, 
         que_out_9__2__15, que_out_9__2__14, que_out_9__2__13, que_out_9__2__12, 
         que_out_9__2__11, que_out_9__2__10, que_out_9__2__9, que_out_9__2__8, 
         que_out_9__2__7, que_out_9__2__6, que_out_9__2__5, que_out_9__2__4, 
         que_out_9__2__3, que_out_9__2__2, que_out_9__2__1, que_out_9__2__0, 
         que_out_9__3__15, que_out_9__3__14, que_out_9__3__13, que_out_9__3__12, 
         que_out_9__3__11, que_out_9__3__10, que_out_9__3__9, que_out_9__3__8, 
         que_out_9__3__7, que_out_9__3__6, que_out_9__3__5, que_out_9__3__4, 
         que_out_9__3__3, que_out_9__3__2, que_out_9__3__1, que_out_9__3__0, 
         que_out_9__4__15, que_out_9__4__14, que_out_9__4__13, que_out_9__4__12, 
         que_out_9__4__11, que_out_9__4__10, que_out_9__4__9, que_out_9__4__8, 
         que_out_9__4__7, que_out_9__4__6, que_out_9__4__5, que_out_9__4__4, 
         que_out_9__4__3, que_out_9__4__2, que_out_9__4__1, que_out_9__4__0, 
         que_out_10__0__15, que_out_10__0__14, que_out_10__0__13, 
         que_out_10__0__12, que_out_10__0__11, que_out_10__0__10, 
         que_out_10__0__9, que_out_10__0__8, que_out_10__0__7, que_out_10__0__6, 
         que_out_10__0__5, que_out_10__0__4, que_out_10__0__3, que_out_10__0__2, 
         que_out_10__0__1, que_out_10__0__0, que_out_10__1__15, 
         que_out_10__1__14, que_out_10__1__13, que_out_10__1__12, 
         que_out_10__1__11, que_out_10__1__10, que_out_10__1__9, 
         que_out_10__1__8, que_out_10__1__7, que_out_10__1__6, que_out_10__1__5, 
         que_out_10__1__4, que_out_10__1__3, que_out_10__1__2, que_out_10__1__1, 
         que_out_10__1__0, que_out_10__2__15, que_out_10__2__14, 
         que_out_10__2__13, que_out_10__2__12, que_out_10__2__11, 
         que_out_10__2__10, que_out_10__2__9, que_out_10__2__8, que_out_10__2__7, 
         que_out_10__2__6, que_out_10__2__5, que_out_10__2__4, que_out_10__2__3, 
         que_out_10__2__2, que_out_10__2__1, que_out_10__2__0, que_out_10__3__15, 
         que_out_10__3__14, que_out_10__3__13, que_out_10__3__12, 
         que_out_10__3__11, que_out_10__3__10, que_out_10__3__9, 
         que_out_10__3__8, que_out_10__3__7, que_out_10__3__6, que_out_10__3__5, 
         que_out_10__3__4, que_out_10__3__3, que_out_10__3__2, que_out_10__3__1, 
         que_out_10__3__0, que_out_10__4__15, que_out_10__4__14, 
         que_out_10__4__13, que_out_10__4__12, que_out_10__4__11, 
         que_out_10__4__10, que_out_10__4__9, que_out_10__4__8, que_out_10__4__7, 
         que_out_10__4__6, que_out_10__4__5, que_out_10__4__4, que_out_10__4__3, 
         que_out_10__4__2, que_out_10__4__1, que_out_10__4__0, que_out_11__0__15, 
         que_out_11__0__14, que_out_11__0__13, que_out_11__0__12, 
         que_out_11__0__11, que_out_11__0__10, que_out_11__0__9, 
         que_out_11__0__8, que_out_11__0__7, que_out_11__0__6, que_out_11__0__5, 
         que_out_11__0__4, que_out_11__0__3, que_out_11__0__2, que_out_11__0__1, 
         que_out_11__0__0, que_out_11__1__15, que_out_11__1__14, 
         que_out_11__1__13, que_out_11__1__12, que_out_11__1__11, 
         que_out_11__1__10, que_out_11__1__9, que_out_11__1__8, que_out_11__1__7, 
         que_out_11__1__6, que_out_11__1__5, que_out_11__1__4, que_out_11__1__3, 
         que_out_11__1__2, que_out_11__1__1, que_out_11__1__0, que_out_11__2__15, 
         que_out_11__2__14, que_out_11__2__13, que_out_11__2__12, 
         que_out_11__2__11, que_out_11__2__10, que_out_11__2__9, 
         que_out_11__2__8, que_out_11__2__7, que_out_11__2__6, que_out_11__2__5, 
         que_out_11__2__4, que_out_11__2__3, que_out_11__2__2, que_out_11__2__1, 
         que_out_11__2__0, que_out_11__3__15, que_out_11__3__14, 
         que_out_11__3__13, que_out_11__3__12, que_out_11__3__11, 
         que_out_11__3__10, que_out_11__3__9, que_out_11__3__8, que_out_11__3__7, 
         que_out_11__3__6, que_out_11__3__5, que_out_11__3__4, que_out_11__3__3, 
         que_out_11__3__2, que_out_11__3__1, que_out_11__3__0, que_out_11__4__15, 
         que_out_11__4__14, que_out_11__4__13, que_out_11__4__12, 
         que_out_11__4__11, que_out_11__4__10, que_out_11__4__9, 
         que_out_11__4__8, que_out_11__4__7, que_out_11__4__6, que_out_11__4__5, 
         que_out_11__4__4, que_out_11__4__3, que_out_11__4__2, que_out_11__4__1, 
         que_out_11__4__0, que_out_12__0__15, que_out_12__0__14, 
         que_out_12__0__13, que_out_12__0__12, que_out_12__0__11, 
         que_out_12__0__10, que_out_12__0__9, que_out_12__0__8, que_out_12__0__7, 
         que_out_12__0__6, que_out_12__0__5, que_out_12__0__4, que_out_12__0__3, 
         que_out_12__0__2, que_out_12__0__1, que_out_12__0__0, que_out_12__1__15, 
         que_out_12__1__14, que_out_12__1__13, que_out_12__1__12, 
         que_out_12__1__11, que_out_12__1__10, que_out_12__1__9, 
         que_out_12__1__8, que_out_12__1__7, que_out_12__1__6, que_out_12__1__5, 
         que_out_12__1__4, que_out_12__1__3, que_out_12__1__2, que_out_12__1__1, 
         que_out_12__1__0, que_out_12__2__15, que_out_12__2__14, 
         que_out_12__2__13, que_out_12__2__12, que_out_12__2__11, 
         que_out_12__2__10, que_out_12__2__9, que_out_12__2__8, que_out_12__2__7, 
         que_out_12__2__6, que_out_12__2__5, que_out_12__2__4, que_out_12__2__3, 
         que_out_12__2__2, que_out_12__2__1, que_out_12__2__0, que_out_12__3__15, 
         que_out_12__3__14, que_out_12__3__13, que_out_12__3__12, 
         que_out_12__3__11, que_out_12__3__10, que_out_12__3__9, 
         que_out_12__3__8, que_out_12__3__7, que_out_12__3__6, que_out_12__3__5, 
         que_out_12__3__4, que_out_12__3__3, que_out_12__3__2, que_out_12__3__1, 
         que_out_12__3__0, que_out_12__4__15, que_out_12__4__14, 
         que_out_12__4__13, que_out_12__4__12, que_out_12__4__11, 
         que_out_12__4__10, que_out_12__4__9, que_out_12__4__8, que_out_12__4__7, 
         que_out_12__4__6, que_out_12__4__5, que_out_12__4__4, que_out_12__4__3, 
         que_out_12__4__2, que_out_12__4__1, que_out_12__4__0, que_out_13__0__15, 
         que_out_13__0__14, que_out_13__0__13, que_out_13__0__12, 
         que_out_13__0__11, que_out_13__0__10, que_out_13__0__9, 
         que_out_13__0__8, que_out_13__0__7, que_out_13__0__6, que_out_13__0__5, 
         que_out_13__0__4, que_out_13__0__3, que_out_13__0__2, que_out_13__0__1, 
         que_out_13__0__0, que_out_13__1__15, que_out_13__1__14, 
         que_out_13__1__13, que_out_13__1__12, que_out_13__1__11, 
         que_out_13__1__10, que_out_13__1__9, que_out_13__1__8, que_out_13__1__7, 
         que_out_13__1__6, que_out_13__1__5, que_out_13__1__4, que_out_13__1__3, 
         que_out_13__1__2, que_out_13__1__1, que_out_13__1__0, que_out_13__2__15, 
         que_out_13__2__14, que_out_13__2__13, que_out_13__2__12, 
         que_out_13__2__11, que_out_13__2__10, que_out_13__2__9, 
         que_out_13__2__8, que_out_13__2__7, que_out_13__2__6, que_out_13__2__5, 
         que_out_13__2__4, que_out_13__2__3, que_out_13__2__2, que_out_13__2__1, 
         que_out_13__2__0, que_out_13__3__15, que_out_13__3__14, 
         que_out_13__3__13, que_out_13__3__12, que_out_13__3__11, 
         que_out_13__3__10, que_out_13__3__9, que_out_13__3__8, que_out_13__3__7, 
         que_out_13__3__6, que_out_13__3__5, que_out_13__3__4, que_out_13__3__3, 
         que_out_13__3__2, que_out_13__3__1, que_out_13__3__0, que_out_13__4__15, 
         que_out_13__4__14, que_out_13__4__13, que_out_13__4__12, 
         que_out_13__4__11, que_out_13__4__10, que_out_13__4__9, 
         que_out_13__4__8, que_out_13__4__7, que_out_13__4__6, que_out_13__4__5, 
         que_out_13__4__4, que_out_13__4__3, que_out_13__4__2, que_out_13__4__1, 
         que_out_13__4__0, que_out_14__0__15, que_out_14__0__14, 
         que_out_14__0__13, que_out_14__0__12, que_out_14__0__11, 
         que_out_14__0__10, que_out_14__0__9, que_out_14__0__8, que_out_14__0__7, 
         que_out_14__0__6, que_out_14__0__5, que_out_14__0__4, que_out_14__0__3, 
         que_out_14__0__2, que_out_14__0__1, que_out_14__0__0, que_out_14__1__15, 
         que_out_14__1__14, que_out_14__1__13, que_out_14__1__12, 
         que_out_14__1__11, que_out_14__1__10, que_out_14__1__9, 
         que_out_14__1__8, que_out_14__1__7, que_out_14__1__6, que_out_14__1__5, 
         que_out_14__1__4, que_out_14__1__3, que_out_14__1__2, que_out_14__1__1, 
         que_out_14__1__0, que_out_14__2__15, que_out_14__2__14, 
         que_out_14__2__13, que_out_14__2__12, que_out_14__2__11, 
         que_out_14__2__10, que_out_14__2__9, que_out_14__2__8, que_out_14__2__7, 
         que_out_14__2__6, que_out_14__2__5, que_out_14__2__4, que_out_14__2__3, 
         que_out_14__2__2, que_out_14__2__1, que_out_14__2__0, que_out_14__3__15, 
         que_out_14__3__14, que_out_14__3__13, que_out_14__3__12, 
         que_out_14__3__11, que_out_14__3__10, que_out_14__3__9, 
         que_out_14__3__8, que_out_14__3__7, que_out_14__3__6, que_out_14__3__5, 
         que_out_14__3__4, que_out_14__3__3, que_out_14__3__2, que_out_14__3__1, 
         que_out_14__3__0, que_out_14__4__15, que_out_14__4__14, 
         que_out_14__4__13, que_out_14__4__12, que_out_14__4__11, 
         que_out_14__4__10, que_out_14__4__9, que_out_14__4__8, que_out_14__4__7, 
         que_out_14__4__6, que_out_14__4__5, que_out_14__4__4, que_out_14__4__3, 
         que_out_14__4__2, que_out_14__4__1, que_out_14__4__0, que_out_15__0__15, 
         que_out_15__0__14, que_out_15__0__13, que_out_15__0__12, 
         que_out_15__0__11, que_out_15__0__10, que_out_15__0__9, 
         que_out_15__0__8, que_out_15__0__7, que_out_15__0__6, que_out_15__0__5, 
         que_out_15__0__4, que_out_15__0__3, que_out_15__0__2, que_out_15__0__1, 
         que_out_15__0__0, que_out_15__1__15, que_out_15__1__14, 
         que_out_15__1__13, que_out_15__1__12, que_out_15__1__11, 
         que_out_15__1__10, que_out_15__1__9, que_out_15__1__8, que_out_15__1__7, 
         que_out_15__1__6, que_out_15__1__5, que_out_15__1__4, que_out_15__1__3, 
         que_out_15__1__2, que_out_15__1__1, que_out_15__1__0, que_out_15__2__15, 
         que_out_15__2__14, que_out_15__2__13, que_out_15__2__12, 
         que_out_15__2__11, que_out_15__2__10, que_out_15__2__9, 
         que_out_15__2__8, que_out_15__2__7, que_out_15__2__6, que_out_15__2__5, 
         que_out_15__2__4, que_out_15__2__3, que_out_15__2__2, que_out_15__2__1, 
         que_out_15__2__0, que_out_15__3__15, que_out_15__3__14, 
         que_out_15__3__13, que_out_15__3__12, que_out_15__3__11, 
         que_out_15__3__10, que_out_15__3__9, que_out_15__3__8, que_out_15__3__7, 
         que_out_15__3__6, que_out_15__3__5, que_out_15__3__4, que_out_15__3__3, 
         que_out_15__3__2, que_out_15__3__1, que_out_15__3__0, que_out_15__4__15, 
         que_out_15__4__14, que_out_15__4__13, que_out_15__4__12, 
         que_out_15__4__11, que_out_15__4__10, que_out_15__4__9, 
         que_out_15__4__8, que_out_15__4__7, que_out_15__4__6, que_out_15__4__5, 
         que_out_15__4__4, que_out_15__4__3, que_out_15__4__2, que_out_15__4__1, 
         que_out_15__4__0, que_out_16__0__15, que_out_16__0__14, 
         que_out_16__0__13, que_out_16__0__12, que_out_16__0__11, 
         que_out_16__0__10, que_out_16__0__9, que_out_16__0__8, que_out_16__0__7, 
         que_out_16__0__6, que_out_16__0__5, que_out_16__0__4, que_out_16__0__3, 
         que_out_16__0__2, que_out_16__0__1, que_out_16__0__0, que_out_16__1__15, 
         que_out_16__1__14, que_out_16__1__13, que_out_16__1__12, 
         que_out_16__1__11, que_out_16__1__10, que_out_16__1__9, 
         que_out_16__1__8, que_out_16__1__7, que_out_16__1__6, que_out_16__1__5, 
         que_out_16__1__4, que_out_16__1__3, que_out_16__1__2, que_out_16__1__1, 
         que_out_16__1__0, que_out_16__2__15, que_out_16__2__14, 
         que_out_16__2__13, que_out_16__2__12, que_out_16__2__11, 
         que_out_16__2__10, que_out_16__2__9, que_out_16__2__8, que_out_16__2__7, 
         que_out_16__2__6, que_out_16__2__5, que_out_16__2__4, que_out_16__2__3, 
         que_out_16__2__2, que_out_16__2__1, que_out_16__2__0, que_out_16__3__15, 
         que_out_16__3__14, que_out_16__3__13, que_out_16__3__12, 
         que_out_16__3__11, que_out_16__3__10, que_out_16__3__9, 
         que_out_16__3__8, que_out_16__3__7, que_out_16__3__6, que_out_16__3__5, 
         que_out_16__3__4, que_out_16__3__3, que_out_16__3__2, que_out_16__3__1, 
         que_out_16__3__0, que_out_16__4__15, que_out_16__4__14, 
         que_out_16__4__13, que_out_16__4__12, que_out_16__4__11, 
         que_out_16__4__10, que_out_16__4__9, que_out_16__4__8, que_out_16__4__7, 
         que_out_16__4__6, que_out_16__4__5, que_out_16__4__4, que_out_16__4__3, 
         que_out_16__4__2, que_out_16__4__1, que_out_16__4__0, que_out_17__0__15, 
         que_out_17__0__14, que_out_17__0__13, que_out_17__0__12, 
         que_out_17__0__11, que_out_17__0__10, que_out_17__0__9, 
         que_out_17__0__8, que_out_17__0__7, que_out_17__0__6, que_out_17__0__5, 
         que_out_17__0__4, que_out_17__0__3, que_out_17__0__2, que_out_17__0__1, 
         que_out_17__0__0, que_out_17__1__15, que_out_17__1__14, 
         que_out_17__1__13, que_out_17__1__12, que_out_17__1__11, 
         que_out_17__1__10, que_out_17__1__9, que_out_17__1__8, que_out_17__1__7, 
         que_out_17__1__6, que_out_17__1__5, que_out_17__1__4, que_out_17__1__3, 
         que_out_17__1__2, que_out_17__1__1, que_out_17__1__0, que_out_17__2__15, 
         que_out_17__2__14, que_out_17__2__13, que_out_17__2__12, 
         que_out_17__2__11, que_out_17__2__10, que_out_17__2__9, 
         que_out_17__2__8, que_out_17__2__7, que_out_17__2__6, que_out_17__2__5, 
         que_out_17__2__4, que_out_17__2__3, que_out_17__2__2, que_out_17__2__1, 
         que_out_17__2__0, que_out_17__3__15, que_out_17__3__14, 
         que_out_17__3__13, que_out_17__3__12, que_out_17__3__11, 
         que_out_17__3__10, que_out_17__3__9, que_out_17__3__8, que_out_17__3__7, 
         que_out_17__3__6, que_out_17__3__5, que_out_17__3__4, que_out_17__3__3, 
         que_out_17__3__2, que_out_17__3__1, que_out_17__3__0, que_out_17__4__15, 
         que_out_17__4__14, que_out_17__4__13, que_out_17__4__12, 
         que_out_17__4__11, que_out_17__4__10, que_out_17__4__9, 
         que_out_17__4__8, que_out_17__4__7, que_out_17__4__6, que_out_17__4__5, 
         que_out_17__4__4, que_out_17__4__3, que_out_17__4__2, que_out_17__4__1, 
         que_out_17__4__0, que_out_18__0__15, que_out_18__0__14, 
         que_out_18__0__13, que_out_18__0__12, que_out_18__0__11, 
         que_out_18__0__10, que_out_18__0__9, que_out_18__0__8, que_out_18__0__7, 
         que_out_18__0__6, que_out_18__0__5, que_out_18__0__4, que_out_18__0__3, 
         que_out_18__0__2, que_out_18__0__1, que_out_18__0__0, que_out_18__1__15, 
         que_out_18__1__14, que_out_18__1__13, que_out_18__1__12, 
         que_out_18__1__11, que_out_18__1__10, que_out_18__1__9, 
         que_out_18__1__8, que_out_18__1__7, que_out_18__1__6, que_out_18__1__5, 
         que_out_18__1__4, que_out_18__1__3, que_out_18__1__2, que_out_18__1__1, 
         que_out_18__1__0, que_out_18__2__15, que_out_18__2__14, 
         que_out_18__2__13, que_out_18__2__12, que_out_18__2__11, 
         que_out_18__2__10, que_out_18__2__9, que_out_18__2__8, que_out_18__2__7, 
         que_out_18__2__6, que_out_18__2__5, que_out_18__2__4, que_out_18__2__3, 
         que_out_18__2__2, que_out_18__2__1, que_out_18__2__0, que_out_18__3__15, 
         que_out_18__3__14, que_out_18__3__13, que_out_18__3__12, 
         que_out_18__3__11, que_out_18__3__10, que_out_18__3__9, 
         que_out_18__3__8, que_out_18__3__7, que_out_18__3__6, que_out_18__3__5, 
         que_out_18__3__4, que_out_18__3__3, que_out_18__3__2, que_out_18__3__1, 
         que_out_18__3__0, que_out_18__4__15, que_out_18__4__14, 
         que_out_18__4__13, que_out_18__4__12, que_out_18__4__11, 
         que_out_18__4__10, que_out_18__4__9, que_out_18__4__8, que_out_18__4__7, 
         que_out_18__4__6, que_out_18__4__5, que_out_18__4__4, que_out_18__4__3, 
         que_out_18__4__2, que_out_18__4__1, que_out_18__4__0, que_out_19__0__15, 
         que_out_19__0__14, que_out_19__0__13, que_out_19__0__12, 
         que_out_19__0__11, que_out_19__0__10, que_out_19__0__9, 
         que_out_19__0__8, que_out_19__0__7, que_out_19__0__6, que_out_19__0__5, 
         que_out_19__0__4, que_out_19__0__3, que_out_19__0__2, que_out_19__0__1, 
         que_out_19__0__0, que_out_19__1__15, que_out_19__1__14, 
         que_out_19__1__13, que_out_19__1__12, que_out_19__1__11, 
         que_out_19__1__10, que_out_19__1__9, que_out_19__1__8, que_out_19__1__7, 
         que_out_19__1__6, que_out_19__1__5, que_out_19__1__4, que_out_19__1__3, 
         que_out_19__1__2, que_out_19__1__1, que_out_19__1__0, que_out_19__2__15, 
         que_out_19__2__14, que_out_19__2__13, que_out_19__2__12, 
         que_out_19__2__11, que_out_19__2__10, que_out_19__2__9, 
         que_out_19__2__8, que_out_19__2__7, que_out_19__2__6, que_out_19__2__5, 
         que_out_19__2__4, que_out_19__2__3, que_out_19__2__2, que_out_19__2__1, 
         que_out_19__2__0, que_out_19__3__15, que_out_19__3__14, 
         que_out_19__3__13, que_out_19__3__12, que_out_19__3__11, 
         que_out_19__3__10, que_out_19__3__9, que_out_19__3__8, que_out_19__3__7, 
         que_out_19__3__6, que_out_19__3__5, que_out_19__3__4, que_out_19__3__3, 
         que_out_19__3__2, que_out_19__3__1, que_out_19__3__0, que_out_19__4__15, 
         que_out_19__4__14, que_out_19__4__13, que_out_19__4__12, 
         que_out_19__4__11, que_out_19__4__10, que_out_19__4__9, 
         que_out_19__4__8, que_out_19__4__7, que_out_19__4__6, que_out_19__4__5, 
         que_out_19__4__4, que_out_19__4__3, que_out_19__4__2, que_out_19__4__1, 
         que_out_19__4__0, que_out_20__0__15, que_out_20__0__14, 
         que_out_20__0__13, que_out_20__0__12, que_out_20__0__11, 
         que_out_20__0__10, que_out_20__0__9, que_out_20__0__8, que_out_20__0__7, 
         que_out_20__0__6, que_out_20__0__5, que_out_20__0__4, que_out_20__0__3, 
         que_out_20__0__2, que_out_20__0__1, que_out_20__0__0, que_out_20__1__15, 
         que_out_20__1__14, que_out_20__1__13, que_out_20__1__12, 
         que_out_20__1__11, que_out_20__1__10, que_out_20__1__9, 
         que_out_20__1__8, que_out_20__1__7, que_out_20__1__6, que_out_20__1__5, 
         que_out_20__1__4, que_out_20__1__3, que_out_20__1__2, que_out_20__1__1, 
         que_out_20__1__0, que_out_20__2__15, que_out_20__2__14, 
         que_out_20__2__13, que_out_20__2__12, que_out_20__2__11, 
         que_out_20__2__10, que_out_20__2__9, que_out_20__2__8, que_out_20__2__7, 
         que_out_20__2__6, que_out_20__2__5, que_out_20__2__4, que_out_20__2__3, 
         que_out_20__2__2, que_out_20__2__1, que_out_20__2__0, que_out_20__3__15, 
         que_out_20__3__14, que_out_20__3__13, que_out_20__3__12, 
         que_out_20__3__11, que_out_20__3__10, que_out_20__3__9, 
         que_out_20__3__8, que_out_20__3__7, que_out_20__3__6, que_out_20__3__5, 
         que_out_20__3__4, que_out_20__3__3, que_out_20__3__2, que_out_20__3__1, 
         que_out_20__3__0, que_out_20__4__15, que_out_20__4__14, 
         que_out_20__4__13, que_out_20__4__12, que_out_20__4__11, 
         que_out_20__4__10, que_out_20__4__9, que_out_20__4__8, que_out_20__4__7, 
         que_out_20__4__6, que_out_20__4__5, que_out_20__4__4, que_out_20__4__3, 
         que_out_20__4__2, que_out_20__4__1, que_out_20__4__0, que_out_21__0__15, 
         que_out_21__0__14, que_out_21__0__13, que_out_21__0__12, 
         que_out_21__0__11, que_out_21__0__10, que_out_21__0__9, 
         que_out_21__0__8, que_out_21__0__7, que_out_21__0__6, que_out_21__0__5, 
         que_out_21__0__4, que_out_21__0__3, que_out_21__0__2, que_out_21__0__1, 
         que_out_21__0__0, que_out_21__1__15, que_out_21__1__14, 
         que_out_21__1__13, que_out_21__1__12, que_out_21__1__11, 
         que_out_21__1__10, que_out_21__1__9, que_out_21__1__8, que_out_21__1__7, 
         que_out_21__1__6, que_out_21__1__5, que_out_21__1__4, que_out_21__1__3, 
         que_out_21__1__2, que_out_21__1__1, que_out_21__1__0, que_out_21__2__15, 
         que_out_21__2__14, que_out_21__2__13, que_out_21__2__12, 
         que_out_21__2__11, que_out_21__2__10, que_out_21__2__9, 
         que_out_21__2__8, que_out_21__2__7, que_out_21__2__6, que_out_21__2__5, 
         que_out_21__2__4, que_out_21__2__3, que_out_21__2__2, que_out_21__2__1, 
         que_out_21__2__0, que_out_21__3__15, que_out_21__3__14, 
         que_out_21__3__13, que_out_21__3__12, que_out_21__3__11, 
         que_out_21__3__10, que_out_21__3__9, que_out_21__3__8, que_out_21__3__7, 
         que_out_21__3__6, que_out_21__3__5, que_out_21__3__4, que_out_21__3__3, 
         que_out_21__3__2, que_out_21__3__1, que_out_21__3__0, que_out_21__4__15, 
         que_out_21__4__14, que_out_21__4__13, que_out_21__4__12, 
         que_out_21__4__11, que_out_21__4__10, que_out_21__4__9, 
         que_out_21__4__8, que_out_21__4__7, que_out_21__4__6, que_out_21__4__5, 
         que_out_21__4__4, que_out_21__4__3, que_out_21__4__2, que_out_21__4__1, 
         que_out_21__4__0, que_out_22__0__15, que_out_22__0__14, 
         que_out_22__0__13, que_out_22__0__12, que_out_22__0__11, 
         que_out_22__0__10, que_out_22__0__9, que_out_22__0__8, que_out_22__0__7, 
         que_out_22__0__6, que_out_22__0__5, que_out_22__0__4, que_out_22__0__3, 
         que_out_22__0__2, que_out_22__0__1, que_out_22__0__0, que_out_22__1__15, 
         que_out_22__1__14, que_out_22__1__13, que_out_22__1__12, 
         que_out_22__1__11, que_out_22__1__10, que_out_22__1__9, 
         que_out_22__1__8, que_out_22__1__7, que_out_22__1__6, que_out_22__1__5, 
         que_out_22__1__4, que_out_22__1__3, que_out_22__1__2, que_out_22__1__1, 
         que_out_22__1__0, que_out_22__2__15, que_out_22__2__14, 
         que_out_22__2__13, que_out_22__2__12, que_out_22__2__11, 
         que_out_22__2__10, que_out_22__2__9, que_out_22__2__8, que_out_22__2__7, 
         que_out_22__2__6, que_out_22__2__5, que_out_22__2__4, que_out_22__2__3, 
         que_out_22__2__2, que_out_22__2__1, que_out_22__2__0, que_out_22__3__15, 
         que_out_22__3__14, que_out_22__3__13, que_out_22__3__12, 
         que_out_22__3__11, que_out_22__3__10, que_out_22__3__9, 
         que_out_22__3__8, que_out_22__3__7, que_out_22__3__6, que_out_22__3__5, 
         que_out_22__3__4, que_out_22__3__3, que_out_22__3__2, que_out_22__3__1, 
         que_out_22__3__0, que_out_22__4__15, que_out_22__4__14, 
         que_out_22__4__13, que_out_22__4__12, que_out_22__4__11, 
         que_out_22__4__10, que_out_22__4__9, que_out_22__4__8, que_out_22__4__7, 
         que_out_22__4__6, que_out_22__4__5, que_out_22__4__4, que_out_22__4__3, 
         que_out_22__4__2, que_out_22__4__1, que_out_22__4__0, que_out_23__0__15, 
         que_out_23__0__14, que_out_23__0__13, que_out_23__0__12, 
         que_out_23__0__11, que_out_23__0__10, que_out_23__0__9, 
         que_out_23__0__8, que_out_23__0__7, que_out_23__0__6, que_out_23__0__5, 
         que_out_23__0__4, que_out_23__0__3, que_out_23__0__2, que_out_23__0__1, 
         que_out_23__0__0, que_out_23__1__15, que_out_23__1__14, 
         que_out_23__1__13, que_out_23__1__12, que_out_23__1__11, 
         que_out_23__1__10, que_out_23__1__9, que_out_23__1__8, que_out_23__1__7, 
         que_out_23__1__6, que_out_23__1__5, que_out_23__1__4, que_out_23__1__3, 
         que_out_23__1__2, que_out_23__1__1, que_out_23__1__0, que_out_23__2__15, 
         que_out_23__2__14, que_out_23__2__13, que_out_23__2__12, 
         que_out_23__2__11, que_out_23__2__10, que_out_23__2__9, 
         que_out_23__2__8, que_out_23__2__7, que_out_23__2__6, que_out_23__2__5, 
         que_out_23__2__4, que_out_23__2__3, que_out_23__2__2, que_out_23__2__1, 
         que_out_23__2__0, que_out_23__3__15, que_out_23__3__14, 
         que_out_23__3__13, que_out_23__3__12, que_out_23__3__11, 
         que_out_23__3__10, que_out_23__3__9, que_out_23__3__8, que_out_23__3__7, 
         que_out_23__3__6, que_out_23__3__5, que_out_23__3__4, que_out_23__3__3, 
         que_out_23__3__2, que_out_23__3__1, que_out_23__3__0, que_out_23__4__15, 
         que_out_23__4__14, que_out_23__4__13, que_out_23__4__12, 
         que_out_23__4__11, que_out_23__4__10, que_out_23__4__9, 
         que_out_23__4__8, que_out_23__4__7, que_out_23__4__6, que_out_23__4__5, 
         que_out_23__4__4, que_out_23__4__3, que_out_23__4__2, que_out_23__4__1, 
         que_out_23__4__0, que_out_24__0__15, que_out_24__0__14, 
         que_out_24__0__13, que_out_24__0__12, que_out_24__0__11, 
         que_out_24__0__10, que_out_24__0__9, que_out_24__0__8, que_out_24__0__7, 
         que_out_24__0__6, que_out_24__0__5, que_out_24__0__4, que_out_24__0__3, 
         que_out_24__0__2, que_out_24__0__1, que_out_24__0__0, que_out_24__1__15, 
         que_out_24__1__14, que_out_24__1__13, que_out_24__1__12, 
         que_out_24__1__11, que_out_24__1__10, que_out_24__1__9, 
         que_out_24__1__8, que_out_24__1__7, que_out_24__1__6, que_out_24__1__5, 
         que_out_24__1__4, que_out_24__1__3, que_out_24__1__2, que_out_24__1__1, 
         que_out_24__1__0, que_out_24__2__15, que_out_24__2__14, 
         que_out_24__2__13, que_out_24__2__12, que_out_24__2__11, 
         que_out_24__2__10, que_out_24__2__9, que_out_24__2__8, que_out_24__2__7, 
         que_out_24__2__6, que_out_24__2__5, que_out_24__2__4, que_out_24__2__3, 
         que_out_24__2__2, que_out_24__2__1, que_out_24__2__0, que_out_24__3__15, 
         que_out_24__3__14, que_out_24__3__13, que_out_24__3__12, 
         que_out_24__3__11, que_out_24__3__10, que_out_24__3__9, 
         que_out_24__3__8, que_out_24__3__7, que_out_24__3__6, que_out_24__3__5, 
         que_out_24__3__4, que_out_24__3__3, que_out_24__3__2, que_out_24__3__1, 
         que_out_24__3__0, que_out_24__4__15, que_out_24__4__14, 
         que_out_24__4__13, que_out_24__4__12, que_out_24__4__11, 
         que_out_24__4__10, que_out_24__4__9, que_out_24__4__8, que_out_24__4__7, 
         que_out_24__4__6, que_out_24__4__5, que_out_24__4__4, que_out_24__4__3, 
         que_out_24__4__2, que_out_24__4__1, que_out_24__4__0, que_out_25__0__15, 
         que_out_25__0__14, que_out_25__0__13, que_out_25__0__12, 
         que_out_25__0__11, que_out_25__0__10, que_out_25__0__9, 
         que_out_25__0__8, que_out_25__0__7, que_out_25__0__6, que_out_25__0__5, 
         que_out_25__0__4, que_out_25__0__3, que_out_25__0__2, que_out_25__0__1, 
         que_out_25__0__0, que_out_25__1__15, que_out_25__1__14, 
         que_out_25__1__13, que_out_25__1__12, que_out_25__1__11, 
         que_out_25__1__10, que_out_25__1__9, que_out_25__1__8, que_out_25__1__7, 
         que_out_25__1__6, que_out_25__1__5, que_out_25__1__4, que_out_25__1__3, 
         que_out_25__1__2, que_out_25__1__1, que_out_25__1__0, que_out_25__2__15, 
         que_out_25__2__14, que_out_25__2__13, que_out_25__2__12, 
         que_out_25__2__11, que_out_25__2__10, que_out_25__2__9, 
         que_out_25__2__8, que_out_25__2__7, que_out_25__2__6, que_out_25__2__5, 
         que_out_25__2__4, que_out_25__2__3, que_out_25__2__2, que_out_25__2__1, 
         que_out_25__2__0, que_out_25__3__15, que_out_25__3__14, 
         que_out_25__3__13, que_out_25__3__12, que_out_25__3__11, 
         que_out_25__3__10, que_out_25__3__9, que_out_25__3__8, que_out_25__3__7, 
         que_out_25__3__6, que_out_25__3__5, que_out_25__3__4, que_out_25__3__3, 
         que_out_25__3__2, que_out_25__3__1, que_out_25__3__0, que_out_25__4__15, 
         que_out_25__4__14, que_out_25__4__13, que_out_25__4__12, 
         que_out_25__4__11, que_out_25__4__10, que_out_25__4__9, 
         que_out_25__4__8, que_out_25__4__7, que_out_25__4__6, que_out_25__4__5, 
         que_out_25__4__4, que_out_25__4__3, que_out_25__4__2, que_out_25__4__1, 
         que_out_25__4__0, que_out_26__0__15, que_out_26__0__14, 
         que_out_26__0__13, que_out_26__0__12, que_out_26__0__11, 
         que_out_26__0__10, que_out_26__0__9, que_out_26__0__8, que_out_26__0__7, 
         que_out_26__0__6, que_out_26__0__5, que_out_26__0__4, que_out_26__0__3, 
         que_out_26__0__2, que_out_26__0__1, que_out_26__0__0, que_out_26__1__15, 
         que_out_26__1__14, que_out_26__1__13, que_out_26__1__12, 
         que_out_26__1__11, que_out_26__1__10, que_out_26__1__9, 
         que_out_26__1__8, que_out_26__1__7, que_out_26__1__6, que_out_26__1__5, 
         que_out_26__1__4, que_out_26__1__3, que_out_26__1__2, que_out_26__1__1, 
         que_out_26__1__0, que_out_26__2__15, que_out_26__2__14, 
         que_out_26__2__13, que_out_26__2__12, que_out_26__2__11, 
         que_out_26__2__10, que_out_26__2__9, que_out_26__2__8, que_out_26__2__7, 
         que_out_26__2__6, que_out_26__2__5, que_out_26__2__4, que_out_26__2__3, 
         que_out_26__2__2, que_out_26__2__1, que_out_26__2__0, que_out_26__3__15, 
         que_out_26__3__14, que_out_26__3__13, que_out_26__3__12, 
         que_out_26__3__11, que_out_26__3__10, que_out_26__3__9, 
         que_out_26__3__8, que_out_26__3__7, que_out_26__3__6, que_out_26__3__5, 
         que_out_26__3__4, que_out_26__3__3, que_out_26__3__2, que_out_26__3__1, 
         que_out_26__3__0, que_out_26__4__15, que_out_26__4__14, 
         que_out_26__4__13, que_out_26__4__12, que_out_26__4__11, 
         que_out_26__4__10, que_out_26__4__9, que_out_26__4__8, que_out_26__4__7, 
         que_out_26__4__6, que_out_26__4__5, que_out_26__4__4, que_out_26__4__3, 
         que_out_26__4__2, que_out_26__4__1, que_out_26__4__0, que_out_27__0__15, 
         que_out_27__0__14, que_out_27__0__13, que_out_27__0__12, 
         que_out_27__0__11, que_out_27__0__10, que_out_27__0__9, 
         que_out_27__0__8, que_out_27__0__7, que_out_27__0__6, que_out_27__0__5, 
         que_out_27__0__4, que_out_27__0__3, que_out_27__0__2, que_out_27__0__1, 
         que_out_27__0__0, que_out_27__1__15, que_out_27__1__14, 
         que_out_27__1__13, que_out_27__1__12, que_out_27__1__11, 
         que_out_27__1__10, que_out_27__1__9, que_out_27__1__8, que_out_27__1__7, 
         que_out_27__1__6, que_out_27__1__5, que_out_27__1__4, que_out_27__1__3, 
         que_out_27__1__2, que_out_27__1__1, que_out_27__1__0, que_out_27__2__15, 
         que_out_27__2__14, que_out_27__2__13, que_out_27__2__12, 
         que_out_27__2__11, que_out_27__2__10, que_out_27__2__9, 
         que_out_27__2__8, que_out_27__2__7, que_out_27__2__6, que_out_27__2__5, 
         que_out_27__2__4, que_out_27__2__3, que_out_27__2__2, que_out_27__2__1, 
         que_out_27__2__0, que_out_27__3__15, que_out_27__3__14, 
         que_out_27__3__13, que_out_27__3__12, que_out_27__3__11, 
         que_out_27__3__10, que_out_27__3__9, que_out_27__3__8, que_out_27__3__7, 
         que_out_27__3__6, que_out_27__3__5, que_out_27__3__4, que_out_27__3__3, 
         que_out_27__3__2, que_out_27__3__1, que_out_27__3__0, que_out_27__4__15, 
         que_out_27__4__14, que_out_27__4__13, que_out_27__4__12, 
         que_out_27__4__11, que_out_27__4__10, que_out_27__4__9, 
         que_out_27__4__8, que_out_27__4__7, que_out_27__4__6, que_out_27__4__5, 
         que_out_27__4__4, que_out_27__4__3, que_out_27__4__2, que_out_27__4__1, 
         que_out_27__4__0, sel_que_27, sel_que_26, sel_que_25, sel_que_24, 
         sel_que_23, sel_que_22, sel_que_21, sel_que_20, sel_que_19, sel_que_18, 
         sel_que_17, sel_que_16, sel_que_15, sel_que_14, sel_que_13, sel_que_12, 
         sel_que_11, sel_que_10, sel_que_9, sel_que_8, sel_que_7, sel_que_6, 
         sel_que_5, sel_que_4, sel_que_3, sel_que_2, sel_que_1, sel_que_0, nx12, 
         nx14, nx28, nx30, nx42, nx48, nx62, nx64, nx68, nx74, nx82, nx88, nx90, 
         nx94, nx100, nx104, nx114, nx118, nx122, nx130, nx136, nx144, nx150, 
         nx158, nx166, nx172, nx180, nx188, nx192, nx200, nx206, nx214, nx222, 
         nx226, nx230, nx238, nx268, nx294, nx322, nx348, nx378, nx404, nx432, 
         nx458, nx488, nx514, nx542, nx568, nx598, nx624, nx652, nx678, nx708, 
         nx734, nx762, nx788, nx818, nx844, nx872, nx898, nx928, nx954, nx982, 
         nx1008, nx1038, nx1064, nx1092, nx1118, nx1148, nx1174, nx1202, nx1228, 
         nx1258, nx1284, nx1312, nx1338, nx1368, nx1394, nx1422, nx1448, nx1478, 
         nx1504, nx1532, nx1558, nx1588, nx1614, nx1642, nx1668, nx1698, nx1724, 
         nx1752, nx1778, nx1808, nx1834, nx1862, nx1888, nx1918, nx1944, nx1972, 
         nx1998, nx2028, nx2054, nx2082, nx2108, nx2138, nx2164, nx2192, nx2218, 
         nx2248, nx2274, nx2302, nx2328, nx2358, nx2384, nx2412, nx2438, nx2468, 
         nx2494, nx2522, nx2548, nx2578, nx2604, nx2632, nx2658, nx2688, nx2714, 
         nx2742, nx2768, nx2798, nx2824, nx2852, nx2878, nx2908, nx2934, nx2962, 
         nx2988, nx3018, nx3044, nx3072, nx3098, nx3128, nx3154, nx3182, nx3208, 
         nx3238, nx3264, nx3292, nx3318, nx3348, nx3374, nx3402, nx3428, nx3458, 
         nx3484, nx3512, nx3538, nx3568, nx3594, nx3622, nx3648, nx3678, nx3704, 
         nx3732, nx3758, nx3788, nx3814, nx3842, nx3868, nx3898, nx3924, nx3952, 
         nx3978, nx4008, nx4034, nx4062, nx4088, nx4118, nx4144, nx4172, nx4198, 
         nx4228, nx4254, nx4282, nx4308, nx4338, nx4364, nx4392, nx4418, nx4448, 
         nx4474, nx4502, nx4528, nx4558, nx4584, nx4612, nx4638, nx4668, nx4694, 
         nx4722, nx4748, nx4778, nx4804, nx4832, nx4858, nx4888, nx4914, nx4942, 
         nx4968, nx4998, nx5024, nx5052, nx5078, nx5108, nx5134, nx5162, nx5188, 
         nx5218, nx5244, nx5272, nx5298, nx5328, nx5354, nx5382, nx5408, nx5438, 
         nx5464, nx5492, nx5518, nx5548, nx5574, nx5602, nx5628, nx5658, nx5684, 
         nx5712, nx5738, nx5768, nx5794, nx5822, nx5848, nx5878, nx5904, nx5932, 
         nx5958, nx5988, nx6014, nx6042, nx6068, nx6098, nx6124, nx6152, nx6178, 
         nx6208, nx6234, nx6262, nx6288, nx6318, nx6344, nx6372, nx6398, nx6428, 
         nx6454, nx6482, nx6508, nx6538, nx6564, nx6592, nx6618, nx6648, nx6674, 
         nx6702, nx6728, nx6758, nx6784, nx6812, nx6838, nx6868, nx6894, nx6922, 
         nx6948, nx6978, nx7004, nx7032, nx7058, nx7088, nx7114, nx7142, nx7168, 
         nx7198, nx7224, nx7252, nx7278, nx7308, nx7334, nx7362, nx7388, nx7418, 
         nx7444, nx7472, nx7498, nx7528, nx7554, nx7582, nx7608, nx7638, nx7664, 
         nx7692, nx7718, nx7748, nx7774, nx7802, nx7828, nx7858, nx7884, nx7912, 
         nx7938, nx7968, nx7994, nx8022, nx8048, nx8078, nx8104, nx8132, nx8158, 
         nx8188, nx8214, nx8242, nx8268, nx8298, nx8324, nx8352, nx8378, nx8408, 
         nx8434, nx8462, nx8488, nx8518, nx8544, nx8572, nx8598, nx8628, nx8654, 
         nx8682, nx8708, nx8738, nx8764, nx8792, nx8818, nx8848, nx8874, nx8902, 
         nx8928, nx8938, nx9038, nx6829, nx6833, nx6835, nx6839, nx6843, nx6847, 
         nx6875, nx6885, nx6889, nx6893, nx6897, nx6901, nx6905, nx6915, nx6927, 
         nx6931, nx6933, nx6937, nx6939, nx6943, nx6945, nx6949, nx6951, nx6955, 
         nx6957, nx6961, nx6965, nx6967, nx6971, nx6977, nx6985, nx6991, nx6999, 
         nx7007, nx7017, nx7029, nx7037, nx7043, nx7053, nx7055, nx7057, nx7061, 
         nx7063, nx7065, nx7069, nx7071, nx7073, nx7077, nx7079, nx7081, nx7087, 
         nx7089, nx7091, nx7095, nx7097, nx7099, nx7103, nx7105, nx7107, nx7111, 
         nx7113, nx7115, nx7121, nx7123, nx7125, nx7129, nx7131, nx7133, nx7137, 
         nx7139, nx7141, nx7145, nx7147, nx7149, nx7155, nx7157, nx7159, nx7163, 
         nx7165, nx7167, nx7171, nx7173, nx7175, nx7179, nx7181, nx7183, nx7189, 
         nx7191, nx7193, nx7197, nx7199, nx7201, nx7205, nx7207, nx7209, nx7213, 
         nx7215, nx7217, nx7223, nx7225, nx7227, nx7231, nx7233, nx7235, nx7239, 
         nx7241, nx7243, nx7247, nx7249, nx7251, nx7257, nx7259, nx7261, nx7265, 
         nx7267, nx7269, nx7273, nx7275, nx7277, nx7281, nx7283, nx7285, nx7291, 
         nx7293, nx7295, nx7299, nx7301, nx7303, nx7307, nx7309, nx7311, nx7315, 
         nx7317, nx7319, nx7325, nx7327, nx7329, nx7333, nx7335, nx7337, nx7341, 
         nx7343, nx7345, nx7349, nx7351, nx7353, nx7359, nx7361, nx7363, nx7367, 
         nx7369, nx7371, nx7375, nx7377, nx7379, nx7383, nx7385, nx7387, nx7393, 
         nx7395, nx7397, nx7401, nx7403, nx7405, nx7409, nx7411, nx7413, nx7417, 
         nx7419, nx7421, nx7427, nx7429, nx7431, nx7435, nx7437, nx7439, nx7443, 
         nx7445, nx7447, nx7451, nx7453, nx7455, nx7461, nx7463, nx7465, nx7469, 
         nx7471, nx7473, nx7477, nx7479, nx7481, nx7485, nx7487, nx7489, nx7495, 
         nx7497, nx7499, nx7503, nx7505, nx7507, nx7511, nx7513, nx7515, nx7519, 
         nx7521, nx7523, nx7529, nx7531, nx7533, nx7537, nx7539, nx7541, nx7545, 
         nx7547, nx7549, nx7553, nx7555, nx7557, nx7563, nx7565, nx7567, nx7571, 
         nx7573, nx7575, nx7579, nx7581, nx7583, nx7587, nx7589, nx7591, nx7597, 
         nx7599, nx7601, nx7605, nx7607, nx7609, nx7613, nx7615, nx7617, nx7621, 
         nx7623, nx7625, nx7631, nx7633, nx7635, nx7639, nx7641, nx7643, nx7647, 
         nx7649, nx7651, nx7655, nx7657, nx7659, nx7665, nx7667, nx7669, nx7673, 
         nx7675, nx7677, nx7681, nx7683, nx7685, nx7689, nx7691, nx7693, nx7699, 
         nx7701, nx7703, nx7707, nx7709, nx7711, nx7715, nx7717, nx7719, nx7723, 
         nx7725, nx7727, nx7733, nx7735, nx7737, nx7741, nx7743, nx7745, nx7749, 
         nx7751, nx7753, nx7757, nx7759, nx7761, nx7767, nx7769, nx7771, nx7775, 
         nx7777, nx7779, nx7783, nx7785, nx7787, nx7791, nx7793, nx7795, nx7801, 
         nx7803, nx7805, nx7809, nx7811, nx7813, nx7817, nx7819, nx7821, nx7825, 
         nx7827, nx7829, nx7835, nx7837, nx7839, nx7843, nx7845, nx7847, nx7851, 
         nx7853, nx7855, nx7859, nx7861, nx7863, nx7869, nx7871, nx7873, nx7877, 
         nx7879, nx7881, nx7885, nx7887, nx7889, nx7893, nx7895, nx7897, nx7903, 
         nx7905, nx7907, nx7911, nx7913, nx7915, nx7919, nx7921, nx7923, nx7927, 
         nx7929, nx7931, nx7937, nx7939, nx7941, nx7945, nx7947, nx7949, nx7953, 
         nx7955, nx7957, nx7961, nx7963, nx7965, nx7971, nx7973, nx7975, nx7979, 
         nx7981, nx7983, nx7987, nx7989, nx7991, nx7995, nx7997, nx7999, nx8005, 
         nx8007, nx8009, nx8013, nx8015, nx8017, nx8021, nx8023, nx8025, nx8029, 
         nx8031, nx8033, nx8039, nx8041, nx8043, nx8047, nx8049, nx8051, nx8055, 
         nx8057, nx8059, nx8063, nx8065, nx8067, nx8073, nx8075, nx8077, nx8081, 
         nx8083, nx8085, nx8089, nx8091, nx8093, nx8097, nx8099, nx8101, nx8107, 
         nx8109, nx8111, nx8115, nx8117, nx8119, nx8123, nx8125, nx8127, nx8131, 
         nx8133, nx8135, nx8141, nx8143, nx8145, nx8149, nx8151, nx8153, nx8157, 
         nx8159, nx8161, nx8165, nx8167, nx8169, nx8175, nx8177, nx8179, nx8183, 
         nx8185, nx8187, nx8191, nx8193, nx8195, nx8199, nx8201, nx8203, nx8209, 
         nx8211, nx8213, nx8217, nx8219, nx8221, nx8225, nx8227, nx8229, nx8233, 
         nx8235, nx8237, nx8243, nx8245, nx8247, nx8251, nx8253, nx8255, nx8259, 
         nx8261, nx8263, nx8267, nx8269, nx8271, nx8277, nx8279, nx8281, nx8285, 
         nx8287, nx8289, nx8293, nx8295, nx8297, nx8301, nx8303, nx8305, nx8311, 
         nx8313, nx8315, nx8319, nx8321, nx8323, nx8327, nx8329, nx8331, nx8335, 
         nx8337, nx8339, nx8345, nx8347, nx8349, nx8353, nx8355, nx8357, nx8361, 
         nx8363, nx8365, nx8369, nx8371, nx8373, nx8379, nx8381, nx8383, nx8387, 
         nx8389, nx8391, nx8395, nx8397, nx8399, nx8403, nx8405, nx8407, nx8413, 
         nx8415, nx8417, nx8421, nx8423, nx8425, nx8429, nx8431, nx8433, nx8437, 
         nx8439, nx8441, nx8447, nx8449, nx8451, nx8455, nx8457, nx8459, nx8463, 
         nx8465, nx8467, nx8471, nx8473, nx8475, nx8481, nx8483, nx8485, nx8489, 
         nx8491, nx8493, nx8497, nx8499, nx8501, nx8505, nx8507, nx8509, nx8515, 
         nx8517, nx8519, nx8523, nx8525, nx8527, nx8531, nx8533, nx8535, nx8539, 
         nx8541, nx8543, nx8549, nx8551, nx8553, nx8557, nx8559, nx8561, nx8565, 
         nx8567, nx8569, nx8573, nx8575, nx8577, nx8583, nx8585, nx8587, nx8591, 
         nx8593, nx8595, nx8599, nx8601, nx8603, nx8607, nx8609, nx8611, nx8617, 
         nx8619, nx8621, nx8625, nx8627, nx8629, nx8633, nx8635, nx8637, nx8641, 
         nx8643, nx8645, nx8651, nx8653, nx8655, nx8659, nx8661, nx8663, nx8667, 
         nx8669, nx8671, nx8675, nx8677, nx8679, nx8685, nx8687, nx8689, nx8693, 
         nx8695, nx8697, nx8701, nx8703, nx8705, nx8709, nx8711, nx8713, nx8719, 
         nx8721, nx8723, nx8727, nx8729, nx8731, nx8735, nx8737, nx8739, nx8743, 
         nx8745, nx8747, nx8753, nx8755, nx8757, nx8761, nx8763, nx8765, nx8769, 
         nx8771, nx8773, nx8777, nx8779, nx8781, nx8787, nx8789, nx8791, nx8795, 
         nx8797, nx8799, nx8803, nx8805, nx8807, nx8811, nx8813, nx8815, nx8821, 
         nx8823, nx8825, nx8829, nx8831, nx8833, nx8837, nx8839, nx8841, nx8845, 
         nx8847, nx8849, nx8855, nx8857, nx8859, nx8863, nx8865, nx8867, nx8871, 
         nx8873, nx8875, nx8879, nx8881, nx8883, nx8889, nx8891, nx8893, nx8897, 
         nx8899, nx8901, nx8905, nx8907, nx8909, nx8913, nx8915, nx8917, nx8923, 
         nx8925, nx8927, nx8931, nx8933, nx8935, nx8939, nx8941, nx8943, nx8947, 
         nx8949, nx8951, nx8955, nx8957, nx8959, nx8963, nx8965, nx8967, nx8970, 
         nx8973, nx8975, nx8978, nx8981, nx8983, nx8989, nx8991, nx8993, nx8997, 
         nx8999, nx9001, nx9005, nx9007, nx9009, nx9013, nx9015, nx9017, nx9023, 
         nx9025, nx9027, nx9031, nx9033, nx9035, nx9039, nx9041, nx9043, nx9047, 
         nx9049, nx9051, nx9057, nx9059, nx9061, nx9065, nx9067, nx9069, nx9073, 
         nx9075, nx9077, nx9081, nx9083, nx9085, nx9090, nx9093, nx9095, nx9098, 
         nx9101, nx9103, nx9106, nx9108, nx9110, nx9113, nx9115, nx9117, nx9121, 
         nx9123, nx9125, nx9128, nx9130, nx9132, nx9135, nx9137, nx9139, nx9142, 
         nx9144, nx9146, nx9150, nx9152, nx9154, nx9157, nx9159, nx9161, nx9164, 
         nx9166, nx9168, nx9171, nx9173, nx9175, nx9179, nx9181, nx9183, nx9186, 
         nx9188, nx9190, nx9193, nx9195, nx9197, nx9200, nx9202, nx9204, nx9208, 
         nx9210, nx9212, nx9215, nx9217, nx9219, nx9222, nx9224, nx9226, nx9229, 
         nx9231, nx9233, nx9237, nx9239, nx9241, nx9244, nx9246, nx9248, nx9251, 
         nx9253, nx9255, nx9258, nx9260, nx9262, nx9266, nx9268, nx9270, nx9273, 
         nx9275, nx9277, nx9280, nx9282, nx9284, nx9287, nx9289, nx9291, nx9295, 
         nx9297, nx9299, nx9302, nx9304, nx9306, nx9309, nx9311, nx9313, nx9316, 
         nx9318, nx9320, nx9324, nx9326, nx9328, nx9331, nx9333, nx9335, nx9338, 
         nx9340, nx9342, nx9345, nx9347, nx9349, nx9353, nx9355, nx9357, nx9360, 
         nx9362, nx9364, nx9367, nx9369, nx9371, nx9374, nx9376, nx9378, nx9382, 
         nx9384, nx9386, nx9389, nx9391, nx9393, nx9396, nx9398, nx9400, nx9403, 
         nx9405, nx9407, nx9411, nx9413, nx9415, nx9418, nx9420, nx9422, nx9425, 
         nx9427, nx9429, nx9432, nx9434, nx9436, nx9440, nx9442, nx9444, nx9447, 
         nx9449, nx9451, nx9454, nx9456, nx9458, nx9461, nx9463, nx9465, nx9469, 
         nx9471, nx9473, nx9476, nx9478, nx9480, nx9483, nx9485, nx9487, nx9490, 
         nx9492, nx9494, nx9498, nx9500, nx9502, nx9505, nx9507, nx9509, nx9512, 
         nx9514, nx9516, nx9519, nx9521, nx9523, nx9527, nx9529, nx9531, nx9534, 
         nx9536, nx9538, nx9541, nx9543, nx9545, nx9548, nx9550, nx9552, nx9556, 
         nx9558, nx9560, nx9563, nx9565, nx9567, nx9570, nx9572, nx9574, nx9577, 
         nx9579, nx9581, nx9585, nx9587, nx9589, nx9592, nx9594, nx9596, nx9599, 
         nx9601, nx9603, nx9606, nx9608, nx9610, nx9614, nx9616, nx9618, nx9621, 
         nx9623, nx9625, nx9628, nx9630, nx9632, nx9635, nx9637, nx9639, nx9648, 
         nx9650, nx9652, nx9654, nx9656, nx9658, nx9660, nx9662, nx9664, nx9666, 
         nx9668, nx9670, nx9674, nx9676, nx9678, nx9680, nx9682, nx9684, nx9686, 
         nx9688, nx9690, nx9692, nx9694, nx9696, nx9700, nx9702, nx9704, nx9706, 
         nx9708, nx9710, nx9712, nx9714, nx9716, nx9718, nx9720, nx9722, nx9726, 
         nx9728, nx9730, nx9732, nx9734, nx9736, nx9738, nx9740, nx9742, nx9744, 
         nx9746, nx9748, nx9752, nx9754, nx9756, nx9758, nx9760, nx9762, nx9764, 
         nx9766, nx9768, nx9770, nx9772, nx9774, nx9778, nx9780, nx9782, nx9784, 
         nx9786, nx9788, nx9790, nx9792, nx9794, nx9796, nx9798, nx9800, nx9804, 
         nx9806, nx9808, nx9810, nx9812, nx9814, nx9816, nx9818, nx9820, nx9822, 
         nx9824, nx9826, nx9830, nx9832, nx9834, nx9836, nx9838, nx9840, nx9842, 
         nx9844, nx9846, nx9848, nx9850, nx9852, nx9856, nx9858, nx9860, nx9862, 
         nx9864, nx9866, nx9868, nx9870, nx9872, nx9874, nx9876, nx9878, nx9882, 
         nx9884, nx9886, nx9888, nx9890, nx9892, nx9894, nx9896, nx9898, nx9900, 
         nx9902, nx9904, nx9908, nx9910, nx9912, nx9914, nx9916, nx9918, nx9920, 
         nx9922, nx9924, nx9926, nx9928, nx9930, nx9934, nx9936, nx9938, nx9940, 
         nx9942, nx9944, nx9946, nx9948, nx9950, nx9952, nx9954, nx9956, nx9960, 
         nx9962, nx9964, nx9966, nx9968, nx9970, nx9972, nx9974, nx9976, nx9978, 
         nx9980, nx9982, nx9986, nx9988, nx9990, nx9992, nx9994, nx9996, nx9998, 
         nx10000, nx10002, nx10004, nx10006, nx10008, nx10012, nx10014, nx10016, 
         nx10018, nx10020, nx10022, nx10024, nx10026, nx10028, nx10030, nx10032, 
         nx10034, nx10038, nx10040, nx10042, nx10044, nx10046, nx10048, nx10050, 
         nx10052, nx10054, nx10056, nx10058, nx10060, nx10064, nx10066, nx10068, 
         nx10070, nx10072, nx10074, nx10076, nx10078, nx10080, nx10082, nx10084, 
         nx10086, nx10090, nx10092, nx10094, nx10096, nx10098, nx10100, nx10102, 
         nx10104, nx10106, nx10108, nx10110, nx10112, nx10116, nx10118, nx10120, 
         nx10122, nx10124, nx10126, nx10128, nx10130, nx10132, nx10134, nx10136, 
         nx10138, nx10142, nx10144, nx10146, nx10148, nx10150, nx10152, nx10154, 
         nx10156, nx10158, nx10160, nx10162, nx10164, nx10168, nx10170, nx10172, 
         nx10174, nx10176, nx10178, nx10180, nx10182, nx10184, nx10186, nx10188, 
         nx10190, nx10194, nx10196, nx10198, nx10200, nx10202, nx10204, nx10206, 
         nx10208, nx10210, nx10212, nx10214, nx10216, nx10220, nx10222, nx10224, 
         nx10226, nx10228, nx10230, nx10232, nx10234, nx10236, nx10238, nx10240, 
         nx10242, nx10246, nx10248, nx10250, nx10252, nx10254, nx10256, nx10258, 
         nx10260, nx10262, nx10264, nx10266, nx10268, nx10272, nx10274, nx10276, 
         nx10278, nx10280, nx10282, nx10284, nx10286, nx10288, nx10290, nx10292, 
         nx10294, nx10298, nx10300, nx10302, nx10304, nx10306, nx10308, nx10310, 
         nx10312, nx10314, nx10316, nx10318, nx10320, nx10324, nx10326, nx10328, 
         nx10330, nx10332, nx10334, nx10336, nx10338, nx10340, nx10342, nx10344, 
         nx10346, nx10350, nx10352, nx10354, nx10356, nx10358, nx10360, nx10362, 
         nx10364, nx10366, nx10368, nx10370, nx10372, nx10374, nx10376, nx10378, 
         nx10380, nx10382, nx10384, nx10386, nx10388, nx10390, nx10392, nx10394, 
         nx10396, nx10398, nx10400, nx10402, nx10404, nx10406, nx10408, nx10410, 
         nx10412, nx10414, nx10416, nx10418, nx10420, nx10422, nx10424, nx10426, 
         nx10428, nx10430, nx10432, nx10434, nx10436, nx10438, nx10440, nx10442, 
         nx10444, nx10446, nx10448, nx10450, nx10452, nx10454, nx10456, nx10458, 
         nx10460, nx10462, nx10464, nx10466, nx10468, nx10470, nx10472, nx10474, 
         nx10476, nx10478, nx10480, nx10482, nx10484, nx10486, nx10488, nx10494, 
         nx10496, nx10498, nx10500, nx10502, nx10504, nx10506, nx10508, nx10510, 
         nx10512, nx10514, nx10516, nx10518, nx10520, nx10522, nx10524, nx10526, 
         nx10528, nx10530, nx10532, nx10534, nx10536, nx10538, nx10540, nx10542, 
         nx10544, nx10546, nx10548, nx10550, nx10552, nx10554, nx10556, nx10558, 
         nx10560, nx10562, nx10564, nx10566, nx10568, nx10570, nx10572, nx10574, 
         nx10576, nx10578, nx10580, nx10582, nx10584, nx10586, nx10588, nx10590, 
         nx10592, nx10594, nx10596, nx10598, nx10600, nx10602, nx10604, nx10606, 
         nx10608, nx10610, nx10612, nx10614, nx10616, nx10618, nx10620, nx10622, 
         nx10624, nx10626, nx10628, nx10630, nx10632, nx10634, nx10636, nx10638, 
         nx10640, nx10642, nx10644, nx10646, nx10648, nx10650, nx10652, nx10654, 
         nx10656, nx10658, nx10660, nx10662, nx10664, nx10666, nx10668, nx10690, 
         nx10692, nx10694, nx10696, nx10698, nx10700, nx10702, nx10704, nx10706, 
         nx10708, nx10710, nx10712, nx10714, nx10716, nx10718, nx10720, nx10722, 
         nx10724, nx10726, nx10728, nx10730, nx10732, nx10734, nx10736, nx10742, 
         nx10744, nx10746, nx10748;



    Queue_5 gen_queues_0_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_0__0__15), .q_0__14 (
            que_out_0__0__14), .q_0__13 (que_out_0__0__13), .q_0__12 (
            que_out_0__0__12), .q_0__11 (que_out_0__0__11), .q_0__10 (
            que_out_0__0__10), .q_0__9 (que_out_0__0__9), .q_0__8 (
            que_out_0__0__8), .q_0__7 (que_out_0__0__7), .q_0__6 (
            que_out_0__0__6), .q_0__5 (que_out_0__0__5), .q_0__4 (
            que_out_0__0__4), .q_0__3 (que_out_0__0__3), .q_0__2 (
            que_out_0__0__2), .q_0__1 (que_out_0__0__1), .q_0__0 (
            que_out_0__0__0), .q_1__15 (que_out_0__1__15), .q_1__14 (
            que_out_0__1__14), .q_1__13 (que_out_0__1__13), .q_1__12 (
            que_out_0__1__12), .q_1__11 (que_out_0__1__11), .q_1__10 (
            que_out_0__1__10), .q_1__9 (que_out_0__1__9), .q_1__8 (
            que_out_0__1__8), .q_1__7 (que_out_0__1__7), .q_1__6 (
            que_out_0__1__6), .q_1__5 (que_out_0__1__5), .q_1__4 (
            que_out_0__1__4), .q_1__3 (que_out_0__1__3), .q_1__2 (
            que_out_0__1__2), .q_1__1 (que_out_0__1__1), .q_1__0 (
            que_out_0__1__0), .q_2__15 (que_out_0__2__15), .q_2__14 (
            que_out_0__2__14), .q_2__13 (que_out_0__2__13), .q_2__12 (
            que_out_0__2__12), .q_2__11 (que_out_0__2__11), .q_2__10 (
            que_out_0__2__10), .q_2__9 (que_out_0__2__9), .q_2__8 (
            que_out_0__2__8), .q_2__7 (que_out_0__2__7), .q_2__6 (
            que_out_0__2__6), .q_2__5 (que_out_0__2__5), .q_2__4 (
            que_out_0__2__4), .q_2__3 (que_out_0__2__3), .q_2__2 (
            que_out_0__2__2), .q_2__1 (que_out_0__2__1), .q_2__0 (
            que_out_0__2__0), .q_3__15 (que_out_0__3__15), .q_3__14 (
            que_out_0__3__14), .q_3__13 (que_out_0__3__13), .q_3__12 (
            que_out_0__3__12), .q_3__11 (que_out_0__3__11), .q_3__10 (
            que_out_0__3__10), .q_3__9 (que_out_0__3__9), .q_3__8 (
            que_out_0__3__8), .q_3__7 (que_out_0__3__7), .q_3__6 (
            que_out_0__3__6), .q_3__5 (que_out_0__3__5), .q_3__4 (
            que_out_0__3__4), .q_3__3 (que_out_0__3__3), .q_3__2 (
            que_out_0__3__2), .q_3__1 (que_out_0__3__1), .q_3__0 (
            que_out_0__3__0), .q_4__15 (que_out_0__4__15), .q_4__14 (
            que_out_0__4__14), .q_4__13 (que_out_0__4__13), .q_4__12 (
            que_out_0__4__12), .q_4__11 (que_out_0__4__11), .q_4__10 (
            que_out_0__4__10), .q_4__9 (que_out_0__4__9), .q_4__8 (
            que_out_0__4__8), .q_4__7 (que_out_0__4__7), .q_4__6 (
            que_out_0__4__6), .q_4__5 (que_out_0__4__5), .q_4__4 (
            que_out_0__4__4), .q_4__3 (que_out_0__4__3), .q_4__2 (
            que_out_0__4__2), .q_4__1 (que_out_0__4__1), .q_4__0 (
            que_out_0__4__0), .clk (nx10714), .load (sel_que_0), .reset (nx10690
            )) ;
    Queue_5 gen_queues_1_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_1__0__15), .q_0__14 (
            que_out_1__0__14), .q_0__13 (que_out_1__0__13), .q_0__12 (
            que_out_1__0__12), .q_0__11 (que_out_1__0__11), .q_0__10 (
            que_out_1__0__10), .q_0__9 (que_out_1__0__9), .q_0__8 (
            que_out_1__0__8), .q_0__7 (que_out_1__0__7), .q_0__6 (
            que_out_1__0__6), .q_0__5 (que_out_1__0__5), .q_0__4 (
            que_out_1__0__4), .q_0__3 (que_out_1__0__3), .q_0__2 (
            que_out_1__0__2), .q_0__1 (que_out_1__0__1), .q_0__0 (
            que_out_1__0__0), .q_1__15 (que_out_1__1__15), .q_1__14 (
            que_out_1__1__14), .q_1__13 (que_out_1__1__13), .q_1__12 (
            que_out_1__1__12), .q_1__11 (que_out_1__1__11), .q_1__10 (
            que_out_1__1__10), .q_1__9 (que_out_1__1__9), .q_1__8 (
            que_out_1__1__8), .q_1__7 (que_out_1__1__7), .q_1__6 (
            que_out_1__1__6), .q_1__5 (que_out_1__1__5), .q_1__4 (
            que_out_1__1__4), .q_1__3 (que_out_1__1__3), .q_1__2 (
            que_out_1__1__2), .q_1__1 (que_out_1__1__1), .q_1__0 (
            que_out_1__1__0), .q_2__15 (que_out_1__2__15), .q_2__14 (
            que_out_1__2__14), .q_2__13 (que_out_1__2__13), .q_2__12 (
            que_out_1__2__12), .q_2__11 (que_out_1__2__11), .q_2__10 (
            que_out_1__2__10), .q_2__9 (que_out_1__2__9), .q_2__8 (
            que_out_1__2__8), .q_2__7 (que_out_1__2__7), .q_2__6 (
            que_out_1__2__6), .q_2__5 (que_out_1__2__5), .q_2__4 (
            que_out_1__2__4), .q_2__3 (que_out_1__2__3), .q_2__2 (
            que_out_1__2__2), .q_2__1 (que_out_1__2__1), .q_2__0 (
            que_out_1__2__0), .q_3__15 (que_out_1__3__15), .q_3__14 (
            que_out_1__3__14), .q_3__13 (que_out_1__3__13), .q_3__12 (
            que_out_1__3__12), .q_3__11 (que_out_1__3__11), .q_3__10 (
            que_out_1__3__10), .q_3__9 (que_out_1__3__9), .q_3__8 (
            que_out_1__3__8), .q_3__7 (que_out_1__3__7), .q_3__6 (
            que_out_1__3__6), .q_3__5 (que_out_1__3__5), .q_3__4 (
            que_out_1__3__4), .q_3__3 (que_out_1__3__3), .q_3__2 (
            que_out_1__3__2), .q_3__1 (que_out_1__3__1), .q_3__0 (
            que_out_1__3__0), .q_4__15 (que_out_1__4__15), .q_4__14 (
            que_out_1__4__14), .q_4__13 (que_out_1__4__13), .q_4__12 (
            que_out_1__4__12), .q_4__11 (que_out_1__4__11), .q_4__10 (
            que_out_1__4__10), .q_4__9 (que_out_1__4__9), .q_4__8 (
            que_out_1__4__8), .q_4__7 (que_out_1__4__7), .q_4__6 (
            que_out_1__4__6), .q_4__5 (que_out_1__4__5), .q_4__4 (
            que_out_1__4__4), .q_4__3 (que_out_1__4__3), .q_4__2 (
            que_out_1__4__2), .q_4__1 (que_out_1__4__1), .q_4__0 (
            que_out_1__4__0), .clk (nx10714), .load (sel_que_1), .reset (nx10690
            )) ;
    Queue_5 gen_queues_2_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_2__0__15), .q_0__14 (
            que_out_2__0__14), .q_0__13 (que_out_2__0__13), .q_0__12 (
            que_out_2__0__12), .q_0__11 (que_out_2__0__11), .q_0__10 (
            que_out_2__0__10), .q_0__9 (que_out_2__0__9), .q_0__8 (
            que_out_2__0__8), .q_0__7 (que_out_2__0__7), .q_0__6 (
            que_out_2__0__6), .q_0__5 (que_out_2__0__5), .q_0__4 (
            que_out_2__0__4), .q_0__3 (que_out_2__0__3), .q_0__2 (
            que_out_2__0__2), .q_0__1 (que_out_2__0__1), .q_0__0 (
            que_out_2__0__0), .q_1__15 (que_out_2__1__15), .q_1__14 (
            que_out_2__1__14), .q_1__13 (que_out_2__1__13), .q_1__12 (
            que_out_2__1__12), .q_1__11 (que_out_2__1__11), .q_1__10 (
            que_out_2__1__10), .q_1__9 (que_out_2__1__9), .q_1__8 (
            que_out_2__1__8), .q_1__7 (que_out_2__1__7), .q_1__6 (
            que_out_2__1__6), .q_1__5 (que_out_2__1__5), .q_1__4 (
            que_out_2__1__4), .q_1__3 (que_out_2__1__3), .q_1__2 (
            que_out_2__1__2), .q_1__1 (que_out_2__1__1), .q_1__0 (
            que_out_2__1__0), .q_2__15 (que_out_2__2__15), .q_2__14 (
            que_out_2__2__14), .q_2__13 (que_out_2__2__13), .q_2__12 (
            que_out_2__2__12), .q_2__11 (que_out_2__2__11), .q_2__10 (
            que_out_2__2__10), .q_2__9 (que_out_2__2__9), .q_2__8 (
            que_out_2__2__8), .q_2__7 (que_out_2__2__7), .q_2__6 (
            que_out_2__2__6), .q_2__5 (que_out_2__2__5), .q_2__4 (
            que_out_2__2__4), .q_2__3 (que_out_2__2__3), .q_2__2 (
            que_out_2__2__2), .q_2__1 (que_out_2__2__1), .q_2__0 (
            que_out_2__2__0), .q_3__15 (que_out_2__3__15), .q_3__14 (
            que_out_2__3__14), .q_3__13 (que_out_2__3__13), .q_3__12 (
            que_out_2__3__12), .q_3__11 (que_out_2__3__11), .q_3__10 (
            que_out_2__3__10), .q_3__9 (que_out_2__3__9), .q_3__8 (
            que_out_2__3__8), .q_3__7 (que_out_2__3__7), .q_3__6 (
            que_out_2__3__6), .q_3__5 (que_out_2__3__5), .q_3__4 (
            que_out_2__3__4), .q_3__3 (que_out_2__3__3), .q_3__2 (
            que_out_2__3__2), .q_3__1 (que_out_2__3__1), .q_3__0 (
            que_out_2__3__0), .q_4__15 (que_out_2__4__15), .q_4__14 (
            que_out_2__4__14), .q_4__13 (que_out_2__4__13), .q_4__12 (
            que_out_2__4__12), .q_4__11 (que_out_2__4__11), .q_4__10 (
            que_out_2__4__10), .q_4__9 (que_out_2__4__9), .q_4__8 (
            que_out_2__4__8), .q_4__7 (que_out_2__4__7), .q_4__6 (
            que_out_2__4__6), .q_4__5 (que_out_2__4__5), .q_4__4 (
            que_out_2__4__4), .q_4__3 (que_out_2__4__3), .q_4__2 (
            que_out_2__4__2), .q_4__1 (que_out_2__4__1), .q_4__0 (
            que_out_2__4__0), .clk (nx10714), .load (sel_que_2), .reset (nx10690
            )) ;
    Queue_5 gen_queues_3_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_3__0__15), .q_0__14 (
            que_out_3__0__14), .q_0__13 (que_out_3__0__13), .q_0__12 (
            que_out_3__0__12), .q_0__11 (que_out_3__0__11), .q_0__10 (
            que_out_3__0__10), .q_0__9 (que_out_3__0__9), .q_0__8 (
            que_out_3__0__8), .q_0__7 (que_out_3__0__7), .q_0__6 (
            que_out_3__0__6), .q_0__5 (que_out_3__0__5), .q_0__4 (
            que_out_3__0__4), .q_0__3 (que_out_3__0__3), .q_0__2 (
            que_out_3__0__2), .q_0__1 (que_out_3__0__1), .q_0__0 (
            que_out_3__0__0), .q_1__15 (que_out_3__1__15), .q_1__14 (
            que_out_3__1__14), .q_1__13 (que_out_3__1__13), .q_1__12 (
            que_out_3__1__12), .q_1__11 (que_out_3__1__11), .q_1__10 (
            que_out_3__1__10), .q_1__9 (que_out_3__1__9), .q_1__8 (
            que_out_3__1__8), .q_1__7 (que_out_3__1__7), .q_1__6 (
            que_out_3__1__6), .q_1__5 (que_out_3__1__5), .q_1__4 (
            que_out_3__1__4), .q_1__3 (que_out_3__1__3), .q_1__2 (
            que_out_3__1__2), .q_1__1 (que_out_3__1__1), .q_1__0 (
            que_out_3__1__0), .q_2__15 (que_out_3__2__15), .q_2__14 (
            que_out_3__2__14), .q_2__13 (que_out_3__2__13), .q_2__12 (
            que_out_3__2__12), .q_2__11 (que_out_3__2__11), .q_2__10 (
            que_out_3__2__10), .q_2__9 (que_out_3__2__9), .q_2__8 (
            que_out_3__2__8), .q_2__7 (que_out_3__2__7), .q_2__6 (
            que_out_3__2__6), .q_2__5 (que_out_3__2__5), .q_2__4 (
            que_out_3__2__4), .q_2__3 (que_out_3__2__3), .q_2__2 (
            que_out_3__2__2), .q_2__1 (que_out_3__2__1), .q_2__0 (
            que_out_3__2__0), .q_3__15 (que_out_3__3__15), .q_3__14 (
            que_out_3__3__14), .q_3__13 (que_out_3__3__13), .q_3__12 (
            que_out_3__3__12), .q_3__11 (que_out_3__3__11), .q_3__10 (
            que_out_3__3__10), .q_3__9 (que_out_3__3__9), .q_3__8 (
            que_out_3__3__8), .q_3__7 (que_out_3__3__7), .q_3__6 (
            que_out_3__3__6), .q_3__5 (que_out_3__3__5), .q_3__4 (
            que_out_3__3__4), .q_3__3 (que_out_3__3__3), .q_3__2 (
            que_out_3__3__2), .q_3__1 (que_out_3__3__1), .q_3__0 (
            que_out_3__3__0), .q_4__15 (que_out_3__4__15), .q_4__14 (
            que_out_3__4__14), .q_4__13 (que_out_3__4__13), .q_4__12 (
            que_out_3__4__12), .q_4__11 (que_out_3__4__11), .q_4__10 (
            que_out_3__4__10), .q_4__9 (que_out_3__4__9), .q_4__8 (
            que_out_3__4__8), .q_4__7 (que_out_3__4__7), .q_4__6 (
            que_out_3__4__6), .q_4__5 (que_out_3__4__5), .q_4__4 (
            que_out_3__4__4), .q_4__3 (que_out_3__4__3), .q_4__2 (
            que_out_3__4__2), .q_4__1 (que_out_3__4__1), .q_4__0 (
            que_out_3__4__0), .clk (nx10716), .load (sel_que_3), .reset (nx10692
            )) ;
    Queue_5 gen_queues_4_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_4__0__15), .q_0__14 (
            que_out_4__0__14), .q_0__13 (que_out_4__0__13), .q_0__12 (
            que_out_4__0__12), .q_0__11 (que_out_4__0__11), .q_0__10 (
            que_out_4__0__10), .q_0__9 (que_out_4__0__9), .q_0__8 (
            que_out_4__0__8), .q_0__7 (que_out_4__0__7), .q_0__6 (
            que_out_4__0__6), .q_0__5 (que_out_4__0__5), .q_0__4 (
            que_out_4__0__4), .q_0__3 (que_out_4__0__3), .q_0__2 (
            que_out_4__0__2), .q_0__1 (que_out_4__0__1), .q_0__0 (
            que_out_4__0__0), .q_1__15 (que_out_4__1__15), .q_1__14 (
            que_out_4__1__14), .q_1__13 (que_out_4__1__13), .q_1__12 (
            que_out_4__1__12), .q_1__11 (que_out_4__1__11), .q_1__10 (
            que_out_4__1__10), .q_1__9 (que_out_4__1__9), .q_1__8 (
            que_out_4__1__8), .q_1__7 (que_out_4__1__7), .q_1__6 (
            que_out_4__1__6), .q_1__5 (que_out_4__1__5), .q_1__4 (
            que_out_4__1__4), .q_1__3 (que_out_4__1__3), .q_1__2 (
            que_out_4__1__2), .q_1__1 (que_out_4__1__1), .q_1__0 (
            que_out_4__1__0), .q_2__15 (que_out_4__2__15), .q_2__14 (
            que_out_4__2__14), .q_2__13 (que_out_4__2__13), .q_2__12 (
            que_out_4__2__12), .q_2__11 (que_out_4__2__11), .q_2__10 (
            que_out_4__2__10), .q_2__9 (que_out_4__2__9), .q_2__8 (
            que_out_4__2__8), .q_2__7 (que_out_4__2__7), .q_2__6 (
            que_out_4__2__6), .q_2__5 (que_out_4__2__5), .q_2__4 (
            que_out_4__2__4), .q_2__3 (que_out_4__2__3), .q_2__2 (
            que_out_4__2__2), .q_2__1 (que_out_4__2__1), .q_2__0 (
            que_out_4__2__0), .q_3__15 (que_out_4__3__15), .q_3__14 (
            que_out_4__3__14), .q_3__13 (que_out_4__3__13), .q_3__12 (
            que_out_4__3__12), .q_3__11 (que_out_4__3__11), .q_3__10 (
            que_out_4__3__10), .q_3__9 (que_out_4__3__9), .q_3__8 (
            que_out_4__3__8), .q_3__7 (que_out_4__3__7), .q_3__6 (
            que_out_4__3__6), .q_3__5 (que_out_4__3__5), .q_3__4 (
            que_out_4__3__4), .q_3__3 (que_out_4__3__3), .q_3__2 (
            que_out_4__3__2), .q_3__1 (que_out_4__3__1), .q_3__0 (
            que_out_4__3__0), .q_4__15 (que_out_4__4__15), .q_4__14 (
            que_out_4__4__14), .q_4__13 (que_out_4__4__13), .q_4__12 (
            que_out_4__4__12), .q_4__11 (que_out_4__4__11), .q_4__10 (
            que_out_4__4__10), .q_4__9 (que_out_4__4__9), .q_4__8 (
            que_out_4__4__8), .q_4__7 (que_out_4__4__7), .q_4__6 (
            que_out_4__4__6), .q_4__5 (que_out_4__4__5), .q_4__4 (
            que_out_4__4__4), .q_4__3 (que_out_4__4__3), .q_4__2 (
            que_out_4__4__2), .q_4__1 (que_out_4__4__1), .q_4__0 (
            que_out_4__4__0), .clk (nx10716), .load (sel_que_4), .reset (nx10692
            )) ;
    Queue_5 gen_queues_5_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_5__0__15), .q_0__14 (
            que_out_5__0__14), .q_0__13 (que_out_5__0__13), .q_0__12 (
            que_out_5__0__12), .q_0__11 (que_out_5__0__11), .q_0__10 (
            que_out_5__0__10), .q_0__9 (que_out_5__0__9), .q_0__8 (
            que_out_5__0__8), .q_0__7 (que_out_5__0__7), .q_0__6 (
            que_out_5__0__6), .q_0__5 (que_out_5__0__5), .q_0__4 (
            que_out_5__0__4), .q_0__3 (que_out_5__0__3), .q_0__2 (
            que_out_5__0__2), .q_0__1 (que_out_5__0__1), .q_0__0 (
            que_out_5__0__0), .q_1__15 (que_out_5__1__15), .q_1__14 (
            que_out_5__1__14), .q_1__13 (que_out_5__1__13), .q_1__12 (
            que_out_5__1__12), .q_1__11 (que_out_5__1__11), .q_1__10 (
            que_out_5__1__10), .q_1__9 (que_out_5__1__9), .q_1__8 (
            que_out_5__1__8), .q_1__7 (que_out_5__1__7), .q_1__6 (
            que_out_5__1__6), .q_1__5 (que_out_5__1__5), .q_1__4 (
            que_out_5__1__4), .q_1__3 (que_out_5__1__3), .q_1__2 (
            que_out_5__1__2), .q_1__1 (que_out_5__1__1), .q_1__0 (
            que_out_5__1__0), .q_2__15 (que_out_5__2__15), .q_2__14 (
            que_out_5__2__14), .q_2__13 (que_out_5__2__13), .q_2__12 (
            que_out_5__2__12), .q_2__11 (que_out_5__2__11), .q_2__10 (
            que_out_5__2__10), .q_2__9 (que_out_5__2__9), .q_2__8 (
            que_out_5__2__8), .q_2__7 (que_out_5__2__7), .q_2__6 (
            que_out_5__2__6), .q_2__5 (que_out_5__2__5), .q_2__4 (
            que_out_5__2__4), .q_2__3 (que_out_5__2__3), .q_2__2 (
            que_out_5__2__2), .q_2__1 (que_out_5__2__1), .q_2__0 (
            que_out_5__2__0), .q_3__15 (que_out_5__3__15), .q_3__14 (
            que_out_5__3__14), .q_3__13 (que_out_5__3__13), .q_3__12 (
            que_out_5__3__12), .q_3__11 (que_out_5__3__11), .q_3__10 (
            que_out_5__3__10), .q_3__9 (que_out_5__3__9), .q_3__8 (
            que_out_5__3__8), .q_3__7 (que_out_5__3__7), .q_3__6 (
            que_out_5__3__6), .q_3__5 (que_out_5__3__5), .q_3__4 (
            que_out_5__3__4), .q_3__3 (que_out_5__3__3), .q_3__2 (
            que_out_5__3__2), .q_3__1 (que_out_5__3__1), .q_3__0 (
            que_out_5__3__0), .q_4__15 (que_out_5__4__15), .q_4__14 (
            que_out_5__4__14), .q_4__13 (que_out_5__4__13), .q_4__12 (
            que_out_5__4__12), .q_4__11 (que_out_5__4__11), .q_4__10 (
            que_out_5__4__10), .q_4__9 (que_out_5__4__9), .q_4__8 (
            que_out_5__4__8), .q_4__7 (que_out_5__4__7), .q_4__6 (
            que_out_5__4__6), .q_4__5 (que_out_5__4__5), .q_4__4 (
            que_out_5__4__4), .q_4__3 (que_out_5__4__3), .q_4__2 (
            que_out_5__4__2), .q_4__1 (que_out_5__4__1), .q_4__0 (
            que_out_5__4__0), .clk (nx10716), .load (sel_que_5), .reset (nx10692
            )) ;
    Queue_5 gen_queues_6_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_6__0__15), .q_0__14 (
            que_out_6__0__14), .q_0__13 (que_out_6__0__13), .q_0__12 (
            que_out_6__0__12), .q_0__11 (que_out_6__0__11), .q_0__10 (
            que_out_6__0__10), .q_0__9 (que_out_6__0__9), .q_0__8 (
            que_out_6__0__8), .q_0__7 (que_out_6__0__7), .q_0__6 (
            que_out_6__0__6), .q_0__5 (que_out_6__0__5), .q_0__4 (
            que_out_6__0__4), .q_0__3 (que_out_6__0__3), .q_0__2 (
            que_out_6__0__2), .q_0__1 (que_out_6__0__1), .q_0__0 (
            que_out_6__0__0), .q_1__15 (que_out_6__1__15), .q_1__14 (
            que_out_6__1__14), .q_1__13 (que_out_6__1__13), .q_1__12 (
            que_out_6__1__12), .q_1__11 (que_out_6__1__11), .q_1__10 (
            que_out_6__1__10), .q_1__9 (que_out_6__1__9), .q_1__8 (
            que_out_6__1__8), .q_1__7 (que_out_6__1__7), .q_1__6 (
            que_out_6__1__6), .q_1__5 (que_out_6__1__5), .q_1__4 (
            que_out_6__1__4), .q_1__3 (que_out_6__1__3), .q_1__2 (
            que_out_6__1__2), .q_1__1 (que_out_6__1__1), .q_1__0 (
            que_out_6__1__0), .q_2__15 (que_out_6__2__15), .q_2__14 (
            que_out_6__2__14), .q_2__13 (que_out_6__2__13), .q_2__12 (
            que_out_6__2__12), .q_2__11 (que_out_6__2__11), .q_2__10 (
            que_out_6__2__10), .q_2__9 (que_out_6__2__9), .q_2__8 (
            que_out_6__2__8), .q_2__7 (que_out_6__2__7), .q_2__6 (
            que_out_6__2__6), .q_2__5 (que_out_6__2__5), .q_2__4 (
            que_out_6__2__4), .q_2__3 (que_out_6__2__3), .q_2__2 (
            que_out_6__2__2), .q_2__1 (que_out_6__2__1), .q_2__0 (
            que_out_6__2__0), .q_3__15 (que_out_6__3__15), .q_3__14 (
            que_out_6__3__14), .q_3__13 (que_out_6__3__13), .q_3__12 (
            que_out_6__3__12), .q_3__11 (que_out_6__3__11), .q_3__10 (
            que_out_6__3__10), .q_3__9 (que_out_6__3__9), .q_3__8 (
            que_out_6__3__8), .q_3__7 (que_out_6__3__7), .q_3__6 (
            que_out_6__3__6), .q_3__5 (que_out_6__3__5), .q_3__4 (
            que_out_6__3__4), .q_3__3 (que_out_6__3__3), .q_3__2 (
            que_out_6__3__2), .q_3__1 (que_out_6__3__1), .q_3__0 (
            que_out_6__3__0), .q_4__15 (que_out_6__4__15), .q_4__14 (
            que_out_6__4__14), .q_4__13 (que_out_6__4__13), .q_4__12 (
            que_out_6__4__12), .q_4__11 (que_out_6__4__11), .q_4__10 (
            que_out_6__4__10), .q_4__9 (que_out_6__4__9), .q_4__8 (
            que_out_6__4__8), .q_4__7 (que_out_6__4__7), .q_4__6 (
            que_out_6__4__6), .q_4__5 (que_out_6__4__5), .q_4__4 (
            que_out_6__4__4), .q_4__3 (que_out_6__4__3), .q_4__2 (
            que_out_6__4__2), .q_4__1 (que_out_6__4__1), .q_4__0 (
            que_out_6__4__0), .clk (nx10718), .load (sel_que_6), .reset (nx10694
            )) ;
    Queue_5 gen_queues_7_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_7__0__15), .q_0__14 (
            que_out_7__0__14), .q_0__13 (que_out_7__0__13), .q_0__12 (
            que_out_7__0__12), .q_0__11 (que_out_7__0__11), .q_0__10 (
            que_out_7__0__10), .q_0__9 (que_out_7__0__9), .q_0__8 (
            que_out_7__0__8), .q_0__7 (que_out_7__0__7), .q_0__6 (
            que_out_7__0__6), .q_0__5 (que_out_7__0__5), .q_0__4 (
            que_out_7__0__4), .q_0__3 (que_out_7__0__3), .q_0__2 (
            que_out_7__0__2), .q_0__1 (que_out_7__0__1), .q_0__0 (
            que_out_7__0__0), .q_1__15 (que_out_7__1__15), .q_1__14 (
            que_out_7__1__14), .q_1__13 (que_out_7__1__13), .q_1__12 (
            que_out_7__1__12), .q_1__11 (que_out_7__1__11), .q_1__10 (
            que_out_7__1__10), .q_1__9 (que_out_7__1__9), .q_1__8 (
            que_out_7__1__8), .q_1__7 (que_out_7__1__7), .q_1__6 (
            que_out_7__1__6), .q_1__5 (que_out_7__1__5), .q_1__4 (
            que_out_7__1__4), .q_1__3 (que_out_7__1__3), .q_1__2 (
            que_out_7__1__2), .q_1__1 (que_out_7__1__1), .q_1__0 (
            que_out_7__1__0), .q_2__15 (que_out_7__2__15), .q_2__14 (
            que_out_7__2__14), .q_2__13 (que_out_7__2__13), .q_2__12 (
            que_out_7__2__12), .q_2__11 (que_out_7__2__11), .q_2__10 (
            que_out_7__2__10), .q_2__9 (que_out_7__2__9), .q_2__8 (
            que_out_7__2__8), .q_2__7 (que_out_7__2__7), .q_2__6 (
            que_out_7__2__6), .q_2__5 (que_out_7__2__5), .q_2__4 (
            que_out_7__2__4), .q_2__3 (que_out_7__2__3), .q_2__2 (
            que_out_7__2__2), .q_2__1 (que_out_7__2__1), .q_2__0 (
            que_out_7__2__0), .q_3__15 (que_out_7__3__15), .q_3__14 (
            que_out_7__3__14), .q_3__13 (que_out_7__3__13), .q_3__12 (
            que_out_7__3__12), .q_3__11 (que_out_7__3__11), .q_3__10 (
            que_out_7__3__10), .q_3__9 (que_out_7__3__9), .q_3__8 (
            que_out_7__3__8), .q_3__7 (que_out_7__3__7), .q_3__6 (
            que_out_7__3__6), .q_3__5 (que_out_7__3__5), .q_3__4 (
            que_out_7__3__4), .q_3__3 (que_out_7__3__3), .q_3__2 (
            que_out_7__3__2), .q_3__1 (que_out_7__3__1), .q_3__0 (
            que_out_7__3__0), .q_4__15 (que_out_7__4__15), .q_4__14 (
            que_out_7__4__14), .q_4__13 (que_out_7__4__13), .q_4__12 (
            que_out_7__4__12), .q_4__11 (que_out_7__4__11), .q_4__10 (
            que_out_7__4__10), .q_4__9 (que_out_7__4__9), .q_4__8 (
            que_out_7__4__8), .q_4__7 (que_out_7__4__7), .q_4__6 (
            que_out_7__4__6), .q_4__5 (que_out_7__4__5), .q_4__4 (
            que_out_7__4__4), .q_4__3 (que_out_7__4__3), .q_4__2 (
            que_out_7__4__2), .q_4__1 (que_out_7__4__1), .q_4__0 (
            que_out_7__4__0), .clk (nx10720), .load (sel_que_7), .reset (nx10696
            )) ;
    Queue_5 gen_queues_8_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_8__0__15), .q_0__14 (
            que_out_8__0__14), .q_0__13 (que_out_8__0__13), .q_0__12 (
            que_out_8__0__12), .q_0__11 (que_out_8__0__11), .q_0__10 (
            que_out_8__0__10), .q_0__9 (que_out_8__0__9), .q_0__8 (
            que_out_8__0__8), .q_0__7 (que_out_8__0__7), .q_0__6 (
            que_out_8__0__6), .q_0__5 (que_out_8__0__5), .q_0__4 (
            que_out_8__0__4), .q_0__3 (que_out_8__0__3), .q_0__2 (
            que_out_8__0__2), .q_0__1 (que_out_8__0__1), .q_0__0 (
            que_out_8__0__0), .q_1__15 (que_out_8__1__15), .q_1__14 (
            que_out_8__1__14), .q_1__13 (que_out_8__1__13), .q_1__12 (
            que_out_8__1__12), .q_1__11 (que_out_8__1__11), .q_1__10 (
            que_out_8__1__10), .q_1__9 (que_out_8__1__9), .q_1__8 (
            que_out_8__1__8), .q_1__7 (que_out_8__1__7), .q_1__6 (
            que_out_8__1__6), .q_1__5 (que_out_8__1__5), .q_1__4 (
            que_out_8__1__4), .q_1__3 (que_out_8__1__3), .q_1__2 (
            que_out_8__1__2), .q_1__1 (que_out_8__1__1), .q_1__0 (
            que_out_8__1__0), .q_2__15 (que_out_8__2__15), .q_2__14 (
            que_out_8__2__14), .q_2__13 (que_out_8__2__13), .q_2__12 (
            que_out_8__2__12), .q_2__11 (que_out_8__2__11), .q_2__10 (
            que_out_8__2__10), .q_2__9 (que_out_8__2__9), .q_2__8 (
            que_out_8__2__8), .q_2__7 (que_out_8__2__7), .q_2__6 (
            que_out_8__2__6), .q_2__5 (que_out_8__2__5), .q_2__4 (
            que_out_8__2__4), .q_2__3 (que_out_8__2__3), .q_2__2 (
            que_out_8__2__2), .q_2__1 (que_out_8__2__1), .q_2__0 (
            que_out_8__2__0), .q_3__15 (que_out_8__3__15), .q_3__14 (
            que_out_8__3__14), .q_3__13 (que_out_8__3__13), .q_3__12 (
            que_out_8__3__12), .q_3__11 (que_out_8__3__11), .q_3__10 (
            que_out_8__3__10), .q_3__9 (que_out_8__3__9), .q_3__8 (
            que_out_8__3__8), .q_3__7 (que_out_8__3__7), .q_3__6 (
            que_out_8__3__6), .q_3__5 (que_out_8__3__5), .q_3__4 (
            que_out_8__3__4), .q_3__3 (que_out_8__3__3), .q_3__2 (
            que_out_8__3__2), .q_3__1 (que_out_8__3__1), .q_3__0 (
            que_out_8__3__0), .q_4__15 (que_out_8__4__15), .q_4__14 (
            que_out_8__4__14), .q_4__13 (que_out_8__4__13), .q_4__12 (
            que_out_8__4__12), .q_4__11 (que_out_8__4__11), .q_4__10 (
            que_out_8__4__10), .q_4__9 (que_out_8__4__9), .q_4__8 (
            que_out_8__4__8), .q_4__7 (que_out_8__4__7), .q_4__6 (
            que_out_8__4__6), .q_4__5 (que_out_8__4__5), .q_4__4 (
            que_out_8__4__4), .q_4__3 (que_out_8__4__3), .q_4__2 (
            que_out_8__4__2), .q_4__1 (que_out_8__4__1), .q_4__0 (
            que_out_8__4__0), .clk (nx10720), .load (sel_que_8), .reset (nx10696
            )) ;
    Queue_5 gen_queues_9_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_9__0__15), .q_0__14 (
            que_out_9__0__14), .q_0__13 (que_out_9__0__13), .q_0__12 (
            que_out_9__0__12), .q_0__11 (que_out_9__0__11), .q_0__10 (
            que_out_9__0__10), .q_0__9 (que_out_9__0__9), .q_0__8 (
            que_out_9__0__8), .q_0__7 (que_out_9__0__7), .q_0__6 (
            que_out_9__0__6), .q_0__5 (que_out_9__0__5), .q_0__4 (
            que_out_9__0__4), .q_0__3 (que_out_9__0__3), .q_0__2 (
            que_out_9__0__2), .q_0__1 (que_out_9__0__1), .q_0__0 (
            que_out_9__0__0), .q_1__15 (que_out_9__1__15), .q_1__14 (
            que_out_9__1__14), .q_1__13 (que_out_9__1__13), .q_1__12 (
            que_out_9__1__12), .q_1__11 (que_out_9__1__11), .q_1__10 (
            que_out_9__1__10), .q_1__9 (que_out_9__1__9), .q_1__8 (
            que_out_9__1__8), .q_1__7 (que_out_9__1__7), .q_1__6 (
            que_out_9__1__6), .q_1__5 (que_out_9__1__5), .q_1__4 (
            que_out_9__1__4), .q_1__3 (que_out_9__1__3), .q_1__2 (
            que_out_9__1__2), .q_1__1 (que_out_9__1__1), .q_1__0 (
            que_out_9__1__0), .q_2__15 (que_out_9__2__15), .q_2__14 (
            que_out_9__2__14), .q_2__13 (que_out_9__2__13), .q_2__12 (
            que_out_9__2__12), .q_2__11 (que_out_9__2__11), .q_2__10 (
            que_out_9__2__10), .q_2__9 (que_out_9__2__9), .q_2__8 (
            que_out_9__2__8), .q_2__7 (que_out_9__2__7), .q_2__6 (
            que_out_9__2__6), .q_2__5 (que_out_9__2__5), .q_2__4 (
            que_out_9__2__4), .q_2__3 (que_out_9__2__3), .q_2__2 (
            que_out_9__2__2), .q_2__1 (que_out_9__2__1), .q_2__0 (
            que_out_9__2__0), .q_3__15 (que_out_9__3__15), .q_3__14 (
            que_out_9__3__14), .q_3__13 (que_out_9__3__13), .q_3__12 (
            que_out_9__3__12), .q_3__11 (que_out_9__3__11), .q_3__10 (
            que_out_9__3__10), .q_3__9 (que_out_9__3__9), .q_3__8 (
            que_out_9__3__8), .q_3__7 (que_out_9__3__7), .q_3__6 (
            que_out_9__3__6), .q_3__5 (que_out_9__3__5), .q_3__4 (
            que_out_9__3__4), .q_3__3 (que_out_9__3__3), .q_3__2 (
            que_out_9__3__2), .q_3__1 (que_out_9__3__1), .q_3__0 (
            que_out_9__3__0), .q_4__15 (que_out_9__4__15), .q_4__14 (
            que_out_9__4__14), .q_4__13 (que_out_9__4__13), .q_4__12 (
            que_out_9__4__12), .q_4__11 (que_out_9__4__11), .q_4__10 (
            que_out_9__4__10), .q_4__9 (que_out_9__4__9), .q_4__8 (
            que_out_9__4__8), .q_4__7 (que_out_9__4__7), .q_4__6 (
            que_out_9__4__6), .q_4__5 (que_out_9__4__5), .q_4__4 (
            que_out_9__4__4), .q_4__3 (que_out_9__4__3), .q_4__2 (
            que_out_9__4__2), .q_4__1 (que_out_9__4__1), .q_4__0 (
            que_out_9__4__0), .clk (nx10720), .load (sel_que_9), .reset (nx10696
            )) ;
    Queue_5 gen_queues_10_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_10__0__15), .q_0__14 (
            que_out_10__0__14), .q_0__13 (que_out_10__0__13), .q_0__12 (
            que_out_10__0__12), .q_0__11 (que_out_10__0__11), .q_0__10 (
            que_out_10__0__10), .q_0__9 (que_out_10__0__9), .q_0__8 (
            que_out_10__0__8), .q_0__7 (que_out_10__0__7), .q_0__6 (
            que_out_10__0__6), .q_0__5 (que_out_10__0__5), .q_0__4 (
            que_out_10__0__4), .q_0__3 (que_out_10__0__3), .q_0__2 (
            que_out_10__0__2), .q_0__1 (que_out_10__0__1), .q_0__0 (
            que_out_10__0__0), .q_1__15 (que_out_10__1__15), .q_1__14 (
            que_out_10__1__14), .q_1__13 (que_out_10__1__13), .q_1__12 (
            que_out_10__1__12), .q_1__11 (que_out_10__1__11), .q_1__10 (
            que_out_10__1__10), .q_1__9 (que_out_10__1__9), .q_1__8 (
            que_out_10__1__8), .q_1__7 (que_out_10__1__7), .q_1__6 (
            que_out_10__1__6), .q_1__5 (que_out_10__1__5), .q_1__4 (
            que_out_10__1__4), .q_1__3 (que_out_10__1__3), .q_1__2 (
            que_out_10__1__2), .q_1__1 (que_out_10__1__1), .q_1__0 (
            que_out_10__1__0), .q_2__15 (que_out_10__2__15), .q_2__14 (
            que_out_10__2__14), .q_2__13 (que_out_10__2__13), .q_2__12 (
            que_out_10__2__12), .q_2__11 (que_out_10__2__11), .q_2__10 (
            que_out_10__2__10), .q_2__9 (que_out_10__2__9), .q_2__8 (
            que_out_10__2__8), .q_2__7 (que_out_10__2__7), .q_2__6 (
            que_out_10__2__6), .q_2__5 (que_out_10__2__5), .q_2__4 (
            que_out_10__2__4), .q_2__3 (que_out_10__2__3), .q_2__2 (
            que_out_10__2__2), .q_2__1 (que_out_10__2__1), .q_2__0 (
            que_out_10__2__0), .q_3__15 (que_out_10__3__15), .q_3__14 (
            que_out_10__3__14), .q_3__13 (que_out_10__3__13), .q_3__12 (
            que_out_10__3__12), .q_3__11 (que_out_10__3__11), .q_3__10 (
            que_out_10__3__10), .q_3__9 (que_out_10__3__9), .q_3__8 (
            que_out_10__3__8), .q_3__7 (que_out_10__3__7), .q_3__6 (
            que_out_10__3__6), .q_3__5 (que_out_10__3__5), .q_3__4 (
            que_out_10__3__4), .q_3__3 (que_out_10__3__3), .q_3__2 (
            que_out_10__3__2), .q_3__1 (que_out_10__3__1), .q_3__0 (
            que_out_10__3__0), .q_4__15 (que_out_10__4__15), .q_4__14 (
            que_out_10__4__14), .q_4__13 (que_out_10__4__13), .q_4__12 (
            que_out_10__4__12), .q_4__11 (que_out_10__4__11), .q_4__10 (
            que_out_10__4__10), .q_4__9 (que_out_10__4__9), .q_4__8 (
            que_out_10__4__8), .q_4__7 (que_out_10__4__7), .q_4__6 (
            que_out_10__4__6), .q_4__5 (que_out_10__4__5), .q_4__4 (
            que_out_10__4__4), .q_4__3 (que_out_10__4__3), .q_4__2 (
            que_out_10__4__2), .q_4__1 (que_out_10__4__1), .q_4__0 (
            que_out_10__4__0), .clk (nx10722), .load (sel_que_10), .reset (
            nx10698)) ;
    Queue_5 gen_queues_11_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_11__0__15), .q_0__14 (
            que_out_11__0__14), .q_0__13 (que_out_11__0__13), .q_0__12 (
            que_out_11__0__12), .q_0__11 (que_out_11__0__11), .q_0__10 (
            que_out_11__0__10), .q_0__9 (que_out_11__0__9), .q_0__8 (
            que_out_11__0__8), .q_0__7 (que_out_11__0__7), .q_0__6 (
            que_out_11__0__6), .q_0__5 (que_out_11__0__5), .q_0__4 (
            que_out_11__0__4), .q_0__3 (que_out_11__0__3), .q_0__2 (
            que_out_11__0__2), .q_0__1 (que_out_11__0__1), .q_0__0 (
            que_out_11__0__0), .q_1__15 (que_out_11__1__15), .q_1__14 (
            que_out_11__1__14), .q_1__13 (que_out_11__1__13), .q_1__12 (
            que_out_11__1__12), .q_1__11 (que_out_11__1__11), .q_1__10 (
            que_out_11__1__10), .q_1__9 (que_out_11__1__9), .q_1__8 (
            que_out_11__1__8), .q_1__7 (que_out_11__1__7), .q_1__6 (
            que_out_11__1__6), .q_1__5 (que_out_11__1__5), .q_1__4 (
            que_out_11__1__4), .q_1__3 (que_out_11__1__3), .q_1__2 (
            que_out_11__1__2), .q_1__1 (que_out_11__1__1), .q_1__0 (
            que_out_11__1__0), .q_2__15 (que_out_11__2__15), .q_2__14 (
            que_out_11__2__14), .q_2__13 (que_out_11__2__13), .q_2__12 (
            que_out_11__2__12), .q_2__11 (que_out_11__2__11), .q_2__10 (
            que_out_11__2__10), .q_2__9 (que_out_11__2__9), .q_2__8 (
            que_out_11__2__8), .q_2__7 (que_out_11__2__7), .q_2__6 (
            que_out_11__2__6), .q_2__5 (que_out_11__2__5), .q_2__4 (
            que_out_11__2__4), .q_2__3 (que_out_11__2__3), .q_2__2 (
            que_out_11__2__2), .q_2__1 (que_out_11__2__1), .q_2__0 (
            que_out_11__2__0), .q_3__15 (que_out_11__3__15), .q_3__14 (
            que_out_11__3__14), .q_3__13 (que_out_11__3__13), .q_3__12 (
            que_out_11__3__12), .q_3__11 (que_out_11__3__11), .q_3__10 (
            que_out_11__3__10), .q_3__9 (que_out_11__3__9), .q_3__8 (
            que_out_11__3__8), .q_3__7 (que_out_11__3__7), .q_3__6 (
            que_out_11__3__6), .q_3__5 (que_out_11__3__5), .q_3__4 (
            que_out_11__3__4), .q_3__3 (que_out_11__3__3), .q_3__2 (
            que_out_11__3__2), .q_3__1 (que_out_11__3__1), .q_3__0 (
            que_out_11__3__0), .q_4__15 (que_out_11__4__15), .q_4__14 (
            que_out_11__4__14), .q_4__13 (que_out_11__4__13), .q_4__12 (
            que_out_11__4__12), .q_4__11 (que_out_11__4__11), .q_4__10 (
            que_out_11__4__10), .q_4__9 (que_out_11__4__9), .q_4__8 (
            que_out_11__4__8), .q_4__7 (que_out_11__4__7), .q_4__6 (
            que_out_11__4__6), .q_4__5 (que_out_11__4__5), .q_4__4 (
            que_out_11__4__4), .q_4__3 (que_out_11__4__3), .q_4__2 (
            que_out_11__4__2), .q_4__1 (que_out_11__4__1), .q_4__0 (
            que_out_11__4__0), .clk (nx10722), .load (sel_que_11), .reset (
            nx10698)) ;
    Queue_5 gen_queues_12_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_12__0__15), .q_0__14 (
            que_out_12__0__14), .q_0__13 (que_out_12__0__13), .q_0__12 (
            que_out_12__0__12), .q_0__11 (que_out_12__0__11), .q_0__10 (
            que_out_12__0__10), .q_0__9 (que_out_12__0__9), .q_0__8 (
            que_out_12__0__8), .q_0__7 (que_out_12__0__7), .q_0__6 (
            que_out_12__0__6), .q_0__5 (que_out_12__0__5), .q_0__4 (
            que_out_12__0__4), .q_0__3 (que_out_12__0__3), .q_0__2 (
            que_out_12__0__2), .q_0__1 (que_out_12__0__1), .q_0__0 (
            que_out_12__0__0), .q_1__15 (que_out_12__1__15), .q_1__14 (
            que_out_12__1__14), .q_1__13 (que_out_12__1__13), .q_1__12 (
            que_out_12__1__12), .q_1__11 (que_out_12__1__11), .q_1__10 (
            que_out_12__1__10), .q_1__9 (que_out_12__1__9), .q_1__8 (
            que_out_12__1__8), .q_1__7 (que_out_12__1__7), .q_1__6 (
            que_out_12__1__6), .q_1__5 (que_out_12__1__5), .q_1__4 (
            que_out_12__1__4), .q_1__3 (que_out_12__1__3), .q_1__2 (
            que_out_12__1__2), .q_1__1 (que_out_12__1__1), .q_1__0 (
            que_out_12__1__0), .q_2__15 (que_out_12__2__15), .q_2__14 (
            que_out_12__2__14), .q_2__13 (que_out_12__2__13), .q_2__12 (
            que_out_12__2__12), .q_2__11 (que_out_12__2__11), .q_2__10 (
            que_out_12__2__10), .q_2__9 (que_out_12__2__9), .q_2__8 (
            que_out_12__2__8), .q_2__7 (que_out_12__2__7), .q_2__6 (
            que_out_12__2__6), .q_2__5 (que_out_12__2__5), .q_2__4 (
            que_out_12__2__4), .q_2__3 (que_out_12__2__3), .q_2__2 (
            que_out_12__2__2), .q_2__1 (que_out_12__2__1), .q_2__0 (
            que_out_12__2__0), .q_3__15 (que_out_12__3__15), .q_3__14 (
            que_out_12__3__14), .q_3__13 (que_out_12__3__13), .q_3__12 (
            que_out_12__3__12), .q_3__11 (que_out_12__3__11), .q_3__10 (
            que_out_12__3__10), .q_3__9 (que_out_12__3__9), .q_3__8 (
            que_out_12__3__8), .q_3__7 (que_out_12__3__7), .q_3__6 (
            que_out_12__3__6), .q_3__5 (que_out_12__3__5), .q_3__4 (
            que_out_12__3__4), .q_3__3 (que_out_12__3__3), .q_3__2 (
            que_out_12__3__2), .q_3__1 (que_out_12__3__1), .q_3__0 (
            que_out_12__3__0), .q_4__15 (que_out_12__4__15), .q_4__14 (
            que_out_12__4__14), .q_4__13 (que_out_12__4__13), .q_4__12 (
            que_out_12__4__12), .q_4__11 (que_out_12__4__11), .q_4__10 (
            que_out_12__4__10), .q_4__9 (que_out_12__4__9), .q_4__8 (
            que_out_12__4__8), .q_4__7 (que_out_12__4__7), .q_4__6 (
            que_out_12__4__6), .q_4__5 (que_out_12__4__5), .q_4__4 (
            que_out_12__4__4), .q_4__3 (que_out_12__4__3), .q_4__2 (
            que_out_12__4__2), .q_4__1 (que_out_12__4__1), .q_4__0 (
            que_out_12__4__0), .clk (nx10722), .load (sel_que_12), .reset (
            nx10698)) ;
    Queue_5 gen_queues_13_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_13__0__15), .q_0__14 (
            que_out_13__0__14), .q_0__13 (que_out_13__0__13), .q_0__12 (
            que_out_13__0__12), .q_0__11 (que_out_13__0__11), .q_0__10 (
            que_out_13__0__10), .q_0__9 (que_out_13__0__9), .q_0__8 (
            que_out_13__0__8), .q_0__7 (que_out_13__0__7), .q_0__6 (
            que_out_13__0__6), .q_0__5 (que_out_13__0__5), .q_0__4 (
            que_out_13__0__4), .q_0__3 (que_out_13__0__3), .q_0__2 (
            que_out_13__0__2), .q_0__1 (que_out_13__0__1), .q_0__0 (
            que_out_13__0__0), .q_1__15 (que_out_13__1__15), .q_1__14 (
            que_out_13__1__14), .q_1__13 (que_out_13__1__13), .q_1__12 (
            que_out_13__1__12), .q_1__11 (que_out_13__1__11), .q_1__10 (
            que_out_13__1__10), .q_1__9 (que_out_13__1__9), .q_1__8 (
            que_out_13__1__8), .q_1__7 (que_out_13__1__7), .q_1__6 (
            que_out_13__1__6), .q_1__5 (que_out_13__1__5), .q_1__4 (
            que_out_13__1__4), .q_1__3 (que_out_13__1__3), .q_1__2 (
            que_out_13__1__2), .q_1__1 (que_out_13__1__1), .q_1__0 (
            que_out_13__1__0), .q_2__15 (que_out_13__2__15), .q_2__14 (
            que_out_13__2__14), .q_2__13 (que_out_13__2__13), .q_2__12 (
            que_out_13__2__12), .q_2__11 (que_out_13__2__11), .q_2__10 (
            que_out_13__2__10), .q_2__9 (que_out_13__2__9), .q_2__8 (
            que_out_13__2__8), .q_2__7 (que_out_13__2__7), .q_2__6 (
            que_out_13__2__6), .q_2__5 (que_out_13__2__5), .q_2__4 (
            que_out_13__2__4), .q_2__3 (que_out_13__2__3), .q_2__2 (
            que_out_13__2__2), .q_2__1 (que_out_13__2__1), .q_2__0 (
            que_out_13__2__0), .q_3__15 (que_out_13__3__15), .q_3__14 (
            que_out_13__3__14), .q_3__13 (que_out_13__3__13), .q_3__12 (
            que_out_13__3__12), .q_3__11 (que_out_13__3__11), .q_3__10 (
            que_out_13__3__10), .q_3__9 (que_out_13__3__9), .q_3__8 (
            que_out_13__3__8), .q_3__7 (que_out_13__3__7), .q_3__6 (
            que_out_13__3__6), .q_3__5 (que_out_13__3__5), .q_3__4 (
            que_out_13__3__4), .q_3__3 (que_out_13__3__3), .q_3__2 (
            que_out_13__3__2), .q_3__1 (que_out_13__3__1), .q_3__0 (
            que_out_13__3__0), .q_4__15 (que_out_13__4__15), .q_4__14 (
            que_out_13__4__14), .q_4__13 (que_out_13__4__13), .q_4__12 (
            que_out_13__4__12), .q_4__11 (que_out_13__4__11), .q_4__10 (
            que_out_13__4__10), .q_4__9 (que_out_13__4__9), .q_4__8 (
            que_out_13__4__8), .q_4__7 (que_out_13__4__7), .q_4__6 (
            que_out_13__4__6), .q_4__5 (que_out_13__4__5), .q_4__4 (
            que_out_13__4__4), .q_4__3 (que_out_13__4__3), .q_4__2 (
            que_out_13__4__2), .q_4__1 (que_out_13__4__1), .q_4__0 (
            que_out_13__4__0), .clk (nx10724), .load (sel_que_13), .reset (
            nx10700)) ;
    Queue_5 gen_queues_14_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_14__0__15), .q_0__14 (
            que_out_14__0__14), .q_0__13 (que_out_14__0__13), .q_0__12 (
            que_out_14__0__12), .q_0__11 (que_out_14__0__11), .q_0__10 (
            que_out_14__0__10), .q_0__9 (que_out_14__0__9), .q_0__8 (
            que_out_14__0__8), .q_0__7 (que_out_14__0__7), .q_0__6 (
            que_out_14__0__6), .q_0__5 (que_out_14__0__5), .q_0__4 (
            que_out_14__0__4), .q_0__3 (que_out_14__0__3), .q_0__2 (
            que_out_14__0__2), .q_0__1 (que_out_14__0__1), .q_0__0 (
            que_out_14__0__0), .q_1__15 (que_out_14__1__15), .q_1__14 (
            que_out_14__1__14), .q_1__13 (que_out_14__1__13), .q_1__12 (
            que_out_14__1__12), .q_1__11 (que_out_14__1__11), .q_1__10 (
            que_out_14__1__10), .q_1__9 (que_out_14__1__9), .q_1__8 (
            que_out_14__1__8), .q_1__7 (que_out_14__1__7), .q_1__6 (
            que_out_14__1__6), .q_1__5 (que_out_14__1__5), .q_1__4 (
            que_out_14__1__4), .q_1__3 (que_out_14__1__3), .q_1__2 (
            que_out_14__1__2), .q_1__1 (que_out_14__1__1), .q_1__0 (
            que_out_14__1__0), .q_2__15 (que_out_14__2__15), .q_2__14 (
            que_out_14__2__14), .q_2__13 (que_out_14__2__13), .q_2__12 (
            que_out_14__2__12), .q_2__11 (que_out_14__2__11), .q_2__10 (
            que_out_14__2__10), .q_2__9 (que_out_14__2__9), .q_2__8 (
            que_out_14__2__8), .q_2__7 (que_out_14__2__7), .q_2__6 (
            que_out_14__2__6), .q_2__5 (que_out_14__2__5), .q_2__4 (
            que_out_14__2__4), .q_2__3 (que_out_14__2__3), .q_2__2 (
            que_out_14__2__2), .q_2__1 (que_out_14__2__1), .q_2__0 (
            que_out_14__2__0), .q_3__15 (que_out_14__3__15), .q_3__14 (
            que_out_14__3__14), .q_3__13 (que_out_14__3__13), .q_3__12 (
            que_out_14__3__12), .q_3__11 (que_out_14__3__11), .q_3__10 (
            que_out_14__3__10), .q_3__9 (que_out_14__3__9), .q_3__8 (
            que_out_14__3__8), .q_3__7 (que_out_14__3__7), .q_3__6 (
            que_out_14__3__6), .q_3__5 (que_out_14__3__5), .q_3__4 (
            que_out_14__3__4), .q_3__3 (que_out_14__3__3), .q_3__2 (
            que_out_14__3__2), .q_3__1 (que_out_14__3__1), .q_3__0 (
            que_out_14__3__0), .q_4__15 (que_out_14__4__15), .q_4__14 (
            que_out_14__4__14), .q_4__13 (que_out_14__4__13), .q_4__12 (
            que_out_14__4__12), .q_4__11 (que_out_14__4__11), .q_4__10 (
            que_out_14__4__10), .q_4__9 (que_out_14__4__9), .q_4__8 (
            que_out_14__4__8), .q_4__7 (que_out_14__4__7), .q_4__6 (
            que_out_14__4__6), .q_4__5 (que_out_14__4__5), .q_4__4 (
            que_out_14__4__4), .q_4__3 (que_out_14__4__3), .q_4__2 (
            que_out_14__4__2), .q_4__1 (que_out_14__4__1), .q_4__0 (
            que_out_14__4__0), .clk (nx10726), .load (sel_que_14), .reset (
            nx10702)) ;
    Queue_5 gen_queues_15_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_15__0__15), .q_0__14 (
            que_out_15__0__14), .q_0__13 (que_out_15__0__13), .q_0__12 (
            que_out_15__0__12), .q_0__11 (que_out_15__0__11), .q_0__10 (
            que_out_15__0__10), .q_0__9 (que_out_15__0__9), .q_0__8 (
            que_out_15__0__8), .q_0__7 (que_out_15__0__7), .q_0__6 (
            que_out_15__0__6), .q_0__5 (que_out_15__0__5), .q_0__4 (
            que_out_15__0__4), .q_0__3 (que_out_15__0__3), .q_0__2 (
            que_out_15__0__2), .q_0__1 (que_out_15__0__1), .q_0__0 (
            que_out_15__0__0), .q_1__15 (que_out_15__1__15), .q_1__14 (
            que_out_15__1__14), .q_1__13 (que_out_15__1__13), .q_1__12 (
            que_out_15__1__12), .q_1__11 (que_out_15__1__11), .q_1__10 (
            que_out_15__1__10), .q_1__9 (que_out_15__1__9), .q_1__8 (
            que_out_15__1__8), .q_1__7 (que_out_15__1__7), .q_1__6 (
            que_out_15__1__6), .q_1__5 (que_out_15__1__5), .q_1__4 (
            que_out_15__1__4), .q_1__3 (que_out_15__1__3), .q_1__2 (
            que_out_15__1__2), .q_1__1 (que_out_15__1__1), .q_1__0 (
            que_out_15__1__0), .q_2__15 (que_out_15__2__15), .q_2__14 (
            que_out_15__2__14), .q_2__13 (que_out_15__2__13), .q_2__12 (
            que_out_15__2__12), .q_2__11 (que_out_15__2__11), .q_2__10 (
            que_out_15__2__10), .q_2__9 (que_out_15__2__9), .q_2__8 (
            que_out_15__2__8), .q_2__7 (que_out_15__2__7), .q_2__6 (
            que_out_15__2__6), .q_2__5 (que_out_15__2__5), .q_2__4 (
            que_out_15__2__4), .q_2__3 (que_out_15__2__3), .q_2__2 (
            que_out_15__2__2), .q_2__1 (que_out_15__2__1), .q_2__0 (
            que_out_15__2__0), .q_3__15 (que_out_15__3__15), .q_3__14 (
            que_out_15__3__14), .q_3__13 (que_out_15__3__13), .q_3__12 (
            que_out_15__3__12), .q_3__11 (que_out_15__3__11), .q_3__10 (
            que_out_15__3__10), .q_3__9 (que_out_15__3__9), .q_3__8 (
            que_out_15__3__8), .q_3__7 (que_out_15__3__7), .q_3__6 (
            que_out_15__3__6), .q_3__5 (que_out_15__3__5), .q_3__4 (
            que_out_15__3__4), .q_3__3 (que_out_15__3__3), .q_3__2 (
            que_out_15__3__2), .q_3__1 (que_out_15__3__1), .q_3__0 (
            que_out_15__3__0), .q_4__15 (que_out_15__4__15), .q_4__14 (
            que_out_15__4__14), .q_4__13 (que_out_15__4__13), .q_4__12 (
            que_out_15__4__12), .q_4__11 (que_out_15__4__11), .q_4__10 (
            que_out_15__4__10), .q_4__9 (que_out_15__4__9), .q_4__8 (
            que_out_15__4__8), .q_4__7 (que_out_15__4__7), .q_4__6 (
            que_out_15__4__6), .q_4__5 (que_out_15__4__5), .q_4__4 (
            que_out_15__4__4), .q_4__3 (que_out_15__4__3), .q_4__2 (
            que_out_15__4__2), .q_4__1 (que_out_15__4__1), .q_4__0 (
            que_out_15__4__0), .clk (nx10726), .load (sel_que_15), .reset (
            nx10702)) ;
    Queue_5 gen_queues_16_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_16__0__15), .q_0__14 (
            que_out_16__0__14), .q_0__13 (que_out_16__0__13), .q_0__12 (
            que_out_16__0__12), .q_0__11 (que_out_16__0__11), .q_0__10 (
            que_out_16__0__10), .q_0__9 (que_out_16__0__9), .q_0__8 (
            que_out_16__0__8), .q_0__7 (que_out_16__0__7), .q_0__6 (
            que_out_16__0__6), .q_0__5 (que_out_16__0__5), .q_0__4 (
            que_out_16__0__4), .q_0__3 (que_out_16__0__3), .q_0__2 (
            que_out_16__0__2), .q_0__1 (que_out_16__0__1), .q_0__0 (
            que_out_16__0__0), .q_1__15 (que_out_16__1__15), .q_1__14 (
            que_out_16__1__14), .q_1__13 (que_out_16__1__13), .q_1__12 (
            que_out_16__1__12), .q_1__11 (que_out_16__1__11), .q_1__10 (
            que_out_16__1__10), .q_1__9 (que_out_16__1__9), .q_1__8 (
            que_out_16__1__8), .q_1__7 (que_out_16__1__7), .q_1__6 (
            que_out_16__1__6), .q_1__5 (que_out_16__1__5), .q_1__4 (
            que_out_16__1__4), .q_1__3 (que_out_16__1__3), .q_1__2 (
            que_out_16__1__2), .q_1__1 (que_out_16__1__1), .q_1__0 (
            que_out_16__1__0), .q_2__15 (que_out_16__2__15), .q_2__14 (
            que_out_16__2__14), .q_2__13 (que_out_16__2__13), .q_2__12 (
            que_out_16__2__12), .q_2__11 (que_out_16__2__11), .q_2__10 (
            que_out_16__2__10), .q_2__9 (que_out_16__2__9), .q_2__8 (
            que_out_16__2__8), .q_2__7 (que_out_16__2__7), .q_2__6 (
            que_out_16__2__6), .q_2__5 (que_out_16__2__5), .q_2__4 (
            que_out_16__2__4), .q_2__3 (que_out_16__2__3), .q_2__2 (
            que_out_16__2__2), .q_2__1 (que_out_16__2__1), .q_2__0 (
            que_out_16__2__0), .q_3__15 (que_out_16__3__15), .q_3__14 (
            que_out_16__3__14), .q_3__13 (que_out_16__3__13), .q_3__12 (
            que_out_16__3__12), .q_3__11 (que_out_16__3__11), .q_3__10 (
            que_out_16__3__10), .q_3__9 (que_out_16__3__9), .q_3__8 (
            que_out_16__3__8), .q_3__7 (que_out_16__3__7), .q_3__6 (
            que_out_16__3__6), .q_3__5 (que_out_16__3__5), .q_3__4 (
            que_out_16__3__4), .q_3__3 (que_out_16__3__3), .q_3__2 (
            que_out_16__3__2), .q_3__1 (que_out_16__3__1), .q_3__0 (
            que_out_16__3__0), .q_4__15 (que_out_16__4__15), .q_4__14 (
            que_out_16__4__14), .q_4__13 (que_out_16__4__13), .q_4__12 (
            que_out_16__4__12), .q_4__11 (que_out_16__4__11), .q_4__10 (
            que_out_16__4__10), .q_4__9 (que_out_16__4__9), .q_4__8 (
            que_out_16__4__8), .q_4__7 (que_out_16__4__7), .q_4__6 (
            que_out_16__4__6), .q_4__5 (que_out_16__4__5), .q_4__4 (
            que_out_16__4__4), .q_4__3 (que_out_16__4__3), .q_4__2 (
            que_out_16__4__2), .q_4__1 (que_out_16__4__1), .q_4__0 (
            que_out_16__4__0), .clk (nx10726), .load (sel_que_16), .reset (
            nx10702)) ;
    Queue_5 gen_queues_17_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_17__0__15), .q_0__14 (
            que_out_17__0__14), .q_0__13 (que_out_17__0__13), .q_0__12 (
            que_out_17__0__12), .q_0__11 (que_out_17__0__11), .q_0__10 (
            que_out_17__0__10), .q_0__9 (que_out_17__0__9), .q_0__8 (
            que_out_17__0__8), .q_0__7 (que_out_17__0__7), .q_0__6 (
            que_out_17__0__6), .q_0__5 (que_out_17__0__5), .q_0__4 (
            que_out_17__0__4), .q_0__3 (que_out_17__0__3), .q_0__2 (
            que_out_17__0__2), .q_0__1 (que_out_17__0__1), .q_0__0 (
            que_out_17__0__0), .q_1__15 (que_out_17__1__15), .q_1__14 (
            que_out_17__1__14), .q_1__13 (que_out_17__1__13), .q_1__12 (
            que_out_17__1__12), .q_1__11 (que_out_17__1__11), .q_1__10 (
            que_out_17__1__10), .q_1__9 (que_out_17__1__9), .q_1__8 (
            que_out_17__1__8), .q_1__7 (que_out_17__1__7), .q_1__6 (
            que_out_17__1__6), .q_1__5 (que_out_17__1__5), .q_1__4 (
            que_out_17__1__4), .q_1__3 (que_out_17__1__3), .q_1__2 (
            que_out_17__1__2), .q_1__1 (que_out_17__1__1), .q_1__0 (
            que_out_17__1__0), .q_2__15 (que_out_17__2__15), .q_2__14 (
            que_out_17__2__14), .q_2__13 (que_out_17__2__13), .q_2__12 (
            que_out_17__2__12), .q_2__11 (que_out_17__2__11), .q_2__10 (
            que_out_17__2__10), .q_2__9 (que_out_17__2__9), .q_2__8 (
            que_out_17__2__8), .q_2__7 (que_out_17__2__7), .q_2__6 (
            que_out_17__2__6), .q_2__5 (que_out_17__2__5), .q_2__4 (
            que_out_17__2__4), .q_2__3 (que_out_17__2__3), .q_2__2 (
            que_out_17__2__2), .q_2__1 (que_out_17__2__1), .q_2__0 (
            que_out_17__2__0), .q_3__15 (que_out_17__3__15), .q_3__14 (
            que_out_17__3__14), .q_3__13 (que_out_17__3__13), .q_3__12 (
            que_out_17__3__12), .q_3__11 (que_out_17__3__11), .q_3__10 (
            que_out_17__3__10), .q_3__9 (que_out_17__3__9), .q_3__8 (
            que_out_17__3__8), .q_3__7 (que_out_17__3__7), .q_3__6 (
            que_out_17__3__6), .q_3__5 (que_out_17__3__5), .q_3__4 (
            que_out_17__3__4), .q_3__3 (que_out_17__3__3), .q_3__2 (
            que_out_17__3__2), .q_3__1 (que_out_17__3__1), .q_3__0 (
            que_out_17__3__0), .q_4__15 (que_out_17__4__15), .q_4__14 (
            que_out_17__4__14), .q_4__13 (que_out_17__4__13), .q_4__12 (
            que_out_17__4__12), .q_4__11 (que_out_17__4__11), .q_4__10 (
            que_out_17__4__10), .q_4__9 (que_out_17__4__9), .q_4__8 (
            que_out_17__4__8), .q_4__7 (que_out_17__4__7), .q_4__6 (
            que_out_17__4__6), .q_4__5 (que_out_17__4__5), .q_4__4 (
            que_out_17__4__4), .q_4__3 (que_out_17__4__3), .q_4__2 (
            que_out_17__4__2), .q_4__1 (que_out_17__4__1), .q_4__0 (
            que_out_17__4__0), .clk (nx10728), .load (sel_que_17), .reset (
            nx10704)) ;
    Queue_5 gen_queues_18_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_18__0__15), .q_0__14 (
            que_out_18__0__14), .q_0__13 (que_out_18__0__13), .q_0__12 (
            que_out_18__0__12), .q_0__11 (que_out_18__0__11), .q_0__10 (
            que_out_18__0__10), .q_0__9 (que_out_18__0__9), .q_0__8 (
            que_out_18__0__8), .q_0__7 (que_out_18__0__7), .q_0__6 (
            que_out_18__0__6), .q_0__5 (que_out_18__0__5), .q_0__4 (
            que_out_18__0__4), .q_0__3 (que_out_18__0__3), .q_0__2 (
            que_out_18__0__2), .q_0__1 (que_out_18__0__1), .q_0__0 (
            que_out_18__0__0), .q_1__15 (que_out_18__1__15), .q_1__14 (
            que_out_18__1__14), .q_1__13 (que_out_18__1__13), .q_1__12 (
            que_out_18__1__12), .q_1__11 (que_out_18__1__11), .q_1__10 (
            que_out_18__1__10), .q_1__9 (que_out_18__1__9), .q_1__8 (
            que_out_18__1__8), .q_1__7 (que_out_18__1__7), .q_1__6 (
            que_out_18__1__6), .q_1__5 (que_out_18__1__5), .q_1__4 (
            que_out_18__1__4), .q_1__3 (que_out_18__1__3), .q_1__2 (
            que_out_18__1__2), .q_1__1 (que_out_18__1__1), .q_1__0 (
            que_out_18__1__0), .q_2__15 (que_out_18__2__15), .q_2__14 (
            que_out_18__2__14), .q_2__13 (que_out_18__2__13), .q_2__12 (
            que_out_18__2__12), .q_2__11 (que_out_18__2__11), .q_2__10 (
            que_out_18__2__10), .q_2__9 (que_out_18__2__9), .q_2__8 (
            que_out_18__2__8), .q_2__7 (que_out_18__2__7), .q_2__6 (
            que_out_18__2__6), .q_2__5 (que_out_18__2__5), .q_2__4 (
            que_out_18__2__4), .q_2__3 (que_out_18__2__3), .q_2__2 (
            que_out_18__2__2), .q_2__1 (que_out_18__2__1), .q_2__0 (
            que_out_18__2__0), .q_3__15 (que_out_18__3__15), .q_3__14 (
            que_out_18__3__14), .q_3__13 (que_out_18__3__13), .q_3__12 (
            que_out_18__3__12), .q_3__11 (que_out_18__3__11), .q_3__10 (
            que_out_18__3__10), .q_3__9 (que_out_18__3__9), .q_3__8 (
            que_out_18__3__8), .q_3__7 (que_out_18__3__7), .q_3__6 (
            que_out_18__3__6), .q_3__5 (que_out_18__3__5), .q_3__4 (
            que_out_18__3__4), .q_3__3 (que_out_18__3__3), .q_3__2 (
            que_out_18__3__2), .q_3__1 (que_out_18__3__1), .q_3__0 (
            que_out_18__3__0), .q_4__15 (que_out_18__4__15), .q_4__14 (
            que_out_18__4__14), .q_4__13 (que_out_18__4__13), .q_4__12 (
            que_out_18__4__12), .q_4__11 (que_out_18__4__11), .q_4__10 (
            que_out_18__4__10), .q_4__9 (que_out_18__4__9), .q_4__8 (
            que_out_18__4__8), .q_4__7 (que_out_18__4__7), .q_4__6 (
            que_out_18__4__6), .q_4__5 (que_out_18__4__5), .q_4__4 (
            que_out_18__4__4), .q_4__3 (que_out_18__4__3), .q_4__2 (
            que_out_18__4__2), .q_4__1 (que_out_18__4__1), .q_4__0 (
            que_out_18__4__0), .clk (nx10728), .load (sel_que_18), .reset (
            nx10704)) ;
    Queue_5 gen_queues_19_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_19__0__15), .q_0__14 (
            que_out_19__0__14), .q_0__13 (que_out_19__0__13), .q_0__12 (
            que_out_19__0__12), .q_0__11 (que_out_19__0__11), .q_0__10 (
            que_out_19__0__10), .q_0__9 (que_out_19__0__9), .q_0__8 (
            que_out_19__0__8), .q_0__7 (que_out_19__0__7), .q_0__6 (
            que_out_19__0__6), .q_0__5 (que_out_19__0__5), .q_0__4 (
            que_out_19__0__4), .q_0__3 (que_out_19__0__3), .q_0__2 (
            que_out_19__0__2), .q_0__1 (que_out_19__0__1), .q_0__0 (
            que_out_19__0__0), .q_1__15 (que_out_19__1__15), .q_1__14 (
            que_out_19__1__14), .q_1__13 (que_out_19__1__13), .q_1__12 (
            que_out_19__1__12), .q_1__11 (que_out_19__1__11), .q_1__10 (
            que_out_19__1__10), .q_1__9 (que_out_19__1__9), .q_1__8 (
            que_out_19__1__8), .q_1__7 (que_out_19__1__7), .q_1__6 (
            que_out_19__1__6), .q_1__5 (que_out_19__1__5), .q_1__4 (
            que_out_19__1__4), .q_1__3 (que_out_19__1__3), .q_1__2 (
            que_out_19__1__2), .q_1__1 (que_out_19__1__1), .q_1__0 (
            que_out_19__1__0), .q_2__15 (que_out_19__2__15), .q_2__14 (
            que_out_19__2__14), .q_2__13 (que_out_19__2__13), .q_2__12 (
            que_out_19__2__12), .q_2__11 (que_out_19__2__11), .q_2__10 (
            que_out_19__2__10), .q_2__9 (que_out_19__2__9), .q_2__8 (
            que_out_19__2__8), .q_2__7 (que_out_19__2__7), .q_2__6 (
            que_out_19__2__6), .q_2__5 (que_out_19__2__5), .q_2__4 (
            que_out_19__2__4), .q_2__3 (que_out_19__2__3), .q_2__2 (
            que_out_19__2__2), .q_2__1 (que_out_19__2__1), .q_2__0 (
            que_out_19__2__0), .q_3__15 (que_out_19__3__15), .q_3__14 (
            que_out_19__3__14), .q_3__13 (que_out_19__3__13), .q_3__12 (
            que_out_19__3__12), .q_3__11 (que_out_19__3__11), .q_3__10 (
            que_out_19__3__10), .q_3__9 (que_out_19__3__9), .q_3__8 (
            que_out_19__3__8), .q_3__7 (que_out_19__3__7), .q_3__6 (
            que_out_19__3__6), .q_3__5 (que_out_19__3__5), .q_3__4 (
            que_out_19__3__4), .q_3__3 (que_out_19__3__3), .q_3__2 (
            que_out_19__3__2), .q_3__1 (que_out_19__3__1), .q_3__0 (
            que_out_19__3__0), .q_4__15 (que_out_19__4__15), .q_4__14 (
            que_out_19__4__14), .q_4__13 (que_out_19__4__13), .q_4__12 (
            que_out_19__4__12), .q_4__11 (que_out_19__4__11), .q_4__10 (
            que_out_19__4__10), .q_4__9 (que_out_19__4__9), .q_4__8 (
            que_out_19__4__8), .q_4__7 (que_out_19__4__7), .q_4__6 (
            que_out_19__4__6), .q_4__5 (que_out_19__4__5), .q_4__4 (
            que_out_19__4__4), .q_4__3 (que_out_19__4__3), .q_4__2 (
            que_out_19__4__2), .q_4__1 (que_out_19__4__1), .q_4__0 (
            que_out_19__4__0), .clk (nx10728), .load (sel_que_19), .reset (
            nx10704)) ;
    Queue_5 gen_queues_20_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_20__0__15), .q_0__14 (
            que_out_20__0__14), .q_0__13 (que_out_20__0__13), .q_0__12 (
            que_out_20__0__12), .q_0__11 (que_out_20__0__11), .q_0__10 (
            que_out_20__0__10), .q_0__9 (que_out_20__0__9), .q_0__8 (
            que_out_20__0__8), .q_0__7 (que_out_20__0__7), .q_0__6 (
            que_out_20__0__6), .q_0__5 (que_out_20__0__5), .q_0__4 (
            que_out_20__0__4), .q_0__3 (que_out_20__0__3), .q_0__2 (
            que_out_20__0__2), .q_0__1 (que_out_20__0__1), .q_0__0 (
            que_out_20__0__0), .q_1__15 (que_out_20__1__15), .q_1__14 (
            que_out_20__1__14), .q_1__13 (que_out_20__1__13), .q_1__12 (
            que_out_20__1__12), .q_1__11 (que_out_20__1__11), .q_1__10 (
            que_out_20__1__10), .q_1__9 (que_out_20__1__9), .q_1__8 (
            que_out_20__1__8), .q_1__7 (que_out_20__1__7), .q_1__6 (
            que_out_20__1__6), .q_1__5 (que_out_20__1__5), .q_1__4 (
            que_out_20__1__4), .q_1__3 (que_out_20__1__3), .q_1__2 (
            que_out_20__1__2), .q_1__1 (que_out_20__1__1), .q_1__0 (
            que_out_20__1__0), .q_2__15 (que_out_20__2__15), .q_2__14 (
            que_out_20__2__14), .q_2__13 (que_out_20__2__13), .q_2__12 (
            que_out_20__2__12), .q_2__11 (que_out_20__2__11), .q_2__10 (
            que_out_20__2__10), .q_2__9 (que_out_20__2__9), .q_2__8 (
            que_out_20__2__8), .q_2__7 (que_out_20__2__7), .q_2__6 (
            que_out_20__2__6), .q_2__5 (que_out_20__2__5), .q_2__4 (
            que_out_20__2__4), .q_2__3 (que_out_20__2__3), .q_2__2 (
            que_out_20__2__2), .q_2__1 (que_out_20__2__1), .q_2__0 (
            que_out_20__2__0), .q_3__15 (que_out_20__3__15), .q_3__14 (
            que_out_20__3__14), .q_3__13 (que_out_20__3__13), .q_3__12 (
            que_out_20__3__12), .q_3__11 (que_out_20__3__11), .q_3__10 (
            que_out_20__3__10), .q_3__9 (que_out_20__3__9), .q_3__8 (
            que_out_20__3__8), .q_3__7 (que_out_20__3__7), .q_3__6 (
            que_out_20__3__6), .q_3__5 (que_out_20__3__5), .q_3__4 (
            que_out_20__3__4), .q_3__3 (que_out_20__3__3), .q_3__2 (
            que_out_20__3__2), .q_3__1 (que_out_20__3__1), .q_3__0 (
            que_out_20__3__0), .q_4__15 (que_out_20__4__15), .q_4__14 (
            que_out_20__4__14), .q_4__13 (que_out_20__4__13), .q_4__12 (
            que_out_20__4__12), .q_4__11 (que_out_20__4__11), .q_4__10 (
            que_out_20__4__10), .q_4__9 (que_out_20__4__9), .q_4__8 (
            que_out_20__4__8), .q_4__7 (que_out_20__4__7), .q_4__6 (
            que_out_20__4__6), .q_4__5 (que_out_20__4__5), .q_4__4 (
            que_out_20__4__4), .q_4__3 (que_out_20__4__3), .q_4__2 (
            que_out_20__4__2), .q_4__1 (que_out_20__4__1), .q_4__0 (
            que_out_20__4__0), .clk (nx10730), .load (sel_que_20), .reset (
            nx10706)) ;
    Queue_5 gen_queues_21_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_21__0__15), .q_0__14 (
            que_out_21__0__14), .q_0__13 (que_out_21__0__13), .q_0__12 (
            que_out_21__0__12), .q_0__11 (que_out_21__0__11), .q_0__10 (
            que_out_21__0__10), .q_0__9 (que_out_21__0__9), .q_0__8 (
            que_out_21__0__8), .q_0__7 (que_out_21__0__7), .q_0__6 (
            que_out_21__0__6), .q_0__5 (que_out_21__0__5), .q_0__4 (
            que_out_21__0__4), .q_0__3 (que_out_21__0__3), .q_0__2 (
            que_out_21__0__2), .q_0__1 (que_out_21__0__1), .q_0__0 (
            que_out_21__0__0), .q_1__15 (que_out_21__1__15), .q_1__14 (
            que_out_21__1__14), .q_1__13 (que_out_21__1__13), .q_1__12 (
            que_out_21__1__12), .q_1__11 (que_out_21__1__11), .q_1__10 (
            que_out_21__1__10), .q_1__9 (que_out_21__1__9), .q_1__8 (
            que_out_21__1__8), .q_1__7 (que_out_21__1__7), .q_1__6 (
            que_out_21__1__6), .q_1__5 (que_out_21__1__5), .q_1__4 (
            que_out_21__1__4), .q_1__3 (que_out_21__1__3), .q_1__2 (
            que_out_21__1__2), .q_1__1 (que_out_21__1__1), .q_1__0 (
            que_out_21__1__0), .q_2__15 (que_out_21__2__15), .q_2__14 (
            que_out_21__2__14), .q_2__13 (que_out_21__2__13), .q_2__12 (
            que_out_21__2__12), .q_2__11 (que_out_21__2__11), .q_2__10 (
            que_out_21__2__10), .q_2__9 (que_out_21__2__9), .q_2__8 (
            que_out_21__2__8), .q_2__7 (que_out_21__2__7), .q_2__6 (
            que_out_21__2__6), .q_2__5 (que_out_21__2__5), .q_2__4 (
            que_out_21__2__4), .q_2__3 (que_out_21__2__3), .q_2__2 (
            que_out_21__2__2), .q_2__1 (que_out_21__2__1), .q_2__0 (
            que_out_21__2__0), .q_3__15 (que_out_21__3__15), .q_3__14 (
            que_out_21__3__14), .q_3__13 (que_out_21__3__13), .q_3__12 (
            que_out_21__3__12), .q_3__11 (que_out_21__3__11), .q_3__10 (
            que_out_21__3__10), .q_3__9 (que_out_21__3__9), .q_3__8 (
            que_out_21__3__8), .q_3__7 (que_out_21__3__7), .q_3__6 (
            que_out_21__3__6), .q_3__5 (que_out_21__3__5), .q_3__4 (
            que_out_21__3__4), .q_3__3 (que_out_21__3__3), .q_3__2 (
            que_out_21__3__2), .q_3__1 (que_out_21__3__1), .q_3__0 (
            que_out_21__3__0), .q_4__15 (que_out_21__4__15), .q_4__14 (
            que_out_21__4__14), .q_4__13 (que_out_21__4__13), .q_4__12 (
            que_out_21__4__12), .q_4__11 (que_out_21__4__11), .q_4__10 (
            que_out_21__4__10), .q_4__9 (que_out_21__4__9), .q_4__8 (
            que_out_21__4__8), .q_4__7 (que_out_21__4__7), .q_4__6 (
            que_out_21__4__6), .q_4__5 (que_out_21__4__5), .q_4__4 (
            que_out_21__4__4), .q_4__3 (que_out_21__4__3), .q_4__2 (
            que_out_21__4__2), .q_4__1 (que_out_21__4__1), .q_4__0 (
            que_out_21__4__0), .clk (nx10732), .load (sel_que_21), .reset (
            nx10708)) ;
    Queue_5 gen_queues_22_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_22__0__15), .q_0__14 (
            que_out_22__0__14), .q_0__13 (que_out_22__0__13), .q_0__12 (
            que_out_22__0__12), .q_0__11 (que_out_22__0__11), .q_0__10 (
            que_out_22__0__10), .q_0__9 (que_out_22__0__9), .q_0__8 (
            que_out_22__0__8), .q_0__7 (que_out_22__0__7), .q_0__6 (
            que_out_22__0__6), .q_0__5 (que_out_22__0__5), .q_0__4 (
            que_out_22__0__4), .q_0__3 (que_out_22__0__3), .q_0__2 (
            que_out_22__0__2), .q_0__1 (que_out_22__0__1), .q_0__0 (
            que_out_22__0__0), .q_1__15 (que_out_22__1__15), .q_1__14 (
            que_out_22__1__14), .q_1__13 (que_out_22__1__13), .q_1__12 (
            que_out_22__1__12), .q_1__11 (que_out_22__1__11), .q_1__10 (
            que_out_22__1__10), .q_1__9 (que_out_22__1__9), .q_1__8 (
            que_out_22__1__8), .q_1__7 (que_out_22__1__7), .q_1__6 (
            que_out_22__1__6), .q_1__5 (que_out_22__1__5), .q_1__4 (
            que_out_22__1__4), .q_1__3 (que_out_22__1__3), .q_1__2 (
            que_out_22__1__2), .q_1__1 (que_out_22__1__1), .q_1__0 (
            que_out_22__1__0), .q_2__15 (que_out_22__2__15), .q_2__14 (
            que_out_22__2__14), .q_2__13 (que_out_22__2__13), .q_2__12 (
            que_out_22__2__12), .q_2__11 (que_out_22__2__11), .q_2__10 (
            que_out_22__2__10), .q_2__9 (que_out_22__2__9), .q_2__8 (
            que_out_22__2__8), .q_2__7 (que_out_22__2__7), .q_2__6 (
            que_out_22__2__6), .q_2__5 (que_out_22__2__5), .q_2__4 (
            que_out_22__2__4), .q_2__3 (que_out_22__2__3), .q_2__2 (
            que_out_22__2__2), .q_2__1 (que_out_22__2__1), .q_2__0 (
            que_out_22__2__0), .q_3__15 (que_out_22__3__15), .q_3__14 (
            que_out_22__3__14), .q_3__13 (que_out_22__3__13), .q_3__12 (
            que_out_22__3__12), .q_3__11 (que_out_22__3__11), .q_3__10 (
            que_out_22__3__10), .q_3__9 (que_out_22__3__9), .q_3__8 (
            que_out_22__3__8), .q_3__7 (que_out_22__3__7), .q_3__6 (
            que_out_22__3__6), .q_3__5 (que_out_22__3__5), .q_3__4 (
            que_out_22__3__4), .q_3__3 (que_out_22__3__3), .q_3__2 (
            que_out_22__3__2), .q_3__1 (que_out_22__3__1), .q_3__0 (
            que_out_22__3__0), .q_4__15 (que_out_22__4__15), .q_4__14 (
            que_out_22__4__14), .q_4__13 (que_out_22__4__13), .q_4__12 (
            que_out_22__4__12), .q_4__11 (que_out_22__4__11), .q_4__10 (
            que_out_22__4__10), .q_4__9 (que_out_22__4__9), .q_4__8 (
            que_out_22__4__8), .q_4__7 (que_out_22__4__7), .q_4__6 (
            que_out_22__4__6), .q_4__5 (que_out_22__4__5), .q_4__4 (
            que_out_22__4__4), .q_4__3 (que_out_22__4__3), .q_4__2 (
            que_out_22__4__2), .q_4__1 (que_out_22__4__1), .q_4__0 (
            que_out_22__4__0), .clk (nx10732), .load (sel_que_22), .reset (
            nx10708)) ;
    Queue_5 gen_queues_23_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_23__0__15), .q_0__14 (
            que_out_23__0__14), .q_0__13 (que_out_23__0__13), .q_0__12 (
            que_out_23__0__12), .q_0__11 (que_out_23__0__11), .q_0__10 (
            que_out_23__0__10), .q_0__9 (que_out_23__0__9), .q_0__8 (
            que_out_23__0__8), .q_0__7 (que_out_23__0__7), .q_0__6 (
            que_out_23__0__6), .q_0__5 (que_out_23__0__5), .q_0__4 (
            que_out_23__0__4), .q_0__3 (que_out_23__0__3), .q_0__2 (
            que_out_23__0__2), .q_0__1 (que_out_23__0__1), .q_0__0 (
            que_out_23__0__0), .q_1__15 (que_out_23__1__15), .q_1__14 (
            que_out_23__1__14), .q_1__13 (que_out_23__1__13), .q_1__12 (
            que_out_23__1__12), .q_1__11 (que_out_23__1__11), .q_1__10 (
            que_out_23__1__10), .q_1__9 (que_out_23__1__9), .q_1__8 (
            que_out_23__1__8), .q_1__7 (que_out_23__1__7), .q_1__6 (
            que_out_23__1__6), .q_1__5 (que_out_23__1__5), .q_1__4 (
            que_out_23__1__4), .q_1__3 (que_out_23__1__3), .q_1__2 (
            que_out_23__1__2), .q_1__1 (que_out_23__1__1), .q_1__0 (
            que_out_23__1__0), .q_2__15 (que_out_23__2__15), .q_2__14 (
            que_out_23__2__14), .q_2__13 (que_out_23__2__13), .q_2__12 (
            que_out_23__2__12), .q_2__11 (que_out_23__2__11), .q_2__10 (
            que_out_23__2__10), .q_2__9 (que_out_23__2__9), .q_2__8 (
            que_out_23__2__8), .q_2__7 (que_out_23__2__7), .q_2__6 (
            que_out_23__2__6), .q_2__5 (que_out_23__2__5), .q_2__4 (
            que_out_23__2__4), .q_2__3 (que_out_23__2__3), .q_2__2 (
            que_out_23__2__2), .q_2__1 (que_out_23__2__1), .q_2__0 (
            que_out_23__2__0), .q_3__15 (que_out_23__3__15), .q_3__14 (
            que_out_23__3__14), .q_3__13 (que_out_23__3__13), .q_3__12 (
            que_out_23__3__12), .q_3__11 (que_out_23__3__11), .q_3__10 (
            que_out_23__3__10), .q_3__9 (que_out_23__3__9), .q_3__8 (
            que_out_23__3__8), .q_3__7 (que_out_23__3__7), .q_3__6 (
            que_out_23__3__6), .q_3__5 (que_out_23__3__5), .q_3__4 (
            que_out_23__3__4), .q_3__3 (que_out_23__3__3), .q_3__2 (
            que_out_23__3__2), .q_3__1 (que_out_23__3__1), .q_3__0 (
            que_out_23__3__0), .q_4__15 (que_out_23__4__15), .q_4__14 (
            que_out_23__4__14), .q_4__13 (que_out_23__4__13), .q_4__12 (
            que_out_23__4__12), .q_4__11 (que_out_23__4__11), .q_4__10 (
            que_out_23__4__10), .q_4__9 (que_out_23__4__9), .q_4__8 (
            que_out_23__4__8), .q_4__7 (que_out_23__4__7), .q_4__6 (
            que_out_23__4__6), .q_4__5 (que_out_23__4__5), .q_4__4 (
            que_out_23__4__4), .q_4__3 (que_out_23__4__3), .q_4__2 (
            que_out_23__4__2), .q_4__1 (que_out_23__4__1), .q_4__0 (
            que_out_23__4__0), .clk (nx10732), .load (sel_que_23), .reset (
            nx10708)) ;
    Queue_5 gen_queues_24_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_24__0__15), .q_0__14 (
            que_out_24__0__14), .q_0__13 (que_out_24__0__13), .q_0__12 (
            que_out_24__0__12), .q_0__11 (que_out_24__0__11), .q_0__10 (
            que_out_24__0__10), .q_0__9 (que_out_24__0__9), .q_0__8 (
            que_out_24__0__8), .q_0__7 (que_out_24__0__7), .q_0__6 (
            que_out_24__0__6), .q_0__5 (que_out_24__0__5), .q_0__4 (
            que_out_24__0__4), .q_0__3 (que_out_24__0__3), .q_0__2 (
            que_out_24__0__2), .q_0__1 (que_out_24__0__1), .q_0__0 (
            que_out_24__0__0), .q_1__15 (que_out_24__1__15), .q_1__14 (
            que_out_24__1__14), .q_1__13 (que_out_24__1__13), .q_1__12 (
            que_out_24__1__12), .q_1__11 (que_out_24__1__11), .q_1__10 (
            que_out_24__1__10), .q_1__9 (que_out_24__1__9), .q_1__8 (
            que_out_24__1__8), .q_1__7 (que_out_24__1__7), .q_1__6 (
            que_out_24__1__6), .q_1__5 (que_out_24__1__5), .q_1__4 (
            que_out_24__1__4), .q_1__3 (que_out_24__1__3), .q_1__2 (
            que_out_24__1__2), .q_1__1 (que_out_24__1__1), .q_1__0 (
            que_out_24__1__0), .q_2__15 (que_out_24__2__15), .q_2__14 (
            que_out_24__2__14), .q_2__13 (que_out_24__2__13), .q_2__12 (
            que_out_24__2__12), .q_2__11 (que_out_24__2__11), .q_2__10 (
            que_out_24__2__10), .q_2__9 (que_out_24__2__9), .q_2__8 (
            que_out_24__2__8), .q_2__7 (que_out_24__2__7), .q_2__6 (
            que_out_24__2__6), .q_2__5 (que_out_24__2__5), .q_2__4 (
            que_out_24__2__4), .q_2__3 (que_out_24__2__3), .q_2__2 (
            que_out_24__2__2), .q_2__1 (que_out_24__2__1), .q_2__0 (
            que_out_24__2__0), .q_3__15 (que_out_24__3__15), .q_3__14 (
            que_out_24__3__14), .q_3__13 (que_out_24__3__13), .q_3__12 (
            que_out_24__3__12), .q_3__11 (que_out_24__3__11), .q_3__10 (
            que_out_24__3__10), .q_3__9 (que_out_24__3__9), .q_3__8 (
            que_out_24__3__8), .q_3__7 (que_out_24__3__7), .q_3__6 (
            que_out_24__3__6), .q_3__5 (que_out_24__3__5), .q_3__4 (
            que_out_24__3__4), .q_3__3 (que_out_24__3__3), .q_3__2 (
            que_out_24__3__2), .q_3__1 (que_out_24__3__1), .q_3__0 (
            que_out_24__3__0), .q_4__15 (que_out_24__4__15), .q_4__14 (
            que_out_24__4__14), .q_4__13 (que_out_24__4__13), .q_4__12 (
            que_out_24__4__12), .q_4__11 (que_out_24__4__11), .q_4__10 (
            que_out_24__4__10), .q_4__9 (que_out_24__4__9), .q_4__8 (
            que_out_24__4__8), .q_4__7 (que_out_24__4__7), .q_4__6 (
            que_out_24__4__6), .q_4__5 (que_out_24__4__5), .q_4__4 (
            que_out_24__4__4), .q_4__3 (que_out_24__4__3), .q_4__2 (
            que_out_24__4__2), .q_4__1 (que_out_24__4__1), .q_4__0 (
            que_out_24__4__0), .clk (nx10734), .load (sel_que_24), .reset (
            nx10710)) ;
    Queue_5 gen_queues_25_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_25__0__15), .q_0__14 (
            que_out_25__0__14), .q_0__13 (que_out_25__0__13), .q_0__12 (
            que_out_25__0__12), .q_0__11 (que_out_25__0__11), .q_0__10 (
            que_out_25__0__10), .q_0__9 (que_out_25__0__9), .q_0__8 (
            que_out_25__0__8), .q_0__7 (que_out_25__0__7), .q_0__6 (
            que_out_25__0__6), .q_0__5 (que_out_25__0__5), .q_0__4 (
            que_out_25__0__4), .q_0__3 (que_out_25__0__3), .q_0__2 (
            que_out_25__0__2), .q_0__1 (que_out_25__0__1), .q_0__0 (
            que_out_25__0__0), .q_1__15 (que_out_25__1__15), .q_1__14 (
            que_out_25__1__14), .q_1__13 (que_out_25__1__13), .q_1__12 (
            que_out_25__1__12), .q_1__11 (que_out_25__1__11), .q_1__10 (
            que_out_25__1__10), .q_1__9 (que_out_25__1__9), .q_1__8 (
            que_out_25__1__8), .q_1__7 (que_out_25__1__7), .q_1__6 (
            que_out_25__1__6), .q_1__5 (que_out_25__1__5), .q_1__4 (
            que_out_25__1__4), .q_1__3 (que_out_25__1__3), .q_1__2 (
            que_out_25__1__2), .q_1__1 (que_out_25__1__1), .q_1__0 (
            que_out_25__1__0), .q_2__15 (que_out_25__2__15), .q_2__14 (
            que_out_25__2__14), .q_2__13 (que_out_25__2__13), .q_2__12 (
            que_out_25__2__12), .q_2__11 (que_out_25__2__11), .q_2__10 (
            que_out_25__2__10), .q_2__9 (que_out_25__2__9), .q_2__8 (
            que_out_25__2__8), .q_2__7 (que_out_25__2__7), .q_2__6 (
            que_out_25__2__6), .q_2__5 (que_out_25__2__5), .q_2__4 (
            que_out_25__2__4), .q_2__3 (que_out_25__2__3), .q_2__2 (
            que_out_25__2__2), .q_2__1 (que_out_25__2__1), .q_2__0 (
            que_out_25__2__0), .q_3__15 (que_out_25__3__15), .q_3__14 (
            que_out_25__3__14), .q_3__13 (que_out_25__3__13), .q_3__12 (
            que_out_25__3__12), .q_3__11 (que_out_25__3__11), .q_3__10 (
            que_out_25__3__10), .q_3__9 (que_out_25__3__9), .q_3__8 (
            que_out_25__3__8), .q_3__7 (que_out_25__3__7), .q_3__6 (
            que_out_25__3__6), .q_3__5 (que_out_25__3__5), .q_3__4 (
            que_out_25__3__4), .q_3__3 (que_out_25__3__3), .q_3__2 (
            que_out_25__3__2), .q_3__1 (que_out_25__3__1), .q_3__0 (
            que_out_25__3__0), .q_4__15 (que_out_25__4__15), .q_4__14 (
            que_out_25__4__14), .q_4__13 (que_out_25__4__13), .q_4__12 (
            que_out_25__4__12), .q_4__11 (que_out_25__4__11), .q_4__10 (
            que_out_25__4__10), .q_4__9 (que_out_25__4__9), .q_4__8 (
            que_out_25__4__8), .q_4__7 (que_out_25__4__7), .q_4__6 (
            que_out_25__4__6), .q_4__5 (que_out_25__4__5), .q_4__4 (
            que_out_25__4__4), .q_4__3 (que_out_25__4__3), .q_4__2 (
            que_out_25__4__2), .q_4__1 (que_out_25__4__1), .q_4__0 (
            que_out_25__4__0), .clk (nx10734), .load (sel_que_25), .reset (
            nx10710)) ;
    Queue_5 gen_queues_26_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_26__0__15), .q_0__14 (
            que_out_26__0__14), .q_0__13 (que_out_26__0__13), .q_0__12 (
            que_out_26__0__12), .q_0__11 (que_out_26__0__11), .q_0__10 (
            que_out_26__0__10), .q_0__9 (que_out_26__0__9), .q_0__8 (
            que_out_26__0__8), .q_0__7 (que_out_26__0__7), .q_0__6 (
            que_out_26__0__6), .q_0__5 (que_out_26__0__5), .q_0__4 (
            que_out_26__0__4), .q_0__3 (que_out_26__0__3), .q_0__2 (
            que_out_26__0__2), .q_0__1 (que_out_26__0__1), .q_0__0 (
            que_out_26__0__0), .q_1__15 (que_out_26__1__15), .q_1__14 (
            que_out_26__1__14), .q_1__13 (que_out_26__1__13), .q_1__12 (
            que_out_26__1__12), .q_1__11 (que_out_26__1__11), .q_1__10 (
            que_out_26__1__10), .q_1__9 (que_out_26__1__9), .q_1__8 (
            que_out_26__1__8), .q_1__7 (que_out_26__1__7), .q_1__6 (
            que_out_26__1__6), .q_1__5 (que_out_26__1__5), .q_1__4 (
            que_out_26__1__4), .q_1__3 (que_out_26__1__3), .q_1__2 (
            que_out_26__1__2), .q_1__1 (que_out_26__1__1), .q_1__0 (
            que_out_26__1__0), .q_2__15 (que_out_26__2__15), .q_2__14 (
            que_out_26__2__14), .q_2__13 (que_out_26__2__13), .q_2__12 (
            que_out_26__2__12), .q_2__11 (que_out_26__2__11), .q_2__10 (
            que_out_26__2__10), .q_2__9 (que_out_26__2__9), .q_2__8 (
            que_out_26__2__8), .q_2__7 (que_out_26__2__7), .q_2__6 (
            que_out_26__2__6), .q_2__5 (que_out_26__2__5), .q_2__4 (
            que_out_26__2__4), .q_2__3 (que_out_26__2__3), .q_2__2 (
            que_out_26__2__2), .q_2__1 (que_out_26__2__1), .q_2__0 (
            que_out_26__2__0), .q_3__15 (que_out_26__3__15), .q_3__14 (
            que_out_26__3__14), .q_3__13 (que_out_26__3__13), .q_3__12 (
            que_out_26__3__12), .q_3__11 (que_out_26__3__11), .q_3__10 (
            que_out_26__3__10), .q_3__9 (que_out_26__3__9), .q_3__8 (
            que_out_26__3__8), .q_3__7 (que_out_26__3__7), .q_3__6 (
            que_out_26__3__6), .q_3__5 (que_out_26__3__5), .q_3__4 (
            que_out_26__3__4), .q_3__3 (que_out_26__3__3), .q_3__2 (
            que_out_26__3__2), .q_3__1 (que_out_26__3__1), .q_3__0 (
            que_out_26__3__0), .q_4__15 (que_out_26__4__15), .q_4__14 (
            que_out_26__4__14), .q_4__13 (que_out_26__4__13), .q_4__12 (
            que_out_26__4__12), .q_4__11 (que_out_26__4__11), .q_4__10 (
            que_out_26__4__10), .q_4__9 (que_out_26__4__9), .q_4__8 (
            que_out_26__4__8), .q_4__7 (que_out_26__4__7), .q_4__6 (
            que_out_26__4__6), .q_4__5 (que_out_26__4__5), .q_4__4 (
            que_out_26__4__4), .q_4__3 (que_out_26__4__3), .q_4__2 (
            que_out_26__4__2), .q_4__1 (que_out_26__4__1), .q_4__0 (
            que_out_26__4__0), .clk (nx10734), .load (sel_que_26), .reset (
            nx10710)) ;
    Queue_5 gen_queues_27_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_27__0__15), .q_0__14 (
            que_out_27__0__14), .q_0__13 (que_out_27__0__13), .q_0__12 (
            que_out_27__0__12), .q_0__11 (que_out_27__0__11), .q_0__10 (
            que_out_27__0__10), .q_0__9 (que_out_27__0__9), .q_0__8 (
            que_out_27__0__8), .q_0__7 (que_out_27__0__7), .q_0__6 (
            que_out_27__0__6), .q_0__5 (que_out_27__0__5), .q_0__4 (
            que_out_27__0__4), .q_0__3 (que_out_27__0__3), .q_0__2 (
            que_out_27__0__2), .q_0__1 (que_out_27__0__1), .q_0__0 (
            que_out_27__0__0), .q_1__15 (que_out_27__1__15), .q_1__14 (
            que_out_27__1__14), .q_1__13 (que_out_27__1__13), .q_1__12 (
            que_out_27__1__12), .q_1__11 (que_out_27__1__11), .q_1__10 (
            que_out_27__1__10), .q_1__9 (que_out_27__1__9), .q_1__8 (
            que_out_27__1__8), .q_1__7 (que_out_27__1__7), .q_1__6 (
            que_out_27__1__6), .q_1__5 (que_out_27__1__5), .q_1__4 (
            que_out_27__1__4), .q_1__3 (que_out_27__1__3), .q_1__2 (
            que_out_27__1__2), .q_1__1 (que_out_27__1__1), .q_1__0 (
            que_out_27__1__0), .q_2__15 (que_out_27__2__15), .q_2__14 (
            que_out_27__2__14), .q_2__13 (que_out_27__2__13), .q_2__12 (
            que_out_27__2__12), .q_2__11 (que_out_27__2__11), .q_2__10 (
            que_out_27__2__10), .q_2__9 (que_out_27__2__9), .q_2__8 (
            que_out_27__2__8), .q_2__7 (que_out_27__2__7), .q_2__6 (
            que_out_27__2__6), .q_2__5 (que_out_27__2__5), .q_2__4 (
            que_out_27__2__4), .q_2__3 (que_out_27__2__3), .q_2__2 (
            que_out_27__2__2), .q_2__1 (que_out_27__2__1), .q_2__0 (
            que_out_27__2__0), .q_3__15 (que_out_27__3__15), .q_3__14 (
            que_out_27__3__14), .q_3__13 (que_out_27__3__13), .q_3__12 (
            que_out_27__3__12), .q_3__11 (que_out_27__3__11), .q_3__10 (
            que_out_27__3__10), .q_3__9 (que_out_27__3__9), .q_3__8 (
            que_out_27__3__8), .q_3__7 (que_out_27__3__7), .q_3__6 (
            que_out_27__3__6), .q_3__5 (que_out_27__3__5), .q_3__4 (
            que_out_27__3__4), .q_3__3 (que_out_27__3__3), .q_3__2 (
            que_out_27__3__2), .q_3__1 (que_out_27__3__1), .q_3__0 (
            que_out_27__3__0), .q_4__15 (que_out_27__4__15), .q_4__14 (
            que_out_27__4__14), .q_4__13 (que_out_27__4__13), .q_4__12 (
            que_out_27__4__12), .q_4__11 (que_out_27__4__11), .q_4__10 (
            que_out_27__4__10), .q_4__9 (que_out_27__4__9), .q_4__8 (
            que_out_27__4__8), .q_4__7 (que_out_27__4__7), .q_4__6 (
            que_out_27__4__6), .q_4__5 (que_out_27__4__5), .q_4__4 (
            que_out_27__4__4), .q_4__3 (que_out_27__4__3), .q_4__2 (
            que_out_27__4__2), .q_4__1 (que_out_27__4__1), .q_4__0 (
            que_out_27__4__0), .clk (nx10736), .load (sel_que_27), .reset (
            nx10712)) ;
    nand03 ix6830 (.Y (nx6829), .A0 (nx8938), .A1 (nx6833), .A2 (nx6835)) ;
    nor02ii ix8939 (.Y (nx8938), .A0 (cache_in_sel[4]), .A1 (decoder_enable)) ;
    inv01 ix6834 (.Y (nx6833), .A (cache_in_sel[1])) ;
    inv01 ix6836 (.Y (nx6835), .A (cache_in_sel[0])) ;
    nand03 ix6840 (.Y (nx6839), .A0 (nx8938), .A1 (nx6833), .A2 (nx10508)) ;
    nand03 ix6844 (.Y (nx6843), .A0 (nx8938), .A1 (nx10506), .A2 (nx6835)) ;
    nand03 ix6848 (.Y (nx6847), .A0 (nx8938), .A1 (nx10506), .A2 (nx10508)) ;
    nor02_2x ix9023 (.Y (sel_que_12), .A0 (nx6875), .A1 (nx6829)) ;
    nand02 ix6876 (.Y (nx6875), .A0 (cache_in_sel[3]), .A1 (cache_in_sel[2])) ;
    nor02_2x ix9025 (.Y (sel_que_13), .A0 (nx6875), .A1 (nx6839)) ;
    nor02_2x ix9027 (.Y (sel_que_14), .A0 (nx6843), .A1 (nx6875)) ;
    nor02_2x ix9029 (.Y (sel_que_15), .A0 (nx6875), .A1 (nx6847)) ;
    and02 ix9043 (.Y (sel_que_16), .A0 (nx6885), .A1 (nx9038)) ;
    nor02_2x ix6886 (.Y (nx6885), .A0 (cache_in_sel[2]), .A1 (cache_in_sel[3])
             ) ;
    nor03_2x ix9039 (.Y (nx9038), .A0 (nx6889), .A1 (nx10506), .A2 (nx10508)) ;
    nand02 ix6890 (.Y (nx6889), .A0 (cache_in_sel[4]), .A1 (decoder_enable)) ;
    nand04 ix6894 (.Y (nx6893), .A0 (cache_in_sel[4]), .A1 (decoder_enable), .A2 (
           nx6833), .A3 (nx10508)) ;
    nand04 ix6898 (.Y (nx6897), .A0 (cache_in_sel[4]), .A1 (decoder_enable), .A2 (
           nx10506), .A3 (nx6835)) ;
    nand04 ix6902 (.Y (nx6901), .A0 (cache_in_sel[4]), .A1 (decoder_enable), .A2 (
           nx10506), .A3 (nx10508)) ;
    and02 ix9075 (.Y (sel_que_20), .A0 (nx6905), .A1 (nx9038)) ;
    and02 ix9091 (.Y (sel_que_24), .A0 (nx6915), .A1 (nx9038)) ;
    or04 ix243 (.Y (out_column_4__0), .A0 (nx238), .A1 (nx188), .A2 (nx130), .A3 (
         nx82)) ;
    nand03 ix239 (.Y (nx238), .A0 (nx6927), .A1 (nx6951), .A2 (nx6967)) ;
    aoi222 ix6928 (.Y (nx6927), .A0 (que_out_10__4__0), .A1 (nx10298), .B0 (
           que_out_6__4__0), .B1 (nx10350), .C0 (que_out_9__4__0), .C1 (nx10324)
           ) ;
    nand02_2x ix6932 (.Y (nx6931), .A0 (cache_out_sel[3]), .A1 (nx6933)) ;
    inv01 ix6934 (.Y (nx6933), .A (cache_out_sel[0])) ;
    inv01 ix6938 (.Y (nx6937), .A (cache_out_sel[4])) ;
    inv02 ix6940 (.Y (nx6939), .A (cache_out_sel[2])) ;
    nand03 ix6946 (.Y (nx6945), .A0 (nx10502), .A1 (nx6937), .A2 (nx10498)) ;
    nor04 ix227 (.Y (nx226), .A0 (nx6949), .A1 (nx10502), .A2 (nx10494), .A3 (
          nx10498)) ;
    nand02_2x ix6950 (.Y (nx6949), .A0 (cache_out_sel[3]), .A1 (cache_out_sel[0]
              )) ;
    aoi22 ix6952 (.Y (nx6951), .A0 (que_out_5__4__0), .A1 (nx10246), .B0 (
          que_out_18__4__0), .B1 (nx10272)) ;
    nand02 ix6956 (.Y (nx6955), .A0 (nx6957), .A1 (cache_out_sel[0])) ;
    inv01 ix6958 (.Y (nx6957), .A (cache_out_sel[3])) ;
    inv01 ix6962 (.Y (nx6961), .A (cache_out_sel[1])) ;
    nor03_2x ix215 (.Y (nx214), .A0 (nx6965), .A1 (nx10498), .A2 (nx6943)) ;
    nand02_2x ix6966 (.Y (nx6965), .A0 (nx10494), .A1 (nx10504)) ;
    aoi22 ix6968 (.Y (nx6967), .A0 (que_out_17__4__0), .A1 (nx10220), .B0 (
          que_out_20__4__0), .B1 (nx10194)) ;
    nor03_2x ix201 (.Y (nx200), .A0 (nx6971), .A1 (nx10498), .A2 (nx10374)) ;
    nand02_2x ix6972 (.Y (nx6971), .A0 (nx10496), .A1 (nx6961)) ;
    nor03_2x ix193 (.Y (nx192), .A0 (nx6971), .A1 (nx6939), .A2 (nx6943)) ;
    nand03 ix189 (.Y (nx188), .A0 (nx6977), .A1 (nx6985), .A2 (nx6991)) ;
    aoi222 ix6978 (.Y (nx6977), .A0 (que_out_19__4__0), .A1 (nx10168), .B0 (
           que_out_21__4__0), .B1 (nx10142), .C0 (que_out_8__4__0), .C1 (nx10116
           )) ;
    nor03_2x ix181 (.Y (nx180), .A0 (nx6965), .A1 (nx10498), .A2 (nx10374)) ;
    nor03_2x ix173 (.Y (nx172), .A0 (nx6971), .A1 (nx6939), .A2 (nx10374)) ;
    nor04 ix167 (.Y (nx166), .A0 (nx6931), .A1 (nx10502), .A2 (nx10494), .A3 (
          nx10498)) ;
    aoi22 ix6986 (.Y (nx6985), .A0 (que_out_25__4__0), .A1 (nx10064), .B0 (
          que_out_16__4__0), .B1 (nx10090)) ;
    nor02_2x ix151 (.Y (nx150), .A0 (nx6949), .A1 (nx6971)) ;
    nor03_2x ix159 (.Y (nx158), .A0 (nx6971), .A1 (nx10498), .A2 (nx6943)) ;
    aoi22 ix6992 (.Y (nx6991), .A0 (que_out_24__4__0), .A1 (nx10038), .B0 (
          que_out_22__4__0), .B1 (nx10012)) ;
    nor02_2x ix145 (.Y (nx144), .A0 (nx6971), .A1 (nx6931)) ;
    nor03_2x ix137 (.Y (nx136), .A0 (nx6965), .A1 (nx6939), .A2 (nx6943)) ;
    nand03 ix131 (.Y (nx130), .A0 (nx6999), .A1 (nx7007), .A2 (nx7017)) ;
    aoi222 ix7000 (.Y (nx6999), .A0 (que_out_15__4__0), .A1 (nx9960), .B0 (
           que_out_3__4__0), .B1 (nx9986), .C0 (que_out_23__4__0), .C1 (nx9934)
           ) ;
    nor02_2x ix119 (.Y (nx118), .A0 (nx6949), .A1 (nx6945)) ;
    nor03_2x ix115 (.Y (nx114), .A0 (nx6965), .A1 (nx6939), .A2 (nx10374)) ;
    aoi22 ix7008 (.Y (nx7007), .A0 (que_out_27__4__0), .A1 (nx9908), .B0 (
          que_out_4__4__0), .B1 (nx9882)) ;
    nor02_2x ix105 (.Y (nx104), .A0 (nx6949), .A1 (nx6965)) ;
    and02 ix101 (.Y (nx100), .A0 (nx88), .A1 (nx28)) ;
    nor02_2x ix89 (.Y (nx88), .A0 (cache_out_sel[3]), .A1 (cache_out_sel[0])) ;
    nor03_2x ix29 (.Y (nx28), .A0 (nx10502), .A1 (nx10494), .A2 (nx6939)) ;
    aoi22 ix7018 (.Y (nx7017), .A0 (que_out_0__4__0), .A1 (nx9830), .B0 (
          que_out_2__4__0), .B1 (nx9856)) ;
    and02 ix91 (.Y (nx90), .A0 (nx88), .A1 (nx12)) ;
    nor03_2x ix13 (.Y (nx12), .A0 (nx10504), .A1 (nx10494), .A2 (nx10500)) ;
    and02 ix95 (.Y (nx94), .A0 (nx88), .A1 (nx62)) ;
    nor03_2x ix63 (.Y (nx62), .A0 (nx6961), .A1 (nx10494), .A2 (nx10500)) ;
    nand03 ix83 (.Y (nx82), .A0 (nx7029), .A1 (nx7037), .A2 (nx7043)) ;
    aoi222 ix7030 (.Y (nx7029), .A0 (que_out_26__4__0), .A1 (nx9804), .B0 (
           que_out_14__4__0), .B1 (nx9778), .C0 (que_out_11__4__0), .C1 (nx9752)
           ) ;
    nor02_2x ix75 (.Y (nx74), .A0 (nx6965), .A1 (nx6931)) ;
    nor02_2x ix69 (.Y (nx68), .A0 (nx6931), .A1 (nx6945)) ;
    aoi22 ix7038 (.Y (nx7037), .A0 (que_out_13__4__0), .A1 (nx9726), .B0 (
          que_out_7__4__0), .B1 (nx9700)) ;
    nor02_2x ix43 (.Y (nx42), .A0 (nx10374), .A1 (nx6945)) ;
    aoi22 ix7044 (.Y (nx7043), .A0 (que_out_12__4__0), .A1 (nx9674), .B0 (
          que_out_1__4__0), .B1 (nx9648)) ;
    nor04 ix15 (.Y (nx14), .A0 (nx10376), .A1 (nx10504), .A2 (nx10494), .A3 (
          nx10500)) ;
    or04 ix353 (.Y (out_column_4__1), .A0 (nx348), .A1 (nx322), .A2 (nx294), .A3 (
         nx268)) ;
    nand03 ix349 (.Y (nx348), .A0 (nx7053), .A1 (nx7055), .A2 (nx7057)) ;
    aoi222 ix7054 (.Y (nx7053), .A0 (que_out_10__4__1), .A1 (nx10298), .B0 (
           que_out_6__4__1), .B1 (nx10350), .C0 (que_out_9__4__1), .C1 (nx10324)
           ) ;
    aoi22 ix7056 (.Y (nx7055), .A0 (que_out_5__4__1), .A1 (nx10246), .B0 (
          que_out_18__4__1), .B1 (nx10272)) ;
    aoi22 ix7058 (.Y (nx7057), .A0 (que_out_17__4__1), .A1 (nx10220), .B0 (
          que_out_20__4__1), .B1 (nx10194)) ;
    nand03 ix323 (.Y (nx322), .A0 (nx7061), .A1 (nx7063), .A2 (nx7065)) ;
    aoi222 ix7062 (.Y (nx7061), .A0 (que_out_19__4__1), .A1 (nx10168), .B0 (
           que_out_21__4__1), .B1 (nx10142), .C0 (que_out_8__4__1), .C1 (nx10116
           )) ;
    aoi22 ix7064 (.Y (nx7063), .A0 (que_out_25__4__1), .A1 (nx10064), .B0 (
          que_out_16__4__1), .B1 (nx10090)) ;
    aoi22 ix7066 (.Y (nx7065), .A0 (que_out_24__4__1), .A1 (nx10038), .B0 (
          que_out_22__4__1), .B1 (nx10012)) ;
    nand03 ix295 (.Y (nx294), .A0 (nx7069), .A1 (nx7071), .A2 (nx7073)) ;
    aoi222 ix7070 (.Y (nx7069), .A0 (que_out_15__4__1), .A1 (nx9960), .B0 (
           que_out_3__4__1), .B1 (nx9986), .C0 (que_out_23__4__1), .C1 (nx9934)
           ) ;
    aoi22 ix7072 (.Y (nx7071), .A0 (que_out_27__4__1), .A1 (nx9908), .B0 (
          que_out_4__4__1), .B1 (nx9882)) ;
    aoi22 ix7074 (.Y (nx7073), .A0 (que_out_0__4__1), .A1 (nx9830), .B0 (
          que_out_2__4__1), .B1 (nx9856)) ;
    nand03 ix269 (.Y (nx268), .A0 (nx7077), .A1 (nx7079), .A2 (nx7081)) ;
    aoi222 ix7078 (.Y (nx7077), .A0 (que_out_26__4__1), .A1 (nx9804), .B0 (
           que_out_14__4__1), .B1 (nx9778), .C0 (que_out_11__4__1), .C1 (nx9752)
           ) ;
    aoi22 ix7080 (.Y (nx7079), .A0 (que_out_13__4__1), .A1 (nx9726), .B0 (
          que_out_7__4__1), .B1 (nx9700)) ;
    aoi22 ix7082 (.Y (nx7081), .A0 (que_out_12__4__1), .A1 (nx9674), .B0 (
          que_out_1__4__1), .B1 (nx9648)) ;
    or04 ix463 (.Y (out_column_4__2), .A0 (nx458), .A1 (nx432), .A2 (nx404), .A3 (
         nx378)) ;
    nand03 ix459 (.Y (nx458), .A0 (nx7087), .A1 (nx7089), .A2 (nx7091)) ;
    aoi222 ix7088 (.Y (nx7087), .A0 (que_out_10__4__2), .A1 (nx10298), .B0 (
           que_out_6__4__2), .B1 (nx10350), .C0 (que_out_9__4__2), .C1 (nx10324)
           ) ;
    aoi22 ix7090 (.Y (nx7089), .A0 (que_out_5__4__2), .A1 (nx10246), .B0 (
          que_out_18__4__2), .B1 (nx10272)) ;
    aoi22 ix7092 (.Y (nx7091), .A0 (que_out_17__4__2), .A1 (nx10220), .B0 (
          que_out_20__4__2), .B1 (nx10194)) ;
    nand03 ix433 (.Y (nx432), .A0 (nx7095), .A1 (nx7097), .A2 (nx7099)) ;
    aoi222 ix7096 (.Y (nx7095), .A0 (que_out_19__4__2), .A1 (nx10168), .B0 (
           que_out_21__4__2), .B1 (nx10142), .C0 (que_out_8__4__2), .C1 (nx10116
           )) ;
    aoi22 ix7098 (.Y (nx7097), .A0 (que_out_25__4__2), .A1 (nx10064), .B0 (
          que_out_16__4__2), .B1 (nx10090)) ;
    aoi22 ix7100 (.Y (nx7099), .A0 (que_out_24__4__2), .A1 (nx10038), .B0 (
          que_out_22__4__2), .B1 (nx10012)) ;
    nand03 ix405 (.Y (nx404), .A0 (nx7103), .A1 (nx7105), .A2 (nx7107)) ;
    aoi222 ix7104 (.Y (nx7103), .A0 (que_out_15__4__2), .A1 (nx9960), .B0 (
           que_out_3__4__2), .B1 (nx9986), .C0 (que_out_23__4__2), .C1 (nx9934)
           ) ;
    aoi22 ix7106 (.Y (nx7105), .A0 (que_out_27__4__2), .A1 (nx9908), .B0 (
          que_out_4__4__2), .B1 (nx9882)) ;
    aoi22 ix7108 (.Y (nx7107), .A0 (que_out_0__4__2), .A1 (nx9830), .B0 (
          que_out_2__4__2), .B1 (nx9856)) ;
    nand03 ix379 (.Y (nx378), .A0 (nx7111), .A1 (nx7113), .A2 (nx7115)) ;
    aoi222 ix7112 (.Y (nx7111), .A0 (que_out_26__4__2), .A1 (nx9804), .B0 (
           que_out_14__4__2), .B1 (nx9778), .C0 (que_out_11__4__2), .C1 (nx9752)
           ) ;
    aoi22 ix7114 (.Y (nx7113), .A0 (que_out_13__4__2), .A1 (nx9726), .B0 (
          que_out_7__4__2), .B1 (nx9700)) ;
    aoi22 ix7116 (.Y (nx7115), .A0 (que_out_12__4__2), .A1 (nx9674), .B0 (
          que_out_1__4__2), .B1 (nx9648)) ;
    or04 ix573 (.Y (out_column_4__3), .A0 (nx568), .A1 (nx542), .A2 (nx514), .A3 (
         nx488)) ;
    nand03 ix569 (.Y (nx568), .A0 (nx7121), .A1 (nx7123), .A2 (nx7125)) ;
    aoi222 ix7122 (.Y (nx7121), .A0 (que_out_10__4__3), .A1 (nx10298), .B0 (
           que_out_6__4__3), .B1 (nx10350), .C0 (que_out_9__4__3), .C1 (nx10324)
           ) ;
    aoi22 ix7124 (.Y (nx7123), .A0 (que_out_5__4__3), .A1 (nx10246), .B0 (
          que_out_18__4__3), .B1 (nx10272)) ;
    aoi22 ix7126 (.Y (nx7125), .A0 (que_out_17__4__3), .A1 (nx10220), .B0 (
          que_out_20__4__3), .B1 (nx10194)) ;
    nand03 ix543 (.Y (nx542), .A0 (nx7129), .A1 (nx7131), .A2 (nx7133)) ;
    aoi222 ix7130 (.Y (nx7129), .A0 (que_out_19__4__3), .A1 (nx10168), .B0 (
           que_out_21__4__3), .B1 (nx10142), .C0 (que_out_8__4__3), .C1 (nx10116
           )) ;
    aoi22 ix7132 (.Y (nx7131), .A0 (que_out_25__4__3), .A1 (nx10064), .B0 (
          que_out_16__4__3), .B1 (nx10090)) ;
    aoi22 ix7134 (.Y (nx7133), .A0 (que_out_24__4__3), .A1 (nx10038), .B0 (
          que_out_22__4__3), .B1 (nx10012)) ;
    nand03 ix515 (.Y (nx514), .A0 (nx7137), .A1 (nx7139), .A2 (nx7141)) ;
    aoi222 ix7138 (.Y (nx7137), .A0 (que_out_15__4__3), .A1 (nx9960), .B0 (
           que_out_3__4__3), .B1 (nx9986), .C0 (que_out_23__4__3), .C1 (nx9934)
           ) ;
    aoi22 ix7140 (.Y (nx7139), .A0 (que_out_27__4__3), .A1 (nx9908), .B0 (
          que_out_4__4__3), .B1 (nx9882)) ;
    aoi22 ix7142 (.Y (nx7141), .A0 (que_out_0__4__3), .A1 (nx9830), .B0 (
          que_out_2__4__3), .B1 (nx9856)) ;
    nand03 ix489 (.Y (nx488), .A0 (nx7145), .A1 (nx7147), .A2 (nx7149)) ;
    aoi222 ix7146 (.Y (nx7145), .A0 (que_out_26__4__3), .A1 (nx9804), .B0 (
           que_out_14__4__3), .B1 (nx9778), .C0 (que_out_11__4__3), .C1 (nx9752)
           ) ;
    aoi22 ix7148 (.Y (nx7147), .A0 (que_out_13__4__3), .A1 (nx9726), .B0 (
          que_out_7__4__3), .B1 (nx9700)) ;
    aoi22 ix7150 (.Y (nx7149), .A0 (que_out_12__4__3), .A1 (nx9674), .B0 (
          que_out_1__4__3), .B1 (nx9648)) ;
    or04 ix683 (.Y (out_column_4__4), .A0 (nx678), .A1 (nx652), .A2 (nx624), .A3 (
         nx598)) ;
    nand03 ix679 (.Y (nx678), .A0 (nx7155), .A1 (nx7157), .A2 (nx7159)) ;
    aoi222 ix7156 (.Y (nx7155), .A0 (que_out_10__4__4), .A1 (nx10298), .B0 (
           que_out_6__4__4), .B1 (nx10350), .C0 (que_out_9__4__4), .C1 (nx10324)
           ) ;
    aoi22 ix7158 (.Y (nx7157), .A0 (que_out_5__4__4), .A1 (nx10246), .B0 (
          que_out_18__4__4), .B1 (nx10272)) ;
    aoi22 ix7160 (.Y (nx7159), .A0 (que_out_17__4__4), .A1 (nx10220), .B0 (
          que_out_20__4__4), .B1 (nx10194)) ;
    nand03 ix653 (.Y (nx652), .A0 (nx7163), .A1 (nx7165), .A2 (nx7167)) ;
    aoi222 ix7164 (.Y (nx7163), .A0 (que_out_19__4__4), .A1 (nx10168), .B0 (
           que_out_21__4__4), .B1 (nx10142), .C0 (que_out_8__4__4), .C1 (nx10116
           )) ;
    aoi22 ix7166 (.Y (nx7165), .A0 (que_out_25__4__4), .A1 (nx10064), .B0 (
          que_out_16__4__4), .B1 (nx10090)) ;
    aoi22 ix7168 (.Y (nx7167), .A0 (que_out_24__4__4), .A1 (nx10038), .B0 (
          que_out_22__4__4), .B1 (nx10012)) ;
    nand03 ix625 (.Y (nx624), .A0 (nx7171), .A1 (nx7173), .A2 (nx7175)) ;
    aoi222 ix7172 (.Y (nx7171), .A0 (que_out_15__4__4), .A1 (nx9960), .B0 (
           que_out_3__4__4), .B1 (nx9986), .C0 (que_out_23__4__4), .C1 (nx9934)
           ) ;
    aoi22 ix7174 (.Y (nx7173), .A0 (que_out_27__4__4), .A1 (nx9908), .B0 (
          que_out_4__4__4), .B1 (nx9882)) ;
    aoi22 ix7176 (.Y (nx7175), .A0 (que_out_0__4__4), .A1 (nx9830), .B0 (
          que_out_2__4__4), .B1 (nx9856)) ;
    nand03 ix599 (.Y (nx598), .A0 (nx7179), .A1 (nx7181), .A2 (nx7183)) ;
    aoi222 ix7180 (.Y (nx7179), .A0 (que_out_26__4__4), .A1 (nx9804), .B0 (
           que_out_14__4__4), .B1 (nx9778), .C0 (que_out_11__4__4), .C1 (nx9752)
           ) ;
    aoi22 ix7182 (.Y (nx7181), .A0 (que_out_13__4__4), .A1 (nx9726), .B0 (
          que_out_7__4__4), .B1 (nx9700)) ;
    aoi22 ix7184 (.Y (nx7183), .A0 (que_out_12__4__4), .A1 (nx9674), .B0 (
          que_out_1__4__4), .B1 (nx9648)) ;
    or04 ix793 (.Y (out_column_4__5), .A0 (nx788), .A1 (nx762), .A2 (nx734), .A3 (
         nx708)) ;
    nand03 ix789 (.Y (nx788), .A0 (nx7189), .A1 (nx7191), .A2 (nx7193)) ;
    aoi222 ix7190 (.Y (nx7189), .A0 (que_out_10__4__5), .A1 (nx10298), .B0 (
           que_out_6__4__5), .B1 (nx10350), .C0 (que_out_9__4__5), .C1 (nx10324)
           ) ;
    aoi22 ix7192 (.Y (nx7191), .A0 (que_out_5__4__5), .A1 (nx10246), .B0 (
          que_out_18__4__5), .B1 (nx10272)) ;
    aoi22 ix7194 (.Y (nx7193), .A0 (que_out_17__4__5), .A1 (nx10220), .B0 (
          que_out_20__4__5), .B1 (nx10194)) ;
    nand03 ix763 (.Y (nx762), .A0 (nx7197), .A1 (nx7199), .A2 (nx7201)) ;
    aoi222 ix7198 (.Y (nx7197), .A0 (que_out_19__4__5), .A1 (nx10168), .B0 (
           que_out_21__4__5), .B1 (nx10142), .C0 (que_out_8__4__5), .C1 (nx10116
           )) ;
    aoi22 ix7200 (.Y (nx7199), .A0 (que_out_25__4__5), .A1 (nx10064), .B0 (
          que_out_16__4__5), .B1 (nx10090)) ;
    aoi22 ix7202 (.Y (nx7201), .A0 (que_out_24__4__5), .A1 (nx10038), .B0 (
          que_out_22__4__5), .B1 (nx10012)) ;
    nand03 ix735 (.Y (nx734), .A0 (nx7205), .A1 (nx7207), .A2 (nx7209)) ;
    aoi222 ix7206 (.Y (nx7205), .A0 (que_out_15__4__5), .A1 (nx9960), .B0 (
           que_out_3__4__5), .B1 (nx9986), .C0 (que_out_23__4__5), .C1 (nx9934)
           ) ;
    aoi22 ix7208 (.Y (nx7207), .A0 (que_out_27__4__5), .A1 (nx9908), .B0 (
          que_out_4__4__5), .B1 (nx9882)) ;
    aoi22 ix7210 (.Y (nx7209), .A0 (que_out_0__4__5), .A1 (nx9830), .B0 (
          que_out_2__4__5), .B1 (nx9856)) ;
    nand03 ix709 (.Y (nx708), .A0 (nx7213), .A1 (nx7215), .A2 (nx7217)) ;
    aoi222 ix7214 (.Y (nx7213), .A0 (que_out_26__4__5), .A1 (nx9804), .B0 (
           que_out_14__4__5), .B1 (nx9778), .C0 (que_out_11__4__5), .C1 (nx9752)
           ) ;
    aoi22 ix7216 (.Y (nx7215), .A0 (que_out_13__4__5), .A1 (nx9726), .B0 (
          que_out_7__4__5), .B1 (nx9700)) ;
    aoi22 ix7218 (.Y (nx7217), .A0 (que_out_12__4__5), .A1 (nx9674), .B0 (
          que_out_1__4__5), .B1 (nx9648)) ;
    or04 ix903 (.Y (out_column_4__6), .A0 (nx898), .A1 (nx872), .A2 (nx844), .A3 (
         nx818)) ;
    nand03 ix899 (.Y (nx898), .A0 (nx7223), .A1 (nx7225), .A2 (nx7227)) ;
    aoi222 ix7224 (.Y (nx7223), .A0 (que_out_10__4__6), .A1 (nx10298), .B0 (
           que_out_6__4__6), .B1 (nx10350), .C0 (que_out_9__4__6), .C1 (nx10324)
           ) ;
    aoi22 ix7226 (.Y (nx7225), .A0 (que_out_5__4__6), .A1 (nx10246), .B0 (
          que_out_18__4__6), .B1 (nx10272)) ;
    aoi22 ix7228 (.Y (nx7227), .A0 (que_out_17__4__6), .A1 (nx10220), .B0 (
          que_out_20__4__6), .B1 (nx10194)) ;
    nand03 ix873 (.Y (nx872), .A0 (nx7231), .A1 (nx7233), .A2 (nx7235)) ;
    aoi222 ix7232 (.Y (nx7231), .A0 (que_out_19__4__6), .A1 (nx10168), .B0 (
           que_out_21__4__6), .B1 (nx10142), .C0 (que_out_8__4__6), .C1 (nx10116
           )) ;
    aoi22 ix7234 (.Y (nx7233), .A0 (que_out_25__4__6), .A1 (nx10064), .B0 (
          que_out_16__4__6), .B1 (nx10090)) ;
    aoi22 ix7236 (.Y (nx7235), .A0 (que_out_24__4__6), .A1 (nx10038), .B0 (
          que_out_22__4__6), .B1 (nx10012)) ;
    nand03 ix845 (.Y (nx844), .A0 (nx7239), .A1 (nx7241), .A2 (nx7243)) ;
    aoi222 ix7240 (.Y (nx7239), .A0 (que_out_15__4__6), .A1 (nx9960), .B0 (
           que_out_3__4__6), .B1 (nx9986), .C0 (que_out_23__4__6), .C1 (nx9934)
           ) ;
    aoi22 ix7242 (.Y (nx7241), .A0 (que_out_27__4__6), .A1 (nx9908), .B0 (
          que_out_4__4__6), .B1 (nx9882)) ;
    aoi22 ix7244 (.Y (nx7243), .A0 (que_out_0__4__6), .A1 (nx9830), .B0 (
          que_out_2__4__6), .B1 (nx9856)) ;
    nand03 ix819 (.Y (nx818), .A0 (nx7247), .A1 (nx7249), .A2 (nx7251)) ;
    aoi222 ix7248 (.Y (nx7247), .A0 (que_out_26__4__6), .A1 (nx9804), .B0 (
           que_out_14__4__6), .B1 (nx9778), .C0 (que_out_11__4__6), .C1 (nx9752)
           ) ;
    aoi22 ix7250 (.Y (nx7249), .A0 (que_out_13__4__6), .A1 (nx9726), .B0 (
          que_out_7__4__6), .B1 (nx9700)) ;
    aoi22 ix7252 (.Y (nx7251), .A0 (que_out_12__4__6), .A1 (nx9674), .B0 (
          que_out_1__4__6), .B1 (nx9648)) ;
    or04 ix1013 (.Y (out_column_4__7), .A0 (nx1008), .A1 (nx982), .A2 (nx954), .A3 (
         nx928)) ;
    nand03 ix1009 (.Y (nx1008), .A0 (nx7257), .A1 (nx7259), .A2 (nx7261)) ;
    aoi222 ix7258 (.Y (nx7257), .A0 (que_out_10__4__7), .A1 (nx10300), .B0 (
           que_out_6__4__7), .B1 (nx10352), .C0 (que_out_9__4__7), .C1 (nx10326)
           ) ;
    aoi22 ix7260 (.Y (nx7259), .A0 (que_out_5__4__7), .A1 (nx10248), .B0 (
          que_out_18__4__7), .B1 (nx10274)) ;
    aoi22 ix7262 (.Y (nx7261), .A0 (que_out_17__4__7), .A1 (nx10222), .B0 (
          que_out_20__4__7), .B1 (nx10196)) ;
    nand03 ix983 (.Y (nx982), .A0 (nx7265), .A1 (nx7267), .A2 (nx7269)) ;
    aoi222 ix7266 (.Y (nx7265), .A0 (que_out_19__4__7), .A1 (nx10170), .B0 (
           que_out_21__4__7), .B1 (nx10144), .C0 (que_out_8__4__7), .C1 (nx10118
           )) ;
    aoi22 ix7268 (.Y (nx7267), .A0 (que_out_25__4__7), .A1 (nx10066), .B0 (
          que_out_16__4__7), .B1 (nx10092)) ;
    aoi22 ix7270 (.Y (nx7269), .A0 (que_out_24__4__7), .A1 (nx10040), .B0 (
          que_out_22__4__7), .B1 (nx10014)) ;
    nand03 ix955 (.Y (nx954), .A0 (nx7273), .A1 (nx7275), .A2 (nx7277)) ;
    aoi222 ix7274 (.Y (nx7273), .A0 (que_out_15__4__7), .A1 (nx9962), .B0 (
           que_out_3__4__7), .B1 (nx9988), .C0 (que_out_23__4__7), .C1 (nx9936)
           ) ;
    aoi22 ix7276 (.Y (nx7275), .A0 (que_out_27__4__7), .A1 (nx9910), .B0 (
          que_out_4__4__7), .B1 (nx9884)) ;
    aoi22 ix7278 (.Y (nx7277), .A0 (que_out_0__4__7), .A1 (nx9832), .B0 (
          que_out_2__4__7), .B1 (nx9858)) ;
    nand03 ix929 (.Y (nx928), .A0 (nx7281), .A1 (nx7283), .A2 (nx7285)) ;
    aoi222 ix7282 (.Y (nx7281), .A0 (que_out_26__4__7), .A1 (nx9806), .B0 (
           que_out_14__4__7), .B1 (nx9780), .C0 (que_out_11__4__7), .C1 (nx9754)
           ) ;
    aoi22 ix7284 (.Y (nx7283), .A0 (que_out_13__4__7), .A1 (nx9728), .B0 (
          que_out_7__4__7), .B1 (nx9702)) ;
    aoi22 ix7286 (.Y (nx7285), .A0 (que_out_12__4__7), .A1 (nx9676), .B0 (
          que_out_1__4__7), .B1 (nx9650)) ;
    or04 ix1123 (.Y (out_column_4__8), .A0 (nx1118), .A1 (nx1092), .A2 (nx1064)
         , .A3 (nx1038)) ;
    nand03 ix1119 (.Y (nx1118), .A0 (nx7291), .A1 (nx7293), .A2 (nx7295)) ;
    aoi222 ix7292 (.Y (nx7291), .A0 (que_out_10__4__8), .A1 (nx10300), .B0 (
           que_out_6__4__8), .B1 (nx10352), .C0 (que_out_9__4__8), .C1 (nx10326)
           ) ;
    aoi22 ix7294 (.Y (nx7293), .A0 (que_out_5__4__8), .A1 (nx10248), .B0 (
          que_out_18__4__8), .B1 (nx10274)) ;
    aoi22 ix7296 (.Y (nx7295), .A0 (que_out_17__4__8), .A1 (nx10222), .B0 (
          que_out_20__4__8), .B1 (nx10196)) ;
    nand03 ix1093 (.Y (nx1092), .A0 (nx7299), .A1 (nx7301), .A2 (nx7303)) ;
    aoi222 ix7300 (.Y (nx7299), .A0 (que_out_19__4__8), .A1 (nx10170), .B0 (
           que_out_21__4__8), .B1 (nx10144), .C0 (que_out_8__4__8), .C1 (nx10118
           )) ;
    aoi22 ix7302 (.Y (nx7301), .A0 (que_out_25__4__8), .A1 (nx10066), .B0 (
          que_out_16__4__8), .B1 (nx10092)) ;
    aoi22 ix7304 (.Y (nx7303), .A0 (que_out_24__4__8), .A1 (nx10040), .B0 (
          que_out_22__4__8), .B1 (nx10014)) ;
    nand03 ix1065 (.Y (nx1064), .A0 (nx7307), .A1 (nx7309), .A2 (nx7311)) ;
    aoi222 ix7308 (.Y (nx7307), .A0 (que_out_15__4__8), .A1 (nx9962), .B0 (
           que_out_3__4__8), .B1 (nx9988), .C0 (que_out_23__4__8), .C1 (nx9936)
           ) ;
    aoi22 ix7310 (.Y (nx7309), .A0 (que_out_27__4__8), .A1 (nx9910), .B0 (
          que_out_4__4__8), .B1 (nx9884)) ;
    aoi22 ix7312 (.Y (nx7311), .A0 (que_out_0__4__8), .A1 (nx9832), .B0 (
          que_out_2__4__8), .B1 (nx9858)) ;
    nand03 ix1039 (.Y (nx1038), .A0 (nx7315), .A1 (nx7317), .A2 (nx7319)) ;
    aoi222 ix7316 (.Y (nx7315), .A0 (que_out_26__4__8), .A1 (nx9806), .B0 (
           que_out_14__4__8), .B1 (nx9780), .C0 (que_out_11__4__8), .C1 (nx9754)
           ) ;
    aoi22 ix7318 (.Y (nx7317), .A0 (que_out_13__4__8), .A1 (nx9728), .B0 (
          que_out_7__4__8), .B1 (nx9702)) ;
    aoi22 ix7320 (.Y (nx7319), .A0 (que_out_12__4__8), .A1 (nx9676), .B0 (
          que_out_1__4__8), .B1 (nx9650)) ;
    or04 ix1233 (.Y (out_column_4__9), .A0 (nx1228), .A1 (nx1202), .A2 (nx1174)
         , .A3 (nx1148)) ;
    nand03 ix1229 (.Y (nx1228), .A0 (nx7325), .A1 (nx7327), .A2 (nx7329)) ;
    aoi222 ix7326 (.Y (nx7325), .A0 (que_out_10__4__9), .A1 (nx10300), .B0 (
           que_out_6__4__9), .B1 (nx10352), .C0 (que_out_9__4__9), .C1 (nx10326)
           ) ;
    aoi22 ix7328 (.Y (nx7327), .A0 (que_out_5__4__9), .A1 (nx10248), .B0 (
          que_out_18__4__9), .B1 (nx10274)) ;
    aoi22 ix7330 (.Y (nx7329), .A0 (que_out_17__4__9), .A1 (nx10222), .B0 (
          que_out_20__4__9), .B1 (nx10196)) ;
    nand03 ix1203 (.Y (nx1202), .A0 (nx7333), .A1 (nx7335), .A2 (nx7337)) ;
    aoi222 ix7334 (.Y (nx7333), .A0 (que_out_19__4__9), .A1 (nx10170), .B0 (
           que_out_21__4__9), .B1 (nx10144), .C0 (que_out_8__4__9), .C1 (nx10118
           )) ;
    aoi22 ix7336 (.Y (nx7335), .A0 (que_out_25__4__9), .A1 (nx10066), .B0 (
          que_out_16__4__9), .B1 (nx10092)) ;
    aoi22 ix7338 (.Y (nx7337), .A0 (que_out_24__4__9), .A1 (nx10040), .B0 (
          que_out_22__4__9), .B1 (nx10014)) ;
    nand03 ix1175 (.Y (nx1174), .A0 (nx7341), .A1 (nx7343), .A2 (nx7345)) ;
    aoi222 ix7342 (.Y (nx7341), .A0 (que_out_15__4__9), .A1 (nx9962), .B0 (
           que_out_3__4__9), .B1 (nx9988), .C0 (que_out_23__4__9), .C1 (nx9936)
           ) ;
    aoi22 ix7344 (.Y (nx7343), .A0 (que_out_27__4__9), .A1 (nx9910), .B0 (
          que_out_4__4__9), .B1 (nx9884)) ;
    aoi22 ix7346 (.Y (nx7345), .A0 (que_out_0__4__9), .A1 (nx9832), .B0 (
          que_out_2__4__9), .B1 (nx9858)) ;
    nand03 ix1149 (.Y (nx1148), .A0 (nx7349), .A1 (nx7351), .A2 (nx7353)) ;
    aoi222 ix7350 (.Y (nx7349), .A0 (que_out_26__4__9), .A1 (nx9806), .B0 (
           que_out_14__4__9), .B1 (nx9780), .C0 (que_out_11__4__9), .C1 (nx9754)
           ) ;
    aoi22 ix7352 (.Y (nx7351), .A0 (que_out_13__4__9), .A1 (nx9728), .B0 (
          que_out_7__4__9), .B1 (nx9702)) ;
    aoi22 ix7354 (.Y (nx7353), .A0 (que_out_12__4__9), .A1 (nx9676), .B0 (
          que_out_1__4__9), .B1 (nx9650)) ;
    or04 ix1343 (.Y (out_column_4__10), .A0 (nx1338), .A1 (nx1312), .A2 (nx1284)
         , .A3 (nx1258)) ;
    nand03 ix1339 (.Y (nx1338), .A0 (nx7359), .A1 (nx7361), .A2 (nx7363)) ;
    aoi222 ix7360 (.Y (nx7359), .A0 (que_out_10__4__10), .A1 (nx10300), .B0 (
           que_out_6__4__10), .B1 (nx10352), .C0 (que_out_9__4__10), .C1 (
           nx10326)) ;
    aoi22 ix7362 (.Y (nx7361), .A0 (que_out_5__4__10), .A1 (nx10248), .B0 (
          que_out_18__4__10), .B1 (nx10274)) ;
    aoi22 ix7364 (.Y (nx7363), .A0 (que_out_17__4__10), .A1 (nx10222), .B0 (
          que_out_20__4__10), .B1 (nx10196)) ;
    nand03 ix1313 (.Y (nx1312), .A0 (nx7367), .A1 (nx7369), .A2 (nx7371)) ;
    aoi222 ix7368 (.Y (nx7367), .A0 (que_out_19__4__10), .A1 (nx10170), .B0 (
           que_out_21__4__10), .B1 (nx10144), .C0 (que_out_8__4__10), .C1 (
           nx10118)) ;
    aoi22 ix7370 (.Y (nx7369), .A0 (que_out_25__4__10), .A1 (nx10066), .B0 (
          que_out_16__4__10), .B1 (nx10092)) ;
    aoi22 ix7372 (.Y (nx7371), .A0 (que_out_24__4__10), .A1 (nx10040), .B0 (
          que_out_22__4__10), .B1 (nx10014)) ;
    nand03 ix1285 (.Y (nx1284), .A0 (nx7375), .A1 (nx7377), .A2 (nx7379)) ;
    aoi222 ix7376 (.Y (nx7375), .A0 (que_out_15__4__10), .A1 (nx9962), .B0 (
           que_out_3__4__10), .B1 (nx9988), .C0 (que_out_23__4__10), .C1 (nx9936
           )) ;
    aoi22 ix7378 (.Y (nx7377), .A0 (que_out_27__4__10), .A1 (nx9910), .B0 (
          que_out_4__4__10), .B1 (nx9884)) ;
    aoi22 ix7380 (.Y (nx7379), .A0 (que_out_0__4__10), .A1 (nx9832), .B0 (
          que_out_2__4__10), .B1 (nx9858)) ;
    nand03 ix1259 (.Y (nx1258), .A0 (nx7383), .A1 (nx7385), .A2 (nx7387)) ;
    aoi222 ix7384 (.Y (nx7383), .A0 (que_out_26__4__10), .A1 (nx9806), .B0 (
           que_out_14__4__10), .B1 (nx9780), .C0 (que_out_11__4__10), .C1 (
           nx9754)) ;
    aoi22 ix7386 (.Y (nx7385), .A0 (que_out_13__4__10), .A1 (nx9728), .B0 (
          que_out_7__4__10), .B1 (nx9702)) ;
    aoi22 ix7388 (.Y (nx7387), .A0 (que_out_12__4__10), .A1 (nx9676), .B0 (
          que_out_1__4__10), .B1 (nx9650)) ;
    or04 ix1453 (.Y (out_column_4__11), .A0 (nx1448), .A1 (nx1422), .A2 (nx1394)
         , .A3 (nx1368)) ;
    nand03 ix1449 (.Y (nx1448), .A0 (nx7393), .A1 (nx7395), .A2 (nx7397)) ;
    aoi222 ix7394 (.Y (nx7393), .A0 (que_out_10__4__11), .A1 (nx10300), .B0 (
           que_out_6__4__11), .B1 (nx10352), .C0 (que_out_9__4__11), .C1 (
           nx10326)) ;
    aoi22 ix7396 (.Y (nx7395), .A0 (que_out_5__4__11), .A1 (nx10248), .B0 (
          que_out_18__4__11), .B1 (nx10274)) ;
    aoi22 ix7398 (.Y (nx7397), .A0 (que_out_17__4__11), .A1 (nx10222), .B0 (
          que_out_20__4__11), .B1 (nx10196)) ;
    nand03 ix1423 (.Y (nx1422), .A0 (nx7401), .A1 (nx7403), .A2 (nx7405)) ;
    aoi222 ix7402 (.Y (nx7401), .A0 (que_out_19__4__11), .A1 (nx10170), .B0 (
           que_out_21__4__11), .B1 (nx10144), .C0 (que_out_8__4__11), .C1 (
           nx10118)) ;
    aoi22 ix7404 (.Y (nx7403), .A0 (que_out_25__4__11), .A1 (nx10066), .B0 (
          que_out_16__4__11), .B1 (nx10092)) ;
    aoi22 ix7406 (.Y (nx7405), .A0 (que_out_24__4__11), .A1 (nx10040), .B0 (
          que_out_22__4__11), .B1 (nx10014)) ;
    nand03 ix1395 (.Y (nx1394), .A0 (nx7409), .A1 (nx7411), .A2 (nx7413)) ;
    aoi222 ix7410 (.Y (nx7409), .A0 (que_out_15__4__11), .A1 (nx9962), .B0 (
           que_out_3__4__11), .B1 (nx9988), .C0 (que_out_23__4__11), .C1 (nx9936
           )) ;
    aoi22 ix7412 (.Y (nx7411), .A0 (que_out_27__4__11), .A1 (nx9910), .B0 (
          que_out_4__4__11), .B1 (nx9884)) ;
    aoi22 ix7414 (.Y (nx7413), .A0 (que_out_0__4__11), .A1 (nx9832), .B0 (
          que_out_2__4__11), .B1 (nx9858)) ;
    nand03 ix1369 (.Y (nx1368), .A0 (nx7417), .A1 (nx7419), .A2 (nx7421)) ;
    aoi222 ix7418 (.Y (nx7417), .A0 (que_out_26__4__11), .A1 (nx9806), .B0 (
           que_out_14__4__11), .B1 (nx9780), .C0 (que_out_11__4__11), .C1 (
           nx9754)) ;
    aoi22 ix7420 (.Y (nx7419), .A0 (que_out_13__4__11), .A1 (nx9728), .B0 (
          que_out_7__4__11), .B1 (nx9702)) ;
    aoi22 ix7422 (.Y (nx7421), .A0 (que_out_12__4__11), .A1 (nx9676), .B0 (
          que_out_1__4__11), .B1 (nx9650)) ;
    or04 ix1563 (.Y (out_column_4__12), .A0 (nx1558), .A1 (nx1532), .A2 (nx1504)
         , .A3 (nx1478)) ;
    nand03 ix1559 (.Y (nx1558), .A0 (nx7427), .A1 (nx7429), .A2 (nx7431)) ;
    aoi222 ix7428 (.Y (nx7427), .A0 (que_out_10__4__12), .A1 (nx10300), .B0 (
           que_out_6__4__12), .B1 (nx10352), .C0 (que_out_9__4__12), .C1 (
           nx10326)) ;
    aoi22 ix7430 (.Y (nx7429), .A0 (que_out_5__4__12), .A1 (nx10248), .B0 (
          que_out_18__4__12), .B1 (nx10274)) ;
    aoi22 ix7432 (.Y (nx7431), .A0 (que_out_17__4__12), .A1 (nx10222), .B0 (
          que_out_20__4__12), .B1 (nx10196)) ;
    nand03 ix1533 (.Y (nx1532), .A0 (nx7435), .A1 (nx7437), .A2 (nx7439)) ;
    aoi222 ix7436 (.Y (nx7435), .A0 (que_out_19__4__12), .A1 (nx10170), .B0 (
           que_out_21__4__12), .B1 (nx10144), .C0 (que_out_8__4__12), .C1 (
           nx10118)) ;
    aoi22 ix7438 (.Y (nx7437), .A0 (que_out_25__4__12), .A1 (nx10066), .B0 (
          que_out_16__4__12), .B1 (nx10092)) ;
    aoi22 ix7440 (.Y (nx7439), .A0 (que_out_24__4__12), .A1 (nx10040), .B0 (
          que_out_22__4__12), .B1 (nx10014)) ;
    nand03 ix1505 (.Y (nx1504), .A0 (nx7443), .A1 (nx7445), .A2 (nx7447)) ;
    aoi222 ix7444 (.Y (nx7443), .A0 (que_out_15__4__12), .A1 (nx9962), .B0 (
           que_out_3__4__12), .B1 (nx9988), .C0 (que_out_23__4__12), .C1 (nx9936
           )) ;
    aoi22 ix7446 (.Y (nx7445), .A0 (que_out_27__4__12), .A1 (nx9910), .B0 (
          que_out_4__4__12), .B1 (nx9884)) ;
    aoi22 ix7448 (.Y (nx7447), .A0 (que_out_0__4__12), .A1 (nx9832), .B0 (
          que_out_2__4__12), .B1 (nx9858)) ;
    nand03 ix1479 (.Y (nx1478), .A0 (nx7451), .A1 (nx7453), .A2 (nx7455)) ;
    aoi222 ix7452 (.Y (nx7451), .A0 (que_out_26__4__12), .A1 (nx9806), .B0 (
           que_out_14__4__12), .B1 (nx9780), .C0 (que_out_11__4__12), .C1 (
           nx9754)) ;
    aoi22 ix7454 (.Y (nx7453), .A0 (que_out_13__4__12), .A1 (nx9728), .B0 (
          que_out_7__4__12), .B1 (nx9702)) ;
    aoi22 ix7456 (.Y (nx7455), .A0 (que_out_12__4__12), .A1 (nx9676), .B0 (
          que_out_1__4__12), .B1 (nx9650)) ;
    or04 ix1673 (.Y (out_column_4__13), .A0 (nx1668), .A1 (nx1642), .A2 (nx1614)
         , .A3 (nx1588)) ;
    nand03 ix1669 (.Y (nx1668), .A0 (nx7461), .A1 (nx7463), .A2 (nx7465)) ;
    aoi222 ix7462 (.Y (nx7461), .A0 (que_out_10__4__13), .A1 (nx10300), .B0 (
           que_out_6__4__13), .B1 (nx10352), .C0 (que_out_9__4__13), .C1 (
           nx10326)) ;
    aoi22 ix7464 (.Y (nx7463), .A0 (que_out_5__4__13), .A1 (nx10248), .B0 (
          que_out_18__4__13), .B1 (nx10274)) ;
    aoi22 ix7466 (.Y (nx7465), .A0 (que_out_17__4__13), .A1 (nx10222), .B0 (
          que_out_20__4__13), .B1 (nx10196)) ;
    nand03 ix1643 (.Y (nx1642), .A0 (nx7469), .A1 (nx7471), .A2 (nx7473)) ;
    aoi222 ix7470 (.Y (nx7469), .A0 (que_out_19__4__13), .A1 (nx10170), .B0 (
           que_out_21__4__13), .B1 (nx10144), .C0 (que_out_8__4__13), .C1 (
           nx10118)) ;
    aoi22 ix7472 (.Y (nx7471), .A0 (que_out_25__4__13), .A1 (nx10066), .B0 (
          que_out_16__4__13), .B1 (nx10092)) ;
    aoi22 ix7474 (.Y (nx7473), .A0 (que_out_24__4__13), .A1 (nx10040), .B0 (
          que_out_22__4__13), .B1 (nx10014)) ;
    nand03 ix1615 (.Y (nx1614), .A0 (nx7477), .A1 (nx7479), .A2 (nx7481)) ;
    aoi222 ix7478 (.Y (nx7477), .A0 (que_out_15__4__13), .A1 (nx9962), .B0 (
           que_out_3__4__13), .B1 (nx9988), .C0 (que_out_23__4__13), .C1 (nx9936
           )) ;
    aoi22 ix7480 (.Y (nx7479), .A0 (que_out_27__4__13), .A1 (nx9910), .B0 (
          que_out_4__4__13), .B1 (nx9884)) ;
    aoi22 ix7482 (.Y (nx7481), .A0 (que_out_0__4__13), .A1 (nx9832), .B0 (
          que_out_2__4__13), .B1 (nx9858)) ;
    nand03 ix1589 (.Y (nx1588), .A0 (nx7485), .A1 (nx7487), .A2 (nx7489)) ;
    aoi222 ix7486 (.Y (nx7485), .A0 (que_out_26__4__13), .A1 (nx9806), .B0 (
           que_out_14__4__13), .B1 (nx9780), .C0 (que_out_11__4__13), .C1 (
           nx9754)) ;
    aoi22 ix7488 (.Y (nx7487), .A0 (que_out_13__4__13), .A1 (nx9728), .B0 (
          que_out_7__4__13), .B1 (nx9702)) ;
    aoi22 ix7490 (.Y (nx7489), .A0 (que_out_12__4__13), .A1 (nx9676), .B0 (
          que_out_1__4__13), .B1 (nx9650)) ;
    or04 ix1783 (.Y (out_column_4__14), .A0 (nx1778), .A1 (nx1752), .A2 (nx1724)
         , .A3 (nx1698)) ;
    nand03 ix1779 (.Y (nx1778), .A0 (nx7495), .A1 (nx7497), .A2 (nx7499)) ;
    aoi222 ix7496 (.Y (nx7495), .A0 (que_out_10__4__14), .A1 (nx10302), .B0 (
           que_out_6__4__14), .B1 (nx10354), .C0 (que_out_9__4__14), .C1 (
           nx10328)) ;
    aoi22 ix7498 (.Y (nx7497), .A0 (que_out_5__4__14), .A1 (nx10250), .B0 (
          que_out_18__4__14), .B1 (nx10276)) ;
    aoi22 ix7500 (.Y (nx7499), .A0 (que_out_17__4__14), .A1 (nx10224), .B0 (
          que_out_20__4__14), .B1 (nx10198)) ;
    nand03 ix1753 (.Y (nx1752), .A0 (nx7503), .A1 (nx7505), .A2 (nx7507)) ;
    aoi222 ix7504 (.Y (nx7503), .A0 (que_out_19__4__14), .A1 (nx10172), .B0 (
           que_out_21__4__14), .B1 (nx10146), .C0 (que_out_8__4__14), .C1 (
           nx10120)) ;
    aoi22 ix7506 (.Y (nx7505), .A0 (que_out_25__4__14), .A1 (nx10068), .B0 (
          que_out_16__4__14), .B1 (nx10094)) ;
    aoi22 ix7508 (.Y (nx7507), .A0 (que_out_24__4__14), .A1 (nx10042), .B0 (
          que_out_22__4__14), .B1 (nx10016)) ;
    nand03 ix1725 (.Y (nx1724), .A0 (nx7511), .A1 (nx7513), .A2 (nx7515)) ;
    aoi222 ix7512 (.Y (nx7511), .A0 (que_out_15__4__14), .A1 (nx9964), .B0 (
           que_out_3__4__14), .B1 (nx9990), .C0 (que_out_23__4__14), .C1 (nx9938
           )) ;
    aoi22 ix7514 (.Y (nx7513), .A0 (que_out_27__4__14), .A1 (nx9912), .B0 (
          que_out_4__4__14), .B1 (nx9886)) ;
    aoi22 ix7516 (.Y (nx7515), .A0 (que_out_0__4__14), .A1 (nx9834), .B0 (
          que_out_2__4__14), .B1 (nx9860)) ;
    nand03 ix1699 (.Y (nx1698), .A0 (nx7519), .A1 (nx7521), .A2 (nx7523)) ;
    aoi222 ix7520 (.Y (nx7519), .A0 (que_out_26__4__14), .A1 (nx9808), .B0 (
           que_out_14__4__14), .B1 (nx9782), .C0 (que_out_11__4__14), .C1 (
           nx9756)) ;
    aoi22 ix7522 (.Y (nx7521), .A0 (que_out_13__4__14), .A1 (nx9730), .B0 (
          que_out_7__4__14), .B1 (nx9704)) ;
    aoi22 ix7524 (.Y (nx7523), .A0 (que_out_12__4__14), .A1 (nx9678), .B0 (
          que_out_1__4__14), .B1 (nx9652)) ;
    or04 ix1893 (.Y (out_column_4__15), .A0 (nx1888), .A1 (nx1862), .A2 (nx1834)
         , .A3 (nx1808)) ;
    nand03 ix1889 (.Y (nx1888), .A0 (nx7529), .A1 (nx7531), .A2 (nx7533)) ;
    aoi222 ix7530 (.Y (nx7529), .A0 (que_out_10__4__15), .A1 (nx10302), .B0 (
           que_out_6__4__15), .B1 (nx10354), .C0 (que_out_9__4__15), .C1 (
           nx10328)) ;
    aoi22 ix7532 (.Y (nx7531), .A0 (que_out_5__4__15), .A1 (nx10250), .B0 (
          que_out_18__4__15), .B1 (nx10276)) ;
    aoi22 ix7534 (.Y (nx7533), .A0 (que_out_17__4__15), .A1 (nx10224), .B0 (
          que_out_20__4__15), .B1 (nx10198)) ;
    nand03 ix1863 (.Y (nx1862), .A0 (nx7537), .A1 (nx7539), .A2 (nx7541)) ;
    aoi222 ix7538 (.Y (nx7537), .A0 (que_out_19__4__15), .A1 (nx10172), .B0 (
           que_out_21__4__15), .B1 (nx10146), .C0 (que_out_8__4__15), .C1 (
           nx10120)) ;
    aoi22 ix7540 (.Y (nx7539), .A0 (que_out_25__4__15), .A1 (nx10068), .B0 (
          que_out_16__4__15), .B1 (nx10094)) ;
    aoi22 ix7542 (.Y (nx7541), .A0 (que_out_24__4__15), .A1 (nx10042), .B0 (
          que_out_22__4__15), .B1 (nx10016)) ;
    nand03 ix1835 (.Y (nx1834), .A0 (nx7545), .A1 (nx7547), .A2 (nx7549)) ;
    aoi222 ix7546 (.Y (nx7545), .A0 (que_out_15__4__15), .A1 (nx9964), .B0 (
           que_out_3__4__15), .B1 (nx9990), .C0 (que_out_23__4__15), .C1 (nx9938
           )) ;
    aoi22 ix7548 (.Y (nx7547), .A0 (que_out_27__4__15), .A1 (nx9912), .B0 (
          que_out_4__4__15), .B1 (nx9886)) ;
    aoi22 ix7550 (.Y (nx7549), .A0 (que_out_0__4__15), .A1 (nx9834), .B0 (
          que_out_2__4__15), .B1 (nx9860)) ;
    nand03 ix1809 (.Y (nx1808), .A0 (nx7553), .A1 (nx7555), .A2 (nx7557)) ;
    aoi222 ix7554 (.Y (nx7553), .A0 (que_out_26__4__15), .A1 (nx9808), .B0 (
           que_out_14__4__15), .B1 (nx9782), .C0 (que_out_11__4__15), .C1 (
           nx9756)) ;
    aoi22 ix7556 (.Y (nx7555), .A0 (que_out_13__4__15), .A1 (nx9730), .B0 (
          que_out_7__4__15), .B1 (nx9704)) ;
    aoi22 ix7558 (.Y (nx7557), .A0 (que_out_12__4__15), .A1 (nx9678), .B0 (
          que_out_1__4__15), .B1 (nx9652)) ;
    or04 ix2003 (.Y (out_column_3__0), .A0 (nx1998), .A1 (nx1972), .A2 (nx1944)
         , .A3 (nx1918)) ;
    nand03 ix1999 (.Y (nx1998), .A0 (nx7563), .A1 (nx7565), .A2 (nx7567)) ;
    aoi222 ix7564 (.Y (nx7563), .A0 (que_out_10__3__0), .A1 (nx10302), .B0 (
           que_out_6__3__0), .B1 (nx10354), .C0 (que_out_9__3__0), .C1 (nx10328)
           ) ;
    aoi22 ix7566 (.Y (nx7565), .A0 (que_out_5__3__0), .A1 (nx10250), .B0 (
          que_out_18__3__0), .B1 (nx10276)) ;
    aoi22 ix7568 (.Y (nx7567), .A0 (que_out_17__3__0), .A1 (nx10224), .B0 (
          que_out_20__3__0), .B1 (nx10198)) ;
    nand03 ix1973 (.Y (nx1972), .A0 (nx7571), .A1 (nx7573), .A2 (nx7575)) ;
    aoi222 ix7572 (.Y (nx7571), .A0 (que_out_19__3__0), .A1 (nx10172), .B0 (
           que_out_21__3__0), .B1 (nx10146), .C0 (que_out_8__3__0), .C1 (nx10120
           )) ;
    aoi22 ix7574 (.Y (nx7573), .A0 (que_out_25__3__0), .A1 (nx10068), .B0 (
          que_out_16__3__0), .B1 (nx10094)) ;
    aoi22 ix7576 (.Y (nx7575), .A0 (que_out_24__3__0), .A1 (nx10042), .B0 (
          que_out_22__3__0), .B1 (nx10016)) ;
    nand03 ix1945 (.Y (nx1944), .A0 (nx7579), .A1 (nx7581), .A2 (nx7583)) ;
    aoi222 ix7580 (.Y (nx7579), .A0 (que_out_15__3__0), .A1 (nx9964), .B0 (
           que_out_3__3__0), .B1 (nx9990), .C0 (que_out_23__3__0), .C1 (nx9938)
           ) ;
    aoi22 ix7582 (.Y (nx7581), .A0 (que_out_27__3__0), .A1 (nx9912), .B0 (
          que_out_4__3__0), .B1 (nx9886)) ;
    aoi22 ix7584 (.Y (nx7583), .A0 (que_out_0__3__0), .A1 (nx9834), .B0 (
          que_out_2__3__0), .B1 (nx9860)) ;
    nand03 ix1919 (.Y (nx1918), .A0 (nx7587), .A1 (nx7589), .A2 (nx7591)) ;
    aoi222 ix7588 (.Y (nx7587), .A0 (que_out_26__3__0), .A1 (nx9808), .B0 (
           que_out_14__3__0), .B1 (nx9782), .C0 (que_out_11__3__0), .C1 (nx9756)
           ) ;
    aoi22 ix7590 (.Y (nx7589), .A0 (que_out_13__3__0), .A1 (nx9730), .B0 (
          que_out_7__3__0), .B1 (nx9704)) ;
    aoi22 ix7592 (.Y (nx7591), .A0 (que_out_12__3__0), .A1 (nx9678), .B0 (
          que_out_1__3__0), .B1 (nx9652)) ;
    or04 ix2113 (.Y (out_column_3__1), .A0 (nx2108), .A1 (nx2082), .A2 (nx2054)
         , .A3 (nx2028)) ;
    nand03 ix2109 (.Y (nx2108), .A0 (nx7597), .A1 (nx7599), .A2 (nx7601)) ;
    aoi222 ix7598 (.Y (nx7597), .A0 (que_out_10__3__1), .A1 (nx10302), .B0 (
           que_out_6__3__1), .B1 (nx10354), .C0 (que_out_9__3__1), .C1 (nx10328)
           ) ;
    aoi22 ix7600 (.Y (nx7599), .A0 (que_out_5__3__1), .A1 (nx10250), .B0 (
          que_out_18__3__1), .B1 (nx10276)) ;
    aoi22 ix7602 (.Y (nx7601), .A0 (que_out_17__3__1), .A1 (nx10224), .B0 (
          que_out_20__3__1), .B1 (nx10198)) ;
    nand03 ix2083 (.Y (nx2082), .A0 (nx7605), .A1 (nx7607), .A2 (nx7609)) ;
    aoi222 ix7606 (.Y (nx7605), .A0 (que_out_19__3__1), .A1 (nx10172), .B0 (
           que_out_21__3__1), .B1 (nx10146), .C0 (que_out_8__3__1), .C1 (nx10120
           )) ;
    aoi22 ix7608 (.Y (nx7607), .A0 (que_out_25__3__1), .A1 (nx10068), .B0 (
          que_out_16__3__1), .B1 (nx10094)) ;
    aoi22 ix7610 (.Y (nx7609), .A0 (que_out_24__3__1), .A1 (nx10042), .B0 (
          que_out_22__3__1), .B1 (nx10016)) ;
    nand03 ix2055 (.Y (nx2054), .A0 (nx7613), .A1 (nx7615), .A2 (nx7617)) ;
    aoi222 ix7614 (.Y (nx7613), .A0 (que_out_15__3__1), .A1 (nx9964), .B0 (
           que_out_3__3__1), .B1 (nx9990), .C0 (que_out_23__3__1), .C1 (nx9938)
           ) ;
    aoi22 ix7616 (.Y (nx7615), .A0 (que_out_27__3__1), .A1 (nx9912), .B0 (
          que_out_4__3__1), .B1 (nx9886)) ;
    aoi22 ix7618 (.Y (nx7617), .A0 (que_out_0__3__1), .A1 (nx9834), .B0 (
          que_out_2__3__1), .B1 (nx9860)) ;
    nand03 ix2029 (.Y (nx2028), .A0 (nx7621), .A1 (nx7623), .A2 (nx7625)) ;
    aoi222 ix7622 (.Y (nx7621), .A0 (que_out_26__3__1), .A1 (nx9808), .B0 (
           que_out_14__3__1), .B1 (nx9782), .C0 (que_out_11__3__1), .C1 (nx9756)
           ) ;
    aoi22 ix7624 (.Y (nx7623), .A0 (que_out_13__3__1), .A1 (nx9730), .B0 (
          que_out_7__3__1), .B1 (nx9704)) ;
    aoi22 ix7626 (.Y (nx7625), .A0 (que_out_12__3__1), .A1 (nx9678), .B0 (
          que_out_1__3__1), .B1 (nx9652)) ;
    or04 ix2223 (.Y (out_column_3__2), .A0 (nx2218), .A1 (nx2192), .A2 (nx2164)
         , .A3 (nx2138)) ;
    nand03 ix2219 (.Y (nx2218), .A0 (nx7631), .A1 (nx7633), .A2 (nx7635)) ;
    aoi222 ix7632 (.Y (nx7631), .A0 (que_out_10__3__2), .A1 (nx10302), .B0 (
           que_out_6__3__2), .B1 (nx10354), .C0 (que_out_9__3__2), .C1 (nx10328)
           ) ;
    aoi22 ix7634 (.Y (nx7633), .A0 (que_out_5__3__2), .A1 (nx10250), .B0 (
          que_out_18__3__2), .B1 (nx10276)) ;
    aoi22 ix7636 (.Y (nx7635), .A0 (que_out_17__3__2), .A1 (nx10224), .B0 (
          que_out_20__3__2), .B1 (nx10198)) ;
    nand03 ix2193 (.Y (nx2192), .A0 (nx7639), .A1 (nx7641), .A2 (nx7643)) ;
    aoi222 ix7640 (.Y (nx7639), .A0 (que_out_19__3__2), .A1 (nx10172), .B0 (
           que_out_21__3__2), .B1 (nx10146), .C0 (que_out_8__3__2), .C1 (nx10120
           )) ;
    aoi22 ix7642 (.Y (nx7641), .A0 (que_out_25__3__2), .A1 (nx10068), .B0 (
          que_out_16__3__2), .B1 (nx10094)) ;
    aoi22 ix7644 (.Y (nx7643), .A0 (que_out_24__3__2), .A1 (nx10042), .B0 (
          que_out_22__3__2), .B1 (nx10016)) ;
    nand03 ix2165 (.Y (nx2164), .A0 (nx7647), .A1 (nx7649), .A2 (nx7651)) ;
    aoi222 ix7648 (.Y (nx7647), .A0 (que_out_15__3__2), .A1 (nx9964), .B0 (
           que_out_3__3__2), .B1 (nx9990), .C0 (que_out_23__3__2), .C1 (nx9938)
           ) ;
    aoi22 ix7650 (.Y (nx7649), .A0 (que_out_27__3__2), .A1 (nx9912), .B0 (
          que_out_4__3__2), .B1 (nx9886)) ;
    aoi22 ix7652 (.Y (nx7651), .A0 (que_out_0__3__2), .A1 (nx9834), .B0 (
          que_out_2__3__2), .B1 (nx9860)) ;
    nand03 ix2139 (.Y (nx2138), .A0 (nx7655), .A1 (nx7657), .A2 (nx7659)) ;
    aoi222 ix7656 (.Y (nx7655), .A0 (que_out_26__3__2), .A1 (nx9808), .B0 (
           que_out_14__3__2), .B1 (nx9782), .C0 (que_out_11__3__2), .C1 (nx9756)
           ) ;
    aoi22 ix7658 (.Y (nx7657), .A0 (que_out_13__3__2), .A1 (nx9730), .B0 (
          que_out_7__3__2), .B1 (nx9704)) ;
    aoi22 ix7660 (.Y (nx7659), .A0 (que_out_12__3__2), .A1 (nx9678), .B0 (
          que_out_1__3__2), .B1 (nx9652)) ;
    or04 ix2333 (.Y (out_column_3__3), .A0 (nx2328), .A1 (nx2302), .A2 (nx2274)
         , .A3 (nx2248)) ;
    nand03 ix2329 (.Y (nx2328), .A0 (nx7665), .A1 (nx7667), .A2 (nx7669)) ;
    aoi222 ix7666 (.Y (nx7665), .A0 (que_out_10__3__3), .A1 (nx10302), .B0 (
           que_out_6__3__3), .B1 (nx10354), .C0 (que_out_9__3__3), .C1 (nx10328)
           ) ;
    aoi22 ix7668 (.Y (nx7667), .A0 (que_out_5__3__3), .A1 (nx10250), .B0 (
          que_out_18__3__3), .B1 (nx10276)) ;
    aoi22 ix7670 (.Y (nx7669), .A0 (que_out_17__3__3), .A1 (nx10224), .B0 (
          que_out_20__3__3), .B1 (nx10198)) ;
    nand03 ix2303 (.Y (nx2302), .A0 (nx7673), .A1 (nx7675), .A2 (nx7677)) ;
    aoi222 ix7674 (.Y (nx7673), .A0 (que_out_19__3__3), .A1 (nx10172), .B0 (
           que_out_21__3__3), .B1 (nx10146), .C0 (que_out_8__3__3), .C1 (nx10120
           )) ;
    aoi22 ix7676 (.Y (nx7675), .A0 (que_out_25__3__3), .A1 (nx10068), .B0 (
          que_out_16__3__3), .B1 (nx10094)) ;
    aoi22 ix7678 (.Y (nx7677), .A0 (que_out_24__3__3), .A1 (nx10042), .B0 (
          que_out_22__3__3), .B1 (nx10016)) ;
    nand03 ix2275 (.Y (nx2274), .A0 (nx7681), .A1 (nx7683), .A2 (nx7685)) ;
    aoi222 ix7682 (.Y (nx7681), .A0 (que_out_15__3__3), .A1 (nx9964), .B0 (
           que_out_3__3__3), .B1 (nx9990), .C0 (que_out_23__3__3), .C1 (nx9938)
           ) ;
    aoi22 ix7684 (.Y (nx7683), .A0 (que_out_27__3__3), .A1 (nx9912), .B0 (
          que_out_4__3__3), .B1 (nx9886)) ;
    aoi22 ix7686 (.Y (nx7685), .A0 (que_out_0__3__3), .A1 (nx9834), .B0 (
          que_out_2__3__3), .B1 (nx9860)) ;
    nand03 ix2249 (.Y (nx2248), .A0 (nx7689), .A1 (nx7691), .A2 (nx7693)) ;
    aoi222 ix7690 (.Y (nx7689), .A0 (que_out_26__3__3), .A1 (nx9808), .B0 (
           que_out_14__3__3), .B1 (nx9782), .C0 (que_out_11__3__3), .C1 (nx9756)
           ) ;
    aoi22 ix7692 (.Y (nx7691), .A0 (que_out_13__3__3), .A1 (nx9730), .B0 (
          que_out_7__3__3), .B1 (nx9704)) ;
    aoi22 ix7694 (.Y (nx7693), .A0 (que_out_12__3__3), .A1 (nx9678), .B0 (
          que_out_1__3__3), .B1 (nx9652)) ;
    or04 ix2443 (.Y (out_column_3__4), .A0 (nx2438), .A1 (nx2412), .A2 (nx2384)
         , .A3 (nx2358)) ;
    nand03 ix2439 (.Y (nx2438), .A0 (nx7699), .A1 (nx7701), .A2 (nx7703)) ;
    aoi222 ix7700 (.Y (nx7699), .A0 (que_out_10__3__4), .A1 (nx10302), .B0 (
           que_out_6__3__4), .B1 (nx10354), .C0 (que_out_9__3__4), .C1 (nx10328)
           ) ;
    aoi22 ix7702 (.Y (nx7701), .A0 (que_out_5__3__4), .A1 (nx10250), .B0 (
          que_out_18__3__4), .B1 (nx10276)) ;
    aoi22 ix7704 (.Y (nx7703), .A0 (que_out_17__3__4), .A1 (nx10224), .B0 (
          que_out_20__3__4), .B1 (nx10198)) ;
    nand03 ix2413 (.Y (nx2412), .A0 (nx7707), .A1 (nx7709), .A2 (nx7711)) ;
    aoi222 ix7708 (.Y (nx7707), .A0 (que_out_19__3__4), .A1 (nx10172), .B0 (
           que_out_21__3__4), .B1 (nx10146), .C0 (que_out_8__3__4), .C1 (nx10120
           )) ;
    aoi22 ix7710 (.Y (nx7709), .A0 (que_out_25__3__4), .A1 (nx10068), .B0 (
          que_out_16__3__4), .B1 (nx10094)) ;
    aoi22 ix7712 (.Y (nx7711), .A0 (que_out_24__3__4), .A1 (nx10042), .B0 (
          que_out_22__3__4), .B1 (nx10016)) ;
    nand03 ix2385 (.Y (nx2384), .A0 (nx7715), .A1 (nx7717), .A2 (nx7719)) ;
    aoi222 ix7716 (.Y (nx7715), .A0 (que_out_15__3__4), .A1 (nx9964), .B0 (
           que_out_3__3__4), .B1 (nx9990), .C0 (que_out_23__3__4), .C1 (nx9938)
           ) ;
    aoi22 ix7718 (.Y (nx7717), .A0 (que_out_27__3__4), .A1 (nx9912), .B0 (
          que_out_4__3__4), .B1 (nx9886)) ;
    aoi22 ix7720 (.Y (nx7719), .A0 (que_out_0__3__4), .A1 (nx9834), .B0 (
          que_out_2__3__4), .B1 (nx9860)) ;
    nand03 ix2359 (.Y (nx2358), .A0 (nx7723), .A1 (nx7725), .A2 (nx7727)) ;
    aoi222 ix7724 (.Y (nx7723), .A0 (que_out_26__3__4), .A1 (nx9808), .B0 (
           que_out_14__3__4), .B1 (nx9782), .C0 (que_out_11__3__4), .C1 (nx9756)
           ) ;
    aoi22 ix7726 (.Y (nx7725), .A0 (que_out_13__3__4), .A1 (nx9730), .B0 (
          que_out_7__3__4), .B1 (nx9704)) ;
    aoi22 ix7728 (.Y (nx7727), .A0 (que_out_12__3__4), .A1 (nx9678), .B0 (
          que_out_1__3__4), .B1 (nx9652)) ;
    or04 ix2553 (.Y (out_column_3__5), .A0 (nx2548), .A1 (nx2522), .A2 (nx2494)
         , .A3 (nx2468)) ;
    nand03 ix2549 (.Y (nx2548), .A0 (nx7733), .A1 (nx7735), .A2 (nx7737)) ;
    aoi222 ix7734 (.Y (nx7733), .A0 (que_out_10__3__5), .A1 (nx10304), .B0 (
           que_out_6__3__5), .B1 (nx10356), .C0 (que_out_9__3__5), .C1 (nx10330)
           ) ;
    aoi22 ix7736 (.Y (nx7735), .A0 (que_out_5__3__5), .A1 (nx10252), .B0 (
          que_out_18__3__5), .B1 (nx10278)) ;
    aoi22 ix7738 (.Y (nx7737), .A0 (que_out_17__3__5), .A1 (nx10226), .B0 (
          que_out_20__3__5), .B1 (nx10200)) ;
    nand03 ix2523 (.Y (nx2522), .A0 (nx7741), .A1 (nx7743), .A2 (nx7745)) ;
    aoi222 ix7742 (.Y (nx7741), .A0 (que_out_19__3__5), .A1 (nx10174), .B0 (
           que_out_21__3__5), .B1 (nx10148), .C0 (que_out_8__3__5), .C1 (nx10122
           )) ;
    aoi22 ix7744 (.Y (nx7743), .A0 (que_out_25__3__5), .A1 (nx10070), .B0 (
          que_out_16__3__5), .B1 (nx10096)) ;
    aoi22 ix7746 (.Y (nx7745), .A0 (que_out_24__3__5), .A1 (nx10044), .B0 (
          que_out_22__3__5), .B1 (nx10018)) ;
    nand03 ix2495 (.Y (nx2494), .A0 (nx7749), .A1 (nx7751), .A2 (nx7753)) ;
    aoi222 ix7750 (.Y (nx7749), .A0 (que_out_15__3__5), .A1 (nx9966), .B0 (
           que_out_3__3__5), .B1 (nx9992), .C0 (que_out_23__3__5), .C1 (nx9940)
           ) ;
    aoi22 ix7752 (.Y (nx7751), .A0 (que_out_27__3__5), .A1 (nx9914), .B0 (
          que_out_4__3__5), .B1 (nx9888)) ;
    aoi22 ix7754 (.Y (nx7753), .A0 (que_out_0__3__5), .A1 (nx9836), .B0 (
          que_out_2__3__5), .B1 (nx9862)) ;
    nand03 ix2469 (.Y (nx2468), .A0 (nx7757), .A1 (nx7759), .A2 (nx7761)) ;
    aoi222 ix7758 (.Y (nx7757), .A0 (que_out_26__3__5), .A1 (nx9810), .B0 (
           que_out_14__3__5), .B1 (nx9784), .C0 (que_out_11__3__5), .C1 (nx9758)
           ) ;
    aoi22 ix7760 (.Y (nx7759), .A0 (que_out_13__3__5), .A1 (nx9732), .B0 (
          que_out_7__3__5), .B1 (nx9706)) ;
    aoi22 ix7762 (.Y (nx7761), .A0 (que_out_12__3__5), .A1 (nx9680), .B0 (
          que_out_1__3__5), .B1 (nx9654)) ;
    or04 ix2663 (.Y (out_column_3__6), .A0 (nx2658), .A1 (nx2632), .A2 (nx2604)
         , .A3 (nx2578)) ;
    nand03 ix2659 (.Y (nx2658), .A0 (nx7767), .A1 (nx7769), .A2 (nx7771)) ;
    aoi222 ix7768 (.Y (nx7767), .A0 (que_out_10__3__6), .A1 (nx10304), .B0 (
           que_out_6__3__6), .B1 (nx10356), .C0 (que_out_9__3__6), .C1 (nx10330)
           ) ;
    aoi22 ix7770 (.Y (nx7769), .A0 (que_out_5__3__6), .A1 (nx10252), .B0 (
          que_out_18__3__6), .B1 (nx10278)) ;
    aoi22 ix7772 (.Y (nx7771), .A0 (que_out_17__3__6), .A1 (nx10226), .B0 (
          que_out_20__3__6), .B1 (nx10200)) ;
    nand03 ix2633 (.Y (nx2632), .A0 (nx7775), .A1 (nx7777), .A2 (nx7779)) ;
    aoi222 ix7776 (.Y (nx7775), .A0 (que_out_19__3__6), .A1 (nx10174), .B0 (
           que_out_21__3__6), .B1 (nx10148), .C0 (que_out_8__3__6), .C1 (nx10122
           )) ;
    aoi22 ix7778 (.Y (nx7777), .A0 (que_out_25__3__6), .A1 (nx10070), .B0 (
          que_out_16__3__6), .B1 (nx10096)) ;
    aoi22 ix7780 (.Y (nx7779), .A0 (que_out_24__3__6), .A1 (nx10044), .B0 (
          que_out_22__3__6), .B1 (nx10018)) ;
    nand03 ix2605 (.Y (nx2604), .A0 (nx7783), .A1 (nx7785), .A2 (nx7787)) ;
    aoi222 ix7784 (.Y (nx7783), .A0 (que_out_15__3__6), .A1 (nx9966), .B0 (
           que_out_3__3__6), .B1 (nx9992), .C0 (que_out_23__3__6), .C1 (nx9940)
           ) ;
    aoi22 ix7786 (.Y (nx7785), .A0 (que_out_27__3__6), .A1 (nx9914), .B0 (
          que_out_4__3__6), .B1 (nx9888)) ;
    aoi22 ix7788 (.Y (nx7787), .A0 (que_out_0__3__6), .A1 (nx9836), .B0 (
          que_out_2__3__6), .B1 (nx9862)) ;
    nand03 ix2579 (.Y (nx2578), .A0 (nx7791), .A1 (nx7793), .A2 (nx7795)) ;
    aoi222 ix7792 (.Y (nx7791), .A0 (que_out_26__3__6), .A1 (nx9810), .B0 (
           que_out_14__3__6), .B1 (nx9784), .C0 (que_out_11__3__6), .C1 (nx9758)
           ) ;
    aoi22 ix7794 (.Y (nx7793), .A0 (que_out_13__3__6), .A1 (nx9732), .B0 (
          que_out_7__3__6), .B1 (nx9706)) ;
    aoi22 ix7796 (.Y (nx7795), .A0 (que_out_12__3__6), .A1 (nx9680), .B0 (
          que_out_1__3__6), .B1 (nx9654)) ;
    or04 ix2773 (.Y (out_column_3__7), .A0 (nx2768), .A1 (nx2742), .A2 (nx2714)
         , .A3 (nx2688)) ;
    nand03 ix2769 (.Y (nx2768), .A0 (nx7801), .A1 (nx7803), .A2 (nx7805)) ;
    aoi222 ix7802 (.Y (nx7801), .A0 (que_out_10__3__7), .A1 (nx10304), .B0 (
           que_out_6__3__7), .B1 (nx10356), .C0 (que_out_9__3__7), .C1 (nx10330)
           ) ;
    aoi22 ix7804 (.Y (nx7803), .A0 (que_out_5__3__7), .A1 (nx10252), .B0 (
          que_out_18__3__7), .B1 (nx10278)) ;
    aoi22 ix7806 (.Y (nx7805), .A0 (que_out_17__3__7), .A1 (nx10226), .B0 (
          que_out_20__3__7), .B1 (nx10200)) ;
    nand03 ix2743 (.Y (nx2742), .A0 (nx7809), .A1 (nx7811), .A2 (nx7813)) ;
    aoi222 ix7810 (.Y (nx7809), .A0 (que_out_19__3__7), .A1 (nx10174), .B0 (
           que_out_21__3__7), .B1 (nx10148), .C0 (que_out_8__3__7), .C1 (nx10122
           )) ;
    aoi22 ix7812 (.Y (nx7811), .A0 (que_out_25__3__7), .A1 (nx10070), .B0 (
          que_out_16__3__7), .B1 (nx10096)) ;
    aoi22 ix7814 (.Y (nx7813), .A0 (que_out_24__3__7), .A1 (nx10044), .B0 (
          que_out_22__3__7), .B1 (nx10018)) ;
    nand03 ix2715 (.Y (nx2714), .A0 (nx7817), .A1 (nx7819), .A2 (nx7821)) ;
    aoi222 ix7818 (.Y (nx7817), .A0 (que_out_15__3__7), .A1 (nx9966), .B0 (
           que_out_3__3__7), .B1 (nx9992), .C0 (que_out_23__3__7), .C1 (nx9940)
           ) ;
    aoi22 ix7820 (.Y (nx7819), .A0 (que_out_27__3__7), .A1 (nx9914), .B0 (
          que_out_4__3__7), .B1 (nx9888)) ;
    aoi22 ix7822 (.Y (nx7821), .A0 (que_out_0__3__7), .A1 (nx9836), .B0 (
          que_out_2__3__7), .B1 (nx9862)) ;
    nand03 ix2689 (.Y (nx2688), .A0 (nx7825), .A1 (nx7827), .A2 (nx7829)) ;
    aoi222 ix7826 (.Y (nx7825), .A0 (que_out_26__3__7), .A1 (nx9810), .B0 (
           que_out_14__3__7), .B1 (nx9784), .C0 (que_out_11__3__7), .C1 (nx9758)
           ) ;
    aoi22 ix7828 (.Y (nx7827), .A0 (que_out_13__3__7), .A1 (nx9732), .B0 (
          que_out_7__3__7), .B1 (nx9706)) ;
    aoi22 ix7830 (.Y (nx7829), .A0 (que_out_12__3__7), .A1 (nx9680), .B0 (
          que_out_1__3__7), .B1 (nx9654)) ;
    or04 ix2883 (.Y (out_column_3__8), .A0 (nx2878), .A1 (nx2852), .A2 (nx2824)
         , .A3 (nx2798)) ;
    nand03 ix2879 (.Y (nx2878), .A0 (nx7835), .A1 (nx7837), .A2 (nx7839)) ;
    aoi222 ix7836 (.Y (nx7835), .A0 (que_out_10__3__8), .A1 (nx10304), .B0 (
           que_out_6__3__8), .B1 (nx10356), .C0 (que_out_9__3__8), .C1 (nx10330)
           ) ;
    aoi22 ix7838 (.Y (nx7837), .A0 (que_out_5__3__8), .A1 (nx10252), .B0 (
          que_out_18__3__8), .B1 (nx10278)) ;
    aoi22 ix7840 (.Y (nx7839), .A0 (que_out_17__3__8), .A1 (nx10226), .B0 (
          que_out_20__3__8), .B1 (nx10200)) ;
    nand03 ix2853 (.Y (nx2852), .A0 (nx7843), .A1 (nx7845), .A2 (nx7847)) ;
    aoi222 ix7844 (.Y (nx7843), .A0 (que_out_19__3__8), .A1 (nx10174), .B0 (
           que_out_21__3__8), .B1 (nx10148), .C0 (que_out_8__3__8), .C1 (nx10122
           )) ;
    aoi22 ix7846 (.Y (nx7845), .A0 (que_out_25__3__8), .A1 (nx10070), .B0 (
          que_out_16__3__8), .B1 (nx10096)) ;
    aoi22 ix7848 (.Y (nx7847), .A0 (que_out_24__3__8), .A1 (nx10044), .B0 (
          que_out_22__3__8), .B1 (nx10018)) ;
    nand03 ix2825 (.Y (nx2824), .A0 (nx7851), .A1 (nx7853), .A2 (nx7855)) ;
    aoi222 ix7852 (.Y (nx7851), .A0 (que_out_15__3__8), .A1 (nx9966), .B0 (
           que_out_3__3__8), .B1 (nx9992), .C0 (que_out_23__3__8), .C1 (nx9940)
           ) ;
    aoi22 ix7854 (.Y (nx7853), .A0 (que_out_27__3__8), .A1 (nx9914), .B0 (
          que_out_4__3__8), .B1 (nx9888)) ;
    aoi22 ix7856 (.Y (nx7855), .A0 (que_out_0__3__8), .A1 (nx9836), .B0 (
          que_out_2__3__8), .B1 (nx9862)) ;
    nand03 ix2799 (.Y (nx2798), .A0 (nx7859), .A1 (nx7861), .A2 (nx7863)) ;
    aoi222 ix7860 (.Y (nx7859), .A0 (que_out_26__3__8), .A1 (nx9810), .B0 (
           que_out_14__3__8), .B1 (nx9784), .C0 (que_out_11__3__8), .C1 (nx9758)
           ) ;
    aoi22 ix7862 (.Y (nx7861), .A0 (que_out_13__3__8), .A1 (nx9732), .B0 (
          que_out_7__3__8), .B1 (nx9706)) ;
    aoi22 ix7864 (.Y (nx7863), .A0 (que_out_12__3__8), .A1 (nx9680), .B0 (
          que_out_1__3__8), .B1 (nx9654)) ;
    or04 ix2993 (.Y (out_column_3__9), .A0 (nx2988), .A1 (nx2962), .A2 (nx2934)
         , .A3 (nx2908)) ;
    nand03 ix2989 (.Y (nx2988), .A0 (nx7869), .A1 (nx7871), .A2 (nx7873)) ;
    aoi222 ix7870 (.Y (nx7869), .A0 (que_out_10__3__9), .A1 (nx10304), .B0 (
           que_out_6__3__9), .B1 (nx10356), .C0 (que_out_9__3__9), .C1 (nx10330)
           ) ;
    aoi22 ix7872 (.Y (nx7871), .A0 (que_out_5__3__9), .A1 (nx10252), .B0 (
          que_out_18__3__9), .B1 (nx10278)) ;
    aoi22 ix7874 (.Y (nx7873), .A0 (que_out_17__3__9), .A1 (nx10226), .B0 (
          que_out_20__3__9), .B1 (nx10200)) ;
    nand03 ix2963 (.Y (nx2962), .A0 (nx7877), .A1 (nx7879), .A2 (nx7881)) ;
    aoi222 ix7878 (.Y (nx7877), .A0 (que_out_19__3__9), .A1 (nx10174), .B0 (
           que_out_21__3__9), .B1 (nx10148), .C0 (que_out_8__3__9), .C1 (nx10122
           )) ;
    aoi22 ix7880 (.Y (nx7879), .A0 (que_out_25__3__9), .A1 (nx10070), .B0 (
          que_out_16__3__9), .B1 (nx10096)) ;
    aoi22 ix7882 (.Y (nx7881), .A0 (que_out_24__3__9), .A1 (nx10044), .B0 (
          que_out_22__3__9), .B1 (nx10018)) ;
    nand03 ix2935 (.Y (nx2934), .A0 (nx7885), .A1 (nx7887), .A2 (nx7889)) ;
    aoi222 ix7886 (.Y (nx7885), .A0 (que_out_15__3__9), .A1 (nx9966), .B0 (
           que_out_3__3__9), .B1 (nx9992), .C0 (que_out_23__3__9), .C1 (nx9940)
           ) ;
    aoi22 ix7888 (.Y (nx7887), .A0 (que_out_27__3__9), .A1 (nx9914), .B0 (
          que_out_4__3__9), .B1 (nx9888)) ;
    aoi22 ix7890 (.Y (nx7889), .A0 (que_out_0__3__9), .A1 (nx9836), .B0 (
          que_out_2__3__9), .B1 (nx9862)) ;
    nand03 ix2909 (.Y (nx2908), .A0 (nx7893), .A1 (nx7895), .A2 (nx7897)) ;
    aoi222 ix7894 (.Y (nx7893), .A0 (que_out_26__3__9), .A1 (nx9810), .B0 (
           que_out_14__3__9), .B1 (nx9784), .C0 (que_out_11__3__9), .C1 (nx9758)
           ) ;
    aoi22 ix7896 (.Y (nx7895), .A0 (que_out_13__3__9), .A1 (nx9732), .B0 (
          que_out_7__3__9), .B1 (nx9706)) ;
    aoi22 ix7898 (.Y (nx7897), .A0 (que_out_12__3__9), .A1 (nx9680), .B0 (
          que_out_1__3__9), .B1 (nx9654)) ;
    or04 ix3103 (.Y (out_column_3__10), .A0 (nx3098), .A1 (nx3072), .A2 (nx3044)
         , .A3 (nx3018)) ;
    nand03 ix3099 (.Y (nx3098), .A0 (nx7903), .A1 (nx7905), .A2 (nx7907)) ;
    aoi222 ix7904 (.Y (nx7903), .A0 (que_out_10__3__10), .A1 (nx10304), .B0 (
           que_out_6__3__10), .B1 (nx10356), .C0 (que_out_9__3__10), .C1 (
           nx10330)) ;
    aoi22 ix7906 (.Y (nx7905), .A0 (que_out_5__3__10), .A1 (nx10252), .B0 (
          que_out_18__3__10), .B1 (nx10278)) ;
    aoi22 ix7908 (.Y (nx7907), .A0 (que_out_17__3__10), .A1 (nx10226), .B0 (
          que_out_20__3__10), .B1 (nx10200)) ;
    nand03 ix3073 (.Y (nx3072), .A0 (nx7911), .A1 (nx7913), .A2 (nx7915)) ;
    aoi222 ix7912 (.Y (nx7911), .A0 (que_out_19__3__10), .A1 (nx10174), .B0 (
           que_out_21__3__10), .B1 (nx10148), .C0 (que_out_8__3__10), .C1 (
           nx10122)) ;
    aoi22 ix7914 (.Y (nx7913), .A0 (que_out_25__3__10), .A1 (nx10070), .B0 (
          que_out_16__3__10), .B1 (nx10096)) ;
    aoi22 ix7916 (.Y (nx7915), .A0 (que_out_24__3__10), .A1 (nx10044), .B0 (
          que_out_22__3__10), .B1 (nx10018)) ;
    nand03 ix3045 (.Y (nx3044), .A0 (nx7919), .A1 (nx7921), .A2 (nx7923)) ;
    aoi222 ix7920 (.Y (nx7919), .A0 (que_out_15__3__10), .A1 (nx9966), .B0 (
           que_out_3__3__10), .B1 (nx9992), .C0 (que_out_23__3__10), .C1 (nx9940
           )) ;
    aoi22 ix7922 (.Y (nx7921), .A0 (que_out_27__3__10), .A1 (nx9914), .B0 (
          que_out_4__3__10), .B1 (nx9888)) ;
    aoi22 ix7924 (.Y (nx7923), .A0 (que_out_0__3__10), .A1 (nx9836), .B0 (
          que_out_2__3__10), .B1 (nx9862)) ;
    nand03 ix3019 (.Y (nx3018), .A0 (nx7927), .A1 (nx7929), .A2 (nx7931)) ;
    aoi222 ix7928 (.Y (nx7927), .A0 (que_out_26__3__10), .A1 (nx9810), .B0 (
           que_out_14__3__10), .B1 (nx9784), .C0 (que_out_11__3__10), .C1 (
           nx9758)) ;
    aoi22 ix7930 (.Y (nx7929), .A0 (que_out_13__3__10), .A1 (nx9732), .B0 (
          que_out_7__3__10), .B1 (nx9706)) ;
    aoi22 ix7932 (.Y (nx7931), .A0 (que_out_12__3__10), .A1 (nx9680), .B0 (
          que_out_1__3__10), .B1 (nx9654)) ;
    or04 ix3213 (.Y (out_column_3__11), .A0 (nx3208), .A1 (nx3182), .A2 (nx3154)
         , .A3 (nx3128)) ;
    nand03 ix3209 (.Y (nx3208), .A0 (nx7937), .A1 (nx7939), .A2 (nx7941)) ;
    aoi222 ix7938 (.Y (nx7937), .A0 (que_out_10__3__11), .A1 (nx10304), .B0 (
           que_out_6__3__11), .B1 (nx10356), .C0 (que_out_9__3__11), .C1 (
           nx10330)) ;
    aoi22 ix7940 (.Y (nx7939), .A0 (que_out_5__3__11), .A1 (nx10252), .B0 (
          que_out_18__3__11), .B1 (nx10278)) ;
    aoi22 ix7942 (.Y (nx7941), .A0 (que_out_17__3__11), .A1 (nx10226), .B0 (
          que_out_20__3__11), .B1 (nx10200)) ;
    nand03 ix3183 (.Y (nx3182), .A0 (nx7945), .A1 (nx7947), .A2 (nx7949)) ;
    aoi222 ix7946 (.Y (nx7945), .A0 (que_out_19__3__11), .A1 (nx10174), .B0 (
           que_out_21__3__11), .B1 (nx10148), .C0 (que_out_8__3__11), .C1 (
           nx10122)) ;
    aoi22 ix7948 (.Y (nx7947), .A0 (que_out_25__3__11), .A1 (nx10070), .B0 (
          que_out_16__3__11), .B1 (nx10096)) ;
    aoi22 ix7950 (.Y (nx7949), .A0 (que_out_24__3__11), .A1 (nx10044), .B0 (
          que_out_22__3__11), .B1 (nx10018)) ;
    nand03 ix3155 (.Y (nx3154), .A0 (nx7953), .A1 (nx7955), .A2 (nx7957)) ;
    aoi222 ix7954 (.Y (nx7953), .A0 (que_out_15__3__11), .A1 (nx9966), .B0 (
           que_out_3__3__11), .B1 (nx9992), .C0 (que_out_23__3__11), .C1 (nx9940
           )) ;
    aoi22 ix7956 (.Y (nx7955), .A0 (que_out_27__3__11), .A1 (nx9914), .B0 (
          que_out_4__3__11), .B1 (nx9888)) ;
    aoi22 ix7958 (.Y (nx7957), .A0 (que_out_0__3__11), .A1 (nx9836), .B0 (
          que_out_2__3__11), .B1 (nx9862)) ;
    nand03 ix3129 (.Y (nx3128), .A0 (nx7961), .A1 (nx7963), .A2 (nx7965)) ;
    aoi222 ix7962 (.Y (nx7961), .A0 (que_out_26__3__11), .A1 (nx9810), .B0 (
           que_out_14__3__11), .B1 (nx9784), .C0 (que_out_11__3__11), .C1 (
           nx9758)) ;
    aoi22 ix7964 (.Y (nx7963), .A0 (que_out_13__3__11), .A1 (nx9732), .B0 (
          que_out_7__3__11), .B1 (nx9706)) ;
    aoi22 ix7966 (.Y (nx7965), .A0 (que_out_12__3__11), .A1 (nx9680), .B0 (
          que_out_1__3__11), .B1 (nx9654)) ;
    or04 ix3323 (.Y (out_column_3__12), .A0 (nx3318), .A1 (nx3292), .A2 (nx3264)
         , .A3 (nx3238)) ;
    nand03 ix3319 (.Y (nx3318), .A0 (nx7971), .A1 (nx7973), .A2 (nx7975)) ;
    aoi222 ix7972 (.Y (nx7971), .A0 (que_out_10__3__12), .A1 (nx10306), .B0 (
           que_out_6__3__12), .B1 (nx10358), .C0 (que_out_9__3__12), .C1 (
           nx10332)) ;
    aoi22 ix7974 (.Y (nx7973), .A0 (que_out_5__3__12), .A1 (nx10254), .B0 (
          que_out_18__3__12), .B1 (nx10280)) ;
    aoi22 ix7976 (.Y (nx7975), .A0 (que_out_17__3__12), .A1 (nx10228), .B0 (
          que_out_20__3__12), .B1 (nx10202)) ;
    nand03 ix3293 (.Y (nx3292), .A0 (nx7979), .A1 (nx7981), .A2 (nx7983)) ;
    aoi222 ix7980 (.Y (nx7979), .A0 (que_out_19__3__12), .A1 (nx10176), .B0 (
           que_out_21__3__12), .B1 (nx10150), .C0 (que_out_8__3__12), .C1 (
           nx10124)) ;
    aoi22 ix7982 (.Y (nx7981), .A0 (que_out_25__3__12), .A1 (nx10072), .B0 (
          que_out_16__3__12), .B1 (nx10098)) ;
    aoi22 ix7984 (.Y (nx7983), .A0 (que_out_24__3__12), .A1 (nx10046), .B0 (
          que_out_22__3__12), .B1 (nx10020)) ;
    nand03 ix3265 (.Y (nx3264), .A0 (nx7987), .A1 (nx7989), .A2 (nx7991)) ;
    aoi222 ix7988 (.Y (nx7987), .A0 (que_out_15__3__12), .A1 (nx9968), .B0 (
           que_out_3__3__12), .B1 (nx9994), .C0 (que_out_23__3__12), .C1 (nx9942
           )) ;
    aoi22 ix7990 (.Y (nx7989), .A0 (que_out_27__3__12), .A1 (nx9916), .B0 (
          que_out_4__3__12), .B1 (nx9890)) ;
    aoi22 ix7992 (.Y (nx7991), .A0 (que_out_0__3__12), .A1 (nx9838), .B0 (
          que_out_2__3__12), .B1 (nx9864)) ;
    nand03 ix3239 (.Y (nx3238), .A0 (nx7995), .A1 (nx7997), .A2 (nx7999)) ;
    aoi222 ix7996 (.Y (nx7995), .A0 (que_out_26__3__12), .A1 (nx9812), .B0 (
           que_out_14__3__12), .B1 (nx9786), .C0 (que_out_11__3__12), .C1 (
           nx9760)) ;
    aoi22 ix7998 (.Y (nx7997), .A0 (que_out_13__3__12), .A1 (nx9734), .B0 (
          que_out_7__3__12), .B1 (nx9708)) ;
    aoi22 ix8000 (.Y (nx7999), .A0 (que_out_12__3__12), .A1 (nx9682), .B0 (
          que_out_1__3__12), .B1 (nx9656)) ;
    or04 ix3433 (.Y (out_column_3__13), .A0 (nx3428), .A1 (nx3402), .A2 (nx3374)
         , .A3 (nx3348)) ;
    nand03 ix3429 (.Y (nx3428), .A0 (nx8005), .A1 (nx8007), .A2 (nx8009)) ;
    aoi222 ix8006 (.Y (nx8005), .A0 (que_out_10__3__13), .A1 (nx10306), .B0 (
           que_out_6__3__13), .B1 (nx10358), .C0 (que_out_9__3__13), .C1 (
           nx10332)) ;
    aoi22 ix8008 (.Y (nx8007), .A0 (que_out_5__3__13), .A1 (nx10254), .B0 (
          que_out_18__3__13), .B1 (nx10280)) ;
    aoi22 ix8010 (.Y (nx8009), .A0 (que_out_17__3__13), .A1 (nx10228), .B0 (
          que_out_20__3__13), .B1 (nx10202)) ;
    nand03 ix3403 (.Y (nx3402), .A0 (nx8013), .A1 (nx8015), .A2 (nx8017)) ;
    aoi222 ix8014 (.Y (nx8013), .A0 (que_out_19__3__13), .A1 (nx10176), .B0 (
           que_out_21__3__13), .B1 (nx10150), .C0 (que_out_8__3__13), .C1 (
           nx10124)) ;
    aoi22 ix8016 (.Y (nx8015), .A0 (que_out_25__3__13), .A1 (nx10072), .B0 (
          que_out_16__3__13), .B1 (nx10098)) ;
    aoi22 ix8018 (.Y (nx8017), .A0 (que_out_24__3__13), .A1 (nx10046), .B0 (
          que_out_22__3__13), .B1 (nx10020)) ;
    nand03 ix3375 (.Y (nx3374), .A0 (nx8021), .A1 (nx8023), .A2 (nx8025)) ;
    aoi222 ix8022 (.Y (nx8021), .A0 (que_out_15__3__13), .A1 (nx9968), .B0 (
           que_out_3__3__13), .B1 (nx9994), .C0 (que_out_23__3__13), .C1 (nx9942
           )) ;
    aoi22 ix8024 (.Y (nx8023), .A0 (que_out_27__3__13), .A1 (nx9916), .B0 (
          que_out_4__3__13), .B1 (nx9890)) ;
    aoi22 ix8026 (.Y (nx8025), .A0 (que_out_0__3__13), .A1 (nx9838), .B0 (
          que_out_2__3__13), .B1 (nx9864)) ;
    nand03 ix3349 (.Y (nx3348), .A0 (nx8029), .A1 (nx8031), .A2 (nx8033)) ;
    aoi222 ix8030 (.Y (nx8029), .A0 (que_out_26__3__13), .A1 (nx9812), .B0 (
           que_out_14__3__13), .B1 (nx9786), .C0 (que_out_11__3__13), .C1 (
           nx9760)) ;
    aoi22 ix8032 (.Y (nx8031), .A0 (que_out_13__3__13), .A1 (nx9734), .B0 (
          que_out_7__3__13), .B1 (nx9708)) ;
    aoi22 ix8034 (.Y (nx8033), .A0 (que_out_12__3__13), .A1 (nx9682), .B0 (
          que_out_1__3__13), .B1 (nx9656)) ;
    or04 ix3543 (.Y (out_column_3__14), .A0 (nx3538), .A1 (nx3512), .A2 (nx3484)
         , .A3 (nx3458)) ;
    nand03 ix3539 (.Y (nx3538), .A0 (nx8039), .A1 (nx8041), .A2 (nx8043)) ;
    aoi222 ix8040 (.Y (nx8039), .A0 (que_out_10__3__14), .A1 (nx10306), .B0 (
           que_out_6__3__14), .B1 (nx10358), .C0 (que_out_9__3__14), .C1 (
           nx10332)) ;
    aoi22 ix8042 (.Y (nx8041), .A0 (que_out_5__3__14), .A1 (nx10254), .B0 (
          que_out_18__3__14), .B1 (nx10280)) ;
    aoi22 ix8044 (.Y (nx8043), .A0 (que_out_17__3__14), .A1 (nx10228), .B0 (
          que_out_20__3__14), .B1 (nx10202)) ;
    nand03 ix3513 (.Y (nx3512), .A0 (nx8047), .A1 (nx8049), .A2 (nx8051)) ;
    aoi222 ix8048 (.Y (nx8047), .A0 (que_out_19__3__14), .A1 (nx10176), .B0 (
           que_out_21__3__14), .B1 (nx10150), .C0 (que_out_8__3__14), .C1 (
           nx10124)) ;
    aoi22 ix8050 (.Y (nx8049), .A0 (que_out_25__3__14), .A1 (nx10072), .B0 (
          que_out_16__3__14), .B1 (nx10098)) ;
    aoi22 ix8052 (.Y (nx8051), .A0 (que_out_24__3__14), .A1 (nx10046), .B0 (
          que_out_22__3__14), .B1 (nx10020)) ;
    nand03 ix3485 (.Y (nx3484), .A0 (nx8055), .A1 (nx8057), .A2 (nx8059)) ;
    aoi222 ix8056 (.Y (nx8055), .A0 (que_out_15__3__14), .A1 (nx9968), .B0 (
           que_out_3__3__14), .B1 (nx9994), .C0 (que_out_23__3__14), .C1 (nx9942
           )) ;
    aoi22 ix8058 (.Y (nx8057), .A0 (que_out_27__3__14), .A1 (nx9916), .B0 (
          que_out_4__3__14), .B1 (nx9890)) ;
    aoi22 ix8060 (.Y (nx8059), .A0 (que_out_0__3__14), .A1 (nx9838), .B0 (
          que_out_2__3__14), .B1 (nx9864)) ;
    nand03 ix3459 (.Y (nx3458), .A0 (nx8063), .A1 (nx8065), .A2 (nx8067)) ;
    aoi222 ix8064 (.Y (nx8063), .A0 (que_out_26__3__14), .A1 (nx9812), .B0 (
           que_out_14__3__14), .B1 (nx9786), .C0 (que_out_11__3__14), .C1 (
           nx9760)) ;
    aoi22 ix8066 (.Y (nx8065), .A0 (que_out_13__3__14), .A1 (nx9734), .B0 (
          que_out_7__3__14), .B1 (nx9708)) ;
    aoi22 ix8068 (.Y (nx8067), .A0 (que_out_12__3__14), .A1 (nx9682), .B0 (
          que_out_1__3__14), .B1 (nx9656)) ;
    or04 ix3653 (.Y (out_column_3__15), .A0 (nx3648), .A1 (nx3622), .A2 (nx3594)
         , .A3 (nx3568)) ;
    nand03 ix3649 (.Y (nx3648), .A0 (nx8073), .A1 (nx8075), .A2 (nx8077)) ;
    aoi222 ix8074 (.Y (nx8073), .A0 (que_out_10__3__15), .A1 (nx10306), .B0 (
           que_out_6__3__15), .B1 (nx10358), .C0 (que_out_9__3__15), .C1 (
           nx10332)) ;
    aoi22 ix8076 (.Y (nx8075), .A0 (que_out_5__3__15), .A1 (nx10254), .B0 (
          que_out_18__3__15), .B1 (nx10280)) ;
    aoi22 ix8078 (.Y (nx8077), .A0 (que_out_17__3__15), .A1 (nx10228), .B0 (
          que_out_20__3__15), .B1 (nx10202)) ;
    nand03 ix3623 (.Y (nx3622), .A0 (nx8081), .A1 (nx8083), .A2 (nx8085)) ;
    aoi222 ix8082 (.Y (nx8081), .A0 (que_out_19__3__15), .A1 (nx10176), .B0 (
           que_out_21__3__15), .B1 (nx10150), .C0 (que_out_8__3__15), .C1 (
           nx10124)) ;
    aoi22 ix8084 (.Y (nx8083), .A0 (que_out_25__3__15), .A1 (nx10072), .B0 (
          que_out_16__3__15), .B1 (nx10098)) ;
    aoi22 ix8086 (.Y (nx8085), .A0 (que_out_24__3__15), .A1 (nx10046), .B0 (
          que_out_22__3__15), .B1 (nx10020)) ;
    nand03 ix3595 (.Y (nx3594), .A0 (nx8089), .A1 (nx8091), .A2 (nx8093)) ;
    aoi222 ix8090 (.Y (nx8089), .A0 (que_out_15__3__15), .A1 (nx9968), .B0 (
           que_out_3__3__15), .B1 (nx9994), .C0 (que_out_23__3__15), .C1 (nx9942
           )) ;
    aoi22 ix8092 (.Y (nx8091), .A0 (que_out_27__3__15), .A1 (nx9916), .B0 (
          que_out_4__3__15), .B1 (nx9890)) ;
    aoi22 ix8094 (.Y (nx8093), .A0 (que_out_0__3__15), .A1 (nx9838), .B0 (
          que_out_2__3__15), .B1 (nx9864)) ;
    nand03 ix3569 (.Y (nx3568), .A0 (nx8097), .A1 (nx8099), .A2 (nx8101)) ;
    aoi222 ix8098 (.Y (nx8097), .A0 (que_out_26__3__15), .A1 (nx9812), .B0 (
           que_out_14__3__15), .B1 (nx9786), .C0 (que_out_11__3__15), .C1 (
           nx9760)) ;
    aoi22 ix8100 (.Y (nx8099), .A0 (que_out_13__3__15), .A1 (nx9734), .B0 (
          que_out_7__3__15), .B1 (nx9708)) ;
    aoi22 ix8102 (.Y (nx8101), .A0 (que_out_12__3__15), .A1 (nx9682), .B0 (
          que_out_1__3__15), .B1 (nx9656)) ;
    or04 ix3763 (.Y (out_column_2__0), .A0 (nx3758), .A1 (nx3732), .A2 (nx3704)
         , .A3 (nx3678)) ;
    nand03 ix3759 (.Y (nx3758), .A0 (nx8107), .A1 (nx8109), .A2 (nx8111)) ;
    aoi222 ix8108 (.Y (nx8107), .A0 (que_out_10__2__0), .A1 (nx10306), .B0 (
           que_out_6__2__0), .B1 (nx10358), .C0 (que_out_9__2__0), .C1 (nx10332)
           ) ;
    aoi22 ix8110 (.Y (nx8109), .A0 (que_out_5__2__0), .A1 (nx10254), .B0 (
          que_out_18__2__0), .B1 (nx10280)) ;
    aoi22 ix8112 (.Y (nx8111), .A0 (que_out_17__2__0), .A1 (nx10228), .B0 (
          que_out_20__2__0), .B1 (nx10202)) ;
    nand03 ix3733 (.Y (nx3732), .A0 (nx8115), .A1 (nx8117), .A2 (nx8119)) ;
    aoi222 ix8116 (.Y (nx8115), .A0 (que_out_19__2__0), .A1 (nx10176), .B0 (
           que_out_21__2__0), .B1 (nx10150), .C0 (que_out_8__2__0), .C1 (nx10124
           )) ;
    aoi22 ix8118 (.Y (nx8117), .A0 (que_out_25__2__0), .A1 (nx10072), .B0 (
          que_out_16__2__0), .B1 (nx10098)) ;
    aoi22 ix8120 (.Y (nx8119), .A0 (que_out_24__2__0), .A1 (nx10046), .B0 (
          que_out_22__2__0), .B1 (nx10020)) ;
    nand03 ix3705 (.Y (nx3704), .A0 (nx8123), .A1 (nx8125), .A2 (nx8127)) ;
    aoi222 ix8124 (.Y (nx8123), .A0 (que_out_15__2__0), .A1 (nx9968), .B0 (
           que_out_3__2__0), .B1 (nx9994), .C0 (que_out_23__2__0), .C1 (nx9942)
           ) ;
    aoi22 ix8126 (.Y (nx8125), .A0 (que_out_27__2__0), .A1 (nx9916), .B0 (
          que_out_4__2__0), .B1 (nx9890)) ;
    aoi22 ix8128 (.Y (nx8127), .A0 (que_out_0__2__0), .A1 (nx9838), .B0 (
          que_out_2__2__0), .B1 (nx9864)) ;
    nand03 ix3679 (.Y (nx3678), .A0 (nx8131), .A1 (nx8133), .A2 (nx8135)) ;
    aoi222 ix8132 (.Y (nx8131), .A0 (que_out_26__2__0), .A1 (nx9812), .B0 (
           que_out_14__2__0), .B1 (nx9786), .C0 (que_out_11__2__0), .C1 (nx9760)
           ) ;
    aoi22 ix8134 (.Y (nx8133), .A0 (que_out_13__2__0), .A1 (nx9734), .B0 (
          que_out_7__2__0), .B1 (nx9708)) ;
    aoi22 ix8136 (.Y (nx8135), .A0 (que_out_12__2__0), .A1 (nx9682), .B0 (
          que_out_1__2__0), .B1 (nx9656)) ;
    or04 ix3873 (.Y (out_column_2__1), .A0 (nx3868), .A1 (nx3842), .A2 (nx3814)
         , .A3 (nx3788)) ;
    nand03 ix3869 (.Y (nx3868), .A0 (nx8141), .A1 (nx8143), .A2 (nx8145)) ;
    aoi222 ix8142 (.Y (nx8141), .A0 (que_out_10__2__1), .A1 (nx10306), .B0 (
           que_out_6__2__1), .B1 (nx10358), .C0 (que_out_9__2__1), .C1 (nx10332)
           ) ;
    aoi22 ix8144 (.Y (nx8143), .A0 (que_out_5__2__1), .A1 (nx10254), .B0 (
          que_out_18__2__1), .B1 (nx10280)) ;
    aoi22 ix8146 (.Y (nx8145), .A0 (que_out_17__2__1), .A1 (nx10228), .B0 (
          que_out_20__2__1), .B1 (nx10202)) ;
    nand03 ix3843 (.Y (nx3842), .A0 (nx8149), .A1 (nx8151), .A2 (nx8153)) ;
    aoi222 ix8150 (.Y (nx8149), .A0 (que_out_19__2__1), .A1 (nx10176), .B0 (
           que_out_21__2__1), .B1 (nx10150), .C0 (que_out_8__2__1), .C1 (nx10124
           )) ;
    aoi22 ix8152 (.Y (nx8151), .A0 (que_out_25__2__1), .A1 (nx10072), .B0 (
          que_out_16__2__1), .B1 (nx10098)) ;
    aoi22 ix8154 (.Y (nx8153), .A0 (que_out_24__2__1), .A1 (nx10046), .B0 (
          que_out_22__2__1), .B1 (nx10020)) ;
    nand03 ix3815 (.Y (nx3814), .A0 (nx8157), .A1 (nx8159), .A2 (nx8161)) ;
    aoi222 ix8158 (.Y (nx8157), .A0 (que_out_15__2__1), .A1 (nx9968), .B0 (
           que_out_3__2__1), .B1 (nx9994), .C0 (que_out_23__2__1), .C1 (nx9942)
           ) ;
    aoi22 ix8160 (.Y (nx8159), .A0 (que_out_27__2__1), .A1 (nx9916), .B0 (
          que_out_4__2__1), .B1 (nx9890)) ;
    aoi22 ix8162 (.Y (nx8161), .A0 (que_out_0__2__1), .A1 (nx9838), .B0 (
          que_out_2__2__1), .B1 (nx9864)) ;
    nand03 ix3789 (.Y (nx3788), .A0 (nx8165), .A1 (nx8167), .A2 (nx8169)) ;
    aoi222 ix8166 (.Y (nx8165), .A0 (que_out_26__2__1), .A1 (nx9812), .B0 (
           que_out_14__2__1), .B1 (nx9786), .C0 (que_out_11__2__1), .C1 (nx9760)
           ) ;
    aoi22 ix8168 (.Y (nx8167), .A0 (que_out_13__2__1), .A1 (nx9734), .B0 (
          que_out_7__2__1), .B1 (nx9708)) ;
    aoi22 ix8170 (.Y (nx8169), .A0 (que_out_12__2__1), .A1 (nx9682), .B0 (
          que_out_1__2__1), .B1 (nx9656)) ;
    or04 ix3983 (.Y (out_column_2__2), .A0 (nx3978), .A1 (nx3952), .A2 (nx3924)
         , .A3 (nx3898)) ;
    nand03 ix3979 (.Y (nx3978), .A0 (nx8175), .A1 (nx8177), .A2 (nx8179)) ;
    aoi222 ix8176 (.Y (nx8175), .A0 (que_out_10__2__2), .A1 (nx10306), .B0 (
           que_out_6__2__2), .B1 (nx10358), .C0 (que_out_9__2__2), .C1 (nx10332)
           ) ;
    aoi22 ix8178 (.Y (nx8177), .A0 (que_out_5__2__2), .A1 (nx10254), .B0 (
          que_out_18__2__2), .B1 (nx10280)) ;
    aoi22 ix8180 (.Y (nx8179), .A0 (que_out_17__2__2), .A1 (nx10228), .B0 (
          que_out_20__2__2), .B1 (nx10202)) ;
    nand03 ix3953 (.Y (nx3952), .A0 (nx8183), .A1 (nx8185), .A2 (nx8187)) ;
    aoi222 ix8184 (.Y (nx8183), .A0 (que_out_19__2__2), .A1 (nx10176), .B0 (
           que_out_21__2__2), .B1 (nx10150), .C0 (que_out_8__2__2), .C1 (nx10124
           )) ;
    aoi22 ix8186 (.Y (nx8185), .A0 (que_out_25__2__2), .A1 (nx10072), .B0 (
          que_out_16__2__2), .B1 (nx10098)) ;
    aoi22 ix8188 (.Y (nx8187), .A0 (que_out_24__2__2), .A1 (nx10046), .B0 (
          que_out_22__2__2), .B1 (nx10020)) ;
    nand03 ix3925 (.Y (nx3924), .A0 (nx8191), .A1 (nx8193), .A2 (nx8195)) ;
    aoi222 ix8192 (.Y (nx8191), .A0 (que_out_15__2__2), .A1 (nx9968), .B0 (
           que_out_3__2__2), .B1 (nx9994), .C0 (que_out_23__2__2), .C1 (nx9942)
           ) ;
    aoi22 ix8194 (.Y (nx8193), .A0 (que_out_27__2__2), .A1 (nx9916), .B0 (
          que_out_4__2__2), .B1 (nx9890)) ;
    aoi22 ix8196 (.Y (nx8195), .A0 (que_out_0__2__2), .A1 (nx9838), .B0 (
          que_out_2__2__2), .B1 (nx9864)) ;
    nand03 ix3899 (.Y (nx3898), .A0 (nx8199), .A1 (nx8201), .A2 (nx8203)) ;
    aoi222 ix8200 (.Y (nx8199), .A0 (que_out_26__2__2), .A1 (nx9812), .B0 (
           que_out_14__2__2), .B1 (nx9786), .C0 (que_out_11__2__2), .C1 (nx9760)
           ) ;
    aoi22 ix8202 (.Y (nx8201), .A0 (que_out_13__2__2), .A1 (nx9734), .B0 (
          que_out_7__2__2), .B1 (nx9708)) ;
    aoi22 ix8204 (.Y (nx8203), .A0 (que_out_12__2__2), .A1 (nx9682), .B0 (
          que_out_1__2__2), .B1 (nx9656)) ;
    or04 ix4093 (.Y (out_column_2__3), .A0 (nx4088), .A1 (nx4062), .A2 (nx4034)
         , .A3 (nx4008)) ;
    nand03 ix4089 (.Y (nx4088), .A0 (nx8209), .A1 (nx8211), .A2 (nx8213)) ;
    aoi222 ix8210 (.Y (nx8209), .A0 (que_out_10__2__3), .A1 (nx10308), .B0 (
           que_out_6__2__3), .B1 (nx10360), .C0 (que_out_9__2__3), .C1 (nx10334)
           ) ;
    aoi22 ix8212 (.Y (nx8211), .A0 (que_out_5__2__3), .A1 (nx10256), .B0 (
          que_out_18__2__3), .B1 (nx10282)) ;
    aoi22 ix8214 (.Y (nx8213), .A0 (que_out_17__2__3), .A1 (nx10230), .B0 (
          que_out_20__2__3), .B1 (nx10204)) ;
    nand03 ix4063 (.Y (nx4062), .A0 (nx8217), .A1 (nx8219), .A2 (nx8221)) ;
    aoi222 ix8218 (.Y (nx8217), .A0 (que_out_19__2__3), .A1 (nx10178), .B0 (
           que_out_21__2__3), .B1 (nx10152), .C0 (que_out_8__2__3), .C1 (nx10126
           )) ;
    aoi22 ix8220 (.Y (nx8219), .A0 (que_out_25__2__3), .A1 (nx10074), .B0 (
          que_out_16__2__3), .B1 (nx10100)) ;
    aoi22 ix8222 (.Y (nx8221), .A0 (que_out_24__2__3), .A1 (nx10048), .B0 (
          que_out_22__2__3), .B1 (nx10022)) ;
    nand03 ix4035 (.Y (nx4034), .A0 (nx8225), .A1 (nx8227), .A2 (nx8229)) ;
    aoi222 ix8226 (.Y (nx8225), .A0 (que_out_15__2__3), .A1 (nx9970), .B0 (
           que_out_3__2__3), .B1 (nx9996), .C0 (que_out_23__2__3), .C1 (nx9944)
           ) ;
    aoi22 ix8228 (.Y (nx8227), .A0 (que_out_27__2__3), .A1 (nx9918), .B0 (
          que_out_4__2__3), .B1 (nx9892)) ;
    aoi22 ix8230 (.Y (nx8229), .A0 (que_out_0__2__3), .A1 (nx9840), .B0 (
          que_out_2__2__3), .B1 (nx9866)) ;
    nand03 ix4009 (.Y (nx4008), .A0 (nx8233), .A1 (nx8235), .A2 (nx8237)) ;
    aoi222 ix8234 (.Y (nx8233), .A0 (que_out_26__2__3), .A1 (nx9814), .B0 (
           que_out_14__2__3), .B1 (nx9788), .C0 (que_out_11__2__3), .C1 (nx9762)
           ) ;
    aoi22 ix8236 (.Y (nx8235), .A0 (que_out_13__2__3), .A1 (nx9736), .B0 (
          que_out_7__2__3), .B1 (nx9710)) ;
    aoi22 ix8238 (.Y (nx8237), .A0 (que_out_12__2__3), .A1 (nx9684), .B0 (
          que_out_1__2__3), .B1 (nx9658)) ;
    or04 ix4203 (.Y (out_column_2__4), .A0 (nx4198), .A1 (nx4172), .A2 (nx4144)
         , .A3 (nx4118)) ;
    nand03 ix4199 (.Y (nx4198), .A0 (nx8243), .A1 (nx8245), .A2 (nx8247)) ;
    aoi222 ix8244 (.Y (nx8243), .A0 (que_out_10__2__4), .A1 (nx10308), .B0 (
           que_out_6__2__4), .B1 (nx10360), .C0 (que_out_9__2__4), .C1 (nx10334)
           ) ;
    aoi22 ix8246 (.Y (nx8245), .A0 (que_out_5__2__4), .A1 (nx10256), .B0 (
          que_out_18__2__4), .B1 (nx10282)) ;
    aoi22 ix8248 (.Y (nx8247), .A0 (que_out_17__2__4), .A1 (nx10230), .B0 (
          que_out_20__2__4), .B1 (nx10204)) ;
    nand03 ix4173 (.Y (nx4172), .A0 (nx8251), .A1 (nx8253), .A2 (nx8255)) ;
    aoi222 ix8252 (.Y (nx8251), .A0 (que_out_19__2__4), .A1 (nx10178), .B0 (
           que_out_21__2__4), .B1 (nx10152), .C0 (que_out_8__2__4), .C1 (nx10126
           )) ;
    aoi22 ix8254 (.Y (nx8253), .A0 (que_out_25__2__4), .A1 (nx10074), .B0 (
          que_out_16__2__4), .B1 (nx10100)) ;
    aoi22 ix8256 (.Y (nx8255), .A0 (que_out_24__2__4), .A1 (nx10048), .B0 (
          que_out_22__2__4), .B1 (nx10022)) ;
    nand03 ix4145 (.Y (nx4144), .A0 (nx8259), .A1 (nx8261), .A2 (nx8263)) ;
    aoi222 ix8260 (.Y (nx8259), .A0 (que_out_15__2__4), .A1 (nx9970), .B0 (
           que_out_3__2__4), .B1 (nx9996), .C0 (que_out_23__2__4), .C1 (nx9944)
           ) ;
    aoi22 ix8262 (.Y (nx8261), .A0 (que_out_27__2__4), .A1 (nx9918), .B0 (
          que_out_4__2__4), .B1 (nx9892)) ;
    aoi22 ix8264 (.Y (nx8263), .A0 (que_out_0__2__4), .A1 (nx9840), .B0 (
          que_out_2__2__4), .B1 (nx9866)) ;
    nand03 ix4119 (.Y (nx4118), .A0 (nx8267), .A1 (nx8269), .A2 (nx8271)) ;
    aoi222 ix8268 (.Y (nx8267), .A0 (que_out_26__2__4), .A1 (nx9814), .B0 (
           que_out_14__2__4), .B1 (nx9788), .C0 (que_out_11__2__4), .C1 (nx9762)
           ) ;
    aoi22 ix8270 (.Y (nx8269), .A0 (que_out_13__2__4), .A1 (nx9736), .B0 (
          que_out_7__2__4), .B1 (nx9710)) ;
    aoi22 ix8272 (.Y (nx8271), .A0 (que_out_12__2__4), .A1 (nx9684), .B0 (
          que_out_1__2__4), .B1 (nx9658)) ;
    or04 ix4313 (.Y (out_column_2__5), .A0 (nx4308), .A1 (nx4282), .A2 (nx4254)
         , .A3 (nx4228)) ;
    nand03 ix4309 (.Y (nx4308), .A0 (nx8277), .A1 (nx8279), .A2 (nx8281)) ;
    aoi222 ix8278 (.Y (nx8277), .A0 (que_out_10__2__5), .A1 (nx10308), .B0 (
           que_out_6__2__5), .B1 (nx10360), .C0 (que_out_9__2__5), .C1 (nx10334)
           ) ;
    aoi22 ix8280 (.Y (nx8279), .A0 (que_out_5__2__5), .A1 (nx10256), .B0 (
          que_out_18__2__5), .B1 (nx10282)) ;
    aoi22 ix8282 (.Y (nx8281), .A0 (que_out_17__2__5), .A1 (nx10230), .B0 (
          que_out_20__2__5), .B1 (nx10204)) ;
    nand03 ix4283 (.Y (nx4282), .A0 (nx8285), .A1 (nx8287), .A2 (nx8289)) ;
    aoi222 ix8286 (.Y (nx8285), .A0 (que_out_19__2__5), .A1 (nx10178), .B0 (
           que_out_21__2__5), .B1 (nx10152), .C0 (que_out_8__2__5), .C1 (nx10126
           )) ;
    aoi22 ix8288 (.Y (nx8287), .A0 (que_out_25__2__5), .A1 (nx10074), .B0 (
          que_out_16__2__5), .B1 (nx10100)) ;
    aoi22 ix8290 (.Y (nx8289), .A0 (que_out_24__2__5), .A1 (nx10048), .B0 (
          que_out_22__2__5), .B1 (nx10022)) ;
    nand03 ix4255 (.Y (nx4254), .A0 (nx8293), .A1 (nx8295), .A2 (nx8297)) ;
    aoi222 ix8294 (.Y (nx8293), .A0 (que_out_15__2__5), .A1 (nx9970), .B0 (
           que_out_3__2__5), .B1 (nx9996), .C0 (que_out_23__2__5), .C1 (nx9944)
           ) ;
    aoi22 ix8296 (.Y (nx8295), .A0 (que_out_27__2__5), .A1 (nx9918), .B0 (
          que_out_4__2__5), .B1 (nx9892)) ;
    aoi22 ix8298 (.Y (nx8297), .A0 (que_out_0__2__5), .A1 (nx9840), .B0 (
          que_out_2__2__5), .B1 (nx9866)) ;
    nand03 ix4229 (.Y (nx4228), .A0 (nx8301), .A1 (nx8303), .A2 (nx8305)) ;
    aoi222 ix8302 (.Y (nx8301), .A0 (que_out_26__2__5), .A1 (nx9814), .B0 (
           que_out_14__2__5), .B1 (nx9788), .C0 (que_out_11__2__5), .C1 (nx9762)
           ) ;
    aoi22 ix8304 (.Y (nx8303), .A0 (que_out_13__2__5), .A1 (nx9736), .B0 (
          que_out_7__2__5), .B1 (nx9710)) ;
    aoi22 ix8306 (.Y (nx8305), .A0 (que_out_12__2__5), .A1 (nx9684), .B0 (
          que_out_1__2__5), .B1 (nx9658)) ;
    or04 ix4423 (.Y (out_column_2__6), .A0 (nx4418), .A1 (nx4392), .A2 (nx4364)
         , .A3 (nx4338)) ;
    nand03 ix4419 (.Y (nx4418), .A0 (nx8311), .A1 (nx8313), .A2 (nx8315)) ;
    aoi222 ix8312 (.Y (nx8311), .A0 (que_out_10__2__6), .A1 (nx10308), .B0 (
           que_out_6__2__6), .B1 (nx10360), .C0 (que_out_9__2__6), .C1 (nx10334)
           ) ;
    aoi22 ix8314 (.Y (nx8313), .A0 (que_out_5__2__6), .A1 (nx10256), .B0 (
          que_out_18__2__6), .B1 (nx10282)) ;
    aoi22 ix8316 (.Y (nx8315), .A0 (que_out_17__2__6), .A1 (nx10230), .B0 (
          que_out_20__2__6), .B1 (nx10204)) ;
    nand03 ix4393 (.Y (nx4392), .A0 (nx8319), .A1 (nx8321), .A2 (nx8323)) ;
    aoi222 ix8320 (.Y (nx8319), .A0 (que_out_19__2__6), .A1 (nx10178), .B0 (
           que_out_21__2__6), .B1 (nx10152), .C0 (que_out_8__2__6), .C1 (nx10126
           )) ;
    aoi22 ix8322 (.Y (nx8321), .A0 (que_out_25__2__6), .A1 (nx10074), .B0 (
          que_out_16__2__6), .B1 (nx10100)) ;
    aoi22 ix8324 (.Y (nx8323), .A0 (que_out_24__2__6), .A1 (nx10048), .B0 (
          que_out_22__2__6), .B1 (nx10022)) ;
    nand03 ix4365 (.Y (nx4364), .A0 (nx8327), .A1 (nx8329), .A2 (nx8331)) ;
    aoi222 ix8328 (.Y (nx8327), .A0 (que_out_15__2__6), .A1 (nx9970), .B0 (
           que_out_3__2__6), .B1 (nx9996), .C0 (que_out_23__2__6), .C1 (nx9944)
           ) ;
    aoi22 ix8330 (.Y (nx8329), .A0 (que_out_27__2__6), .A1 (nx9918), .B0 (
          que_out_4__2__6), .B1 (nx9892)) ;
    aoi22 ix8332 (.Y (nx8331), .A0 (que_out_0__2__6), .A1 (nx9840), .B0 (
          que_out_2__2__6), .B1 (nx9866)) ;
    nand03 ix4339 (.Y (nx4338), .A0 (nx8335), .A1 (nx8337), .A2 (nx8339)) ;
    aoi222 ix8336 (.Y (nx8335), .A0 (que_out_26__2__6), .A1 (nx9814), .B0 (
           que_out_14__2__6), .B1 (nx9788), .C0 (que_out_11__2__6), .C1 (nx9762)
           ) ;
    aoi22 ix8338 (.Y (nx8337), .A0 (que_out_13__2__6), .A1 (nx9736), .B0 (
          que_out_7__2__6), .B1 (nx9710)) ;
    aoi22 ix8340 (.Y (nx8339), .A0 (que_out_12__2__6), .A1 (nx9684), .B0 (
          que_out_1__2__6), .B1 (nx9658)) ;
    or04 ix4533 (.Y (out_column_2__7), .A0 (nx4528), .A1 (nx4502), .A2 (nx4474)
         , .A3 (nx4448)) ;
    nand03 ix4529 (.Y (nx4528), .A0 (nx8345), .A1 (nx8347), .A2 (nx8349)) ;
    aoi222 ix8346 (.Y (nx8345), .A0 (que_out_10__2__7), .A1 (nx10308), .B0 (
           que_out_6__2__7), .B1 (nx10360), .C0 (que_out_9__2__7), .C1 (nx10334)
           ) ;
    aoi22 ix8348 (.Y (nx8347), .A0 (que_out_5__2__7), .A1 (nx10256), .B0 (
          que_out_18__2__7), .B1 (nx10282)) ;
    aoi22 ix8350 (.Y (nx8349), .A0 (que_out_17__2__7), .A1 (nx10230), .B0 (
          que_out_20__2__7), .B1 (nx10204)) ;
    nand03 ix4503 (.Y (nx4502), .A0 (nx8353), .A1 (nx8355), .A2 (nx8357)) ;
    aoi222 ix8354 (.Y (nx8353), .A0 (que_out_19__2__7), .A1 (nx10178), .B0 (
           que_out_21__2__7), .B1 (nx10152), .C0 (que_out_8__2__7), .C1 (nx10126
           )) ;
    aoi22 ix8356 (.Y (nx8355), .A0 (que_out_25__2__7), .A1 (nx10074), .B0 (
          que_out_16__2__7), .B1 (nx10100)) ;
    aoi22 ix8358 (.Y (nx8357), .A0 (que_out_24__2__7), .A1 (nx10048), .B0 (
          que_out_22__2__7), .B1 (nx10022)) ;
    nand03 ix4475 (.Y (nx4474), .A0 (nx8361), .A1 (nx8363), .A2 (nx8365)) ;
    aoi222 ix8362 (.Y (nx8361), .A0 (que_out_15__2__7), .A1 (nx9970), .B0 (
           que_out_3__2__7), .B1 (nx9996), .C0 (que_out_23__2__7), .C1 (nx9944)
           ) ;
    aoi22 ix8364 (.Y (nx8363), .A0 (que_out_27__2__7), .A1 (nx9918), .B0 (
          que_out_4__2__7), .B1 (nx9892)) ;
    aoi22 ix8366 (.Y (nx8365), .A0 (que_out_0__2__7), .A1 (nx9840), .B0 (
          que_out_2__2__7), .B1 (nx9866)) ;
    nand03 ix4449 (.Y (nx4448), .A0 (nx8369), .A1 (nx8371), .A2 (nx8373)) ;
    aoi222 ix8370 (.Y (nx8369), .A0 (que_out_26__2__7), .A1 (nx9814), .B0 (
           que_out_14__2__7), .B1 (nx9788), .C0 (que_out_11__2__7), .C1 (nx9762)
           ) ;
    aoi22 ix8372 (.Y (nx8371), .A0 (que_out_13__2__7), .A1 (nx9736), .B0 (
          que_out_7__2__7), .B1 (nx9710)) ;
    aoi22 ix8374 (.Y (nx8373), .A0 (que_out_12__2__7), .A1 (nx9684), .B0 (
          que_out_1__2__7), .B1 (nx9658)) ;
    or04 ix4643 (.Y (out_column_2__8), .A0 (nx4638), .A1 (nx4612), .A2 (nx4584)
         , .A3 (nx4558)) ;
    nand03 ix4639 (.Y (nx4638), .A0 (nx8379), .A1 (nx8381), .A2 (nx8383)) ;
    aoi222 ix8380 (.Y (nx8379), .A0 (que_out_10__2__8), .A1 (nx10308), .B0 (
           que_out_6__2__8), .B1 (nx10360), .C0 (que_out_9__2__8), .C1 (nx10334)
           ) ;
    aoi22 ix8382 (.Y (nx8381), .A0 (que_out_5__2__8), .A1 (nx10256), .B0 (
          que_out_18__2__8), .B1 (nx10282)) ;
    aoi22 ix8384 (.Y (nx8383), .A0 (que_out_17__2__8), .A1 (nx10230), .B0 (
          que_out_20__2__8), .B1 (nx10204)) ;
    nand03 ix4613 (.Y (nx4612), .A0 (nx8387), .A1 (nx8389), .A2 (nx8391)) ;
    aoi222 ix8388 (.Y (nx8387), .A0 (que_out_19__2__8), .A1 (nx10178), .B0 (
           que_out_21__2__8), .B1 (nx10152), .C0 (que_out_8__2__8), .C1 (nx10126
           )) ;
    aoi22 ix8390 (.Y (nx8389), .A0 (que_out_25__2__8), .A1 (nx10074), .B0 (
          que_out_16__2__8), .B1 (nx10100)) ;
    aoi22 ix8392 (.Y (nx8391), .A0 (que_out_24__2__8), .A1 (nx10048), .B0 (
          que_out_22__2__8), .B1 (nx10022)) ;
    nand03 ix4585 (.Y (nx4584), .A0 (nx8395), .A1 (nx8397), .A2 (nx8399)) ;
    aoi222 ix8396 (.Y (nx8395), .A0 (que_out_15__2__8), .A1 (nx9970), .B0 (
           que_out_3__2__8), .B1 (nx9996), .C0 (que_out_23__2__8), .C1 (nx9944)
           ) ;
    aoi22 ix8398 (.Y (nx8397), .A0 (que_out_27__2__8), .A1 (nx9918), .B0 (
          que_out_4__2__8), .B1 (nx9892)) ;
    aoi22 ix8400 (.Y (nx8399), .A0 (que_out_0__2__8), .A1 (nx9840), .B0 (
          que_out_2__2__8), .B1 (nx9866)) ;
    nand03 ix4559 (.Y (nx4558), .A0 (nx8403), .A1 (nx8405), .A2 (nx8407)) ;
    aoi222 ix8404 (.Y (nx8403), .A0 (que_out_26__2__8), .A1 (nx9814), .B0 (
           que_out_14__2__8), .B1 (nx9788), .C0 (que_out_11__2__8), .C1 (nx9762)
           ) ;
    aoi22 ix8406 (.Y (nx8405), .A0 (que_out_13__2__8), .A1 (nx9736), .B0 (
          que_out_7__2__8), .B1 (nx9710)) ;
    aoi22 ix8408 (.Y (nx8407), .A0 (que_out_12__2__8), .A1 (nx9684), .B0 (
          que_out_1__2__8), .B1 (nx9658)) ;
    or04 ix4753 (.Y (out_column_2__9), .A0 (nx4748), .A1 (nx4722), .A2 (nx4694)
         , .A3 (nx4668)) ;
    nand03 ix4749 (.Y (nx4748), .A0 (nx8413), .A1 (nx8415), .A2 (nx8417)) ;
    aoi222 ix8414 (.Y (nx8413), .A0 (que_out_10__2__9), .A1 (nx10308), .B0 (
           que_out_6__2__9), .B1 (nx10360), .C0 (que_out_9__2__9), .C1 (nx10334)
           ) ;
    aoi22 ix8416 (.Y (nx8415), .A0 (que_out_5__2__9), .A1 (nx10256), .B0 (
          que_out_18__2__9), .B1 (nx10282)) ;
    aoi22 ix8418 (.Y (nx8417), .A0 (que_out_17__2__9), .A1 (nx10230), .B0 (
          que_out_20__2__9), .B1 (nx10204)) ;
    nand03 ix4723 (.Y (nx4722), .A0 (nx8421), .A1 (nx8423), .A2 (nx8425)) ;
    aoi222 ix8422 (.Y (nx8421), .A0 (que_out_19__2__9), .A1 (nx10178), .B0 (
           que_out_21__2__9), .B1 (nx10152), .C0 (que_out_8__2__9), .C1 (nx10126
           )) ;
    aoi22 ix8424 (.Y (nx8423), .A0 (que_out_25__2__9), .A1 (nx10074), .B0 (
          que_out_16__2__9), .B1 (nx10100)) ;
    aoi22 ix8426 (.Y (nx8425), .A0 (que_out_24__2__9), .A1 (nx10048), .B0 (
          que_out_22__2__9), .B1 (nx10022)) ;
    nand03 ix4695 (.Y (nx4694), .A0 (nx8429), .A1 (nx8431), .A2 (nx8433)) ;
    aoi222 ix8430 (.Y (nx8429), .A0 (que_out_15__2__9), .A1 (nx9970), .B0 (
           que_out_3__2__9), .B1 (nx9996), .C0 (que_out_23__2__9), .C1 (nx9944)
           ) ;
    aoi22 ix8432 (.Y (nx8431), .A0 (que_out_27__2__9), .A1 (nx9918), .B0 (
          que_out_4__2__9), .B1 (nx9892)) ;
    aoi22 ix8434 (.Y (nx8433), .A0 (que_out_0__2__9), .A1 (nx9840), .B0 (
          que_out_2__2__9), .B1 (nx9866)) ;
    nand03 ix4669 (.Y (nx4668), .A0 (nx8437), .A1 (nx8439), .A2 (nx8441)) ;
    aoi222 ix8438 (.Y (nx8437), .A0 (que_out_26__2__9), .A1 (nx9814), .B0 (
           que_out_14__2__9), .B1 (nx9788), .C0 (que_out_11__2__9), .C1 (nx9762)
           ) ;
    aoi22 ix8440 (.Y (nx8439), .A0 (que_out_13__2__9), .A1 (nx9736), .B0 (
          que_out_7__2__9), .B1 (nx9710)) ;
    aoi22 ix8442 (.Y (nx8441), .A0 (que_out_12__2__9), .A1 (nx9684), .B0 (
          que_out_1__2__9), .B1 (nx9658)) ;
    or04 ix4863 (.Y (out_column_2__10), .A0 (nx4858), .A1 (nx4832), .A2 (nx4804)
         , .A3 (nx4778)) ;
    nand03 ix4859 (.Y (nx4858), .A0 (nx8447), .A1 (nx8449), .A2 (nx8451)) ;
    aoi222 ix8448 (.Y (nx8447), .A0 (que_out_10__2__10), .A1 (nx10310), .B0 (
           que_out_6__2__10), .B1 (nx10362), .C0 (que_out_9__2__10), .C1 (
           nx10336)) ;
    aoi22 ix8450 (.Y (nx8449), .A0 (que_out_5__2__10), .A1 (nx10258), .B0 (
          que_out_18__2__10), .B1 (nx10284)) ;
    aoi22 ix8452 (.Y (nx8451), .A0 (que_out_17__2__10), .A1 (nx10232), .B0 (
          que_out_20__2__10), .B1 (nx10206)) ;
    nand03 ix4833 (.Y (nx4832), .A0 (nx8455), .A1 (nx8457), .A2 (nx8459)) ;
    aoi222 ix8456 (.Y (nx8455), .A0 (que_out_19__2__10), .A1 (nx10180), .B0 (
           que_out_21__2__10), .B1 (nx10154), .C0 (que_out_8__2__10), .C1 (
           nx10128)) ;
    aoi22 ix8458 (.Y (nx8457), .A0 (que_out_25__2__10), .A1 (nx10076), .B0 (
          que_out_16__2__10), .B1 (nx10102)) ;
    aoi22 ix8460 (.Y (nx8459), .A0 (que_out_24__2__10), .A1 (nx10050), .B0 (
          que_out_22__2__10), .B1 (nx10024)) ;
    nand03 ix4805 (.Y (nx4804), .A0 (nx8463), .A1 (nx8465), .A2 (nx8467)) ;
    aoi222 ix8464 (.Y (nx8463), .A0 (que_out_15__2__10), .A1 (nx9972), .B0 (
           que_out_3__2__10), .B1 (nx9998), .C0 (que_out_23__2__10), .C1 (nx9946
           )) ;
    aoi22 ix8466 (.Y (nx8465), .A0 (que_out_27__2__10), .A1 (nx9920), .B0 (
          que_out_4__2__10), .B1 (nx9894)) ;
    aoi22 ix8468 (.Y (nx8467), .A0 (que_out_0__2__10), .A1 (nx9842), .B0 (
          que_out_2__2__10), .B1 (nx9868)) ;
    nand03 ix4779 (.Y (nx4778), .A0 (nx8471), .A1 (nx8473), .A2 (nx8475)) ;
    aoi222 ix8472 (.Y (nx8471), .A0 (que_out_26__2__10), .A1 (nx9816), .B0 (
           que_out_14__2__10), .B1 (nx9790), .C0 (que_out_11__2__10), .C1 (
           nx9764)) ;
    aoi22 ix8474 (.Y (nx8473), .A0 (que_out_13__2__10), .A1 (nx9738), .B0 (
          que_out_7__2__10), .B1 (nx9712)) ;
    aoi22 ix8476 (.Y (nx8475), .A0 (que_out_12__2__10), .A1 (nx9686), .B0 (
          que_out_1__2__10), .B1 (nx9660)) ;
    or04 ix4973 (.Y (out_column_2__11), .A0 (nx4968), .A1 (nx4942), .A2 (nx4914)
         , .A3 (nx4888)) ;
    nand03 ix4969 (.Y (nx4968), .A0 (nx8481), .A1 (nx8483), .A2 (nx8485)) ;
    aoi222 ix8482 (.Y (nx8481), .A0 (que_out_10__2__11), .A1 (nx10310), .B0 (
           que_out_6__2__11), .B1 (nx10362), .C0 (que_out_9__2__11), .C1 (
           nx10336)) ;
    aoi22 ix8484 (.Y (nx8483), .A0 (que_out_5__2__11), .A1 (nx10258), .B0 (
          que_out_18__2__11), .B1 (nx10284)) ;
    aoi22 ix8486 (.Y (nx8485), .A0 (que_out_17__2__11), .A1 (nx10232), .B0 (
          que_out_20__2__11), .B1 (nx10206)) ;
    nand03 ix4943 (.Y (nx4942), .A0 (nx8489), .A1 (nx8491), .A2 (nx8493)) ;
    aoi222 ix8490 (.Y (nx8489), .A0 (que_out_19__2__11), .A1 (nx10180), .B0 (
           que_out_21__2__11), .B1 (nx10154), .C0 (que_out_8__2__11), .C1 (
           nx10128)) ;
    aoi22 ix8492 (.Y (nx8491), .A0 (que_out_25__2__11), .A1 (nx10076), .B0 (
          que_out_16__2__11), .B1 (nx10102)) ;
    aoi22 ix8494 (.Y (nx8493), .A0 (que_out_24__2__11), .A1 (nx10050), .B0 (
          que_out_22__2__11), .B1 (nx10024)) ;
    nand03 ix4915 (.Y (nx4914), .A0 (nx8497), .A1 (nx8499), .A2 (nx8501)) ;
    aoi222 ix8498 (.Y (nx8497), .A0 (que_out_15__2__11), .A1 (nx9972), .B0 (
           que_out_3__2__11), .B1 (nx9998), .C0 (que_out_23__2__11), .C1 (nx9946
           )) ;
    aoi22 ix8500 (.Y (nx8499), .A0 (que_out_27__2__11), .A1 (nx9920), .B0 (
          que_out_4__2__11), .B1 (nx9894)) ;
    aoi22 ix8502 (.Y (nx8501), .A0 (que_out_0__2__11), .A1 (nx9842), .B0 (
          que_out_2__2__11), .B1 (nx9868)) ;
    nand03 ix4889 (.Y (nx4888), .A0 (nx8505), .A1 (nx8507), .A2 (nx8509)) ;
    aoi222 ix8506 (.Y (nx8505), .A0 (que_out_26__2__11), .A1 (nx9816), .B0 (
           que_out_14__2__11), .B1 (nx9790), .C0 (que_out_11__2__11), .C1 (
           nx9764)) ;
    aoi22 ix8508 (.Y (nx8507), .A0 (que_out_13__2__11), .A1 (nx9738), .B0 (
          que_out_7__2__11), .B1 (nx9712)) ;
    aoi22 ix8510 (.Y (nx8509), .A0 (que_out_12__2__11), .A1 (nx9686), .B0 (
          que_out_1__2__11), .B1 (nx9660)) ;
    or04 ix5083 (.Y (out_column_2__12), .A0 (nx5078), .A1 (nx5052), .A2 (nx5024)
         , .A3 (nx4998)) ;
    nand03 ix5079 (.Y (nx5078), .A0 (nx8515), .A1 (nx8517), .A2 (nx8519)) ;
    aoi222 ix8516 (.Y (nx8515), .A0 (que_out_10__2__12), .A1 (nx10310), .B0 (
           que_out_6__2__12), .B1 (nx10362), .C0 (que_out_9__2__12), .C1 (
           nx10336)) ;
    aoi22 ix8518 (.Y (nx8517), .A0 (que_out_5__2__12), .A1 (nx10258), .B0 (
          que_out_18__2__12), .B1 (nx10284)) ;
    aoi22 ix8520 (.Y (nx8519), .A0 (que_out_17__2__12), .A1 (nx10232), .B0 (
          que_out_20__2__12), .B1 (nx10206)) ;
    nand03 ix5053 (.Y (nx5052), .A0 (nx8523), .A1 (nx8525), .A2 (nx8527)) ;
    aoi222 ix8524 (.Y (nx8523), .A0 (que_out_19__2__12), .A1 (nx10180), .B0 (
           que_out_21__2__12), .B1 (nx10154), .C0 (que_out_8__2__12), .C1 (
           nx10128)) ;
    aoi22 ix8526 (.Y (nx8525), .A0 (que_out_25__2__12), .A1 (nx10076), .B0 (
          que_out_16__2__12), .B1 (nx10102)) ;
    aoi22 ix8528 (.Y (nx8527), .A0 (que_out_24__2__12), .A1 (nx10050), .B0 (
          que_out_22__2__12), .B1 (nx10024)) ;
    nand03 ix5025 (.Y (nx5024), .A0 (nx8531), .A1 (nx8533), .A2 (nx8535)) ;
    aoi222 ix8532 (.Y (nx8531), .A0 (que_out_15__2__12), .A1 (nx9972), .B0 (
           que_out_3__2__12), .B1 (nx9998), .C0 (que_out_23__2__12), .C1 (nx9946
           )) ;
    aoi22 ix8534 (.Y (nx8533), .A0 (que_out_27__2__12), .A1 (nx9920), .B0 (
          que_out_4__2__12), .B1 (nx9894)) ;
    aoi22 ix8536 (.Y (nx8535), .A0 (que_out_0__2__12), .A1 (nx9842), .B0 (
          que_out_2__2__12), .B1 (nx9868)) ;
    nand03 ix4999 (.Y (nx4998), .A0 (nx8539), .A1 (nx8541), .A2 (nx8543)) ;
    aoi222 ix8540 (.Y (nx8539), .A0 (que_out_26__2__12), .A1 (nx9816), .B0 (
           que_out_14__2__12), .B1 (nx9790), .C0 (que_out_11__2__12), .C1 (
           nx9764)) ;
    aoi22 ix8542 (.Y (nx8541), .A0 (que_out_13__2__12), .A1 (nx9738), .B0 (
          que_out_7__2__12), .B1 (nx9712)) ;
    aoi22 ix8544 (.Y (nx8543), .A0 (que_out_12__2__12), .A1 (nx9686), .B0 (
          que_out_1__2__12), .B1 (nx9660)) ;
    or04 ix5193 (.Y (out_column_2__13), .A0 (nx5188), .A1 (nx5162), .A2 (nx5134)
         , .A3 (nx5108)) ;
    nand03 ix5189 (.Y (nx5188), .A0 (nx8549), .A1 (nx8551), .A2 (nx8553)) ;
    aoi222 ix8550 (.Y (nx8549), .A0 (que_out_10__2__13), .A1 (nx10310), .B0 (
           que_out_6__2__13), .B1 (nx10362), .C0 (que_out_9__2__13), .C1 (
           nx10336)) ;
    aoi22 ix8552 (.Y (nx8551), .A0 (que_out_5__2__13), .A1 (nx10258), .B0 (
          que_out_18__2__13), .B1 (nx10284)) ;
    aoi22 ix8554 (.Y (nx8553), .A0 (que_out_17__2__13), .A1 (nx10232), .B0 (
          que_out_20__2__13), .B1 (nx10206)) ;
    nand03 ix5163 (.Y (nx5162), .A0 (nx8557), .A1 (nx8559), .A2 (nx8561)) ;
    aoi222 ix8558 (.Y (nx8557), .A0 (que_out_19__2__13), .A1 (nx10180), .B0 (
           que_out_21__2__13), .B1 (nx10154), .C0 (que_out_8__2__13), .C1 (
           nx10128)) ;
    aoi22 ix8560 (.Y (nx8559), .A0 (que_out_25__2__13), .A1 (nx10076), .B0 (
          que_out_16__2__13), .B1 (nx10102)) ;
    aoi22 ix8562 (.Y (nx8561), .A0 (que_out_24__2__13), .A1 (nx10050), .B0 (
          que_out_22__2__13), .B1 (nx10024)) ;
    nand03 ix5135 (.Y (nx5134), .A0 (nx8565), .A1 (nx8567), .A2 (nx8569)) ;
    aoi222 ix8566 (.Y (nx8565), .A0 (que_out_15__2__13), .A1 (nx9972), .B0 (
           que_out_3__2__13), .B1 (nx9998), .C0 (que_out_23__2__13), .C1 (nx9946
           )) ;
    aoi22 ix8568 (.Y (nx8567), .A0 (que_out_27__2__13), .A1 (nx9920), .B0 (
          que_out_4__2__13), .B1 (nx9894)) ;
    aoi22 ix8570 (.Y (nx8569), .A0 (que_out_0__2__13), .A1 (nx9842), .B0 (
          que_out_2__2__13), .B1 (nx9868)) ;
    nand03 ix5109 (.Y (nx5108), .A0 (nx8573), .A1 (nx8575), .A2 (nx8577)) ;
    aoi222 ix8574 (.Y (nx8573), .A0 (que_out_26__2__13), .A1 (nx9816), .B0 (
           que_out_14__2__13), .B1 (nx9790), .C0 (que_out_11__2__13), .C1 (
           nx9764)) ;
    aoi22 ix8576 (.Y (nx8575), .A0 (que_out_13__2__13), .A1 (nx9738), .B0 (
          que_out_7__2__13), .B1 (nx9712)) ;
    aoi22 ix8578 (.Y (nx8577), .A0 (que_out_12__2__13), .A1 (nx9686), .B0 (
          que_out_1__2__13), .B1 (nx9660)) ;
    or04 ix5303 (.Y (out_column_2__14), .A0 (nx5298), .A1 (nx5272), .A2 (nx5244)
         , .A3 (nx5218)) ;
    nand03 ix5299 (.Y (nx5298), .A0 (nx8583), .A1 (nx8585), .A2 (nx8587)) ;
    aoi222 ix8584 (.Y (nx8583), .A0 (que_out_10__2__14), .A1 (nx10310), .B0 (
           que_out_6__2__14), .B1 (nx10362), .C0 (que_out_9__2__14), .C1 (
           nx10336)) ;
    aoi22 ix8586 (.Y (nx8585), .A0 (que_out_5__2__14), .A1 (nx10258), .B0 (
          que_out_18__2__14), .B1 (nx10284)) ;
    aoi22 ix8588 (.Y (nx8587), .A0 (que_out_17__2__14), .A1 (nx10232), .B0 (
          que_out_20__2__14), .B1 (nx10206)) ;
    nand03 ix5273 (.Y (nx5272), .A0 (nx8591), .A1 (nx8593), .A2 (nx8595)) ;
    aoi222 ix8592 (.Y (nx8591), .A0 (que_out_19__2__14), .A1 (nx10180), .B0 (
           que_out_21__2__14), .B1 (nx10154), .C0 (que_out_8__2__14), .C1 (
           nx10128)) ;
    aoi22 ix8594 (.Y (nx8593), .A0 (que_out_25__2__14), .A1 (nx10076), .B0 (
          que_out_16__2__14), .B1 (nx10102)) ;
    aoi22 ix8596 (.Y (nx8595), .A0 (que_out_24__2__14), .A1 (nx10050), .B0 (
          que_out_22__2__14), .B1 (nx10024)) ;
    nand03 ix5245 (.Y (nx5244), .A0 (nx8599), .A1 (nx8601), .A2 (nx8603)) ;
    aoi222 ix8600 (.Y (nx8599), .A0 (que_out_15__2__14), .A1 (nx9972), .B0 (
           que_out_3__2__14), .B1 (nx9998), .C0 (que_out_23__2__14), .C1 (nx9946
           )) ;
    aoi22 ix8602 (.Y (nx8601), .A0 (que_out_27__2__14), .A1 (nx9920), .B0 (
          que_out_4__2__14), .B1 (nx9894)) ;
    aoi22 ix8604 (.Y (nx8603), .A0 (que_out_0__2__14), .A1 (nx9842), .B0 (
          que_out_2__2__14), .B1 (nx9868)) ;
    nand03 ix5219 (.Y (nx5218), .A0 (nx8607), .A1 (nx8609), .A2 (nx8611)) ;
    aoi222 ix8608 (.Y (nx8607), .A0 (que_out_26__2__14), .A1 (nx9816), .B0 (
           que_out_14__2__14), .B1 (nx9790), .C0 (que_out_11__2__14), .C1 (
           nx9764)) ;
    aoi22 ix8610 (.Y (nx8609), .A0 (que_out_13__2__14), .A1 (nx9738), .B0 (
          que_out_7__2__14), .B1 (nx9712)) ;
    aoi22 ix8612 (.Y (nx8611), .A0 (que_out_12__2__14), .A1 (nx9686), .B0 (
          que_out_1__2__14), .B1 (nx9660)) ;
    or04 ix5413 (.Y (out_column_2__15), .A0 (nx5408), .A1 (nx5382), .A2 (nx5354)
         , .A3 (nx5328)) ;
    nand03 ix5409 (.Y (nx5408), .A0 (nx8617), .A1 (nx8619), .A2 (nx8621)) ;
    aoi222 ix8618 (.Y (nx8617), .A0 (que_out_10__2__15), .A1 (nx10310), .B0 (
           que_out_6__2__15), .B1 (nx10362), .C0 (que_out_9__2__15), .C1 (
           nx10336)) ;
    aoi22 ix8620 (.Y (nx8619), .A0 (que_out_5__2__15), .A1 (nx10258), .B0 (
          que_out_18__2__15), .B1 (nx10284)) ;
    aoi22 ix8622 (.Y (nx8621), .A0 (que_out_17__2__15), .A1 (nx10232), .B0 (
          que_out_20__2__15), .B1 (nx10206)) ;
    nand03 ix5383 (.Y (nx5382), .A0 (nx8625), .A1 (nx8627), .A2 (nx8629)) ;
    aoi222 ix8626 (.Y (nx8625), .A0 (que_out_19__2__15), .A1 (nx10180), .B0 (
           que_out_21__2__15), .B1 (nx10154), .C0 (que_out_8__2__15), .C1 (
           nx10128)) ;
    aoi22 ix8628 (.Y (nx8627), .A0 (que_out_25__2__15), .A1 (nx10076), .B0 (
          que_out_16__2__15), .B1 (nx10102)) ;
    aoi22 ix8630 (.Y (nx8629), .A0 (que_out_24__2__15), .A1 (nx10050), .B0 (
          que_out_22__2__15), .B1 (nx10024)) ;
    nand03 ix5355 (.Y (nx5354), .A0 (nx8633), .A1 (nx8635), .A2 (nx8637)) ;
    aoi222 ix8634 (.Y (nx8633), .A0 (que_out_15__2__15), .A1 (nx9972), .B0 (
           que_out_3__2__15), .B1 (nx9998), .C0 (que_out_23__2__15), .C1 (nx9946
           )) ;
    aoi22 ix8636 (.Y (nx8635), .A0 (que_out_27__2__15), .A1 (nx9920), .B0 (
          que_out_4__2__15), .B1 (nx9894)) ;
    aoi22 ix8638 (.Y (nx8637), .A0 (que_out_0__2__15), .A1 (nx9842), .B0 (
          que_out_2__2__15), .B1 (nx9868)) ;
    nand03 ix5329 (.Y (nx5328), .A0 (nx8641), .A1 (nx8643), .A2 (nx8645)) ;
    aoi222 ix8642 (.Y (nx8641), .A0 (que_out_26__2__15), .A1 (nx9816), .B0 (
           que_out_14__2__15), .B1 (nx9790), .C0 (que_out_11__2__15), .C1 (
           nx9764)) ;
    aoi22 ix8644 (.Y (nx8643), .A0 (que_out_13__2__15), .A1 (nx9738), .B0 (
          que_out_7__2__15), .B1 (nx9712)) ;
    aoi22 ix8646 (.Y (nx8645), .A0 (que_out_12__2__15), .A1 (nx9686), .B0 (
          que_out_1__2__15), .B1 (nx9660)) ;
    or04 ix5523 (.Y (out_column_1__0), .A0 (nx5518), .A1 (nx5492), .A2 (nx5464)
         , .A3 (nx5438)) ;
    nand03 ix5519 (.Y (nx5518), .A0 (nx8651), .A1 (nx8653), .A2 (nx8655)) ;
    aoi222 ix8652 (.Y (nx8651), .A0 (que_out_10__1__0), .A1 (nx10310), .B0 (
           que_out_6__1__0), .B1 (nx10362), .C0 (que_out_9__1__0), .C1 (nx10336)
           ) ;
    aoi22 ix8654 (.Y (nx8653), .A0 (que_out_5__1__0), .A1 (nx10258), .B0 (
          que_out_18__1__0), .B1 (nx10284)) ;
    aoi22 ix8656 (.Y (nx8655), .A0 (que_out_17__1__0), .A1 (nx10232), .B0 (
          que_out_20__1__0), .B1 (nx10206)) ;
    nand03 ix5493 (.Y (nx5492), .A0 (nx8659), .A1 (nx8661), .A2 (nx8663)) ;
    aoi222 ix8660 (.Y (nx8659), .A0 (que_out_19__1__0), .A1 (nx10180), .B0 (
           que_out_21__1__0), .B1 (nx10154), .C0 (que_out_8__1__0), .C1 (nx10128
           )) ;
    aoi22 ix8662 (.Y (nx8661), .A0 (que_out_25__1__0), .A1 (nx10076), .B0 (
          que_out_16__1__0), .B1 (nx10102)) ;
    aoi22 ix8664 (.Y (nx8663), .A0 (que_out_24__1__0), .A1 (nx10050), .B0 (
          que_out_22__1__0), .B1 (nx10024)) ;
    nand03 ix5465 (.Y (nx5464), .A0 (nx8667), .A1 (nx8669), .A2 (nx8671)) ;
    aoi222 ix8668 (.Y (nx8667), .A0 (que_out_15__1__0), .A1 (nx9972), .B0 (
           que_out_3__1__0), .B1 (nx9998), .C0 (que_out_23__1__0), .C1 (nx9946)
           ) ;
    aoi22 ix8670 (.Y (nx8669), .A0 (que_out_27__1__0), .A1 (nx9920), .B0 (
          que_out_4__1__0), .B1 (nx9894)) ;
    aoi22 ix8672 (.Y (nx8671), .A0 (que_out_0__1__0), .A1 (nx9842), .B0 (
          que_out_2__1__0), .B1 (nx9868)) ;
    nand03 ix5439 (.Y (nx5438), .A0 (nx8675), .A1 (nx8677), .A2 (nx8679)) ;
    aoi222 ix8676 (.Y (nx8675), .A0 (que_out_26__1__0), .A1 (nx9816), .B0 (
           que_out_14__1__0), .B1 (nx9790), .C0 (que_out_11__1__0), .C1 (nx9764)
           ) ;
    aoi22 ix8678 (.Y (nx8677), .A0 (que_out_13__1__0), .A1 (nx9738), .B0 (
          que_out_7__1__0), .B1 (nx9712)) ;
    aoi22 ix8680 (.Y (nx8679), .A0 (que_out_12__1__0), .A1 (nx9686), .B0 (
          que_out_1__1__0), .B1 (nx9660)) ;
    or04 ix5633 (.Y (out_column_1__1), .A0 (nx5628), .A1 (nx5602), .A2 (nx5574)
         , .A3 (nx5548)) ;
    nand03 ix5629 (.Y (nx5628), .A0 (nx8685), .A1 (nx8687), .A2 (nx8689)) ;
    aoi222 ix8686 (.Y (nx8685), .A0 (que_out_10__1__1), .A1 (nx10312), .B0 (
           que_out_6__1__1), .B1 (nx10364), .C0 (que_out_9__1__1), .C1 (nx10338)
           ) ;
    aoi22 ix8688 (.Y (nx8687), .A0 (que_out_5__1__1), .A1 (nx10260), .B0 (
          que_out_18__1__1), .B1 (nx10286)) ;
    aoi22 ix8690 (.Y (nx8689), .A0 (que_out_17__1__1), .A1 (nx10234), .B0 (
          que_out_20__1__1), .B1 (nx10208)) ;
    nand03 ix5603 (.Y (nx5602), .A0 (nx8693), .A1 (nx8695), .A2 (nx8697)) ;
    aoi222 ix8694 (.Y (nx8693), .A0 (que_out_19__1__1), .A1 (nx10182), .B0 (
           que_out_21__1__1), .B1 (nx10156), .C0 (que_out_8__1__1), .C1 (nx10130
           )) ;
    aoi22 ix8696 (.Y (nx8695), .A0 (que_out_25__1__1), .A1 (nx10078), .B0 (
          que_out_16__1__1), .B1 (nx10104)) ;
    aoi22 ix8698 (.Y (nx8697), .A0 (que_out_24__1__1), .A1 (nx10052), .B0 (
          que_out_22__1__1), .B1 (nx10026)) ;
    nand03 ix5575 (.Y (nx5574), .A0 (nx8701), .A1 (nx8703), .A2 (nx8705)) ;
    aoi222 ix8702 (.Y (nx8701), .A0 (que_out_15__1__1), .A1 (nx9974), .B0 (
           que_out_3__1__1), .B1 (nx10000), .C0 (que_out_23__1__1), .C1 (nx9948)
           ) ;
    aoi22 ix8704 (.Y (nx8703), .A0 (que_out_27__1__1), .A1 (nx9922), .B0 (
          que_out_4__1__1), .B1 (nx9896)) ;
    aoi22 ix8706 (.Y (nx8705), .A0 (que_out_0__1__1), .A1 (nx9844), .B0 (
          que_out_2__1__1), .B1 (nx9870)) ;
    nand03 ix5549 (.Y (nx5548), .A0 (nx8709), .A1 (nx8711), .A2 (nx8713)) ;
    aoi222 ix8710 (.Y (nx8709), .A0 (que_out_26__1__1), .A1 (nx9818), .B0 (
           que_out_14__1__1), .B1 (nx9792), .C0 (que_out_11__1__1), .C1 (nx9766)
           ) ;
    aoi22 ix8712 (.Y (nx8711), .A0 (que_out_13__1__1), .A1 (nx9740), .B0 (
          que_out_7__1__1), .B1 (nx9714)) ;
    aoi22 ix8714 (.Y (nx8713), .A0 (que_out_12__1__1), .A1 (nx9688), .B0 (
          que_out_1__1__1), .B1 (nx9662)) ;
    or04 ix5743 (.Y (out_column_1__2), .A0 (nx5738), .A1 (nx5712), .A2 (nx5684)
         , .A3 (nx5658)) ;
    nand03 ix5739 (.Y (nx5738), .A0 (nx8719), .A1 (nx8721), .A2 (nx8723)) ;
    aoi222 ix8720 (.Y (nx8719), .A0 (que_out_10__1__2), .A1 (nx10312), .B0 (
           que_out_6__1__2), .B1 (nx10364), .C0 (que_out_9__1__2), .C1 (nx10338)
           ) ;
    aoi22 ix8722 (.Y (nx8721), .A0 (que_out_5__1__2), .A1 (nx10260), .B0 (
          que_out_18__1__2), .B1 (nx10286)) ;
    aoi22 ix8724 (.Y (nx8723), .A0 (que_out_17__1__2), .A1 (nx10234), .B0 (
          que_out_20__1__2), .B1 (nx10208)) ;
    nand03 ix5713 (.Y (nx5712), .A0 (nx8727), .A1 (nx8729), .A2 (nx8731)) ;
    aoi222 ix8728 (.Y (nx8727), .A0 (que_out_19__1__2), .A1 (nx10182), .B0 (
           que_out_21__1__2), .B1 (nx10156), .C0 (que_out_8__1__2), .C1 (nx10130
           )) ;
    aoi22 ix8730 (.Y (nx8729), .A0 (que_out_25__1__2), .A1 (nx10078), .B0 (
          que_out_16__1__2), .B1 (nx10104)) ;
    aoi22 ix8732 (.Y (nx8731), .A0 (que_out_24__1__2), .A1 (nx10052), .B0 (
          que_out_22__1__2), .B1 (nx10026)) ;
    nand03 ix5685 (.Y (nx5684), .A0 (nx8735), .A1 (nx8737), .A2 (nx8739)) ;
    aoi222 ix8736 (.Y (nx8735), .A0 (que_out_15__1__2), .A1 (nx9974), .B0 (
           que_out_3__1__2), .B1 (nx10000), .C0 (que_out_23__1__2), .C1 (nx9948)
           ) ;
    aoi22 ix8738 (.Y (nx8737), .A0 (que_out_27__1__2), .A1 (nx9922), .B0 (
          que_out_4__1__2), .B1 (nx9896)) ;
    aoi22 ix8740 (.Y (nx8739), .A0 (que_out_0__1__2), .A1 (nx9844), .B0 (
          que_out_2__1__2), .B1 (nx9870)) ;
    nand03 ix5659 (.Y (nx5658), .A0 (nx8743), .A1 (nx8745), .A2 (nx8747)) ;
    aoi222 ix8744 (.Y (nx8743), .A0 (que_out_26__1__2), .A1 (nx9818), .B0 (
           que_out_14__1__2), .B1 (nx9792), .C0 (que_out_11__1__2), .C1 (nx9766)
           ) ;
    aoi22 ix8746 (.Y (nx8745), .A0 (que_out_13__1__2), .A1 (nx9740), .B0 (
          que_out_7__1__2), .B1 (nx9714)) ;
    aoi22 ix8748 (.Y (nx8747), .A0 (que_out_12__1__2), .A1 (nx9688), .B0 (
          que_out_1__1__2), .B1 (nx9662)) ;
    or04 ix5853 (.Y (out_column_1__3), .A0 (nx5848), .A1 (nx5822), .A2 (nx5794)
         , .A3 (nx5768)) ;
    nand03 ix5849 (.Y (nx5848), .A0 (nx8753), .A1 (nx8755), .A2 (nx8757)) ;
    aoi222 ix8754 (.Y (nx8753), .A0 (que_out_10__1__3), .A1 (nx10312), .B0 (
           que_out_6__1__3), .B1 (nx10364), .C0 (que_out_9__1__3), .C1 (nx10338)
           ) ;
    aoi22 ix8756 (.Y (nx8755), .A0 (que_out_5__1__3), .A1 (nx10260), .B0 (
          que_out_18__1__3), .B1 (nx10286)) ;
    aoi22 ix8758 (.Y (nx8757), .A0 (que_out_17__1__3), .A1 (nx10234), .B0 (
          que_out_20__1__3), .B1 (nx10208)) ;
    nand03 ix5823 (.Y (nx5822), .A0 (nx8761), .A1 (nx8763), .A2 (nx8765)) ;
    aoi222 ix8762 (.Y (nx8761), .A0 (que_out_19__1__3), .A1 (nx10182), .B0 (
           que_out_21__1__3), .B1 (nx10156), .C0 (que_out_8__1__3), .C1 (nx10130
           )) ;
    aoi22 ix8764 (.Y (nx8763), .A0 (que_out_25__1__3), .A1 (nx10078), .B0 (
          que_out_16__1__3), .B1 (nx10104)) ;
    aoi22 ix8766 (.Y (nx8765), .A0 (que_out_24__1__3), .A1 (nx10052), .B0 (
          que_out_22__1__3), .B1 (nx10026)) ;
    nand03 ix5795 (.Y (nx5794), .A0 (nx8769), .A1 (nx8771), .A2 (nx8773)) ;
    aoi222 ix8770 (.Y (nx8769), .A0 (que_out_15__1__3), .A1 (nx9974), .B0 (
           que_out_3__1__3), .B1 (nx10000), .C0 (que_out_23__1__3), .C1 (nx9948)
           ) ;
    aoi22 ix8772 (.Y (nx8771), .A0 (que_out_27__1__3), .A1 (nx9922), .B0 (
          que_out_4__1__3), .B1 (nx9896)) ;
    aoi22 ix8774 (.Y (nx8773), .A0 (que_out_0__1__3), .A1 (nx9844), .B0 (
          que_out_2__1__3), .B1 (nx9870)) ;
    nand03 ix5769 (.Y (nx5768), .A0 (nx8777), .A1 (nx8779), .A2 (nx8781)) ;
    aoi222 ix8778 (.Y (nx8777), .A0 (que_out_26__1__3), .A1 (nx9818), .B0 (
           que_out_14__1__3), .B1 (nx9792), .C0 (que_out_11__1__3), .C1 (nx9766)
           ) ;
    aoi22 ix8780 (.Y (nx8779), .A0 (que_out_13__1__3), .A1 (nx9740), .B0 (
          que_out_7__1__3), .B1 (nx9714)) ;
    aoi22 ix8782 (.Y (nx8781), .A0 (que_out_12__1__3), .A1 (nx9688), .B0 (
          que_out_1__1__3), .B1 (nx9662)) ;
    or04 ix5963 (.Y (out_column_1__4), .A0 (nx5958), .A1 (nx5932), .A2 (nx5904)
         , .A3 (nx5878)) ;
    nand03 ix5959 (.Y (nx5958), .A0 (nx8787), .A1 (nx8789), .A2 (nx8791)) ;
    aoi222 ix8788 (.Y (nx8787), .A0 (que_out_10__1__4), .A1 (nx10312), .B0 (
           que_out_6__1__4), .B1 (nx10364), .C0 (que_out_9__1__4), .C1 (nx10338)
           ) ;
    aoi22 ix8790 (.Y (nx8789), .A0 (que_out_5__1__4), .A1 (nx10260), .B0 (
          que_out_18__1__4), .B1 (nx10286)) ;
    aoi22 ix8792 (.Y (nx8791), .A0 (que_out_17__1__4), .A1 (nx10234), .B0 (
          que_out_20__1__4), .B1 (nx10208)) ;
    nand03 ix5933 (.Y (nx5932), .A0 (nx8795), .A1 (nx8797), .A2 (nx8799)) ;
    aoi222 ix8796 (.Y (nx8795), .A0 (que_out_19__1__4), .A1 (nx10182), .B0 (
           que_out_21__1__4), .B1 (nx10156), .C0 (que_out_8__1__4), .C1 (nx10130
           )) ;
    aoi22 ix8798 (.Y (nx8797), .A0 (que_out_25__1__4), .A1 (nx10078), .B0 (
          que_out_16__1__4), .B1 (nx10104)) ;
    aoi22 ix8800 (.Y (nx8799), .A0 (que_out_24__1__4), .A1 (nx10052), .B0 (
          que_out_22__1__4), .B1 (nx10026)) ;
    nand03 ix5905 (.Y (nx5904), .A0 (nx8803), .A1 (nx8805), .A2 (nx8807)) ;
    aoi222 ix8804 (.Y (nx8803), .A0 (que_out_15__1__4), .A1 (nx9974), .B0 (
           que_out_3__1__4), .B1 (nx10000), .C0 (que_out_23__1__4), .C1 (nx9948)
           ) ;
    aoi22 ix8806 (.Y (nx8805), .A0 (que_out_27__1__4), .A1 (nx9922), .B0 (
          que_out_4__1__4), .B1 (nx9896)) ;
    aoi22 ix8808 (.Y (nx8807), .A0 (que_out_0__1__4), .A1 (nx9844), .B0 (
          que_out_2__1__4), .B1 (nx9870)) ;
    nand03 ix5879 (.Y (nx5878), .A0 (nx8811), .A1 (nx8813), .A2 (nx8815)) ;
    aoi222 ix8812 (.Y (nx8811), .A0 (que_out_26__1__4), .A1 (nx9818), .B0 (
           que_out_14__1__4), .B1 (nx9792), .C0 (que_out_11__1__4), .C1 (nx9766)
           ) ;
    aoi22 ix8814 (.Y (nx8813), .A0 (que_out_13__1__4), .A1 (nx9740), .B0 (
          que_out_7__1__4), .B1 (nx9714)) ;
    aoi22 ix8816 (.Y (nx8815), .A0 (que_out_12__1__4), .A1 (nx9688), .B0 (
          que_out_1__1__4), .B1 (nx9662)) ;
    or04 ix6073 (.Y (out_column_1__5), .A0 (nx6068), .A1 (nx6042), .A2 (nx6014)
         , .A3 (nx5988)) ;
    nand03 ix6069 (.Y (nx6068), .A0 (nx8821), .A1 (nx8823), .A2 (nx8825)) ;
    aoi222 ix8822 (.Y (nx8821), .A0 (que_out_10__1__5), .A1 (nx10312), .B0 (
           que_out_6__1__5), .B1 (nx10364), .C0 (que_out_9__1__5), .C1 (nx10338)
           ) ;
    aoi22 ix8824 (.Y (nx8823), .A0 (que_out_5__1__5), .A1 (nx10260), .B0 (
          que_out_18__1__5), .B1 (nx10286)) ;
    aoi22 ix8826 (.Y (nx8825), .A0 (que_out_17__1__5), .A1 (nx10234), .B0 (
          que_out_20__1__5), .B1 (nx10208)) ;
    nand03 ix6043 (.Y (nx6042), .A0 (nx8829), .A1 (nx8831), .A2 (nx8833)) ;
    aoi222 ix8830 (.Y (nx8829), .A0 (que_out_19__1__5), .A1 (nx10182), .B0 (
           que_out_21__1__5), .B1 (nx10156), .C0 (que_out_8__1__5), .C1 (nx10130
           )) ;
    aoi22 ix8832 (.Y (nx8831), .A0 (que_out_25__1__5), .A1 (nx10078), .B0 (
          que_out_16__1__5), .B1 (nx10104)) ;
    aoi22 ix8834 (.Y (nx8833), .A0 (que_out_24__1__5), .A1 (nx10052), .B0 (
          que_out_22__1__5), .B1 (nx10026)) ;
    nand03 ix6015 (.Y (nx6014), .A0 (nx8837), .A1 (nx8839), .A2 (nx8841)) ;
    aoi222 ix8838 (.Y (nx8837), .A0 (que_out_15__1__5), .A1 (nx9974), .B0 (
           que_out_3__1__5), .B1 (nx10000), .C0 (que_out_23__1__5), .C1 (nx9948)
           ) ;
    aoi22 ix8840 (.Y (nx8839), .A0 (que_out_27__1__5), .A1 (nx9922), .B0 (
          que_out_4__1__5), .B1 (nx9896)) ;
    aoi22 ix8842 (.Y (nx8841), .A0 (que_out_0__1__5), .A1 (nx9844), .B0 (
          que_out_2__1__5), .B1 (nx9870)) ;
    nand03 ix5989 (.Y (nx5988), .A0 (nx8845), .A1 (nx8847), .A2 (nx8849)) ;
    aoi222 ix8846 (.Y (nx8845), .A0 (que_out_26__1__5), .A1 (nx9818), .B0 (
           que_out_14__1__5), .B1 (nx9792), .C0 (que_out_11__1__5), .C1 (nx9766)
           ) ;
    aoi22 ix8848 (.Y (nx8847), .A0 (que_out_13__1__5), .A1 (nx9740), .B0 (
          que_out_7__1__5), .B1 (nx9714)) ;
    aoi22 ix8850 (.Y (nx8849), .A0 (que_out_12__1__5), .A1 (nx9688), .B0 (
          que_out_1__1__5), .B1 (nx9662)) ;
    or04 ix6183 (.Y (out_column_1__6), .A0 (nx6178), .A1 (nx6152), .A2 (nx6124)
         , .A3 (nx6098)) ;
    nand03 ix6179 (.Y (nx6178), .A0 (nx8855), .A1 (nx8857), .A2 (nx8859)) ;
    aoi222 ix8856 (.Y (nx8855), .A0 (que_out_10__1__6), .A1 (nx10312), .B0 (
           que_out_6__1__6), .B1 (nx10364), .C0 (que_out_9__1__6), .C1 (nx10338)
           ) ;
    aoi22 ix8858 (.Y (nx8857), .A0 (que_out_5__1__6), .A1 (nx10260), .B0 (
          que_out_18__1__6), .B1 (nx10286)) ;
    aoi22 ix8860 (.Y (nx8859), .A0 (que_out_17__1__6), .A1 (nx10234), .B0 (
          que_out_20__1__6), .B1 (nx10208)) ;
    nand03 ix6153 (.Y (nx6152), .A0 (nx8863), .A1 (nx8865), .A2 (nx8867)) ;
    aoi222 ix8864 (.Y (nx8863), .A0 (que_out_19__1__6), .A1 (nx10182), .B0 (
           que_out_21__1__6), .B1 (nx10156), .C0 (que_out_8__1__6), .C1 (nx10130
           )) ;
    aoi22 ix8866 (.Y (nx8865), .A0 (que_out_25__1__6), .A1 (nx10078), .B0 (
          que_out_16__1__6), .B1 (nx10104)) ;
    aoi22 ix8868 (.Y (nx8867), .A0 (que_out_24__1__6), .A1 (nx10052), .B0 (
          que_out_22__1__6), .B1 (nx10026)) ;
    nand03 ix6125 (.Y (nx6124), .A0 (nx8871), .A1 (nx8873), .A2 (nx8875)) ;
    aoi222 ix8872 (.Y (nx8871), .A0 (que_out_15__1__6), .A1 (nx9974), .B0 (
           que_out_3__1__6), .B1 (nx10000), .C0 (que_out_23__1__6), .C1 (nx9948)
           ) ;
    aoi22 ix8874 (.Y (nx8873), .A0 (que_out_27__1__6), .A1 (nx9922), .B0 (
          que_out_4__1__6), .B1 (nx9896)) ;
    aoi22 ix8876 (.Y (nx8875), .A0 (que_out_0__1__6), .A1 (nx9844), .B0 (
          que_out_2__1__6), .B1 (nx9870)) ;
    nand03 ix6099 (.Y (nx6098), .A0 (nx8879), .A1 (nx8881), .A2 (nx8883)) ;
    aoi222 ix8880 (.Y (nx8879), .A0 (que_out_26__1__6), .A1 (nx9818), .B0 (
           que_out_14__1__6), .B1 (nx9792), .C0 (que_out_11__1__6), .C1 (nx9766)
           ) ;
    aoi22 ix8882 (.Y (nx8881), .A0 (que_out_13__1__6), .A1 (nx9740), .B0 (
          que_out_7__1__6), .B1 (nx9714)) ;
    aoi22 ix8884 (.Y (nx8883), .A0 (que_out_12__1__6), .A1 (nx9688), .B0 (
          que_out_1__1__6), .B1 (nx9662)) ;
    or04 ix6293 (.Y (out_column_1__7), .A0 (nx6288), .A1 (nx6262), .A2 (nx6234)
         , .A3 (nx6208)) ;
    nand03 ix6289 (.Y (nx6288), .A0 (nx8889), .A1 (nx8891), .A2 (nx8893)) ;
    aoi222 ix8890 (.Y (nx8889), .A0 (que_out_10__1__7), .A1 (nx10312), .B0 (
           que_out_6__1__7), .B1 (nx10364), .C0 (que_out_9__1__7), .C1 (nx10338)
           ) ;
    aoi22 ix8892 (.Y (nx8891), .A0 (que_out_5__1__7), .A1 (nx10260), .B0 (
          que_out_18__1__7), .B1 (nx10286)) ;
    aoi22 ix8894 (.Y (nx8893), .A0 (que_out_17__1__7), .A1 (nx10234), .B0 (
          que_out_20__1__7), .B1 (nx10208)) ;
    nand03 ix6263 (.Y (nx6262), .A0 (nx8897), .A1 (nx8899), .A2 (nx8901)) ;
    aoi222 ix8898 (.Y (nx8897), .A0 (que_out_19__1__7), .A1 (nx10182), .B0 (
           que_out_21__1__7), .B1 (nx10156), .C0 (que_out_8__1__7), .C1 (nx10130
           )) ;
    aoi22 ix8900 (.Y (nx8899), .A0 (que_out_25__1__7), .A1 (nx10078), .B0 (
          que_out_16__1__7), .B1 (nx10104)) ;
    aoi22 ix8902 (.Y (nx8901), .A0 (que_out_24__1__7), .A1 (nx10052), .B0 (
          que_out_22__1__7), .B1 (nx10026)) ;
    nand03 ix6235 (.Y (nx6234), .A0 (nx8905), .A1 (nx8907), .A2 (nx8909)) ;
    aoi222 ix8906 (.Y (nx8905), .A0 (que_out_15__1__7), .A1 (nx9974), .B0 (
           que_out_3__1__7), .B1 (nx10000), .C0 (que_out_23__1__7), .C1 (nx9948)
           ) ;
    aoi22 ix8908 (.Y (nx8907), .A0 (que_out_27__1__7), .A1 (nx9922), .B0 (
          que_out_4__1__7), .B1 (nx9896)) ;
    aoi22 ix8910 (.Y (nx8909), .A0 (que_out_0__1__7), .A1 (nx9844), .B0 (
          que_out_2__1__7), .B1 (nx9870)) ;
    nand03 ix6209 (.Y (nx6208), .A0 (nx8913), .A1 (nx8915), .A2 (nx8917)) ;
    aoi222 ix8914 (.Y (nx8913), .A0 (que_out_26__1__7), .A1 (nx9818), .B0 (
           que_out_14__1__7), .B1 (nx9792), .C0 (que_out_11__1__7), .C1 (nx9766)
           ) ;
    aoi22 ix8916 (.Y (nx8915), .A0 (que_out_13__1__7), .A1 (nx9740), .B0 (
          que_out_7__1__7), .B1 (nx9714)) ;
    aoi22 ix8918 (.Y (nx8917), .A0 (que_out_12__1__7), .A1 (nx9688), .B0 (
          que_out_1__1__7), .B1 (nx9662)) ;
    or04 ix6403 (.Y (out_column_1__8), .A0 (nx6398), .A1 (nx6372), .A2 (nx6344)
         , .A3 (nx6318)) ;
    nand03 ix6399 (.Y (nx6398), .A0 (nx8923), .A1 (nx8925), .A2 (nx8927)) ;
    aoi222 ix8924 (.Y (nx8923), .A0 (que_out_10__1__8), .A1 (nx10314), .B0 (
           que_out_6__1__8), .B1 (nx10366), .C0 (que_out_9__1__8), .C1 (nx10340)
           ) ;
    aoi22 ix8926 (.Y (nx8925), .A0 (que_out_5__1__8), .A1 (nx10262), .B0 (
          que_out_18__1__8), .B1 (nx10288)) ;
    aoi22 ix8928 (.Y (nx8927), .A0 (que_out_17__1__8), .A1 (nx10236), .B0 (
          que_out_20__1__8), .B1 (nx10210)) ;
    nand03 ix6373 (.Y (nx6372), .A0 (nx8931), .A1 (nx8933), .A2 (nx8935)) ;
    aoi222 ix8932 (.Y (nx8931), .A0 (que_out_19__1__8), .A1 (nx10184), .B0 (
           que_out_21__1__8), .B1 (nx10158), .C0 (que_out_8__1__8), .C1 (nx10132
           )) ;
    aoi22 ix8934 (.Y (nx8933), .A0 (que_out_25__1__8), .A1 (nx10080), .B0 (
          que_out_16__1__8), .B1 (nx10106)) ;
    aoi22 ix8936 (.Y (nx8935), .A0 (que_out_24__1__8), .A1 (nx10054), .B0 (
          que_out_22__1__8), .B1 (nx10028)) ;
    nand03 ix6345 (.Y (nx6344), .A0 (nx8939), .A1 (nx8941), .A2 (nx8943)) ;
    aoi222 ix8940 (.Y (nx8939), .A0 (que_out_15__1__8), .A1 (nx9976), .B0 (
           que_out_3__1__8), .B1 (nx10002), .C0 (que_out_23__1__8), .C1 (nx9950)
           ) ;
    aoi22 ix8942 (.Y (nx8941), .A0 (que_out_27__1__8), .A1 (nx9924), .B0 (
          que_out_4__1__8), .B1 (nx9898)) ;
    aoi22 ix8944 (.Y (nx8943), .A0 (que_out_0__1__8), .A1 (nx9846), .B0 (
          que_out_2__1__8), .B1 (nx9872)) ;
    nand03 ix6319 (.Y (nx6318), .A0 (nx8947), .A1 (nx8949), .A2 (nx8951)) ;
    aoi222 ix8948 (.Y (nx8947), .A0 (que_out_26__1__8), .A1 (nx9820), .B0 (
           que_out_14__1__8), .B1 (nx9794), .C0 (que_out_11__1__8), .C1 (nx9768)
           ) ;
    aoi22 ix8950 (.Y (nx8949), .A0 (que_out_13__1__8), .A1 (nx9742), .B0 (
          que_out_7__1__8), .B1 (nx9716)) ;
    aoi22 ix8952 (.Y (nx8951), .A0 (que_out_12__1__8), .A1 (nx9690), .B0 (
          que_out_1__1__8), .B1 (nx9664)) ;
    or04 ix6513 (.Y (out_column_1__9), .A0 (nx6508), .A1 (nx6482), .A2 (nx6454)
         , .A3 (nx6428)) ;
    nand03 ix6509 (.Y (nx6508), .A0 (nx8955), .A1 (nx8957), .A2 (nx8959)) ;
    aoi222 ix8956 (.Y (nx8955), .A0 (que_out_10__1__9), .A1 (nx10314), .B0 (
           que_out_6__1__9), .B1 (nx10366), .C0 (que_out_9__1__9), .C1 (nx10340)
           ) ;
    aoi22 ix8958 (.Y (nx8957), .A0 (que_out_5__1__9), .A1 (nx10262), .B0 (
          que_out_18__1__9), .B1 (nx10288)) ;
    aoi22 ix8960 (.Y (nx8959), .A0 (que_out_17__1__9), .A1 (nx10236), .B0 (
          que_out_20__1__9), .B1 (nx10210)) ;
    nand03 ix6483 (.Y (nx6482), .A0 (nx8963), .A1 (nx8965), .A2 (nx8967)) ;
    aoi222 ix8964 (.Y (nx8963), .A0 (que_out_19__1__9), .A1 (nx10184), .B0 (
           que_out_21__1__9), .B1 (nx10158), .C0 (que_out_8__1__9), .C1 (nx10132
           )) ;
    aoi22 ix8966 (.Y (nx8965), .A0 (que_out_25__1__9), .A1 (nx10080), .B0 (
          que_out_16__1__9), .B1 (nx10106)) ;
    aoi22 ix8968 (.Y (nx8967), .A0 (que_out_24__1__9), .A1 (nx10054), .B0 (
          que_out_22__1__9), .B1 (nx10028)) ;
    nand03 ix6455 (.Y (nx6454), .A0 (nx8970), .A1 (nx8973), .A2 (nx8975)) ;
    aoi222 ix8972 (.Y (nx8970), .A0 (que_out_15__1__9), .A1 (nx9976), .B0 (
           que_out_3__1__9), .B1 (nx10002), .C0 (que_out_23__1__9), .C1 (nx9950)
           ) ;
    aoi22 ix8974 (.Y (nx8973), .A0 (que_out_27__1__9), .A1 (nx9924), .B0 (
          que_out_4__1__9), .B1 (nx9898)) ;
    aoi22 ix8976 (.Y (nx8975), .A0 (que_out_0__1__9), .A1 (nx9846), .B0 (
          que_out_2__1__9), .B1 (nx9872)) ;
    nand03 ix6429 (.Y (nx6428), .A0 (nx8978), .A1 (nx8981), .A2 (nx8983)) ;
    aoi222 ix8980 (.Y (nx8978), .A0 (que_out_26__1__9), .A1 (nx9820), .B0 (
           que_out_14__1__9), .B1 (nx9794), .C0 (que_out_11__1__9), .C1 (nx9768)
           ) ;
    aoi22 ix8982 (.Y (nx8981), .A0 (que_out_13__1__9), .A1 (nx9742), .B0 (
          que_out_7__1__9), .B1 (nx9716)) ;
    aoi22 ix8984 (.Y (nx8983), .A0 (que_out_12__1__9), .A1 (nx9690), .B0 (
          que_out_1__1__9), .B1 (nx9664)) ;
    or04 ix6623 (.Y (out_column_1__10), .A0 (nx6618), .A1 (nx6592), .A2 (nx6564)
         , .A3 (nx6538)) ;
    nand03 ix6619 (.Y (nx6618), .A0 (nx8989), .A1 (nx8991), .A2 (nx8993)) ;
    aoi222 ix8990 (.Y (nx8989), .A0 (que_out_10__1__10), .A1 (nx10314), .B0 (
           que_out_6__1__10), .B1 (nx10366), .C0 (que_out_9__1__10), .C1 (
           nx10340)) ;
    aoi22 ix8992 (.Y (nx8991), .A0 (que_out_5__1__10), .A1 (nx10262), .B0 (
          que_out_18__1__10), .B1 (nx10288)) ;
    aoi22 ix8994 (.Y (nx8993), .A0 (que_out_17__1__10), .A1 (nx10236), .B0 (
          que_out_20__1__10), .B1 (nx10210)) ;
    nand03 ix6593 (.Y (nx6592), .A0 (nx8997), .A1 (nx8999), .A2 (nx9001)) ;
    aoi222 ix8998 (.Y (nx8997), .A0 (que_out_19__1__10), .A1 (nx10184), .B0 (
           que_out_21__1__10), .B1 (nx10158), .C0 (que_out_8__1__10), .C1 (
           nx10132)) ;
    aoi22 ix9000 (.Y (nx8999), .A0 (que_out_25__1__10), .A1 (nx10080), .B0 (
          que_out_16__1__10), .B1 (nx10106)) ;
    aoi22 ix9002 (.Y (nx9001), .A0 (que_out_24__1__10), .A1 (nx10054), .B0 (
          que_out_22__1__10), .B1 (nx10028)) ;
    nand03 ix6565 (.Y (nx6564), .A0 (nx9005), .A1 (nx9007), .A2 (nx9009)) ;
    aoi222 ix9006 (.Y (nx9005), .A0 (que_out_15__1__10), .A1 (nx9976), .B0 (
           que_out_3__1__10), .B1 (nx10002), .C0 (que_out_23__1__10), .C1 (
           nx9950)) ;
    aoi22 ix9008 (.Y (nx9007), .A0 (que_out_27__1__10), .A1 (nx9924), .B0 (
          que_out_4__1__10), .B1 (nx9898)) ;
    aoi22 ix9010 (.Y (nx9009), .A0 (que_out_0__1__10), .A1 (nx9846), .B0 (
          que_out_2__1__10), .B1 (nx9872)) ;
    nand03 ix6539 (.Y (nx6538), .A0 (nx9013), .A1 (nx9015), .A2 (nx9017)) ;
    aoi222 ix9014 (.Y (nx9013), .A0 (que_out_26__1__10), .A1 (nx9820), .B0 (
           que_out_14__1__10), .B1 (nx9794), .C0 (que_out_11__1__10), .C1 (
           nx9768)) ;
    aoi22 ix9016 (.Y (nx9015), .A0 (que_out_13__1__10), .A1 (nx9742), .B0 (
          que_out_7__1__10), .B1 (nx9716)) ;
    aoi22 ix9018 (.Y (nx9017), .A0 (que_out_12__1__10), .A1 (nx9690), .B0 (
          que_out_1__1__10), .B1 (nx9664)) ;
    or04 ix6733 (.Y (out_column_1__11), .A0 (nx6728), .A1 (nx6702), .A2 (nx6674)
         , .A3 (nx6648)) ;
    nand03 ix6729 (.Y (nx6728), .A0 (nx9023), .A1 (nx9025), .A2 (nx9027)) ;
    aoi222 ix9024 (.Y (nx9023), .A0 (que_out_10__1__11), .A1 (nx10314), .B0 (
           que_out_6__1__11), .B1 (nx10366), .C0 (que_out_9__1__11), .C1 (
           nx10340)) ;
    aoi22 ix9026 (.Y (nx9025), .A0 (que_out_5__1__11), .A1 (nx10262), .B0 (
          que_out_18__1__11), .B1 (nx10288)) ;
    aoi22 ix9028 (.Y (nx9027), .A0 (que_out_17__1__11), .A1 (nx10236), .B0 (
          que_out_20__1__11), .B1 (nx10210)) ;
    nand03 ix6703 (.Y (nx6702), .A0 (nx9031), .A1 (nx9033), .A2 (nx9035)) ;
    aoi222 ix9032 (.Y (nx9031), .A0 (que_out_19__1__11), .A1 (nx10184), .B0 (
           que_out_21__1__11), .B1 (nx10158), .C0 (que_out_8__1__11), .C1 (
           nx10132)) ;
    aoi22 ix9034 (.Y (nx9033), .A0 (que_out_25__1__11), .A1 (nx10080), .B0 (
          que_out_16__1__11), .B1 (nx10106)) ;
    aoi22 ix9036 (.Y (nx9035), .A0 (que_out_24__1__11), .A1 (nx10054), .B0 (
          que_out_22__1__11), .B1 (nx10028)) ;
    nand03 ix6675 (.Y (nx6674), .A0 (nx9039), .A1 (nx9041), .A2 (nx9043)) ;
    aoi222 ix9040 (.Y (nx9039), .A0 (que_out_15__1__11), .A1 (nx9976), .B0 (
           que_out_3__1__11), .B1 (nx10002), .C0 (que_out_23__1__11), .C1 (
           nx9950)) ;
    aoi22 ix9042 (.Y (nx9041), .A0 (que_out_27__1__11), .A1 (nx9924), .B0 (
          que_out_4__1__11), .B1 (nx9898)) ;
    aoi22 ix9044 (.Y (nx9043), .A0 (que_out_0__1__11), .A1 (nx9846), .B0 (
          que_out_2__1__11), .B1 (nx9872)) ;
    nand03 ix6649 (.Y (nx6648), .A0 (nx9047), .A1 (nx9049), .A2 (nx9051)) ;
    aoi222 ix9048 (.Y (nx9047), .A0 (que_out_26__1__11), .A1 (nx9820), .B0 (
           que_out_14__1__11), .B1 (nx9794), .C0 (que_out_11__1__11), .C1 (
           nx9768)) ;
    aoi22 ix9050 (.Y (nx9049), .A0 (que_out_13__1__11), .A1 (nx9742), .B0 (
          que_out_7__1__11), .B1 (nx9716)) ;
    aoi22 ix9052 (.Y (nx9051), .A0 (que_out_12__1__11), .A1 (nx9690), .B0 (
          que_out_1__1__11), .B1 (nx9664)) ;
    or04 ix6843 (.Y (out_column_1__12), .A0 (nx6838), .A1 (nx6812), .A2 (nx6784)
         , .A3 (nx6758)) ;
    nand03 ix6839 (.Y (nx6838), .A0 (nx9057), .A1 (nx9059), .A2 (nx9061)) ;
    aoi222 ix9058 (.Y (nx9057), .A0 (que_out_10__1__12), .A1 (nx10314), .B0 (
           que_out_6__1__12), .B1 (nx10366), .C0 (que_out_9__1__12), .C1 (
           nx10340)) ;
    aoi22 ix9060 (.Y (nx9059), .A0 (que_out_5__1__12), .A1 (nx10262), .B0 (
          que_out_18__1__12), .B1 (nx10288)) ;
    aoi22 ix9062 (.Y (nx9061), .A0 (que_out_17__1__12), .A1 (nx10236), .B0 (
          que_out_20__1__12), .B1 (nx10210)) ;
    nand03 ix6813 (.Y (nx6812), .A0 (nx9065), .A1 (nx9067), .A2 (nx9069)) ;
    aoi222 ix9066 (.Y (nx9065), .A0 (que_out_19__1__12), .A1 (nx10184), .B0 (
           que_out_21__1__12), .B1 (nx10158), .C0 (que_out_8__1__12), .C1 (
           nx10132)) ;
    aoi22 ix9068 (.Y (nx9067), .A0 (que_out_25__1__12), .A1 (nx10080), .B0 (
          que_out_16__1__12), .B1 (nx10106)) ;
    aoi22 ix9070 (.Y (nx9069), .A0 (que_out_24__1__12), .A1 (nx10054), .B0 (
          que_out_22__1__12), .B1 (nx10028)) ;
    nand03 ix6785 (.Y (nx6784), .A0 (nx9073), .A1 (nx9075), .A2 (nx9077)) ;
    aoi222 ix9074 (.Y (nx9073), .A0 (que_out_15__1__12), .A1 (nx9976), .B0 (
           que_out_3__1__12), .B1 (nx10002), .C0 (que_out_23__1__12), .C1 (
           nx9950)) ;
    aoi22 ix9076 (.Y (nx9075), .A0 (que_out_27__1__12), .A1 (nx9924), .B0 (
          que_out_4__1__12), .B1 (nx9898)) ;
    aoi22 ix9078 (.Y (nx9077), .A0 (que_out_0__1__12), .A1 (nx9846), .B0 (
          que_out_2__1__12), .B1 (nx9872)) ;
    nand03 ix6759 (.Y (nx6758), .A0 (nx9081), .A1 (nx9083), .A2 (nx9085)) ;
    aoi222 ix9082 (.Y (nx9081), .A0 (que_out_26__1__12), .A1 (nx9820), .B0 (
           que_out_14__1__12), .B1 (nx9794), .C0 (que_out_11__1__12), .C1 (
           nx9768)) ;
    aoi22 ix9084 (.Y (nx9083), .A0 (que_out_13__1__12), .A1 (nx9742), .B0 (
          que_out_7__1__12), .B1 (nx9716)) ;
    aoi22 ix9086 (.Y (nx9085), .A0 (que_out_12__1__12), .A1 (nx9690), .B0 (
          que_out_1__1__12), .B1 (nx9664)) ;
    or04 ix6953 (.Y (out_column_1__13), .A0 (nx6948), .A1 (nx6922), .A2 (nx6894)
         , .A3 (nx6868)) ;
    nand03 ix6949 (.Y (nx6948), .A0 (nx9090), .A1 (nx9093), .A2 (nx9095)) ;
    aoi222 ix9092 (.Y (nx9090), .A0 (que_out_10__1__13), .A1 (nx10314), .B0 (
           que_out_6__1__13), .B1 (nx10366), .C0 (que_out_9__1__13), .C1 (
           nx10340)) ;
    aoi22 ix9094 (.Y (nx9093), .A0 (que_out_5__1__13), .A1 (nx10262), .B0 (
          que_out_18__1__13), .B1 (nx10288)) ;
    aoi22 ix9096 (.Y (nx9095), .A0 (que_out_17__1__13), .A1 (nx10236), .B0 (
          que_out_20__1__13), .B1 (nx10210)) ;
    nand03 ix6923 (.Y (nx6922), .A0 (nx9098), .A1 (nx9101), .A2 (nx9103)) ;
    aoi222 ix9100 (.Y (nx9098), .A0 (que_out_19__1__13), .A1 (nx10184), .B0 (
           que_out_21__1__13), .B1 (nx10158), .C0 (que_out_8__1__13), .C1 (
           nx10132)) ;
    aoi22 ix9102 (.Y (nx9101), .A0 (que_out_25__1__13), .A1 (nx10080), .B0 (
          que_out_16__1__13), .B1 (nx10106)) ;
    aoi22 ix9104 (.Y (nx9103), .A0 (que_out_24__1__13), .A1 (nx10054), .B0 (
          que_out_22__1__13), .B1 (nx10028)) ;
    nand03 ix6895 (.Y (nx6894), .A0 (nx9106), .A1 (nx9108), .A2 (nx9110)) ;
    aoi222 ix9107 (.Y (nx9106), .A0 (que_out_15__1__13), .A1 (nx9976), .B0 (
           que_out_3__1__13), .B1 (nx10002), .C0 (que_out_23__1__13), .C1 (
           nx9950)) ;
    aoi22 ix9109 (.Y (nx9108), .A0 (que_out_27__1__13), .A1 (nx9924), .B0 (
          que_out_4__1__13), .B1 (nx9898)) ;
    aoi22 ix9111 (.Y (nx9110), .A0 (que_out_0__1__13), .A1 (nx9846), .B0 (
          que_out_2__1__13), .B1 (nx9872)) ;
    nand03 ix6869 (.Y (nx6868), .A0 (nx9113), .A1 (nx9115), .A2 (nx9117)) ;
    aoi222 ix9114 (.Y (nx9113), .A0 (que_out_26__1__13), .A1 (nx9820), .B0 (
           que_out_14__1__13), .B1 (nx9794), .C0 (que_out_11__1__13), .C1 (
           nx9768)) ;
    aoi22 ix9116 (.Y (nx9115), .A0 (que_out_13__1__13), .A1 (nx9742), .B0 (
          que_out_7__1__13), .B1 (nx9716)) ;
    aoi22 ix9118 (.Y (nx9117), .A0 (que_out_12__1__13), .A1 (nx9690), .B0 (
          que_out_1__1__13), .B1 (nx9664)) ;
    or04 ix7063 (.Y (out_column_1__14), .A0 (nx7058), .A1 (nx7032), .A2 (nx7004)
         , .A3 (nx6978)) ;
    nand03 ix7059 (.Y (nx7058), .A0 (nx9121), .A1 (nx9123), .A2 (nx9125)) ;
    aoi222 ix9122 (.Y (nx9121), .A0 (que_out_10__1__14), .A1 (nx10314), .B0 (
           que_out_6__1__14), .B1 (nx10366), .C0 (que_out_9__1__14), .C1 (
           nx10340)) ;
    aoi22 ix9124 (.Y (nx9123), .A0 (que_out_5__1__14), .A1 (nx10262), .B0 (
          que_out_18__1__14), .B1 (nx10288)) ;
    aoi22 ix9126 (.Y (nx9125), .A0 (que_out_17__1__14), .A1 (nx10236), .B0 (
          que_out_20__1__14), .B1 (nx10210)) ;
    nand03 ix7033 (.Y (nx7032), .A0 (nx9128), .A1 (nx9130), .A2 (nx9132)) ;
    aoi222 ix9129 (.Y (nx9128), .A0 (que_out_19__1__14), .A1 (nx10184), .B0 (
           que_out_21__1__14), .B1 (nx10158), .C0 (que_out_8__1__14), .C1 (
           nx10132)) ;
    aoi22 ix9131 (.Y (nx9130), .A0 (que_out_25__1__14), .A1 (nx10080), .B0 (
          que_out_16__1__14), .B1 (nx10106)) ;
    aoi22 ix9133 (.Y (nx9132), .A0 (que_out_24__1__14), .A1 (nx10054), .B0 (
          que_out_22__1__14), .B1 (nx10028)) ;
    nand03 ix7005 (.Y (nx7004), .A0 (nx9135), .A1 (nx9137), .A2 (nx9139)) ;
    aoi222 ix9136 (.Y (nx9135), .A0 (que_out_15__1__14), .A1 (nx9976), .B0 (
           que_out_3__1__14), .B1 (nx10002), .C0 (que_out_23__1__14), .C1 (
           nx9950)) ;
    aoi22 ix9138 (.Y (nx9137), .A0 (que_out_27__1__14), .A1 (nx9924), .B0 (
          que_out_4__1__14), .B1 (nx9898)) ;
    aoi22 ix9140 (.Y (nx9139), .A0 (que_out_0__1__14), .A1 (nx9846), .B0 (
          que_out_2__1__14), .B1 (nx9872)) ;
    nand03 ix6979 (.Y (nx6978), .A0 (nx9142), .A1 (nx9144), .A2 (nx9146)) ;
    aoi222 ix9143 (.Y (nx9142), .A0 (que_out_26__1__14), .A1 (nx9820), .B0 (
           que_out_14__1__14), .B1 (nx9794), .C0 (que_out_11__1__14), .C1 (
           nx9768)) ;
    aoi22 ix9145 (.Y (nx9144), .A0 (que_out_13__1__14), .A1 (nx9742), .B0 (
          que_out_7__1__14), .B1 (nx9716)) ;
    aoi22 ix9147 (.Y (nx9146), .A0 (que_out_12__1__14), .A1 (nx9690), .B0 (
          que_out_1__1__14), .B1 (nx9664)) ;
    or04 ix7173 (.Y (out_column_1__15), .A0 (nx7168), .A1 (nx7142), .A2 (nx7114)
         , .A3 (nx7088)) ;
    nand03 ix7169 (.Y (nx7168), .A0 (nx9150), .A1 (nx9152), .A2 (nx9154)) ;
    aoi222 ix9151 (.Y (nx9150), .A0 (que_out_10__1__15), .A1 (nx10316), .B0 (
           que_out_6__1__15), .B1 (nx10368), .C0 (que_out_9__1__15), .C1 (
           nx10342)) ;
    aoi22 ix9153 (.Y (nx9152), .A0 (que_out_5__1__15), .A1 (nx10264), .B0 (
          que_out_18__1__15), .B1 (nx10290)) ;
    aoi22 ix9155 (.Y (nx9154), .A0 (que_out_17__1__15), .A1 (nx10238), .B0 (
          que_out_20__1__15), .B1 (nx10212)) ;
    nand03 ix7143 (.Y (nx7142), .A0 (nx9157), .A1 (nx9159), .A2 (nx9161)) ;
    aoi222 ix9158 (.Y (nx9157), .A0 (que_out_19__1__15), .A1 (nx10186), .B0 (
           que_out_21__1__15), .B1 (nx10160), .C0 (que_out_8__1__15), .C1 (
           nx10134)) ;
    aoi22 ix9160 (.Y (nx9159), .A0 (que_out_25__1__15), .A1 (nx10082), .B0 (
          que_out_16__1__15), .B1 (nx10108)) ;
    aoi22 ix9162 (.Y (nx9161), .A0 (que_out_24__1__15), .A1 (nx10056), .B0 (
          que_out_22__1__15), .B1 (nx10030)) ;
    nand03 ix7115 (.Y (nx7114), .A0 (nx9164), .A1 (nx9166), .A2 (nx9168)) ;
    aoi222 ix9165 (.Y (nx9164), .A0 (que_out_15__1__15), .A1 (nx9978), .B0 (
           que_out_3__1__15), .B1 (nx10004), .C0 (que_out_23__1__15), .C1 (
           nx9952)) ;
    aoi22 ix9167 (.Y (nx9166), .A0 (que_out_27__1__15), .A1 (nx9926), .B0 (
          que_out_4__1__15), .B1 (nx9900)) ;
    aoi22 ix9169 (.Y (nx9168), .A0 (que_out_0__1__15), .A1 (nx9848), .B0 (
          que_out_2__1__15), .B1 (nx9874)) ;
    nand03 ix7089 (.Y (nx7088), .A0 (nx9171), .A1 (nx9173), .A2 (nx9175)) ;
    aoi222 ix9172 (.Y (nx9171), .A0 (que_out_26__1__15), .A1 (nx9822), .B0 (
           que_out_14__1__15), .B1 (nx9796), .C0 (que_out_11__1__15), .C1 (
           nx9770)) ;
    aoi22 ix9174 (.Y (nx9173), .A0 (que_out_13__1__15), .A1 (nx9744), .B0 (
          que_out_7__1__15), .B1 (nx9718)) ;
    aoi22 ix9176 (.Y (nx9175), .A0 (que_out_12__1__15), .A1 (nx9692), .B0 (
          que_out_1__1__15), .B1 (nx9666)) ;
    or04 ix7283 (.Y (out_column_0__0), .A0 (nx7278), .A1 (nx7252), .A2 (nx7224)
         , .A3 (nx7198)) ;
    nand03 ix7279 (.Y (nx7278), .A0 (nx9179), .A1 (nx9181), .A2 (nx9183)) ;
    aoi222 ix9180 (.Y (nx9179), .A0 (que_out_10__0__0), .A1 (nx10316), .B0 (
           que_out_6__0__0), .B1 (nx10368), .C0 (que_out_9__0__0), .C1 (nx10342)
           ) ;
    aoi22 ix9182 (.Y (nx9181), .A0 (que_out_5__0__0), .A1 (nx10264), .B0 (
          que_out_18__0__0), .B1 (nx10290)) ;
    aoi22 ix9184 (.Y (nx9183), .A0 (que_out_17__0__0), .A1 (nx10238), .B0 (
          que_out_20__0__0), .B1 (nx10212)) ;
    nand03 ix7253 (.Y (nx7252), .A0 (nx9186), .A1 (nx9188), .A2 (nx9190)) ;
    aoi222 ix9187 (.Y (nx9186), .A0 (que_out_19__0__0), .A1 (nx10186), .B0 (
           que_out_21__0__0), .B1 (nx10160), .C0 (que_out_8__0__0), .C1 (nx10134
           )) ;
    aoi22 ix9189 (.Y (nx9188), .A0 (que_out_25__0__0), .A1 (nx10082), .B0 (
          que_out_16__0__0), .B1 (nx10108)) ;
    aoi22 ix9191 (.Y (nx9190), .A0 (que_out_24__0__0), .A1 (nx10056), .B0 (
          que_out_22__0__0), .B1 (nx10030)) ;
    nand03 ix7225 (.Y (nx7224), .A0 (nx9193), .A1 (nx9195), .A2 (nx9197)) ;
    aoi222 ix9194 (.Y (nx9193), .A0 (que_out_15__0__0), .A1 (nx9978), .B0 (
           que_out_3__0__0), .B1 (nx10004), .C0 (que_out_23__0__0), .C1 (nx9952)
           ) ;
    aoi22 ix9196 (.Y (nx9195), .A0 (que_out_27__0__0), .A1 (nx9926), .B0 (
          que_out_4__0__0), .B1 (nx9900)) ;
    aoi22 ix9198 (.Y (nx9197), .A0 (que_out_0__0__0), .A1 (nx9848), .B0 (
          que_out_2__0__0), .B1 (nx9874)) ;
    nand03 ix7199 (.Y (nx7198), .A0 (nx9200), .A1 (nx9202), .A2 (nx9204)) ;
    aoi222 ix9201 (.Y (nx9200), .A0 (que_out_26__0__0), .A1 (nx9822), .B0 (
           que_out_14__0__0), .B1 (nx9796), .C0 (que_out_11__0__0), .C1 (nx9770)
           ) ;
    aoi22 ix9203 (.Y (nx9202), .A0 (que_out_13__0__0), .A1 (nx9744), .B0 (
          que_out_7__0__0), .B1 (nx9718)) ;
    aoi22 ix9205 (.Y (nx9204), .A0 (que_out_12__0__0), .A1 (nx9692), .B0 (
          que_out_1__0__0), .B1 (nx9666)) ;
    or04 ix7393 (.Y (out_column_0__1), .A0 (nx7388), .A1 (nx7362), .A2 (nx7334)
         , .A3 (nx7308)) ;
    nand03 ix7389 (.Y (nx7388), .A0 (nx9208), .A1 (nx9210), .A2 (nx9212)) ;
    aoi222 ix9209 (.Y (nx9208), .A0 (que_out_10__0__1), .A1 (nx10316), .B0 (
           que_out_6__0__1), .B1 (nx10368), .C0 (que_out_9__0__1), .C1 (nx10342)
           ) ;
    aoi22 ix9211 (.Y (nx9210), .A0 (que_out_5__0__1), .A1 (nx10264), .B0 (
          que_out_18__0__1), .B1 (nx10290)) ;
    aoi22 ix9213 (.Y (nx9212), .A0 (que_out_17__0__1), .A1 (nx10238), .B0 (
          que_out_20__0__1), .B1 (nx10212)) ;
    nand03 ix7363 (.Y (nx7362), .A0 (nx9215), .A1 (nx9217), .A2 (nx9219)) ;
    aoi222 ix9216 (.Y (nx9215), .A0 (que_out_19__0__1), .A1 (nx10186), .B0 (
           que_out_21__0__1), .B1 (nx10160), .C0 (que_out_8__0__1), .C1 (nx10134
           )) ;
    aoi22 ix9218 (.Y (nx9217), .A0 (que_out_25__0__1), .A1 (nx10082), .B0 (
          que_out_16__0__1), .B1 (nx10108)) ;
    aoi22 ix9220 (.Y (nx9219), .A0 (que_out_24__0__1), .A1 (nx10056), .B0 (
          que_out_22__0__1), .B1 (nx10030)) ;
    nand03 ix7335 (.Y (nx7334), .A0 (nx9222), .A1 (nx9224), .A2 (nx9226)) ;
    aoi222 ix9223 (.Y (nx9222), .A0 (que_out_15__0__1), .A1 (nx9978), .B0 (
           que_out_3__0__1), .B1 (nx10004), .C0 (que_out_23__0__1), .C1 (nx9952)
           ) ;
    aoi22 ix9225 (.Y (nx9224), .A0 (que_out_27__0__1), .A1 (nx9926), .B0 (
          que_out_4__0__1), .B1 (nx9900)) ;
    aoi22 ix9227 (.Y (nx9226), .A0 (que_out_0__0__1), .A1 (nx9848), .B0 (
          que_out_2__0__1), .B1 (nx9874)) ;
    nand03 ix7309 (.Y (nx7308), .A0 (nx9229), .A1 (nx9231), .A2 (nx9233)) ;
    aoi222 ix9230 (.Y (nx9229), .A0 (que_out_26__0__1), .A1 (nx9822), .B0 (
           que_out_14__0__1), .B1 (nx9796), .C0 (que_out_11__0__1), .C1 (nx9770)
           ) ;
    aoi22 ix9232 (.Y (nx9231), .A0 (que_out_13__0__1), .A1 (nx9744), .B0 (
          que_out_7__0__1), .B1 (nx9718)) ;
    aoi22 ix9234 (.Y (nx9233), .A0 (que_out_12__0__1), .A1 (nx9692), .B0 (
          que_out_1__0__1), .B1 (nx9666)) ;
    or04 ix7503 (.Y (out_column_0__2), .A0 (nx7498), .A1 (nx7472), .A2 (nx7444)
         , .A3 (nx7418)) ;
    nand03 ix7499 (.Y (nx7498), .A0 (nx9237), .A1 (nx9239), .A2 (nx9241)) ;
    aoi222 ix9238 (.Y (nx9237), .A0 (que_out_10__0__2), .A1 (nx10316), .B0 (
           que_out_6__0__2), .B1 (nx10368), .C0 (que_out_9__0__2), .C1 (nx10342)
           ) ;
    aoi22 ix9240 (.Y (nx9239), .A0 (que_out_5__0__2), .A1 (nx10264), .B0 (
          que_out_18__0__2), .B1 (nx10290)) ;
    aoi22 ix9242 (.Y (nx9241), .A0 (que_out_17__0__2), .A1 (nx10238), .B0 (
          que_out_20__0__2), .B1 (nx10212)) ;
    nand03 ix7473 (.Y (nx7472), .A0 (nx9244), .A1 (nx9246), .A2 (nx9248)) ;
    aoi222 ix9245 (.Y (nx9244), .A0 (que_out_19__0__2), .A1 (nx10186), .B0 (
           que_out_21__0__2), .B1 (nx10160), .C0 (que_out_8__0__2), .C1 (nx10134
           )) ;
    aoi22 ix9247 (.Y (nx9246), .A0 (que_out_25__0__2), .A1 (nx10082), .B0 (
          que_out_16__0__2), .B1 (nx10108)) ;
    aoi22 ix9249 (.Y (nx9248), .A0 (que_out_24__0__2), .A1 (nx10056), .B0 (
          que_out_22__0__2), .B1 (nx10030)) ;
    nand03 ix7445 (.Y (nx7444), .A0 (nx9251), .A1 (nx9253), .A2 (nx9255)) ;
    aoi222 ix9252 (.Y (nx9251), .A0 (que_out_15__0__2), .A1 (nx9978), .B0 (
           que_out_3__0__2), .B1 (nx10004), .C0 (que_out_23__0__2), .C1 (nx9952)
           ) ;
    aoi22 ix9254 (.Y (nx9253), .A0 (que_out_27__0__2), .A1 (nx9926), .B0 (
          que_out_4__0__2), .B1 (nx9900)) ;
    aoi22 ix9256 (.Y (nx9255), .A0 (que_out_0__0__2), .A1 (nx9848), .B0 (
          que_out_2__0__2), .B1 (nx9874)) ;
    nand03 ix7419 (.Y (nx7418), .A0 (nx9258), .A1 (nx9260), .A2 (nx9262)) ;
    aoi222 ix9259 (.Y (nx9258), .A0 (que_out_26__0__2), .A1 (nx9822), .B0 (
           que_out_14__0__2), .B1 (nx9796), .C0 (que_out_11__0__2), .C1 (nx9770)
           ) ;
    aoi22 ix9261 (.Y (nx9260), .A0 (que_out_13__0__2), .A1 (nx9744), .B0 (
          que_out_7__0__2), .B1 (nx9718)) ;
    aoi22 ix9263 (.Y (nx9262), .A0 (que_out_12__0__2), .A1 (nx9692), .B0 (
          que_out_1__0__2), .B1 (nx9666)) ;
    or04 ix7613 (.Y (out_column_0__3), .A0 (nx7608), .A1 (nx7582), .A2 (nx7554)
         , .A3 (nx7528)) ;
    nand03 ix7609 (.Y (nx7608), .A0 (nx9266), .A1 (nx9268), .A2 (nx9270)) ;
    aoi222 ix9267 (.Y (nx9266), .A0 (que_out_10__0__3), .A1 (nx10316), .B0 (
           que_out_6__0__3), .B1 (nx10368), .C0 (que_out_9__0__3), .C1 (nx10342)
           ) ;
    aoi22 ix9269 (.Y (nx9268), .A0 (que_out_5__0__3), .A1 (nx10264), .B0 (
          que_out_18__0__3), .B1 (nx10290)) ;
    aoi22 ix9271 (.Y (nx9270), .A0 (que_out_17__0__3), .A1 (nx10238), .B0 (
          que_out_20__0__3), .B1 (nx10212)) ;
    nand03 ix7583 (.Y (nx7582), .A0 (nx9273), .A1 (nx9275), .A2 (nx9277)) ;
    aoi222 ix9274 (.Y (nx9273), .A0 (que_out_19__0__3), .A1 (nx10186), .B0 (
           que_out_21__0__3), .B1 (nx10160), .C0 (que_out_8__0__3), .C1 (nx10134
           )) ;
    aoi22 ix9276 (.Y (nx9275), .A0 (que_out_25__0__3), .A1 (nx10082), .B0 (
          que_out_16__0__3), .B1 (nx10108)) ;
    aoi22 ix9278 (.Y (nx9277), .A0 (que_out_24__0__3), .A1 (nx10056), .B0 (
          que_out_22__0__3), .B1 (nx10030)) ;
    nand03 ix7555 (.Y (nx7554), .A0 (nx9280), .A1 (nx9282), .A2 (nx9284)) ;
    aoi222 ix9281 (.Y (nx9280), .A0 (que_out_15__0__3), .A1 (nx9978), .B0 (
           que_out_3__0__3), .B1 (nx10004), .C0 (que_out_23__0__3), .C1 (nx9952)
           ) ;
    aoi22 ix9283 (.Y (nx9282), .A0 (que_out_27__0__3), .A1 (nx9926), .B0 (
          que_out_4__0__3), .B1 (nx9900)) ;
    aoi22 ix9285 (.Y (nx9284), .A0 (que_out_0__0__3), .A1 (nx9848), .B0 (
          que_out_2__0__3), .B1 (nx9874)) ;
    nand03 ix7529 (.Y (nx7528), .A0 (nx9287), .A1 (nx9289), .A2 (nx9291)) ;
    aoi222 ix9288 (.Y (nx9287), .A0 (que_out_26__0__3), .A1 (nx9822), .B0 (
           que_out_14__0__3), .B1 (nx9796), .C0 (que_out_11__0__3), .C1 (nx9770)
           ) ;
    aoi22 ix9290 (.Y (nx9289), .A0 (que_out_13__0__3), .A1 (nx9744), .B0 (
          que_out_7__0__3), .B1 (nx9718)) ;
    aoi22 ix9292 (.Y (nx9291), .A0 (que_out_12__0__3), .A1 (nx9692), .B0 (
          que_out_1__0__3), .B1 (nx9666)) ;
    or04 ix7723 (.Y (out_column_0__4), .A0 (nx7718), .A1 (nx7692), .A2 (nx7664)
         , .A3 (nx7638)) ;
    nand03 ix7719 (.Y (nx7718), .A0 (nx9295), .A1 (nx9297), .A2 (nx9299)) ;
    aoi222 ix9296 (.Y (nx9295), .A0 (que_out_10__0__4), .A1 (nx10316), .B0 (
           que_out_6__0__4), .B1 (nx10368), .C0 (que_out_9__0__4), .C1 (nx10342)
           ) ;
    aoi22 ix9298 (.Y (nx9297), .A0 (que_out_5__0__4), .A1 (nx10264), .B0 (
          que_out_18__0__4), .B1 (nx10290)) ;
    aoi22 ix9300 (.Y (nx9299), .A0 (que_out_17__0__4), .A1 (nx10238), .B0 (
          que_out_20__0__4), .B1 (nx10212)) ;
    nand03 ix7693 (.Y (nx7692), .A0 (nx9302), .A1 (nx9304), .A2 (nx9306)) ;
    aoi222 ix9303 (.Y (nx9302), .A0 (que_out_19__0__4), .A1 (nx10186), .B0 (
           que_out_21__0__4), .B1 (nx10160), .C0 (que_out_8__0__4), .C1 (nx10134
           )) ;
    aoi22 ix9305 (.Y (nx9304), .A0 (que_out_25__0__4), .A1 (nx10082), .B0 (
          que_out_16__0__4), .B1 (nx10108)) ;
    aoi22 ix9307 (.Y (nx9306), .A0 (que_out_24__0__4), .A1 (nx10056), .B0 (
          que_out_22__0__4), .B1 (nx10030)) ;
    nand03 ix7665 (.Y (nx7664), .A0 (nx9309), .A1 (nx9311), .A2 (nx9313)) ;
    aoi222 ix9310 (.Y (nx9309), .A0 (que_out_15__0__4), .A1 (nx9978), .B0 (
           que_out_3__0__4), .B1 (nx10004), .C0 (que_out_23__0__4), .C1 (nx9952)
           ) ;
    aoi22 ix9312 (.Y (nx9311), .A0 (que_out_27__0__4), .A1 (nx9926), .B0 (
          que_out_4__0__4), .B1 (nx9900)) ;
    aoi22 ix9314 (.Y (nx9313), .A0 (que_out_0__0__4), .A1 (nx9848), .B0 (
          que_out_2__0__4), .B1 (nx9874)) ;
    nand03 ix7639 (.Y (nx7638), .A0 (nx9316), .A1 (nx9318), .A2 (nx9320)) ;
    aoi222 ix9317 (.Y (nx9316), .A0 (que_out_26__0__4), .A1 (nx9822), .B0 (
           que_out_14__0__4), .B1 (nx9796), .C0 (que_out_11__0__4), .C1 (nx9770)
           ) ;
    aoi22 ix9319 (.Y (nx9318), .A0 (que_out_13__0__4), .A1 (nx9744), .B0 (
          que_out_7__0__4), .B1 (nx9718)) ;
    aoi22 ix9321 (.Y (nx9320), .A0 (que_out_12__0__4), .A1 (nx9692), .B0 (
          que_out_1__0__4), .B1 (nx9666)) ;
    or04 ix7833 (.Y (out_column_0__5), .A0 (nx7828), .A1 (nx7802), .A2 (nx7774)
         , .A3 (nx7748)) ;
    nand03 ix7829 (.Y (nx7828), .A0 (nx9324), .A1 (nx9326), .A2 (nx9328)) ;
    aoi222 ix9325 (.Y (nx9324), .A0 (que_out_10__0__5), .A1 (nx10316), .B0 (
           que_out_6__0__5), .B1 (nx10368), .C0 (que_out_9__0__5), .C1 (nx10342)
           ) ;
    aoi22 ix9327 (.Y (nx9326), .A0 (que_out_5__0__5), .A1 (nx10264), .B0 (
          que_out_18__0__5), .B1 (nx10290)) ;
    aoi22 ix9329 (.Y (nx9328), .A0 (que_out_17__0__5), .A1 (nx10238), .B0 (
          que_out_20__0__5), .B1 (nx10212)) ;
    nand03 ix7803 (.Y (nx7802), .A0 (nx9331), .A1 (nx9333), .A2 (nx9335)) ;
    aoi222 ix9332 (.Y (nx9331), .A0 (que_out_19__0__5), .A1 (nx10186), .B0 (
           que_out_21__0__5), .B1 (nx10160), .C0 (que_out_8__0__5), .C1 (nx10134
           )) ;
    aoi22 ix9334 (.Y (nx9333), .A0 (que_out_25__0__5), .A1 (nx10082), .B0 (
          que_out_16__0__5), .B1 (nx10108)) ;
    aoi22 ix9336 (.Y (nx9335), .A0 (que_out_24__0__5), .A1 (nx10056), .B0 (
          que_out_22__0__5), .B1 (nx10030)) ;
    nand03 ix7775 (.Y (nx7774), .A0 (nx9338), .A1 (nx9340), .A2 (nx9342)) ;
    aoi222 ix9339 (.Y (nx9338), .A0 (que_out_15__0__5), .A1 (nx9978), .B0 (
           que_out_3__0__5), .B1 (nx10004), .C0 (que_out_23__0__5), .C1 (nx9952)
           ) ;
    aoi22 ix9341 (.Y (nx9340), .A0 (que_out_27__0__5), .A1 (nx9926), .B0 (
          que_out_4__0__5), .B1 (nx9900)) ;
    aoi22 ix9343 (.Y (nx9342), .A0 (que_out_0__0__5), .A1 (nx9848), .B0 (
          que_out_2__0__5), .B1 (nx9874)) ;
    nand03 ix7749 (.Y (nx7748), .A0 (nx9345), .A1 (nx9347), .A2 (nx9349)) ;
    aoi222 ix9346 (.Y (nx9345), .A0 (que_out_26__0__5), .A1 (nx9822), .B0 (
           que_out_14__0__5), .B1 (nx9796), .C0 (que_out_11__0__5), .C1 (nx9770)
           ) ;
    aoi22 ix9348 (.Y (nx9347), .A0 (que_out_13__0__5), .A1 (nx9744), .B0 (
          que_out_7__0__5), .B1 (nx9718)) ;
    aoi22 ix9350 (.Y (nx9349), .A0 (que_out_12__0__5), .A1 (nx9692), .B0 (
          que_out_1__0__5), .B1 (nx9666)) ;
    or04 ix7943 (.Y (out_column_0__6), .A0 (nx7938), .A1 (nx7912), .A2 (nx7884)
         , .A3 (nx7858)) ;
    nand03 ix7939 (.Y (nx7938), .A0 (nx9353), .A1 (nx9355), .A2 (nx9357)) ;
    aoi222 ix9354 (.Y (nx9353), .A0 (que_out_10__0__6), .A1 (nx10318), .B0 (
           que_out_6__0__6), .B1 (nx10370), .C0 (que_out_9__0__6), .C1 (nx10344)
           ) ;
    aoi22 ix9356 (.Y (nx9355), .A0 (que_out_5__0__6), .A1 (nx10266), .B0 (
          que_out_18__0__6), .B1 (nx10292)) ;
    aoi22 ix9358 (.Y (nx9357), .A0 (que_out_17__0__6), .A1 (nx10240), .B0 (
          que_out_20__0__6), .B1 (nx10214)) ;
    nand03 ix7913 (.Y (nx7912), .A0 (nx9360), .A1 (nx9362), .A2 (nx9364)) ;
    aoi222 ix9361 (.Y (nx9360), .A0 (que_out_19__0__6), .A1 (nx10188), .B0 (
           que_out_21__0__6), .B1 (nx10162), .C0 (que_out_8__0__6), .C1 (nx10136
           )) ;
    aoi22 ix9363 (.Y (nx9362), .A0 (que_out_25__0__6), .A1 (nx10084), .B0 (
          que_out_16__0__6), .B1 (nx10110)) ;
    aoi22 ix9365 (.Y (nx9364), .A0 (que_out_24__0__6), .A1 (nx10058), .B0 (
          que_out_22__0__6), .B1 (nx10032)) ;
    nand03 ix7885 (.Y (nx7884), .A0 (nx9367), .A1 (nx9369), .A2 (nx9371)) ;
    aoi222 ix9368 (.Y (nx9367), .A0 (que_out_15__0__6), .A1 (nx9980), .B0 (
           que_out_3__0__6), .B1 (nx10006), .C0 (que_out_23__0__6), .C1 (nx9954)
           ) ;
    aoi22 ix9370 (.Y (nx9369), .A0 (que_out_27__0__6), .A1 (nx9928), .B0 (
          que_out_4__0__6), .B1 (nx9902)) ;
    aoi22 ix9372 (.Y (nx9371), .A0 (que_out_0__0__6), .A1 (nx9850), .B0 (
          que_out_2__0__6), .B1 (nx9876)) ;
    nand03 ix7859 (.Y (nx7858), .A0 (nx9374), .A1 (nx9376), .A2 (nx9378)) ;
    aoi222 ix9375 (.Y (nx9374), .A0 (que_out_26__0__6), .A1 (nx9824), .B0 (
           que_out_14__0__6), .B1 (nx9798), .C0 (que_out_11__0__6), .C1 (nx9772)
           ) ;
    aoi22 ix9377 (.Y (nx9376), .A0 (que_out_13__0__6), .A1 (nx9746), .B0 (
          que_out_7__0__6), .B1 (nx9720)) ;
    aoi22 ix9379 (.Y (nx9378), .A0 (que_out_12__0__6), .A1 (nx9694), .B0 (
          que_out_1__0__6), .B1 (nx9668)) ;
    or04 ix8053 (.Y (out_column_0__7), .A0 (nx8048), .A1 (nx8022), .A2 (nx7994)
         , .A3 (nx7968)) ;
    nand03 ix8049 (.Y (nx8048), .A0 (nx9382), .A1 (nx9384), .A2 (nx9386)) ;
    aoi222 ix9383 (.Y (nx9382), .A0 (que_out_10__0__7), .A1 (nx10318), .B0 (
           que_out_6__0__7), .B1 (nx10370), .C0 (que_out_9__0__7), .C1 (nx10344)
           ) ;
    aoi22 ix9385 (.Y (nx9384), .A0 (que_out_5__0__7), .A1 (nx10266), .B0 (
          que_out_18__0__7), .B1 (nx10292)) ;
    aoi22 ix9387 (.Y (nx9386), .A0 (que_out_17__0__7), .A1 (nx10240), .B0 (
          que_out_20__0__7), .B1 (nx10214)) ;
    nand03 ix8023 (.Y (nx8022), .A0 (nx9389), .A1 (nx9391), .A2 (nx9393)) ;
    aoi222 ix9390 (.Y (nx9389), .A0 (que_out_19__0__7), .A1 (nx10188), .B0 (
           que_out_21__0__7), .B1 (nx10162), .C0 (que_out_8__0__7), .C1 (nx10136
           )) ;
    aoi22 ix9392 (.Y (nx9391), .A0 (que_out_25__0__7), .A1 (nx10084), .B0 (
          que_out_16__0__7), .B1 (nx10110)) ;
    aoi22 ix9394 (.Y (nx9393), .A0 (que_out_24__0__7), .A1 (nx10058), .B0 (
          que_out_22__0__7), .B1 (nx10032)) ;
    nand03 ix7995 (.Y (nx7994), .A0 (nx9396), .A1 (nx9398), .A2 (nx9400)) ;
    aoi222 ix9397 (.Y (nx9396), .A0 (que_out_15__0__7), .A1 (nx9980), .B0 (
           que_out_3__0__7), .B1 (nx10006), .C0 (que_out_23__0__7), .C1 (nx9954)
           ) ;
    aoi22 ix9399 (.Y (nx9398), .A0 (que_out_27__0__7), .A1 (nx9928), .B0 (
          que_out_4__0__7), .B1 (nx9902)) ;
    aoi22 ix9401 (.Y (nx9400), .A0 (que_out_0__0__7), .A1 (nx9850), .B0 (
          que_out_2__0__7), .B1 (nx9876)) ;
    nand03 ix7969 (.Y (nx7968), .A0 (nx9403), .A1 (nx9405), .A2 (nx9407)) ;
    aoi222 ix9404 (.Y (nx9403), .A0 (que_out_26__0__7), .A1 (nx9824), .B0 (
           que_out_14__0__7), .B1 (nx9798), .C0 (que_out_11__0__7), .C1 (nx9772)
           ) ;
    aoi22 ix9406 (.Y (nx9405), .A0 (que_out_13__0__7), .A1 (nx9746), .B0 (
          que_out_7__0__7), .B1 (nx9720)) ;
    aoi22 ix9408 (.Y (nx9407), .A0 (que_out_12__0__7), .A1 (nx9694), .B0 (
          que_out_1__0__7), .B1 (nx9668)) ;
    or04 ix8163 (.Y (out_column_0__8), .A0 (nx8158), .A1 (nx8132), .A2 (nx8104)
         , .A3 (nx8078)) ;
    nand03 ix8159 (.Y (nx8158), .A0 (nx9411), .A1 (nx9413), .A2 (nx9415)) ;
    aoi222 ix9412 (.Y (nx9411), .A0 (que_out_10__0__8), .A1 (nx10318), .B0 (
           que_out_6__0__8), .B1 (nx10370), .C0 (que_out_9__0__8), .C1 (nx10344)
           ) ;
    aoi22 ix9414 (.Y (nx9413), .A0 (que_out_5__0__8), .A1 (nx10266), .B0 (
          que_out_18__0__8), .B1 (nx10292)) ;
    aoi22 ix9416 (.Y (nx9415), .A0 (que_out_17__0__8), .A1 (nx10240), .B0 (
          que_out_20__0__8), .B1 (nx10214)) ;
    nand03 ix8133 (.Y (nx8132), .A0 (nx9418), .A1 (nx9420), .A2 (nx9422)) ;
    aoi222 ix9419 (.Y (nx9418), .A0 (que_out_19__0__8), .A1 (nx10188), .B0 (
           que_out_21__0__8), .B1 (nx10162), .C0 (que_out_8__0__8), .C1 (nx10136
           )) ;
    aoi22 ix9421 (.Y (nx9420), .A0 (que_out_25__0__8), .A1 (nx10084), .B0 (
          que_out_16__0__8), .B1 (nx10110)) ;
    aoi22 ix9423 (.Y (nx9422), .A0 (que_out_24__0__8), .A1 (nx10058), .B0 (
          que_out_22__0__8), .B1 (nx10032)) ;
    nand03 ix8105 (.Y (nx8104), .A0 (nx9425), .A1 (nx9427), .A2 (nx9429)) ;
    aoi222 ix9426 (.Y (nx9425), .A0 (que_out_15__0__8), .A1 (nx9980), .B0 (
           que_out_3__0__8), .B1 (nx10006), .C0 (que_out_23__0__8), .C1 (nx9954)
           ) ;
    aoi22 ix9428 (.Y (nx9427), .A0 (que_out_27__0__8), .A1 (nx9928), .B0 (
          que_out_4__0__8), .B1 (nx9902)) ;
    aoi22 ix9430 (.Y (nx9429), .A0 (que_out_0__0__8), .A1 (nx9850), .B0 (
          que_out_2__0__8), .B1 (nx9876)) ;
    nand03 ix8079 (.Y (nx8078), .A0 (nx9432), .A1 (nx9434), .A2 (nx9436)) ;
    aoi222 ix9433 (.Y (nx9432), .A0 (que_out_26__0__8), .A1 (nx9824), .B0 (
           que_out_14__0__8), .B1 (nx9798), .C0 (que_out_11__0__8), .C1 (nx9772)
           ) ;
    aoi22 ix9435 (.Y (nx9434), .A0 (que_out_13__0__8), .A1 (nx9746), .B0 (
          que_out_7__0__8), .B1 (nx9720)) ;
    aoi22 ix9437 (.Y (nx9436), .A0 (que_out_12__0__8), .A1 (nx9694), .B0 (
          que_out_1__0__8), .B1 (nx9668)) ;
    or04 ix8273 (.Y (out_column_0__9), .A0 (nx8268), .A1 (nx8242), .A2 (nx8214)
         , .A3 (nx8188)) ;
    nand03 ix8269 (.Y (nx8268), .A0 (nx9440), .A1 (nx9442), .A2 (nx9444)) ;
    aoi222 ix9441 (.Y (nx9440), .A0 (que_out_10__0__9), .A1 (nx10318), .B0 (
           que_out_6__0__9), .B1 (nx10370), .C0 (que_out_9__0__9), .C1 (nx10344)
           ) ;
    aoi22 ix9443 (.Y (nx9442), .A0 (que_out_5__0__9), .A1 (nx10266), .B0 (
          que_out_18__0__9), .B1 (nx10292)) ;
    aoi22 ix9445 (.Y (nx9444), .A0 (que_out_17__0__9), .A1 (nx10240), .B0 (
          que_out_20__0__9), .B1 (nx10214)) ;
    nand03 ix8243 (.Y (nx8242), .A0 (nx9447), .A1 (nx9449), .A2 (nx9451)) ;
    aoi222 ix9448 (.Y (nx9447), .A0 (que_out_19__0__9), .A1 (nx10188), .B0 (
           que_out_21__0__9), .B1 (nx10162), .C0 (que_out_8__0__9), .C1 (nx10136
           )) ;
    aoi22 ix9450 (.Y (nx9449), .A0 (que_out_25__0__9), .A1 (nx10084), .B0 (
          que_out_16__0__9), .B1 (nx10110)) ;
    aoi22 ix9452 (.Y (nx9451), .A0 (que_out_24__0__9), .A1 (nx10058), .B0 (
          que_out_22__0__9), .B1 (nx10032)) ;
    nand03 ix8215 (.Y (nx8214), .A0 (nx9454), .A1 (nx9456), .A2 (nx9458)) ;
    aoi222 ix9455 (.Y (nx9454), .A0 (que_out_15__0__9), .A1 (nx9980), .B0 (
           que_out_3__0__9), .B1 (nx10006), .C0 (que_out_23__0__9), .C1 (nx9954)
           ) ;
    aoi22 ix9457 (.Y (nx9456), .A0 (que_out_27__0__9), .A1 (nx9928), .B0 (
          que_out_4__0__9), .B1 (nx9902)) ;
    aoi22 ix9459 (.Y (nx9458), .A0 (que_out_0__0__9), .A1 (nx9850), .B0 (
          que_out_2__0__9), .B1 (nx9876)) ;
    nand03 ix8189 (.Y (nx8188), .A0 (nx9461), .A1 (nx9463), .A2 (nx9465)) ;
    aoi222 ix9462 (.Y (nx9461), .A0 (que_out_26__0__9), .A1 (nx9824), .B0 (
           que_out_14__0__9), .B1 (nx9798), .C0 (que_out_11__0__9), .C1 (nx9772)
           ) ;
    aoi22 ix9464 (.Y (nx9463), .A0 (que_out_13__0__9), .A1 (nx9746), .B0 (
          que_out_7__0__9), .B1 (nx9720)) ;
    aoi22 ix9466 (.Y (nx9465), .A0 (que_out_12__0__9), .A1 (nx9694), .B0 (
          que_out_1__0__9), .B1 (nx9668)) ;
    or04 ix8383 (.Y (out_column_0__10), .A0 (nx8378), .A1 (nx8352), .A2 (nx8324)
         , .A3 (nx8298)) ;
    nand03 ix8379 (.Y (nx8378), .A0 (nx9469), .A1 (nx9471), .A2 (nx9473)) ;
    aoi222 ix9470 (.Y (nx9469), .A0 (que_out_10__0__10), .A1 (nx10318), .B0 (
           que_out_6__0__10), .B1 (nx10370), .C0 (que_out_9__0__10), .C1 (
           nx10344)) ;
    aoi22 ix9472 (.Y (nx9471), .A0 (que_out_5__0__10), .A1 (nx10266), .B0 (
          que_out_18__0__10), .B1 (nx10292)) ;
    aoi22 ix9474 (.Y (nx9473), .A0 (que_out_17__0__10), .A1 (nx10240), .B0 (
          que_out_20__0__10), .B1 (nx10214)) ;
    nand03 ix8353 (.Y (nx8352), .A0 (nx9476), .A1 (nx9478), .A2 (nx9480)) ;
    aoi222 ix9477 (.Y (nx9476), .A0 (que_out_19__0__10), .A1 (nx10188), .B0 (
           que_out_21__0__10), .B1 (nx10162), .C0 (que_out_8__0__10), .C1 (
           nx10136)) ;
    aoi22 ix9479 (.Y (nx9478), .A0 (que_out_25__0__10), .A1 (nx10084), .B0 (
          que_out_16__0__10), .B1 (nx10110)) ;
    aoi22 ix9481 (.Y (nx9480), .A0 (que_out_24__0__10), .A1 (nx10058), .B0 (
          que_out_22__0__10), .B1 (nx10032)) ;
    nand03 ix8325 (.Y (nx8324), .A0 (nx9483), .A1 (nx9485), .A2 (nx9487)) ;
    aoi222 ix9484 (.Y (nx9483), .A0 (que_out_15__0__10), .A1 (nx9980), .B0 (
           que_out_3__0__10), .B1 (nx10006), .C0 (que_out_23__0__10), .C1 (
           nx9954)) ;
    aoi22 ix9486 (.Y (nx9485), .A0 (que_out_27__0__10), .A1 (nx9928), .B0 (
          que_out_4__0__10), .B1 (nx9902)) ;
    aoi22 ix9488 (.Y (nx9487), .A0 (que_out_0__0__10), .A1 (nx9850), .B0 (
          que_out_2__0__10), .B1 (nx9876)) ;
    nand03 ix8299 (.Y (nx8298), .A0 (nx9490), .A1 (nx9492), .A2 (nx9494)) ;
    aoi222 ix9491 (.Y (nx9490), .A0 (que_out_26__0__10), .A1 (nx9824), .B0 (
           que_out_14__0__10), .B1 (nx9798), .C0 (que_out_11__0__10), .C1 (
           nx9772)) ;
    aoi22 ix9493 (.Y (nx9492), .A0 (que_out_13__0__10), .A1 (nx9746), .B0 (
          que_out_7__0__10), .B1 (nx9720)) ;
    aoi22 ix9495 (.Y (nx9494), .A0 (que_out_12__0__10), .A1 (nx9694), .B0 (
          que_out_1__0__10), .B1 (nx9668)) ;
    or04 ix8493 (.Y (out_column_0__11), .A0 (nx8488), .A1 (nx8462), .A2 (nx8434)
         , .A3 (nx8408)) ;
    nand03 ix8489 (.Y (nx8488), .A0 (nx9498), .A1 (nx9500), .A2 (nx9502)) ;
    aoi222 ix9499 (.Y (nx9498), .A0 (que_out_10__0__11), .A1 (nx10318), .B0 (
           que_out_6__0__11), .B1 (nx10370), .C0 (que_out_9__0__11), .C1 (
           nx10344)) ;
    aoi22 ix9501 (.Y (nx9500), .A0 (que_out_5__0__11), .A1 (nx10266), .B0 (
          que_out_18__0__11), .B1 (nx10292)) ;
    aoi22 ix9503 (.Y (nx9502), .A0 (que_out_17__0__11), .A1 (nx10240), .B0 (
          que_out_20__0__11), .B1 (nx10214)) ;
    nand03 ix8463 (.Y (nx8462), .A0 (nx9505), .A1 (nx9507), .A2 (nx9509)) ;
    aoi222 ix9506 (.Y (nx9505), .A0 (que_out_19__0__11), .A1 (nx10188), .B0 (
           que_out_21__0__11), .B1 (nx10162), .C0 (que_out_8__0__11), .C1 (
           nx10136)) ;
    aoi22 ix9508 (.Y (nx9507), .A0 (que_out_25__0__11), .A1 (nx10084), .B0 (
          que_out_16__0__11), .B1 (nx10110)) ;
    aoi22 ix9510 (.Y (nx9509), .A0 (que_out_24__0__11), .A1 (nx10058), .B0 (
          que_out_22__0__11), .B1 (nx10032)) ;
    nand03 ix8435 (.Y (nx8434), .A0 (nx9512), .A1 (nx9514), .A2 (nx9516)) ;
    aoi222 ix9513 (.Y (nx9512), .A0 (que_out_15__0__11), .A1 (nx9980), .B0 (
           que_out_3__0__11), .B1 (nx10006), .C0 (que_out_23__0__11), .C1 (
           nx9954)) ;
    aoi22 ix9515 (.Y (nx9514), .A0 (que_out_27__0__11), .A1 (nx9928), .B0 (
          que_out_4__0__11), .B1 (nx9902)) ;
    aoi22 ix9517 (.Y (nx9516), .A0 (que_out_0__0__11), .A1 (nx9850), .B0 (
          que_out_2__0__11), .B1 (nx9876)) ;
    nand03 ix8409 (.Y (nx8408), .A0 (nx9519), .A1 (nx9521), .A2 (nx9523)) ;
    aoi222 ix9520 (.Y (nx9519), .A0 (que_out_26__0__11), .A1 (nx9824), .B0 (
           que_out_14__0__11), .B1 (nx9798), .C0 (que_out_11__0__11), .C1 (
           nx9772)) ;
    aoi22 ix9522 (.Y (nx9521), .A0 (que_out_13__0__11), .A1 (nx9746), .B0 (
          que_out_7__0__11), .B1 (nx9720)) ;
    aoi22 ix9524 (.Y (nx9523), .A0 (que_out_12__0__11), .A1 (nx9694), .B0 (
          que_out_1__0__11), .B1 (nx9668)) ;
    or04 ix8603 (.Y (out_column_0__12), .A0 (nx8598), .A1 (nx8572), .A2 (nx8544)
         , .A3 (nx8518)) ;
    nand03 ix8599 (.Y (nx8598), .A0 (nx9527), .A1 (nx9529), .A2 (nx9531)) ;
    aoi222 ix9528 (.Y (nx9527), .A0 (que_out_10__0__12), .A1 (nx10318), .B0 (
           que_out_6__0__12), .B1 (nx10370), .C0 (que_out_9__0__12), .C1 (
           nx10344)) ;
    aoi22 ix9530 (.Y (nx9529), .A0 (que_out_5__0__12), .A1 (nx10266), .B0 (
          que_out_18__0__12), .B1 (nx10292)) ;
    aoi22 ix9532 (.Y (nx9531), .A0 (que_out_17__0__12), .A1 (nx10240), .B0 (
          que_out_20__0__12), .B1 (nx10214)) ;
    nand03 ix8573 (.Y (nx8572), .A0 (nx9534), .A1 (nx9536), .A2 (nx9538)) ;
    aoi222 ix9535 (.Y (nx9534), .A0 (que_out_19__0__12), .A1 (nx10188), .B0 (
           que_out_21__0__12), .B1 (nx10162), .C0 (que_out_8__0__12), .C1 (
           nx10136)) ;
    aoi22 ix9537 (.Y (nx9536), .A0 (que_out_25__0__12), .A1 (nx10084), .B0 (
          que_out_16__0__12), .B1 (nx10110)) ;
    aoi22 ix9539 (.Y (nx9538), .A0 (que_out_24__0__12), .A1 (nx10058), .B0 (
          que_out_22__0__12), .B1 (nx10032)) ;
    nand03 ix8545 (.Y (nx8544), .A0 (nx9541), .A1 (nx9543), .A2 (nx9545)) ;
    aoi222 ix9542 (.Y (nx9541), .A0 (que_out_15__0__12), .A1 (nx9980), .B0 (
           que_out_3__0__12), .B1 (nx10006), .C0 (que_out_23__0__12), .C1 (
           nx9954)) ;
    aoi22 ix9544 (.Y (nx9543), .A0 (que_out_27__0__12), .A1 (nx9928), .B0 (
          que_out_4__0__12), .B1 (nx9902)) ;
    aoi22 ix9546 (.Y (nx9545), .A0 (que_out_0__0__12), .A1 (nx9850), .B0 (
          que_out_2__0__12), .B1 (nx9876)) ;
    nand03 ix8519 (.Y (nx8518), .A0 (nx9548), .A1 (nx9550), .A2 (nx9552)) ;
    aoi222 ix9549 (.Y (nx9548), .A0 (que_out_26__0__12), .A1 (nx9824), .B0 (
           que_out_14__0__12), .B1 (nx9798), .C0 (que_out_11__0__12), .C1 (
           nx9772)) ;
    aoi22 ix9551 (.Y (nx9550), .A0 (que_out_13__0__12), .A1 (nx9746), .B0 (
          que_out_7__0__12), .B1 (nx9720)) ;
    aoi22 ix9553 (.Y (nx9552), .A0 (que_out_12__0__12), .A1 (nx9694), .B0 (
          que_out_1__0__12), .B1 (nx9668)) ;
    or04 ix8713 (.Y (out_column_0__13), .A0 (nx8708), .A1 (nx8682), .A2 (nx8654)
         , .A3 (nx8628)) ;
    nand03 ix8709 (.Y (nx8708), .A0 (nx9556), .A1 (nx9558), .A2 (nx9560)) ;
    aoi222 ix9557 (.Y (nx9556), .A0 (que_out_10__0__13), .A1 (nx10320), .B0 (
           que_out_6__0__13), .B1 (nx10372), .C0 (que_out_9__0__13), .C1 (
           nx10346)) ;
    aoi22 ix9559 (.Y (nx9558), .A0 (que_out_5__0__13), .A1 (nx10268), .B0 (
          que_out_18__0__13), .B1 (nx10294)) ;
    aoi22 ix9561 (.Y (nx9560), .A0 (que_out_17__0__13), .A1 (nx10242), .B0 (
          que_out_20__0__13), .B1 (nx10216)) ;
    nand03 ix8683 (.Y (nx8682), .A0 (nx9563), .A1 (nx9565), .A2 (nx9567)) ;
    aoi222 ix9564 (.Y (nx9563), .A0 (que_out_19__0__13), .A1 (nx10190), .B0 (
           que_out_21__0__13), .B1 (nx10164), .C0 (que_out_8__0__13), .C1 (
           nx10138)) ;
    aoi22 ix9566 (.Y (nx9565), .A0 (que_out_25__0__13), .A1 (nx10086), .B0 (
          que_out_16__0__13), .B1 (nx10112)) ;
    aoi22 ix9568 (.Y (nx9567), .A0 (que_out_24__0__13), .A1 (nx10060), .B0 (
          que_out_22__0__13), .B1 (nx10034)) ;
    nand03 ix8655 (.Y (nx8654), .A0 (nx9570), .A1 (nx9572), .A2 (nx9574)) ;
    aoi222 ix9571 (.Y (nx9570), .A0 (que_out_15__0__13), .A1 (nx9982), .B0 (
           que_out_3__0__13), .B1 (nx10008), .C0 (que_out_23__0__13), .C1 (
           nx9956)) ;
    aoi22 ix9573 (.Y (nx9572), .A0 (que_out_27__0__13), .A1 (nx9930), .B0 (
          que_out_4__0__13), .B1 (nx9904)) ;
    aoi22 ix9575 (.Y (nx9574), .A0 (que_out_0__0__13), .A1 (nx9852), .B0 (
          que_out_2__0__13), .B1 (nx9878)) ;
    nand03 ix8629 (.Y (nx8628), .A0 (nx9577), .A1 (nx9579), .A2 (nx9581)) ;
    aoi222 ix9578 (.Y (nx9577), .A0 (que_out_26__0__13), .A1 (nx9826), .B0 (
           que_out_14__0__13), .B1 (nx9800), .C0 (que_out_11__0__13), .C1 (
           nx9774)) ;
    aoi22 ix9580 (.Y (nx9579), .A0 (que_out_13__0__13), .A1 (nx9748), .B0 (
          que_out_7__0__13), .B1 (nx9722)) ;
    aoi22 ix9582 (.Y (nx9581), .A0 (que_out_12__0__13), .A1 (nx9696), .B0 (
          que_out_1__0__13), .B1 (nx9670)) ;
    or04 ix8823 (.Y (out_column_0__14), .A0 (nx8818), .A1 (nx8792), .A2 (nx8764)
         , .A3 (nx8738)) ;
    nand03 ix8819 (.Y (nx8818), .A0 (nx9585), .A1 (nx9587), .A2 (nx9589)) ;
    aoi222 ix9586 (.Y (nx9585), .A0 (que_out_10__0__14), .A1 (nx10320), .B0 (
           que_out_6__0__14), .B1 (nx10372), .C0 (que_out_9__0__14), .C1 (
           nx10346)) ;
    aoi22 ix9588 (.Y (nx9587), .A0 (que_out_5__0__14), .A1 (nx10268), .B0 (
          que_out_18__0__14), .B1 (nx10294)) ;
    aoi22 ix9590 (.Y (nx9589), .A0 (que_out_17__0__14), .A1 (nx10242), .B0 (
          que_out_20__0__14), .B1 (nx10216)) ;
    nand03 ix8793 (.Y (nx8792), .A0 (nx9592), .A1 (nx9594), .A2 (nx9596)) ;
    aoi222 ix9593 (.Y (nx9592), .A0 (que_out_19__0__14), .A1 (nx10190), .B0 (
           que_out_21__0__14), .B1 (nx10164), .C0 (que_out_8__0__14), .C1 (
           nx10138)) ;
    aoi22 ix9595 (.Y (nx9594), .A0 (que_out_25__0__14), .A1 (nx10086), .B0 (
          que_out_16__0__14), .B1 (nx10112)) ;
    aoi22 ix9597 (.Y (nx9596), .A0 (que_out_24__0__14), .A1 (nx10060), .B0 (
          que_out_22__0__14), .B1 (nx10034)) ;
    nand03 ix8765 (.Y (nx8764), .A0 (nx9599), .A1 (nx9601), .A2 (nx9603)) ;
    aoi222 ix9600 (.Y (nx9599), .A0 (que_out_15__0__14), .A1 (nx9982), .B0 (
           que_out_3__0__14), .B1 (nx10008), .C0 (que_out_23__0__14), .C1 (
           nx9956)) ;
    aoi22 ix9602 (.Y (nx9601), .A0 (que_out_27__0__14), .A1 (nx9930), .B0 (
          que_out_4__0__14), .B1 (nx9904)) ;
    aoi22 ix9604 (.Y (nx9603), .A0 (que_out_0__0__14), .A1 (nx9852), .B0 (
          que_out_2__0__14), .B1 (nx9878)) ;
    nand03 ix8739 (.Y (nx8738), .A0 (nx9606), .A1 (nx9608), .A2 (nx9610)) ;
    aoi222 ix9607 (.Y (nx9606), .A0 (que_out_26__0__14), .A1 (nx9826), .B0 (
           que_out_14__0__14), .B1 (nx9800), .C0 (que_out_11__0__14), .C1 (
           nx9774)) ;
    aoi22 ix9609 (.Y (nx9608), .A0 (que_out_13__0__14), .A1 (nx9748), .B0 (
          que_out_7__0__14), .B1 (nx9722)) ;
    aoi22 ix9611 (.Y (nx9610), .A0 (que_out_12__0__14), .A1 (nx9696), .B0 (
          que_out_1__0__14), .B1 (nx9670)) ;
    or04 ix8933 (.Y (out_column_0__15), .A0 (nx8928), .A1 (nx8902), .A2 (nx8874)
         , .A3 (nx8848)) ;
    nand03 ix8929 (.Y (nx8928), .A0 (nx9614), .A1 (nx9616), .A2 (nx9618)) ;
    aoi222 ix9615 (.Y (nx9614), .A0 (que_out_10__0__15), .A1 (nx10320), .B0 (
           que_out_6__0__15), .B1 (nx10372), .C0 (que_out_9__0__15), .C1 (
           nx10346)) ;
    aoi22 ix9617 (.Y (nx9616), .A0 (que_out_5__0__15), .A1 (nx10268), .B0 (
          que_out_18__0__15), .B1 (nx10294)) ;
    aoi22 ix9619 (.Y (nx9618), .A0 (que_out_17__0__15), .A1 (nx10242), .B0 (
          que_out_20__0__15), .B1 (nx10216)) ;
    nand03 ix8903 (.Y (nx8902), .A0 (nx9621), .A1 (nx9623), .A2 (nx9625)) ;
    aoi222 ix9622 (.Y (nx9621), .A0 (que_out_19__0__15), .A1 (nx10190), .B0 (
           que_out_21__0__15), .B1 (nx10164), .C0 (que_out_8__0__15), .C1 (
           nx10138)) ;
    aoi22 ix9624 (.Y (nx9623), .A0 (que_out_25__0__15), .A1 (nx10086), .B0 (
          que_out_16__0__15), .B1 (nx10112)) ;
    aoi22 ix9626 (.Y (nx9625), .A0 (que_out_24__0__15), .A1 (nx10060), .B0 (
          que_out_22__0__15), .B1 (nx10034)) ;
    nand03 ix8875 (.Y (nx8874), .A0 (nx9628), .A1 (nx9630), .A2 (nx9632)) ;
    aoi222 ix9629 (.Y (nx9628), .A0 (que_out_15__0__15), .A1 (nx9982), .B0 (
           que_out_3__0__15), .B1 (nx10008), .C0 (que_out_23__0__15), .C1 (
           nx9956)) ;
    aoi22 ix9631 (.Y (nx9630), .A0 (que_out_27__0__15), .A1 (nx9930), .B0 (
          que_out_4__0__15), .B1 (nx9904)) ;
    aoi22 ix9633 (.Y (nx9632), .A0 (que_out_0__0__15), .A1 (nx9852), .B0 (
          que_out_2__0__15), .B1 (nx9878)) ;
    nand03 ix8849 (.Y (nx8848), .A0 (nx9635), .A1 (nx9637), .A2 (nx9639)) ;
    aoi222 ix9636 (.Y (nx9635), .A0 (que_out_26__0__15), .A1 (nx9826), .B0 (
           que_out_14__0__15), .B1 (nx9800), .C0 (que_out_11__0__15), .C1 (
           nx9774)) ;
    aoi22 ix9638 (.Y (nx9637), .A0 (que_out_13__0__15), .A1 (nx9748), .B0 (
          que_out_7__0__15), .B1 (nx9722)) ;
    aoi22 ix9640 (.Y (nx9639), .A0 (que_out_12__0__15), .A1 (nx9696), .B0 (
          que_out_1__0__15), .B1 (nx9670)) ;
    inv02 ix6944 (.Y (nx6943), .A (nx88)) ;
    inv02 ix9647 (.Y (nx9648), .A (nx10378)) ;
    inv02 ix9649 (.Y (nx9650), .A (nx10378)) ;
    inv02 ix9651 (.Y (nx9652), .A (nx10378)) ;
    inv02 ix9653 (.Y (nx9654), .A (nx10378)) ;
    inv02 ix9655 (.Y (nx9656), .A (nx10378)) ;
    inv02 ix9657 (.Y (nx9658), .A (nx10378)) ;
    inv02 ix9659 (.Y (nx9660), .A (nx10378)) ;
    inv02 ix9661 (.Y (nx9662), .A (nx10380)) ;
    inv02 ix9663 (.Y (nx9664), .A (nx10380)) ;
    inv02 ix9665 (.Y (nx9666), .A (nx10380)) ;
    inv02 ix9667 (.Y (nx9668), .A (nx10380)) ;
    inv02 ix9669 (.Y (nx9670), .A (nx10380)) ;
    inv02 ix9673 (.Y (nx9674), .A (nx10382)) ;
    inv02 ix9675 (.Y (nx9676), .A (nx10382)) ;
    inv02 ix9677 (.Y (nx9678), .A (nx10382)) ;
    inv02 ix9679 (.Y (nx9680), .A (nx10382)) ;
    inv02 ix9681 (.Y (nx9682), .A (nx10382)) ;
    inv02 ix9683 (.Y (nx9684), .A (nx10382)) ;
    inv02 ix9685 (.Y (nx9686), .A (nx10382)) ;
    inv02 ix9687 (.Y (nx9688), .A (nx10384)) ;
    inv02 ix9689 (.Y (nx9690), .A (nx10384)) ;
    inv02 ix9691 (.Y (nx9692), .A (nx10384)) ;
    inv02 ix9693 (.Y (nx9694), .A (nx10384)) ;
    inv02 ix9695 (.Y (nx9696), .A (nx10384)) ;
    inv02 ix9699 (.Y (nx9700), .A (nx10386)) ;
    inv02 ix9701 (.Y (nx9702), .A (nx10386)) ;
    inv02 ix9703 (.Y (nx9704), .A (nx10386)) ;
    inv02 ix9705 (.Y (nx9706), .A (nx10386)) ;
    inv02 ix9707 (.Y (nx9708), .A (nx10386)) ;
    inv02 ix9709 (.Y (nx9710), .A (nx10386)) ;
    inv02 ix9711 (.Y (nx9712), .A (nx10386)) ;
    inv02 ix9713 (.Y (nx9714), .A (nx10388)) ;
    inv02 ix9715 (.Y (nx9716), .A (nx10388)) ;
    inv02 ix9717 (.Y (nx9718), .A (nx10388)) ;
    inv02 ix9719 (.Y (nx9720), .A (nx10388)) ;
    inv02 ix9721 (.Y (nx9722), .A (nx10388)) ;
    inv02 ix9725 (.Y (nx9726), .A (nx10390)) ;
    inv02 ix9727 (.Y (nx9728), .A (nx10390)) ;
    inv02 ix9729 (.Y (nx9730), .A (nx10390)) ;
    inv02 ix9731 (.Y (nx9732), .A (nx10390)) ;
    inv02 ix9733 (.Y (nx9734), .A (nx10390)) ;
    inv02 ix9735 (.Y (nx9736), .A (nx10390)) ;
    inv02 ix9737 (.Y (nx9738), .A (nx10390)) ;
    inv02 ix9739 (.Y (nx9740), .A (nx10392)) ;
    inv02 ix9741 (.Y (nx9742), .A (nx10392)) ;
    inv02 ix9743 (.Y (nx9744), .A (nx10392)) ;
    inv02 ix9745 (.Y (nx9746), .A (nx10392)) ;
    inv02 ix9747 (.Y (nx9748), .A (nx10392)) ;
    inv02 ix9751 (.Y (nx9752), .A (nx10394)) ;
    inv02 ix9753 (.Y (nx9754), .A (nx10394)) ;
    inv02 ix9755 (.Y (nx9756), .A (nx10394)) ;
    inv02 ix9757 (.Y (nx9758), .A (nx10394)) ;
    inv02 ix9759 (.Y (nx9760), .A (nx10394)) ;
    inv02 ix9761 (.Y (nx9762), .A (nx10394)) ;
    inv02 ix9763 (.Y (nx9764), .A (nx10394)) ;
    inv02 ix9765 (.Y (nx9766), .A (nx10396)) ;
    inv02 ix9767 (.Y (nx9768), .A (nx10396)) ;
    inv02 ix9769 (.Y (nx9770), .A (nx10396)) ;
    inv02 ix9771 (.Y (nx9772), .A (nx10396)) ;
    inv02 ix9773 (.Y (nx9774), .A (nx10396)) ;
    inv02 ix9777 (.Y (nx9778), .A (nx10398)) ;
    inv02 ix9779 (.Y (nx9780), .A (nx10398)) ;
    inv02 ix9781 (.Y (nx9782), .A (nx10398)) ;
    inv02 ix9783 (.Y (nx9784), .A (nx10398)) ;
    inv02 ix9785 (.Y (nx9786), .A (nx10398)) ;
    inv02 ix9787 (.Y (nx9788), .A (nx10398)) ;
    inv02 ix9789 (.Y (nx9790), .A (nx10398)) ;
    inv02 ix9791 (.Y (nx9792), .A (nx10400)) ;
    inv02 ix9793 (.Y (nx9794), .A (nx10400)) ;
    inv02 ix9795 (.Y (nx9796), .A (nx10400)) ;
    inv02 ix9797 (.Y (nx9798), .A (nx10400)) ;
    inv02 ix9799 (.Y (nx9800), .A (nx10400)) ;
    inv02 ix9803 (.Y (nx9804), .A (nx10402)) ;
    inv02 ix9805 (.Y (nx9806), .A (nx10402)) ;
    inv02 ix9807 (.Y (nx9808), .A (nx10402)) ;
    inv02 ix9809 (.Y (nx9810), .A (nx10402)) ;
    inv02 ix9811 (.Y (nx9812), .A (nx10402)) ;
    inv02 ix9813 (.Y (nx9814), .A (nx10402)) ;
    inv02 ix9815 (.Y (nx9816), .A (nx10402)) ;
    inv02 ix9817 (.Y (nx9818), .A (nx10404)) ;
    inv02 ix9819 (.Y (nx9820), .A (nx10404)) ;
    inv02 ix9821 (.Y (nx9822), .A (nx10404)) ;
    inv02 ix9823 (.Y (nx9824), .A (nx10404)) ;
    inv02 ix9825 (.Y (nx9826), .A (nx10404)) ;
    inv02 ix9829 (.Y (nx9830), .A (nx10406)) ;
    inv02 ix9831 (.Y (nx9832), .A (nx10406)) ;
    inv02 ix9833 (.Y (nx9834), .A (nx10406)) ;
    inv02 ix9835 (.Y (nx9836), .A (nx10406)) ;
    inv02 ix9837 (.Y (nx9838), .A (nx10406)) ;
    inv02 ix9839 (.Y (nx9840), .A (nx10406)) ;
    inv02 ix9841 (.Y (nx9842), .A (nx10406)) ;
    inv02 ix9843 (.Y (nx9844), .A (nx10408)) ;
    inv02 ix9845 (.Y (nx9846), .A (nx10408)) ;
    inv02 ix9847 (.Y (nx9848), .A (nx10408)) ;
    inv02 ix9849 (.Y (nx9850), .A (nx10408)) ;
    inv02 ix9851 (.Y (nx9852), .A (nx10408)) ;
    inv02 ix9855 (.Y (nx9856), .A (nx10410)) ;
    inv02 ix9857 (.Y (nx9858), .A (nx10410)) ;
    inv02 ix9859 (.Y (nx9860), .A (nx10410)) ;
    inv02 ix9861 (.Y (nx9862), .A (nx10410)) ;
    inv02 ix9863 (.Y (nx9864), .A (nx10410)) ;
    inv02 ix9865 (.Y (nx9866), .A (nx10410)) ;
    inv02 ix9867 (.Y (nx9868), .A (nx10410)) ;
    inv02 ix9869 (.Y (nx9870), .A (nx10412)) ;
    inv02 ix9871 (.Y (nx9872), .A (nx10412)) ;
    inv02 ix9873 (.Y (nx9874), .A (nx10412)) ;
    inv02 ix9875 (.Y (nx9876), .A (nx10412)) ;
    inv02 ix9877 (.Y (nx9878), .A (nx10412)) ;
    inv02 ix9881 (.Y (nx9882), .A (nx10414)) ;
    inv02 ix9883 (.Y (nx9884), .A (nx10414)) ;
    inv02 ix9885 (.Y (nx9886), .A (nx10414)) ;
    inv02 ix9887 (.Y (nx9888), .A (nx10414)) ;
    inv02 ix9889 (.Y (nx9890), .A (nx10414)) ;
    inv02 ix9891 (.Y (nx9892), .A (nx10414)) ;
    inv02 ix9893 (.Y (nx9894), .A (nx10414)) ;
    inv02 ix9895 (.Y (nx9896), .A (nx10416)) ;
    inv02 ix9897 (.Y (nx9898), .A (nx10416)) ;
    inv02 ix9899 (.Y (nx9900), .A (nx10416)) ;
    inv02 ix9901 (.Y (nx9902), .A (nx10416)) ;
    inv02 ix9903 (.Y (nx9904), .A (nx10416)) ;
    inv02 ix9907 (.Y (nx9908), .A (nx10418)) ;
    inv02 ix9909 (.Y (nx9910), .A (nx10418)) ;
    inv02 ix9911 (.Y (nx9912), .A (nx10418)) ;
    inv02 ix9913 (.Y (nx9914), .A (nx10418)) ;
    inv02 ix9915 (.Y (nx9916), .A (nx10418)) ;
    inv02 ix9917 (.Y (nx9918), .A (nx10418)) ;
    inv02 ix9919 (.Y (nx9920), .A (nx10418)) ;
    inv02 ix9921 (.Y (nx9922), .A (nx10420)) ;
    inv02 ix9923 (.Y (nx9924), .A (nx10420)) ;
    inv02 ix9925 (.Y (nx9926), .A (nx10420)) ;
    inv02 ix9927 (.Y (nx9928), .A (nx10420)) ;
    inv02 ix9929 (.Y (nx9930), .A (nx10420)) ;
    inv02 ix9933 (.Y (nx9934), .A (nx10422)) ;
    inv02 ix9935 (.Y (nx9936), .A (nx10422)) ;
    inv02 ix9937 (.Y (nx9938), .A (nx10422)) ;
    inv02 ix9939 (.Y (nx9940), .A (nx10422)) ;
    inv02 ix9941 (.Y (nx9942), .A (nx10422)) ;
    inv02 ix9943 (.Y (nx9944), .A (nx10422)) ;
    inv02 ix9945 (.Y (nx9946), .A (nx10422)) ;
    inv02 ix9947 (.Y (nx9948), .A (nx10424)) ;
    inv02 ix9949 (.Y (nx9950), .A (nx10424)) ;
    inv02 ix9951 (.Y (nx9952), .A (nx10424)) ;
    inv02 ix9953 (.Y (nx9954), .A (nx10424)) ;
    inv02 ix9955 (.Y (nx9956), .A (nx10424)) ;
    inv02 ix9959 (.Y (nx9960), .A (nx10426)) ;
    inv02 ix9961 (.Y (nx9962), .A (nx10426)) ;
    inv02 ix9963 (.Y (nx9964), .A (nx10426)) ;
    inv02 ix9965 (.Y (nx9966), .A (nx10426)) ;
    inv02 ix9967 (.Y (nx9968), .A (nx10426)) ;
    inv02 ix9969 (.Y (nx9970), .A (nx10426)) ;
    inv02 ix9971 (.Y (nx9972), .A (nx10426)) ;
    inv02 ix9973 (.Y (nx9974), .A (nx10428)) ;
    inv02 ix9975 (.Y (nx9976), .A (nx10428)) ;
    inv02 ix9977 (.Y (nx9978), .A (nx10428)) ;
    inv02 ix9979 (.Y (nx9980), .A (nx10428)) ;
    inv02 ix9981 (.Y (nx9982), .A (nx10428)) ;
    inv02 ix9985 (.Y (nx9986), .A (nx10430)) ;
    inv02 ix9987 (.Y (nx9988), .A (nx10430)) ;
    inv02 ix9989 (.Y (nx9990), .A (nx10430)) ;
    inv02 ix9991 (.Y (nx9992), .A (nx10430)) ;
    inv02 ix9993 (.Y (nx9994), .A (nx10430)) ;
    inv02 ix9995 (.Y (nx9996), .A (nx10430)) ;
    inv02 ix9997 (.Y (nx9998), .A (nx10430)) ;
    inv02 ix9999 (.Y (nx10000), .A (nx10432)) ;
    inv02 ix10001 (.Y (nx10002), .A (nx10432)) ;
    inv02 ix10003 (.Y (nx10004), .A (nx10432)) ;
    inv02 ix10005 (.Y (nx10006), .A (nx10432)) ;
    inv02 ix10007 (.Y (nx10008), .A (nx10432)) ;
    inv02 ix10011 (.Y (nx10012), .A (nx10434)) ;
    inv02 ix10013 (.Y (nx10014), .A (nx10434)) ;
    inv02 ix10015 (.Y (nx10016), .A (nx10434)) ;
    inv02 ix10017 (.Y (nx10018), .A (nx10434)) ;
    inv02 ix10019 (.Y (nx10020), .A (nx10434)) ;
    inv02 ix10021 (.Y (nx10022), .A (nx10434)) ;
    inv02 ix10023 (.Y (nx10024), .A (nx10434)) ;
    inv02 ix10025 (.Y (nx10026), .A (nx10436)) ;
    inv02 ix10027 (.Y (nx10028), .A (nx10436)) ;
    inv02 ix10029 (.Y (nx10030), .A (nx10436)) ;
    inv02 ix10031 (.Y (nx10032), .A (nx10436)) ;
    inv02 ix10033 (.Y (nx10034), .A (nx10436)) ;
    inv02 ix10037 (.Y (nx10038), .A (nx10438)) ;
    inv02 ix10039 (.Y (nx10040), .A (nx10438)) ;
    inv02 ix10041 (.Y (nx10042), .A (nx10438)) ;
    inv02 ix10043 (.Y (nx10044), .A (nx10438)) ;
    inv02 ix10045 (.Y (nx10046), .A (nx10438)) ;
    inv02 ix10047 (.Y (nx10048), .A (nx10438)) ;
    inv02 ix10049 (.Y (nx10050), .A (nx10438)) ;
    inv02 ix10051 (.Y (nx10052), .A (nx10440)) ;
    inv02 ix10053 (.Y (nx10054), .A (nx10440)) ;
    inv02 ix10055 (.Y (nx10056), .A (nx10440)) ;
    inv02 ix10057 (.Y (nx10058), .A (nx10440)) ;
    inv02 ix10059 (.Y (nx10060), .A (nx10440)) ;
    inv02 ix10063 (.Y (nx10064), .A (nx10442)) ;
    inv02 ix10065 (.Y (nx10066), .A (nx10442)) ;
    inv02 ix10067 (.Y (nx10068), .A (nx10442)) ;
    inv02 ix10069 (.Y (nx10070), .A (nx10442)) ;
    inv02 ix10071 (.Y (nx10072), .A (nx10442)) ;
    inv02 ix10073 (.Y (nx10074), .A (nx10442)) ;
    inv02 ix10075 (.Y (nx10076), .A (nx10442)) ;
    inv02 ix10077 (.Y (nx10078), .A (nx10444)) ;
    inv02 ix10079 (.Y (nx10080), .A (nx10444)) ;
    inv02 ix10081 (.Y (nx10082), .A (nx10444)) ;
    inv02 ix10083 (.Y (nx10084), .A (nx10444)) ;
    inv02 ix10085 (.Y (nx10086), .A (nx10444)) ;
    inv02 ix10089 (.Y (nx10090), .A (nx10446)) ;
    inv02 ix10091 (.Y (nx10092), .A (nx10446)) ;
    inv02 ix10093 (.Y (nx10094), .A (nx10446)) ;
    inv02 ix10095 (.Y (nx10096), .A (nx10446)) ;
    inv02 ix10097 (.Y (nx10098), .A (nx10446)) ;
    inv02 ix10099 (.Y (nx10100), .A (nx10446)) ;
    inv02 ix10101 (.Y (nx10102), .A (nx10446)) ;
    inv02 ix10103 (.Y (nx10104), .A (nx10448)) ;
    inv02 ix10105 (.Y (nx10106), .A (nx10448)) ;
    inv02 ix10107 (.Y (nx10108), .A (nx10448)) ;
    inv02 ix10109 (.Y (nx10110), .A (nx10448)) ;
    inv02 ix10111 (.Y (nx10112), .A (nx10448)) ;
    inv02 ix10115 (.Y (nx10116), .A (nx10450)) ;
    inv02 ix10117 (.Y (nx10118), .A (nx10450)) ;
    inv02 ix10119 (.Y (nx10120), .A (nx10450)) ;
    inv02 ix10121 (.Y (nx10122), .A (nx10450)) ;
    inv02 ix10123 (.Y (nx10124), .A (nx10450)) ;
    inv02 ix10125 (.Y (nx10126), .A (nx10450)) ;
    inv02 ix10127 (.Y (nx10128), .A (nx10450)) ;
    inv02 ix10129 (.Y (nx10130), .A (nx10452)) ;
    inv02 ix10131 (.Y (nx10132), .A (nx10452)) ;
    inv02 ix10133 (.Y (nx10134), .A (nx10452)) ;
    inv02 ix10135 (.Y (nx10136), .A (nx10452)) ;
    inv02 ix10137 (.Y (nx10138), .A (nx10452)) ;
    inv02 ix10141 (.Y (nx10142), .A (nx10454)) ;
    inv02 ix10143 (.Y (nx10144), .A (nx10454)) ;
    inv02 ix10145 (.Y (nx10146), .A (nx10454)) ;
    inv02 ix10147 (.Y (nx10148), .A (nx10454)) ;
    inv02 ix10149 (.Y (nx10150), .A (nx10454)) ;
    inv02 ix10151 (.Y (nx10152), .A (nx10454)) ;
    inv02 ix10153 (.Y (nx10154), .A (nx10454)) ;
    inv02 ix10155 (.Y (nx10156), .A (nx10456)) ;
    inv02 ix10157 (.Y (nx10158), .A (nx10456)) ;
    inv02 ix10159 (.Y (nx10160), .A (nx10456)) ;
    inv02 ix10161 (.Y (nx10162), .A (nx10456)) ;
    inv02 ix10163 (.Y (nx10164), .A (nx10456)) ;
    inv02 ix10167 (.Y (nx10168), .A (nx10458)) ;
    inv02 ix10169 (.Y (nx10170), .A (nx10458)) ;
    inv02 ix10171 (.Y (nx10172), .A (nx10458)) ;
    inv02 ix10173 (.Y (nx10174), .A (nx10458)) ;
    inv02 ix10175 (.Y (nx10176), .A (nx10458)) ;
    inv02 ix10177 (.Y (nx10178), .A (nx10458)) ;
    inv02 ix10179 (.Y (nx10180), .A (nx10458)) ;
    inv02 ix10181 (.Y (nx10182), .A (nx10460)) ;
    inv02 ix10183 (.Y (nx10184), .A (nx10460)) ;
    inv02 ix10185 (.Y (nx10186), .A (nx10460)) ;
    inv02 ix10187 (.Y (nx10188), .A (nx10460)) ;
    inv02 ix10189 (.Y (nx10190), .A (nx10460)) ;
    inv02 ix10193 (.Y (nx10194), .A (nx10462)) ;
    inv02 ix10195 (.Y (nx10196), .A (nx10462)) ;
    inv02 ix10197 (.Y (nx10198), .A (nx10462)) ;
    inv02 ix10199 (.Y (nx10200), .A (nx10462)) ;
    inv02 ix10201 (.Y (nx10202), .A (nx10462)) ;
    inv02 ix10203 (.Y (nx10204), .A (nx10462)) ;
    inv02 ix10205 (.Y (nx10206), .A (nx10462)) ;
    inv02 ix10207 (.Y (nx10208), .A (nx10464)) ;
    inv02 ix10209 (.Y (nx10210), .A (nx10464)) ;
    inv02 ix10211 (.Y (nx10212), .A (nx10464)) ;
    inv02 ix10213 (.Y (nx10214), .A (nx10464)) ;
    inv02 ix10215 (.Y (nx10216), .A (nx10464)) ;
    inv02 ix10219 (.Y (nx10220), .A (nx10466)) ;
    inv02 ix10221 (.Y (nx10222), .A (nx10466)) ;
    inv02 ix10223 (.Y (nx10224), .A (nx10466)) ;
    inv02 ix10225 (.Y (nx10226), .A (nx10466)) ;
    inv02 ix10227 (.Y (nx10228), .A (nx10466)) ;
    inv02 ix10229 (.Y (nx10230), .A (nx10466)) ;
    inv02 ix10231 (.Y (nx10232), .A (nx10466)) ;
    inv02 ix10233 (.Y (nx10234), .A (nx10468)) ;
    inv02 ix10235 (.Y (nx10236), .A (nx10468)) ;
    inv02 ix10237 (.Y (nx10238), .A (nx10468)) ;
    inv02 ix10239 (.Y (nx10240), .A (nx10468)) ;
    inv02 ix10241 (.Y (nx10242), .A (nx10468)) ;
    inv02 ix10245 (.Y (nx10246), .A (nx10470)) ;
    inv02 ix10247 (.Y (nx10248), .A (nx10470)) ;
    inv02 ix10249 (.Y (nx10250), .A (nx10470)) ;
    inv02 ix10251 (.Y (nx10252), .A (nx10470)) ;
    inv02 ix10253 (.Y (nx10254), .A (nx10470)) ;
    inv02 ix10255 (.Y (nx10256), .A (nx10470)) ;
    inv02 ix10257 (.Y (nx10258), .A (nx10470)) ;
    inv02 ix10259 (.Y (nx10260), .A (nx10472)) ;
    inv02 ix10261 (.Y (nx10262), .A (nx10472)) ;
    inv02 ix10263 (.Y (nx10264), .A (nx10472)) ;
    inv02 ix10265 (.Y (nx10266), .A (nx10472)) ;
    inv02 ix10267 (.Y (nx10268), .A (nx10472)) ;
    inv02 ix10271 (.Y (nx10272), .A (nx10474)) ;
    inv02 ix10273 (.Y (nx10274), .A (nx10474)) ;
    inv02 ix10275 (.Y (nx10276), .A (nx10474)) ;
    inv02 ix10277 (.Y (nx10278), .A (nx10474)) ;
    inv02 ix10279 (.Y (nx10280), .A (nx10474)) ;
    inv02 ix10281 (.Y (nx10282), .A (nx10474)) ;
    inv02 ix10283 (.Y (nx10284), .A (nx10474)) ;
    inv02 ix10285 (.Y (nx10286), .A (nx10476)) ;
    inv02 ix10287 (.Y (nx10288), .A (nx10476)) ;
    inv02 ix10289 (.Y (nx10290), .A (nx10476)) ;
    inv02 ix10291 (.Y (nx10292), .A (nx10476)) ;
    inv02 ix10293 (.Y (nx10294), .A (nx10476)) ;
    inv02 ix10297 (.Y (nx10298), .A (nx10478)) ;
    inv02 ix10299 (.Y (nx10300), .A (nx10478)) ;
    inv02 ix10301 (.Y (nx10302), .A (nx10478)) ;
    inv02 ix10303 (.Y (nx10304), .A (nx10478)) ;
    inv02 ix10305 (.Y (nx10306), .A (nx10478)) ;
    inv02 ix10307 (.Y (nx10308), .A (nx10478)) ;
    inv02 ix10309 (.Y (nx10310), .A (nx10478)) ;
    inv02 ix10311 (.Y (nx10312), .A (nx10480)) ;
    inv02 ix10313 (.Y (nx10314), .A (nx10480)) ;
    inv02 ix10315 (.Y (nx10316), .A (nx10480)) ;
    inv02 ix10317 (.Y (nx10318), .A (nx10480)) ;
    inv02 ix10319 (.Y (nx10320), .A (nx10480)) ;
    inv02 ix10323 (.Y (nx10324), .A (nx10482)) ;
    inv02 ix10325 (.Y (nx10326), .A (nx10482)) ;
    inv02 ix10327 (.Y (nx10328), .A (nx10482)) ;
    inv02 ix10329 (.Y (nx10330), .A (nx10482)) ;
    inv02 ix10331 (.Y (nx10332), .A (nx10482)) ;
    inv02 ix10333 (.Y (nx10334), .A (nx10482)) ;
    inv02 ix10335 (.Y (nx10336), .A (nx10482)) ;
    inv02 ix10337 (.Y (nx10338), .A (nx10484)) ;
    inv02 ix10339 (.Y (nx10340), .A (nx10484)) ;
    inv02 ix10341 (.Y (nx10342), .A (nx10484)) ;
    inv02 ix10343 (.Y (nx10344), .A (nx10484)) ;
    inv02 ix10345 (.Y (nx10346), .A (nx10484)) ;
    inv02 ix10349 (.Y (nx10350), .A (nx10486)) ;
    inv02 ix10351 (.Y (nx10352), .A (nx10486)) ;
    inv02 ix10353 (.Y (nx10354), .A (nx10486)) ;
    inv02 ix10355 (.Y (nx10356), .A (nx10486)) ;
    inv02 ix10357 (.Y (nx10358), .A (nx10486)) ;
    inv02 ix10359 (.Y (nx10360), .A (nx10486)) ;
    inv02 ix10361 (.Y (nx10362), .A (nx10486)) ;
    inv02 ix10363 (.Y (nx10364), .A (nx10488)) ;
    inv02 ix10365 (.Y (nx10366), .A (nx10488)) ;
    inv02 ix10367 (.Y (nx10368), .A (nx10488)) ;
    inv02 ix10369 (.Y (nx10370), .A (nx10488)) ;
    inv02 ix10371 (.Y (nx10372), .A (nx10488)) ;
    buf02 ix10373 (.Y (nx10374), .A (nx6955)) ;
    buf02 ix10375 (.Y (nx10376), .A (nx6955)) ;
    inv02 ix10377 (.Y (nx10378), .A (nx14)) ;
    inv02 ix10379 (.Y (nx10380), .A (nx14)) ;
    inv02 ix10381 (.Y (nx10382), .A (nx30)) ;
    inv02 ix10383 (.Y (nx10384), .A (nx30)) ;
    inv02 ix10385 (.Y (nx10386), .A (nx42)) ;
    inv02 ix10387 (.Y (nx10388), .A (nx42)) ;
    inv02 ix10389 (.Y (nx10390), .A (nx48)) ;
    inv02 ix10391 (.Y (nx10392), .A (nx48)) ;
    inv02 ix10393 (.Y (nx10394), .A (nx64)) ;
    inv02 ix10395 (.Y (nx10396), .A (nx64)) ;
    inv02 ix10397 (.Y (nx10398), .A (nx68)) ;
    inv02 ix10399 (.Y (nx10400), .A (nx68)) ;
    inv02 ix10401 (.Y (nx10402), .A (nx74)) ;
    inv02 ix10403 (.Y (nx10404), .A (nx74)) ;
    inv02 ix10405 (.Y (nx10406), .A (nx90)) ;
    inv02 ix10407 (.Y (nx10408), .A (nx90)) ;
    inv02 ix10409 (.Y (nx10410), .A (nx94)) ;
    inv02 ix10411 (.Y (nx10412), .A (nx94)) ;
    inv02 ix10413 (.Y (nx10414), .A (nx100)) ;
    inv02 ix10415 (.Y (nx10416), .A (nx100)) ;
    inv02 ix10417 (.Y (nx10418), .A (nx104)) ;
    inv02 ix10419 (.Y (nx10420), .A (nx104)) ;
    inv02 ix10421 (.Y (nx10422), .A (nx114)) ;
    inv02 ix10423 (.Y (nx10424), .A (nx114)) ;
    inv02 ix10425 (.Y (nx10426), .A (nx118)) ;
    inv02 ix10427 (.Y (nx10428), .A (nx118)) ;
    inv02 ix10429 (.Y (nx10430), .A (nx122)) ;
    inv02 ix10431 (.Y (nx10432), .A (nx122)) ;
    inv02 ix10433 (.Y (nx10434), .A (nx136)) ;
    inv02 ix10435 (.Y (nx10436), .A (nx136)) ;
    inv02 ix10437 (.Y (nx10438), .A (nx144)) ;
    inv02 ix10439 (.Y (nx10440), .A (nx144)) ;
    inv02 ix10441 (.Y (nx10442), .A (nx150)) ;
    inv02 ix10443 (.Y (nx10444), .A (nx150)) ;
    inv02 ix10445 (.Y (nx10446), .A (nx158)) ;
    inv02 ix10447 (.Y (nx10448), .A (nx158)) ;
    inv02 ix10449 (.Y (nx10450), .A (nx166)) ;
    inv02 ix10451 (.Y (nx10452), .A (nx166)) ;
    inv02 ix10453 (.Y (nx10454), .A (nx172)) ;
    inv02 ix10455 (.Y (nx10456), .A (nx172)) ;
    inv02 ix10457 (.Y (nx10458), .A (nx180)) ;
    inv02 ix10459 (.Y (nx10460), .A (nx180)) ;
    inv02 ix10461 (.Y (nx10462), .A (nx192)) ;
    inv02 ix10463 (.Y (nx10464), .A (nx192)) ;
    inv02 ix10465 (.Y (nx10466), .A (nx200)) ;
    inv02 ix10467 (.Y (nx10468), .A (nx200)) ;
    inv02 ix10469 (.Y (nx10470), .A (nx206)) ;
    inv02 ix10471 (.Y (nx10472), .A (nx206)) ;
    inv02 ix10473 (.Y (nx10474), .A (nx214)) ;
    inv02 ix10475 (.Y (nx10476), .A (nx214)) ;
    inv02 ix10477 (.Y (nx10478), .A (nx222)) ;
    inv02 ix10479 (.Y (nx10480), .A (nx222)) ;
    inv02 ix10481 (.Y (nx10482), .A (nx226)) ;
    inv02 ix10483 (.Y (nx10484), .A (nx226)) ;
    inv02 ix10485 (.Y (nx10486), .A (nx230)) ;
    inv02 ix10487 (.Y (nx10488), .A (nx230)) ;
    nor02ii ix8951 (.Y (sel_que_0), .A0 (nx6829), .A1 (nx6885)) ;
    nor02ii ix8961 (.Y (sel_que_1), .A0 (nx6839), .A1 (nx6885)) ;
    nor02ii ix8971 (.Y (sel_que_2), .A0 (nx6843), .A1 (nx6885)) ;
    nor02ii ix8979 (.Y (sel_que_3), .A0 (nx6847), .A1 (nx6885)) ;
    nor02ii ix8987 (.Y (sel_que_4), .A0 (nx6829), .A1 (nx6905)) ;
    nor02ii ix8991 (.Y (sel_que_5), .A0 (nx6839), .A1 (nx6905)) ;
    nor02ii ix8995 (.Y (sel_que_6), .A0 (nx6843), .A1 (nx6905)) ;
    nor02ii ix8999 (.Y (sel_que_7), .A0 (nx6847), .A1 (nx6905)) ;
    nor02ii ix9007 (.Y (sel_que_8), .A0 (nx6829), .A1 (nx6915)) ;
    nor02ii ix9011 (.Y (sel_que_9), .A0 (nx6839), .A1 (nx6915)) ;
    nor02ii ix9015 (.Y (sel_que_10), .A0 (nx6843), .A1 (nx6915)) ;
    nor02ii ix9019 (.Y (sel_que_11), .A0 (nx6847), .A1 (nx6915)) ;
    nor02ii ix9053 (.Y (sel_que_17), .A0 (nx6893), .A1 (nx6885)) ;
    nor02ii ix9063 (.Y (sel_que_18), .A0 (nx6897), .A1 (nx6885)) ;
    nor02ii ix9071 (.Y (sel_que_19), .A0 (nx6901), .A1 (nx6885)) ;
    nor02ii ix6906 (.Y (nx6905), .A0 (cache_in_sel[3]), .A1 (cache_in_sel[2])) ;
    nor02ii ix9079 (.Y (sel_que_21), .A0 (nx6893), .A1 (nx6905)) ;
    nor02ii ix9083 (.Y (sel_que_22), .A0 (nx6897), .A1 (nx6905)) ;
    nor02ii ix9087 (.Y (sel_que_23), .A0 (nx6901), .A1 (nx6905)) ;
    nor02ii ix6916 (.Y (nx6915), .A0 (cache_in_sel[2]), .A1 (cache_in_sel[3])) ;
    nor02ii ix9095 (.Y (sel_que_25), .A0 (nx6893), .A1 (nx6915)) ;
    nor02ii ix9099 (.Y (sel_que_26), .A0 (nx6897), .A1 (nx6915)) ;
    nor02ii ix9103 (.Y (sel_que_27), .A0 (nx6901), .A1 (nx6915)) ;
    nor02ii ix223 (.Y (nx222), .A0 (nx6931), .A1 (nx62)) ;
    nor02ii ix231 (.Y (nx230), .A0 (nx6945), .A1 (nx88)) ;
    nor02ii ix207 (.Y (nx206), .A0 (nx10374), .A1 (nx28)) ;
    nor02ii ix123 (.Y (nx122), .A0 (nx10374), .A1 (nx62)) ;
    nor02ii ix65 (.Y (nx64), .A0 (nx6949), .A1 (nx62)) ;
    nor02ii ix49 (.Y (nx48), .A0 (nx6949), .A1 (nx28)) ;
    nor02ii ix31 (.Y (nx30), .A0 (nx6931), .A1 (nx28)) ;
    inv02 ix10493 (.Y (nx10494), .A (nx6937)) ;
    inv02 ix10495 (.Y (nx10496), .A (nx6937)) ;
    inv02 ix10497 (.Y (nx10498), .A (nx6939)) ;
    inv02 ix10499 (.Y (nx10500), .A (nx6939)) ;
    inv01 ix10501 (.Y (nx10502), .A (nx6961)) ;
    inv01 ix10503 (.Y (nx10504), .A (nx6961)) ;
    inv02 ix10505 (.Y (nx10506), .A (nx6833)) ;
    inv02 ix10507 (.Y (nx10508), .A (nx6835)) ;
    inv01 ix10509 (.Y (nx10510), .A (in_word[15])) ;
    inv01 ix10511 (.Y (nx10512), .A (nx10510)) ;
    inv01 ix10513 (.Y (nx10514), .A (nx10510)) ;
    inv01 ix10515 (.Y (nx10516), .A (nx10510)) ;
    inv01 ix10517 (.Y (nx10518), .A (nx10510)) ;
    inv01 ix10519 (.Y (nx10520), .A (in_word[14])) ;
    inv01 ix10521 (.Y (nx10522), .A (nx10520)) ;
    inv01 ix10523 (.Y (nx10524), .A (nx10520)) ;
    inv01 ix10525 (.Y (nx10526), .A (nx10520)) ;
    inv01 ix10527 (.Y (nx10528), .A (nx10520)) ;
    inv01 ix10529 (.Y (nx10530), .A (in_word[13])) ;
    inv01 ix10531 (.Y (nx10532), .A (nx10530)) ;
    inv01 ix10533 (.Y (nx10534), .A (nx10530)) ;
    inv01 ix10535 (.Y (nx10536), .A (nx10530)) ;
    inv01 ix10537 (.Y (nx10538), .A (nx10530)) ;
    inv01 ix10539 (.Y (nx10540), .A (in_word[12])) ;
    inv01 ix10541 (.Y (nx10542), .A (nx10540)) ;
    inv01 ix10543 (.Y (nx10544), .A (nx10540)) ;
    inv01 ix10545 (.Y (nx10546), .A (nx10540)) ;
    inv01 ix10547 (.Y (nx10548), .A (nx10540)) ;
    inv01 ix10549 (.Y (nx10550), .A (in_word[11])) ;
    inv01 ix10551 (.Y (nx10552), .A (nx10550)) ;
    inv01 ix10553 (.Y (nx10554), .A (nx10550)) ;
    inv01 ix10555 (.Y (nx10556), .A (nx10550)) ;
    inv01 ix10557 (.Y (nx10558), .A (nx10550)) ;
    inv01 ix10559 (.Y (nx10560), .A (in_word[10])) ;
    inv01 ix10561 (.Y (nx10562), .A (nx10560)) ;
    inv01 ix10563 (.Y (nx10564), .A (nx10560)) ;
    inv01 ix10565 (.Y (nx10566), .A (nx10560)) ;
    inv01 ix10567 (.Y (nx10568), .A (nx10560)) ;
    inv01 ix10569 (.Y (nx10570), .A (in_word[9])) ;
    inv01 ix10571 (.Y (nx10572), .A (nx10570)) ;
    inv01 ix10573 (.Y (nx10574), .A (nx10570)) ;
    inv01 ix10575 (.Y (nx10576), .A (nx10570)) ;
    inv01 ix10577 (.Y (nx10578), .A (nx10570)) ;
    inv01 ix10579 (.Y (nx10580), .A (in_word[8])) ;
    inv01 ix10581 (.Y (nx10582), .A (nx10580)) ;
    inv01 ix10583 (.Y (nx10584), .A (nx10580)) ;
    inv01 ix10585 (.Y (nx10586), .A (nx10580)) ;
    inv01 ix10587 (.Y (nx10588), .A (nx10580)) ;
    inv01 ix10589 (.Y (nx10590), .A (in_word[7])) ;
    inv01 ix10591 (.Y (nx10592), .A (nx10590)) ;
    inv01 ix10593 (.Y (nx10594), .A (nx10590)) ;
    inv01 ix10595 (.Y (nx10596), .A (nx10590)) ;
    inv01 ix10597 (.Y (nx10598), .A (nx10590)) ;
    inv01 ix10599 (.Y (nx10600), .A (in_word[6])) ;
    inv01 ix10601 (.Y (nx10602), .A (nx10600)) ;
    inv01 ix10603 (.Y (nx10604), .A (nx10600)) ;
    inv01 ix10605 (.Y (nx10606), .A (nx10600)) ;
    inv01 ix10607 (.Y (nx10608), .A (nx10600)) ;
    inv01 ix10609 (.Y (nx10610), .A (in_word[5])) ;
    inv01 ix10611 (.Y (nx10612), .A (nx10610)) ;
    inv01 ix10613 (.Y (nx10614), .A (nx10610)) ;
    inv01 ix10615 (.Y (nx10616), .A (nx10610)) ;
    inv01 ix10617 (.Y (nx10618), .A (nx10610)) ;
    inv01 ix10619 (.Y (nx10620), .A (in_word[4])) ;
    inv01 ix10621 (.Y (nx10622), .A (nx10620)) ;
    inv01 ix10623 (.Y (nx10624), .A (nx10620)) ;
    inv01 ix10625 (.Y (nx10626), .A (nx10620)) ;
    inv01 ix10627 (.Y (nx10628), .A (nx10620)) ;
    inv01 ix10629 (.Y (nx10630), .A (in_word[3])) ;
    inv01 ix10631 (.Y (nx10632), .A (nx10630)) ;
    inv01 ix10633 (.Y (nx10634), .A (nx10630)) ;
    inv01 ix10635 (.Y (nx10636), .A (nx10630)) ;
    inv01 ix10637 (.Y (nx10638), .A (nx10630)) ;
    inv01 ix10639 (.Y (nx10640), .A (in_word[2])) ;
    inv01 ix10641 (.Y (nx10642), .A (nx10640)) ;
    inv01 ix10643 (.Y (nx10644), .A (nx10640)) ;
    inv01 ix10645 (.Y (nx10646), .A (nx10640)) ;
    inv01 ix10647 (.Y (nx10648), .A (nx10640)) ;
    inv01 ix10649 (.Y (nx10650), .A (in_word[1])) ;
    inv01 ix10651 (.Y (nx10652), .A (nx10650)) ;
    inv01 ix10653 (.Y (nx10654), .A (nx10650)) ;
    inv01 ix10655 (.Y (nx10656), .A (nx10650)) ;
    inv01 ix10657 (.Y (nx10658), .A (nx10650)) ;
    inv01 ix10659 (.Y (nx10660), .A (in_word[0])) ;
    inv01 ix10661 (.Y (nx10662), .A (nx10660)) ;
    inv01 ix10663 (.Y (nx10664), .A (nx10660)) ;
    inv01 ix10665 (.Y (nx10666), .A (nx10660)) ;
    inv01 ix10667 (.Y (nx10668), .A (nx10660)) ;
    inv02 ix10689 (.Y (nx10690), .A (nx10742)) ;
    inv02 ix10691 (.Y (nx10692), .A (nx10742)) ;
    inv02 ix10693 (.Y (nx10694), .A (nx10742)) ;
    inv02 ix10695 (.Y (nx10696), .A (nx10742)) ;
    inv02 ix10697 (.Y (nx10698), .A (nx10742)) ;
    inv02 ix10699 (.Y (nx10700), .A (nx10742)) ;
    inv02 ix10701 (.Y (nx10702), .A (nx10742)) ;
    inv02 ix10703 (.Y (nx10704), .A (nx10744)) ;
    inv02 ix10705 (.Y (nx10706), .A (nx10744)) ;
    inv02 ix10707 (.Y (nx10708), .A (nx10744)) ;
    inv02 ix10709 (.Y (nx10710), .A (nx10744)) ;
    inv02 ix10711 (.Y (nx10712), .A (nx10744)) ;
    inv02 ix10713 (.Y (nx10714), .A (nx10746)) ;
    inv02 ix10715 (.Y (nx10716), .A (nx10746)) ;
    inv02 ix10717 (.Y (nx10718), .A (nx10746)) ;
    inv02 ix10719 (.Y (nx10720), .A (nx10746)) ;
    inv02 ix10721 (.Y (nx10722), .A (nx10746)) ;
    inv02 ix10723 (.Y (nx10724), .A (nx10746)) ;
    inv02 ix10725 (.Y (nx10726), .A (nx10746)) ;
    inv02 ix10727 (.Y (nx10728), .A (nx10748)) ;
    inv02 ix10729 (.Y (nx10730), .A (nx10748)) ;
    inv02 ix10731 (.Y (nx10732), .A (nx10748)) ;
    inv02 ix10733 (.Y (nx10734), .A (nx10748)) ;
    inv02 ix10735 (.Y (nx10736), .A (nx10748)) ;
    inv02 ix10741 (.Y (nx10742), .A (reset)) ;
    inv02 ix10743 (.Y (nx10744), .A (reset)) ;
    inv02 ix10745 (.Y (nx10746), .A (clk)) ;
    inv02 ix10747 (.Y (nx10748), .A (clk)) ;
endmodule


module Queue_5 ( d, q_0__15, q_0__14, q_0__13, q_0__12, q_0__11, q_0__10, q_0__9, 
                 q_0__8, q_0__7, q_0__6, q_0__5, q_0__4, q_0__3, q_0__2, q_0__1, 
                 q_0__0, q_1__15, q_1__14, q_1__13, q_1__12, q_1__11, q_1__10, 
                 q_1__9, q_1__8, q_1__7, q_1__6, q_1__5, q_1__4, q_1__3, q_1__2, 
                 q_1__1, q_1__0, q_2__15, q_2__14, q_2__13, q_2__12, q_2__11, 
                 q_2__10, q_2__9, q_2__8, q_2__7, q_2__6, q_2__5, q_2__4, q_2__3, 
                 q_2__2, q_2__1, q_2__0, q_3__15, q_3__14, q_3__13, q_3__12, 
                 q_3__11, q_3__10, q_3__9, q_3__8, q_3__7, q_3__6, q_3__5, 
                 q_3__4, q_3__3, q_3__2, q_3__1, q_3__0, q_4__15, q_4__14, 
                 q_4__13, q_4__12, q_4__11, q_4__10, q_4__9, q_4__8, q_4__7, 
                 q_4__6, q_4__5, q_4__4, q_4__3, q_4__2, q_4__1, q_4__0, clk, 
                 load, reset ) ;

    input [15:0]d ;
    output q_0__15 ;
    output q_0__14 ;
    output q_0__13 ;
    output q_0__12 ;
    output q_0__11 ;
    output q_0__10 ;
    output q_0__9 ;
    output q_0__8 ;
    output q_0__7 ;
    output q_0__6 ;
    output q_0__5 ;
    output q_0__4 ;
    output q_0__3 ;
    output q_0__2 ;
    output q_0__1 ;
    output q_0__0 ;
    output q_1__15 ;
    output q_1__14 ;
    output q_1__13 ;
    output q_1__12 ;
    output q_1__11 ;
    output q_1__10 ;
    output q_1__9 ;
    output q_1__8 ;
    output q_1__7 ;
    output q_1__6 ;
    output q_1__5 ;
    output q_1__4 ;
    output q_1__3 ;
    output q_1__2 ;
    output q_1__1 ;
    output q_1__0 ;
    output q_2__15 ;
    output q_2__14 ;
    output q_2__13 ;
    output q_2__12 ;
    output q_2__11 ;
    output q_2__10 ;
    output q_2__9 ;
    output q_2__8 ;
    output q_2__7 ;
    output q_2__6 ;
    output q_2__5 ;
    output q_2__4 ;
    output q_2__3 ;
    output q_2__2 ;
    output q_2__1 ;
    output q_2__0 ;
    output q_3__15 ;
    output q_3__14 ;
    output q_3__13 ;
    output q_3__12 ;
    output q_3__11 ;
    output q_3__10 ;
    output q_3__9 ;
    output q_3__8 ;
    output q_3__7 ;
    output q_3__6 ;
    output q_3__5 ;
    output q_3__4 ;
    output q_3__3 ;
    output q_3__2 ;
    output q_3__1 ;
    output q_3__0 ;
    output q_4__15 ;
    output q_4__14 ;
    output q_4__13 ;
    output q_4__12 ;
    output q_4__11 ;
    output q_4__10 ;
    output q_4__9 ;
    output q_4__8 ;
    output q_4__7 ;
    output q_4__6 ;
    output q_4__5 ;
    output q_4__4 ;
    output q_4__3 ;
    output q_4__2 ;
    output q_4__1 ;
    output q_4__0 ;
    input clk ;
    input load ;
    input reset ;

    wire nx393, nx403, nx413, nx423, nx433, nx443, nx453, nx463, nx473, nx483, 
         nx493, nx503, nx513, nx523, nx533, nx543, nx553, nx563, nx573, nx583, 
         nx593, nx603, nx613, nx623, nx633, nx643, nx653, nx663, nx673, nx683, 
         nx693, nx703, nx713, nx723, nx733, nx743, nx753, nx763, nx773, nx783, 
         nx793, nx803, nx813, nx823, nx833, nx843, nx853, nx863, nx873, nx883, 
         nx893, nx903, nx913, nx923, nx933, nx943, nx953, nx963, nx973, nx983, 
         nx993, nx1003, nx1013, nx1023, nx1033, nx1043, nx1053, nx1063, nx1073, 
         nx1083, nx1093, nx1103, nx1113, nx1123, nx1133, nx1143, nx1153, nx1163, 
         nx1173, nx1183, nx1440, nx1442, nx1444, nx1446, nx1448, nx1450, nx1452, 
         nx1454, nx1456, nx1458, nx1460, nx1462, nx1466, nx1468, nx1470, nx1472, 
         nx1474, nx1476, nx1478, nx1480, nx1482, nx1484, nx1486, nx1488, nx1492, 
         nx1494, nx1496, nx1498, nx1500, nx1502, nx1504, nx1506, nx1508, nx1510, 
         nx1512, nx1514, nx1516, nx1518, nx1520, nx1522, nx1524, nx1526;
    wire [79:0] \$dummy ;




    dffr gen_regs_4_regi_reg_q_0 (.Q (q_4__0), .QB (\$dummy [0]), .D (nx433), .CLK (
         nx1492), .R (nx1466)) ;
    mux21_ni ix434 (.Y (nx433), .A0 (q_4__0), .A1 (q_3__0), .S0 (nx1440)) ;
    dffr gen_regs_3_regi_reg_q_0 (.Q (q_3__0), .QB (\$dummy [1]), .D (nx423), .CLK (
         nx1492), .R (nx1466)) ;
    mux21_ni ix424 (.Y (nx423), .A0 (q_3__0), .A1 (q_2__0), .S0 (nx1440)) ;
    dffr gen_regs_2_regi_reg_q_0 (.Q (q_2__0), .QB (\$dummy [2]), .D (nx413), .CLK (
         nx1492), .R (nx1466)) ;
    mux21_ni ix414 (.Y (nx413), .A0 (q_2__0), .A1 (q_1__0), .S0 (nx1440)) ;
    dffr gen_regs_1_regi_reg_q_0 (.Q (q_1__0), .QB (\$dummy [3]), .D (nx403), .CLK (
         nx1492), .R (nx1466)) ;
    mux21_ni ix404 (.Y (nx403), .A0 (q_1__0), .A1 (q_0__0), .S0 (nx1440)) ;
    dffr reg0_reg_q_0 (.Q (q_0__0), .QB (\$dummy [4]), .D (nx393), .CLK (nx1492)
         , .R (nx1466)) ;
    mux21_ni ix394 (.Y (nx393), .A0 (q_0__0), .A1 (d[0]), .S0 (nx1440)) ;
    dffr gen_regs_4_regi_reg_q_1 (.Q (q_4__1), .QB (\$dummy [5]), .D (nx483), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix484 (.Y (nx483), .A0 (q_4__1), .A1 (q_3__1), .S0 (nx1442)) ;
    dffr gen_regs_3_regi_reg_q_1 (.Q (q_3__1), .QB (\$dummy [6]), .D (nx473), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix474 (.Y (nx473), .A0 (q_3__1), .A1 (q_2__1), .S0 (nx1442)) ;
    dffr gen_regs_2_regi_reg_q_1 (.Q (q_2__1), .QB (\$dummy [7]), .D (nx463), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix464 (.Y (nx463), .A0 (q_2__1), .A1 (q_1__1), .S0 (nx1442)) ;
    dffr gen_regs_1_regi_reg_q_1 (.Q (q_1__1), .QB (\$dummy [8]), .D (nx453), .CLK (
         nx1492), .R (nx1466)) ;
    mux21_ni ix454 (.Y (nx453), .A0 (q_1__1), .A1 (q_0__1), .S0 (nx1440)) ;
    dffr reg0_reg_q_1 (.Q (q_0__1), .QB (\$dummy [9]), .D (nx443), .CLK (nx1492)
         , .R (nx1466)) ;
    mux21_ni ix444 (.Y (nx443), .A0 (q_0__1), .A1 (d[1]), .S0 (nx1440)) ;
    dffr gen_regs_4_regi_reg_q_2 (.Q (q_4__2), .QB (\$dummy [10]), .D (nx533), .CLK (
         nx1496), .R (nx1470)) ;
    mux21_ni ix534 (.Y (nx533), .A0 (q_4__2), .A1 (q_3__2), .S0 (nx1444)) ;
    dffr gen_regs_3_regi_reg_q_2 (.Q (q_3__2), .QB (\$dummy [11]), .D (nx523), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix524 (.Y (nx523), .A0 (q_3__2), .A1 (q_2__2), .S0 (nx1442)) ;
    dffr gen_regs_2_regi_reg_q_2 (.Q (q_2__2), .QB (\$dummy [12]), .D (nx513), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix514 (.Y (nx513), .A0 (q_2__2), .A1 (q_1__2), .S0 (nx1442)) ;
    dffr gen_regs_1_regi_reg_q_2 (.Q (q_1__2), .QB (\$dummy [13]), .D (nx503), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix504 (.Y (nx503), .A0 (q_1__2), .A1 (q_0__2), .S0 (nx1442)) ;
    dffr reg0_reg_q_2 (.Q (q_0__2), .QB (\$dummy [14]), .D (nx493), .CLK (nx1494
         ), .R (nx1468)) ;
    mux21_ni ix494 (.Y (nx493), .A0 (q_0__2), .A1 (d[2]), .S0 (nx1442)) ;
    dffr gen_regs_4_regi_reg_q_3 (.Q (q_4__3), .QB (\$dummy [15]), .D (nx583), .CLK (
         nx1496), .R (nx1470)) ;
    mux21_ni ix584 (.Y (nx583), .A0 (q_4__3), .A1 (q_3__3), .S0 (nx1444)) ;
    dffr gen_regs_3_regi_reg_q_3 (.Q (q_3__3), .QB (\$dummy [16]), .D (nx573), .CLK (
         nx1496), .R (nx1470)) ;
    mux21_ni ix574 (.Y (nx573), .A0 (q_3__3), .A1 (q_2__3), .S0 (nx1444)) ;
    dffr gen_regs_2_regi_reg_q_3 (.Q (q_2__3), .QB (\$dummy [17]), .D (nx563), .CLK (
         nx1496), .R (nx1470)) ;
    mux21_ni ix564 (.Y (nx563), .A0 (q_2__3), .A1 (q_1__3), .S0 (nx1444)) ;
    dffr gen_regs_1_regi_reg_q_3 (.Q (q_1__3), .QB (\$dummy [18]), .D (nx553), .CLK (
         nx1496), .R (nx1470)) ;
    mux21_ni ix554 (.Y (nx553), .A0 (q_1__3), .A1 (q_0__3), .S0 (nx1444)) ;
    dffr reg0_reg_q_3 (.Q (q_0__3), .QB (\$dummy [19]), .D (nx543), .CLK (nx1496
         ), .R (nx1470)) ;
    mux21_ni ix544 (.Y (nx543), .A0 (q_0__3), .A1 (d[3]), .S0 (nx1444)) ;
    dffr gen_regs_4_regi_reg_q_4 (.Q (q_4__4), .QB (\$dummy [20]), .D (nx633), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix634 (.Y (nx633), .A0 (q_4__4), .A1 (q_3__4), .S0 (nx1446)) ;
    dffr gen_regs_3_regi_reg_q_4 (.Q (q_3__4), .QB (\$dummy [21]), .D (nx623), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix624 (.Y (nx623), .A0 (q_3__4), .A1 (q_2__4), .S0 (nx1446)) ;
    dffr gen_regs_2_regi_reg_q_4 (.Q (q_2__4), .QB (\$dummy [22]), .D (nx613), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix614 (.Y (nx613), .A0 (q_2__4), .A1 (q_1__4), .S0 (nx1446)) ;
    dffr gen_regs_1_regi_reg_q_4 (.Q (q_1__4), .QB (\$dummy [23]), .D (nx603), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix604 (.Y (nx603), .A0 (q_1__4), .A1 (q_0__4), .S0 (nx1446)) ;
    dffr reg0_reg_q_4 (.Q (q_0__4), .QB (\$dummy [24]), .D (nx593), .CLK (nx1496
         ), .R (nx1470)) ;
    mux21_ni ix594 (.Y (nx593), .A0 (q_0__4), .A1 (d[4]), .S0 (nx1444)) ;
    dffr gen_regs_4_regi_reg_q_5 (.Q (q_4__5), .QB (\$dummy [25]), .D (nx683), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix684 (.Y (nx683), .A0 (q_4__5), .A1 (q_3__5), .S0 (nx1448)) ;
    dffr gen_regs_3_regi_reg_q_5 (.Q (q_3__5), .QB (\$dummy [26]), .D (nx673), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix674 (.Y (nx673), .A0 (q_3__5), .A1 (q_2__5), .S0 (nx1448)) ;
    dffr gen_regs_2_regi_reg_q_5 (.Q (q_2__5), .QB (\$dummy [27]), .D (nx663), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix664 (.Y (nx663), .A0 (q_2__5), .A1 (q_1__5), .S0 (nx1446)) ;
    dffr gen_regs_1_regi_reg_q_5 (.Q (q_1__5), .QB (\$dummy [28]), .D (nx653), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix654 (.Y (nx653), .A0 (q_1__5), .A1 (q_0__5), .S0 (nx1446)) ;
    dffr reg0_reg_q_5 (.Q (q_0__5), .QB (\$dummy [29]), .D (nx643), .CLK (nx1498
         ), .R (nx1472)) ;
    mux21_ni ix644 (.Y (nx643), .A0 (q_0__5), .A1 (d[5]), .S0 (nx1446)) ;
    dffr gen_regs_4_regi_reg_q_6 (.Q (q_4__6), .QB (\$dummy [30]), .D (nx733), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix734 (.Y (nx733), .A0 (q_4__6), .A1 (q_3__6), .S0 (nx1448)) ;
    dffr gen_regs_3_regi_reg_q_6 (.Q (q_3__6), .QB (\$dummy [31]), .D (nx723), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix724 (.Y (nx723), .A0 (q_3__6), .A1 (q_2__6), .S0 (nx1448)) ;
    dffr gen_regs_2_regi_reg_q_6 (.Q (q_2__6), .QB (\$dummy [32]), .D (nx713), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix714 (.Y (nx713), .A0 (q_2__6), .A1 (q_1__6), .S0 (nx1448)) ;
    dffr gen_regs_1_regi_reg_q_6 (.Q (q_1__6), .QB (\$dummy [33]), .D (nx703), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix704 (.Y (nx703), .A0 (q_1__6), .A1 (q_0__6), .S0 (nx1448)) ;
    dffr reg0_reg_q_6 (.Q (q_0__6), .QB (\$dummy [34]), .D (nx693), .CLK (nx1500
         ), .R (nx1474)) ;
    mux21_ni ix694 (.Y (nx693), .A0 (q_0__6), .A1 (d[6]), .S0 (nx1448)) ;
    dffr gen_regs_4_regi_reg_q_7 (.Q (q_4__7), .QB (\$dummy [35]), .D (nx783), .CLK (
         nx1502), .R (nx1476)) ;
    mux21_ni ix784 (.Y (nx783), .A0 (q_4__7), .A1 (q_3__7), .S0 (nx1450)) ;
    dffr gen_regs_3_regi_reg_q_7 (.Q (q_3__7), .QB (\$dummy [36]), .D (nx773), .CLK (
         nx1502), .R (nx1476)) ;
    mux21_ni ix774 (.Y (nx773), .A0 (q_3__7), .A1 (q_2__7), .S0 (nx1450)) ;
    dffr gen_regs_2_regi_reg_q_7 (.Q (q_2__7), .QB (\$dummy [37]), .D (nx763), .CLK (
         nx1502), .R (nx1476)) ;
    mux21_ni ix764 (.Y (nx763), .A0 (q_2__7), .A1 (q_1__7), .S0 (nx1450)) ;
    dffr gen_regs_1_regi_reg_q_7 (.Q (q_1__7), .QB (\$dummy [38]), .D (nx753), .CLK (
         nx1502), .R (nx1476)) ;
    mux21_ni ix754 (.Y (nx753), .A0 (q_1__7), .A1 (q_0__7), .S0 (nx1450)) ;
    dffr reg0_reg_q_7 (.Q (q_0__7), .QB (\$dummy [39]), .D (nx743), .CLK (nx1502
         ), .R (nx1476)) ;
    mux21_ni ix744 (.Y (nx743), .A0 (q_0__7), .A1 (d[7]), .S0 (nx1450)) ;
    dffr gen_regs_4_regi_reg_q_8 (.Q (q_4__8), .QB (\$dummy [40]), .D (nx833), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix834 (.Y (nx833), .A0 (q_4__8), .A1 (q_3__8), .S0 (nx1452)) ;
    dffr gen_regs_3_regi_reg_q_8 (.Q (q_3__8), .QB (\$dummy [41]), .D (nx823), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix824 (.Y (nx823), .A0 (q_3__8), .A1 (q_2__8), .S0 (nx1452)) ;
    dffr gen_regs_2_regi_reg_q_8 (.Q (q_2__8), .QB (\$dummy [42]), .D (nx813), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix814 (.Y (nx813), .A0 (q_2__8), .A1 (q_1__8), .S0 (nx1452)) ;
    dffr gen_regs_1_regi_reg_q_8 (.Q (q_1__8), .QB (\$dummy [43]), .D (nx803), .CLK (
         nx1502), .R (nx1476)) ;
    mux21_ni ix804 (.Y (nx803), .A0 (q_1__8), .A1 (q_0__8), .S0 (nx1450)) ;
    dffr reg0_reg_q_8 (.Q (q_0__8), .QB (\$dummy [44]), .D (nx793), .CLK (nx1502
         ), .R (nx1476)) ;
    mux21_ni ix794 (.Y (nx793), .A0 (q_0__8), .A1 (d[8]), .S0 (nx1450)) ;
    dffr gen_regs_4_regi_reg_q_9 (.Q (q_4__9), .QB (\$dummy [45]), .D (nx883), .CLK (
         nx1506), .R (nx1480)) ;
    mux21_ni ix884 (.Y (nx883), .A0 (q_4__9), .A1 (q_3__9), .S0 (nx1454)) ;
    dffr gen_regs_3_regi_reg_q_9 (.Q (q_3__9), .QB (\$dummy [46]), .D (nx873), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix874 (.Y (nx873), .A0 (q_3__9), .A1 (q_2__9), .S0 (nx1452)) ;
    dffr gen_regs_2_regi_reg_q_9 (.Q (q_2__9), .QB (\$dummy [47]), .D (nx863), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix864 (.Y (nx863), .A0 (q_2__9), .A1 (q_1__9), .S0 (nx1452)) ;
    dffr gen_regs_1_regi_reg_q_9 (.Q (q_1__9), .QB (\$dummy [48]), .D (nx853), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix854 (.Y (nx853), .A0 (q_1__9), .A1 (q_0__9), .S0 (nx1452)) ;
    dffr reg0_reg_q_9 (.Q (q_0__9), .QB (\$dummy [49]), .D (nx843), .CLK (nx1504
         ), .R (nx1478)) ;
    mux21_ni ix844 (.Y (nx843), .A0 (q_0__9), .A1 (d[9]), .S0 (nx1452)) ;
    dffr gen_regs_4_regi_reg_q_10 (.Q (q_4__10), .QB (\$dummy [50]), .D (nx933)
         , .CLK (nx1506), .R (nx1480)) ;
    mux21_ni ix934 (.Y (nx933), .A0 (q_4__10), .A1 (q_3__10), .S0 (nx1454)) ;
    dffr gen_regs_3_regi_reg_q_10 (.Q (q_3__10), .QB (\$dummy [51]), .D (nx923)
         , .CLK (nx1506), .R (nx1480)) ;
    mux21_ni ix924 (.Y (nx923), .A0 (q_3__10), .A1 (q_2__10), .S0 (nx1454)) ;
    dffr gen_regs_2_regi_reg_q_10 (.Q (q_2__10), .QB (\$dummy [52]), .D (nx913)
         , .CLK (nx1506), .R (nx1480)) ;
    mux21_ni ix914 (.Y (nx913), .A0 (q_2__10), .A1 (q_1__10), .S0 (nx1454)) ;
    dffr gen_regs_1_regi_reg_q_10 (.Q (q_1__10), .QB (\$dummy [53]), .D (nx903)
         , .CLK (nx1506), .R (nx1480)) ;
    mux21_ni ix904 (.Y (nx903), .A0 (q_1__10), .A1 (q_0__10), .S0 (nx1454)) ;
    dffr reg0_reg_q_10 (.Q (q_0__10), .QB (\$dummy [54]), .D (nx893), .CLK (
         nx1506), .R (nx1480)) ;
    mux21_ni ix894 (.Y (nx893), .A0 (q_0__10), .A1 (d[10]), .S0 (nx1454)) ;
    dffr gen_regs_4_regi_reg_q_11 (.Q (q_4__11), .QB (\$dummy [55]), .D (nx983)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix984 (.Y (nx983), .A0 (q_4__11), .A1 (q_3__11), .S0 (nx1456)) ;
    dffr gen_regs_3_regi_reg_q_11 (.Q (q_3__11), .QB (\$dummy [56]), .D (nx973)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix974 (.Y (nx973), .A0 (q_3__11), .A1 (q_2__11), .S0 (nx1456)) ;
    dffr gen_regs_2_regi_reg_q_11 (.Q (q_2__11), .QB (\$dummy [57]), .D (nx963)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix964 (.Y (nx963), .A0 (q_2__11), .A1 (q_1__11), .S0 (nx1456)) ;
    dffr gen_regs_1_regi_reg_q_11 (.Q (q_1__11), .QB (\$dummy [58]), .D (nx953)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix954 (.Y (nx953), .A0 (q_1__11), .A1 (q_0__11), .S0 (nx1456)) ;
    dffr reg0_reg_q_11 (.Q (q_0__11), .QB (\$dummy [59]), .D (nx943), .CLK (
         nx1506), .R (nx1480)) ;
    mux21_ni ix944 (.Y (nx943), .A0 (q_0__11), .A1 (d[11]), .S0 (nx1454)) ;
    dffr gen_regs_4_regi_reg_q_12 (.Q (q_4__12), .QB (\$dummy [60]), .D (nx1033)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1034 (.Y (nx1033), .A0 (q_4__12), .A1 (q_3__12), .S0 (nx1458)) ;
    dffr gen_regs_3_regi_reg_q_12 (.Q (q_3__12), .QB (\$dummy [61]), .D (nx1023)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1024 (.Y (nx1023), .A0 (q_3__12), .A1 (q_2__12), .S0 (nx1458)) ;
    dffr gen_regs_2_regi_reg_q_12 (.Q (q_2__12), .QB (\$dummy [62]), .D (nx1013)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix1014 (.Y (nx1013), .A0 (q_2__12), .A1 (q_1__12), .S0 (nx1456)) ;
    dffr gen_regs_1_regi_reg_q_12 (.Q (q_1__12), .QB (\$dummy [63]), .D (nx1003)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix1004 (.Y (nx1003), .A0 (q_1__12), .A1 (q_0__12), .S0 (nx1456)) ;
    dffr reg0_reg_q_12 (.Q (q_0__12), .QB (\$dummy [64]), .D (nx993), .CLK (
         nx1508), .R (nx1482)) ;
    mux21_ni ix994 (.Y (nx993), .A0 (q_0__12), .A1 (d[12]), .S0 (nx1456)) ;
    dffr gen_regs_4_regi_reg_q_13 (.Q (q_4__13), .QB (\$dummy [65]), .D (nx1083)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1084 (.Y (nx1083), .A0 (q_4__13), .A1 (q_3__13), .S0 (nx1458)) ;
    dffr gen_regs_3_regi_reg_q_13 (.Q (q_3__13), .QB (\$dummy [66]), .D (nx1073)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1074 (.Y (nx1073), .A0 (q_3__13), .A1 (q_2__13), .S0 (nx1458)) ;
    dffr gen_regs_2_regi_reg_q_13 (.Q (q_2__13), .QB (\$dummy [67]), .D (nx1063)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1064 (.Y (nx1063), .A0 (q_2__13), .A1 (q_1__13), .S0 (nx1458)) ;
    dffr gen_regs_1_regi_reg_q_13 (.Q (q_1__13), .QB (\$dummy [68]), .D (nx1053)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1054 (.Y (nx1053), .A0 (q_1__13), .A1 (q_0__13), .S0 (nx1458)) ;
    dffr reg0_reg_q_13 (.Q (q_0__13), .QB (\$dummy [69]), .D (nx1043), .CLK (
         nx1510), .R (nx1484)) ;
    mux21_ni ix1044 (.Y (nx1043), .A0 (q_0__13), .A1 (d[13]), .S0 (nx1458)) ;
    dffr gen_regs_4_regi_reg_q_14 (.Q (q_4__14), .QB (\$dummy [70]), .D (nx1133)
         , .CLK (nx1512), .R (nx1486)) ;
    mux21_ni ix1134 (.Y (nx1133), .A0 (q_4__14), .A1 (q_3__14), .S0 (nx1460)) ;
    dffr gen_regs_3_regi_reg_q_14 (.Q (q_3__14), .QB (\$dummy [71]), .D (nx1123)
         , .CLK (nx1512), .R (nx1486)) ;
    mux21_ni ix1124 (.Y (nx1123), .A0 (q_3__14), .A1 (q_2__14), .S0 (nx1460)) ;
    dffr gen_regs_2_regi_reg_q_14 (.Q (q_2__14), .QB (\$dummy [72]), .D (nx1113)
         , .CLK (nx1512), .R (nx1486)) ;
    mux21_ni ix1114 (.Y (nx1113), .A0 (q_2__14), .A1 (q_1__14), .S0 (nx1460)) ;
    dffr gen_regs_1_regi_reg_q_14 (.Q (q_1__14), .QB (\$dummy [73]), .D (nx1103)
         , .CLK (nx1512), .R (nx1486)) ;
    mux21_ni ix1104 (.Y (nx1103), .A0 (q_1__14), .A1 (q_0__14), .S0 (nx1460)) ;
    dffr reg0_reg_q_14 (.Q (q_0__14), .QB (\$dummy [74]), .D (nx1093), .CLK (
         nx1512), .R (nx1486)) ;
    mux21_ni ix1094 (.Y (nx1093), .A0 (q_0__14), .A1 (d[14]), .S0 (nx1460)) ;
    dffr gen_regs_4_regi_reg_q_15 (.Q (q_4__15), .QB (\$dummy [75]), .D (nx1183)
         , .CLK (nx1514), .R (nx1488)) ;
    mux21_ni ix1184 (.Y (nx1183), .A0 (q_4__15), .A1 (q_3__15), .S0 (nx1462)) ;
    dffr gen_regs_3_regi_reg_q_15 (.Q (q_3__15), .QB (\$dummy [76]), .D (nx1173)
         , .CLK (nx1514), .R (nx1488)) ;
    mux21_ni ix1174 (.Y (nx1173), .A0 (q_3__15), .A1 (q_2__15), .S0 (nx1462)) ;
    dffr gen_regs_2_regi_reg_q_15 (.Q (q_2__15), .QB (\$dummy [77]), .D (nx1163)
         , .CLK (nx1514), .R (nx1488)) ;
    mux21_ni ix1164 (.Y (nx1163), .A0 (q_2__15), .A1 (q_1__15), .S0 (nx1462)) ;
    dffr gen_regs_1_regi_reg_q_15 (.Q (q_1__15), .QB (\$dummy [78]), .D (nx1153)
         , .CLK (nx1512), .R (nx1486)) ;
    mux21_ni ix1154 (.Y (nx1153), .A0 (q_1__15), .A1 (q_0__15), .S0 (nx1460)) ;
    dffr reg0_reg_q_15 (.Q (q_0__15), .QB (\$dummy [79]), .D (nx1143), .CLK (
         nx1512), .R (nx1486)) ;
    mux21_ni ix1144 (.Y (nx1143), .A0 (q_0__15), .A1 (d[15]), .S0 (nx1460)) ;
    inv02 ix1439 (.Y (nx1440), .A (nx1516)) ;
    inv02 ix1441 (.Y (nx1442), .A (nx1516)) ;
    inv02 ix1443 (.Y (nx1444), .A (nx1516)) ;
    inv02 ix1445 (.Y (nx1446), .A (nx1516)) ;
    inv02 ix1447 (.Y (nx1448), .A (nx1516)) ;
    inv02 ix1449 (.Y (nx1450), .A (nx1516)) ;
    inv02 ix1451 (.Y (nx1452), .A (nx1516)) ;
    inv02 ix1453 (.Y (nx1454), .A (nx1518)) ;
    inv02 ix1455 (.Y (nx1456), .A (nx1518)) ;
    inv02 ix1457 (.Y (nx1458), .A (nx1518)) ;
    inv02 ix1459 (.Y (nx1460), .A (nx1518)) ;
    inv02 ix1461 (.Y (nx1462), .A (nx1518)) ;
    inv02 ix1465 (.Y (nx1466), .A (nx1520)) ;
    inv02 ix1467 (.Y (nx1468), .A (nx1520)) ;
    inv02 ix1469 (.Y (nx1470), .A (nx1520)) ;
    inv02 ix1471 (.Y (nx1472), .A (nx1520)) ;
    inv02 ix1473 (.Y (nx1474), .A (nx1520)) ;
    inv02 ix1475 (.Y (nx1476), .A (nx1520)) ;
    inv02 ix1477 (.Y (nx1478), .A (nx1520)) ;
    inv02 ix1479 (.Y (nx1480), .A (nx1522)) ;
    inv02 ix1481 (.Y (nx1482), .A (nx1522)) ;
    inv02 ix1483 (.Y (nx1484), .A (nx1522)) ;
    inv02 ix1485 (.Y (nx1486), .A (nx1522)) ;
    inv02 ix1487 (.Y (nx1488), .A (nx1522)) ;
    inv02 ix1491 (.Y (nx1492), .A (nx1524)) ;
    inv02 ix1493 (.Y (nx1494), .A (nx1524)) ;
    inv02 ix1495 (.Y (nx1496), .A (nx1524)) ;
    inv02 ix1497 (.Y (nx1498), .A (nx1524)) ;
    inv02 ix1499 (.Y (nx1500), .A (nx1524)) ;
    inv02 ix1501 (.Y (nx1502), .A (nx1524)) ;
    inv02 ix1503 (.Y (nx1504), .A (nx1524)) ;
    inv02 ix1505 (.Y (nx1506), .A (nx1526)) ;
    inv02 ix1507 (.Y (nx1508), .A (nx1526)) ;
    inv02 ix1509 (.Y (nx1510), .A (nx1526)) ;
    inv02 ix1511 (.Y (nx1512), .A (nx1526)) ;
    inv02 ix1513 (.Y (nx1514), .A (nx1526)) ;
    inv02 ix1515 (.Y (nx1516), .A (load)) ;
    inv02 ix1517 (.Y (nx1518), .A (load)) ;
    inv02 ix1519 (.Y (nx1520), .A (reset)) ;
    inv02 ix1521 (.Y (nx1522), .A (reset)) ;
    inv02 ix1523 (.Y (nx1524), .A (clk)) ;
    inv02 ix1525 (.Y (nx1526), .A (clk)) ;
endmodule

