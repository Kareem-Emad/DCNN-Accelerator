* SPICE NETLIST
***************************************

.SUBCKT mux21_ni S0 A1 A0 Y GND VDD
** N=24 EP=6 IP=0 FDC=12
M0 GND S0 7 GND N L=4e-07 W=1e-06 AD=2.4e-12 AS=1.1e-12 $X=11500 $Y=31000 $D=1
M1 21 S0 GND GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.4e-12 $X=20000 $Y=26000 $D=1
M2 8 A1 21 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=25000 $Y=26000 $D=1
M3 22 A0 8 GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.4e-12 $X=33000 $Y=26000 $D=1
M4 GND 7 22 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=38000 $Y=26000 $D=1
M5 Y 8 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=2.4e-12 $X=46500 $Y=31000 $D=1
M6 VDD S0 7 VDD P L=4e-07 W=1.8e-06 AD=4.32e-12 AS=1.58e-12 $X=11500 $Y=71000 $D=0
M7 23 S0 VDD VDD P L=4e-07 W=3.6e-06 AD=2.16e-12 AS=4.32e-12 $X=20000 $Y=71000 $D=0
M8 8 A0 23 VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=2.16e-12 $X=25000 $Y=71000 $D=0
M9 24 A1 8 VDD P L=4e-07 W=3.6e-06 AD=2.16e-12 AS=4.32e-12 $X=33000 $Y=71000 $D=0
M10 VDD 7 24 VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=2.16e-12 $X=38000 $Y=71000 $D=0
M11 Y 8 VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=4.32e-12 $X=46500 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT nwell_contact
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT inv01 A Y GND VDD
** N=6 EP=4 IP=1 FDC=2
M0 Y A GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.1e-12 $X=11500 $Y=26000 $D=1
M1 Y A VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=1.58e-12 $X=11500 $Y=80000 $D=0
.ENDS
***************************************
.SUBCKT inv02 A Y GND VDD
** N=6 EP=4 IP=1 FDC=2
M0 Y A GND GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 Y A VDD VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=3.66e-12 $X=11500 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT nand02 A1 A0 Y GND VDD
** N=10 EP=5 IP=2 FDC=4
M0 10 A1 GND GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 Y A0 10 GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=1.2e-12 $X=16500 $Y=26000 $D=1
M2 Y A1 VDD VDD P L=4e-07 W=2.4e-06 AD=2.88e-12 AS=2.44e-12 $X=11500 $Y=77000 $D=0
M3 VDD A0 Y VDD P L=4e-07 W=2.4e-06 AD=2.44e-12 AS=2.88e-12 $X=19500 $Y=77000 $D=0
.ENDS
***************************************
.SUBCKT dffr D CLK R Q GND VDD
** N=59 EP=6 IP=9 FDC=34
M0 52 D GND GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.3e-12 $X=11500 $Y=26000 $D=1
M1 8 12 52 GND N L=4e-07 W=3e-06 AD=3.5e-12 AS=1.8e-12 $X=16500 $Y=26000 $D=1
M2 53 11 8 GND N L=4e-07 W=1e-06 AD=6e-13 AS=3.5e-12 $X=25000 $Y=31000 $D=1
M3 GND 9 53 GND N L=4e-07 W=1e-06 AD=2.4e-12 AS=6e-13 $X=30000 $Y=31000 $D=1
M4 9 8 GND GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=38500 $Y=26000 $D=1
M5 GND R 9 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=46500 $Y=26000 $D=1
M6 10 9 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=2.4e-12 $X=55000 $Y=31000 $D=1
M7 GND 12 11 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=76000 $Y=31000 $D=1
M8 12 CLK GND GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=84000 $Y=31000 $D=1
M9 54 10 GND GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.3e-12 $X=100000 $Y=26000 $D=1
M10 13 11 54 GND N L=4e-07 W=3e-06 AD=3.5e-12 AS=1.8e-12 $X=105000 $Y=26000 $D=1
M11 14 12 13 GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=3.5e-12 $X=113500 $Y=26000 $D=1
M12 14 R GND GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.1e-12 $X=130500 $Y=26000 $D=1
M13 GND 15 14 GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.2e-12 $X=138500 $Y=26000 $D=1
M14 15 13 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.2e-12 $X=146500 $Y=26000 $D=1
M15 GND 13 QB GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=162500 $Y=31000 $D=1
M16 Q QB GND GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=170500 $Y=31000 $D=1
M17 55 11 VDD VDD P L=4e-07 W=5.4e-06 AD=3.24e-12 AS=5.74e-12 $X=11500 $Y=62000 $D=0
M18 8 D 55 VDD P L=4e-07 W=5.4e-06 AD=6.14e-12 AS=3.24e-12 $X=16500 $Y=62000 $D=0
M19 56 12 8 VDD P L=4e-07 W=1e-06 AD=6e-13 AS=6.14e-12 $X=25000 $Y=62000 $D=0
M20 VDD 9 56 VDD P L=4e-07 W=1e-06 AD=1.1e-12 AS=6e-13 $X=30000 $Y=62000 $D=0
M21 57 8 9 VDD P L=4e-07 W=2.4e-06 AD=1.44e-12 AS=2.44e-12 $X=46000 $Y=62000 $D=0
M22 VDD R 57 VDD P L=4e-07 W=2.4e-06 AD=3e-12 AS=1.44e-12 $X=51000 $Y=62000 $D=0
M23 10 9 VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=3e-12 $X=59500 $Y=62000 $D=0
M24 VDD 12 11 VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=3.66e-12 $X=76000 $Y=62000 $D=0
M25 12 CLK VDD VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=4.32e-12 $X=84000 $Y=62000 $D=0
M26 58 10 VDD VDD P L=4e-07 W=5.4e-06 AD=3.24e-12 AS=5.74e-12 $X=100000 $Y=53000 $D=0
M27 13 12 58 VDD P L=4e-07 W=5.4e-06 AD=6.14e-12 AS=3.24e-12 $X=105000 $Y=53000 $D=0
M28 14 11 13 VDD P L=4e-07 W=1e-06 AD=1.2e-12 AS=6.14e-12 $X=113500 $Y=68000 $D=0
M29 59 R 14 VDD P L=4e-07 W=1e-06 AD=6e-13 AS=1.2e-12 $X=121500 $Y=68000 $D=0
M30 VDD 15 59 VDD P L=4e-07 W=1e-06 AD=1.2e-12 AS=6e-13 $X=126500 $Y=68000 $D=0
M31 15 13 VDD VDD P L=4e-07 W=1e-06 AD=1.1e-12 AS=1.2e-12 $X=134500 $Y=68000 $D=0
M32 VDD 13 QB VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=3.66e-12 $X=162500 $Y=62000 $D=0
M33 Q QB VDD VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=4.32e-12 $X=170500 $Y=62000 $D=0
.ENDS
***************************************
.SUBCKT DCNNChip
** N=202 EP=0 IP=453 FDC=844
X0 10 33 27 138 136 137 mux21_ni $T=212000 72000 1 180 $X=152000 $Y=72000
X1 10 32 38 139 136 137 mux21_ni $T=152000 232000 0 0 $X=152000 $Y=232000
X2 39 34 28 140 136 137 mux21_ni $T=152000 392000 0 0 $X=152000 $Y=392000
X3 2 35 29 141 136 137 mux21_ni $T=152000 552000 0 0 $X=152000 $Y=552000
X4 1 36 30 142 136 137 mux21_ni $T=152000 712000 0 0 $X=152000 $Y=712000
X5 3 37 31 143 136 137 mux21_ni $T=152000 872000 0 0 $X=152000 $Y=872000
X6 39 27 33 144 136 137 mux21_ni $T=216000 72000 0 0 $X=216000 $Y=72000
X7 39 38 32 145 136 137 mux21_ni $T=276000 232000 1 180 $X=216000 $Y=232000
X8 10 28 34 146 136 137 mux21_ni $T=216000 392000 0 0 $X=216000 $Y=392000
X9 3 29 35 147 136 137 mux21_ni $T=216000 552000 0 0 $X=216000 $Y=552000
X10 3 30 36 148 136 137 mux21_ni $T=216000 712000 0 0 $X=216000 $Y=712000
X11 1 31 37 149 136 137 mux21_ni $T=216000 872000 0 0 $X=216000 $Y=872000
X12 39 46 40 150 136 137 mux21_ni $T=280000 72000 0 0 $X=280000 $Y=72000
X13 12 47 41 151 136 137 mux21_ni $T=280000 232000 0 0 $X=280000 $Y=232000
X14 12 48 42 152 136 137 mux21_ni $T=280000 392000 0 0 $X=280000 $Y=392000
X15 1 49 43 153 136 137 mux21_ni $T=280000 552000 0 0 $X=280000 $Y=552000
X16 2 50 44 154 136 137 mux21_ni $T=280000 712000 0 0 $X=280000 $Y=712000
X17 1 51 45 155 136 137 mux21_ni $T=280000 872000 0 0 $X=280000 $Y=872000
X18 5 40 46 156 136 137 mux21_ni $T=344000 72000 0 0 $X=344000 $Y=72000
X19 52 41 47 157 136 137 mux21_ni $T=344000 232000 0 0 $X=344000 $Y=232000
X20 10 42 48 158 136 137 mux21_ni $T=344000 392000 0 0 $X=344000 $Y=392000
X21 4 43 49 159 136 137 mux21_ni $T=344000 552000 0 0 $X=344000 $Y=552000
X22 3 44 50 160 136 137 mux21_ni $T=344000 712000 0 0 $X=344000 $Y=712000
X23 4 45 51 161 136 137 mux21_ni $T=344000 872000 0 0 $X=344000 $Y=872000
X24 52 58 53 162 136 137 mux21_ni $T=408000 72000 0 0 $X=408000 $Y=72000
X25 10 59 54 163 136 137 mux21_ni $T=408000 232000 0 0 $X=408000 $Y=232000
X26 4 57 55 164 136 137 mux21_ni $T=408000 552000 0 0 $X=408000 $Y=552000
X27 4 62 61 165 136 137 mux21_ni $T=408000 712000 0 0 $X=408000 $Y=712000
X28 12 60 56 166 136 137 mux21_ni $T=408000 872000 0 0 $X=408000 $Y=872000
X29 5 53 58 167 136 137 mux21_ni $T=472000 72000 0 0 $X=472000 $Y=72000
X30 12 54 59 168 136 137 mux21_ni $T=472000 392000 0 0 $X=472000 $Y=392000
X31 1 55 57 169 136 137 mux21_ni $T=472000 712000 0 0 $X=472000 $Y=712000
X32 52 56 60 170 136 137 mux21_ni $T=472000 872000 0 0 $X=472000 $Y=872000
X33 4 68 63 171 136 137 mux21_ni $T=536000 72000 0 0 $X=536000 $Y=72000
X34 52 69 64 172 136 137 mux21_ni $T=536000 232000 0 0 $X=536000 $Y=232000
X35 52 70 65 173 136 137 mux21_ni $T=536000 392000 0 0 $X=536000 $Y=392000
X36 83 71 66 174 136 137 mux21_ni $T=536000 552000 0 0 $X=536000 $Y=552000
X37 83 61 62 175 136 137 mux21_ni $T=536000 712000 0 0 $X=536000 $Y=712000
X38 52 72 67 176 136 137 mux21_ni $T=536000 872000 0 0 $X=536000 $Y=872000
X39 1 63 68 177 136 137 mux21_ni $T=600000 72000 0 0 $X=600000 $Y=72000
X40 12 64 69 178 136 137 mux21_ni $T=600000 232000 0 0 $X=600000 $Y=232000
X41 5 65 70 179 136 137 mux21_ni $T=600000 392000 0 0 $X=600000 $Y=392000
X42 4 66 71 180 136 137 mux21_ni $T=600000 552000 0 0 $X=600000 $Y=552000
X43 52 79 76 181 136 137 mux21_ni $T=600000 712000 0 0 $X=600000 $Y=712000
X44 5 67 72 182 136 137 mux21_ni $T=600000 872000 0 0 $X=600000 $Y=872000
X45 1 77 74 183 136 137 mux21_ni $T=664000 72000 0 0 $X=664000 $Y=72000
X46 3 9 13 184 136 137 mux21_ni $T=664000 232000 0 0 $X=664000 $Y=232000
X47 3 78 75 185 136 137 mux21_ni $T=664000 392000 0 0 $X=664000 $Y=392000
X48 2 73 6 186 136 137 mux21_ni $T=664000 552000 0 0 $X=664000 $Y=552000
X49 3 6 73 187 136 137 mux21_ni $T=664000 712000 0 0 $X=664000 $Y=712000
X50 5 81 7 188 136 137 mux21_ni $T=664000 872000 0 0 $X=664000 $Y=872000
X51 4 74 77 189 136 137 mux21_ni $T=728000 72000 0 0 $X=728000 $Y=72000
X52 2 75 78 190 136 137 mux21_ni $T=728000 392000 0 0 $X=728000 $Y=392000
X53 12 76 79 191 136 137 mux21_ni $T=728000 712000 0 0 $X=728000 $Y=712000
X54 2 87 85 192 136 137 mux21_ni $T=760000 232000 0 0 $X=760000 $Y=232000
X55 10 92 90 193 136 137 mux21_ni $T=792000 72000 0 0 $X=792000 $Y=72000
X56 83 95 94 194 136 137 mux21_ni $T=792000 392000 0 0 $X=792000 $Y=392000
X57 39 86 84 195 136 137 mux21_ni $T=824000 232000 0 0 $X=824000 $Y=232000
X58 10 84 86 196 136 137 mux21_ni $T=856000 72000 0 0 $X=856000 $Y=72000
X59 83 85 87 197 136 137 mux21_ni $T=856000 392000 0 0 $X=856000 $Y=392000
X60 2 13 9 198 136 137 mux21_ni $T=888000 232000 0 0 $X=888000 $Y=232000
X61 39 90 92 199 136 137 mux21_ni $T=920000 72000 0 0 $X=920000 $Y=72000
X62 39 7 81 200 136 137 mux21_ni $T=920000 392000 0 0 $X=920000 $Y=392000
X63 201 91 93 96 136 137 mux21_ni $T=920000 712000 0 0 $X=920000 $Y=712000
X64 2 94 95 202 136 137 mux21_ni $T=952000 232000 0 0 $X=952000 $Y=232000
X65 91 82 136 137 inv01 $T=792000 872000 0 0 $X=792000 $Y=872000
X66 88 80 136 137 inv01 $T=921000 872000 1 180 $X=896000 $Y=872000
X67 8 39 136 137 inv02 $T=728000 232000 0 0 $X=728000 $Y=232000
X68 8 52 136 137 inv02 $T=753000 552000 1 180 $X=728000 $Y=552000
X69 80 3 136 137 inv02 $T=753000 872000 1 180 $X=728000 $Y=872000
X70 8 10 136 137 inv02 $T=760000 552000 0 0 $X=760000 $Y=552000
X71 80 1 136 137 inv02 $T=785000 872000 1 180 $X=760000 $Y=872000
X72 8 12 136 137 inv02 $T=792000 552000 0 0 $X=792000 $Y=552000
X73 80 2 136 137 inv02 $T=792000 712000 0 0 $X=792000 $Y=712000
X74 8 5 136 137 inv02 $T=824000 712000 0 0 $X=824000 $Y=712000
X75 80 4 136 137 inv02 $T=849000 872000 1 180 $X=824000 $Y=872000
X76 80 83 136 137 inv02 $T=856000 712000 0 0 $X=856000 $Y=712000
X77 12 93 136 137 inv02 $T=888000 712000 0 0 $X=888000 $Y=712000
X78 82 5 88 136 137 nand02 $T=856000 872000 0 0 $X=856000 $Y=872000
X79 96 89 11 8 136 137 dffr $T=1008000 552000 1 180 $X=824000 $Y=552000
.ENDS
***************************************
