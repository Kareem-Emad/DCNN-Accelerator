library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;

entity ControlUnitTB is
end ControlUnitTB;

architecture TB of ControlUnitTB is
begin
end TB;