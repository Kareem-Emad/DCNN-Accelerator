
-- 
-- Definition of  Controller
-- 
--      Fri May 10 20:13:02 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Queue_5 is
   port (
      d : IN std_logic_vector (15 DOWNTO 0) ;
      q_0_15 : OUT std_logic ;
      q_0_14 : OUT std_logic ;
      q_0_13 : OUT std_logic ;
      q_0_12 : OUT std_logic ;
      q_0_11 : OUT std_logic ;
      q_0_10 : OUT std_logic ;
      q_0_9 : OUT std_logic ;
      q_0_8 : OUT std_logic ;
      q_0_7 : OUT std_logic ;
      q_0_6 : OUT std_logic ;
      q_0_5 : OUT std_logic ;
      q_0_4 : OUT std_logic ;
      q_0_3 : OUT std_logic ;
      q_0_2 : OUT std_logic ;
      q_0_1 : OUT std_logic ;
      q_0_0 : OUT std_logic ;
      q_1_15 : OUT std_logic ;
      q_1_14 : OUT std_logic ;
      q_1_13 : OUT std_logic ;
      q_1_12 : OUT std_logic ;
      q_1_11 : OUT std_logic ;
      q_1_10 : OUT std_logic ;
      q_1_9 : OUT std_logic ;
      q_1_8 : OUT std_logic ;
      q_1_7 : OUT std_logic ;
      q_1_6 : OUT std_logic ;
      q_1_5 : OUT std_logic ;
      q_1_4 : OUT std_logic ;
      q_1_3 : OUT std_logic ;
      q_1_2 : OUT std_logic ;
      q_1_1 : OUT std_logic ;
      q_1_0 : OUT std_logic ;
      q_2_15 : OUT std_logic ;
      q_2_14 : OUT std_logic ;
      q_2_13 : OUT std_logic ;
      q_2_12 : OUT std_logic ;
      q_2_11 : OUT std_logic ;
      q_2_10 : OUT std_logic ;
      q_2_9 : OUT std_logic ;
      q_2_8 : OUT std_logic ;
      q_2_7 : OUT std_logic ;
      q_2_6 : OUT std_logic ;
      q_2_5 : OUT std_logic ;
      q_2_4 : OUT std_logic ;
      q_2_3 : OUT std_logic ;
      q_2_2 : OUT std_logic ;
      q_2_1 : OUT std_logic ;
      q_2_0 : OUT std_logic ;
      q_3_15 : OUT std_logic ;
      q_3_14 : OUT std_logic ;
      q_3_13 : OUT std_logic ;
      q_3_12 : OUT std_logic ;
      q_3_11 : OUT std_logic ;
      q_3_10 : OUT std_logic ;
      q_3_9 : OUT std_logic ;
      q_3_8 : OUT std_logic ;
      q_3_7 : OUT std_logic ;
      q_3_6 : OUT std_logic ;
      q_3_5 : OUT std_logic ;
      q_3_4 : OUT std_logic ;
      q_3_3 : OUT std_logic ;
      q_3_2 : OUT std_logic ;
      q_3_1 : OUT std_logic ;
      q_3_0 : OUT std_logic ;
      q_4_15 : OUT std_logic ;
      q_4_14 : OUT std_logic ;
      q_4_13 : OUT std_logic ;
      q_4_12 : OUT std_logic ;
      q_4_11 : OUT std_logic ;
      q_4_10 : OUT std_logic ;
      q_4_9 : OUT std_logic ;
      q_4_8 : OUT std_logic ;
      q_4_7 : OUT std_logic ;
      q_4_6 : OUT std_logic ;
      q_4_5 : OUT std_logic ;
      q_4_4 : OUT std_logic ;
      q_4_3 : OUT std_logic ;
      q_4_2 : OUT std_logic ;
      q_4_1 : OUT std_logic ;
      q_4_0 : OUT std_logic ;
      clk : IN std_logic ;
      load : IN std_logic ;
      reset : IN std_logic) ;
end Queue_5 ;

architecture Dataflow of Queue_5 is
   signal q_0_15_EXMPLR, q_0_14_EXMPLR, q_0_13_EXMPLR, q_0_12_EXMPLR, 
      q_0_11_EXMPLR, q_0_10_EXMPLR, q_0_9_EXMPLR, q_0_8_EXMPLR, q_0_7_EXMPLR, 
      q_0_6_EXMPLR, q_0_5_EXMPLR, q_0_4_EXMPLR, q_0_3_EXMPLR, q_0_2_EXMPLR, 
      q_0_1_EXMPLR, q_0_0_EXMPLR, q_1_15_EXMPLR, q_1_14_EXMPLR, 
      q_1_13_EXMPLR, q_1_12_EXMPLR, q_1_11_EXMPLR, q_1_10_EXMPLR, 
      q_1_9_EXMPLR, q_1_8_EXMPLR, q_1_7_EXMPLR, q_1_6_EXMPLR, q_1_5_EXMPLR, 
      q_1_4_EXMPLR, q_1_3_EXMPLR, q_1_2_EXMPLR, q_1_1_EXMPLR, q_1_0_EXMPLR, 
      q_2_15_EXMPLR, q_2_14_EXMPLR, q_2_13_EXMPLR, q_2_12_EXMPLR, 
      q_2_11_EXMPLR, q_2_10_EXMPLR, q_2_9_EXMPLR, q_2_8_EXMPLR, q_2_7_EXMPLR, 
      q_2_6_EXMPLR, q_2_5_EXMPLR, q_2_4_EXMPLR, q_2_3_EXMPLR, q_2_2_EXMPLR, 
      q_2_1_EXMPLR, q_2_0_EXMPLR, q_3_15_EXMPLR, q_3_14_EXMPLR, 
      q_3_13_EXMPLR, q_3_12_EXMPLR, q_3_11_EXMPLR, q_3_10_EXMPLR, 
      q_3_9_EXMPLR, q_3_8_EXMPLR, q_3_7_EXMPLR, q_3_6_EXMPLR, q_3_5_EXMPLR, 
      q_3_4_EXMPLR, q_3_3_EXMPLR, q_3_2_EXMPLR, q_3_1_EXMPLR, q_3_0_EXMPLR, 
      q_4_15_EXMPLR, q_4_14_EXMPLR, q_4_13_EXMPLR, q_4_12_EXMPLR, 
      q_4_11_EXMPLR, q_4_10_EXMPLR, q_4_9_EXMPLR, q_4_8_EXMPLR, q_4_7_EXMPLR, 
      q_4_6_EXMPLR, q_4_5_EXMPLR, q_4_4_EXMPLR, q_4_3_EXMPLR, q_4_2_EXMPLR, 
      q_4_1_EXMPLR, q_4_0_EXMPLR, nx393, nx403, nx413, nx423, nx433, nx443, 
      nx453, nx463, nx473, nx483, nx493, nx503, nx513, nx523, nx533, nx543, 
      nx553, nx563, nx573, nx583, nx593, nx603, nx613, nx623, nx633, nx643, 
      nx653, nx663, nx673, nx683, nx693, nx703, nx713, nx723, nx733, nx743, 
      nx753, nx763, nx773, nx783, nx793, nx803, nx813, nx823, nx833, nx843, 
      nx853, nx863, nx873, nx883, nx893, nx903, nx913, nx923, nx933, nx943, 
      nx953, nx963, nx973, nx983, nx993, nx1003, nx1013, nx1023, nx1033, 
      nx1043, nx1053, nx1063, nx1073, nx1083, nx1093, nx1103, nx1113, nx1123, 
      nx1133, nx1143, nx1153, nx1163, nx1173, nx1183, nx1440, nx1442, nx1444, 
      nx1446, nx1448, nx1450, nx1452, nx1454, nx1456, nx1458, nx1460, nx1462, 
      nx1466, nx1468, nx1470, nx1472, nx1474, nx1476, nx1478, nx1480, nx1482, 
      nx1484, nx1486, nx1488, nx1492, nx1494, nx1496, nx1498, nx1500, nx1502, 
      nx1504, nx1506, nx1508, nx1510, nx1512, nx1514, nx1516, nx1518, nx1520, 
      nx1522, nx1524, nx1526: std_logic ;

begin
   q_0_15 <= q_0_15_EXMPLR ;
   q_0_14 <= q_0_14_EXMPLR ;
   q_0_13 <= q_0_13_EXMPLR ;
   q_0_12 <= q_0_12_EXMPLR ;
   q_0_11 <= q_0_11_EXMPLR ;
   q_0_10 <= q_0_10_EXMPLR ;
   q_0_9 <= q_0_9_EXMPLR ;
   q_0_8 <= q_0_8_EXMPLR ;
   q_0_7 <= q_0_7_EXMPLR ;
   q_0_6 <= q_0_6_EXMPLR ;
   q_0_5 <= q_0_5_EXMPLR ;
   q_0_4 <= q_0_4_EXMPLR ;
   q_0_3 <= q_0_3_EXMPLR ;
   q_0_2 <= q_0_2_EXMPLR ;
   q_0_1 <= q_0_1_EXMPLR ;
   q_0_0 <= q_0_0_EXMPLR ;
   q_1_15 <= q_1_15_EXMPLR ;
   q_1_14 <= q_1_14_EXMPLR ;
   q_1_13 <= q_1_13_EXMPLR ;
   q_1_12 <= q_1_12_EXMPLR ;
   q_1_11 <= q_1_11_EXMPLR ;
   q_1_10 <= q_1_10_EXMPLR ;
   q_1_9 <= q_1_9_EXMPLR ;
   q_1_8 <= q_1_8_EXMPLR ;
   q_1_7 <= q_1_7_EXMPLR ;
   q_1_6 <= q_1_6_EXMPLR ;
   q_1_5 <= q_1_5_EXMPLR ;
   q_1_4 <= q_1_4_EXMPLR ;
   q_1_3 <= q_1_3_EXMPLR ;
   q_1_2 <= q_1_2_EXMPLR ;
   q_1_1 <= q_1_1_EXMPLR ;
   q_1_0 <= q_1_0_EXMPLR ;
   q_2_15 <= q_2_15_EXMPLR ;
   q_2_14 <= q_2_14_EXMPLR ;
   q_2_13 <= q_2_13_EXMPLR ;
   q_2_12 <= q_2_12_EXMPLR ;
   q_2_11 <= q_2_11_EXMPLR ;
   q_2_10 <= q_2_10_EXMPLR ;
   q_2_9 <= q_2_9_EXMPLR ;
   q_2_8 <= q_2_8_EXMPLR ;
   q_2_7 <= q_2_7_EXMPLR ;
   q_2_6 <= q_2_6_EXMPLR ;
   q_2_5 <= q_2_5_EXMPLR ;
   q_2_4 <= q_2_4_EXMPLR ;
   q_2_3 <= q_2_3_EXMPLR ;
   q_2_2 <= q_2_2_EXMPLR ;
   q_2_1 <= q_2_1_EXMPLR ;
   q_2_0 <= q_2_0_EXMPLR ;
   q_3_15 <= q_3_15_EXMPLR ;
   q_3_14 <= q_3_14_EXMPLR ;
   q_3_13 <= q_3_13_EXMPLR ;
   q_3_12 <= q_3_12_EXMPLR ;
   q_3_11 <= q_3_11_EXMPLR ;
   q_3_10 <= q_3_10_EXMPLR ;
   q_3_9 <= q_3_9_EXMPLR ;
   q_3_8 <= q_3_8_EXMPLR ;
   q_3_7 <= q_3_7_EXMPLR ;
   q_3_6 <= q_3_6_EXMPLR ;
   q_3_5 <= q_3_5_EXMPLR ;
   q_3_4 <= q_3_4_EXMPLR ;
   q_3_3 <= q_3_3_EXMPLR ;
   q_3_2 <= q_3_2_EXMPLR ;
   q_3_1 <= q_3_1_EXMPLR ;
   q_3_0 <= q_3_0_EXMPLR ;
   q_4_15 <= q_4_15_EXMPLR ;
   q_4_14 <= q_4_14_EXMPLR ;
   q_4_13 <= q_4_13_EXMPLR ;
   q_4_12 <= q_4_12_EXMPLR ;
   q_4_11 <= q_4_11_EXMPLR ;
   q_4_10 <= q_4_10_EXMPLR ;
   q_4_9 <= q_4_9_EXMPLR ;
   q_4_8 <= q_4_8_EXMPLR ;
   q_4_7 <= q_4_7_EXMPLR ;
   q_4_6 <= q_4_6_EXMPLR ;
   q_4_5 <= q_4_5_EXMPLR ;
   q_4_4 <= q_4_4_EXMPLR ;
   q_4_3 <= q_4_3_EXMPLR ;
   q_4_2 <= q_4_2_EXMPLR ;
   q_4_1 <= q_4_1_EXMPLR ;
   q_4_0 <= q_4_0_EXMPLR ;
   gen_regs_4_regi_reg_q_0 : dffr port map ( Q=>q_4_0_EXMPLR, QB=>OPEN, D=>
      nx433, CLK=>nx1492, R=>nx1466);
   ix434 : mux21_ni port map ( Y=>nx433, A0=>q_4_0_EXMPLR, A1=>q_3_0_EXMPLR, 
      S0=>nx1440);
   gen_regs_3_regi_reg_q_0 : dffr port map ( Q=>q_3_0_EXMPLR, QB=>OPEN, D=>
      nx423, CLK=>nx1492, R=>nx1466);
   ix424 : mux21_ni port map ( Y=>nx423, A0=>q_3_0_EXMPLR, A1=>q_2_0_EXMPLR, 
      S0=>nx1440);
   gen_regs_2_regi_reg_q_0 : dffr port map ( Q=>q_2_0_EXMPLR, QB=>OPEN, D=>
      nx413, CLK=>nx1492, R=>nx1466);
   ix414 : mux21_ni port map ( Y=>nx413, A0=>q_2_0_EXMPLR, A1=>q_1_0_EXMPLR, 
      S0=>nx1440);
   gen_regs_1_regi_reg_q_0 : dffr port map ( Q=>q_1_0_EXMPLR, QB=>OPEN, D=>
      nx403, CLK=>nx1492, R=>nx1466);
   ix404 : mux21_ni port map ( Y=>nx403, A0=>q_1_0_EXMPLR, A1=>q_0_0_EXMPLR, 
      S0=>nx1440);
   reg0_reg_q_0 : dffr port map ( Q=>q_0_0_EXMPLR, QB=>OPEN, D=>nx393, CLK=>
      nx1492, R=>nx1466);
   ix394 : mux21_ni port map ( Y=>nx393, A0=>q_0_0_EXMPLR, A1=>d(0), S0=>
      nx1440);
   gen_regs_4_regi_reg_q_1 : dffr port map ( Q=>q_4_1_EXMPLR, QB=>OPEN, D=>
      nx483, CLK=>nx1494, R=>nx1468);
   ix484 : mux21_ni port map ( Y=>nx483, A0=>q_4_1_EXMPLR, A1=>q_3_1_EXMPLR, 
      S0=>nx1442);
   gen_regs_3_regi_reg_q_1 : dffr port map ( Q=>q_3_1_EXMPLR, QB=>OPEN, D=>
      nx473, CLK=>nx1494, R=>nx1468);
   ix474 : mux21_ni port map ( Y=>nx473, A0=>q_3_1_EXMPLR, A1=>q_2_1_EXMPLR, 
      S0=>nx1442);
   gen_regs_2_regi_reg_q_1 : dffr port map ( Q=>q_2_1_EXMPLR, QB=>OPEN, D=>
      nx463, CLK=>nx1494, R=>nx1468);
   ix464 : mux21_ni port map ( Y=>nx463, A0=>q_2_1_EXMPLR, A1=>q_1_1_EXMPLR, 
      S0=>nx1442);
   gen_regs_1_regi_reg_q_1 : dffr port map ( Q=>q_1_1_EXMPLR, QB=>OPEN, D=>
      nx453, CLK=>nx1492, R=>nx1466);
   ix454 : mux21_ni port map ( Y=>nx453, A0=>q_1_1_EXMPLR, A1=>q_0_1_EXMPLR, 
      S0=>nx1440);
   reg0_reg_q_1 : dffr port map ( Q=>q_0_1_EXMPLR, QB=>OPEN, D=>nx443, CLK=>
      nx1492, R=>nx1466);
   ix444 : mux21_ni port map ( Y=>nx443, A0=>q_0_1_EXMPLR, A1=>d(1), S0=>
      nx1440);
   gen_regs_4_regi_reg_q_2 : dffr port map ( Q=>q_4_2_EXMPLR, QB=>OPEN, D=>
      nx533, CLK=>nx1496, R=>nx1470);
   ix534 : mux21_ni port map ( Y=>nx533, A0=>q_4_2_EXMPLR, A1=>q_3_2_EXMPLR, 
      S0=>nx1444);
   gen_regs_3_regi_reg_q_2 : dffr port map ( Q=>q_3_2_EXMPLR, QB=>OPEN, D=>
      nx523, CLK=>nx1494, R=>nx1468);
   ix524 : mux21_ni port map ( Y=>nx523, A0=>q_3_2_EXMPLR, A1=>q_2_2_EXMPLR, 
      S0=>nx1442);
   gen_regs_2_regi_reg_q_2 : dffr port map ( Q=>q_2_2_EXMPLR, QB=>OPEN, D=>
      nx513, CLK=>nx1494, R=>nx1468);
   ix514 : mux21_ni port map ( Y=>nx513, A0=>q_2_2_EXMPLR, A1=>q_1_2_EXMPLR, 
      S0=>nx1442);
   gen_regs_1_regi_reg_q_2 : dffr port map ( Q=>q_1_2_EXMPLR, QB=>OPEN, D=>
      nx503, CLK=>nx1494, R=>nx1468);
   ix504 : mux21_ni port map ( Y=>nx503, A0=>q_1_2_EXMPLR, A1=>q_0_2_EXMPLR, 
      S0=>nx1442);
   reg0_reg_q_2 : dffr port map ( Q=>q_0_2_EXMPLR, QB=>OPEN, D=>nx493, CLK=>
      nx1494, R=>nx1468);
   ix494 : mux21_ni port map ( Y=>nx493, A0=>q_0_2_EXMPLR, A1=>d(2), S0=>
      nx1442);
   gen_regs_4_regi_reg_q_3 : dffr port map ( Q=>q_4_3_EXMPLR, QB=>OPEN, D=>
      nx583, CLK=>nx1496, R=>nx1470);
   ix584 : mux21_ni port map ( Y=>nx583, A0=>q_4_3_EXMPLR, A1=>q_3_3_EXMPLR, 
      S0=>nx1444);
   gen_regs_3_regi_reg_q_3 : dffr port map ( Q=>q_3_3_EXMPLR, QB=>OPEN, D=>
      nx573, CLK=>nx1496, R=>nx1470);
   ix574 : mux21_ni port map ( Y=>nx573, A0=>q_3_3_EXMPLR, A1=>q_2_3_EXMPLR, 
      S0=>nx1444);
   gen_regs_2_regi_reg_q_3 : dffr port map ( Q=>q_2_3_EXMPLR, QB=>OPEN, D=>
      nx563, CLK=>nx1496, R=>nx1470);
   ix564 : mux21_ni port map ( Y=>nx563, A0=>q_2_3_EXMPLR, A1=>q_1_3_EXMPLR, 
      S0=>nx1444);
   gen_regs_1_regi_reg_q_3 : dffr port map ( Q=>q_1_3_EXMPLR, QB=>OPEN, D=>
      nx553, CLK=>nx1496, R=>nx1470);
   ix554 : mux21_ni port map ( Y=>nx553, A0=>q_1_3_EXMPLR, A1=>q_0_3_EXMPLR, 
      S0=>nx1444);
   reg0_reg_q_3 : dffr port map ( Q=>q_0_3_EXMPLR, QB=>OPEN, D=>nx543, CLK=>
      nx1496, R=>nx1470);
   ix544 : mux21_ni port map ( Y=>nx543, A0=>q_0_3_EXMPLR, A1=>d(3), S0=>
      nx1444);
   gen_regs_4_regi_reg_q_4 : dffr port map ( Q=>q_4_4_EXMPLR, QB=>OPEN, D=>
      nx633, CLK=>nx1498, R=>nx1472);
   ix634 : mux21_ni port map ( Y=>nx633, A0=>q_4_4_EXMPLR, A1=>q_3_4_EXMPLR, 
      S0=>nx1446);
   gen_regs_3_regi_reg_q_4 : dffr port map ( Q=>q_3_4_EXMPLR, QB=>OPEN, D=>
      nx623, CLK=>nx1498, R=>nx1472);
   ix624 : mux21_ni port map ( Y=>nx623, A0=>q_3_4_EXMPLR, A1=>q_2_4_EXMPLR, 
      S0=>nx1446);
   gen_regs_2_regi_reg_q_4 : dffr port map ( Q=>q_2_4_EXMPLR, QB=>OPEN, D=>
      nx613, CLK=>nx1498, R=>nx1472);
   ix614 : mux21_ni port map ( Y=>nx613, A0=>q_2_4_EXMPLR, A1=>q_1_4_EXMPLR, 
      S0=>nx1446);
   gen_regs_1_regi_reg_q_4 : dffr port map ( Q=>q_1_4_EXMPLR, QB=>OPEN, D=>
      nx603, CLK=>nx1498, R=>nx1472);
   ix604 : mux21_ni port map ( Y=>nx603, A0=>q_1_4_EXMPLR, A1=>q_0_4_EXMPLR, 
      S0=>nx1446);
   reg0_reg_q_4 : dffr port map ( Q=>q_0_4_EXMPLR, QB=>OPEN, D=>nx593, CLK=>
      nx1496, R=>nx1470);
   ix594 : mux21_ni port map ( Y=>nx593, A0=>q_0_4_EXMPLR, A1=>d(4), S0=>
      nx1444);
   gen_regs_4_regi_reg_q_5 : dffr port map ( Q=>q_4_5_EXMPLR, QB=>OPEN, D=>
      nx683, CLK=>nx1500, R=>nx1474);
   ix684 : mux21_ni port map ( Y=>nx683, A0=>q_4_5_EXMPLR, A1=>q_3_5_EXMPLR, 
      S0=>nx1448);
   gen_regs_3_regi_reg_q_5 : dffr port map ( Q=>q_3_5_EXMPLR, QB=>OPEN, D=>
      nx673, CLK=>nx1500, R=>nx1474);
   ix674 : mux21_ni port map ( Y=>nx673, A0=>q_3_5_EXMPLR, A1=>q_2_5_EXMPLR, 
      S0=>nx1448);
   gen_regs_2_regi_reg_q_5 : dffr port map ( Q=>q_2_5_EXMPLR, QB=>OPEN, D=>
      nx663, CLK=>nx1498, R=>nx1472);
   ix664 : mux21_ni port map ( Y=>nx663, A0=>q_2_5_EXMPLR, A1=>q_1_5_EXMPLR, 
      S0=>nx1446);
   gen_regs_1_regi_reg_q_5 : dffr port map ( Q=>q_1_5_EXMPLR, QB=>OPEN, D=>
      nx653, CLK=>nx1498, R=>nx1472);
   ix654 : mux21_ni port map ( Y=>nx653, A0=>q_1_5_EXMPLR, A1=>q_0_5_EXMPLR, 
      S0=>nx1446);
   reg0_reg_q_5 : dffr port map ( Q=>q_0_5_EXMPLR, QB=>OPEN, D=>nx643, CLK=>
      nx1498, R=>nx1472);
   ix644 : mux21_ni port map ( Y=>nx643, A0=>q_0_5_EXMPLR, A1=>d(5), S0=>
      nx1446);
   gen_regs_4_regi_reg_q_6 : dffr port map ( Q=>q_4_6_EXMPLR, QB=>OPEN, D=>
      nx733, CLK=>nx1500, R=>nx1474);
   ix734 : mux21_ni port map ( Y=>nx733, A0=>q_4_6_EXMPLR, A1=>q_3_6_EXMPLR, 
      S0=>nx1448);
   gen_regs_3_regi_reg_q_6 : dffr port map ( Q=>q_3_6_EXMPLR, QB=>OPEN, D=>
      nx723, CLK=>nx1500, R=>nx1474);
   ix724 : mux21_ni port map ( Y=>nx723, A0=>q_3_6_EXMPLR, A1=>q_2_6_EXMPLR, 
      S0=>nx1448);
   gen_regs_2_regi_reg_q_6 : dffr port map ( Q=>q_2_6_EXMPLR, QB=>OPEN, D=>
      nx713, CLK=>nx1500, R=>nx1474);
   ix714 : mux21_ni port map ( Y=>nx713, A0=>q_2_6_EXMPLR, A1=>q_1_6_EXMPLR, 
      S0=>nx1448);
   gen_regs_1_regi_reg_q_6 : dffr port map ( Q=>q_1_6_EXMPLR, QB=>OPEN, D=>
      nx703, CLK=>nx1500, R=>nx1474);
   ix704 : mux21_ni port map ( Y=>nx703, A0=>q_1_6_EXMPLR, A1=>q_0_6_EXMPLR, 
      S0=>nx1448);
   reg0_reg_q_6 : dffr port map ( Q=>q_0_6_EXMPLR, QB=>OPEN, D=>nx693, CLK=>
      nx1500, R=>nx1474);
   ix694 : mux21_ni port map ( Y=>nx693, A0=>q_0_6_EXMPLR, A1=>d(6), S0=>
      nx1448);
   gen_regs_4_regi_reg_q_7 : dffr port map ( Q=>q_4_7_EXMPLR, QB=>OPEN, D=>
      nx783, CLK=>nx1502, R=>nx1476);
   ix784 : mux21_ni port map ( Y=>nx783, A0=>q_4_7_EXMPLR, A1=>q_3_7_EXMPLR, 
      S0=>nx1450);
   gen_regs_3_regi_reg_q_7 : dffr port map ( Q=>q_3_7_EXMPLR, QB=>OPEN, D=>
      nx773, CLK=>nx1502, R=>nx1476);
   ix774 : mux21_ni port map ( Y=>nx773, A0=>q_3_7_EXMPLR, A1=>q_2_7_EXMPLR, 
      S0=>nx1450);
   gen_regs_2_regi_reg_q_7 : dffr port map ( Q=>q_2_7_EXMPLR, QB=>OPEN, D=>
      nx763, CLK=>nx1502, R=>nx1476);
   ix764 : mux21_ni port map ( Y=>nx763, A0=>q_2_7_EXMPLR, A1=>q_1_7_EXMPLR, 
      S0=>nx1450);
   gen_regs_1_regi_reg_q_7 : dffr port map ( Q=>q_1_7_EXMPLR, QB=>OPEN, D=>
      nx753, CLK=>nx1502, R=>nx1476);
   ix754 : mux21_ni port map ( Y=>nx753, A0=>q_1_7_EXMPLR, A1=>q_0_7_EXMPLR, 
      S0=>nx1450);
   reg0_reg_q_7 : dffr port map ( Q=>q_0_7_EXMPLR, QB=>OPEN, D=>nx743, CLK=>
      nx1502, R=>nx1476);
   ix744 : mux21_ni port map ( Y=>nx743, A0=>q_0_7_EXMPLR, A1=>d(7), S0=>
      nx1450);
   gen_regs_4_regi_reg_q_8 : dffr port map ( Q=>q_4_8_EXMPLR, QB=>OPEN, D=>
      nx833, CLK=>nx1504, R=>nx1478);
   ix834 : mux21_ni port map ( Y=>nx833, A0=>q_4_8_EXMPLR, A1=>q_3_8_EXMPLR, 
      S0=>nx1452);
   gen_regs_3_regi_reg_q_8 : dffr port map ( Q=>q_3_8_EXMPLR, QB=>OPEN, D=>
      nx823, CLK=>nx1504, R=>nx1478);
   ix824 : mux21_ni port map ( Y=>nx823, A0=>q_3_8_EXMPLR, A1=>q_2_8_EXMPLR, 
      S0=>nx1452);
   gen_regs_2_regi_reg_q_8 : dffr port map ( Q=>q_2_8_EXMPLR, QB=>OPEN, D=>
      nx813, CLK=>nx1504, R=>nx1478);
   ix814 : mux21_ni port map ( Y=>nx813, A0=>q_2_8_EXMPLR, A1=>q_1_8_EXMPLR, 
      S0=>nx1452);
   gen_regs_1_regi_reg_q_8 : dffr port map ( Q=>q_1_8_EXMPLR, QB=>OPEN, D=>
      nx803, CLK=>nx1502, R=>nx1476);
   ix804 : mux21_ni port map ( Y=>nx803, A0=>q_1_8_EXMPLR, A1=>q_0_8_EXMPLR, 
      S0=>nx1450);
   reg0_reg_q_8 : dffr port map ( Q=>q_0_8_EXMPLR, QB=>OPEN, D=>nx793, CLK=>
      nx1502, R=>nx1476);
   ix794 : mux21_ni port map ( Y=>nx793, A0=>q_0_8_EXMPLR, A1=>d(8), S0=>
      nx1450);
   gen_regs_4_regi_reg_q_9 : dffr port map ( Q=>q_4_9_EXMPLR, QB=>OPEN, D=>
      nx883, CLK=>nx1506, R=>nx1480);
   ix884 : mux21_ni port map ( Y=>nx883, A0=>q_4_9_EXMPLR, A1=>q_3_9_EXMPLR, 
      S0=>nx1454);
   gen_regs_3_regi_reg_q_9 : dffr port map ( Q=>q_3_9_EXMPLR, QB=>OPEN, D=>
      nx873, CLK=>nx1504, R=>nx1478);
   ix874 : mux21_ni port map ( Y=>nx873, A0=>q_3_9_EXMPLR, A1=>q_2_9_EXMPLR, 
      S0=>nx1452);
   gen_regs_2_regi_reg_q_9 : dffr port map ( Q=>q_2_9_EXMPLR, QB=>OPEN, D=>
      nx863, CLK=>nx1504, R=>nx1478);
   ix864 : mux21_ni port map ( Y=>nx863, A0=>q_2_9_EXMPLR, A1=>q_1_9_EXMPLR, 
      S0=>nx1452);
   gen_regs_1_regi_reg_q_9 : dffr port map ( Q=>q_1_9_EXMPLR, QB=>OPEN, D=>
      nx853, CLK=>nx1504, R=>nx1478);
   ix854 : mux21_ni port map ( Y=>nx853, A0=>q_1_9_EXMPLR, A1=>q_0_9_EXMPLR, 
      S0=>nx1452);
   reg0_reg_q_9 : dffr port map ( Q=>q_0_9_EXMPLR, QB=>OPEN, D=>nx843, CLK=>
      nx1504, R=>nx1478);
   ix844 : mux21_ni port map ( Y=>nx843, A0=>q_0_9_EXMPLR, A1=>d(9), S0=>
      nx1452);
   gen_regs_4_regi_reg_q_10 : dffr port map ( Q=>q_4_10_EXMPLR, QB=>OPEN, D
      =>nx933, CLK=>nx1506, R=>nx1480);
   ix934 : mux21_ni port map ( Y=>nx933, A0=>q_4_10_EXMPLR, A1=>
      q_3_10_EXMPLR, S0=>nx1454);
   gen_regs_3_regi_reg_q_10 : dffr port map ( Q=>q_3_10_EXMPLR, QB=>OPEN, D
      =>nx923, CLK=>nx1506, R=>nx1480);
   ix924 : mux21_ni port map ( Y=>nx923, A0=>q_3_10_EXMPLR, A1=>
      q_2_10_EXMPLR, S0=>nx1454);
   gen_regs_2_regi_reg_q_10 : dffr port map ( Q=>q_2_10_EXMPLR, QB=>OPEN, D
      =>nx913, CLK=>nx1506, R=>nx1480);
   ix914 : mux21_ni port map ( Y=>nx913, A0=>q_2_10_EXMPLR, A1=>
      q_1_10_EXMPLR, S0=>nx1454);
   gen_regs_1_regi_reg_q_10 : dffr port map ( Q=>q_1_10_EXMPLR, QB=>OPEN, D
      =>nx903, CLK=>nx1506, R=>nx1480);
   ix904 : mux21_ni port map ( Y=>nx903, A0=>q_1_10_EXMPLR, A1=>
      q_0_10_EXMPLR, S0=>nx1454);
   reg0_reg_q_10 : dffr port map ( Q=>q_0_10_EXMPLR, QB=>OPEN, D=>nx893, CLK
      =>nx1506, R=>nx1480);
   ix894 : mux21_ni port map ( Y=>nx893, A0=>q_0_10_EXMPLR, A1=>d(10), S0=>
      nx1454);
   gen_regs_4_regi_reg_q_11 : dffr port map ( Q=>q_4_11_EXMPLR, QB=>OPEN, D
      =>nx983, CLK=>nx1508, R=>nx1482);
   ix984 : mux21_ni port map ( Y=>nx983, A0=>q_4_11_EXMPLR, A1=>
      q_3_11_EXMPLR, S0=>nx1456);
   gen_regs_3_regi_reg_q_11 : dffr port map ( Q=>q_3_11_EXMPLR, QB=>OPEN, D
      =>nx973, CLK=>nx1508, R=>nx1482);
   ix974 : mux21_ni port map ( Y=>nx973, A0=>q_3_11_EXMPLR, A1=>
      q_2_11_EXMPLR, S0=>nx1456);
   gen_regs_2_regi_reg_q_11 : dffr port map ( Q=>q_2_11_EXMPLR, QB=>OPEN, D
      =>nx963, CLK=>nx1508, R=>nx1482);
   ix964 : mux21_ni port map ( Y=>nx963, A0=>q_2_11_EXMPLR, A1=>
      q_1_11_EXMPLR, S0=>nx1456);
   gen_regs_1_regi_reg_q_11 : dffr port map ( Q=>q_1_11_EXMPLR, QB=>OPEN, D
      =>nx953, CLK=>nx1508, R=>nx1482);
   ix954 : mux21_ni port map ( Y=>nx953, A0=>q_1_11_EXMPLR, A1=>
      q_0_11_EXMPLR, S0=>nx1456);
   reg0_reg_q_11 : dffr port map ( Q=>q_0_11_EXMPLR, QB=>OPEN, D=>nx943, CLK
      =>nx1506, R=>nx1480);
   ix944 : mux21_ni port map ( Y=>nx943, A0=>q_0_11_EXMPLR, A1=>d(11), S0=>
      nx1454);
   gen_regs_4_regi_reg_q_12 : dffr port map ( Q=>q_4_12_EXMPLR, QB=>OPEN, D
      =>nx1033, CLK=>nx1510, R=>nx1484);
   ix1034 : mux21_ni port map ( Y=>nx1033, A0=>q_4_12_EXMPLR, A1=>
      q_3_12_EXMPLR, S0=>nx1458);
   gen_regs_3_regi_reg_q_12 : dffr port map ( Q=>q_3_12_EXMPLR, QB=>OPEN, D
      =>nx1023, CLK=>nx1510, R=>nx1484);
   ix1024 : mux21_ni port map ( Y=>nx1023, A0=>q_3_12_EXMPLR, A1=>
      q_2_12_EXMPLR, S0=>nx1458);
   gen_regs_2_regi_reg_q_12 : dffr port map ( Q=>q_2_12_EXMPLR, QB=>OPEN, D
      =>nx1013, CLK=>nx1508, R=>nx1482);
   ix1014 : mux21_ni port map ( Y=>nx1013, A0=>q_2_12_EXMPLR, A1=>
      q_1_12_EXMPLR, S0=>nx1456);
   gen_regs_1_regi_reg_q_12 : dffr port map ( Q=>q_1_12_EXMPLR, QB=>OPEN, D
      =>nx1003, CLK=>nx1508, R=>nx1482);
   ix1004 : mux21_ni port map ( Y=>nx1003, A0=>q_1_12_EXMPLR, A1=>
      q_0_12_EXMPLR, S0=>nx1456);
   reg0_reg_q_12 : dffr port map ( Q=>q_0_12_EXMPLR, QB=>OPEN, D=>nx993, CLK
      =>nx1508, R=>nx1482);
   ix994 : mux21_ni port map ( Y=>nx993, A0=>q_0_12_EXMPLR, A1=>d(12), S0=>
      nx1456);
   gen_regs_4_regi_reg_q_13 : dffr port map ( Q=>q_4_13_EXMPLR, QB=>OPEN, D
      =>nx1083, CLK=>nx1510, R=>nx1484);
   ix1084 : mux21_ni port map ( Y=>nx1083, A0=>q_4_13_EXMPLR, A1=>
      q_3_13_EXMPLR, S0=>nx1458);
   gen_regs_3_regi_reg_q_13 : dffr port map ( Q=>q_3_13_EXMPLR, QB=>OPEN, D
      =>nx1073, CLK=>nx1510, R=>nx1484);
   ix1074 : mux21_ni port map ( Y=>nx1073, A0=>q_3_13_EXMPLR, A1=>
      q_2_13_EXMPLR, S0=>nx1458);
   gen_regs_2_regi_reg_q_13 : dffr port map ( Q=>q_2_13_EXMPLR, QB=>OPEN, D
      =>nx1063, CLK=>nx1510, R=>nx1484);
   ix1064 : mux21_ni port map ( Y=>nx1063, A0=>q_2_13_EXMPLR, A1=>
      q_1_13_EXMPLR, S0=>nx1458);
   gen_regs_1_regi_reg_q_13 : dffr port map ( Q=>q_1_13_EXMPLR, QB=>OPEN, D
      =>nx1053, CLK=>nx1510, R=>nx1484);
   ix1054 : mux21_ni port map ( Y=>nx1053, A0=>q_1_13_EXMPLR, A1=>
      q_0_13_EXMPLR, S0=>nx1458);
   reg0_reg_q_13 : dffr port map ( Q=>q_0_13_EXMPLR, QB=>OPEN, D=>nx1043, 
      CLK=>nx1510, R=>nx1484);
   ix1044 : mux21_ni port map ( Y=>nx1043, A0=>q_0_13_EXMPLR, A1=>d(13), S0
      =>nx1458);
   gen_regs_4_regi_reg_q_14 : dffr port map ( Q=>q_4_14_EXMPLR, QB=>OPEN, D
      =>nx1133, CLK=>nx1512, R=>nx1486);
   ix1134 : mux21_ni port map ( Y=>nx1133, A0=>q_4_14_EXMPLR, A1=>
      q_3_14_EXMPLR, S0=>nx1460);
   gen_regs_3_regi_reg_q_14 : dffr port map ( Q=>q_3_14_EXMPLR, QB=>OPEN, D
      =>nx1123, CLK=>nx1512, R=>nx1486);
   ix1124 : mux21_ni port map ( Y=>nx1123, A0=>q_3_14_EXMPLR, A1=>
      q_2_14_EXMPLR, S0=>nx1460);
   gen_regs_2_regi_reg_q_14 : dffr port map ( Q=>q_2_14_EXMPLR, QB=>OPEN, D
      =>nx1113, CLK=>nx1512, R=>nx1486);
   ix1114 : mux21_ni port map ( Y=>nx1113, A0=>q_2_14_EXMPLR, A1=>
      q_1_14_EXMPLR, S0=>nx1460);
   gen_regs_1_regi_reg_q_14 : dffr port map ( Q=>q_1_14_EXMPLR, QB=>OPEN, D
      =>nx1103, CLK=>nx1512, R=>nx1486);
   ix1104 : mux21_ni port map ( Y=>nx1103, A0=>q_1_14_EXMPLR, A1=>
      q_0_14_EXMPLR, S0=>nx1460);
   reg0_reg_q_14 : dffr port map ( Q=>q_0_14_EXMPLR, QB=>OPEN, D=>nx1093, 
      CLK=>nx1512, R=>nx1486);
   ix1094 : mux21_ni port map ( Y=>nx1093, A0=>q_0_14_EXMPLR, A1=>d(14), S0
      =>nx1460);
   gen_regs_4_regi_reg_q_15 : dffr port map ( Q=>q_4_15_EXMPLR, QB=>OPEN, D
      =>nx1183, CLK=>nx1514, R=>nx1488);
   ix1184 : mux21_ni port map ( Y=>nx1183, A0=>q_4_15_EXMPLR, A1=>
      q_3_15_EXMPLR, S0=>nx1462);
   gen_regs_3_regi_reg_q_15 : dffr port map ( Q=>q_3_15_EXMPLR, QB=>OPEN, D
      =>nx1173, CLK=>nx1514, R=>nx1488);
   ix1174 : mux21_ni port map ( Y=>nx1173, A0=>q_3_15_EXMPLR, A1=>
      q_2_15_EXMPLR, S0=>nx1462);
   gen_regs_2_regi_reg_q_15 : dffr port map ( Q=>q_2_15_EXMPLR, QB=>OPEN, D
      =>nx1163, CLK=>nx1514, R=>nx1488);
   ix1164 : mux21_ni port map ( Y=>nx1163, A0=>q_2_15_EXMPLR, A1=>
      q_1_15_EXMPLR, S0=>nx1462);
   gen_regs_1_regi_reg_q_15 : dffr port map ( Q=>q_1_15_EXMPLR, QB=>OPEN, D
      =>nx1153, CLK=>nx1512, R=>nx1486);
   ix1154 : mux21_ni port map ( Y=>nx1153, A0=>q_1_15_EXMPLR, A1=>
      q_0_15_EXMPLR, S0=>nx1460);
   reg0_reg_q_15 : dffr port map ( Q=>q_0_15_EXMPLR, QB=>OPEN, D=>nx1143, 
      CLK=>nx1512, R=>nx1486);
   ix1144 : mux21_ni port map ( Y=>nx1143, A0=>q_0_15_EXMPLR, A1=>d(15), S0
      =>nx1460);
   ix1439 : inv02 port map ( Y=>nx1440, A=>nx1516);
   ix1441 : inv02 port map ( Y=>nx1442, A=>nx1516);
   ix1443 : inv02 port map ( Y=>nx1444, A=>nx1516);
   ix1445 : inv02 port map ( Y=>nx1446, A=>nx1516);
   ix1447 : inv02 port map ( Y=>nx1448, A=>nx1516);
   ix1449 : inv02 port map ( Y=>nx1450, A=>nx1516);
   ix1451 : inv02 port map ( Y=>nx1452, A=>nx1516);
   ix1453 : inv02 port map ( Y=>nx1454, A=>nx1518);
   ix1455 : inv02 port map ( Y=>nx1456, A=>nx1518);
   ix1457 : inv02 port map ( Y=>nx1458, A=>nx1518);
   ix1459 : inv02 port map ( Y=>nx1460, A=>nx1518);
   ix1461 : inv02 port map ( Y=>nx1462, A=>nx1518);
   ix1465 : inv02 port map ( Y=>nx1466, A=>nx1520);
   ix1467 : inv02 port map ( Y=>nx1468, A=>nx1520);
   ix1469 : inv02 port map ( Y=>nx1470, A=>nx1520);
   ix1471 : inv02 port map ( Y=>nx1472, A=>nx1520);
   ix1473 : inv02 port map ( Y=>nx1474, A=>nx1520);
   ix1475 : inv02 port map ( Y=>nx1476, A=>nx1520);
   ix1477 : inv02 port map ( Y=>nx1478, A=>nx1520);
   ix1479 : inv02 port map ( Y=>nx1480, A=>nx1522);
   ix1481 : inv02 port map ( Y=>nx1482, A=>nx1522);
   ix1483 : inv02 port map ( Y=>nx1484, A=>nx1522);
   ix1485 : inv02 port map ( Y=>nx1486, A=>nx1522);
   ix1487 : inv02 port map ( Y=>nx1488, A=>nx1522);
   ix1491 : inv02 port map ( Y=>nx1492, A=>nx1524);
   ix1493 : inv02 port map ( Y=>nx1494, A=>nx1524);
   ix1495 : inv02 port map ( Y=>nx1496, A=>nx1524);
   ix1497 : inv02 port map ( Y=>nx1498, A=>nx1524);
   ix1499 : inv02 port map ( Y=>nx1500, A=>nx1524);
   ix1501 : inv02 port map ( Y=>nx1502, A=>nx1524);
   ix1503 : inv02 port map ( Y=>nx1504, A=>nx1524);
   ix1505 : inv02 port map ( Y=>nx1506, A=>nx1526);
   ix1507 : inv02 port map ( Y=>nx1508, A=>nx1526);
   ix1509 : inv02 port map ( Y=>nx1510, A=>nx1526);
   ix1511 : inv02 port map ( Y=>nx1512, A=>nx1526);
   ix1513 : inv02 port map ( Y=>nx1514, A=>nx1526);
   ix1515 : inv02 port map ( Y=>nx1516, A=>load);
   ix1517 : inv02 port map ( Y=>nx1518, A=>load);
   ix1519 : inv02 port map ( Y=>nx1520, A=>reset);
   ix1521 : inv02 port map ( Y=>nx1522, A=>reset);
   ix1523 : inv02 port map ( Y=>nx1524, A=>clk);
   ix1525 : inv02 port map ( Y=>nx1526, A=>clk);
end Dataflow ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Cache_5_16_28_5 is
   port (
      in_word : IN std_logic_vector (15 DOWNTO 0) ;
      cache_in_sel : IN std_logic_vector (4 DOWNTO 0) ;
      cache_out_sel : IN std_logic_vector (4 DOWNTO 0) ;
      decoder_enable : IN std_logic ;
      out_column_0_15 : OUT std_logic ;
      out_column_0_14 : OUT std_logic ;
      out_column_0_13 : OUT std_logic ;
      out_column_0_12 : OUT std_logic ;
      out_column_0_11 : OUT std_logic ;
      out_column_0_10 : OUT std_logic ;
      out_column_0_9 : OUT std_logic ;
      out_column_0_8 : OUT std_logic ;
      out_column_0_7 : OUT std_logic ;
      out_column_0_6 : OUT std_logic ;
      out_column_0_5 : OUT std_logic ;
      out_column_0_4 : OUT std_logic ;
      out_column_0_3 : OUT std_logic ;
      out_column_0_2 : OUT std_logic ;
      out_column_0_1 : OUT std_logic ;
      out_column_0_0 : OUT std_logic ;
      out_column_1_15 : OUT std_logic ;
      out_column_1_14 : OUT std_logic ;
      out_column_1_13 : OUT std_logic ;
      out_column_1_12 : OUT std_logic ;
      out_column_1_11 : OUT std_logic ;
      out_column_1_10 : OUT std_logic ;
      out_column_1_9 : OUT std_logic ;
      out_column_1_8 : OUT std_logic ;
      out_column_1_7 : OUT std_logic ;
      out_column_1_6 : OUT std_logic ;
      out_column_1_5 : OUT std_logic ;
      out_column_1_4 : OUT std_logic ;
      out_column_1_3 : OUT std_logic ;
      out_column_1_2 : OUT std_logic ;
      out_column_1_1 : OUT std_logic ;
      out_column_1_0 : OUT std_logic ;
      out_column_2_15 : OUT std_logic ;
      out_column_2_14 : OUT std_logic ;
      out_column_2_13 : OUT std_logic ;
      out_column_2_12 : OUT std_logic ;
      out_column_2_11 : OUT std_logic ;
      out_column_2_10 : OUT std_logic ;
      out_column_2_9 : OUT std_logic ;
      out_column_2_8 : OUT std_logic ;
      out_column_2_7 : OUT std_logic ;
      out_column_2_6 : OUT std_logic ;
      out_column_2_5 : OUT std_logic ;
      out_column_2_4 : OUT std_logic ;
      out_column_2_3 : OUT std_logic ;
      out_column_2_2 : OUT std_logic ;
      out_column_2_1 : OUT std_logic ;
      out_column_2_0 : OUT std_logic ;
      out_column_3_15 : OUT std_logic ;
      out_column_3_14 : OUT std_logic ;
      out_column_3_13 : OUT std_logic ;
      out_column_3_12 : OUT std_logic ;
      out_column_3_11 : OUT std_logic ;
      out_column_3_10 : OUT std_logic ;
      out_column_3_9 : OUT std_logic ;
      out_column_3_8 : OUT std_logic ;
      out_column_3_7 : OUT std_logic ;
      out_column_3_6 : OUT std_logic ;
      out_column_3_5 : OUT std_logic ;
      out_column_3_4 : OUT std_logic ;
      out_column_3_3 : OUT std_logic ;
      out_column_3_2 : OUT std_logic ;
      out_column_3_1 : OUT std_logic ;
      out_column_3_0 : OUT std_logic ;
      out_column_4_15 : OUT std_logic ;
      out_column_4_14 : OUT std_logic ;
      out_column_4_13 : OUT std_logic ;
      out_column_4_12 : OUT std_logic ;
      out_column_4_11 : OUT std_logic ;
      out_column_4_10 : OUT std_logic ;
      out_column_4_9 : OUT std_logic ;
      out_column_4_8 : OUT std_logic ;
      out_column_4_7 : OUT std_logic ;
      out_column_4_6 : OUT std_logic ;
      out_column_4_5 : OUT std_logic ;
      out_column_4_4 : OUT std_logic ;
      out_column_4_3 : OUT std_logic ;
      out_column_4_2 : OUT std_logic ;
      out_column_4_1 : OUT std_logic ;
      out_column_4_0 : OUT std_logic ;
      clk : IN std_logic ;
      reset : IN std_logic) ;
end Cache_5_16_28_5 ;

architecture Dataflow of Cache_5_16_28_5 is
   component Queue_5
      port (
         d : IN std_logic_vector (15 DOWNTO 0) ;
         q_0_15 : OUT std_logic ;
         q_0_14 : OUT std_logic ;
         q_0_13 : OUT std_logic ;
         q_0_12 : OUT std_logic ;
         q_0_11 : OUT std_logic ;
         q_0_10 : OUT std_logic ;
         q_0_9 : OUT std_logic ;
         q_0_8 : OUT std_logic ;
         q_0_7 : OUT std_logic ;
         q_0_6 : OUT std_logic ;
         q_0_5 : OUT std_logic ;
         q_0_4 : OUT std_logic ;
         q_0_3 : OUT std_logic ;
         q_0_2 : OUT std_logic ;
         q_0_1 : OUT std_logic ;
         q_0_0 : OUT std_logic ;
         q_1_15 : OUT std_logic ;
         q_1_14 : OUT std_logic ;
         q_1_13 : OUT std_logic ;
         q_1_12 : OUT std_logic ;
         q_1_11 : OUT std_logic ;
         q_1_10 : OUT std_logic ;
         q_1_9 : OUT std_logic ;
         q_1_8 : OUT std_logic ;
         q_1_7 : OUT std_logic ;
         q_1_6 : OUT std_logic ;
         q_1_5 : OUT std_logic ;
         q_1_4 : OUT std_logic ;
         q_1_3 : OUT std_logic ;
         q_1_2 : OUT std_logic ;
         q_1_1 : OUT std_logic ;
         q_1_0 : OUT std_logic ;
         q_2_15 : OUT std_logic ;
         q_2_14 : OUT std_logic ;
         q_2_13 : OUT std_logic ;
         q_2_12 : OUT std_logic ;
         q_2_11 : OUT std_logic ;
         q_2_10 : OUT std_logic ;
         q_2_9 : OUT std_logic ;
         q_2_8 : OUT std_logic ;
         q_2_7 : OUT std_logic ;
         q_2_6 : OUT std_logic ;
         q_2_5 : OUT std_logic ;
         q_2_4 : OUT std_logic ;
         q_2_3 : OUT std_logic ;
         q_2_2 : OUT std_logic ;
         q_2_1 : OUT std_logic ;
         q_2_0 : OUT std_logic ;
         q_3_15 : OUT std_logic ;
         q_3_14 : OUT std_logic ;
         q_3_13 : OUT std_logic ;
         q_3_12 : OUT std_logic ;
         q_3_11 : OUT std_logic ;
         q_3_10 : OUT std_logic ;
         q_3_9 : OUT std_logic ;
         q_3_8 : OUT std_logic ;
         q_3_7 : OUT std_logic ;
         q_3_6 : OUT std_logic ;
         q_3_5 : OUT std_logic ;
         q_3_4 : OUT std_logic ;
         q_3_3 : OUT std_logic ;
         q_3_2 : OUT std_logic ;
         q_3_1 : OUT std_logic ;
         q_3_0 : OUT std_logic ;
         q_4_15 : OUT std_logic ;
         q_4_14 : OUT std_logic ;
         q_4_13 : OUT std_logic ;
         q_4_12 : OUT std_logic ;
         q_4_11 : OUT std_logic ;
         q_4_10 : OUT std_logic ;
         q_4_9 : OUT std_logic ;
         q_4_8 : OUT std_logic ;
         q_4_7 : OUT std_logic ;
         q_4_6 : OUT std_logic ;
         q_4_5 : OUT std_logic ;
         q_4_4 : OUT std_logic ;
         q_4_3 : OUT std_logic ;
         q_4_2 : OUT std_logic ;
         q_4_1 : OUT std_logic ;
         q_4_0 : OUT std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         reset : IN std_logic) ;
   end component ;
   signal que_out_0_0_15, que_out_0_0_14, que_out_0_0_13, que_out_0_0_12, 
      que_out_0_0_11, que_out_0_0_10, que_out_0_0_9, que_out_0_0_8, 
      que_out_0_0_7, que_out_0_0_6, que_out_0_0_5, que_out_0_0_4, 
      que_out_0_0_3, que_out_0_0_2, que_out_0_0_1, que_out_0_0_0, 
      que_out_0_1_15, que_out_0_1_14, que_out_0_1_13, que_out_0_1_12, 
      que_out_0_1_11, que_out_0_1_10, que_out_0_1_9, que_out_0_1_8, 
      que_out_0_1_7, que_out_0_1_6, que_out_0_1_5, que_out_0_1_4, 
      que_out_0_1_3, que_out_0_1_2, que_out_0_1_1, que_out_0_1_0, 
      que_out_0_2_15, que_out_0_2_14, que_out_0_2_13, que_out_0_2_12, 
      que_out_0_2_11, que_out_0_2_10, que_out_0_2_9, que_out_0_2_8, 
      que_out_0_2_7, que_out_0_2_6, que_out_0_2_5, que_out_0_2_4, 
      que_out_0_2_3, que_out_0_2_2, que_out_0_2_1, que_out_0_2_0, 
      que_out_0_3_15, que_out_0_3_14, que_out_0_3_13, que_out_0_3_12, 
      que_out_0_3_11, que_out_0_3_10, que_out_0_3_9, que_out_0_3_8, 
      que_out_0_3_7, que_out_0_3_6, que_out_0_3_5, que_out_0_3_4, 
      que_out_0_3_3, que_out_0_3_2, que_out_0_3_1, que_out_0_3_0, 
      que_out_0_4_15, que_out_0_4_14, que_out_0_4_13, que_out_0_4_12, 
      que_out_0_4_11, que_out_0_4_10, que_out_0_4_9, que_out_0_4_8, 
      que_out_0_4_7, que_out_0_4_6, que_out_0_4_5, que_out_0_4_4, 
      que_out_0_4_3, que_out_0_4_2, que_out_0_4_1, que_out_0_4_0, 
      que_out_1_0_15, que_out_1_0_14, que_out_1_0_13, que_out_1_0_12, 
      que_out_1_0_11, que_out_1_0_10, que_out_1_0_9, que_out_1_0_8, 
      que_out_1_0_7, que_out_1_0_6, que_out_1_0_5, que_out_1_0_4, 
      que_out_1_0_3, que_out_1_0_2, que_out_1_0_1, que_out_1_0_0, 
      que_out_1_1_15, que_out_1_1_14, que_out_1_1_13, que_out_1_1_12, 
      que_out_1_1_11, que_out_1_1_10, que_out_1_1_9, que_out_1_1_8, 
      que_out_1_1_7, que_out_1_1_6, que_out_1_1_5, que_out_1_1_4, 
      que_out_1_1_3, que_out_1_1_2, que_out_1_1_1, que_out_1_1_0, 
      que_out_1_2_15, que_out_1_2_14, que_out_1_2_13, que_out_1_2_12, 
      que_out_1_2_11, que_out_1_2_10, que_out_1_2_9, que_out_1_2_8, 
      que_out_1_2_7, que_out_1_2_6, que_out_1_2_5, que_out_1_2_4, 
      que_out_1_2_3, que_out_1_2_2, que_out_1_2_1, que_out_1_2_0, 
      que_out_1_3_15, que_out_1_3_14, que_out_1_3_13, que_out_1_3_12, 
      que_out_1_3_11, que_out_1_3_10, que_out_1_3_9, que_out_1_3_8, 
      que_out_1_3_7, que_out_1_3_6, que_out_1_3_5, que_out_1_3_4, 
      que_out_1_3_3, que_out_1_3_2, que_out_1_3_1, que_out_1_3_0, 
      que_out_1_4_15, que_out_1_4_14, que_out_1_4_13, que_out_1_4_12, 
      que_out_1_4_11, que_out_1_4_10, que_out_1_4_9, que_out_1_4_8, 
      que_out_1_4_7, que_out_1_4_6, que_out_1_4_5, que_out_1_4_4, 
      que_out_1_4_3, que_out_1_4_2, que_out_1_4_1, que_out_1_4_0, 
      que_out_2_0_15, que_out_2_0_14, que_out_2_0_13, que_out_2_0_12, 
      que_out_2_0_11, que_out_2_0_10, que_out_2_0_9, que_out_2_0_8, 
      que_out_2_0_7, que_out_2_0_6, que_out_2_0_5, que_out_2_0_4, 
      que_out_2_0_3, que_out_2_0_2, que_out_2_0_1, que_out_2_0_0, 
      que_out_2_1_15, que_out_2_1_14, que_out_2_1_13, que_out_2_1_12, 
      que_out_2_1_11, que_out_2_1_10, que_out_2_1_9, que_out_2_1_8, 
      que_out_2_1_7, que_out_2_1_6, que_out_2_1_5, que_out_2_1_4, 
      que_out_2_1_3, que_out_2_1_2, que_out_2_1_1, que_out_2_1_0, 
      que_out_2_2_15, que_out_2_2_14, que_out_2_2_13, que_out_2_2_12, 
      que_out_2_2_11, que_out_2_2_10, que_out_2_2_9, que_out_2_2_8, 
      que_out_2_2_7, que_out_2_2_6, que_out_2_2_5, que_out_2_2_4, 
      que_out_2_2_3, que_out_2_2_2, que_out_2_2_1, que_out_2_2_0, 
      que_out_2_3_15, que_out_2_3_14, que_out_2_3_13, que_out_2_3_12, 
      que_out_2_3_11, que_out_2_3_10, que_out_2_3_9, que_out_2_3_8, 
      que_out_2_3_7, que_out_2_3_6, que_out_2_3_5, que_out_2_3_4, 
      que_out_2_3_3, que_out_2_3_2, que_out_2_3_1, que_out_2_3_0, 
      que_out_2_4_15, que_out_2_4_14, que_out_2_4_13, que_out_2_4_12, 
      que_out_2_4_11, que_out_2_4_10, que_out_2_4_9, que_out_2_4_8, 
      que_out_2_4_7, que_out_2_4_6, que_out_2_4_5, que_out_2_4_4, 
      que_out_2_4_3, que_out_2_4_2, que_out_2_4_1, que_out_2_4_0, 
      que_out_3_0_15, que_out_3_0_14, que_out_3_0_13, que_out_3_0_12, 
      que_out_3_0_11, que_out_3_0_10, que_out_3_0_9, que_out_3_0_8, 
      que_out_3_0_7, que_out_3_0_6, que_out_3_0_5, que_out_3_0_4, 
      que_out_3_0_3, que_out_3_0_2, que_out_3_0_1, que_out_3_0_0, 
      que_out_3_1_15, que_out_3_1_14, que_out_3_1_13, que_out_3_1_12, 
      que_out_3_1_11, que_out_3_1_10, que_out_3_1_9, que_out_3_1_8, 
      que_out_3_1_7, que_out_3_1_6, que_out_3_1_5, que_out_3_1_4, 
      que_out_3_1_3, que_out_3_1_2, que_out_3_1_1, que_out_3_1_0, 
      que_out_3_2_15, que_out_3_2_14, que_out_3_2_13, que_out_3_2_12, 
      que_out_3_2_11, que_out_3_2_10, que_out_3_2_9, que_out_3_2_8, 
      que_out_3_2_7, que_out_3_2_6, que_out_3_2_5, que_out_3_2_4, 
      que_out_3_2_3, que_out_3_2_2, que_out_3_2_1, que_out_3_2_0, 
      que_out_3_3_15, que_out_3_3_14, que_out_3_3_13, que_out_3_3_12, 
      que_out_3_3_11, que_out_3_3_10, que_out_3_3_9, que_out_3_3_8, 
      que_out_3_3_7, que_out_3_3_6, que_out_3_3_5, que_out_3_3_4, 
      que_out_3_3_3, que_out_3_3_2, que_out_3_3_1, que_out_3_3_0, 
      que_out_3_4_15, que_out_3_4_14, que_out_3_4_13, que_out_3_4_12, 
      que_out_3_4_11, que_out_3_4_10, que_out_3_4_9, que_out_3_4_8, 
      que_out_3_4_7, que_out_3_4_6, que_out_3_4_5, que_out_3_4_4, 
      que_out_3_4_3, que_out_3_4_2, que_out_3_4_1, que_out_3_4_0, 
      que_out_4_0_15, que_out_4_0_14, que_out_4_0_13, que_out_4_0_12, 
      que_out_4_0_11, que_out_4_0_10, que_out_4_0_9, que_out_4_0_8, 
      que_out_4_0_7, que_out_4_0_6, que_out_4_0_5, que_out_4_0_4, 
      que_out_4_0_3, que_out_4_0_2, que_out_4_0_1, que_out_4_0_0, 
      que_out_4_1_15, que_out_4_1_14, que_out_4_1_13, que_out_4_1_12, 
      que_out_4_1_11, que_out_4_1_10, que_out_4_1_9, que_out_4_1_8, 
      que_out_4_1_7, que_out_4_1_6, que_out_4_1_5, que_out_4_1_4, 
      que_out_4_1_3, que_out_4_1_2, que_out_4_1_1, que_out_4_1_0, 
      que_out_4_2_15, que_out_4_2_14, que_out_4_2_13, que_out_4_2_12, 
      que_out_4_2_11, que_out_4_2_10, que_out_4_2_9, que_out_4_2_8, 
      que_out_4_2_7, que_out_4_2_6, que_out_4_2_5, que_out_4_2_4, 
      que_out_4_2_3, que_out_4_2_2, que_out_4_2_1, que_out_4_2_0, 
      que_out_4_3_15, que_out_4_3_14, que_out_4_3_13, que_out_4_3_12, 
      que_out_4_3_11, que_out_4_3_10, que_out_4_3_9, que_out_4_3_8, 
      que_out_4_3_7, que_out_4_3_6, que_out_4_3_5, que_out_4_3_4, 
      que_out_4_3_3, que_out_4_3_2, que_out_4_3_1, que_out_4_3_0, 
      que_out_4_4_15, que_out_4_4_14, que_out_4_4_13, que_out_4_4_12, 
      que_out_4_4_11, que_out_4_4_10, que_out_4_4_9, que_out_4_4_8, 
      que_out_4_4_7, que_out_4_4_6, que_out_4_4_5, que_out_4_4_4, 
      que_out_4_4_3, que_out_4_4_2, que_out_4_4_1, que_out_4_4_0, 
      que_out_5_0_15, que_out_5_0_14, que_out_5_0_13, que_out_5_0_12, 
      que_out_5_0_11, que_out_5_0_10, que_out_5_0_9, que_out_5_0_8, 
      que_out_5_0_7, que_out_5_0_6, que_out_5_0_5, que_out_5_0_4, 
      que_out_5_0_3, que_out_5_0_2, que_out_5_0_1, que_out_5_0_0, 
      que_out_5_1_15, que_out_5_1_14, que_out_5_1_13, que_out_5_1_12, 
      que_out_5_1_11, que_out_5_1_10, que_out_5_1_9, que_out_5_1_8, 
      que_out_5_1_7, que_out_5_1_6, que_out_5_1_5, que_out_5_1_4, 
      que_out_5_1_3, que_out_5_1_2, que_out_5_1_1, que_out_5_1_0, 
      que_out_5_2_15, que_out_5_2_14, que_out_5_2_13, que_out_5_2_12, 
      que_out_5_2_11, que_out_5_2_10, que_out_5_2_9, que_out_5_2_8, 
      que_out_5_2_7, que_out_5_2_6, que_out_5_2_5, que_out_5_2_4, 
      que_out_5_2_3, que_out_5_2_2, que_out_5_2_1, que_out_5_2_0, 
      que_out_5_3_15, que_out_5_3_14, que_out_5_3_13, que_out_5_3_12, 
      que_out_5_3_11, que_out_5_3_10, que_out_5_3_9, que_out_5_3_8, 
      que_out_5_3_7, que_out_5_3_6, que_out_5_3_5, que_out_5_3_4, 
      que_out_5_3_3, que_out_5_3_2, que_out_5_3_1, que_out_5_3_0, 
      que_out_5_4_15, que_out_5_4_14, que_out_5_4_13, que_out_5_4_12, 
      que_out_5_4_11, que_out_5_4_10, que_out_5_4_9, que_out_5_4_8, 
      que_out_5_4_7, que_out_5_4_6, que_out_5_4_5, que_out_5_4_4, 
      que_out_5_4_3, que_out_5_4_2, que_out_5_4_1, que_out_5_4_0, 
      que_out_6_0_15, que_out_6_0_14, que_out_6_0_13, que_out_6_0_12, 
      que_out_6_0_11, que_out_6_0_10, que_out_6_0_9, que_out_6_0_8, 
      que_out_6_0_7, que_out_6_0_6, que_out_6_0_5, que_out_6_0_4, 
      que_out_6_0_3, que_out_6_0_2, que_out_6_0_1, que_out_6_0_0, 
      que_out_6_1_15, que_out_6_1_14, que_out_6_1_13, que_out_6_1_12, 
      que_out_6_1_11, que_out_6_1_10, que_out_6_1_9, que_out_6_1_8, 
      que_out_6_1_7, que_out_6_1_6, que_out_6_1_5, que_out_6_1_4, 
      que_out_6_1_3, que_out_6_1_2, que_out_6_1_1, que_out_6_1_0, 
      que_out_6_2_15, que_out_6_2_14, que_out_6_2_13, que_out_6_2_12, 
      que_out_6_2_11, que_out_6_2_10, que_out_6_2_9, que_out_6_2_8, 
      que_out_6_2_7, que_out_6_2_6, que_out_6_2_5, que_out_6_2_4, 
      que_out_6_2_3, que_out_6_2_2, que_out_6_2_1, que_out_6_2_0, 
      que_out_6_3_15, que_out_6_3_14, que_out_6_3_13, que_out_6_3_12, 
      que_out_6_3_11, que_out_6_3_10, que_out_6_3_9, que_out_6_3_8, 
      que_out_6_3_7, que_out_6_3_6, que_out_6_3_5, que_out_6_3_4, 
      que_out_6_3_3, que_out_6_3_2, que_out_6_3_1, que_out_6_3_0, 
      que_out_6_4_15, que_out_6_4_14, que_out_6_4_13, que_out_6_4_12, 
      que_out_6_4_11, que_out_6_4_10, que_out_6_4_9, que_out_6_4_8, 
      que_out_6_4_7, que_out_6_4_6, que_out_6_4_5, que_out_6_4_4, 
      que_out_6_4_3, que_out_6_4_2, que_out_6_4_1, que_out_6_4_0, 
      que_out_7_0_15, que_out_7_0_14, que_out_7_0_13, que_out_7_0_12, 
      que_out_7_0_11, que_out_7_0_10, que_out_7_0_9, que_out_7_0_8, 
      que_out_7_0_7, que_out_7_0_6, que_out_7_0_5, que_out_7_0_4, 
      que_out_7_0_3, que_out_7_0_2, que_out_7_0_1, que_out_7_0_0, 
      que_out_7_1_15, que_out_7_1_14, que_out_7_1_13, que_out_7_1_12, 
      que_out_7_1_11, que_out_7_1_10, que_out_7_1_9, que_out_7_1_8, 
      que_out_7_1_7, que_out_7_1_6, que_out_7_1_5, que_out_7_1_4, 
      que_out_7_1_3, que_out_7_1_2, que_out_7_1_1, que_out_7_1_0, 
      que_out_7_2_15, que_out_7_2_14, que_out_7_2_13, que_out_7_2_12, 
      que_out_7_2_11, que_out_7_2_10, que_out_7_2_9, que_out_7_2_8, 
      que_out_7_2_7, que_out_7_2_6, que_out_7_2_5, que_out_7_2_4, 
      que_out_7_2_3, que_out_7_2_2, que_out_7_2_1, que_out_7_2_0, 
      que_out_7_3_15, que_out_7_3_14, que_out_7_3_13, que_out_7_3_12, 
      que_out_7_3_11, que_out_7_3_10, que_out_7_3_9, que_out_7_3_8, 
      que_out_7_3_7, que_out_7_3_6, que_out_7_3_5, que_out_7_3_4, 
      que_out_7_3_3, que_out_7_3_2, que_out_7_3_1, que_out_7_3_0, 
      que_out_7_4_15, que_out_7_4_14, que_out_7_4_13, que_out_7_4_12, 
      que_out_7_4_11, que_out_7_4_10, que_out_7_4_9, que_out_7_4_8, 
      que_out_7_4_7, que_out_7_4_6, que_out_7_4_5, que_out_7_4_4, 
      que_out_7_4_3, que_out_7_4_2, que_out_7_4_1, que_out_7_4_0, 
      que_out_8_0_15, que_out_8_0_14, que_out_8_0_13, que_out_8_0_12, 
      que_out_8_0_11, que_out_8_0_10, que_out_8_0_9, que_out_8_0_8, 
      que_out_8_0_7, que_out_8_0_6, que_out_8_0_5, que_out_8_0_4, 
      que_out_8_0_3, que_out_8_0_2, que_out_8_0_1, que_out_8_0_0, 
      que_out_8_1_15, que_out_8_1_14, que_out_8_1_13, que_out_8_1_12, 
      que_out_8_1_11, que_out_8_1_10, que_out_8_1_9, que_out_8_1_8, 
      que_out_8_1_7, que_out_8_1_6, que_out_8_1_5, que_out_8_1_4, 
      que_out_8_1_3, que_out_8_1_2, que_out_8_1_1, que_out_8_1_0, 
      que_out_8_2_15, que_out_8_2_14, que_out_8_2_13, que_out_8_2_12, 
      que_out_8_2_11, que_out_8_2_10, que_out_8_2_9, que_out_8_2_8, 
      que_out_8_2_7, que_out_8_2_6, que_out_8_2_5, que_out_8_2_4, 
      que_out_8_2_3, que_out_8_2_2, que_out_8_2_1, que_out_8_2_0, 
      que_out_8_3_15, que_out_8_3_14, que_out_8_3_13, que_out_8_3_12, 
      que_out_8_3_11, que_out_8_3_10, que_out_8_3_9, que_out_8_3_8, 
      que_out_8_3_7, que_out_8_3_6, que_out_8_3_5, que_out_8_3_4, 
      que_out_8_3_3, que_out_8_3_2, que_out_8_3_1, que_out_8_3_0, 
      que_out_8_4_15, que_out_8_4_14, que_out_8_4_13, que_out_8_4_12, 
      que_out_8_4_11, que_out_8_4_10, que_out_8_4_9, que_out_8_4_8, 
      que_out_8_4_7, que_out_8_4_6, que_out_8_4_5, que_out_8_4_4, 
      que_out_8_4_3, que_out_8_4_2, que_out_8_4_1, que_out_8_4_0, 
      que_out_9_0_15, que_out_9_0_14, que_out_9_0_13, que_out_9_0_12, 
      que_out_9_0_11, que_out_9_0_10, que_out_9_0_9, que_out_9_0_8, 
      que_out_9_0_7, que_out_9_0_6, que_out_9_0_5, que_out_9_0_4, 
      que_out_9_0_3, que_out_9_0_2, que_out_9_0_1, que_out_9_0_0, 
      que_out_9_1_15, que_out_9_1_14, que_out_9_1_13, que_out_9_1_12, 
      que_out_9_1_11, que_out_9_1_10, que_out_9_1_9, que_out_9_1_8, 
      que_out_9_1_7, que_out_9_1_6, que_out_9_1_5, que_out_9_1_4, 
      que_out_9_1_3, que_out_9_1_2, que_out_9_1_1, que_out_9_1_0, 
      que_out_9_2_15, que_out_9_2_14, que_out_9_2_13, que_out_9_2_12, 
      que_out_9_2_11, que_out_9_2_10, que_out_9_2_9, que_out_9_2_8, 
      que_out_9_2_7, que_out_9_2_6, que_out_9_2_5, que_out_9_2_4, 
      que_out_9_2_3, que_out_9_2_2, que_out_9_2_1, que_out_9_2_0, 
      que_out_9_3_15, que_out_9_3_14, que_out_9_3_13, que_out_9_3_12, 
      que_out_9_3_11, que_out_9_3_10, que_out_9_3_9, que_out_9_3_8, 
      que_out_9_3_7, que_out_9_3_6, que_out_9_3_5, que_out_9_3_4, 
      que_out_9_3_3, que_out_9_3_2, que_out_9_3_1, que_out_9_3_0, 
      que_out_9_4_15, que_out_9_4_14, que_out_9_4_13, que_out_9_4_12, 
      que_out_9_4_11, que_out_9_4_10, que_out_9_4_9, que_out_9_4_8, 
      que_out_9_4_7, que_out_9_4_6, que_out_9_4_5, que_out_9_4_4, 
      que_out_9_4_3, que_out_9_4_2, que_out_9_4_1, que_out_9_4_0, 
      que_out_10_0_15, que_out_10_0_14, que_out_10_0_13, que_out_10_0_12, 
      que_out_10_0_11, que_out_10_0_10, que_out_10_0_9, que_out_10_0_8, 
      que_out_10_0_7, que_out_10_0_6, que_out_10_0_5, que_out_10_0_4, 
      que_out_10_0_3, que_out_10_0_2, que_out_10_0_1, que_out_10_0_0, 
      que_out_10_1_15, que_out_10_1_14, que_out_10_1_13, que_out_10_1_12, 
      que_out_10_1_11, que_out_10_1_10, que_out_10_1_9, que_out_10_1_8, 
      que_out_10_1_7, que_out_10_1_6, que_out_10_1_5, que_out_10_1_4, 
      que_out_10_1_3, que_out_10_1_2, que_out_10_1_1, que_out_10_1_0, 
      que_out_10_2_15, que_out_10_2_14, que_out_10_2_13, que_out_10_2_12, 
      que_out_10_2_11, que_out_10_2_10, que_out_10_2_9, que_out_10_2_8, 
      que_out_10_2_7, que_out_10_2_6, que_out_10_2_5, que_out_10_2_4, 
      que_out_10_2_3, que_out_10_2_2, que_out_10_2_1, que_out_10_2_0, 
      que_out_10_3_15, que_out_10_3_14, que_out_10_3_13, que_out_10_3_12, 
      que_out_10_3_11, que_out_10_3_10, que_out_10_3_9, que_out_10_3_8, 
      que_out_10_3_7, que_out_10_3_6, que_out_10_3_5, que_out_10_3_4, 
      que_out_10_3_3, que_out_10_3_2, que_out_10_3_1, que_out_10_3_0, 
      que_out_10_4_15, que_out_10_4_14, que_out_10_4_13, que_out_10_4_12, 
      que_out_10_4_11, que_out_10_4_10, que_out_10_4_9, que_out_10_4_8, 
      que_out_10_4_7, que_out_10_4_6, que_out_10_4_5, que_out_10_4_4, 
      que_out_10_4_3, que_out_10_4_2, que_out_10_4_1, que_out_10_4_0, 
      que_out_11_0_15, que_out_11_0_14, que_out_11_0_13, que_out_11_0_12, 
      que_out_11_0_11, que_out_11_0_10, que_out_11_0_9, que_out_11_0_8, 
      que_out_11_0_7, que_out_11_0_6, que_out_11_0_5, que_out_11_0_4, 
      que_out_11_0_3, que_out_11_0_2, que_out_11_0_1, que_out_11_0_0, 
      que_out_11_1_15, que_out_11_1_14, que_out_11_1_13, que_out_11_1_12, 
      que_out_11_1_11, que_out_11_1_10, que_out_11_1_9, que_out_11_1_8, 
      que_out_11_1_7, que_out_11_1_6, que_out_11_1_5, que_out_11_1_4, 
      que_out_11_1_3, que_out_11_1_2, que_out_11_1_1, que_out_11_1_0, 
      que_out_11_2_15, que_out_11_2_14, que_out_11_2_13, que_out_11_2_12, 
      que_out_11_2_11, que_out_11_2_10, que_out_11_2_9, que_out_11_2_8, 
      que_out_11_2_7, que_out_11_2_6, que_out_11_2_5, que_out_11_2_4, 
      que_out_11_2_3, que_out_11_2_2, que_out_11_2_1, que_out_11_2_0, 
      que_out_11_3_15, que_out_11_3_14, que_out_11_3_13, que_out_11_3_12, 
      que_out_11_3_11, que_out_11_3_10, que_out_11_3_9, que_out_11_3_8, 
      que_out_11_3_7, que_out_11_3_6, que_out_11_3_5, que_out_11_3_4, 
      que_out_11_3_3, que_out_11_3_2, que_out_11_3_1, que_out_11_3_0, 
      que_out_11_4_15, que_out_11_4_14, que_out_11_4_13, que_out_11_4_12, 
      que_out_11_4_11, que_out_11_4_10, que_out_11_4_9, que_out_11_4_8, 
      que_out_11_4_7, que_out_11_4_6, que_out_11_4_5, que_out_11_4_4, 
      que_out_11_4_3, que_out_11_4_2, que_out_11_4_1, que_out_11_4_0, 
      que_out_12_0_15, que_out_12_0_14, que_out_12_0_13, que_out_12_0_12, 
      que_out_12_0_11, que_out_12_0_10, que_out_12_0_9, que_out_12_0_8, 
      que_out_12_0_7, que_out_12_0_6, que_out_12_0_5, que_out_12_0_4, 
      que_out_12_0_3, que_out_12_0_2, que_out_12_0_1, que_out_12_0_0, 
      que_out_12_1_15, que_out_12_1_14, que_out_12_1_13, que_out_12_1_12, 
      que_out_12_1_11, que_out_12_1_10, que_out_12_1_9, que_out_12_1_8, 
      que_out_12_1_7, que_out_12_1_6, que_out_12_1_5, que_out_12_1_4, 
      que_out_12_1_3, que_out_12_1_2, que_out_12_1_1, que_out_12_1_0, 
      que_out_12_2_15, que_out_12_2_14, que_out_12_2_13, que_out_12_2_12, 
      que_out_12_2_11, que_out_12_2_10, que_out_12_2_9, que_out_12_2_8, 
      que_out_12_2_7, que_out_12_2_6, que_out_12_2_5, que_out_12_2_4, 
      que_out_12_2_3, que_out_12_2_2, que_out_12_2_1, que_out_12_2_0, 
      que_out_12_3_15, que_out_12_3_14, que_out_12_3_13, que_out_12_3_12, 
      que_out_12_3_11, que_out_12_3_10, que_out_12_3_9, que_out_12_3_8, 
      que_out_12_3_7, que_out_12_3_6, que_out_12_3_5, que_out_12_3_4, 
      que_out_12_3_3, que_out_12_3_2, que_out_12_3_1, que_out_12_3_0, 
      que_out_12_4_15, que_out_12_4_14, que_out_12_4_13, que_out_12_4_12, 
      que_out_12_4_11, que_out_12_4_10, que_out_12_4_9, que_out_12_4_8, 
      que_out_12_4_7, que_out_12_4_6, que_out_12_4_5, que_out_12_4_4, 
      que_out_12_4_3, que_out_12_4_2, que_out_12_4_1, que_out_12_4_0, 
      que_out_13_0_15, que_out_13_0_14, que_out_13_0_13, que_out_13_0_12, 
      que_out_13_0_11, que_out_13_0_10, que_out_13_0_9, que_out_13_0_8, 
      que_out_13_0_7, que_out_13_0_6, que_out_13_0_5, que_out_13_0_4, 
      que_out_13_0_3, que_out_13_0_2, que_out_13_0_1, que_out_13_0_0, 
      que_out_13_1_15, que_out_13_1_14, que_out_13_1_13, que_out_13_1_12, 
      que_out_13_1_11, que_out_13_1_10, que_out_13_1_9, que_out_13_1_8, 
      que_out_13_1_7, que_out_13_1_6, que_out_13_1_5, que_out_13_1_4, 
      que_out_13_1_3, que_out_13_1_2, que_out_13_1_1, que_out_13_1_0, 
      que_out_13_2_15, que_out_13_2_14, que_out_13_2_13, que_out_13_2_12, 
      que_out_13_2_11, que_out_13_2_10, que_out_13_2_9, que_out_13_2_8, 
      que_out_13_2_7, que_out_13_2_6, que_out_13_2_5, que_out_13_2_4, 
      que_out_13_2_3, que_out_13_2_2, que_out_13_2_1, que_out_13_2_0, 
      que_out_13_3_15, que_out_13_3_14, que_out_13_3_13, que_out_13_3_12, 
      que_out_13_3_11, que_out_13_3_10, que_out_13_3_9, que_out_13_3_8, 
      que_out_13_3_7, que_out_13_3_6, que_out_13_3_5, que_out_13_3_4, 
      que_out_13_3_3, que_out_13_3_2, que_out_13_3_1, que_out_13_3_0, 
      que_out_13_4_15, que_out_13_4_14, que_out_13_4_13, que_out_13_4_12, 
      que_out_13_4_11, que_out_13_4_10, que_out_13_4_9, que_out_13_4_8, 
      que_out_13_4_7, que_out_13_4_6, que_out_13_4_5, que_out_13_4_4, 
      que_out_13_4_3, que_out_13_4_2, que_out_13_4_1, que_out_13_4_0, 
      que_out_14_0_15, que_out_14_0_14, que_out_14_0_13, que_out_14_0_12, 
      que_out_14_0_11, que_out_14_0_10, que_out_14_0_9, que_out_14_0_8, 
      que_out_14_0_7, que_out_14_0_6, que_out_14_0_5, que_out_14_0_4, 
      que_out_14_0_3, que_out_14_0_2, que_out_14_0_1, que_out_14_0_0, 
      que_out_14_1_15, que_out_14_1_14, que_out_14_1_13, que_out_14_1_12, 
      que_out_14_1_11, que_out_14_1_10, que_out_14_1_9, que_out_14_1_8, 
      que_out_14_1_7, que_out_14_1_6, que_out_14_1_5, que_out_14_1_4, 
      que_out_14_1_3, que_out_14_1_2, que_out_14_1_1, que_out_14_1_0, 
      que_out_14_2_15, que_out_14_2_14, que_out_14_2_13, que_out_14_2_12, 
      que_out_14_2_11, que_out_14_2_10, que_out_14_2_9, que_out_14_2_8, 
      que_out_14_2_7, que_out_14_2_6, que_out_14_2_5, que_out_14_2_4, 
      que_out_14_2_3, que_out_14_2_2, que_out_14_2_1, que_out_14_2_0, 
      que_out_14_3_15, que_out_14_3_14, que_out_14_3_13, que_out_14_3_12, 
      que_out_14_3_11, que_out_14_3_10, que_out_14_3_9, que_out_14_3_8, 
      que_out_14_3_7, que_out_14_3_6, que_out_14_3_5, que_out_14_3_4, 
      que_out_14_3_3, que_out_14_3_2, que_out_14_3_1, que_out_14_3_0, 
      que_out_14_4_15, que_out_14_4_14, que_out_14_4_13, que_out_14_4_12, 
      que_out_14_4_11, que_out_14_4_10, que_out_14_4_9, que_out_14_4_8, 
      que_out_14_4_7, que_out_14_4_6, que_out_14_4_5, que_out_14_4_4, 
      que_out_14_4_3, que_out_14_4_2, que_out_14_4_1, que_out_14_4_0, 
      que_out_15_0_15, que_out_15_0_14, que_out_15_0_13, que_out_15_0_12, 
      que_out_15_0_11, que_out_15_0_10, que_out_15_0_9, que_out_15_0_8, 
      que_out_15_0_7, que_out_15_0_6, que_out_15_0_5, que_out_15_0_4, 
      que_out_15_0_3, que_out_15_0_2, que_out_15_0_1, que_out_15_0_0, 
      que_out_15_1_15, que_out_15_1_14, que_out_15_1_13, que_out_15_1_12, 
      que_out_15_1_11, que_out_15_1_10, que_out_15_1_9, que_out_15_1_8, 
      que_out_15_1_7, que_out_15_1_6, que_out_15_1_5, que_out_15_1_4, 
      que_out_15_1_3, que_out_15_1_2, que_out_15_1_1, que_out_15_1_0, 
      que_out_15_2_15, que_out_15_2_14, que_out_15_2_13, que_out_15_2_12, 
      que_out_15_2_11, que_out_15_2_10, que_out_15_2_9, que_out_15_2_8, 
      que_out_15_2_7, que_out_15_2_6, que_out_15_2_5, que_out_15_2_4, 
      que_out_15_2_3, que_out_15_2_2, que_out_15_2_1, que_out_15_2_0, 
      que_out_15_3_15, que_out_15_3_14, que_out_15_3_13, que_out_15_3_12, 
      que_out_15_3_11, que_out_15_3_10, que_out_15_3_9, que_out_15_3_8, 
      que_out_15_3_7, que_out_15_3_6, que_out_15_3_5, que_out_15_3_4, 
      que_out_15_3_3, que_out_15_3_2, que_out_15_3_1, que_out_15_3_0, 
      que_out_15_4_15, que_out_15_4_14, que_out_15_4_13, que_out_15_4_12, 
      que_out_15_4_11, que_out_15_4_10, que_out_15_4_9, que_out_15_4_8, 
      que_out_15_4_7, que_out_15_4_6, que_out_15_4_5, que_out_15_4_4, 
      que_out_15_4_3, que_out_15_4_2, que_out_15_4_1, que_out_15_4_0, 
      que_out_16_0_15, que_out_16_0_14, que_out_16_0_13, que_out_16_0_12, 
      que_out_16_0_11, que_out_16_0_10, que_out_16_0_9, que_out_16_0_8, 
      que_out_16_0_7, que_out_16_0_6, que_out_16_0_5, que_out_16_0_4, 
      que_out_16_0_3, que_out_16_0_2, que_out_16_0_1, que_out_16_0_0, 
      que_out_16_1_15, que_out_16_1_14, que_out_16_1_13, que_out_16_1_12, 
      que_out_16_1_11, que_out_16_1_10, que_out_16_1_9, que_out_16_1_8, 
      que_out_16_1_7, que_out_16_1_6, que_out_16_1_5, que_out_16_1_4, 
      que_out_16_1_3, que_out_16_1_2, que_out_16_1_1, que_out_16_1_0, 
      que_out_16_2_15, que_out_16_2_14, que_out_16_2_13, que_out_16_2_12, 
      que_out_16_2_11, que_out_16_2_10, que_out_16_2_9, que_out_16_2_8, 
      que_out_16_2_7, que_out_16_2_6, que_out_16_2_5, que_out_16_2_4, 
      que_out_16_2_3, que_out_16_2_2, que_out_16_2_1, que_out_16_2_0, 
      que_out_16_3_15, que_out_16_3_14, que_out_16_3_13, que_out_16_3_12, 
      que_out_16_3_11, que_out_16_3_10, que_out_16_3_9, que_out_16_3_8, 
      que_out_16_3_7, que_out_16_3_6, que_out_16_3_5, que_out_16_3_4, 
      que_out_16_3_3, que_out_16_3_2, que_out_16_3_1, que_out_16_3_0, 
      que_out_16_4_15, que_out_16_4_14, que_out_16_4_13, que_out_16_4_12, 
      que_out_16_4_11, que_out_16_4_10, que_out_16_4_9, que_out_16_4_8, 
      que_out_16_4_7, que_out_16_4_6, que_out_16_4_5, que_out_16_4_4, 
      que_out_16_4_3, que_out_16_4_2, que_out_16_4_1, que_out_16_4_0, 
      que_out_17_0_15, que_out_17_0_14, que_out_17_0_13, que_out_17_0_12, 
      que_out_17_0_11, que_out_17_0_10, que_out_17_0_9, que_out_17_0_8, 
      que_out_17_0_7, que_out_17_0_6, que_out_17_0_5, que_out_17_0_4, 
      que_out_17_0_3, que_out_17_0_2, que_out_17_0_1, que_out_17_0_0, 
      que_out_17_1_15, que_out_17_1_14, que_out_17_1_13, que_out_17_1_12, 
      que_out_17_1_11, que_out_17_1_10, que_out_17_1_9, que_out_17_1_8, 
      que_out_17_1_7, que_out_17_1_6, que_out_17_1_5, que_out_17_1_4, 
      que_out_17_1_3, que_out_17_1_2, que_out_17_1_1, que_out_17_1_0, 
      que_out_17_2_15, que_out_17_2_14, que_out_17_2_13, que_out_17_2_12, 
      que_out_17_2_11, que_out_17_2_10, que_out_17_2_9, que_out_17_2_8, 
      que_out_17_2_7, que_out_17_2_6, que_out_17_2_5, que_out_17_2_4, 
      que_out_17_2_3, que_out_17_2_2, que_out_17_2_1, que_out_17_2_0, 
      que_out_17_3_15, que_out_17_3_14, que_out_17_3_13, que_out_17_3_12, 
      que_out_17_3_11, que_out_17_3_10, que_out_17_3_9, que_out_17_3_8, 
      que_out_17_3_7, que_out_17_3_6, que_out_17_3_5, que_out_17_3_4, 
      que_out_17_3_3, que_out_17_3_2, que_out_17_3_1, que_out_17_3_0, 
      que_out_17_4_15, que_out_17_4_14, que_out_17_4_13, que_out_17_4_12, 
      que_out_17_4_11, que_out_17_4_10, que_out_17_4_9, que_out_17_4_8, 
      que_out_17_4_7, que_out_17_4_6, que_out_17_4_5, que_out_17_4_4, 
      que_out_17_4_3, que_out_17_4_2, que_out_17_4_1, que_out_17_4_0, 
      que_out_18_0_15, que_out_18_0_14, que_out_18_0_13, que_out_18_0_12, 
      que_out_18_0_11, que_out_18_0_10, que_out_18_0_9, que_out_18_0_8, 
      que_out_18_0_7, que_out_18_0_6, que_out_18_0_5, que_out_18_0_4, 
      que_out_18_0_3, que_out_18_0_2, que_out_18_0_1, que_out_18_0_0, 
      que_out_18_1_15, que_out_18_1_14, que_out_18_1_13, que_out_18_1_12, 
      que_out_18_1_11, que_out_18_1_10, que_out_18_1_9, que_out_18_1_8, 
      que_out_18_1_7, que_out_18_1_6, que_out_18_1_5, que_out_18_1_4, 
      que_out_18_1_3, que_out_18_1_2, que_out_18_1_1, que_out_18_1_0, 
      que_out_18_2_15, que_out_18_2_14, que_out_18_2_13, que_out_18_2_12, 
      que_out_18_2_11, que_out_18_2_10, que_out_18_2_9, que_out_18_2_8, 
      que_out_18_2_7, que_out_18_2_6, que_out_18_2_5, que_out_18_2_4, 
      que_out_18_2_3, que_out_18_2_2, que_out_18_2_1, que_out_18_2_0, 
      que_out_18_3_15, que_out_18_3_14, que_out_18_3_13, que_out_18_3_12, 
      que_out_18_3_11, que_out_18_3_10, que_out_18_3_9, que_out_18_3_8, 
      que_out_18_3_7, que_out_18_3_6, que_out_18_3_5, que_out_18_3_4, 
      que_out_18_3_3, que_out_18_3_2, que_out_18_3_1, que_out_18_3_0, 
      que_out_18_4_15, que_out_18_4_14, que_out_18_4_13, que_out_18_4_12, 
      que_out_18_4_11, que_out_18_4_10, que_out_18_4_9, que_out_18_4_8, 
      que_out_18_4_7, que_out_18_4_6, que_out_18_4_5, que_out_18_4_4, 
      que_out_18_4_3, que_out_18_4_2, que_out_18_4_1, que_out_18_4_0, 
      que_out_19_0_15, que_out_19_0_14, que_out_19_0_13, que_out_19_0_12, 
      que_out_19_0_11, que_out_19_0_10, que_out_19_0_9, que_out_19_0_8, 
      que_out_19_0_7, que_out_19_0_6, que_out_19_0_5, que_out_19_0_4, 
      que_out_19_0_3, que_out_19_0_2, que_out_19_0_1, que_out_19_0_0, 
      que_out_19_1_15, que_out_19_1_14, que_out_19_1_13, que_out_19_1_12, 
      que_out_19_1_11, que_out_19_1_10, que_out_19_1_9, que_out_19_1_8, 
      que_out_19_1_7, que_out_19_1_6, que_out_19_1_5, que_out_19_1_4, 
      que_out_19_1_3, que_out_19_1_2, que_out_19_1_1, que_out_19_1_0, 
      que_out_19_2_15, que_out_19_2_14, que_out_19_2_13, que_out_19_2_12, 
      que_out_19_2_11, que_out_19_2_10, que_out_19_2_9, que_out_19_2_8, 
      que_out_19_2_7, que_out_19_2_6, que_out_19_2_5, que_out_19_2_4, 
      que_out_19_2_3, que_out_19_2_2, que_out_19_2_1, que_out_19_2_0, 
      que_out_19_3_15, que_out_19_3_14, que_out_19_3_13, que_out_19_3_12, 
      que_out_19_3_11, que_out_19_3_10, que_out_19_3_9, que_out_19_3_8, 
      que_out_19_3_7, que_out_19_3_6, que_out_19_3_5, que_out_19_3_4, 
      que_out_19_3_3, que_out_19_3_2, que_out_19_3_1, que_out_19_3_0, 
      que_out_19_4_15, que_out_19_4_14, que_out_19_4_13, que_out_19_4_12, 
      que_out_19_4_11, que_out_19_4_10, que_out_19_4_9, que_out_19_4_8, 
      que_out_19_4_7, que_out_19_4_6, que_out_19_4_5, que_out_19_4_4, 
      que_out_19_4_3, que_out_19_4_2, que_out_19_4_1, que_out_19_4_0, 
      que_out_20_0_15, que_out_20_0_14, que_out_20_0_13, que_out_20_0_12, 
      que_out_20_0_11, que_out_20_0_10, que_out_20_0_9, que_out_20_0_8, 
      que_out_20_0_7, que_out_20_0_6, que_out_20_0_5, que_out_20_0_4, 
      que_out_20_0_3, que_out_20_0_2, que_out_20_0_1, que_out_20_0_0, 
      que_out_20_1_15, que_out_20_1_14, que_out_20_1_13, que_out_20_1_12, 
      que_out_20_1_11, que_out_20_1_10, que_out_20_1_9, que_out_20_1_8, 
      que_out_20_1_7, que_out_20_1_6, que_out_20_1_5, que_out_20_1_4, 
      que_out_20_1_3, que_out_20_1_2, que_out_20_1_1, que_out_20_1_0, 
      que_out_20_2_15, que_out_20_2_14, que_out_20_2_13, que_out_20_2_12, 
      que_out_20_2_11, que_out_20_2_10, que_out_20_2_9, que_out_20_2_8, 
      que_out_20_2_7, que_out_20_2_6, que_out_20_2_5, que_out_20_2_4, 
      que_out_20_2_3, que_out_20_2_2, que_out_20_2_1, que_out_20_2_0, 
      que_out_20_3_15, que_out_20_3_14, que_out_20_3_13, que_out_20_3_12, 
      que_out_20_3_11, que_out_20_3_10, que_out_20_3_9, que_out_20_3_8, 
      que_out_20_3_7, que_out_20_3_6, que_out_20_3_5, que_out_20_3_4, 
      que_out_20_3_3, que_out_20_3_2, que_out_20_3_1, que_out_20_3_0, 
      que_out_20_4_15, que_out_20_4_14, que_out_20_4_13, que_out_20_4_12, 
      que_out_20_4_11, que_out_20_4_10, que_out_20_4_9, que_out_20_4_8, 
      que_out_20_4_7, que_out_20_4_6, que_out_20_4_5, que_out_20_4_4, 
      que_out_20_4_3, que_out_20_4_2, que_out_20_4_1, que_out_20_4_0, 
      que_out_21_0_15, que_out_21_0_14, que_out_21_0_13, que_out_21_0_12, 
      que_out_21_0_11, que_out_21_0_10, que_out_21_0_9, que_out_21_0_8, 
      que_out_21_0_7, que_out_21_0_6, que_out_21_0_5, que_out_21_0_4, 
      que_out_21_0_3, que_out_21_0_2, que_out_21_0_1, que_out_21_0_0, 
      que_out_21_1_15, que_out_21_1_14, que_out_21_1_13, que_out_21_1_12, 
      que_out_21_1_11, que_out_21_1_10, que_out_21_1_9, que_out_21_1_8, 
      que_out_21_1_7, que_out_21_1_6, que_out_21_1_5, que_out_21_1_4, 
      que_out_21_1_3, que_out_21_1_2, que_out_21_1_1, que_out_21_1_0, 
      que_out_21_2_15, que_out_21_2_14, que_out_21_2_13, que_out_21_2_12, 
      que_out_21_2_11, que_out_21_2_10, que_out_21_2_9, que_out_21_2_8, 
      que_out_21_2_7, que_out_21_2_6, que_out_21_2_5, que_out_21_2_4, 
      que_out_21_2_3, que_out_21_2_2, que_out_21_2_1, que_out_21_2_0, 
      que_out_21_3_15, que_out_21_3_14, que_out_21_3_13, que_out_21_3_12, 
      que_out_21_3_11, que_out_21_3_10, que_out_21_3_9, que_out_21_3_8, 
      que_out_21_3_7, que_out_21_3_6, que_out_21_3_5, que_out_21_3_4, 
      que_out_21_3_3, que_out_21_3_2, que_out_21_3_1, que_out_21_3_0, 
      que_out_21_4_15, que_out_21_4_14, que_out_21_4_13, que_out_21_4_12, 
      que_out_21_4_11, que_out_21_4_10, que_out_21_4_9, que_out_21_4_8, 
      que_out_21_4_7, que_out_21_4_6, que_out_21_4_5, que_out_21_4_4, 
      que_out_21_4_3, que_out_21_4_2, que_out_21_4_1, que_out_21_4_0, 
      que_out_22_0_15, que_out_22_0_14, que_out_22_0_13, que_out_22_0_12, 
      que_out_22_0_11, que_out_22_0_10, que_out_22_0_9, que_out_22_0_8, 
      que_out_22_0_7, que_out_22_0_6, que_out_22_0_5, que_out_22_0_4, 
      que_out_22_0_3, que_out_22_0_2, que_out_22_0_1, que_out_22_0_0, 
      que_out_22_1_15, que_out_22_1_14, que_out_22_1_13, que_out_22_1_12, 
      que_out_22_1_11, que_out_22_1_10, que_out_22_1_9, que_out_22_1_8, 
      que_out_22_1_7, que_out_22_1_6, que_out_22_1_5, que_out_22_1_4, 
      que_out_22_1_3, que_out_22_1_2, que_out_22_1_1, que_out_22_1_0, 
      que_out_22_2_15, que_out_22_2_14, que_out_22_2_13, que_out_22_2_12, 
      que_out_22_2_11, que_out_22_2_10, que_out_22_2_9, que_out_22_2_8, 
      que_out_22_2_7, que_out_22_2_6, que_out_22_2_5, que_out_22_2_4, 
      que_out_22_2_3, que_out_22_2_2, que_out_22_2_1, que_out_22_2_0, 
      que_out_22_3_15, que_out_22_3_14, que_out_22_3_13, que_out_22_3_12, 
      que_out_22_3_11, que_out_22_3_10, que_out_22_3_9, que_out_22_3_8, 
      que_out_22_3_7, que_out_22_3_6, que_out_22_3_5, que_out_22_3_4, 
      que_out_22_3_3, que_out_22_3_2, que_out_22_3_1, que_out_22_3_0, 
      que_out_22_4_15, que_out_22_4_14, que_out_22_4_13, que_out_22_4_12, 
      que_out_22_4_11, que_out_22_4_10, que_out_22_4_9, que_out_22_4_8, 
      que_out_22_4_7, que_out_22_4_6, que_out_22_4_5, que_out_22_4_4, 
      que_out_22_4_3, que_out_22_4_2, que_out_22_4_1, que_out_22_4_0, 
      que_out_23_0_15, que_out_23_0_14, que_out_23_0_13, que_out_23_0_12, 
      que_out_23_0_11, que_out_23_0_10, que_out_23_0_9, que_out_23_0_8, 
      que_out_23_0_7, que_out_23_0_6, que_out_23_0_5, que_out_23_0_4, 
      que_out_23_0_3, que_out_23_0_2, que_out_23_0_1, que_out_23_0_0, 
      que_out_23_1_15, que_out_23_1_14, que_out_23_1_13, que_out_23_1_12, 
      que_out_23_1_11, que_out_23_1_10, que_out_23_1_9, que_out_23_1_8, 
      que_out_23_1_7, que_out_23_1_6, que_out_23_1_5, que_out_23_1_4, 
      que_out_23_1_3, que_out_23_1_2, que_out_23_1_1, que_out_23_1_0, 
      que_out_23_2_15, que_out_23_2_14, que_out_23_2_13, que_out_23_2_12, 
      que_out_23_2_11, que_out_23_2_10, que_out_23_2_9, que_out_23_2_8, 
      que_out_23_2_7, que_out_23_2_6, que_out_23_2_5, que_out_23_2_4, 
      que_out_23_2_3, que_out_23_2_2, que_out_23_2_1, que_out_23_2_0, 
      que_out_23_3_15, que_out_23_3_14, que_out_23_3_13, que_out_23_3_12, 
      que_out_23_3_11, que_out_23_3_10, que_out_23_3_9, que_out_23_3_8, 
      que_out_23_3_7, que_out_23_3_6, que_out_23_3_5, que_out_23_3_4, 
      que_out_23_3_3, que_out_23_3_2, que_out_23_3_1, que_out_23_3_0, 
      que_out_23_4_15, que_out_23_4_14, que_out_23_4_13, que_out_23_4_12, 
      que_out_23_4_11, que_out_23_4_10, que_out_23_4_9, que_out_23_4_8, 
      que_out_23_4_7, que_out_23_4_6, que_out_23_4_5, que_out_23_4_4, 
      que_out_23_4_3, que_out_23_4_2, que_out_23_4_1, que_out_23_4_0, 
      que_out_24_0_15, que_out_24_0_14, que_out_24_0_13, que_out_24_0_12, 
      que_out_24_0_11, que_out_24_0_10, que_out_24_0_9, que_out_24_0_8, 
      que_out_24_0_7, que_out_24_0_6, que_out_24_0_5, que_out_24_0_4, 
      que_out_24_0_3, que_out_24_0_2, que_out_24_0_1, que_out_24_0_0, 
      que_out_24_1_15, que_out_24_1_14, que_out_24_1_13, que_out_24_1_12, 
      que_out_24_1_11, que_out_24_1_10, que_out_24_1_9, que_out_24_1_8, 
      que_out_24_1_7, que_out_24_1_6, que_out_24_1_5, que_out_24_1_4, 
      que_out_24_1_3, que_out_24_1_2, que_out_24_1_1, que_out_24_1_0, 
      que_out_24_2_15, que_out_24_2_14, que_out_24_2_13, que_out_24_2_12, 
      que_out_24_2_11, que_out_24_2_10, que_out_24_2_9, que_out_24_2_8, 
      que_out_24_2_7, que_out_24_2_6, que_out_24_2_5, que_out_24_2_4, 
      que_out_24_2_3, que_out_24_2_2, que_out_24_2_1, que_out_24_2_0, 
      que_out_24_3_15, que_out_24_3_14, que_out_24_3_13, que_out_24_3_12, 
      que_out_24_3_11, que_out_24_3_10, que_out_24_3_9, que_out_24_3_8, 
      que_out_24_3_7, que_out_24_3_6, que_out_24_3_5, que_out_24_3_4, 
      que_out_24_3_3, que_out_24_3_2, que_out_24_3_1, que_out_24_3_0, 
      que_out_24_4_15, que_out_24_4_14, que_out_24_4_13, que_out_24_4_12, 
      que_out_24_4_11, que_out_24_4_10, que_out_24_4_9, que_out_24_4_8, 
      que_out_24_4_7, que_out_24_4_6, que_out_24_4_5, que_out_24_4_4, 
      que_out_24_4_3, que_out_24_4_2, que_out_24_4_1, que_out_24_4_0, 
      que_out_25_0_15, que_out_25_0_14, que_out_25_0_13, que_out_25_0_12, 
      que_out_25_0_11, que_out_25_0_10, que_out_25_0_9, que_out_25_0_8, 
      que_out_25_0_7, que_out_25_0_6, que_out_25_0_5, que_out_25_0_4, 
      que_out_25_0_3, que_out_25_0_2, que_out_25_0_1, que_out_25_0_0, 
      que_out_25_1_15, que_out_25_1_14, que_out_25_1_13, que_out_25_1_12, 
      que_out_25_1_11, que_out_25_1_10, que_out_25_1_9, que_out_25_1_8, 
      que_out_25_1_7, que_out_25_1_6, que_out_25_1_5, que_out_25_1_4, 
      que_out_25_1_3, que_out_25_1_2, que_out_25_1_1, que_out_25_1_0, 
      que_out_25_2_15, que_out_25_2_14, que_out_25_2_13, que_out_25_2_12, 
      que_out_25_2_11, que_out_25_2_10, que_out_25_2_9, que_out_25_2_8, 
      que_out_25_2_7, que_out_25_2_6, que_out_25_2_5, que_out_25_2_4, 
      que_out_25_2_3, que_out_25_2_2, que_out_25_2_1, que_out_25_2_0, 
      que_out_25_3_15, que_out_25_3_14, que_out_25_3_13, que_out_25_3_12, 
      que_out_25_3_11, que_out_25_3_10, que_out_25_3_9, que_out_25_3_8, 
      que_out_25_3_7, que_out_25_3_6, que_out_25_3_5, que_out_25_3_4, 
      que_out_25_3_3, que_out_25_3_2, que_out_25_3_1, que_out_25_3_0, 
      que_out_25_4_15, que_out_25_4_14, que_out_25_4_13, que_out_25_4_12, 
      que_out_25_4_11, que_out_25_4_10, que_out_25_4_9, que_out_25_4_8, 
      que_out_25_4_7, que_out_25_4_6, que_out_25_4_5, que_out_25_4_4, 
      que_out_25_4_3, que_out_25_4_2, que_out_25_4_1, que_out_25_4_0, 
      que_out_26_0_15, que_out_26_0_14, que_out_26_0_13, que_out_26_0_12, 
      que_out_26_0_11, que_out_26_0_10, que_out_26_0_9, que_out_26_0_8, 
      que_out_26_0_7, que_out_26_0_6, que_out_26_0_5, que_out_26_0_4, 
      que_out_26_0_3, que_out_26_0_2, que_out_26_0_1, que_out_26_0_0, 
      que_out_26_1_15, que_out_26_1_14, que_out_26_1_13, que_out_26_1_12, 
      que_out_26_1_11, que_out_26_1_10, que_out_26_1_9, que_out_26_1_8, 
      que_out_26_1_7, que_out_26_1_6, que_out_26_1_5, que_out_26_1_4, 
      que_out_26_1_3, que_out_26_1_2, que_out_26_1_1, que_out_26_1_0, 
      que_out_26_2_15, que_out_26_2_14, que_out_26_2_13, que_out_26_2_12, 
      que_out_26_2_11, que_out_26_2_10, que_out_26_2_9, que_out_26_2_8, 
      que_out_26_2_7, que_out_26_2_6, que_out_26_2_5, que_out_26_2_4, 
      que_out_26_2_3, que_out_26_2_2, que_out_26_2_1, que_out_26_2_0, 
      que_out_26_3_15, que_out_26_3_14, que_out_26_3_13, que_out_26_3_12, 
      que_out_26_3_11, que_out_26_3_10, que_out_26_3_9, que_out_26_3_8, 
      que_out_26_3_7, que_out_26_3_6, que_out_26_3_5, que_out_26_3_4, 
      que_out_26_3_3, que_out_26_3_2, que_out_26_3_1, que_out_26_3_0, 
      que_out_26_4_15, que_out_26_4_14, que_out_26_4_13, que_out_26_4_12, 
      que_out_26_4_11, que_out_26_4_10, que_out_26_4_9, que_out_26_4_8, 
      que_out_26_4_7, que_out_26_4_6, que_out_26_4_5, que_out_26_4_4, 
      que_out_26_4_3, que_out_26_4_2, que_out_26_4_1, que_out_26_4_0, 
      que_out_27_0_15, que_out_27_0_14, que_out_27_0_13, que_out_27_0_12, 
      que_out_27_0_11, que_out_27_0_10, que_out_27_0_9, que_out_27_0_8, 
      que_out_27_0_7, que_out_27_0_6, que_out_27_0_5, que_out_27_0_4, 
      que_out_27_0_3, que_out_27_0_2, que_out_27_0_1, que_out_27_0_0, 
      que_out_27_1_15, que_out_27_1_14, que_out_27_1_13, que_out_27_1_12, 
      que_out_27_1_11, que_out_27_1_10, que_out_27_1_9, que_out_27_1_8, 
      que_out_27_1_7, que_out_27_1_6, que_out_27_1_5, que_out_27_1_4, 
      que_out_27_1_3, que_out_27_1_2, que_out_27_1_1, que_out_27_1_0, 
      que_out_27_2_15, que_out_27_2_14, que_out_27_2_13, que_out_27_2_12, 
      que_out_27_2_11, que_out_27_2_10, que_out_27_2_9, que_out_27_2_8, 
      que_out_27_2_7, que_out_27_2_6, que_out_27_2_5, que_out_27_2_4, 
      que_out_27_2_3, que_out_27_2_2, que_out_27_2_1, que_out_27_2_0, 
      que_out_27_3_15, que_out_27_3_14, que_out_27_3_13, que_out_27_3_12, 
      que_out_27_3_11, que_out_27_3_10, que_out_27_3_9, que_out_27_3_8, 
      que_out_27_3_7, que_out_27_3_6, que_out_27_3_5, que_out_27_3_4, 
      que_out_27_3_3, que_out_27_3_2, que_out_27_3_1, que_out_27_3_0, 
      que_out_27_4_15, que_out_27_4_14, que_out_27_4_13, que_out_27_4_12, 
      que_out_27_4_11, que_out_27_4_10, que_out_27_4_9, que_out_27_4_8, 
      que_out_27_4_7, que_out_27_4_6, que_out_27_4_5, que_out_27_4_4, 
      que_out_27_4_3, que_out_27_4_2, que_out_27_4_1, que_out_27_4_0, 
      sel_que_27, sel_que_26, sel_que_25, sel_que_24, sel_que_23, sel_que_22, 
      sel_que_21, sel_que_20, sel_que_19, sel_que_18, sel_que_17, sel_que_16, 
      sel_que_15, sel_que_14, sel_que_13, sel_que_12, sel_que_11, sel_que_10, 
      sel_que_9, sel_que_8, sel_que_7, sel_que_6, sel_que_5, sel_que_4, 
      sel_que_3, sel_que_2, sel_que_1, sel_que_0, nx12, nx14, nx28, nx30, 
      nx42, nx48, nx62, nx64, nx68, nx74, nx82, nx88, nx90, nx94, nx100, 
      nx104, nx114, nx118, nx122, nx130, nx136, nx144, nx150, nx158, nx166, 
      nx172, nx180, nx188, nx192, nx200, nx206, nx214, nx222, nx226, nx230, 
      nx238, nx268, nx294, nx322, nx348, nx378, nx404, nx432, nx458, nx488, 
      nx514, nx542, nx568, nx598, nx624, nx652, nx678, nx708, nx734, nx762, 
      nx788, nx818, nx844, nx872, nx898, nx928, nx954, nx982, nx1008, nx1038, 
      nx1064, nx1092, nx1118, nx1148, nx1174, nx1202, nx1228, nx1258, nx1284, 
      nx1312, nx1338, nx1368, nx1394, nx1422, nx1448, nx1478, nx1504, nx1532, 
      nx1558, nx1588, nx1614, nx1642, nx1668, nx1698, nx1724, nx1752, nx1778, 
      nx1808, nx1834, nx1862, nx1888, nx1918, nx1944, nx1972, nx1998, nx2028, 
      nx2054, nx2082, nx2108, nx2138, nx2164, nx2192, nx2218, nx2248, nx2274, 
      nx2302, nx2328, nx2358, nx2384, nx2412, nx2438, nx2468, nx2494, nx2522, 
      nx2548, nx2578, nx2604, nx2632, nx2658, nx2688, nx2714, nx2742, nx2768, 
      nx2798, nx2824, nx2852, nx2878, nx2908, nx2934, nx2962, nx2988, nx3018, 
      nx3044, nx3072, nx3098, nx3128, nx3154, nx3182, nx3208, nx3238, nx3264, 
      nx3292, nx3318, nx3348, nx3374, nx3402, nx3428, nx3458, nx3484, nx3512, 
      nx3538, nx3568, nx3594, nx3622, nx3648, nx3678, nx3704, nx3732, nx3758, 
      nx3788, nx3814, nx3842, nx3868, nx3898, nx3924, nx3952, nx3978, nx4008, 
      nx4034, nx4062, nx4088, nx4118, nx4144, nx4172, nx4198, nx4228, nx4254, 
      nx4282, nx4308, nx4338, nx4364, nx4392, nx4418, nx4448, nx4474, nx4502, 
      nx4528, nx4558, nx4584, nx4612, nx4638, nx4668, nx4694, nx4722, nx4748, 
      nx4778, nx4804, nx4832, nx4858, nx4888, nx4914, nx4942, nx4968, nx4998, 
      nx5024, nx5052, nx5078, nx5108, nx5134, nx5162, nx5188, nx5218, nx5244, 
      nx5272, nx5298, nx5328, nx5354, nx5382, nx5408, nx5438, nx5464, nx5492, 
      nx5518, nx5548, nx5574, nx5602, nx5628, nx5658, nx5684, nx5712, nx5738, 
      nx5768, nx5794, nx5822, nx5848, nx5878, nx5904, nx5932, nx5958, nx5988, 
      nx6014, nx6042, nx6068, nx6098, nx6124, nx6152, nx6178, nx6208, nx6234, 
      nx6262, nx6288, nx6318, nx6344, nx6372, nx6398, nx6428, nx6454, nx6482, 
      nx6508, nx6538, nx6564, nx6592, nx6618, nx6648, nx6674, nx6702, nx6728, 
      nx6758, nx6784, nx6812, nx6838, nx6868, nx6894, nx6922, nx6948, nx6978, 
      nx7004, nx7032, nx7058, nx7088, nx7114, nx7142, nx7168, nx7198, nx7224, 
      nx7252, nx7278, nx7308, nx7334, nx7362, nx7388, nx7418, nx7444, nx7472, 
      nx7498, nx7528, nx7554, nx7582, nx7608, nx7638, nx7664, nx7692, nx7718, 
      nx7748, nx7774, nx7802, nx7828, nx7858, nx7884, nx7912, nx7938, nx7968, 
      nx7994, nx8022, nx8048, nx8078, nx8104, nx8132, nx8158, nx8188, nx8214, 
      nx8242, nx8268, nx8298, nx8324, nx8352, nx8378, nx8408, nx8434, nx8462, 
      nx8488, nx8518, nx8544, nx8572, nx8598, nx8628, nx8654, nx8682, nx8708, 
      nx8738, nx8764, nx8792, nx8818, nx8848, nx8874, nx8902, nx8928, nx8938, 
      nx9038, nx6829, nx6833, nx6835, nx6839, nx6843, nx6847, nx6875, nx6885, 
      nx6889, nx6893, nx6897, nx6901, nx6905, nx6915, nx6927, nx6931, nx6933, 
      nx6937, nx6939, nx6943, nx6945, nx6949, nx6951, nx6955, nx6957, nx6961, 
      nx6965, nx6967, nx6971, nx6977, nx6985, nx6991, nx6999, nx7007, nx7017, 
      nx7029, nx7037, nx7043, nx7053, nx7055, nx7057, nx7061, nx7063, nx7065, 
      nx7069, nx7071, nx7073, nx7077, nx7079, nx7081, nx7087, nx7089, nx7091, 
      nx7095, nx7097, nx7099, nx7103, nx7105, nx7107, nx7111, nx7113, nx7115, 
      nx7121, nx7123, nx7125, nx7129, nx7131, nx7133, nx7137, nx7139, nx7141, 
      nx7145, nx7147, nx7149, nx7155, nx7157, nx7159, nx7163, nx7165, nx7167, 
      nx7171, nx7173, nx7175, nx7179, nx7181, nx7183, nx7189, nx7191, nx7193, 
      nx7197, nx7199, nx7201, nx7205, nx7207, nx7209, nx7213, nx7215, nx7217, 
      nx7223, nx7225, nx7227, nx7231, nx7233, nx7235, nx7239, nx7241, nx7243, 
      nx7247, nx7249, nx7251, nx7257, nx7259, nx7261, nx7265, nx7267, nx7269, 
      nx7273, nx7275, nx7277, nx7281, nx7283, nx7285, nx7291, nx7293, nx7295, 
      nx7299, nx7301, nx7303, nx7307, nx7309, nx7311, nx7315, nx7317, nx7319, 
      nx7325, nx7327, nx7329, nx7333, nx7335, nx7337, nx7341, nx7343, nx7345, 
      nx7349, nx7351, nx7353, nx7359, nx7361, nx7363, nx7367, nx7369, nx7371, 
      nx7375, nx7377, nx7379, nx7383, nx7385, nx7387, nx7393, nx7395, nx7397, 
      nx7401, nx7403, nx7405, nx7409, nx7411, nx7413, nx7417, nx7419, nx7421, 
      nx7427, nx7429, nx7431, nx7435, nx7437, nx7439, nx7443, nx7445, nx7447, 
      nx7451, nx7453, nx7455, nx7461, nx7463, nx7465, nx7469, nx7471, nx7473, 
      nx7477, nx7479, nx7481, nx7485, nx7487, nx7489, nx7495, nx7497, nx7499, 
      nx7503, nx7505, nx7507, nx7511, nx7513, nx7515, nx7519, nx7521, nx7523, 
      nx7529, nx7531, nx7533, nx7537, nx7539, nx7541, nx7545, nx7547, nx7549, 
      nx7553, nx7555, nx7557, nx7563, nx7565, nx7567, nx7571, nx7573, nx7575, 
      nx7579, nx7581, nx7583, nx7587, nx7589, nx7591, nx7597, nx7599, nx7601, 
      nx7605, nx7607, nx7609, nx7613, nx7615, nx7617, nx7621, nx7623, nx7625, 
      nx7631, nx7633, nx7635, nx7639, nx7641, nx7643, nx7647, nx7649, nx7651, 
      nx7655, nx7657, nx7659, nx7665, nx7667, nx7669, nx7673, nx7675, nx7677, 
      nx7681, nx7683, nx7685, nx7689, nx7691, nx7693, nx7699, nx7701, nx7703, 
      nx7707, nx7709, nx7711, nx7715, nx7717, nx7719, nx7723, nx7725, nx7727, 
      nx7733, nx7735, nx7737, nx7741, nx7743, nx7745, nx7749, nx7751, nx7753, 
      nx7757, nx7759, nx7761, nx7767, nx7769, nx7771, nx7775, nx7777, nx7779, 
      nx7783, nx7785, nx7787, nx7791, nx7793, nx7795, nx7801, nx7803, nx7805, 
      nx7809, nx7811, nx7813, nx7817, nx7819, nx7821, nx7825, nx7827, nx7829, 
      nx7835, nx7837, nx7839, nx7843, nx7845, nx7847, nx7851, nx7853, nx7855, 
      nx7859, nx7861, nx7863, nx7869, nx7871, nx7873, nx7877, nx7879, nx7881, 
      nx7885, nx7887, nx7889, nx7893, nx7895, nx7897, nx7903, nx7905, nx7907, 
      nx7911, nx7913, nx7915, nx7919, nx7921, nx7923, nx7927, nx7929, nx7931, 
      nx7937, nx7939, nx7941, nx7945, nx7947, nx7949, nx7953, nx7955, nx7957, 
      nx7961, nx7963, nx7965, nx7971, nx7973, nx7975, nx7979, nx7981, nx7983, 
      nx7987, nx7989, nx7991, nx7995, nx7997, nx7999, nx8005, nx8007, nx8009, 
      nx8013, nx8015, nx8017, nx8021, nx8023, nx8025, nx8029, nx8031, nx8033, 
      nx8039, nx8041, nx8043, nx8047, nx8049, nx8051, nx8055, nx8057, nx8059, 
      nx8063, nx8065, nx8067, nx8073, nx8075, nx8077, nx8081, nx8083, nx8085, 
      nx8089, nx8091, nx8093, nx8097, nx8099, nx8101, nx8107, nx8109, nx8111, 
      nx8115, nx8117, nx8119, nx8123, nx8125, nx8127, nx8131, nx8133, nx8135, 
      nx8141, nx8143, nx8145, nx8149, nx8151, nx8153, nx8157, nx8159, nx8161, 
      nx8165, nx8167, nx8169, nx8175, nx8177, nx8179, nx8183, nx8185, nx8187, 
      nx8191, nx8193, nx8195, nx8199, nx8201, nx8203, nx8209, nx8211, nx8213, 
      nx8217, nx8219, nx8221, nx8225, nx8227, nx8229, nx8233, nx8235, nx8237, 
      nx8243, nx8245, nx8247, nx8251, nx8253, nx8255, nx8259, nx8261, nx8263, 
      nx8267, nx8269, nx8271, nx8277, nx8279, nx8281, nx8285, nx8287, nx8289, 
      nx8293, nx8295, nx8297, nx8301, nx8303, nx8305, nx8311, nx8313, nx8315, 
      nx8319, nx8321, nx8323, nx8327, nx8329, nx8331, nx8335, nx8337, nx8339, 
      nx8345, nx8347, nx8349, nx8353, nx8355, nx8357, nx8361, nx8363, nx8365, 
      nx8369, nx8371, nx8373, nx8379, nx8381, nx8383, nx8387, nx8389, nx8391, 
      nx8395, nx8397, nx8399, nx8403, nx8405, nx8407, nx8413, nx8415, nx8417, 
      nx8421, nx8423, nx8425, nx8429, nx8431, nx8433, nx8437, nx8439, nx8441, 
      nx8447, nx8449, nx8451, nx8455, nx8457, nx8459, nx8463, nx8465, nx8467, 
      nx8471, nx8473, nx8475, nx8481, nx8483, nx8485, nx8489, nx8491, nx8493, 
      nx8497, nx8499, nx8501, nx8505, nx8507, nx8509, nx8515, nx8517, nx8519, 
      nx8523, nx8525, nx8527, nx8531, nx8533, nx8535, nx8539, nx8541, nx8543, 
      nx8549, nx8551, nx8553, nx8557, nx8559, nx8561, nx8565, nx8567, nx8569, 
      nx8573, nx8575, nx8577, nx8583, nx8585, nx8587, nx8591, nx8593, nx8595, 
      nx8599, nx8601, nx8603, nx8607, nx8609, nx8611, nx8617, nx8619, nx8621, 
      nx8625, nx8627, nx8629, nx8633, nx8635, nx8637, nx8641, nx8643, nx8645, 
      nx8651, nx8653, nx8655, nx8659, nx8661, nx8663, nx8667, nx8669, nx8671, 
      nx8675, nx8677, nx8679, nx8685, nx8687, nx8689, nx8693, nx8695, nx8697, 
      nx8701, nx8703, nx8705, nx8709, nx8711, nx8713, nx8719, nx8721, nx8723, 
      nx8727, nx8729, nx8731, nx8735, nx8737, nx8739, nx8743, nx8745, nx8747, 
      nx8753, nx8755, nx8757, nx8761, nx8763, nx8765, nx8769, nx8771, nx8773, 
      nx8777, nx8779, nx8781, nx8787, nx8789, nx8791, nx8795, nx8797, nx8799, 
      nx8803, nx8805, nx8807, nx8811, nx8813, nx8815, nx8821, nx8823, nx8825, 
      nx8829, nx8831, nx8833, nx8837, nx8839, nx8841, nx8845, nx8847, nx8849, 
      nx8855, nx8857, nx8859, nx8863, nx8865, nx8867, nx8871, nx8873, nx8875, 
      nx8879, nx8881, nx8883, nx8889, nx8891, nx8893, nx8897, nx8899, nx8901, 
      nx8905, nx8907, nx8909, nx8913, nx8915, nx8917, nx8923, nx8925, nx8927, 
      nx8931, nx8933, nx8935, nx8939, nx8941, nx8943, nx8947, nx8949, nx8951, 
      nx8955, nx8957, nx8959, nx8963, nx8965, nx8967, nx8970, nx8973, nx8975, 
      nx8978, nx8981, nx8983, nx8989, nx8991, nx8993, nx8997, nx8999, nx9001, 
      nx9005, nx9007, nx9009, nx9013, nx9015, nx9017, nx9023, nx9025, nx9027, 
      nx9031, nx9033, nx9035, nx9039, nx9041, nx9043, nx9047, nx9049, nx9051, 
      nx9057, nx9059, nx9061, nx9065, nx9067, nx9069, nx9073, nx9075, nx9077, 
      nx9081, nx9083, nx9085, nx9090, nx9093, nx9095, nx9098, nx9101, nx9103, 
      nx9106, nx9108, nx9110, nx9113, nx9115, nx9117, nx9121, nx9123, nx9125, 
      nx9128, nx9130, nx9132, nx9135, nx9137, nx9139, nx9142, nx9144, nx9146, 
      nx9150, nx9152, nx9154, nx9157, nx9159, nx9161, nx9164, nx9166, nx9168, 
      nx9171, nx9173, nx9175, nx9179, nx9181, nx9183, nx9186, nx9188, nx9190, 
      nx9193, nx9195, nx9197, nx9200, nx9202, nx9204, nx9208, nx9210, nx9212, 
      nx9215, nx9217, nx9219, nx9222, nx9224, nx9226, nx9229, nx9231, nx9233, 
      nx9237, nx9239, nx9241, nx9244, nx9246, nx9248, nx9251, nx9253, nx9255, 
      nx9258, nx9260, nx9262, nx9266, nx9268, nx9270, nx9273, nx9275, nx9277, 
      nx9280, nx9282, nx9284, nx9287, nx9289, nx9291, nx9295, nx9297, nx9299, 
      nx9302, nx9304, nx9306, nx9309, nx9311, nx9313, nx9316, nx9318, nx9320, 
      nx9324, nx9326, nx9328, nx9331, nx9333, nx9335, nx9338, nx9340, nx9342, 
      nx9345, nx9347, nx9349, nx9353, nx9355, nx9357, nx9360, nx9362, nx9364, 
      nx9367, nx9369, nx9371, nx9374, nx9376, nx9378, nx9382, nx9384, nx9386, 
      nx9389, nx9391, nx9393, nx9396, nx9398, nx9400, nx9403, nx9405, nx9407, 
      nx9411, nx9413, nx9415, nx9418, nx9420, nx9422, nx9425, nx9427, nx9429, 
      nx9432, nx9434, nx9436, nx9440, nx9442, nx9444, nx9447, nx9449, nx9451, 
      nx9454, nx9456, nx9458, nx9461, nx9463, nx9465, nx9469, nx9471, nx9473, 
      nx9476, nx9478, nx9480, nx9483, nx9485, nx9487, nx9490, nx9492, nx9494, 
      nx9498, nx9500, nx9502, nx9505, nx9507, nx9509, nx9512, nx9514, nx9516, 
      nx9519, nx9521, nx9523, nx9527, nx9529, nx9531, nx9534, nx9536, nx9538, 
      nx9541, nx9543, nx9545, nx9548, nx9550, nx9552, nx9556, nx9558, nx9560, 
      nx9563, nx9565, nx9567, nx9570, nx9572, nx9574, nx9577, nx9579, nx9581, 
      nx9585, nx9587, nx9589, nx9592, nx9594, nx9596, nx9599, nx9601, nx9603, 
      nx9606, nx9608, nx9610, nx9614, nx9616, nx9618, nx9621, nx9623, nx9625, 
      nx9628, nx9630, nx9632, nx9635, nx9637, nx9639, nx9648, nx9650, nx9652, 
      nx9654, nx9656, nx9658, nx9660, nx9662, nx9664, nx9666, nx9668, nx9670, 
      nx9674, nx9676, nx9678, nx9680, nx9682, nx9684, nx9686, nx9688, nx9690, 
      nx9692, nx9694, nx9696, nx9700, nx9702, nx9704, nx9706, nx9708, nx9710, 
      nx9712, nx9714, nx9716, nx9718, nx9720, nx9722, nx9726, nx9728, nx9730, 
      nx9732, nx9734, nx9736, nx9738, nx9740, nx9742, nx9744, nx9746, nx9748, 
      nx9752, nx9754, nx9756, nx9758, nx9760, nx9762, nx9764, nx9766, nx9768, 
      nx9770, nx9772, nx9774, nx9778, nx9780, nx9782, nx9784, nx9786, nx9788, 
      nx9790, nx9792, nx9794, nx9796, nx9798, nx9800, nx9804, nx9806, nx9808, 
      nx9810, nx9812, nx9814, nx9816, nx9818, nx9820, nx9822, nx9824, nx9826, 
      nx9830, nx9832, nx9834, nx9836, nx9838, nx9840, nx9842, nx9844, nx9846, 
      nx9848, nx9850, nx9852, nx9856, nx9858, nx9860, nx9862, nx9864, nx9866, 
      nx9868, nx9870, nx9872, nx9874, nx9876, nx9878, nx9882, nx9884, nx9886, 
      nx9888, nx9890, nx9892, nx9894, nx9896, nx9898, nx9900, nx9902, nx9904, 
      nx9908, nx9910, nx9912, nx9914, nx9916, nx9918, nx9920, nx9922, nx9924, 
      nx9926, nx9928, nx9930, nx9934, nx9936, nx9938, nx9940, nx9942, nx9944, 
      nx9946, nx9948, nx9950, nx9952, nx9954, nx9956, nx9960, nx9962, nx9964, 
      nx9966, nx9968, nx9970, nx9972, nx9974, nx9976, nx9978, nx9980, nx9982, 
      nx9986, nx9988, nx9990, nx9992, nx9994, nx9996, nx9998, nx10000, 
      nx10002, nx10004, nx10006, nx10008, nx10012, nx10014, nx10016, nx10018, 
      nx10020, nx10022, nx10024, nx10026, nx10028, nx10030, nx10032, nx10034, 
      nx10038, nx10040, nx10042, nx10044, nx10046, nx10048, nx10050, nx10052, 
      nx10054, nx10056, nx10058, nx10060, nx10064, nx10066, nx10068, nx10070, 
      nx10072, nx10074, nx10076, nx10078, nx10080, nx10082, nx10084, nx10086, 
      nx10090, nx10092, nx10094, nx10096, nx10098, nx10100, nx10102, nx10104, 
      nx10106, nx10108, nx10110, nx10112, nx10116, nx10118, nx10120, nx10122, 
      nx10124, nx10126, nx10128, nx10130, nx10132, nx10134, nx10136, nx10138, 
      nx10142, nx10144, nx10146, nx10148, nx10150, nx10152, nx10154, nx10156, 
      nx10158, nx10160, nx10162, nx10164, nx10168, nx10170, nx10172, nx10174, 
      nx10176, nx10178, nx10180, nx10182, nx10184, nx10186, nx10188, nx10190, 
      nx10194, nx10196, nx10198, nx10200, nx10202, nx10204, nx10206, nx10208, 
      nx10210, nx10212, nx10214, nx10216, nx10220, nx10222, nx10224, nx10226, 
      nx10228, nx10230, nx10232, nx10234, nx10236, nx10238, nx10240, nx10242, 
      nx10246, nx10248, nx10250, nx10252, nx10254, nx10256, nx10258, nx10260, 
      nx10262, nx10264, nx10266, nx10268, nx10272, nx10274, nx10276, nx10278, 
      nx10280, nx10282, nx10284, nx10286, nx10288, nx10290, nx10292, nx10294, 
      nx10298, nx10300, nx10302, nx10304, nx10306, nx10308, nx10310, nx10312, 
      nx10314, nx10316, nx10318, nx10320, nx10324, nx10326, nx10328, nx10330, 
      nx10332, nx10334, nx10336, nx10338, nx10340, nx10342, nx10344, nx10346, 
      nx10350, nx10352, nx10354, nx10356, nx10358, nx10360, nx10362, nx10364, 
      nx10366, nx10368, nx10370, nx10372, nx10374, nx10376, nx10378, nx10380, 
      nx10382, nx10384, nx10386, nx10388, nx10390, nx10392, nx10394, nx10396, 
      nx10398, nx10400, nx10402, nx10404, nx10406, nx10408, nx10410, nx10412, 
      nx10414, nx10416, nx10418, nx10420, nx10422, nx10424, nx10426, nx10428, 
      nx10430, nx10432, nx10434, nx10436, nx10438, nx10440, nx10442, nx10444, 
      nx10446, nx10448, nx10450, nx10452, nx10454, nx10456, nx10458, nx10460, 
      nx10462, nx10464, nx10466, nx10468, nx10470, nx10472, nx10474, nx10476, 
      nx10478, nx10480, nx10482, nx10484, nx10486, nx10488, nx10494, nx10496, 
      nx10498, nx10500, nx10502, nx10504, nx10506, nx10508, nx10510, nx10512, 
      nx10514, nx10516, nx10518, nx10520, nx10522, nx10524, nx10526, nx10528, 
      nx10530, nx10532, nx10534, nx10536, nx10538, nx10540, nx10542, nx10544, 
      nx10546, nx10548, nx10550, nx10552, nx10554, nx10556, nx10558, nx10560, 
      nx10562, nx10564, nx10566, nx10568, nx10570, nx10572, nx10574, nx10576, 
      nx10578, nx10580, nx10582, nx10584, nx10586, nx10588, nx10590, nx10592, 
      nx10594, nx10596, nx10598, nx10600, nx10602, nx10604, nx10606, nx10608, 
      nx10610, nx10612, nx10614, nx10616, nx10618, nx10620, nx10622, nx10624, 
      nx10626, nx10628, nx10630, nx10632, nx10634, nx10636, nx10638, nx10640, 
      nx10642, nx10644, nx10646, nx10648, nx10650, nx10652, nx10654, nx10656, 
      nx10658, nx10660, nx10662, nx10664, nx10666, nx10668, nx10690, nx10692, 
      nx10694, nx10696, nx10698, nx10700, nx10702, nx10704, nx10706, nx10708, 
      nx10710, nx10712, nx10714, nx10716, nx10718, nx10720, nx10722, nx10724, 
      nx10726, nx10728, nx10730, nx10732, nx10734, nx10736, nx10742, nx10744, 
      nx10746, nx10748: std_logic ;

begin
   gen_queues_0_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_0_0_15, q_0_14=>que_out_0_0_14, q_0_13=>
      que_out_0_0_13, q_0_12=>que_out_0_0_12, q_0_11=>que_out_0_0_11, q_0_10
      =>que_out_0_0_10, q_0_9=>que_out_0_0_9, q_0_8=>que_out_0_0_8, q_0_7=>
      que_out_0_0_7, q_0_6=>que_out_0_0_6, q_0_5=>que_out_0_0_5, q_0_4=>
      que_out_0_0_4, q_0_3=>que_out_0_0_3, q_0_2=>que_out_0_0_2, q_0_1=>
      que_out_0_0_1, q_0_0=>que_out_0_0_0, q_1_15=>que_out_0_1_15, q_1_14=>
      que_out_0_1_14, q_1_13=>que_out_0_1_13, q_1_12=>que_out_0_1_12, q_1_11
      =>que_out_0_1_11, q_1_10=>que_out_0_1_10, q_1_9=>que_out_0_1_9, q_1_8
      =>que_out_0_1_8, q_1_7=>que_out_0_1_7, q_1_6=>que_out_0_1_6, q_1_5=>
      que_out_0_1_5, q_1_4=>que_out_0_1_4, q_1_3=>que_out_0_1_3, q_1_2=>
      que_out_0_1_2, q_1_1=>que_out_0_1_1, q_1_0=>que_out_0_1_0, q_2_15=>
      que_out_0_2_15, q_2_14=>que_out_0_2_14, q_2_13=>que_out_0_2_13, q_2_12
      =>que_out_0_2_12, q_2_11=>que_out_0_2_11, q_2_10=>que_out_0_2_10, 
      q_2_9=>que_out_0_2_9, q_2_8=>que_out_0_2_8, q_2_7=>que_out_0_2_7, 
      q_2_6=>que_out_0_2_6, q_2_5=>que_out_0_2_5, q_2_4=>que_out_0_2_4, 
      q_2_3=>que_out_0_2_3, q_2_2=>que_out_0_2_2, q_2_1=>que_out_0_2_1, 
      q_2_0=>que_out_0_2_0, q_3_15=>que_out_0_3_15, q_3_14=>que_out_0_3_14, 
      q_3_13=>que_out_0_3_13, q_3_12=>que_out_0_3_12, q_3_11=>que_out_0_3_11, 
      q_3_10=>que_out_0_3_10, q_3_9=>que_out_0_3_9, q_3_8=>que_out_0_3_8, 
      q_3_7=>que_out_0_3_7, q_3_6=>que_out_0_3_6, q_3_5=>que_out_0_3_5, 
      q_3_4=>que_out_0_3_4, q_3_3=>que_out_0_3_3, q_3_2=>que_out_0_3_2, 
      q_3_1=>que_out_0_3_1, q_3_0=>que_out_0_3_0, q_4_15=>que_out_0_4_15, 
      q_4_14=>que_out_0_4_14, q_4_13=>que_out_0_4_13, q_4_12=>que_out_0_4_12, 
      q_4_11=>que_out_0_4_11, q_4_10=>que_out_0_4_10, q_4_9=>que_out_0_4_9, 
      q_4_8=>que_out_0_4_8, q_4_7=>que_out_0_4_7, q_4_6=>que_out_0_4_6, 
      q_4_5=>que_out_0_4_5, q_4_4=>que_out_0_4_4, q_4_3=>que_out_0_4_3, 
      q_4_2=>que_out_0_4_2, q_4_1=>que_out_0_4_1, q_4_0=>que_out_0_4_0, clk
      =>nx10714, load=>sel_que_0, reset=>nx10690);
   gen_queues_1_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_1_0_15, q_0_14=>que_out_1_0_14, q_0_13=>
      que_out_1_0_13, q_0_12=>que_out_1_0_12, q_0_11=>que_out_1_0_11, q_0_10
      =>que_out_1_0_10, q_0_9=>que_out_1_0_9, q_0_8=>que_out_1_0_8, q_0_7=>
      que_out_1_0_7, q_0_6=>que_out_1_0_6, q_0_5=>que_out_1_0_5, q_0_4=>
      que_out_1_0_4, q_0_3=>que_out_1_0_3, q_0_2=>que_out_1_0_2, q_0_1=>
      que_out_1_0_1, q_0_0=>que_out_1_0_0, q_1_15=>que_out_1_1_15, q_1_14=>
      que_out_1_1_14, q_1_13=>que_out_1_1_13, q_1_12=>que_out_1_1_12, q_1_11
      =>que_out_1_1_11, q_1_10=>que_out_1_1_10, q_1_9=>que_out_1_1_9, q_1_8
      =>que_out_1_1_8, q_1_7=>que_out_1_1_7, q_1_6=>que_out_1_1_6, q_1_5=>
      que_out_1_1_5, q_1_4=>que_out_1_1_4, q_1_3=>que_out_1_1_3, q_1_2=>
      que_out_1_1_2, q_1_1=>que_out_1_1_1, q_1_0=>que_out_1_1_0, q_2_15=>
      que_out_1_2_15, q_2_14=>que_out_1_2_14, q_2_13=>que_out_1_2_13, q_2_12
      =>que_out_1_2_12, q_2_11=>que_out_1_2_11, q_2_10=>que_out_1_2_10, 
      q_2_9=>que_out_1_2_9, q_2_8=>que_out_1_2_8, q_2_7=>que_out_1_2_7, 
      q_2_6=>que_out_1_2_6, q_2_5=>que_out_1_2_5, q_2_4=>que_out_1_2_4, 
      q_2_3=>que_out_1_2_3, q_2_2=>que_out_1_2_2, q_2_1=>que_out_1_2_1, 
      q_2_0=>que_out_1_2_0, q_3_15=>que_out_1_3_15, q_3_14=>que_out_1_3_14, 
      q_3_13=>que_out_1_3_13, q_3_12=>que_out_1_3_12, q_3_11=>que_out_1_3_11, 
      q_3_10=>que_out_1_3_10, q_3_9=>que_out_1_3_9, q_3_8=>que_out_1_3_8, 
      q_3_7=>que_out_1_3_7, q_3_6=>que_out_1_3_6, q_3_5=>que_out_1_3_5, 
      q_3_4=>que_out_1_3_4, q_3_3=>que_out_1_3_3, q_3_2=>que_out_1_3_2, 
      q_3_1=>que_out_1_3_1, q_3_0=>que_out_1_3_0, q_4_15=>que_out_1_4_15, 
      q_4_14=>que_out_1_4_14, q_4_13=>que_out_1_4_13, q_4_12=>que_out_1_4_12, 
      q_4_11=>que_out_1_4_11, q_4_10=>que_out_1_4_10, q_4_9=>que_out_1_4_9, 
      q_4_8=>que_out_1_4_8, q_4_7=>que_out_1_4_7, q_4_6=>que_out_1_4_6, 
      q_4_5=>que_out_1_4_5, q_4_4=>que_out_1_4_4, q_4_3=>que_out_1_4_3, 
      q_4_2=>que_out_1_4_2, q_4_1=>que_out_1_4_1, q_4_0=>que_out_1_4_0, clk
      =>nx10714, load=>sel_que_1, reset=>nx10690);
   gen_queues_2_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_2_0_15, q_0_14=>que_out_2_0_14, q_0_13=>
      que_out_2_0_13, q_0_12=>que_out_2_0_12, q_0_11=>que_out_2_0_11, q_0_10
      =>que_out_2_0_10, q_0_9=>que_out_2_0_9, q_0_8=>que_out_2_0_8, q_0_7=>
      que_out_2_0_7, q_0_6=>que_out_2_0_6, q_0_5=>que_out_2_0_5, q_0_4=>
      que_out_2_0_4, q_0_3=>que_out_2_0_3, q_0_2=>que_out_2_0_2, q_0_1=>
      que_out_2_0_1, q_0_0=>que_out_2_0_0, q_1_15=>que_out_2_1_15, q_1_14=>
      que_out_2_1_14, q_1_13=>que_out_2_1_13, q_1_12=>que_out_2_1_12, q_1_11
      =>que_out_2_1_11, q_1_10=>que_out_2_1_10, q_1_9=>que_out_2_1_9, q_1_8
      =>que_out_2_1_8, q_1_7=>que_out_2_1_7, q_1_6=>que_out_2_1_6, q_1_5=>
      que_out_2_1_5, q_1_4=>que_out_2_1_4, q_1_3=>que_out_2_1_3, q_1_2=>
      que_out_2_1_2, q_1_1=>que_out_2_1_1, q_1_0=>que_out_2_1_0, q_2_15=>
      que_out_2_2_15, q_2_14=>que_out_2_2_14, q_2_13=>que_out_2_2_13, q_2_12
      =>que_out_2_2_12, q_2_11=>que_out_2_2_11, q_2_10=>que_out_2_2_10, 
      q_2_9=>que_out_2_2_9, q_2_8=>que_out_2_2_8, q_2_7=>que_out_2_2_7, 
      q_2_6=>que_out_2_2_6, q_2_5=>que_out_2_2_5, q_2_4=>que_out_2_2_4, 
      q_2_3=>que_out_2_2_3, q_2_2=>que_out_2_2_2, q_2_1=>que_out_2_2_1, 
      q_2_0=>que_out_2_2_0, q_3_15=>que_out_2_3_15, q_3_14=>que_out_2_3_14, 
      q_3_13=>que_out_2_3_13, q_3_12=>que_out_2_3_12, q_3_11=>que_out_2_3_11, 
      q_3_10=>que_out_2_3_10, q_3_9=>que_out_2_3_9, q_3_8=>que_out_2_3_8, 
      q_3_7=>que_out_2_3_7, q_3_6=>que_out_2_3_6, q_3_5=>que_out_2_3_5, 
      q_3_4=>que_out_2_3_4, q_3_3=>que_out_2_3_3, q_3_2=>que_out_2_3_2, 
      q_3_1=>que_out_2_3_1, q_3_0=>que_out_2_3_0, q_4_15=>que_out_2_4_15, 
      q_4_14=>que_out_2_4_14, q_4_13=>que_out_2_4_13, q_4_12=>que_out_2_4_12, 
      q_4_11=>que_out_2_4_11, q_4_10=>que_out_2_4_10, q_4_9=>que_out_2_4_9, 
      q_4_8=>que_out_2_4_8, q_4_7=>que_out_2_4_7, q_4_6=>que_out_2_4_6, 
      q_4_5=>que_out_2_4_5, q_4_4=>que_out_2_4_4, q_4_3=>que_out_2_4_3, 
      q_4_2=>que_out_2_4_2, q_4_1=>que_out_2_4_1, q_4_0=>que_out_2_4_0, clk
      =>nx10714, load=>sel_que_2, reset=>nx10690);
   gen_queues_3_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_3_0_15, q_0_14=>que_out_3_0_14, q_0_13=>
      que_out_3_0_13, q_0_12=>que_out_3_0_12, q_0_11=>que_out_3_0_11, q_0_10
      =>que_out_3_0_10, q_0_9=>que_out_3_0_9, q_0_8=>que_out_3_0_8, q_0_7=>
      que_out_3_0_7, q_0_6=>que_out_3_0_6, q_0_5=>que_out_3_0_5, q_0_4=>
      que_out_3_0_4, q_0_3=>que_out_3_0_3, q_0_2=>que_out_3_0_2, q_0_1=>
      que_out_3_0_1, q_0_0=>que_out_3_0_0, q_1_15=>que_out_3_1_15, q_1_14=>
      que_out_3_1_14, q_1_13=>que_out_3_1_13, q_1_12=>que_out_3_1_12, q_1_11
      =>que_out_3_1_11, q_1_10=>que_out_3_1_10, q_1_9=>que_out_3_1_9, q_1_8
      =>que_out_3_1_8, q_1_7=>que_out_3_1_7, q_1_6=>que_out_3_1_6, q_1_5=>
      que_out_3_1_5, q_1_4=>que_out_3_1_4, q_1_3=>que_out_3_1_3, q_1_2=>
      que_out_3_1_2, q_1_1=>que_out_3_1_1, q_1_0=>que_out_3_1_0, q_2_15=>
      que_out_3_2_15, q_2_14=>que_out_3_2_14, q_2_13=>que_out_3_2_13, q_2_12
      =>que_out_3_2_12, q_2_11=>que_out_3_2_11, q_2_10=>que_out_3_2_10, 
      q_2_9=>que_out_3_2_9, q_2_8=>que_out_3_2_8, q_2_7=>que_out_3_2_7, 
      q_2_6=>que_out_3_2_6, q_2_5=>que_out_3_2_5, q_2_4=>que_out_3_2_4, 
      q_2_3=>que_out_3_2_3, q_2_2=>que_out_3_2_2, q_2_1=>que_out_3_2_1, 
      q_2_0=>que_out_3_2_0, q_3_15=>que_out_3_3_15, q_3_14=>que_out_3_3_14, 
      q_3_13=>que_out_3_3_13, q_3_12=>que_out_3_3_12, q_3_11=>que_out_3_3_11, 
      q_3_10=>que_out_3_3_10, q_3_9=>que_out_3_3_9, q_3_8=>que_out_3_3_8, 
      q_3_7=>que_out_3_3_7, q_3_6=>que_out_3_3_6, q_3_5=>que_out_3_3_5, 
      q_3_4=>que_out_3_3_4, q_3_3=>que_out_3_3_3, q_3_2=>que_out_3_3_2, 
      q_3_1=>que_out_3_3_1, q_3_0=>que_out_3_3_0, q_4_15=>que_out_3_4_15, 
      q_4_14=>que_out_3_4_14, q_4_13=>que_out_3_4_13, q_4_12=>que_out_3_4_12, 
      q_4_11=>que_out_3_4_11, q_4_10=>que_out_3_4_10, q_4_9=>que_out_3_4_9, 
      q_4_8=>que_out_3_4_8, q_4_7=>que_out_3_4_7, q_4_6=>que_out_3_4_6, 
      q_4_5=>que_out_3_4_5, q_4_4=>que_out_3_4_4, q_4_3=>que_out_3_4_3, 
      q_4_2=>que_out_3_4_2, q_4_1=>que_out_3_4_1, q_4_0=>que_out_3_4_0, clk
      =>nx10716, load=>sel_que_3, reset=>nx10692);
   gen_queues_4_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_4_0_15, q_0_14=>que_out_4_0_14, q_0_13=>
      que_out_4_0_13, q_0_12=>que_out_4_0_12, q_0_11=>que_out_4_0_11, q_0_10
      =>que_out_4_0_10, q_0_9=>que_out_4_0_9, q_0_8=>que_out_4_0_8, q_0_7=>
      que_out_4_0_7, q_0_6=>que_out_4_0_6, q_0_5=>que_out_4_0_5, q_0_4=>
      que_out_4_0_4, q_0_3=>que_out_4_0_3, q_0_2=>que_out_4_0_2, q_0_1=>
      que_out_4_0_1, q_0_0=>que_out_4_0_0, q_1_15=>que_out_4_1_15, q_1_14=>
      que_out_4_1_14, q_1_13=>que_out_4_1_13, q_1_12=>que_out_4_1_12, q_1_11
      =>que_out_4_1_11, q_1_10=>que_out_4_1_10, q_1_9=>que_out_4_1_9, q_1_8
      =>que_out_4_1_8, q_1_7=>que_out_4_1_7, q_1_6=>que_out_4_1_6, q_1_5=>
      que_out_4_1_5, q_1_4=>que_out_4_1_4, q_1_3=>que_out_4_1_3, q_1_2=>
      que_out_4_1_2, q_1_1=>que_out_4_1_1, q_1_0=>que_out_4_1_0, q_2_15=>
      que_out_4_2_15, q_2_14=>que_out_4_2_14, q_2_13=>que_out_4_2_13, q_2_12
      =>que_out_4_2_12, q_2_11=>que_out_4_2_11, q_2_10=>que_out_4_2_10, 
      q_2_9=>que_out_4_2_9, q_2_8=>que_out_4_2_8, q_2_7=>que_out_4_2_7, 
      q_2_6=>que_out_4_2_6, q_2_5=>que_out_4_2_5, q_2_4=>que_out_4_2_4, 
      q_2_3=>que_out_4_2_3, q_2_2=>que_out_4_2_2, q_2_1=>que_out_4_2_1, 
      q_2_0=>que_out_4_2_0, q_3_15=>que_out_4_3_15, q_3_14=>que_out_4_3_14, 
      q_3_13=>que_out_4_3_13, q_3_12=>que_out_4_3_12, q_3_11=>que_out_4_3_11, 
      q_3_10=>que_out_4_3_10, q_3_9=>que_out_4_3_9, q_3_8=>que_out_4_3_8, 
      q_3_7=>que_out_4_3_7, q_3_6=>que_out_4_3_6, q_3_5=>que_out_4_3_5, 
      q_3_4=>que_out_4_3_4, q_3_3=>que_out_4_3_3, q_3_2=>que_out_4_3_2, 
      q_3_1=>que_out_4_3_1, q_3_0=>que_out_4_3_0, q_4_15=>que_out_4_4_15, 
      q_4_14=>que_out_4_4_14, q_4_13=>que_out_4_4_13, q_4_12=>que_out_4_4_12, 
      q_4_11=>que_out_4_4_11, q_4_10=>que_out_4_4_10, q_4_9=>que_out_4_4_9, 
      q_4_8=>que_out_4_4_8, q_4_7=>que_out_4_4_7, q_4_6=>que_out_4_4_6, 
      q_4_5=>que_out_4_4_5, q_4_4=>que_out_4_4_4, q_4_3=>que_out_4_4_3, 
      q_4_2=>que_out_4_4_2, q_4_1=>que_out_4_4_1, q_4_0=>que_out_4_4_0, clk
      =>nx10716, load=>sel_que_4, reset=>nx10692);
   gen_queues_5_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_5_0_15, q_0_14=>que_out_5_0_14, q_0_13=>
      que_out_5_0_13, q_0_12=>que_out_5_0_12, q_0_11=>que_out_5_0_11, q_0_10
      =>que_out_5_0_10, q_0_9=>que_out_5_0_9, q_0_8=>que_out_5_0_8, q_0_7=>
      que_out_5_0_7, q_0_6=>que_out_5_0_6, q_0_5=>que_out_5_0_5, q_0_4=>
      que_out_5_0_4, q_0_3=>que_out_5_0_3, q_0_2=>que_out_5_0_2, q_0_1=>
      que_out_5_0_1, q_0_0=>que_out_5_0_0, q_1_15=>que_out_5_1_15, q_1_14=>
      que_out_5_1_14, q_1_13=>que_out_5_1_13, q_1_12=>que_out_5_1_12, q_1_11
      =>que_out_5_1_11, q_1_10=>que_out_5_1_10, q_1_9=>que_out_5_1_9, q_1_8
      =>que_out_5_1_8, q_1_7=>que_out_5_1_7, q_1_6=>que_out_5_1_6, q_1_5=>
      que_out_5_1_5, q_1_4=>que_out_5_1_4, q_1_3=>que_out_5_1_3, q_1_2=>
      que_out_5_1_2, q_1_1=>que_out_5_1_1, q_1_0=>que_out_5_1_0, q_2_15=>
      que_out_5_2_15, q_2_14=>que_out_5_2_14, q_2_13=>que_out_5_2_13, q_2_12
      =>que_out_5_2_12, q_2_11=>que_out_5_2_11, q_2_10=>que_out_5_2_10, 
      q_2_9=>que_out_5_2_9, q_2_8=>que_out_5_2_8, q_2_7=>que_out_5_2_7, 
      q_2_6=>que_out_5_2_6, q_2_5=>que_out_5_2_5, q_2_4=>que_out_5_2_4, 
      q_2_3=>que_out_5_2_3, q_2_2=>que_out_5_2_2, q_2_1=>que_out_5_2_1, 
      q_2_0=>que_out_5_2_0, q_3_15=>que_out_5_3_15, q_3_14=>que_out_5_3_14, 
      q_3_13=>que_out_5_3_13, q_3_12=>que_out_5_3_12, q_3_11=>que_out_5_3_11, 
      q_3_10=>que_out_5_3_10, q_3_9=>que_out_5_3_9, q_3_8=>que_out_5_3_8, 
      q_3_7=>que_out_5_3_7, q_3_6=>que_out_5_3_6, q_3_5=>que_out_5_3_5, 
      q_3_4=>que_out_5_3_4, q_3_3=>que_out_5_3_3, q_3_2=>que_out_5_3_2, 
      q_3_1=>que_out_5_3_1, q_3_0=>que_out_5_3_0, q_4_15=>que_out_5_4_15, 
      q_4_14=>que_out_5_4_14, q_4_13=>que_out_5_4_13, q_4_12=>que_out_5_4_12, 
      q_4_11=>que_out_5_4_11, q_4_10=>que_out_5_4_10, q_4_9=>que_out_5_4_9, 
      q_4_8=>que_out_5_4_8, q_4_7=>que_out_5_4_7, q_4_6=>que_out_5_4_6, 
      q_4_5=>que_out_5_4_5, q_4_4=>que_out_5_4_4, q_4_3=>que_out_5_4_3, 
      q_4_2=>que_out_5_4_2, q_4_1=>que_out_5_4_1, q_4_0=>que_out_5_4_0, clk
      =>nx10716, load=>sel_que_5, reset=>nx10692);
   gen_queues_6_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_6_0_15, q_0_14=>que_out_6_0_14, q_0_13=>
      que_out_6_0_13, q_0_12=>que_out_6_0_12, q_0_11=>que_out_6_0_11, q_0_10
      =>que_out_6_0_10, q_0_9=>que_out_6_0_9, q_0_8=>que_out_6_0_8, q_0_7=>
      que_out_6_0_7, q_0_6=>que_out_6_0_6, q_0_5=>que_out_6_0_5, q_0_4=>
      que_out_6_0_4, q_0_3=>que_out_6_0_3, q_0_2=>que_out_6_0_2, q_0_1=>
      que_out_6_0_1, q_0_0=>que_out_6_0_0, q_1_15=>que_out_6_1_15, q_1_14=>
      que_out_6_1_14, q_1_13=>que_out_6_1_13, q_1_12=>que_out_6_1_12, q_1_11
      =>que_out_6_1_11, q_1_10=>que_out_6_1_10, q_1_9=>que_out_6_1_9, q_1_8
      =>que_out_6_1_8, q_1_7=>que_out_6_1_7, q_1_6=>que_out_6_1_6, q_1_5=>
      que_out_6_1_5, q_1_4=>que_out_6_1_4, q_1_3=>que_out_6_1_3, q_1_2=>
      que_out_6_1_2, q_1_1=>que_out_6_1_1, q_1_0=>que_out_6_1_0, q_2_15=>
      que_out_6_2_15, q_2_14=>que_out_6_2_14, q_2_13=>que_out_6_2_13, q_2_12
      =>que_out_6_2_12, q_2_11=>que_out_6_2_11, q_2_10=>que_out_6_2_10, 
      q_2_9=>que_out_6_2_9, q_2_8=>que_out_6_2_8, q_2_7=>que_out_6_2_7, 
      q_2_6=>que_out_6_2_6, q_2_5=>que_out_6_2_5, q_2_4=>que_out_6_2_4, 
      q_2_3=>que_out_6_2_3, q_2_2=>que_out_6_2_2, q_2_1=>que_out_6_2_1, 
      q_2_0=>que_out_6_2_0, q_3_15=>que_out_6_3_15, q_3_14=>que_out_6_3_14, 
      q_3_13=>que_out_6_3_13, q_3_12=>que_out_6_3_12, q_3_11=>que_out_6_3_11, 
      q_3_10=>que_out_6_3_10, q_3_9=>que_out_6_3_9, q_3_8=>que_out_6_3_8, 
      q_3_7=>que_out_6_3_7, q_3_6=>que_out_6_3_6, q_3_5=>que_out_6_3_5, 
      q_3_4=>que_out_6_3_4, q_3_3=>que_out_6_3_3, q_3_2=>que_out_6_3_2, 
      q_3_1=>que_out_6_3_1, q_3_0=>que_out_6_3_0, q_4_15=>que_out_6_4_15, 
      q_4_14=>que_out_6_4_14, q_4_13=>que_out_6_4_13, q_4_12=>que_out_6_4_12, 
      q_4_11=>que_out_6_4_11, q_4_10=>que_out_6_4_10, q_4_9=>que_out_6_4_9, 
      q_4_8=>que_out_6_4_8, q_4_7=>que_out_6_4_7, q_4_6=>que_out_6_4_6, 
      q_4_5=>que_out_6_4_5, q_4_4=>que_out_6_4_4, q_4_3=>que_out_6_4_3, 
      q_4_2=>que_out_6_4_2, q_4_1=>que_out_6_4_1, q_4_0=>que_out_6_4_0, clk
      =>nx10718, load=>sel_que_6, reset=>nx10694);
   gen_queues_7_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_7_0_15, q_0_14=>que_out_7_0_14, q_0_13=>
      que_out_7_0_13, q_0_12=>que_out_7_0_12, q_0_11=>que_out_7_0_11, q_0_10
      =>que_out_7_0_10, q_0_9=>que_out_7_0_9, q_0_8=>que_out_7_0_8, q_0_7=>
      que_out_7_0_7, q_0_6=>que_out_7_0_6, q_0_5=>que_out_7_0_5, q_0_4=>
      que_out_7_0_4, q_0_3=>que_out_7_0_3, q_0_2=>que_out_7_0_2, q_0_1=>
      que_out_7_0_1, q_0_0=>que_out_7_0_0, q_1_15=>que_out_7_1_15, q_1_14=>
      que_out_7_1_14, q_1_13=>que_out_7_1_13, q_1_12=>que_out_7_1_12, q_1_11
      =>que_out_7_1_11, q_1_10=>que_out_7_1_10, q_1_9=>que_out_7_1_9, q_1_8
      =>que_out_7_1_8, q_1_7=>que_out_7_1_7, q_1_6=>que_out_7_1_6, q_1_5=>
      que_out_7_1_5, q_1_4=>que_out_7_1_4, q_1_3=>que_out_7_1_3, q_1_2=>
      que_out_7_1_2, q_1_1=>que_out_7_1_1, q_1_0=>que_out_7_1_0, q_2_15=>
      que_out_7_2_15, q_2_14=>que_out_7_2_14, q_2_13=>que_out_7_2_13, q_2_12
      =>que_out_7_2_12, q_2_11=>que_out_7_2_11, q_2_10=>que_out_7_2_10, 
      q_2_9=>que_out_7_2_9, q_2_8=>que_out_7_2_8, q_2_7=>que_out_7_2_7, 
      q_2_6=>que_out_7_2_6, q_2_5=>que_out_7_2_5, q_2_4=>que_out_7_2_4, 
      q_2_3=>que_out_7_2_3, q_2_2=>que_out_7_2_2, q_2_1=>que_out_7_2_1, 
      q_2_0=>que_out_7_2_0, q_3_15=>que_out_7_3_15, q_3_14=>que_out_7_3_14, 
      q_3_13=>que_out_7_3_13, q_3_12=>que_out_7_3_12, q_3_11=>que_out_7_3_11, 
      q_3_10=>que_out_7_3_10, q_3_9=>que_out_7_3_9, q_3_8=>que_out_7_3_8, 
      q_3_7=>que_out_7_3_7, q_3_6=>que_out_7_3_6, q_3_5=>que_out_7_3_5, 
      q_3_4=>que_out_7_3_4, q_3_3=>que_out_7_3_3, q_3_2=>que_out_7_3_2, 
      q_3_1=>que_out_7_3_1, q_3_0=>que_out_7_3_0, q_4_15=>que_out_7_4_15, 
      q_4_14=>que_out_7_4_14, q_4_13=>que_out_7_4_13, q_4_12=>que_out_7_4_12, 
      q_4_11=>que_out_7_4_11, q_4_10=>que_out_7_4_10, q_4_9=>que_out_7_4_9, 
      q_4_8=>que_out_7_4_8, q_4_7=>que_out_7_4_7, q_4_6=>que_out_7_4_6, 
      q_4_5=>que_out_7_4_5, q_4_4=>que_out_7_4_4, q_4_3=>que_out_7_4_3, 
      q_4_2=>que_out_7_4_2, q_4_1=>que_out_7_4_1, q_4_0=>que_out_7_4_0, clk
      =>nx10720, load=>sel_que_7, reset=>nx10696);
   gen_queues_8_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_8_0_15, q_0_14=>que_out_8_0_14, q_0_13=>
      que_out_8_0_13, q_0_12=>que_out_8_0_12, q_0_11=>que_out_8_0_11, q_0_10
      =>que_out_8_0_10, q_0_9=>que_out_8_0_9, q_0_8=>que_out_8_0_8, q_0_7=>
      que_out_8_0_7, q_0_6=>que_out_8_0_6, q_0_5=>que_out_8_0_5, q_0_4=>
      que_out_8_0_4, q_0_3=>que_out_8_0_3, q_0_2=>que_out_8_0_2, q_0_1=>
      que_out_8_0_1, q_0_0=>que_out_8_0_0, q_1_15=>que_out_8_1_15, q_1_14=>
      que_out_8_1_14, q_1_13=>que_out_8_1_13, q_1_12=>que_out_8_1_12, q_1_11
      =>que_out_8_1_11, q_1_10=>que_out_8_1_10, q_1_9=>que_out_8_1_9, q_1_8
      =>que_out_8_1_8, q_1_7=>que_out_8_1_7, q_1_6=>que_out_8_1_6, q_1_5=>
      que_out_8_1_5, q_1_4=>que_out_8_1_4, q_1_3=>que_out_8_1_3, q_1_2=>
      que_out_8_1_2, q_1_1=>que_out_8_1_1, q_1_0=>que_out_8_1_0, q_2_15=>
      que_out_8_2_15, q_2_14=>que_out_8_2_14, q_2_13=>que_out_8_2_13, q_2_12
      =>que_out_8_2_12, q_2_11=>que_out_8_2_11, q_2_10=>que_out_8_2_10, 
      q_2_9=>que_out_8_2_9, q_2_8=>que_out_8_2_8, q_2_7=>que_out_8_2_7, 
      q_2_6=>que_out_8_2_6, q_2_5=>que_out_8_2_5, q_2_4=>que_out_8_2_4, 
      q_2_3=>que_out_8_2_3, q_2_2=>que_out_8_2_2, q_2_1=>que_out_8_2_1, 
      q_2_0=>que_out_8_2_0, q_3_15=>que_out_8_3_15, q_3_14=>que_out_8_3_14, 
      q_3_13=>que_out_8_3_13, q_3_12=>que_out_8_3_12, q_3_11=>que_out_8_3_11, 
      q_3_10=>que_out_8_3_10, q_3_9=>que_out_8_3_9, q_3_8=>que_out_8_3_8, 
      q_3_7=>que_out_8_3_7, q_3_6=>que_out_8_3_6, q_3_5=>que_out_8_3_5, 
      q_3_4=>que_out_8_3_4, q_3_3=>que_out_8_3_3, q_3_2=>que_out_8_3_2, 
      q_3_1=>que_out_8_3_1, q_3_0=>que_out_8_3_0, q_4_15=>que_out_8_4_15, 
      q_4_14=>que_out_8_4_14, q_4_13=>que_out_8_4_13, q_4_12=>que_out_8_4_12, 
      q_4_11=>que_out_8_4_11, q_4_10=>que_out_8_4_10, q_4_9=>que_out_8_4_9, 
      q_4_8=>que_out_8_4_8, q_4_7=>que_out_8_4_7, q_4_6=>que_out_8_4_6, 
      q_4_5=>que_out_8_4_5, q_4_4=>que_out_8_4_4, q_4_3=>que_out_8_4_3, 
      q_4_2=>que_out_8_4_2, q_4_1=>que_out_8_4_1, q_4_0=>que_out_8_4_0, clk
      =>nx10720, load=>sel_que_8, reset=>nx10696);
   gen_queues_9_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_9_0_15, q_0_14=>que_out_9_0_14, q_0_13=>
      que_out_9_0_13, q_0_12=>que_out_9_0_12, q_0_11=>que_out_9_0_11, q_0_10
      =>que_out_9_0_10, q_0_9=>que_out_9_0_9, q_0_8=>que_out_9_0_8, q_0_7=>
      que_out_9_0_7, q_0_6=>que_out_9_0_6, q_0_5=>que_out_9_0_5, q_0_4=>
      que_out_9_0_4, q_0_3=>que_out_9_0_3, q_0_2=>que_out_9_0_2, q_0_1=>
      que_out_9_0_1, q_0_0=>que_out_9_0_0, q_1_15=>que_out_9_1_15, q_1_14=>
      que_out_9_1_14, q_1_13=>que_out_9_1_13, q_1_12=>que_out_9_1_12, q_1_11
      =>que_out_9_1_11, q_1_10=>que_out_9_1_10, q_1_9=>que_out_9_1_9, q_1_8
      =>que_out_9_1_8, q_1_7=>que_out_9_1_7, q_1_6=>que_out_9_1_6, q_1_5=>
      que_out_9_1_5, q_1_4=>que_out_9_1_4, q_1_3=>que_out_9_1_3, q_1_2=>
      que_out_9_1_2, q_1_1=>que_out_9_1_1, q_1_0=>que_out_9_1_0, q_2_15=>
      que_out_9_2_15, q_2_14=>que_out_9_2_14, q_2_13=>que_out_9_2_13, q_2_12
      =>que_out_9_2_12, q_2_11=>que_out_9_2_11, q_2_10=>que_out_9_2_10, 
      q_2_9=>que_out_9_2_9, q_2_8=>que_out_9_2_8, q_2_7=>que_out_9_2_7, 
      q_2_6=>que_out_9_2_6, q_2_5=>que_out_9_2_5, q_2_4=>que_out_9_2_4, 
      q_2_3=>que_out_9_2_3, q_2_2=>que_out_9_2_2, q_2_1=>que_out_9_2_1, 
      q_2_0=>que_out_9_2_0, q_3_15=>que_out_9_3_15, q_3_14=>que_out_9_3_14, 
      q_3_13=>que_out_9_3_13, q_3_12=>que_out_9_3_12, q_3_11=>que_out_9_3_11, 
      q_3_10=>que_out_9_3_10, q_3_9=>que_out_9_3_9, q_3_8=>que_out_9_3_8, 
      q_3_7=>que_out_9_3_7, q_3_6=>que_out_9_3_6, q_3_5=>que_out_9_3_5, 
      q_3_4=>que_out_9_3_4, q_3_3=>que_out_9_3_3, q_3_2=>que_out_9_3_2, 
      q_3_1=>que_out_9_3_1, q_3_0=>que_out_9_3_0, q_4_15=>que_out_9_4_15, 
      q_4_14=>que_out_9_4_14, q_4_13=>que_out_9_4_13, q_4_12=>que_out_9_4_12, 
      q_4_11=>que_out_9_4_11, q_4_10=>que_out_9_4_10, q_4_9=>que_out_9_4_9, 
      q_4_8=>que_out_9_4_8, q_4_7=>que_out_9_4_7, q_4_6=>que_out_9_4_6, 
      q_4_5=>que_out_9_4_5, q_4_4=>que_out_9_4_4, q_4_3=>que_out_9_4_3, 
      q_4_2=>que_out_9_4_2, q_4_1=>que_out_9_4_1, q_4_0=>que_out_9_4_0, clk
      =>nx10720, load=>sel_que_9, reset=>nx10696);
   gen_queues_10_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_10_0_15, q_0_14=>que_out_10_0_14, q_0_13=>
      que_out_10_0_13, q_0_12=>que_out_10_0_12, q_0_11=>que_out_10_0_11, 
      q_0_10=>que_out_10_0_10, q_0_9=>que_out_10_0_9, q_0_8=>que_out_10_0_8, 
      q_0_7=>que_out_10_0_7, q_0_6=>que_out_10_0_6, q_0_5=>que_out_10_0_5, 
      q_0_4=>que_out_10_0_4, q_0_3=>que_out_10_0_3, q_0_2=>que_out_10_0_2, 
      q_0_1=>que_out_10_0_1, q_0_0=>que_out_10_0_0, q_1_15=>que_out_10_1_15, 
      q_1_14=>que_out_10_1_14, q_1_13=>que_out_10_1_13, q_1_12=>
      que_out_10_1_12, q_1_11=>que_out_10_1_11, q_1_10=>que_out_10_1_10, 
      q_1_9=>que_out_10_1_9, q_1_8=>que_out_10_1_8, q_1_7=>que_out_10_1_7, 
      q_1_6=>que_out_10_1_6, q_1_5=>que_out_10_1_5, q_1_4=>que_out_10_1_4, 
      q_1_3=>que_out_10_1_3, q_1_2=>que_out_10_1_2, q_1_1=>que_out_10_1_1, 
      q_1_0=>que_out_10_1_0, q_2_15=>que_out_10_2_15, q_2_14=>
      que_out_10_2_14, q_2_13=>que_out_10_2_13, q_2_12=>que_out_10_2_12, 
      q_2_11=>que_out_10_2_11, q_2_10=>que_out_10_2_10, q_2_9=>
      que_out_10_2_9, q_2_8=>que_out_10_2_8, q_2_7=>que_out_10_2_7, q_2_6=>
      que_out_10_2_6, q_2_5=>que_out_10_2_5, q_2_4=>que_out_10_2_4, q_2_3=>
      que_out_10_2_3, q_2_2=>que_out_10_2_2, q_2_1=>que_out_10_2_1, q_2_0=>
      que_out_10_2_0, q_3_15=>que_out_10_3_15, q_3_14=>que_out_10_3_14, 
      q_3_13=>que_out_10_3_13, q_3_12=>que_out_10_3_12, q_3_11=>
      que_out_10_3_11, q_3_10=>que_out_10_3_10, q_3_9=>que_out_10_3_9, q_3_8
      =>que_out_10_3_8, q_3_7=>que_out_10_3_7, q_3_6=>que_out_10_3_6, q_3_5
      =>que_out_10_3_5, q_3_4=>que_out_10_3_4, q_3_3=>que_out_10_3_3, q_3_2
      =>que_out_10_3_2, q_3_1=>que_out_10_3_1, q_3_0=>que_out_10_3_0, q_4_15
      =>que_out_10_4_15, q_4_14=>que_out_10_4_14, q_4_13=>que_out_10_4_13, 
      q_4_12=>que_out_10_4_12, q_4_11=>que_out_10_4_11, q_4_10=>
      que_out_10_4_10, q_4_9=>que_out_10_4_9, q_4_8=>que_out_10_4_8, q_4_7=>
      que_out_10_4_7, q_4_6=>que_out_10_4_6, q_4_5=>que_out_10_4_5, q_4_4=>
      que_out_10_4_4, q_4_3=>que_out_10_4_3, q_4_2=>que_out_10_4_2, q_4_1=>
      que_out_10_4_1, q_4_0=>que_out_10_4_0, clk=>nx10722, load=>sel_que_10, 
      reset=>nx10698);
   gen_queues_11_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_11_0_15, q_0_14=>que_out_11_0_14, q_0_13=>
      que_out_11_0_13, q_0_12=>que_out_11_0_12, q_0_11=>que_out_11_0_11, 
      q_0_10=>que_out_11_0_10, q_0_9=>que_out_11_0_9, q_0_8=>que_out_11_0_8, 
      q_0_7=>que_out_11_0_7, q_0_6=>que_out_11_0_6, q_0_5=>que_out_11_0_5, 
      q_0_4=>que_out_11_0_4, q_0_3=>que_out_11_0_3, q_0_2=>que_out_11_0_2, 
      q_0_1=>que_out_11_0_1, q_0_0=>que_out_11_0_0, q_1_15=>que_out_11_1_15, 
      q_1_14=>que_out_11_1_14, q_1_13=>que_out_11_1_13, q_1_12=>
      que_out_11_1_12, q_1_11=>que_out_11_1_11, q_1_10=>que_out_11_1_10, 
      q_1_9=>que_out_11_1_9, q_1_8=>que_out_11_1_8, q_1_7=>que_out_11_1_7, 
      q_1_6=>que_out_11_1_6, q_1_5=>que_out_11_1_5, q_1_4=>que_out_11_1_4, 
      q_1_3=>que_out_11_1_3, q_1_2=>que_out_11_1_2, q_1_1=>que_out_11_1_1, 
      q_1_0=>que_out_11_1_0, q_2_15=>que_out_11_2_15, q_2_14=>
      que_out_11_2_14, q_2_13=>que_out_11_2_13, q_2_12=>que_out_11_2_12, 
      q_2_11=>que_out_11_2_11, q_2_10=>que_out_11_2_10, q_2_9=>
      que_out_11_2_9, q_2_8=>que_out_11_2_8, q_2_7=>que_out_11_2_7, q_2_6=>
      que_out_11_2_6, q_2_5=>que_out_11_2_5, q_2_4=>que_out_11_2_4, q_2_3=>
      que_out_11_2_3, q_2_2=>que_out_11_2_2, q_2_1=>que_out_11_2_1, q_2_0=>
      que_out_11_2_0, q_3_15=>que_out_11_3_15, q_3_14=>que_out_11_3_14, 
      q_3_13=>que_out_11_3_13, q_3_12=>que_out_11_3_12, q_3_11=>
      que_out_11_3_11, q_3_10=>que_out_11_3_10, q_3_9=>que_out_11_3_9, q_3_8
      =>que_out_11_3_8, q_3_7=>que_out_11_3_7, q_3_6=>que_out_11_3_6, q_3_5
      =>que_out_11_3_5, q_3_4=>que_out_11_3_4, q_3_3=>que_out_11_3_3, q_3_2
      =>que_out_11_3_2, q_3_1=>que_out_11_3_1, q_3_0=>que_out_11_3_0, q_4_15
      =>que_out_11_4_15, q_4_14=>que_out_11_4_14, q_4_13=>que_out_11_4_13, 
      q_4_12=>que_out_11_4_12, q_4_11=>que_out_11_4_11, q_4_10=>
      que_out_11_4_10, q_4_9=>que_out_11_4_9, q_4_8=>que_out_11_4_8, q_4_7=>
      que_out_11_4_7, q_4_6=>que_out_11_4_6, q_4_5=>que_out_11_4_5, q_4_4=>
      que_out_11_4_4, q_4_3=>que_out_11_4_3, q_4_2=>que_out_11_4_2, q_4_1=>
      que_out_11_4_1, q_4_0=>que_out_11_4_0, clk=>nx10722, load=>sel_que_11, 
      reset=>nx10698);
   gen_queues_12_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_12_0_15, q_0_14=>que_out_12_0_14, q_0_13=>
      que_out_12_0_13, q_0_12=>que_out_12_0_12, q_0_11=>que_out_12_0_11, 
      q_0_10=>que_out_12_0_10, q_0_9=>que_out_12_0_9, q_0_8=>que_out_12_0_8, 
      q_0_7=>que_out_12_0_7, q_0_6=>que_out_12_0_6, q_0_5=>que_out_12_0_5, 
      q_0_4=>que_out_12_0_4, q_0_3=>que_out_12_0_3, q_0_2=>que_out_12_0_2, 
      q_0_1=>que_out_12_0_1, q_0_0=>que_out_12_0_0, q_1_15=>que_out_12_1_15, 
      q_1_14=>que_out_12_1_14, q_1_13=>que_out_12_1_13, q_1_12=>
      que_out_12_1_12, q_1_11=>que_out_12_1_11, q_1_10=>que_out_12_1_10, 
      q_1_9=>que_out_12_1_9, q_1_8=>que_out_12_1_8, q_1_7=>que_out_12_1_7, 
      q_1_6=>que_out_12_1_6, q_1_5=>que_out_12_1_5, q_1_4=>que_out_12_1_4, 
      q_1_3=>que_out_12_1_3, q_1_2=>que_out_12_1_2, q_1_1=>que_out_12_1_1, 
      q_1_0=>que_out_12_1_0, q_2_15=>que_out_12_2_15, q_2_14=>
      que_out_12_2_14, q_2_13=>que_out_12_2_13, q_2_12=>que_out_12_2_12, 
      q_2_11=>que_out_12_2_11, q_2_10=>que_out_12_2_10, q_2_9=>
      que_out_12_2_9, q_2_8=>que_out_12_2_8, q_2_7=>que_out_12_2_7, q_2_6=>
      que_out_12_2_6, q_2_5=>que_out_12_2_5, q_2_4=>que_out_12_2_4, q_2_3=>
      que_out_12_2_3, q_2_2=>que_out_12_2_2, q_2_1=>que_out_12_2_1, q_2_0=>
      que_out_12_2_0, q_3_15=>que_out_12_3_15, q_3_14=>que_out_12_3_14, 
      q_3_13=>que_out_12_3_13, q_3_12=>que_out_12_3_12, q_3_11=>
      que_out_12_3_11, q_3_10=>que_out_12_3_10, q_3_9=>que_out_12_3_9, q_3_8
      =>que_out_12_3_8, q_3_7=>que_out_12_3_7, q_3_6=>que_out_12_3_6, q_3_5
      =>que_out_12_3_5, q_3_4=>que_out_12_3_4, q_3_3=>que_out_12_3_3, q_3_2
      =>que_out_12_3_2, q_3_1=>que_out_12_3_1, q_3_0=>que_out_12_3_0, q_4_15
      =>que_out_12_4_15, q_4_14=>que_out_12_4_14, q_4_13=>que_out_12_4_13, 
      q_4_12=>que_out_12_4_12, q_4_11=>que_out_12_4_11, q_4_10=>
      que_out_12_4_10, q_4_9=>que_out_12_4_9, q_4_8=>que_out_12_4_8, q_4_7=>
      que_out_12_4_7, q_4_6=>que_out_12_4_6, q_4_5=>que_out_12_4_5, q_4_4=>
      que_out_12_4_4, q_4_3=>que_out_12_4_3, q_4_2=>que_out_12_4_2, q_4_1=>
      que_out_12_4_1, q_4_0=>que_out_12_4_0, clk=>nx10722, load=>sel_que_12, 
      reset=>nx10698);
   gen_queues_13_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_13_0_15, q_0_14=>que_out_13_0_14, q_0_13=>
      que_out_13_0_13, q_0_12=>que_out_13_0_12, q_0_11=>que_out_13_0_11, 
      q_0_10=>que_out_13_0_10, q_0_9=>que_out_13_0_9, q_0_8=>que_out_13_0_8, 
      q_0_7=>que_out_13_0_7, q_0_6=>que_out_13_0_6, q_0_5=>que_out_13_0_5, 
      q_0_4=>que_out_13_0_4, q_0_3=>que_out_13_0_3, q_0_2=>que_out_13_0_2, 
      q_0_1=>que_out_13_0_1, q_0_0=>que_out_13_0_0, q_1_15=>que_out_13_1_15, 
      q_1_14=>que_out_13_1_14, q_1_13=>que_out_13_1_13, q_1_12=>
      que_out_13_1_12, q_1_11=>que_out_13_1_11, q_1_10=>que_out_13_1_10, 
      q_1_9=>que_out_13_1_9, q_1_8=>que_out_13_1_8, q_1_7=>que_out_13_1_7, 
      q_1_6=>que_out_13_1_6, q_1_5=>que_out_13_1_5, q_1_4=>que_out_13_1_4, 
      q_1_3=>que_out_13_1_3, q_1_2=>que_out_13_1_2, q_1_1=>que_out_13_1_1, 
      q_1_0=>que_out_13_1_0, q_2_15=>que_out_13_2_15, q_2_14=>
      que_out_13_2_14, q_2_13=>que_out_13_2_13, q_2_12=>que_out_13_2_12, 
      q_2_11=>que_out_13_2_11, q_2_10=>que_out_13_2_10, q_2_9=>
      que_out_13_2_9, q_2_8=>que_out_13_2_8, q_2_7=>que_out_13_2_7, q_2_6=>
      que_out_13_2_6, q_2_5=>que_out_13_2_5, q_2_4=>que_out_13_2_4, q_2_3=>
      que_out_13_2_3, q_2_2=>que_out_13_2_2, q_2_1=>que_out_13_2_1, q_2_0=>
      que_out_13_2_0, q_3_15=>que_out_13_3_15, q_3_14=>que_out_13_3_14, 
      q_3_13=>que_out_13_3_13, q_3_12=>que_out_13_3_12, q_3_11=>
      que_out_13_3_11, q_3_10=>que_out_13_3_10, q_3_9=>que_out_13_3_9, q_3_8
      =>que_out_13_3_8, q_3_7=>que_out_13_3_7, q_3_6=>que_out_13_3_6, q_3_5
      =>que_out_13_3_5, q_3_4=>que_out_13_3_4, q_3_3=>que_out_13_3_3, q_3_2
      =>que_out_13_3_2, q_3_1=>que_out_13_3_1, q_3_0=>que_out_13_3_0, q_4_15
      =>que_out_13_4_15, q_4_14=>que_out_13_4_14, q_4_13=>que_out_13_4_13, 
      q_4_12=>que_out_13_4_12, q_4_11=>que_out_13_4_11, q_4_10=>
      que_out_13_4_10, q_4_9=>que_out_13_4_9, q_4_8=>que_out_13_4_8, q_4_7=>
      que_out_13_4_7, q_4_6=>que_out_13_4_6, q_4_5=>que_out_13_4_5, q_4_4=>
      que_out_13_4_4, q_4_3=>que_out_13_4_3, q_4_2=>que_out_13_4_2, q_4_1=>
      que_out_13_4_1, q_4_0=>que_out_13_4_0, clk=>nx10724, load=>sel_que_13, 
      reset=>nx10700);
   gen_queues_14_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_14_0_15, q_0_14=>que_out_14_0_14, q_0_13=>
      que_out_14_0_13, q_0_12=>que_out_14_0_12, q_0_11=>que_out_14_0_11, 
      q_0_10=>que_out_14_0_10, q_0_9=>que_out_14_0_9, q_0_8=>que_out_14_0_8, 
      q_0_7=>que_out_14_0_7, q_0_6=>que_out_14_0_6, q_0_5=>que_out_14_0_5, 
      q_0_4=>que_out_14_0_4, q_0_3=>que_out_14_0_3, q_0_2=>que_out_14_0_2, 
      q_0_1=>que_out_14_0_1, q_0_0=>que_out_14_0_0, q_1_15=>que_out_14_1_15, 
      q_1_14=>que_out_14_1_14, q_1_13=>que_out_14_1_13, q_1_12=>
      que_out_14_1_12, q_1_11=>que_out_14_1_11, q_1_10=>que_out_14_1_10, 
      q_1_9=>que_out_14_1_9, q_1_8=>que_out_14_1_8, q_1_7=>que_out_14_1_7, 
      q_1_6=>que_out_14_1_6, q_1_5=>que_out_14_1_5, q_1_4=>que_out_14_1_4, 
      q_1_3=>que_out_14_1_3, q_1_2=>que_out_14_1_2, q_1_1=>que_out_14_1_1, 
      q_1_0=>que_out_14_1_0, q_2_15=>que_out_14_2_15, q_2_14=>
      que_out_14_2_14, q_2_13=>que_out_14_2_13, q_2_12=>que_out_14_2_12, 
      q_2_11=>que_out_14_2_11, q_2_10=>que_out_14_2_10, q_2_9=>
      que_out_14_2_9, q_2_8=>que_out_14_2_8, q_2_7=>que_out_14_2_7, q_2_6=>
      que_out_14_2_6, q_2_5=>que_out_14_2_5, q_2_4=>que_out_14_2_4, q_2_3=>
      que_out_14_2_3, q_2_2=>que_out_14_2_2, q_2_1=>que_out_14_2_1, q_2_0=>
      que_out_14_2_0, q_3_15=>que_out_14_3_15, q_3_14=>que_out_14_3_14, 
      q_3_13=>que_out_14_3_13, q_3_12=>que_out_14_3_12, q_3_11=>
      que_out_14_3_11, q_3_10=>que_out_14_3_10, q_3_9=>que_out_14_3_9, q_3_8
      =>que_out_14_3_8, q_3_7=>que_out_14_3_7, q_3_6=>que_out_14_3_6, q_3_5
      =>que_out_14_3_5, q_3_4=>que_out_14_3_4, q_3_3=>que_out_14_3_3, q_3_2
      =>que_out_14_3_2, q_3_1=>que_out_14_3_1, q_3_0=>que_out_14_3_0, q_4_15
      =>que_out_14_4_15, q_4_14=>que_out_14_4_14, q_4_13=>que_out_14_4_13, 
      q_4_12=>que_out_14_4_12, q_4_11=>que_out_14_4_11, q_4_10=>
      que_out_14_4_10, q_4_9=>que_out_14_4_9, q_4_8=>que_out_14_4_8, q_4_7=>
      que_out_14_4_7, q_4_6=>que_out_14_4_6, q_4_5=>que_out_14_4_5, q_4_4=>
      que_out_14_4_4, q_4_3=>que_out_14_4_3, q_4_2=>que_out_14_4_2, q_4_1=>
      que_out_14_4_1, q_4_0=>que_out_14_4_0, clk=>nx10726, load=>sel_que_14, 
      reset=>nx10702);
   gen_queues_15_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_15_0_15, q_0_14=>que_out_15_0_14, q_0_13=>
      que_out_15_0_13, q_0_12=>que_out_15_0_12, q_0_11=>que_out_15_0_11, 
      q_0_10=>que_out_15_0_10, q_0_9=>que_out_15_0_9, q_0_8=>que_out_15_0_8, 
      q_0_7=>que_out_15_0_7, q_0_6=>que_out_15_0_6, q_0_5=>que_out_15_0_5, 
      q_0_4=>que_out_15_0_4, q_0_3=>que_out_15_0_3, q_0_2=>que_out_15_0_2, 
      q_0_1=>que_out_15_0_1, q_0_0=>que_out_15_0_0, q_1_15=>que_out_15_1_15, 
      q_1_14=>que_out_15_1_14, q_1_13=>que_out_15_1_13, q_1_12=>
      que_out_15_1_12, q_1_11=>que_out_15_1_11, q_1_10=>que_out_15_1_10, 
      q_1_9=>que_out_15_1_9, q_1_8=>que_out_15_1_8, q_1_7=>que_out_15_1_7, 
      q_1_6=>que_out_15_1_6, q_1_5=>que_out_15_1_5, q_1_4=>que_out_15_1_4, 
      q_1_3=>que_out_15_1_3, q_1_2=>que_out_15_1_2, q_1_1=>que_out_15_1_1, 
      q_1_0=>que_out_15_1_0, q_2_15=>que_out_15_2_15, q_2_14=>
      que_out_15_2_14, q_2_13=>que_out_15_2_13, q_2_12=>que_out_15_2_12, 
      q_2_11=>que_out_15_2_11, q_2_10=>que_out_15_2_10, q_2_9=>
      que_out_15_2_9, q_2_8=>que_out_15_2_8, q_2_7=>que_out_15_2_7, q_2_6=>
      que_out_15_2_6, q_2_5=>que_out_15_2_5, q_2_4=>que_out_15_2_4, q_2_3=>
      que_out_15_2_3, q_2_2=>que_out_15_2_2, q_2_1=>que_out_15_2_1, q_2_0=>
      que_out_15_2_0, q_3_15=>que_out_15_3_15, q_3_14=>que_out_15_3_14, 
      q_3_13=>que_out_15_3_13, q_3_12=>que_out_15_3_12, q_3_11=>
      que_out_15_3_11, q_3_10=>que_out_15_3_10, q_3_9=>que_out_15_3_9, q_3_8
      =>que_out_15_3_8, q_3_7=>que_out_15_3_7, q_3_6=>que_out_15_3_6, q_3_5
      =>que_out_15_3_5, q_3_4=>que_out_15_3_4, q_3_3=>que_out_15_3_3, q_3_2
      =>que_out_15_3_2, q_3_1=>que_out_15_3_1, q_3_0=>que_out_15_3_0, q_4_15
      =>que_out_15_4_15, q_4_14=>que_out_15_4_14, q_4_13=>que_out_15_4_13, 
      q_4_12=>que_out_15_4_12, q_4_11=>que_out_15_4_11, q_4_10=>
      que_out_15_4_10, q_4_9=>que_out_15_4_9, q_4_8=>que_out_15_4_8, q_4_7=>
      que_out_15_4_7, q_4_6=>que_out_15_4_6, q_4_5=>que_out_15_4_5, q_4_4=>
      que_out_15_4_4, q_4_3=>que_out_15_4_3, q_4_2=>que_out_15_4_2, q_4_1=>
      que_out_15_4_1, q_4_0=>que_out_15_4_0, clk=>nx10726, load=>sel_que_15, 
      reset=>nx10702);
   gen_queues_16_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_16_0_15, q_0_14=>que_out_16_0_14, q_0_13=>
      que_out_16_0_13, q_0_12=>que_out_16_0_12, q_0_11=>que_out_16_0_11, 
      q_0_10=>que_out_16_0_10, q_0_9=>que_out_16_0_9, q_0_8=>que_out_16_0_8, 
      q_0_7=>que_out_16_0_7, q_0_6=>que_out_16_0_6, q_0_5=>que_out_16_0_5, 
      q_0_4=>que_out_16_0_4, q_0_3=>que_out_16_0_3, q_0_2=>que_out_16_0_2, 
      q_0_1=>que_out_16_0_1, q_0_0=>que_out_16_0_0, q_1_15=>que_out_16_1_15, 
      q_1_14=>que_out_16_1_14, q_1_13=>que_out_16_1_13, q_1_12=>
      que_out_16_1_12, q_1_11=>que_out_16_1_11, q_1_10=>que_out_16_1_10, 
      q_1_9=>que_out_16_1_9, q_1_8=>que_out_16_1_8, q_1_7=>que_out_16_1_7, 
      q_1_6=>que_out_16_1_6, q_1_5=>que_out_16_1_5, q_1_4=>que_out_16_1_4, 
      q_1_3=>que_out_16_1_3, q_1_2=>que_out_16_1_2, q_1_1=>que_out_16_1_1, 
      q_1_0=>que_out_16_1_0, q_2_15=>que_out_16_2_15, q_2_14=>
      que_out_16_2_14, q_2_13=>que_out_16_2_13, q_2_12=>que_out_16_2_12, 
      q_2_11=>que_out_16_2_11, q_2_10=>que_out_16_2_10, q_2_9=>
      que_out_16_2_9, q_2_8=>que_out_16_2_8, q_2_7=>que_out_16_2_7, q_2_6=>
      que_out_16_2_6, q_2_5=>que_out_16_2_5, q_2_4=>que_out_16_2_4, q_2_3=>
      que_out_16_2_3, q_2_2=>que_out_16_2_2, q_2_1=>que_out_16_2_1, q_2_0=>
      que_out_16_2_0, q_3_15=>que_out_16_3_15, q_3_14=>que_out_16_3_14, 
      q_3_13=>que_out_16_3_13, q_3_12=>que_out_16_3_12, q_3_11=>
      que_out_16_3_11, q_3_10=>que_out_16_3_10, q_3_9=>que_out_16_3_9, q_3_8
      =>que_out_16_3_8, q_3_7=>que_out_16_3_7, q_3_6=>que_out_16_3_6, q_3_5
      =>que_out_16_3_5, q_3_4=>que_out_16_3_4, q_3_3=>que_out_16_3_3, q_3_2
      =>que_out_16_3_2, q_3_1=>que_out_16_3_1, q_3_0=>que_out_16_3_0, q_4_15
      =>que_out_16_4_15, q_4_14=>que_out_16_4_14, q_4_13=>que_out_16_4_13, 
      q_4_12=>que_out_16_4_12, q_4_11=>que_out_16_4_11, q_4_10=>
      que_out_16_4_10, q_4_9=>que_out_16_4_9, q_4_8=>que_out_16_4_8, q_4_7=>
      que_out_16_4_7, q_4_6=>que_out_16_4_6, q_4_5=>que_out_16_4_5, q_4_4=>
      que_out_16_4_4, q_4_3=>que_out_16_4_3, q_4_2=>que_out_16_4_2, q_4_1=>
      que_out_16_4_1, q_4_0=>que_out_16_4_0, clk=>nx10726, load=>sel_que_16, 
      reset=>nx10702);
   gen_queues_17_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_17_0_15, q_0_14=>que_out_17_0_14, q_0_13=>
      que_out_17_0_13, q_0_12=>que_out_17_0_12, q_0_11=>que_out_17_0_11, 
      q_0_10=>que_out_17_0_10, q_0_9=>que_out_17_0_9, q_0_8=>que_out_17_0_8, 
      q_0_7=>que_out_17_0_7, q_0_6=>que_out_17_0_6, q_0_5=>que_out_17_0_5, 
      q_0_4=>que_out_17_0_4, q_0_3=>que_out_17_0_3, q_0_2=>que_out_17_0_2, 
      q_0_1=>que_out_17_0_1, q_0_0=>que_out_17_0_0, q_1_15=>que_out_17_1_15, 
      q_1_14=>que_out_17_1_14, q_1_13=>que_out_17_1_13, q_1_12=>
      que_out_17_1_12, q_1_11=>que_out_17_1_11, q_1_10=>que_out_17_1_10, 
      q_1_9=>que_out_17_1_9, q_1_8=>que_out_17_1_8, q_1_7=>que_out_17_1_7, 
      q_1_6=>que_out_17_1_6, q_1_5=>que_out_17_1_5, q_1_4=>que_out_17_1_4, 
      q_1_3=>que_out_17_1_3, q_1_2=>que_out_17_1_2, q_1_1=>que_out_17_1_1, 
      q_1_0=>que_out_17_1_0, q_2_15=>que_out_17_2_15, q_2_14=>
      que_out_17_2_14, q_2_13=>que_out_17_2_13, q_2_12=>que_out_17_2_12, 
      q_2_11=>que_out_17_2_11, q_2_10=>que_out_17_2_10, q_2_9=>
      que_out_17_2_9, q_2_8=>que_out_17_2_8, q_2_7=>que_out_17_2_7, q_2_6=>
      que_out_17_2_6, q_2_5=>que_out_17_2_5, q_2_4=>que_out_17_2_4, q_2_3=>
      que_out_17_2_3, q_2_2=>que_out_17_2_2, q_2_1=>que_out_17_2_1, q_2_0=>
      que_out_17_2_0, q_3_15=>que_out_17_3_15, q_3_14=>que_out_17_3_14, 
      q_3_13=>que_out_17_3_13, q_3_12=>que_out_17_3_12, q_3_11=>
      que_out_17_3_11, q_3_10=>que_out_17_3_10, q_3_9=>que_out_17_3_9, q_3_8
      =>que_out_17_3_8, q_3_7=>que_out_17_3_7, q_3_6=>que_out_17_3_6, q_3_5
      =>que_out_17_3_5, q_3_4=>que_out_17_3_4, q_3_3=>que_out_17_3_3, q_3_2
      =>que_out_17_3_2, q_3_1=>que_out_17_3_1, q_3_0=>que_out_17_3_0, q_4_15
      =>que_out_17_4_15, q_4_14=>que_out_17_4_14, q_4_13=>que_out_17_4_13, 
      q_4_12=>que_out_17_4_12, q_4_11=>que_out_17_4_11, q_4_10=>
      que_out_17_4_10, q_4_9=>que_out_17_4_9, q_4_8=>que_out_17_4_8, q_4_7=>
      que_out_17_4_7, q_4_6=>que_out_17_4_6, q_4_5=>que_out_17_4_5, q_4_4=>
      que_out_17_4_4, q_4_3=>que_out_17_4_3, q_4_2=>que_out_17_4_2, q_4_1=>
      que_out_17_4_1, q_4_0=>que_out_17_4_0, clk=>nx10728, load=>sel_que_17, 
      reset=>nx10704);
   gen_queues_18_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_18_0_15, q_0_14=>que_out_18_0_14, q_0_13=>
      que_out_18_0_13, q_0_12=>que_out_18_0_12, q_0_11=>que_out_18_0_11, 
      q_0_10=>que_out_18_0_10, q_0_9=>que_out_18_0_9, q_0_8=>que_out_18_0_8, 
      q_0_7=>que_out_18_0_7, q_0_6=>que_out_18_0_6, q_0_5=>que_out_18_0_5, 
      q_0_4=>que_out_18_0_4, q_0_3=>que_out_18_0_3, q_0_2=>que_out_18_0_2, 
      q_0_1=>que_out_18_0_1, q_0_0=>que_out_18_0_0, q_1_15=>que_out_18_1_15, 
      q_1_14=>que_out_18_1_14, q_1_13=>que_out_18_1_13, q_1_12=>
      que_out_18_1_12, q_1_11=>que_out_18_1_11, q_1_10=>que_out_18_1_10, 
      q_1_9=>que_out_18_1_9, q_1_8=>que_out_18_1_8, q_1_7=>que_out_18_1_7, 
      q_1_6=>que_out_18_1_6, q_1_5=>que_out_18_1_5, q_1_4=>que_out_18_1_4, 
      q_1_3=>que_out_18_1_3, q_1_2=>que_out_18_1_2, q_1_1=>que_out_18_1_1, 
      q_1_0=>que_out_18_1_0, q_2_15=>que_out_18_2_15, q_2_14=>
      que_out_18_2_14, q_2_13=>que_out_18_2_13, q_2_12=>que_out_18_2_12, 
      q_2_11=>que_out_18_2_11, q_2_10=>que_out_18_2_10, q_2_9=>
      que_out_18_2_9, q_2_8=>que_out_18_2_8, q_2_7=>que_out_18_2_7, q_2_6=>
      que_out_18_2_6, q_2_5=>que_out_18_2_5, q_2_4=>que_out_18_2_4, q_2_3=>
      que_out_18_2_3, q_2_2=>que_out_18_2_2, q_2_1=>que_out_18_2_1, q_2_0=>
      que_out_18_2_0, q_3_15=>que_out_18_3_15, q_3_14=>que_out_18_3_14, 
      q_3_13=>que_out_18_3_13, q_3_12=>que_out_18_3_12, q_3_11=>
      que_out_18_3_11, q_3_10=>que_out_18_3_10, q_3_9=>que_out_18_3_9, q_3_8
      =>que_out_18_3_8, q_3_7=>que_out_18_3_7, q_3_6=>que_out_18_3_6, q_3_5
      =>que_out_18_3_5, q_3_4=>que_out_18_3_4, q_3_3=>que_out_18_3_3, q_3_2
      =>que_out_18_3_2, q_3_1=>que_out_18_3_1, q_3_0=>que_out_18_3_0, q_4_15
      =>que_out_18_4_15, q_4_14=>que_out_18_4_14, q_4_13=>que_out_18_4_13, 
      q_4_12=>que_out_18_4_12, q_4_11=>que_out_18_4_11, q_4_10=>
      que_out_18_4_10, q_4_9=>que_out_18_4_9, q_4_8=>que_out_18_4_8, q_4_7=>
      que_out_18_4_7, q_4_6=>que_out_18_4_6, q_4_5=>que_out_18_4_5, q_4_4=>
      que_out_18_4_4, q_4_3=>que_out_18_4_3, q_4_2=>que_out_18_4_2, q_4_1=>
      que_out_18_4_1, q_4_0=>que_out_18_4_0, clk=>nx10728, load=>sel_que_18, 
      reset=>nx10704);
   gen_queues_19_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_19_0_15, q_0_14=>que_out_19_0_14, q_0_13=>
      que_out_19_0_13, q_0_12=>que_out_19_0_12, q_0_11=>que_out_19_0_11, 
      q_0_10=>que_out_19_0_10, q_0_9=>que_out_19_0_9, q_0_8=>que_out_19_0_8, 
      q_0_7=>que_out_19_0_7, q_0_6=>que_out_19_0_6, q_0_5=>que_out_19_0_5, 
      q_0_4=>que_out_19_0_4, q_0_3=>que_out_19_0_3, q_0_2=>que_out_19_0_2, 
      q_0_1=>que_out_19_0_1, q_0_0=>que_out_19_0_0, q_1_15=>que_out_19_1_15, 
      q_1_14=>que_out_19_1_14, q_1_13=>que_out_19_1_13, q_1_12=>
      que_out_19_1_12, q_1_11=>que_out_19_1_11, q_1_10=>que_out_19_1_10, 
      q_1_9=>que_out_19_1_9, q_1_8=>que_out_19_1_8, q_1_7=>que_out_19_1_7, 
      q_1_6=>que_out_19_1_6, q_1_5=>que_out_19_1_5, q_1_4=>que_out_19_1_4, 
      q_1_3=>que_out_19_1_3, q_1_2=>que_out_19_1_2, q_1_1=>que_out_19_1_1, 
      q_1_0=>que_out_19_1_0, q_2_15=>que_out_19_2_15, q_2_14=>
      que_out_19_2_14, q_2_13=>que_out_19_2_13, q_2_12=>que_out_19_2_12, 
      q_2_11=>que_out_19_2_11, q_2_10=>que_out_19_2_10, q_2_9=>
      que_out_19_2_9, q_2_8=>que_out_19_2_8, q_2_7=>que_out_19_2_7, q_2_6=>
      que_out_19_2_6, q_2_5=>que_out_19_2_5, q_2_4=>que_out_19_2_4, q_2_3=>
      que_out_19_2_3, q_2_2=>que_out_19_2_2, q_2_1=>que_out_19_2_1, q_2_0=>
      que_out_19_2_0, q_3_15=>que_out_19_3_15, q_3_14=>que_out_19_3_14, 
      q_3_13=>que_out_19_3_13, q_3_12=>que_out_19_3_12, q_3_11=>
      que_out_19_3_11, q_3_10=>que_out_19_3_10, q_3_9=>que_out_19_3_9, q_3_8
      =>que_out_19_3_8, q_3_7=>que_out_19_3_7, q_3_6=>que_out_19_3_6, q_3_5
      =>que_out_19_3_5, q_3_4=>que_out_19_3_4, q_3_3=>que_out_19_3_3, q_3_2
      =>que_out_19_3_2, q_3_1=>que_out_19_3_1, q_3_0=>que_out_19_3_0, q_4_15
      =>que_out_19_4_15, q_4_14=>que_out_19_4_14, q_4_13=>que_out_19_4_13, 
      q_4_12=>que_out_19_4_12, q_4_11=>que_out_19_4_11, q_4_10=>
      que_out_19_4_10, q_4_9=>que_out_19_4_9, q_4_8=>que_out_19_4_8, q_4_7=>
      que_out_19_4_7, q_4_6=>que_out_19_4_6, q_4_5=>que_out_19_4_5, q_4_4=>
      que_out_19_4_4, q_4_3=>que_out_19_4_3, q_4_2=>que_out_19_4_2, q_4_1=>
      que_out_19_4_1, q_4_0=>que_out_19_4_0, clk=>nx10728, load=>sel_que_19, 
      reset=>nx10704);
   gen_queues_20_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_20_0_15, q_0_14=>que_out_20_0_14, q_0_13=>
      que_out_20_0_13, q_0_12=>que_out_20_0_12, q_0_11=>que_out_20_0_11, 
      q_0_10=>que_out_20_0_10, q_0_9=>que_out_20_0_9, q_0_8=>que_out_20_0_8, 
      q_0_7=>que_out_20_0_7, q_0_6=>que_out_20_0_6, q_0_5=>que_out_20_0_5, 
      q_0_4=>que_out_20_0_4, q_0_3=>que_out_20_0_3, q_0_2=>que_out_20_0_2, 
      q_0_1=>que_out_20_0_1, q_0_0=>que_out_20_0_0, q_1_15=>que_out_20_1_15, 
      q_1_14=>que_out_20_1_14, q_1_13=>que_out_20_1_13, q_1_12=>
      que_out_20_1_12, q_1_11=>que_out_20_1_11, q_1_10=>que_out_20_1_10, 
      q_1_9=>que_out_20_1_9, q_1_8=>que_out_20_1_8, q_1_7=>que_out_20_1_7, 
      q_1_6=>que_out_20_1_6, q_1_5=>que_out_20_1_5, q_1_4=>que_out_20_1_4, 
      q_1_3=>que_out_20_1_3, q_1_2=>que_out_20_1_2, q_1_1=>que_out_20_1_1, 
      q_1_0=>que_out_20_1_0, q_2_15=>que_out_20_2_15, q_2_14=>
      que_out_20_2_14, q_2_13=>que_out_20_2_13, q_2_12=>que_out_20_2_12, 
      q_2_11=>que_out_20_2_11, q_2_10=>que_out_20_2_10, q_2_9=>
      que_out_20_2_9, q_2_8=>que_out_20_2_8, q_2_7=>que_out_20_2_7, q_2_6=>
      que_out_20_2_6, q_2_5=>que_out_20_2_5, q_2_4=>que_out_20_2_4, q_2_3=>
      que_out_20_2_3, q_2_2=>que_out_20_2_2, q_2_1=>que_out_20_2_1, q_2_0=>
      que_out_20_2_0, q_3_15=>que_out_20_3_15, q_3_14=>que_out_20_3_14, 
      q_3_13=>que_out_20_3_13, q_3_12=>que_out_20_3_12, q_3_11=>
      que_out_20_3_11, q_3_10=>que_out_20_3_10, q_3_9=>que_out_20_3_9, q_3_8
      =>que_out_20_3_8, q_3_7=>que_out_20_3_7, q_3_6=>que_out_20_3_6, q_3_5
      =>que_out_20_3_5, q_3_4=>que_out_20_3_4, q_3_3=>que_out_20_3_3, q_3_2
      =>que_out_20_3_2, q_3_1=>que_out_20_3_1, q_3_0=>que_out_20_3_0, q_4_15
      =>que_out_20_4_15, q_4_14=>que_out_20_4_14, q_4_13=>que_out_20_4_13, 
      q_4_12=>que_out_20_4_12, q_4_11=>que_out_20_4_11, q_4_10=>
      que_out_20_4_10, q_4_9=>que_out_20_4_9, q_4_8=>que_out_20_4_8, q_4_7=>
      que_out_20_4_7, q_4_6=>que_out_20_4_6, q_4_5=>que_out_20_4_5, q_4_4=>
      que_out_20_4_4, q_4_3=>que_out_20_4_3, q_4_2=>que_out_20_4_2, q_4_1=>
      que_out_20_4_1, q_4_0=>que_out_20_4_0, clk=>nx10730, load=>sel_que_20, 
      reset=>nx10706);
   gen_queues_21_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_21_0_15, q_0_14=>que_out_21_0_14, q_0_13=>
      que_out_21_0_13, q_0_12=>que_out_21_0_12, q_0_11=>que_out_21_0_11, 
      q_0_10=>que_out_21_0_10, q_0_9=>que_out_21_0_9, q_0_8=>que_out_21_0_8, 
      q_0_7=>que_out_21_0_7, q_0_6=>que_out_21_0_6, q_0_5=>que_out_21_0_5, 
      q_0_4=>que_out_21_0_4, q_0_3=>que_out_21_0_3, q_0_2=>que_out_21_0_2, 
      q_0_1=>que_out_21_0_1, q_0_0=>que_out_21_0_0, q_1_15=>que_out_21_1_15, 
      q_1_14=>que_out_21_1_14, q_1_13=>que_out_21_1_13, q_1_12=>
      que_out_21_1_12, q_1_11=>que_out_21_1_11, q_1_10=>que_out_21_1_10, 
      q_1_9=>que_out_21_1_9, q_1_8=>que_out_21_1_8, q_1_7=>que_out_21_1_7, 
      q_1_6=>que_out_21_1_6, q_1_5=>que_out_21_1_5, q_1_4=>que_out_21_1_4, 
      q_1_3=>que_out_21_1_3, q_1_2=>que_out_21_1_2, q_1_1=>que_out_21_1_1, 
      q_1_0=>que_out_21_1_0, q_2_15=>que_out_21_2_15, q_2_14=>
      que_out_21_2_14, q_2_13=>que_out_21_2_13, q_2_12=>que_out_21_2_12, 
      q_2_11=>que_out_21_2_11, q_2_10=>que_out_21_2_10, q_2_9=>
      que_out_21_2_9, q_2_8=>que_out_21_2_8, q_2_7=>que_out_21_2_7, q_2_6=>
      que_out_21_2_6, q_2_5=>que_out_21_2_5, q_2_4=>que_out_21_2_4, q_2_3=>
      que_out_21_2_3, q_2_2=>que_out_21_2_2, q_2_1=>que_out_21_2_1, q_2_0=>
      que_out_21_2_0, q_3_15=>que_out_21_3_15, q_3_14=>que_out_21_3_14, 
      q_3_13=>que_out_21_3_13, q_3_12=>que_out_21_3_12, q_3_11=>
      que_out_21_3_11, q_3_10=>que_out_21_3_10, q_3_9=>que_out_21_3_9, q_3_8
      =>que_out_21_3_8, q_3_7=>que_out_21_3_7, q_3_6=>que_out_21_3_6, q_3_5
      =>que_out_21_3_5, q_3_4=>que_out_21_3_4, q_3_3=>que_out_21_3_3, q_3_2
      =>que_out_21_3_2, q_3_1=>que_out_21_3_1, q_3_0=>que_out_21_3_0, q_4_15
      =>que_out_21_4_15, q_4_14=>que_out_21_4_14, q_4_13=>que_out_21_4_13, 
      q_4_12=>que_out_21_4_12, q_4_11=>que_out_21_4_11, q_4_10=>
      que_out_21_4_10, q_4_9=>que_out_21_4_9, q_4_8=>que_out_21_4_8, q_4_7=>
      que_out_21_4_7, q_4_6=>que_out_21_4_6, q_4_5=>que_out_21_4_5, q_4_4=>
      que_out_21_4_4, q_4_3=>que_out_21_4_3, q_4_2=>que_out_21_4_2, q_4_1=>
      que_out_21_4_1, q_4_0=>que_out_21_4_0, clk=>nx10732, load=>sel_que_21, 
      reset=>nx10708);
   gen_queues_22_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_22_0_15, q_0_14=>que_out_22_0_14, q_0_13=>
      que_out_22_0_13, q_0_12=>que_out_22_0_12, q_0_11=>que_out_22_0_11, 
      q_0_10=>que_out_22_0_10, q_0_9=>que_out_22_0_9, q_0_8=>que_out_22_0_8, 
      q_0_7=>que_out_22_0_7, q_0_6=>que_out_22_0_6, q_0_5=>que_out_22_0_5, 
      q_0_4=>que_out_22_0_4, q_0_3=>que_out_22_0_3, q_0_2=>que_out_22_0_2, 
      q_0_1=>que_out_22_0_1, q_0_0=>que_out_22_0_0, q_1_15=>que_out_22_1_15, 
      q_1_14=>que_out_22_1_14, q_1_13=>que_out_22_1_13, q_1_12=>
      que_out_22_1_12, q_1_11=>que_out_22_1_11, q_1_10=>que_out_22_1_10, 
      q_1_9=>que_out_22_1_9, q_1_8=>que_out_22_1_8, q_1_7=>que_out_22_1_7, 
      q_1_6=>que_out_22_1_6, q_1_5=>que_out_22_1_5, q_1_4=>que_out_22_1_4, 
      q_1_3=>que_out_22_1_3, q_1_2=>que_out_22_1_2, q_1_1=>que_out_22_1_1, 
      q_1_0=>que_out_22_1_0, q_2_15=>que_out_22_2_15, q_2_14=>
      que_out_22_2_14, q_2_13=>que_out_22_2_13, q_2_12=>que_out_22_2_12, 
      q_2_11=>que_out_22_2_11, q_2_10=>que_out_22_2_10, q_2_9=>
      que_out_22_2_9, q_2_8=>que_out_22_2_8, q_2_7=>que_out_22_2_7, q_2_6=>
      que_out_22_2_6, q_2_5=>que_out_22_2_5, q_2_4=>que_out_22_2_4, q_2_3=>
      que_out_22_2_3, q_2_2=>que_out_22_2_2, q_2_1=>que_out_22_2_1, q_2_0=>
      que_out_22_2_0, q_3_15=>que_out_22_3_15, q_3_14=>que_out_22_3_14, 
      q_3_13=>que_out_22_3_13, q_3_12=>que_out_22_3_12, q_3_11=>
      que_out_22_3_11, q_3_10=>que_out_22_3_10, q_3_9=>que_out_22_3_9, q_3_8
      =>que_out_22_3_8, q_3_7=>que_out_22_3_7, q_3_6=>que_out_22_3_6, q_3_5
      =>que_out_22_3_5, q_3_4=>que_out_22_3_4, q_3_3=>que_out_22_3_3, q_3_2
      =>que_out_22_3_2, q_3_1=>que_out_22_3_1, q_3_0=>que_out_22_3_0, q_4_15
      =>que_out_22_4_15, q_4_14=>que_out_22_4_14, q_4_13=>que_out_22_4_13, 
      q_4_12=>que_out_22_4_12, q_4_11=>que_out_22_4_11, q_4_10=>
      que_out_22_4_10, q_4_9=>que_out_22_4_9, q_4_8=>que_out_22_4_8, q_4_7=>
      que_out_22_4_7, q_4_6=>que_out_22_4_6, q_4_5=>que_out_22_4_5, q_4_4=>
      que_out_22_4_4, q_4_3=>que_out_22_4_3, q_4_2=>que_out_22_4_2, q_4_1=>
      que_out_22_4_1, q_4_0=>que_out_22_4_0, clk=>nx10732, load=>sel_que_22, 
      reset=>nx10708);
   gen_queues_23_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_23_0_15, q_0_14=>que_out_23_0_14, q_0_13=>
      que_out_23_0_13, q_0_12=>que_out_23_0_12, q_0_11=>que_out_23_0_11, 
      q_0_10=>que_out_23_0_10, q_0_9=>que_out_23_0_9, q_0_8=>que_out_23_0_8, 
      q_0_7=>que_out_23_0_7, q_0_6=>que_out_23_0_6, q_0_5=>que_out_23_0_5, 
      q_0_4=>que_out_23_0_4, q_0_3=>que_out_23_0_3, q_0_2=>que_out_23_0_2, 
      q_0_1=>que_out_23_0_1, q_0_0=>que_out_23_0_0, q_1_15=>que_out_23_1_15, 
      q_1_14=>que_out_23_1_14, q_1_13=>que_out_23_1_13, q_1_12=>
      que_out_23_1_12, q_1_11=>que_out_23_1_11, q_1_10=>que_out_23_1_10, 
      q_1_9=>que_out_23_1_9, q_1_8=>que_out_23_1_8, q_1_7=>que_out_23_1_7, 
      q_1_6=>que_out_23_1_6, q_1_5=>que_out_23_1_5, q_1_4=>que_out_23_1_4, 
      q_1_3=>que_out_23_1_3, q_1_2=>que_out_23_1_2, q_1_1=>que_out_23_1_1, 
      q_1_0=>que_out_23_1_0, q_2_15=>que_out_23_2_15, q_2_14=>
      que_out_23_2_14, q_2_13=>que_out_23_2_13, q_2_12=>que_out_23_2_12, 
      q_2_11=>que_out_23_2_11, q_2_10=>que_out_23_2_10, q_2_9=>
      que_out_23_2_9, q_2_8=>que_out_23_2_8, q_2_7=>que_out_23_2_7, q_2_6=>
      que_out_23_2_6, q_2_5=>que_out_23_2_5, q_2_4=>que_out_23_2_4, q_2_3=>
      que_out_23_2_3, q_2_2=>que_out_23_2_2, q_2_1=>que_out_23_2_1, q_2_0=>
      que_out_23_2_0, q_3_15=>que_out_23_3_15, q_3_14=>que_out_23_3_14, 
      q_3_13=>que_out_23_3_13, q_3_12=>que_out_23_3_12, q_3_11=>
      que_out_23_3_11, q_3_10=>que_out_23_3_10, q_3_9=>que_out_23_3_9, q_3_8
      =>que_out_23_3_8, q_3_7=>que_out_23_3_7, q_3_6=>que_out_23_3_6, q_3_5
      =>que_out_23_3_5, q_3_4=>que_out_23_3_4, q_3_3=>que_out_23_3_3, q_3_2
      =>que_out_23_3_2, q_3_1=>que_out_23_3_1, q_3_0=>que_out_23_3_0, q_4_15
      =>que_out_23_4_15, q_4_14=>que_out_23_4_14, q_4_13=>que_out_23_4_13, 
      q_4_12=>que_out_23_4_12, q_4_11=>que_out_23_4_11, q_4_10=>
      que_out_23_4_10, q_4_9=>que_out_23_4_9, q_4_8=>que_out_23_4_8, q_4_7=>
      que_out_23_4_7, q_4_6=>que_out_23_4_6, q_4_5=>que_out_23_4_5, q_4_4=>
      que_out_23_4_4, q_4_3=>que_out_23_4_3, q_4_2=>que_out_23_4_2, q_4_1=>
      que_out_23_4_1, q_4_0=>que_out_23_4_0, clk=>nx10732, load=>sel_que_23, 
      reset=>nx10708);
   gen_queues_24_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_24_0_15, q_0_14=>que_out_24_0_14, q_0_13=>
      que_out_24_0_13, q_0_12=>que_out_24_0_12, q_0_11=>que_out_24_0_11, 
      q_0_10=>que_out_24_0_10, q_0_9=>que_out_24_0_9, q_0_8=>que_out_24_0_8, 
      q_0_7=>que_out_24_0_7, q_0_6=>que_out_24_0_6, q_0_5=>que_out_24_0_5, 
      q_0_4=>que_out_24_0_4, q_0_3=>que_out_24_0_3, q_0_2=>que_out_24_0_2, 
      q_0_1=>que_out_24_0_1, q_0_0=>que_out_24_0_0, q_1_15=>que_out_24_1_15, 
      q_1_14=>que_out_24_1_14, q_1_13=>que_out_24_1_13, q_1_12=>
      que_out_24_1_12, q_1_11=>que_out_24_1_11, q_1_10=>que_out_24_1_10, 
      q_1_9=>que_out_24_1_9, q_1_8=>que_out_24_1_8, q_1_7=>que_out_24_1_7, 
      q_1_6=>que_out_24_1_6, q_1_5=>que_out_24_1_5, q_1_4=>que_out_24_1_4, 
      q_1_3=>que_out_24_1_3, q_1_2=>que_out_24_1_2, q_1_1=>que_out_24_1_1, 
      q_1_0=>que_out_24_1_0, q_2_15=>que_out_24_2_15, q_2_14=>
      que_out_24_2_14, q_2_13=>que_out_24_2_13, q_2_12=>que_out_24_2_12, 
      q_2_11=>que_out_24_2_11, q_2_10=>que_out_24_2_10, q_2_9=>
      que_out_24_2_9, q_2_8=>que_out_24_2_8, q_2_7=>que_out_24_2_7, q_2_6=>
      que_out_24_2_6, q_2_5=>que_out_24_2_5, q_2_4=>que_out_24_2_4, q_2_3=>
      que_out_24_2_3, q_2_2=>que_out_24_2_2, q_2_1=>que_out_24_2_1, q_2_0=>
      que_out_24_2_0, q_3_15=>que_out_24_3_15, q_3_14=>que_out_24_3_14, 
      q_3_13=>que_out_24_3_13, q_3_12=>que_out_24_3_12, q_3_11=>
      que_out_24_3_11, q_3_10=>que_out_24_3_10, q_3_9=>que_out_24_3_9, q_3_8
      =>que_out_24_3_8, q_3_7=>que_out_24_3_7, q_3_6=>que_out_24_3_6, q_3_5
      =>que_out_24_3_5, q_3_4=>que_out_24_3_4, q_3_3=>que_out_24_3_3, q_3_2
      =>que_out_24_3_2, q_3_1=>que_out_24_3_1, q_3_0=>que_out_24_3_0, q_4_15
      =>que_out_24_4_15, q_4_14=>que_out_24_4_14, q_4_13=>que_out_24_4_13, 
      q_4_12=>que_out_24_4_12, q_4_11=>que_out_24_4_11, q_4_10=>
      que_out_24_4_10, q_4_9=>que_out_24_4_9, q_4_8=>que_out_24_4_8, q_4_7=>
      que_out_24_4_7, q_4_6=>que_out_24_4_6, q_4_5=>que_out_24_4_5, q_4_4=>
      que_out_24_4_4, q_4_3=>que_out_24_4_3, q_4_2=>que_out_24_4_2, q_4_1=>
      que_out_24_4_1, q_4_0=>que_out_24_4_0, clk=>nx10734, load=>sel_que_24, 
      reset=>nx10710);
   gen_queues_25_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_25_0_15, q_0_14=>que_out_25_0_14, q_0_13=>
      que_out_25_0_13, q_0_12=>que_out_25_0_12, q_0_11=>que_out_25_0_11, 
      q_0_10=>que_out_25_0_10, q_0_9=>que_out_25_0_9, q_0_8=>que_out_25_0_8, 
      q_0_7=>que_out_25_0_7, q_0_6=>que_out_25_0_6, q_0_5=>que_out_25_0_5, 
      q_0_4=>que_out_25_0_4, q_0_3=>que_out_25_0_3, q_0_2=>que_out_25_0_2, 
      q_0_1=>que_out_25_0_1, q_0_0=>que_out_25_0_0, q_1_15=>que_out_25_1_15, 
      q_1_14=>que_out_25_1_14, q_1_13=>que_out_25_1_13, q_1_12=>
      que_out_25_1_12, q_1_11=>que_out_25_1_11, q_1_10=>que_out_25_1_10, 
      q_1_9=>que_out_25_1_9, q_1_8=>que_out_25_1_8, q_1_7=>que_out_25_1_7, 
      q_1_6=>que_out_25_1_6, q_1_5=>que_out_25_1_5, q_1_4=>que_out_25_1_4, 
      q_1_3=>que_out_25_1_3, q_1_2=>que_out_25_1_2, q_1_1=>que_out_25_1_1, 
      q_1_0=>que_out_25_1_0, q_2_15=>que_out_25_2_15, q_2_14=>
      que_out_25_2_14, q_2_13=>que_out_25_2_13, q_2_12=>que_out_25_2_12, 
      q_2_11=>que_out_25_2_11, q_2_10=>que_out_25_2_10, q_2_9=>
      que_out_25_2_9, q_2_8=>que_out_25_2_8, q_2_7=>que_out_25_2_7, q_2_6=>
      que_out_25_2_6, q_2_5=>que_out_25_2_5, q_2_4=>que_out_25_2_4, q_2_3=>
      que_out_25_2_3, q_2_2=>que_out_25_2_2, q_2_1=>que_out_25_2_1, q_2_0=>
      que_out_25_2_0, q_3_15=>que_out_25_3_15, q_3_14=>que_out_25_3_14, 
      q_3_13=>que_out_25_3_13, q_3_12=>que_out_25_3_12, q_3_11=>
      que_out_25_3_11, q_3_10=>que_out_25_3_10, q_3_9=>que_out_25_3_9, q_3_8
      =>que_out_25_3_8, q_3_7=>que_out_25_3_7, q_3_6=>que_out_25_3_6, q_3_5
      =>que_out_25_3_5, q_3_4=>que_out_25_3_4, q_3_3=>que_out_25_3_3, q_3_2
      =>que_out_25_3_2, q_3_1=>que_out_25_3_1, q_3_0=>que_out_25_3_0, q_4_15
      =>que_out_25_4_15, q_4_14=>que_out_25_4_14, q_4_13=>que_out_25_4_13, 
      q_4_12=>que_out_25_4_12, q_4_11=>que_out_25_4_11, q_4_10=>
      que_out_25_4_10, q_4_9=>que_out_25_4_9, q_4_8=>que_out_25_4_8, q_4_7=>
      que_out_25_4_7, q_4_6=>que_out_25_4_6, q_4_5=>que_out_25_4_5, q_4_4=>
      que_out_25_4_4, q_4_3=>que_out_25_4_3, q_4_2=>que_out_25_4_2, q_4_1=>
      que_out_25_4_1, q_4_0=>que_out_25_4_0, clk=>nx10734, load=>sel_que_25, 
      reset=>nx10710);
   gen_queues_26_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_26_0_15, q_0_14=>que_out_26_0_14, q_0_13=>
      que_out_26_0_13, q_0_12=>que_out_26_0_12, q_0_11=>que_out_26_0_11, 
      q_0_10=>que_out_26_0_10, q_0_9=>que_out_26_0_9, q_0_8=>que_out_26_0_8, 
      q_0_7=>que_out_26_0_7, q_0_6=>que_out_26_0_6, q_0_5=>que_out_26_0_5, 
      q_0_4=>que_out_26_0_4, q_0_3=>que_out_26_0_3, q_0_2=>que_out_26_0_2, 
      q_0_1=>que_out_26_0_1, q_0_0=>que_out_26_0_0, q_1_15=>que_out_26_1_15, 
      q_1_14=>que_out_26_1_14, q_1_13=>que_out_26_1_13, q_1_12=>
      que_out_26_1_12, q_1_11=>que_out_26_1_11, q_1_10=>que_out_26_1_10, 
      q_1_9=>que_out_26_1_9, q_1_8=>que_out_26_1_8, q_1_7=>que_out_26_1_7, 
      q_1_6=>que_out_26_1_6, q_1_5=>que_out_26_1_5, q_1_4=>que_out_26_1_4, 
      q_1_3=>que_out_26_1_3, q_1_2=>que_out_26_1_2, q_1_1=>que_out_26_1_1, 
      q_1_0=>que_out_26_1_0, q_2_15=>que_out_26_2_15, q_2_14=>
      que_out_26_2_14, q_2_13=>que_out_26_2_13, q_2_12=>que_out_26_2_12, 
      q_2_11=>que_out_26_2_11, q_2_10=>que_out_26_2_10, q_2_9=>
      que_out_26_2_9, q_2_8=>que_out_26_2_8, q_2_7=>que_out_26_2_7, q_2_6=>
      que_out_26_2_6, q_2_5=>que_out_26_2_5, q_2_4=>que_out_26_2_4, q_2_3=>
      que_out_26_2_3, q_2_2=>que_out_26_2_2, q_2_1=>que_out_26_2_1, q_2_0=>
      que_out_26_2_0, q_3_15=>que_out_26_3_15, q_3_14=>que_out_26_3_14, 
      q_3_13=>que_out_26_3_13, q_3_12=>que_out_26_3_12, q_3_11=>
      que_out_26_3_11, q_3_10=>que_out_26_3_10, q_3_9=>que_out_26_3_9, q_3_8
      =>que_out_26_3_8, q_3_7=>que_out_26_3_7, q_3_6=>que_out_26_3_6, q_3_5
      =>que_out_26_3_5, q_3_4=>que_out_26_3_4, q_3_3=>que_out_26_3_3, q_3_2
      =>que_out_26_3_2, q_3_1=>que_out_26_3_1, q_3_0=>que_out_26_3_0, q_4_15
      =>que_out_26_4_15, q_4_14=>que_out_26_4_14, q_4_13=>que_out_26_4_13, 
      q_4_12=>que_out_26_4_12, q_4_11=>que_out_26_4_11, q_4_10=>
      que_out_26_4_10, q_4_9=>que_out_26_4_9, q_4_8=>que_out_26_4_8, q_4_7=>
      que_out_26_4_7, q_4_6=>que_out_26_4_6, q_4_5=>que_out_26_4_5, q_4_4=>
      que_out_26_4_4, q_4_3=>que_out_26_4_3, q_4_2=>que_out_26_4_2, q_4_1=>
      que_out_26_4_1, q_4_0=>que_out_26_4_0, clk=>nx10734, load=>sel_que_26, 
      reset=>nx10710);
   gen_queues_27_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_27_0_15, q_0_14=>que_out_27_0_14, q_0_13=>
      que_out_27_0_13, q_0_12=>que_out_27_0_12, q_0_11=>que_out_27_0_11, 
      q_0_10=>que_out_27_0_10, q_0_9=>que_out_27_0_9, q_0_8=>que_out_27_0_8, 
      q_0_7=>que_out_27_0_7, q_0_6=>que_out_27_0_6, q_0_5=>que_out_27_0_5, 
      q_0_4=>que_out_27_0_4, q_0_3=>que_out_27_0_3, q_0_2=>que_out_27_0_2, 
      q_0_1=>que_out_27_0_1, q_0_0=>que_out_27_0_0, q_1_15=>que_out_27_1_15, 
      q_1_14=>que_out_27_1_14, q_1_13=>que_out_27_1_13, q_1_12=>
      que_out_27_1_12, q_1_11=>que_out_27_1_11, q_1_10=>que_out_27_1_10, 
      q_1_9=>que_out_27_1_9, q_1_8=>que_out_27_1_8, q_1_7=>que_out_27_1_7, 
      q_1_6=>que_out_27_1_6, q_1_5=>que_out_27_1_5, q_1_4=>que_out_27_1_4, 
      q_1_3=>que_out_27_1_3, q_1_2=>que_out_27_1_2, q_1_1=>que_out_27_1_1, 
      q_1_0=>que_out_27_1_0, q_2_15=>que_out_27_2_15, q_2_14=>
      que_out_27_2_14, q_2_13=>que_out_27_2_13, q_2_12=>que_out_27_2_12, 
      q_2_11=>que_out_27_2_11, q_2_10=>que_out_27_2_10, q_2_9=>
      que_out_27_2_9, q_2_8=>que_out_27_2_8, q_2_7=>que_out_27_2_7, q_2_6=>
      que_out_27_2_6, q_2_5=>que_out_27_2_5, q_2_4=>que_out_27_2_4, q_2_3=>
      que_out_27_2_3, q_2_2=>que_out_27_2_2, q_2_1=>que_out_27_2_1, q_2_0=>
      que_out_27_2_0, q_3_15=>que_out_27_3_15, q_3_14=>que_out_27_3_14, 
      q_3_13=>que_out_27_3_13, q_3_12=>que_out_27_3_12, q_3_11=>
      que_out_27_3_11, q_3_10=>que_out_27_3_10, q_3_9=>que_out_27_3_9, q_3_8
      =>que_out_27_3_8, q_3_7=>que_out_27_3_7, q_3_6=>que_out_27_3_6, q_3_5
      =>que_out_27_3_5, q_3_4=>que_out_27_3_4, q_3_3=>que_out_27_3_3, q_3_2
      =>que_out_27_3_2, q_3_1=>que_out_27_3_1, q_3_0=>que_out_27_3_0, q_4_15
      =>que_out_27_4_15, q_4_14=>que_out_27_4_14, q_4_13=>que_out_27_4_13, 
      q_4_12=>que_out_27_4_12, q_4_11=>que_out_27_4_11, q_4_10=>
      que_out_27_4_10, q_4_9=>que_out_27_4_9, q_4_8=>que_out_27_4_8, q_4_7=>
      que_out_27_4_7, q_4_6=>que_out_27_4_6, q_4_5=>que_out_27_4_5, q_4_4=>
      que_out_27_4_4, q_4_3=>que_out_27_4_3, q_4_2=>que_out_27_4_2, q_4_1=>
      que_out_27_4_1, q_4_0=>que_out_27_4_0, clk=>nx10736, load=>sel_que_27, 
      reset=>nx10712);
   ix6830 : nand03 port map ( Y=>nx6829, A0=>nx8938, A1=>nx6833, A2=>nx6835
   );
   ix8939 : nor02ii port map ( Y=>nx8938, A0=>cache_in_sel(4), A1=>
      decoder_enable);
   ix6834 : inv01 port map ( Y=>nx6833, A=>cache_in_sel(1));
   ix6836 : inv01 port map ( Y=>nx6835, A=>cache_in_sel(0));
   ix6840 : nand03 port map ( Y=>nx6839, A0=>nx8938, A1=>nx6833, A2=>nx10508
   );
   ix6844 : nand03 port map ( Y=>nx6843, A0=>nx8938, A1=>nx10506, A2=>nx6835
   );
   ix6848 : nand03 port map ( Y=>nx6847, A0=>nx8938, A1=>nx10506, A2=>
      nx10508);
   ix9023 : nor02_2x port map ( Y=>sel_que_12, A0=>nx6875, A1=>nx6829);
   ix6876 : nand02 port map ( Y=>nx6875, A0=>cache_in_sel(3), A1=>
      cache_in_sel(2));
   ix9025 : nor02_2x port map ( Y=>sel_que_13, A0=>nx6875, A1=>nx6839);
   ix9027 : nor02_2x port map ( Y=>sel_que_14, A0=>nx6843, A1=>nx6875);
   ix9029 : nor02_2x port map ( Y=>sel_que_15, A0=>nx6875, A1=>nx6847);
   ix9043 : and02 port map ( Y=>sel_que_16, A0=>nx6885, A1=>nx9038);
   ix6886 : nor02_2x port map ( Y=>nx6885, A0=>cache_in_sel(2), A1=>
      cache_in_sel(3));
   ix9039 : nor03_2x port map ( Y=>nx9038, A0=>nx6889, A1=>nx10506, A2=>
      nx10508);
   ix6890 : nand02 port map ( Y=>nx6889, A0=>cache_in_sel(4), A1=>
      decoder_enable);
   ix6894 : nand04 port map ( Y=>nx6893, A0=>cache_in_sel(4), A1=>
      decoder_enable, A2=>nx6833, A3=>nx10508);
   ix6898 : nand04 port map ( Y=>nx6897, A0=>cache_in_sel(4), A1=>
      decoder_enable, A2=>nx10506, A3=>nx6835);
   ix6902 : nand04 port map ( Y=>nx6901, A0=>cache_in_sel(4), A1=>
      decoder_enable, A2=>nx10506, A3=>nx10508);
   ix9075 : and02 port map ( Y=>sel_que_20, A0=>nx6905, A1=>nx9038);
   ix9091 : and02 port map ( Y=>sel_que_24, A0=>nx6915, A1=>nx9038);
   ix243 : or04 port map ( Y=>out_column_4_0, A0=>nx238, A1=>nx188, A2=>
      nx130, A3=>nx82);
   ix239 : nand03 port map ( Y=>nx238, A0=>nx6927, A1=>nx6951, A2=>nx6967);
   ix6928 : aoi222 port map ( Y=>nx6927, A0=>que_out_10_4_0, A1=>nx10298, B0
      =>que_out_6_4_0, B1=>nx10350, C0=>que_out_9_4_0, C1=>nx10324);
   ix6932 : nand02_2x port map ( Y=>nx6931, A0=>cache_out_sel(3), A1=>nx6933
   );
   ix6934 : inv01 port map ( Y=>nx6933, A=>cache_out_sel(0));
   ix6938 : inv01 port map ( Y=>nx6937, A=>cache_out_sel(4));
   ix6940 : inv02 port map ( Y=>nx6939, A=>cache_out_sel(2));
   ix6946 : nand03 port map ( Y=>nx6945, A0=>nx10502, A1=>nx6937, A2=>
      nx10498);
   ix227 : nor04 port map ( Y=>nx226, A0=>nx6949, A1=>nx10502, A2=>nx10494, 
      A3=>nx10498);
   ix6950 : nand02_2x port map ( Y=>nx6949, A0=>cache_out_sel(3), A1=>
      cache_out_sel(0));
   ix6952 : aoi22 port map ( Y=>nx6951, A0=>que_out_5_4_0, A1=>nx10246, B0=>
      que_out_18_4_0, B1=>nx10272);
   ix6956 : nand02 port map ( Y=>nx6955, A0=>nx6957, A1=>cache_out_sel(0));
   ix6958 : inv01 port map ( Y=>nx6957, A=>cache_out_sel(3));
   ix6962 : inv01 port map ( Y=>nx6961, A=>cache_out_sel(1));
   ix215 : nor03_2x port map ( Y=>nx214, A0=>nx6965, A1=>nx10498, A2=>nx6943
   );
   ix6966 : nand02_2x port map ( Y=>nx6965, A0=>nx10494, A1=>nx10504);
   ix6968 : aoi22 port map ( Y=>nx6967, A0=>que_out_17_4_0, A1=>nx10220, B0
      =>que_out_20_4_0, B1=>nx10194);
   ix201 : nor03_2x port map ( Y=>nx200, A0=>nx6971, A1=>nx10498, A2=>
      nx10374);
   ix6972 : nand02_2x port map ( Y=>nx6971, A0=>nx10496, A1=>nx6961);
   ix193 : nor03_2x port map ( Y=>nx192, A0=>nx6971, A1=>nx6939, A2=>nx6943
   );
   ix189 : nand03 port map ( Y=>nx188, A0=>nx6977, A1=>nx6985, A2=>nx6991);
   ix6978 : aoi222 port map ( Y=>nx6977, A0=>que_out_19_4_0, A1=>nx10168, B0
      =>que_out_21_4_0, B1=>nx10142, C0=>que_out_8_4_0, C1=>nx10116);
   ix181 : nor03_2x port map ( Y=>nx180, A0=>nx6965, A1=>nx10498, A2=>
      nx10374);
   ix173 : nor03_2x port map ( Y=>nx172, A0=>nx6971, A1=>nx6939, A2=>nx10374
   );
   ix167 : nor04 port map ( Y=>nx166, A0=>nx6931, A1=>nx10502, A2=>nx10494, 
      A3=>nx10498);
   ix6986 : aoi22 port map ( Y=>nx6985, A0=>que_out_25_4_0, A1=>nx10064, B0
      =>que_out_16_4_0, B1=>nx10090);
   ix151 : nor02_2x port map ( Y=>nx150, A0=>nx6949, A1=>nx6971);
   ix159 : nor03_2x port map ( Y=>nx158, A0=>nx6971, A1=>nx10498, A2=>nx6943
   );
   ix6992 : aoi22 port map ( Y=>nx6991, A0=>que_out_24_4_0, A1=>nx10038, B0
      =>que_out_22_4_0, B1=>nx10012);
   ix145 : nor02_2x port map ( Y=>nx144, A0=>nx6971, A1=>nx6931);
   ix137 : nor03_2x port map ( Y=>nx136, A0=>nx6965, A1=>nx6939, A2=>nx6943
   );
   ix131 : nand03 port map ( Y=>nx130, A0=>nx6999, A1=>nx7007, A2=>nx7017);
   ix7000 : aoi222 port map ( Y=>nx6999, A0=>que_out_15_4_0, A1=>nx9960, B0
      =>que_out_3_4_0, B1=>nx9986, C0=>que_out_23_4_0, C1=>nx9934);
   ix119 : nor02_2x port map ( Y=>nx118, A0=>nx6949, A1=>nx6945);
   ix115 : nor03_2x port map ( Y=>nx114, A0=>nx6965, A1=>nx6939, A2=>nx10374
   );
   ix7008 : aoi22 port map ( Y=>nx7007, A0=>que_out_27_4_0, A1=>nx9908, B0=>
      que_out_4_4_0, B1=>nx9882);
   ix105 : nor02_2x port map ( Y=>nx104, A0=>nx6949, A1=>nx6965);
   ix101 : and02 port map ( Y=>nx100, A0=>nx88, A1=>nx28);
   ix89 : nor02_2x port map ( Y=>nx88, A0=>cache_out_sel(3), A1=>
      cache_out_sel(0));
   ix29 : nor03_2x port map ( Y=>nx28, A0=>nx10502, A1=>nx10494, A2=>nx6939
   );
   ix7018 : aoi22 port map ( Y=>nx7017, A0=>que_out_0_4_0, A1=>nx9830, B0=>
      que_out_2_4_0, B1=>nx9856);
   ix91 : and02 port map ( Y=>nx90, A0=>nx88, A1=>nx12);
   ix13 : nor03_2x port map ( Y=>nx12, A0=>nx10504, A1=>nx10494, A2=>nx10500
   );
   ix95 : and02 port map ( Y=>nx94, A0=>nx88, A1=>nx62);
   ix63 : nor03_2x port map ( Y=>nx62, A0=>nx6961, A1=>nx10494, A2=>nx10500
   );
   ix83 : nand03 port map ( Y=>nx82, A0=>nx7029, A1=>nx7037, A2=>nx7043);
   ix7030 : aoi222 port map ( Y=>nx7029, A0=>que_out_26_4_0, A1=>nx9804, B0
      =>que_out_14_4_0, B1=>nx9778, C0=>que_out_11_4_0, C1=>nx9752);
   ix75 : nor02_2x port map ( Y=>nx74, A0=>nx6965, A1=>nx6931);
   ix69 : nor02_2x port map ( Y=>nx68, A0=>nx6931, A1=>nx6945);
   ix7038 : aoi22 port map ( Y=>nx7037, A0=>que_out_13_4_0, A1=>nx9726, B0=>
      que_out_7_4_0, B1=>nx9700);
   ix43 : nor02_2x port map ( Y=>nx42, A0=>nx10374, A1=>nx6945);
   ix7044 : aoi22 port map ( Y=>nx7043, A0=>que_out_12_4_0, A1=>nx9674, B0=>
      que_out_1_4_0, B1=>nx9648);
   ix15 : nor04 port map ( Y=>nx14, A0=>nx10376, A1=>nx10504, A2=>nx10494, 
      A3=>nx10500);
   ix353 : or04 port map ( Y=>out_column_4_1, A0=>nx348, A1=>nx322, A2=>
      nx294, A3=>nx268);
   ix349 : nand03 port map ( Y=>nx348, A0=>nx7053, A1=>nx7055, A2=>nx7057);
   ix7054 : aoi222 port map ( Y=>nx7053, A0=>que_out_10_4_1, A1=>nx10298, B0
      =>que_out_6_4_1, B1=>nx10350, C0=>que_out_9_4_1, C1=>nx10324);
   ix7056 : aoi22 port map ( Y=>nx7055, A0=>que_out_5_4_1, A1=>nx10246, B0=>
      que_out_18_4_1, B1=>nx10272);
   ix7058 : aoi22 port map ( Y=>nx7057, A0=>que_out_17_4_1, A1=>nx10220, B0
      =>que_out_20_4_1, B1=>nx10194);
   ix323 : nand03 port map ( Y=>nx322, A0=>nx7061, A1=>nx7063, A2=>nx7065);
   ix7062 : aoi222 port map ( Y=>nx7061, A0=>que_out_19_4_1, A1=>nx10168, B0
      =>que_out_21_4_1, B1=>nx10142, C0=>que_out_8_4_1, C1=>nx10116);
   ix7064 : aoi22 port map ( Y=>nx7063, A0=>que_out_25_4_1, A1=>nx10064, B0
      =>que_out_16_4_1, B1=>nx10090);
   ix7066 : aoi22 port map ( Y=>nx7065, A0=>que_out_24_4_1, A1=>nx10038, B0
      =>que_out_22_4_1, B1=>nx10012);
   ix295 : nand03 port map ( Y=>nx294, A0=>nx7069, A1=>nx7071, A2=>nx7073);
   ix7070 : aoi222 port map ( Y=>nx7069, A0=>que_out_15_4_1, A1=>nx9960, B0
      =>que_out_3_4_1, B1=>nx9986, C0=>que_out_23_4_1, C1=>nx9934);
   ix7072 : aoi22 port map ( Y=>nx7071, A0=>que_out_27_4_1, A1=>nx9908, B0=>
      que_out_4_4_1, B1=>nx9882);
   ix7074 : aoi22 port map ( Y=>nx7073, A0=>que_out_0_4_1, A1=>nx9830, B0=>
      que_out_2_4_1, B1=>nx9856);
   ix269 : nand03 port map ( Y=>nx268, A0=>nx7077, A1=>nx7079, A2=>nx7081);
   ix7078 : aoi222 port map ( Y=>nx7077, A0=>que_out_26_4_1, A1=>nx9804, B0
      =>que_out_14_4_1, B1=>nx9778, C0=>que_out_11_4_1, C1=>nx9752);
   ix7080 : aoi22 port map ( Y=>nx7079, A0=>que_out_13_4_1, A1=>nx9726, B0=>
      que_out_7_4_1, B1=>nx9700);
   ix7082 : aoi22 port map ( Y=>nx7081, A0=>que_out_12_4_1, A1=>nx9674, B0=>
      que_out_1_4_1, B1=>nx9648);
   ix463 : or04 port map ( Y=>out_column_4_2, A0=>nx458, A1=>nx432, A2=>
      nx404, A3=>nx378);
   ix459 : nand03 port map ( Y=>nx458, A0=>nx7087, A1=>nx7089, A2=>nx7091);
   ix7088 : aoi222 port map ( Y=>nx7087, A0=>que_out_10_4_2, A1=>nx10298, B0
      =>que_out_6_4_2, B1=>nx10350, C0=>que_out_9_4_2, C1=>nx10324);
   ix7090 : aoi22 port map ( Y=>nx7089, A0=>que_out_5_4_2, A1=>nx10246, B0=>
      que_out_18_4_2, B1=>nx10272);
   ix7092 : aoi22 port map ( Y=>nx7091, A0=>que_out_17_4_2, A1=>nx10220, B0
      =>que_out_20_4_2, B1=>nx10194);
   ix433 : nand03 port map ( Y=>nx432, A0=>nx7095, A1=>nx7097, A2=>nx7099);
   ix7096 : aoi222 port map ( Y=>nx7095, A0=>que_out_19_4_2, A1=>nx10168, B0
      =>que_out_21_4_2, B1=>nx10142, C0=>que_out_8_4_2, C1=>nx10116);
   ix7098 : aoi22 port map ( Y=>nx7097, A0=>que_out_25_4_2, A1=>nx10064, B0
      =>que_out_16_4_2, B1=>nx10090);
   ix7100 : aoi22 port map ( Y=>nx7099, A0=>que_out_24_4_2, A1=>nx10038, B0
      =>que_out_22_4_2, B1=>nx10012);
   ix405 : nand03 port map ( Y=>nx404, A0=>nx7103, A1=>nx7105, A2=>nx7107);
   ix7104 : aoi222 port map ( Y=>nx7103, A0=>que_out_15_4_2, A1=>nx9960, B0
      =>que_out_3_4_2, B1=>nx9986, C0=>que_out_23_4_2, C1=>nx9934);
   ix7106 : aoi22 port map ( Y=>nx7105, A0=>que_out_27_4_2, A1=>nx9908, B0=>
      que_out_4_4_2, B1=>nx9882);
   ix7108 : aoi22 port map ( Y=>nx7107, A0=>que_out_0_4_2, A1=>nx9830, B0=>
      que_out_2_4_2, B1=>nx9856);
   ix379 : nand03 port map ( Y=>nx378, A0=>nx7111, A1=>nx7113, A2=>nx7115);
   ix7112 : aoi222 port map ( Y=>nx7111, A0=>que_out_26_4_2, A1=>nx9804, B0
      =>que_out_14_4_2, B1=>nx9778, C0=>que_out_11_4_2, C1=>nx9752);
   ix7114 : aoi22 port map ( Y=>nx7113, A0=>que_out_13_4_2, A1=>nx9726, B0=>
      que_out_7_4_2, B1=>nx9700);
   ix7116 : aoi22 port map ( Y=>nx7115, A0=>que_out_12_4_2, A1=>nx9674, B0=>
      que_out_1_4_2, B1=>nx9648);
   ix573 : or04 port map ( Y=>out_column_4_3, A0=>nx568, A1=>nx542, A2=>
      nx514, A3=>nx488);
   ix569 : nand03 port map ( Y=>nx568, A0=>nx7121, A1=>nx7123, A2=>nx7125);
   ix7122 : aoi222 port map ( Y=>nx7121, A0=>que_out_10_4_3, A1=>nx10298, B0
      =>que_out_6_4_3, B1=>nx10350, C0=>que_out_9_4_3, C1=>nx10324);
   ix7124 : aoi22 port map ( Y=>nx7123, A0=>que_out_5_4_3, A1=>nx10246, B0=>
      que_out_18_4_3, B1=>nx10272);
   ix7126 : aoi22 port map ( Y=>nx7125, A0=>que_out_17_4_3, A1=>nx10220, B0
      =>que_out_20_4_3, B1=>nx10194);
   ix543 : nand03 port map ( Y=>nx542, A0=>nx7129, A1=>nx7131, A2=>nx7133);
   ix7130 : aoi222 port map ( Y=>nx7129, A0=>que_out_19_4_3, A1=>nx10168, B0
      =>que_out_21_4_3, B1=>nx10142, C0=>que_out_8_4_3, C1=>nx10116);
   ix7132 : aoi22 port map ( Y=>nx7131, A0=>que_out_25_4_3, A1=>nx10064, B0
      =>que_out_16_4_3, B1=>nx10090);
   ix7134 : aoi22 port map ( Y=>nx7133, A0=>que_out_24_4_3, A1=>nx10038, B0
      =>que_out_22_4_3, B1=>nx10012);
   ix515 : nand03 port map ( Y=>nx514, A0=>nx7137, A1=>nx7139, A2=>nx7141);
   ix7138 : aoi222 port map ( Y=>nx7137, A0=>que_out_15_4_3, A1=>nx9960, B0
      =>que_out_3_4_3, B1=>nx9986, C0=>que_out_23_4_3, C1=>nx9934);
   ix7140 : aoi22 port map ( Y=>nx7139, A0=>que_out_27_4_3, A1=>nx9908, B0=>
      que_out_4_4_3, B1=>nx9882);
   ix7142 : aoi22 port map ( Y=>nx7141, A0=>que_out_0_4_3, A1=>nx9830, B0=>
      que_out_2_4_3, B1=>nx9856);
   ix489 : nand03 port map ( Y=>nx488, A0=>nx7145, A1=>nx7147, A2=>nx7149);
   ix7146 : aoi222 port map ( Y=>nx7145, A0=>que_out_26_4_3, A1=>nx9804, B0
      =>que_out_14_4_3, B1=>nx9778, C0=>que_out_11_4_3, C1=>nx9752);
   ix7148 : aoi22 port map ( Y=>nx7147, A0=>que_out_13_4_3, A1=>nx9726, B0=>
      que_out_7_4_3, B1=>nx9700);
   ix7150 : aoi22 port map ( Y=>nx7149, A0=>que_out_12_4_3, A1=>nx9674, B0=>
      que_out_1_4_3, B1=>nx9648);
   ix683 : or04 port map ( Y=>out_column_4_4, A0=>nx678, A1=>nx652, A2=>
      nx624, A3=>nx598);
   ix679 : nand03 port map ( Y=>nx678, A0=>nx7155, A1=>nx7157, A2=>nx7159);
   ix7156 : aoi222 port map ( Y=>nx7155, A0=>que_out_10_4_4, A1=>nx10298, B0
      =>que_out_6_4_4, B1=>nx10350, C0=>que_out_9_4_4, C1=>nx10324);
   ix7158 : aoi22 port map ( Y=>nx7157, A0=>que_out_5_4_4, A1=>nx10246, B0=>
      que_out_18_4_4, B1=>nx10272);
   ix7160 : aoi22 port map ( Y=>nx7159, A0=>que_out_17_4_4, A1=>nx10220, B0
      =>que_out_20_4_4, B1=>nx10194);
   ix653 : nand03 port map ( Y=>nx652, A0=>nx7163, A1=>nx7165, A2=>nx7167);
   ix7164 : aoi222 port map ( Y=>nx7163, A0=>que_out_19_4_4, A1=>nx10168, B0
      =>que_out_21_4_4, B1=>nx10142, C0=>que_out_8_4_4, C1=>nx10116);
   ix7166 : aoi22 port map ( Y=>nx7165, A0=>que_out_25_4_4, A1=>nx10064, B0
      =>que_out_16_4_4, B1=>nx10090);
   ix7168 : aoi22 port map ( Y=>nx7167, A0=>que_out_24_4_4, A1=>nx10038, B0
      =>que_out_22_4_4, B1=>nx10012);
   ix625 : nand03 port map ( Y=>nx624, A0=>nx7171, A1=>nx7173, A2=>nx7175);
   ix7172 : aoi222 port map ( Y=>nx7171, A0=>que_out_15_4_4, A1=>nx9960, B0
      =>que_out_3_4_4, B1=>nx9986, C0=>que_out_23_4_4, C1=>nx9934);
   ix7174 : aoi22 port map ( Y=>nx7173, A0=>que_out_27_4_4, A1=>nx9908, B0=>
      que_out_4_4_4, B1=>nx9882);
   ix7176 : aoi22 port map ( Y=>nx7175, A0=>que_out_0_4_4, A1=>nx9830, B0=>
      que_out_2_4_4, B1=>nx9856);
   ix599 : nand03 port map ( Y=>nx598, A0=>nx7179, A1=>nx7181, A2=>nx7183);
   ix7180 : aoi222 port map ( Y=>nx7179, A0=>que_out_26_4_4, A1=>nx9804, B0
      =>que_out_14_4_4, B1=>nx9778, C0=>que_out_11_4_4, C1=>nx9752);
   ix7182 : aoi22 port map ( Y=>nx7181, A0=>que_out_13_4_4, A1=>nx9726, B0=>
      que_out_7_4_4, B1=>nx9700);
   ix7184 : aoi22 port map ( Y=>nx7183, A0=>que_out_12_4_4, A1=>nx9674, B0=>
      que_out_1_4_4, B1=>nx9648);
   ix793 : or04 port map ( Y=>out_column_4_5, A0=>nx788, A1=>nx762, A2=>
      nx734, A3=>nx708);
   ix789 : nand03 port map ( Y=>nx788, A0=>nx7189, A1=>nx7191, A2=>nx7193);
   ix7190 : aoi222 port map ( Y=>nx7189, A0=>que_out_10_4_5, A1=>nx10298, B0
      =>que_out_6_4_5, B1=>nx10350, C0=>que_out_9_4_5, C1=>nx10324);
   ix7192 : aoi22 port map ( Y=>nx7191, A0=>que_out_5_4_5, A1=>nx10246, B0=>
      que_out_18_4_5, B1=>nx10272);
   ix7194 : aoi22 port map ( Y=>nx7193, A0=>que_out_17_4_5, A1=>nx10220, B0
      =>que_out_20_4_5, B1=>nx10194);
   ix763 : nand03 port map ( Y=>nx762, A0=>nx7197, A1=>nx7199, A2=>nx7201);
   ix7198 : aoi222 port map ( Y=>nx7197, A0=>que_out_19_4_5, A1=>nx10168, B0
      =>que_out_21_4_5, B1=>nx10142, C0=>que_out_8_4_5, C1=>nx10116);
   ix7200 : aoi22 port map ( Y=>nx7199, A0=>que_out_25_4_5, A1=>nx10064, B0
      =>que_out_16_4_5, B1=>nx10090);
   ix7202 : aoi22 port map ( Y=>nx7201, A0=>que_out_24_4_5, A1=>nx10038, B0
      =>que_out_22_4_5, B1=>nx10012);
   ix735 : nand03 port map ( Y=>nx734, A0=>nx7205, A1=>nx7207, A2=>nx7209);
   ix7206 : aoi222 port map ( Y=>nx7205, A0=>que_out_15_4_5, A1=>nx9960, B0
      =>que_out_3_4_5, B1=>nx9986, C0=>que_out_23_4_5, C1=>nx9934);
   ix7208 : aoi22 port map ( Y=>nx7207, A0=>que_out_27_4_5, A1=>nx9908, B0=>
      que_out_4_4_5, B1=>nx9882);
   ix7210 : aoi22 port map ( Y=>nx7209, A0=>que_out_0_4_5, A1=>nx9830, B0=>
      que_out_2_4_5, B1=>nx9856);
   ix709 : nand03 port map ( Y=>nx708, A0=>nx7213, A1=>nx7215, A2=>nx7217);
   ix7214 : aoi222 port map ( Y=>nx7213, A0=>que_out_26_4_5, A1=>nx9804, B0
      =>que_out_14_4_5, B1=>nx9778, C0=>que_out_11_4_5, C1=>nx9752);
   ix7216 : aoi22 port map ( Y=>nx7215, A0=>que_out_13_4_5, A1=>nx9726, B0=>
      que_out_7_4_5, B1=>nx9700);
   ix7218 : aoi22 port map ( Y=>nx7217, A0=>que_out_12_4_5, A1=>nx9674, B0=>
      que_out_1_4_5, B1=>nx9648);
   ix903 : or04 port map ( Y=>out_column_4_6, A0=>nx898, A1=>nx872, A2=>
      nx844, A3=>nx818);
   ix899 : nand03 port map ( Y=>nx898, A0=>nx7223, A1=>nx7225, A2=>nx7227);
   ix7224 : aoi222 port map ( Y=>nx7223, A0=>que_out_10_4_6, A1=>nx10298, B0
      =>que_out_6_4_6, B1=>nx10350, C0=>que_out_9_4_6, C1=>nx10324);
   ix7226 : aoi22 port map ( Y=>nx7225, A0=>que_out_5_4_6, A1=>nx10246, B0=>
      que_out_18_4_6, B1=>nx10272);
   ix7228 : aoi22 port map ( Y=>nx7227, A0=>que_out_17_4_6, A1=>nx10220, B0
      =>que_out_20_4_6, B1=>nx10194);
   ix873 : nand03 port map ( Y=>nx872, A0=>nx7231, A1=>nx7233, A2=>nx7235);
   ix7232 : aoi222 port map ( Y=>nx7231, A0=>que_out_19_4_6, A1=>nx10168, B0
      =>que_out_21_4_6, B1=>nx10142, C0=>que_out_8_4_6, C1=>nx10116);
   ix7234 : aoi22 port map ( Y=>nx7233, A0=>que_out_25_4_6, A1=>nx10064, B0
      =>que_out_16_4_6, B1=>nx10090);
   ix7236 : aoi22 port map ( Y=>nx7235, A0=>que_out_24_4_6, A1=>nx10038, B0
      =>que_out_22_4_6, B1=>nx10012);
   ix845 : nand03 port map ( Y=>nx844, A0=>nx7239, A1=>nx7241, A2=>nx7243);
   ix7240 : aoi222 port map ( Y=>nx7239, A0=>que_out_15_4_6, A1=>nx9960, B0
      =>que_out_3_4_6, B1=>nx9986, C0=>que_out_23_4_6, C1=>nx9934);
   ix7242 : aoi22 port map ( Y=>nx7241, A0=>que_out_27_4_6, A1=>nx9908, B0=>
      que_out_4_4_6, B1=>nx9882);
   ix7244 : aoi22 port map ( Y=>nx7243, A0=>que_out_0_4_6, A1=>nx9830, B0=>
      que_out_2_4_6, B1=>nx9856);
   ix819 : nand03 port map ( Y=>nx818, A0=>nx7247, A1=>nx7249, A2=>nx7251);
   ix7248 : aoi222 port map ( Y=>nx7247, A0=>que_out_26_4_6, A1=>nx9804, B0
      =>que_out_14_4_6, B1=>nx9778, C0=>que_out_11_4_6, C1=>nx9752);
   ix7250 : aoi22 port map ( Y=>nx7249, A0=>que_out_13_4_6, A1=>nx9726, B0=>
      que_out_7_4_6, B1=>nx9700);
   ix7252 : aoi22 port map ( Y=>nx7251, A0=>que_out_12_4_6, A1=>nx9674, B0=>
      que_out_1_4_6, B1=>nx9648);
   ix1013 : or04 port map ( Y=>out_column_4_7, A0=>nx1008, A1=>nx982, A2=>
      nx954, A3=>nx928);
   ix1009 : nand03 port map ( Y=>nx1008, A0=>nx7257, A1=>nx7259, A2=>nx7261
   );
   ix7258 : aoi222 port map ( Y=>nx7257, A0=>que_out_10_4_7, A1=>nx10300, B0
      =>que_out_6_4_7, B1=>nx10352, C0=>que_out_9_4_7, C1=>nx10326);
   ix7260 : aoi22 port map ( Y=>nx7259, A0=>que_out_5_4_7, A1=>nx10248, B0=>
      que_out_18_4_7, B1=>nx10274);
   ix7262 : aoi22 port map ( Y=>nx7261, A0=>que_out_17_4_7, A1=>nx10222, B0
      =>que_out_20_4_7, B1=>nx10196);
   ix983 : nand03 port map ( Y=>nx982, A0=>nx7265, A1=>nx7267, A2=>nx7269);
   ix7266 : aoi222 port map ( Y=>nx7265, A0=>que_out_19_4_7, A1=>nx10170, B0
      =>que_out_21_4_7, B1=>nx10144, C0=>que_out_8_4_7, C1=>nx10118);
   ix7268 : aoi22 port map ( Y=>nx7267, A0=>que_out_25_4_7, A1=>nx10066, B0
      =>que_out_16_4_7, B1=>nx10092);
   ix7270 : aoi22 port map ( Y=>nx7269, A0=>que_out_24_4_7, A1=>nx10040, B0
      =>que_out_22_4_7, B1=>nx10014);
   ix955 : nand03 port map ( Y=>nx954, A0=>nx7273, A1=>nx7275, A2=>nx7277);
   ix7274 : aoi222 port map ( Y=>nx7273, A0=>que_out_15_4_7, A1=>nx9962, B0
      =>que_out_3_4_7, B1=>nx9988, C0=>que_out_23_4_7, C1=>nx9936);
   ix7276 : aoi22 port map ( Y=>nx7275, A0=>que_out_27_4_7, A1=>nx9910, B0=>
      que_out_4_4_7, B1=>nx9884);
   ix7278 : aoi22 port map ( Y=>nx7277, A0=>que_out_0_4_7, A1=>nx9832, B0=>
      que_out_2_4_7, B1=>nx9858);
   ix929 : nand03 port map ( Y=>nx928, A0=>nx7281, A1=>nx7283, A2=>nx7285);
   ix7282 : aoi222 port map ( Y=>nx7281, A0=>que_out_26_4_7, A1=>nx9806, B0
      =>que_out_14_4_7, B1=>nx9780, C0=>que_out_11_4_7, C1=>nx9754);
   ix7284 : aoi22 port map ( Y=>nx7283, A0=>que_out_13_4_7, A1=>nx9728, B0=>
      que_out_7_4_7, B1=>nx9702);
   ix7286 : aoi22 port map ( Y=>nx7285, A0=>que_out_12_4_7, A1=>nx9676, B0=>
      que_out_1_4_7, B1=>nx9650);
   ix1123 : or04 port map ( Y=>out_column_4_8, A0=>nx1118, A1=>nx1092, A2=>
      nx1064, A3=>nx1038);
   ix1119 : nand03 port map ( Y=>nx1118, A0=>nx7291, A1=>nx7293, A2=>nx7295
   );
   ix7292 : aoi222 port map ( Y=>nx7291, A0=>que_out_10_4_8, A1=>nx10300, B0
      =>que_out_6_4_8, B1=>nx10352, C0=>que_out_9_4_8, C1=>nx10326);
   ix7294 : aoi22 port map ( Y=>nx7293, A0=>que_out_5_4_8, A1=>nx10248, B0=>
      que_out_18_4_8, B1=>nx10274);
   ix7296 : aoi22 port map ( Y=>nx7295, A0=>que_out_17_4_8, A1=>nx10222, B0
      =>que_out_20_4_8, B1=>nx10196);
   ix1093 : nand03 port map ( Y=>nx1092, A0=>nx7299, A1=>nx7301, A2=>nx7303
   );
   ix7300 : aoi222 port map ( Y=>nx7299, A0=>que_out_19_4_8, A1=>nx10170, B0
      =>que_out_21_4_8, B1=>nx10144, C0=>que_out_8_4_8, C1=>nx10118);
   ix7302 : aoi22 port map ( Y=>nx7301, A0=>que_out_25_4_8, A1=>nx10066, B0
      =>que_out_16_4_8, B1=>nx10092);
   ix7304 : aoi22 port map ( Y=>nx7303, A0=>que_out_24_4_8, A1=>nx10040, B0
      =>que_out_22_4_8, B1=>nx10014);
   ix1065 : nand03 port map ( Y=>nx1064, A0=>nx7307, A1=>nx7309, A2=>nx7311
   );
   ix7308 : aoi222 port map ( Y=>nx7307, A0=>que_out_15_4_8, A1=>nx9962, B0
      =>que_out_3_4_8, B1=>nx9988, C0=>que_out_23_4_8, C1=>nx9936);
   ix7310 : aoi22 port map ( Y=>nx7309, A0=>que_out_27_4_8, A1=>nx9910, B0=>
      que_out_4_4_8, B1=>nx9884);
   ix7312 : aoi22 port map ( Y=>nx7311, A0=>que_out_0_4_8, A1=>nx9832, B0=>
      que_out_2_4_8, B1=>nx9858);
   ix1039 : nand03 port map ( Y=>nx1038, A0=>nx7315, A1=>nx7317, A2=>nx7319
   );
   ix7316 : aoi222 port map ( Y=>nx7315, A0=>que_out_26_4_8, A1=>nx9806, B0
      =>que_out_14_4_8, B1=>nx9780, C0=>que_out_11_4_8, C1=>nx9754);
   ix7318 : aoi22 port map ( Y=>nx7317, A0=>que_out_13_4_8, A1=>nx9728, B0=>
      que_out_7_4_8, B1=>nx9702);
   ix7320 : aoi22 port map ( Y=>nx7319, A0=>que_out_12_4_8, A1=>nx9676, B0=>
      que_out_1_4_8, B1=>nx9650);
   ix1233 : or04 port map ( Y=>out_column_4_9, A0=>nx1228, A1=>nx1202, A2=>
      nx1174, A3=>nx1148);
   ix1229 : nand03 port map ( Y=>nx1228, A0=>nx7325, A1=>nx7327, A2=>nx7329
   );
   ix7326 : aoi222 port map ( Y=>nx7325, A0=>que_out_10_4_9, A1=>nx10300, B0
      =>que_out_6_4_9, B1=>nx10352, C0=>que_out_9_4_9, C1=>nx10326);
   ix7328 : aoi22 port map ( Y=>nx7327, A0=>que_out_5_4_9, A1=>nx10248, B0=>
      que_out_18_4_9, B1=>nx10274);
   ix7330 : aoi22 port map ( Y=>nx7329, A0=>que_out_17_4_9, A1=>nx10222, B0
      =>que_out_20_4_9, B1=>nx10196);
   ix1203 : nand03 port map ( Y=>nx1202, A0=>nx7333, A1=>nx7335, A2=>nx7337
   );
   ix7334 : aoi222 port map ( Y=>nx7333, A0=>que_out_19_4_9, A1=>nx10170, B0
      =>que_out_21_4_9, B1=>nx10144, C0=>que_out_8_4_9, C1=>nx10118);
   ix7336 : aoi22 port map ( Y=>nx7335, A0=>que_out_25_4_9, A1=>nx10066, B0
      =>que_out_16_4_9, B1=>nx10092);
   ix7338 : aoi22 port map ( Y=>nx7337, A0=>que_out_24_4_9, A1=>nx10040, B0
      =>que_out_22_4_9, B1=>nx10014);
   ix1175 : nand03 port map ( Y=>nx1174, A0=>nx7341, A1=>nx7343, A2=>nx7345
   );
   ix7342 : aoi222 port map ( Y=>nx7341, A0=>que_out_15_4_9, A1=>nx9962, B0
      =>que_out_3_4_9, B1=>nx9988, C0=>que_out_23_4_9, C1=>nx9936);
   ix7344 : aoi22 port map ( Y=>nx7343, A0=>que_out_27_4_9, A1=>nx9910, B0=>
      que_out_4_4_9, B1=>nx9884);
   ix7346 : aoi22 port map ( Y=>nx7345, A0=>que_out_0_4_9, A1=>nx9832, B0=>
      que_out_2_4_9, B1=>nx9858);
   ix1149 : nand03 port map ( Y=>nx1148, A0=>nx7349, A1=>nx7351, A2=>nx7353
   );
   ix7350 : aoi222 port map ( Y=>nx7349, A0=>que_out_26_4_9, A1=>nx9806, B0
      =>que_out_14_4_9, B1=>nx9780, C0=>que_out_11_4_9, C1=>nx9754);
   ix7352 : aoi22 port map ( Y=>nx7351, A0=>que_out_13_4_9, A1=>nx9728, B0=>
      que_out_7_4_9, B1=>nx9702);
   ix7354 : aoi22 port map ( Y=>nx7353, A0=>que_out_12_4_9, A1=>nx9676, B0=>
      que_out_1_4_9, B1=>nx9650);
   ix1343 : or04 port map ( Y=>out_column_4_10, A0=>nx1338, A1=>nx1312, A2=>
      nx1284, A3=>nx1258);
   ix1339 : nand03 port map ( Y=>nx1338, A0=>nx7359, A1=>nx7361, A2=>nx7363
   );
   ix7360 : aoi222 port map ( Y=>nx7359, A0=>que_out_10_4_10, A1=>nx10300, 
      B0=>que_out_6_4_10, B1=>nx10352, C0=>que_out_9_4_10, C1=>nx10326);
   ix7362 : aoi22 port map ( Y=>nx7361, A0=>que_out_5_4_10, A1=>nx10248, B0
      =>que_out_18_4_10, B1=>nx10274);
   ix7364 : aoi22 port map ( Y=>nx7363, A0=>que_out_17_4_10, A1=>nx10222, B0
      =>que_out_20_4_10, B1=>nx10196);
   ix1313 : nand03 port map ( Y=>nx1312, A0=>nx7367, A1=>nx7369, A2=>nx7371
   );
   ix7368 : aoi222 port map ( Y=>nx7367, A0=>que_out_19_4_10, A1=>nx10170, 
      B0=>que_out_21_4_10, B1=>nx10144, C0=>que_out_8_4_10, C1=>nx10118);
   ix7370 : aoi22 port map ( Y=>nx7369, A0=>que_out_25_4_10, A1=>nx10066, B0
      =>que_out_16_4_10, B1=>nx10092);
   ix7372 : aoi22 port map ( Y=>nx7371, A0=>que_out_24_4_10, A1=>nx10040, B0
      =>que_out_22_4_10, B1=>nx10014);
   ix1285 : nand03 port map ( Y=>nx1284, A0=>nx7375, A1=>nx7377, A2=>nx7379
   );
   ix7376 : aoi222 port map ( Y=>nx7375, A0=>que_out_15_4_10, A1=>nx9962, B0
      =>que_out_3_4_10, B1=>nx9988, C0=>que_out_23_4_10, C1=>nx9936);
   ix7378 : aoi22 port map ( Y=>nx7377, A0=>que_out_27_4_10, A1=>nx9910, B0
      =>que_out_4_4_10, B1=>nx9884);
   ix7380 : aoi22 port map ( Y=>nx7379, A0=>que_out_0_4_10, A1=>nx9832, B0=>
      que_out_2_4_10, B1=>nx9858);
   ix1259 : nand03 port map ( Y=>nx1258, A0=>nx7383, A1=>nx7385, A2=>nx7387
   );
   ix7384 : aoi222 port map ( Y=>nx7383, A0=>que_out_26_4_10, A1=>nx9806, B0
      =>que_out_14_4_10, B1=>nx9780, C0=>que_out_11_4_10, C1=>nx9754);
   ix7386 : aoi22 port map ( Y=>nx7385, A0=>que_out_13_4_10, A1=>nx9728, B0
      =>que_out_7_4_10, B1=>nx9702);
   ix7388 : aoi22 port map ( Y=>nx7387, A0=>que_out_12_4_10, A1=>nx9676, B0
      =>que_out_1_4_10, B1=>nx9650);
   ix1453 : or04 port map ( Y=>out_column_4_11, A0=>nx1448, A1=>nx1422, A2=>
      nx1394, A3=>nx1368);
   ix1449 : nand03 port map ( Y=>nx1448, A0=>nx7393, A1=>nx7395, A2=>nx7397
   );
   ix7394 : aoi222 port map ( Y=>nx7393, A0=>que_out_10_4_11, A1=>nx10300, 
      B0=>que_out_6_4_11, B1=>nx10352, C0=>que_out_9_4_11, C1=>nx10326);
   ix7396 : aoi22 port map ( Y=>nx7395, A0=>que_out_5_4_11, A1=>nx10248, B0
      =>que_out_18_4_11, B1=>nx10274);
   ix7398 : aoi22 port map ( Y=>nx7397, A0=>que_out_17_4_11, A1=>nx10222, B0
      =>que_out_20_4_11, B1=>nx10196);
   ix1423 : nand03 port map ( Y=>nx1422, A0=>nx7401, A1=>nx7403, A2=>nx7405
   );
   ix7402 : aoi222 port map ( Y=>nx7401, A0=>que_out_19_4_11, A1=>nx10170, 
      B0=>que_out_21_4_11, B1=>nx10144, C0=>que_out_8_4_11, C1=>nx10118);
   ix7404 : aoi22 port map ( Y=>nx7403, A0=>que_out_25_4_11, A1=>nx10066, B0
      =>que_out_16_4_11, B1=>nx10092);
   ix7406 : aoi22 port map ( Y=>nx7405, A0=>que_out_24_4_11, A1=>nx10040, B0
      =>que_out_22_4_11, B1=>nx10014);
   ix1395 : nand03 port map ( Y=>nx1394, A0=>nx7409, A1=>nx7411, A2=>nx7413
   );
   ix7410 : aoi222 port map ( Y=>nx7409, A0=>que_out_15_4_11, A1=>nx9962, B0
      =>que_out_3_4_11, B1=>nx9988, C0=>que_out_23_4_11, C1=>nx9936);
   ix7412 : aoi22 port map ( Y=>nx7411, A0=>que_out_27_4_11, A1=>nx9910, B0
      =>que_out_4_4_11, B1=>nx9884);
   ix7414 : aoi22 port map ( Y=>nx7413, A0=>que_out_0_4_11, A1=>nx9832, B0=>
      que_out_2_4_11, B1=>nx9858);
   ix1369 : nand03 port map ( Y=>nx1368, A0=>nx7417, A1=>nx7419, A2=>nx7421
   );
   ix7418 : aoi222 port map ( Y=>nx7417, A0=>que_out_26_4_11, A1=>nx9806, B0
      =>que_out_14_4_11, B1=>nx9780, C0=>que_out_11_4_11, C1=>nx9754);
   ix7420 : aoi22 port map ( Y=>nx7419, A0=>que_out_13_4_11, A1=>nx9728, B0
      =>que_out_7_4_11, B1=>nx9702);
   ix7422 : aoi22 port map ( Y=>nx7421, A0=>que_out_12_4_11, A1=>nx9676, B0
      =>que_out_1_4_11, B1=>nx9650);
   ix1563 : or04 port map ( Y=>out_column_4_12, A0=>nx1558, A1=>nx1532, A2=>
      nx1504, A3=>nx1478);
   ix1559 : nand03 port map ( Y=>nx1558, A0=>nx7427, A1=>nx7429, A2=>nx7431
   );
   ix7428 : aoi222 port map ( Y=>nx7427, A0=>que_out_10_4_12, A1=>nx10300, 
      B0=>que_out_6_4_12, B1=>nx10352, C0=>que_out_9_4_12, C1=>nx10326);
   ix7430 : aoi22 port map ( Y=>nx7429, A0=>que_out_5_4_12, A1=>nx10248, B0
      =>que_out_18_4_12, B1=>nx10274);
   ix7432 : aoi22 port map ( Y=>nx7431, A0=>que_out_17_4_12, A1=>nx10222, B0
      =>que_out_20_4_12, B1=>nx10196);
   ix1533 : nand03 port map ( Y=>nx1532, A0=>nx7435, A1=>nx7437, A2=>nx7439
   );
   ix7436 : aoi222 port map ( Y=>nx7435, A0=>que_out_19_4_12, A1=>nx10170, 
      B0=>que_out_21_4_12, B1=>nx10144, C0=>que_out_8_4_12, C1=>nx10118);
   ix7438 : aoi22 port map ( Y=>nx7437, A0=>que_out_25_4_12, A1=>nx10066, B0
      =>que_out_16_4_12, B1=>nx10092);
   ix7440 : aoi22 port map ( Y=>nx7439, A0=>que_out_24_4_12, A1=>nx10040, B0
      =>que_out_22_4_12, B1=>nx10014);
   ix1505 : nand03 port map ( Y=>nx1504, A0=>nx7443, A1=>nx7445, A2=>nx7447
   );
   ix7444 : aoi222 port map ( Y=>nx7443, A0=>que_out_15_4_12, A1=>nx9962, B0
      =>que_out_3_4_12, B1=>nx9988, C0=>que_out_23_4_12, C1=>nx9936);
   ix7446 : aoi22 port map ( Y=>nx7445, A0=>que_out_27_4_12, A1=>nx9910, B0
      =>que_out_4_4_12, B1=>nx9884);
   ix7448 : aoi22 port map ( Y=>nx7447, A0=>que_out_0_4_12, A1=>nx9832, B0=>
      que_out_2_4_12, B1=>nx9858);
   ix1479 : nand03 port map ( Y=>nx1478, A0=>nx7451, A1=>nx7453, A2=>nx7455
   );
   ix7452 : aoi222 port map ( Y=>nx7451, A0=>que_out_26_4_12, A1=>nx9806, B0
      =>que_out_14_4_12, B1=>nx9780, C0=>que_out_11_4_12, C1=>nx9754);
   ix7454 : aoi22 port map ( Y=>nx7453, A0=>que_out_13_4_12, A1=>nx9728, B0
      =>que_out_7_4_12, B1=>nx9702);
   ix7456 : aoi22 port map ( Y=>nx7455, A0=>que_out_12_4_12, A1=>nx9676, B0
      =>que_out_1_4_12, B1=>nx9650);
   ix1673 : or04 port map ( Y=>out_column_4_13, A0=>nx1668, A1=>nx1642, A2=>
      nx1614, A3=>nx1588);
   ix1669 : nand03 port map ( Y=>nx1668, A0=>nx7461, A1=>nx7463, A2=>nx7465
   );
   ix7462 : aoi222 port map ( Y=>nx7461, A0=>que_out_10_4_13, A1=>nx10300, 
      B0=>que_out_6_4_13, B1=>nx10352, C0=>que_out_9_4_13, C1=>nx10326);
   ix7464 : aoi22 port map ( Y=>nx7463, A0=>que_out_5_4_13, A1=>nx10248, B0
      =>que_out_18_4_13, B1=>nx10274);
   ix7466 : aoi22 port map ( Y=>nx7465, A0=>que_out_17_4_13, A1=>nx10222, B0
      =>que_out_20_4_13, B1=>nx10196);
   ix1643 : nand03 port map ( Y=>nx1642, A0=>nx7469, A1=>nx7471, A2=>nx7473
   );
   ix7470 : aoi222 port map ( Y=>nx7469, A0=>que_out_19_4_13, A1=>nx10170, 
      B0=>que_out_21_4_13, B1=>nx10144, C0=>que_out_8_4_13, C1=>nx10118);
   ix7472 : aoi22 port map ( Y=>nx7471, A0=>que_out_25_4_13, A1=>nx10066, B0
      =>que_out_16_4_13, B1=>nx10092);
   ix7474 : aoi22 port map ( Y=>nx7473, A0=>que_out_24_4_13, A1=>nx10040, B0
      =>que_out_22_4_13, B1=>nx10014);
   ix1615 : nand03 port map ( Y=>nx1614, A0=>nx7477, A1=>nx7479, A2=>nx7481
   );
   ix7478 : aoi222 port map ( Y=>nx7477, A0=>que_out_15_4_13, A1=>nx9962, B0
      =>que_out_3_4_13, B1=>nx9988, C0=>que_out_23_4_13, C1=>nx9936);
   ix7480 : aoi22 port map ( Y=>nx7479, A0=>que_out_27_4_13, A1=>nx9910, B0
      =>que_out_4_4_13, B1=>nx9884);
   ix7482 : aoi22 port map ( Y=>nx7481, A0=>que_out_0_4_13, A1=>nx9832, B0=>
      que_out_2_4_13, B1=>nx9858);
   ix1589 : nand03 port map ( Y=>nx1588, A0=>nx7485, A1=>nx7487, A2=>nx7489
   );
   ix7486 : aoi222 port map ( Y=>nx7485, A0=>que_out_26_4_13, A1=>nx9806, B0
      =>que_out_14_4_13, B1=>nx9780, C0=>que_out_11_4_13, C1=>nx9754);
   ix7488 : aoi22 port map ( Y=>nx7487, A0=>que_out_13_4_13, A1=>nx9728, B0
      =>que_out_7_4_13, B1=>nx9702);
   ix7490 : aoi22 port map ( Y=>nx7489, A0=>que_out_12_4_13, A1=>nx9676, B0
      =>que_out_1_4_13, B1=>nx9650);
   ix1783 : or04 port map ( Y=>out_column_4_14, A0=>nx1778, A1=>nx1752, A2=>
      nx1724, A3=>nx1698);
   ix1779 : nand03 port map ( Y=>nx1778, A0=>nx7495, A1=>nx7497, A2=>nx7499
   );
   ix7496 : aoi222 port map ( Y=>nx7495, A0=>que_out_10_4_14, A1=>nx10302, 
      B0=>que_out_6_4_14, B1=>nx10354, C0=>que_out_9_4_14, C1=>nx10328);
   ix7498 : aoi22 port map ( Y=>nx7497, A0=>que_out_5_4_14, A1=>nx10250, B0
      =>que_out_18_4_14, B1=>nx10276);
   ix7500 : aoi22 port map ( Y=>nx7499, A0=>que_out_17_4_14, A1=>nx10224, B0
      =>que_out_20_4_14, B1=>nx10198);
   ix1753 : nand03 port map ( Y=>nx1752, A0=>nx7503, A1=>nx7505, A2=>nx7507
   );
   ix7504 : aoi222 port map ( Y=>nx7503, A0=>que_out_19_4_14, A1=>nx10172, 
      B0=>que_out_21_4_14, B1=>nx10146, C0=>que_out_8_4_14, C1=>nx10120);
   ix7506 : aoi22 port map ( Y=>nx7505, A0=>que_out_25_4_14, A1=>nx10068, B0
      =>que_out_16_4_14, B1=>nx10094);
   ix7508 : aoi22 port map ( Y=>nx7507, A0=>que_out_24_4_14, A1=>nx10042, B0
      =>que_out_22_4_14, B1=>nx10016);
   ix1725 : nand03 port map ( Y=>nx1724, A0=>nx7511, A1=>nx7513, A2=>nx7515
   );
   ix7512 : aoi222 port map ( Y=>nx7511, A0=>que_out_15_4_14, A1=>nx9964, B0
      =>que_out_3_4_14, B1=>nx9990, C0=>que_out_23_4_14, C1=>nx9938);
   ix7514 : aoi22 port map ( Y=>nx7513, A0=>que_out_27_4_14, A1=>nx9912, B0
      =>que_out_4_4_14, B1=>nx9886);
   ix7516 : aoi22 port map ( Y=>nx7515, A0=>que_out_0_4_14, A1=>nx9834, B0=>
      que_out_2_4_14, B1=>nx9860);
   ix1699 : nand03 port map ( Y=>nx1698, A0=>nx7519, A1=>nx7521, A2=>nx7523
   );
   ix7520 : aoi222 port map ( Y=>nx7519, A0=>que_out_26_4_14, A1=>nx9808, B0
      =>que_out_14_4_14, B1=>nx9782, C0=>que_out_11_4_14, C1=>nx9756);
   ix7522 : aoi22 port map ( Y=>nx7521, A0=>que_out_13_4_14, A1=>nx9730, B0
      =>que_out_7_4_14, B1=>nx9704);
   ix7524 : aoi22 port map ( Y=>nx7523, A0=>que_out_12_4_14, A1=>nx9678, B0
      =>que_out_1_4_14, B1=>nx9652);
   ix1893 : or04 port map ( Y=>out_column_4_15, A0=>nx1888, A1=>nx1862, A2=>
      nx1834, A3=>nx1808);
   ix1889 : nand03 port map ( Y=>nx1888, A0=>nx7529, A1=>nx7531, A2=>nx7533
   );
   ix7530 : aoi222 port map ( Y=>nx7529, A0=>que_out_10_4_15, A1=>nx10302, 
      B0=>que_out_6_4_15, B1=>nx10354, C0=>que_out_9_4_15, C1=>nx10328);
   ix7532 : aoi22 port map ( Y=>nx7531, A0=>que_out_5_4_15, A1=>nx10250, B0
      =>que_out_18_4_15, B1=>nx10276);
   ix7534 : aoi22 port map ( Y=>nx7533, A0=>que_out_17_4_15, A1=>nx10224, B0
      =>que_out_20_4_15, B1=>nx10198);
   ix1863 : nand03 port map ( Y=>nx1862, A0=>nx7537, A1=>nx7539, A2=>nx7541
   );
   ix7538 : aoi222 port map ( Y=>nx7537, A0=>que_out_19_4_15, A1=>nx10172, 
      B0=>que_out_21_4_15, B1=>nx10146, C0=>que_out_8_4_15, C1=>nx10120);
   ix7540 : aoi22 port map ( Y=>nx7539, A0=>que_out_25_4_15, A1=>nx10068, B0
      =>que_out_16_4_15, B1=>nx10094);
   ix7542 : aoi22 port map ( Y=>nx7541, A0=>que_out_24_4_15, A1=>nx10042, B0
      =>que_out_22_4_15, B1=>nx10016);
   ix1835 : nand03 port map ( Y=>nx1834, A0=>nx7545, A1=>nx7547, A2=>nx7549
   );
   ix7546 : aoi222 port map ( Y=>nx7545, A0=>que_out_15_4_15, A1=>nx9964, B0
      =>que_out_3_4_15, B1=>nx9990, C0=>que_out_23_4_15, C1=>nx9938);
   ix7548 : aoi22 port map ( Y=>nx7547, A0=>que_out_27_4_15, A1=>nx9912, B0
      =>que_out_4_4_15, B1=>nx9886);
   ix7550 : aoi22 port map ( Y=>nx7549, A0=>que_out_0_4_15, A1=>nx9834, B0=>
      que_out_2_4_15, B1=>nx9860);
   ix1809 : nand03 port map ( Y=>nx1808, A0=>nx7553, A1=>nx7555, A2=>nx7557
   );
   ix7554 : aoi222 port map ( Y=>nx7553, A0=>que_out_26_4_15, A1=>nx9808, B0
      =>que_out_14_4_15, B1=>nx9782, C0=>que_out_11_4_15, C1=>nx9756);
   ix7556 : aoi22 port map ( Y=>nx7555, A0=>que_out_13_4_15, A1=>nx9730, B0
      =>que_out_7_4_15, B1=>nx9704);
   ix7558 : aoi22 port map ( Y=>nx7557, A0=>que_out_12_4_15, A1=>nx9678, B0
      =>que_out_1_4_15, B1=>nx9652);
   ix2003 : or04 port map ( Y=>out_column_3_0, A0=>nx1998, A1=>nx1972, A2=>
      nx1944, A3=>nx1918);
   ix1999 : nand03 port map ( Y=>nx1998, A0=>nx7563, A1=>nx7565, A2=>nx7567
   );
   ix7564 : aoi222 port map ( Y=>nx7563, A0=>que_out_10_3_0, A1=>nx10302, B0
      =>que_out_6_3_0, B1=>nx10354, C0=>que_out_9_3_0, C1=>nx10328);
   ix7566 : aoi22 port map ( Y=>nx7565, A0=>que_out_5_3_0, A1=>nx10250, B0=>
      que_out_18_3_0, B1=>nx10276);
   ix7568 : aoi22 port map ( Y=>nx7567, A0=>que_out_17_3_0, A1=>nx10224, B0
      =>que_out_20_3_0, B1=>nx10198);
   ix1973 : nand03 port map ( Y=>nx1972, A0=>nx7571, A1=>nx7573, A2=>nx7575
   );
   ix7572 : aoi222 port map ( Y=>nx7571, A0=>que_out_19_3_0, A1=>nx10172, B0
      =>que_out_21_3_0, B1=>nx10146, C0=>que_out_8_3_0, C1=>nx10120);
   ix7574 : aoi22 port map ( Y=>nx7573, A0=>que_out_25_3_0, A1=>nx10068, B0
      =>que_out_16_3_0, B1=>nx10094);
   ix7576 : aoi22 port map ( Y=>nx7575, A0=>que_out_24_3_0, A1=>nx10042, B0
      =>que_out_22_3_0, B1=>nx10016);
   ix1945 : nand03 port map ( Y=>nx1944, A0=>nx7579, A1=>nx7581, A2=>nx7583
   );
   ix7580 : aoi222 port map ( Y=>nx7579, A0=>que_out_15_3_0, A1=>nx9964, B0
      =>que_out_3_3_0, B1=>nx9990, C0=>que_out_23_3_0, C1=>nx9938);
   ix7582 : aoi22 port map ( Y=>nx7581, A0=>que_out_27_3_0, A1=>nx9912, B0=>
      que_out_4_3_0, B1=>nx9886);
   ix7584 : aoi22 port map ( Y=>nx7583, A0=>que_out_0_3_0, A1=>nx9834, B0=>
      que_out_2_3_0, B1=>nx9860);
   ix1919 : nand03 port map ( Y=>nx1918, A0=>nx7587, A1=>nx7589, A2=>nx7591
   );
   ix7588 : aoi222 port map ( Y=>nx7587, A0=>que_out_26_3_0, A1=>nx9808, B0
      =>que_out_14_3_0, B1=>nx9782, C0=>que_out_11_3_0, C1=>nx9756);
   ix7590 : aoi22 port map ( Y=>nx7589, A0=>que_out_13_3_0, A1=>nx9730, B0=>
      que_out_7_3_0, B1=>nx9704);
   ix7592 : aoi22 port map ( Y=>nx7591, A0=>que_out_12_3_0, A1=>nx9678, B0=>
      que_out_1_3_0, B1=>nx9652);
   ix2113 : or04 port map ( Y=>out_column_3_1, A0=>nx2108, A1=>nx2082, A2=>
      nx2054, A3=>nx2028);
   ix2109 : nand03 port map ( Y=>nx2108, A0=>nx7597, A1=>nx7599, A2=>nx7601
   );
   ix7598 : aoi222 port map ( Y=>nx7597, A0=>que_out_10_3_1, A1=>nx10302, B0
      =>que_out_6_3_1, B1=>nx10354, C0=>que_out_9_3_1, C1=>nx10328);
   ix7600 : aoi22 port map ( Y=>nx7599, A0=>que_out_5_3_1, A1=>nx10250, B0=>
      que_out_18_3_1, B1=>nx10276);
   ix7602 : aoi22 port map ( Y=>nx7601, A0=>que_out_17_3_1, A1=>nx10224, B0
      =>que_out_20_3_1, B1=>nx10198);
   ix2083 : nand03 port map ( Y=>nx2082, A0=>nx7605, A1=>nx7607, A2=>nx7609
   );
   ix7606 : aoi222 port map ( Y=>nx7605, A0=>que_out_19_3_1, A1=>nx10172, B0
      =>que_out_21_3_1, B1=>nx10146, C0=>que_out_8_3_1, C1=>nx10120);
   ix7608 : aoi22 port map ( Y=>nx7607, A0=>que_out_25_3_1, A1=>nx10068, B0
      =>que_out_16_3_1, B1=>nx10094);
   ix7610 : aoi22 port map ( Y=>nx7609, A0=>que_out_24_3_1, A1=>nx10042, B0
      =>que_out_22_3_1, B1=>nx10016);
   ix2055 : nand03 port map ( Y=>nx2054, A0=>nx7613, A1=>nx7615, A2=>nx7617
   );
   ix7614 : aoi222 port map ( Y=>nx7613, A0=>que_out_15_3_1, A1=>nx9964, B0
      =>que_out_3_3_1, B1=>nx9990, C0=>que_out_23_3_1, C1=>nx9938);
   ix7616 : aoi22 port map ( Y=>nx7615, A0=>que_out_27_3_1, A1=>nx9912, B0=>
      que_out_4_3_1, B1=>nx9886);
   ix7618 : aoi22 port map ( Y=>nx7617, A0=>que_out_0_3_1, A1=>nx9834, B0=>
      que_out_2_3_1, B1=>nx9860);
   ix2029 : nand03 port map ( Y=>nx2028, A0=>nx7621, A1=>nx7623, A2=>nx7625
   );
   ix7622 : aoi222 port map ( Y=>nx7621, A0=>que_out_26_3_1, A1=>nx9808, B0
      =>que_out_14_3_1, B1=>nx9782, C0=>que_out_11_3_1, C1=>nx9756);
   ix7624 : aoi22 port map ( Y=>nx7623, A0=>que_out_13_3_1, A1=>nx9730, B0=>
      que_out_7_3_1, B1=>nx9704);
   ix7626 : aoi22 port map ( Y=>nx7625, A0=>que_out_12_3_1, A1=>nx9678, B0=>
      que_out_1_3_1, B1=>nx9652);
   ix2223 : or04 port map ( Y=>out_column_3_2, A0=>nx2218, A1=>nx2192, A2=>
      nx2164, A3=>nx2138);
   ix2219 : nand03 port map ( Y=>nx2218, A0=>nx7631, A1=>nx7633, A2=>nx7635
   );
   ix7632 : aoi222 port map ( Y=>nx7631, A0=>que_out_10_3_2, A1=>nx10302, B0
      =>que_out_6_3_2, B1=>nx10354, C0=>que_out_9_3_2, C1=>nx10328);
   ix7634 : aoi22 port map ( Y=>nx7633, A0=>que_out_5_3_2, A1=>nx10250, B0=>
      que_out_18_3_2, B1=>nx10276);
   ix7636 : aoi22 port map ( Y=>nx7635, A0=>que_out_17_3_2, A1=>nx10224, B0
      =>que_out_20_3_2, B1=>nx10198);
   ix2193 : nand03 port map ( Y=>nx2192, A0=>nx7639, A1=>nx7641, A2=>nx7643
   );
   ix7640 : aoi222 port map ( Y=>nx7639, A0=>que_out_19_3_2, A1=>nx10172, B0
      =>que_out_21_3_2, B1=>nx10146, C0=>que_out_8_3_2, C1=>nx10120);
   ix7642 : aoi22 port map ( Y=>nx7641, A0=>que_out_25_3_2, A1=>nx10068, B0
      =>que_out_16_3_2, B1=>nx10094);
   ix7644 : aoi22 port map ( Y=>nx7643, A0=>que_out_24_3_2, A1=>nx10042, B0
      =>que_out_22_3_2, B1=>nx10016);
   ix2165 : nand03 port map ( Y=>nx2164, A0=>nx7647, A1=>nx7649, A2=>nx7651
   );
   ix7648 : aoi222 port map ( Y=>nx7647, A0=>que_out_15_3_2, A1=>nx9964, B0
      =>que_out_3_3_2, B1=>nx9990, C0=>que_out_23_3_2, C1=>nx9938);
   ix7650 : aoi22 port map ( Y=>nx7649, A0=>que_out_27_3_2, A1=>nx9912, B0=>
      que_out_4_3_2, B1=>nx9886);
   ix7652 : aoi22 port map ( Y=>nx7651, A0=>que_out_0_3_2, A1=>nx9834, B0=>
      que_out_2_3_2, B1=>nx9860);
   ix2139 : nand03 port map ( Y=>nx2138, A0=>nx7655, A1=>nx7657, A2=>nx7659
   );
   ix7656 : aoi222 port map ( Y=>nx7655, A0=>que_out_26_3_2, A1=>nx9808, B0
      =>que_out_14_3_2, B1=>nx9782, C0=>que_out_11_3_2, C1=>nx9756);
   ix7658 : aoi22 port map ( Y=>nx7657, A0=>que_out_13_3_2, A1=>nx9730, B0=>
      que_out_7_3_2, B1=>nx9704);
   ix7660 : aoi22 port map ( Y=>nx7659, A0=>que_out_12_3_2, A1=>nx9678, B0=>
      que_out_1_3_2, B1=>nx9652);
   ix2333 : or04 port map ( Y=>out_column_3_3, A0=>nx2328, A1=>nx2302, A2=>
      nx2274, A3=>nx2248);
   ix2329 : nand03 port map ( Y=>nx2328, A0=>nx7665, A1=>nx7667, A2=>nx7669
   );
   ix7666 : aoi222 port map ( Y=>nx7665, A0=>que_out_10_3_3, A1=>nx10302, B0
      =>que_out_6_3_3, B1=>nx10354, C0=>que_out_9_3_3, C1=>nx10328);
   ix7668 : aoi22 port map ( Y=>nx7667, A0=>que_out_5_3_3, A1=>nx10250, B0=>
      que_out_18_3_3, B1=>nx10276);
   ix7670 : aoi22 port map ( Y=>nx7669, A0=>que_out_17_3_3, A1=>nx10224, B0
      =>que_out_20_3_3, B1=>nx10198);
   ix2303 : nand03 port map ( Y=>nx2302, A0=>nx7673, A1=>nx7675, A2=>nx7677
   );
   ix7674 : aoi222 port map ( Y=>nx7673, A0=>que_out_19_3_3, A1=>nx10172, B0
      =>que_out_21_3_3, B1=>nx10146, C0=>que_out_8_3_3, C1=>nx10120);
   ix7676 : aoi22 port map ( Y=>nx7675, A0=>que_out_25_3_3, A1=>nx10068, B0
      =>que_out_16_3_3, B1=>nx10094);
   ix7678 : aoi22 port map ( Y=>nx7677, A0=>que_out_24_3_3, A1=>nx10042, B0
      =>que_out_22_3_3, B1=>nx10016);
   ix2275 : nand03 port map ( Y=>nx2274, A0=>nx7681, A1=>nx7683, A2=>nx7685
   );
   ix7682 : aoi222 port map ( Y=>nx7681, A0=>que_out_15_3_3, A1=>nx9964, B0
      =>que_out_3_3_3, B1=>nx9990, C0=>que_out_23_3_3, C1=>nx9938);
   ix7684 : aoi22 port map ( Y=>nx7683, A0=>que_out_27_3_3, A1=>nx9912, B0=>
      que_out_4_3_3, B1=>nx9886);
   ix7686 : aoi22 port map ( Y=>nx7685, A0=>que_out_0_3_3, A1=>nx9834, B0=>
      que_out_2_3_3, B1=>nx9860);
   ix2249 : nand03 port map ( Y=>nx2248, A0=>nx7689, A1=>nx7691, A2=>nx7693
   );
   ix7690 : aoi222 port map ( Y=>nx7689, A0=>que_out_26_3_3, A1=>nx9808, B0
      =>que_out_14_3_3, B1=>nx9782, C0=>que_out_11_3_3, C1=>nx9756);
   ix7692 : aoi22 port map ( Y=>nx7691, A0=>que_out_13_3_3, A1=>nx9730, B0=>
      que_out_7_3_3, B1=>nx9704);
   ix7694 : aoi22 port map ( Y=>nx7693, A0=>que_out_12_3_3, A1=>nx9678, B0=>
      que_out_1_3_3, B1=>nx9652);
   ix2443 : or04 port map ( Y=>out_column_3_4, A0=>nx2438, A1=>nx2412, A2=>
      nx2384, A3=>nx2358);
   ix2439 : nand03 port map ( Y=>nx2438, A0=>nx7699, A1=>nx7701, A2=>nx7703
   );
   ix7700 : aoi222 port map ( Y=>nx7699, A0=>que_out_10_3_4, A1=>nx10302, B0
      =>que_out_6_3_4, B1=>nx10354, C0=>que_out_9_3_4, C1=>nx10328);
   ix7702 : aoi22 port map ( Y=>nx7701, A0=>que_out_5_3_4, A1=>nx10250, B0=>
      que_out_18_3_4, B1=>nx10276);
   ix7704 : aoi22 port map ( Y=>nx7703, A0=>que_out_17_3_4, A1=>nx10224, B0
      =>que_out_20_3_4, B1=>nx10198);
   ix2413 : nand03 port map ( Y=>nx2412, A0=>nx7707, A1=>nx7709, A2=>nx7711
   );
   ix7708 : aoi222 port map ( Y=>nx7707, A0=>que_out_19_3_4, A1=>nx10172, B0
      =>que_out_21_3_4, B1=>nx10146, C0=>que_out_8_3_4, C1=>nx10120);
   ix7710 : aoi22 port map ( Y=>nx7709, A0=>que_out_25_3_4, A1=>nx10068, B0
      =>que_out_16_3_4, B1=>nx10094);
   ix7712 : aoi22 port map ( Y=>nx7711, A0=>que_out_24_3_4, A1=>nx10042, B0
      =>que_out_22_3_4, B1=>nx10016);
   ix2385 : nand03 port map ( Y=>nx2384, A0=>nx7715, A1=>nx7717, A2=>nx7719
   );
   ix7716 : aoi222 port map ( Y=>nx7715, A0=>que_out_15_3_4, A1=>nx9964, B0
      =>que_out_3_3_4, B1=>nx9990, C0=>que_out_23_3_4, C1=>nx9938);
   ix7718 : aoi22 port map ( Y=>nx7717, A0=>que_out_27_3_4, A1=>nx9912, B0=>
      que_out_4_3_4, B1=>nx9886);
   ix7720 : aoi22 port map ( Y=>nx7719, A0=>que_out_0_3_4, A1=>nx9834, B0=>
      que_out_2_3_4, B1=>nx9860);
   ix2359 : nand03 port map ( Y=>nx2358, A0=>nx7723, A1=>nx7725, A2=>nx7727
   );
   ix7724 : aoi222 port map ( Y=>nx7723, A0=>que_out_26_3_4, A1=>nx9808, B0
      =>que_out_14_3_4, B1=>nx9782, C0=>que_out_11_3_4, C1=>nx9756);
   ix7726 : aoi22 port map ( Y=>nx7725, A0=>que_out_13_3_4, A1=>nx9730, B0=>
      que_out_7_3_4, B1=>nx9704);
   ix7728 : aoi22 port map ( Y=>nx7727, A0=>que_out_12_3_4, A1=>nx9678, B0=>
      que_out_1_3_4, B1=>nx9652);
   ix2553 : or04 port map ( Y=>out_column_3_5, A0=>nx2548, A1=>nx2522, A2=>
      nx2494, A3=>nx2468);
   ix2549 : nand03 port map ( Y=>nx2548, A0=>nx7733, A1=>nx7735, A2=>nx7737
   );
   ix7734 : aoi222 port map ( Y=>nx7733, A0=>que_out_10_3_5, A1=>nx10304, B0
      =>que_out_6_3_5, B1=>nx10356, C0=>que_out_9_3_5, C1=>nx10330);
   ix7736 : aoi22 port map ( Y=>nx7735, A0=>que_out_5_3_5, A1=>nx10252, B0=>
      que_out_18_3_5, B1=>nx10278);
   ix7738 : aoi22 port map ( Y=>nx7737, A0=>que_out_17_3_5, A1=>nx10226, B0
      =>que_out_20_3_5, B1=>nx10200);
   ix2523 : nand03 port map ( Y=>nx2522, A0=>nx7741, A1=>nx7743, A2=>nx7745
   );
   ix7742 : aoi222 port map ( Y=>nx7741, A0=>que_out_19_3_5, A1=>nx10174, B0
      =>que_out_21_3_5, B1=>nx10148, C0=>que_out_8_3_5, C1=>nx10122);
   ix7744 : aoi22 port map ( Y=>nx7743, A0=>que_out_25_3_5, A1=>nx10070, B0
      =>que_out_16_3_5, B1=>nx10096);
   ix7746 : aoi22 port map ( Y=>nx7745, A0=>que_out_24_3_5, A1=>nx10044, B0
      =>que_out_22_3_5, B1=>nx10018);
   ix2495 : nand03 port map ( Y=>nx2494, A0=>nx7749, A1=>nx7751, A2=>nx7753
   );
   ix7750 : aoi222 port map ( Y=>nx7749, A0=>que_out_15_3_5, A1=>nx9966, B0
      =>que_out_3_3_5, B1=>nx9992, C0=>que_out_23_3_5, C1=>nx9940);
   ix7752 : aoi22 port map ( Y=>nx7751, A0=>que_out_27_3_5, A1=>nx9914, B0=>
      que_out_4_3_5, B1=>nx9888);
   ix7754 : aoi22 port map ( Y=>nx7753, A0=>que_out_0_3_5, A1=>nx9836, B0=>
      que_out_2_3_5, B1=>nx9862);
   ix2469 : nand03 port map ( Y=>nx2468, A0=>nx7757, A1=>nx7759, A2=>nx7761
   );
   ix7758 : aoi222 port map ( Y=>nx7757, A0=>que_out_26_3_5, A1=>nx9810, B0
      =>que_out_14_3_5, B1=>nx9784, C0=>que_out_11_3_5, C1=>nx9758);
   ix7760 : aoi22 port map ( Y=>nx7759, A0=>que_out_13_3_5, A1=>nx9732, B0=>
      que_out_7_3_5, B1=>nx9706);
   ix7762 : aoi22 port map ( Y=>nx7761, A0=>que_out_12_3_5, A1=>nx9680, B0=>
      que_out_1_3_5, B1=>nx9654);
   ix2663 : or04 port map ( Y=>out_column_3_6, A0=>nx2658, A1=>nx2632, A2=>
      nx2604, A3=>nx2578);
   ix2659 : nand03 port map ( Y=>nx2658, A0=>nx7767, A1=>nx7769, A2=>nx7771
   );
   ix7768 : aoi222 port map ( Y=>nx7767, A0=>que_out_10_3_6, A1=>nx10304, B0
      =>que_out_6_3_6, B1=>nx10356, C0=>que_out_9_3_6, C1=>nx10330);
   ix7770 : aoi22 port map ( Y=>nx7769, A0=>que_out_5_3_6, A1=>nx10252, B0=>
      que_out_18_3_6, B1=>nx10278);
   ix7772 : aoi22 port map ( Y=>nx7771, A0=>que_out_17_3_6, A1=>nx10226, B0
      =>que_out_20_3_6, B1=>nx10200);
   ix2633 : nand03 port map ( Y=>nx2632, A0=>nx7775, A1=>nx7777, A2=>nx7779
   );
   ix7776 : aoi222 port map ( Y=>nx7775, A0=>que_out_19_3_6, A1=>nx10174, B0
      =>que_out_21_3_6, B1=>nx10148, C0=>que_out_8_3_6, C1=>nx10122);
   ix7778 : aoi22 port map ( Y=>nx7777, A0=>que_out_25_3_6, A1=>nx10070, B0
      =>que_out_16_3_6, B1=>nx10096);
   ix7780 : aoi22 port map ( Y=>nx7779, A0=>que_out_24_3_6, A1=>nx10044, B0
      =>que_out_22_3_6, B1=>nx10018);
   ix2605 : nand03 port map ( Y=>nx2604, A0=>nx7783, A1=>nx7785, A2=>nx7787
   );
   ix7784 : aoi222 port map ( Y=>nx7783, A0=>que_out_15_3_6, A1=>nx9966, B0
      =>que_out_3_3_6, B1=>nx9992, C0=>que_out_23_3_6, C1=>nx9940);
   ix7786 : aoi22 port map ( Y=>nx7785, A0=>que_out_27_3_6, A1=>nx9914, B0=>
      que_out_4_3_6, B1=>nx9888);
   ix7788 : aoi22 port map ( Y=>nx7787, A0=>que_out_0_3_6, A1=>nx9836, B0=>
      que_out_2_3_6, B1=>nx9862);
   ix2579 : nand03 port map ( Y=>nx2578, A0=>nx7791, A1=>nx7793, A2=>nx7795
   );
   ix7792 : aoi222 port map ( Y=>nx7791, A0=>que_out_26_3_6, A1=>nx9810, B0
      =>que_out_14_3_6, B1=>nx9784, C0=>que_out_11_3_6, C1=>nx9758);
   ix7794 : aoi22 port map ( Y=>nx7793, A0=>que_out_13_3_6, A1=>nx9732, B0=>
      que_out_7_3_6, B1=>nx9706);
   ix7796 : aoi22 port map ( Y=>nx7795, A0=>que_out_12_3_6, A1=>nx9680, B0=>
      que_out_1_3_6, B1=>nx9654);
   ix2773 : or04 port map ( Y=>out_column_3_7, A0=>nx2768, A1=>nx2742, A2=>
      nx2714, A3=>nx2688);
   ix2769 : nand03 port map ( Y=>nx2768, A0=>nx7801, A1=>nx7803, A2=>nx7805
   );
   ix7802 : aoi222 port map ( Y=>nx7801, A0=>que_out_10_3_7, A1=>nx10304, B0
      =>que_out_6_3_7, B1=>nx10356, C0=>que_out_9_3_7, C1=>nx10330);
   ix7804 : aoi22 port map ( Y=>nx7803, A0=>que_out_5_3_7, A1=>nx10252, B0=>
      que_out_18_3_7, B1=>nx10278);
   ix7806 : aoi22 port map ( Y=>nx7805, A0=>que_out_17_3_7, A1=>nx10226, B0
      =>que_out_20_3_7, B1=>nx10200);
   ix2743 : nand03 port map ( Y=>nx2742, A0=>nx7809, A1=>nx7811, A2=>nx7813
   );
   ix7810 : aoi222 port map ( Y=>nx7809, A0=>que_out_19_3_7, A1=>nx10174, B0
      =>que_out_21_3_7, B1=>nx10148, C0=>que_out_8_3_7, C1=>nx10122);
   ix7812 : aoi22 port map ( Y=>nx7811, A0=>que_out_25_3_7, A1=>nx10070, B0
      =>que_out_16_3_7, B1=>nx10096);
   ix7814 : aoi22 port map ( Y=>nx7813, A0=>que_out_24_3_7, A1=>nx10044, B0
      =>que_out_22_3_7, B1=>nx10018);
   ix2715 : nand03 port map ( Y=>nx2714, A0=>nx7817, A1=>nx7819, A2=>nx7821
   );
   ix7818 : aoi222 port map ( Y=>nx7817, A0=>que_out_15_3_7, A1=>nx9966, B0
      =>que_out_3_3_7, B1=>nx9992, C0=>que_out_23_3_7, C1=>nx9940);
   ix7820 : aoi22 port map ( Y=>nx7819, A0=>que_out_27_3_7, A1=>nx9914, B0=>
      que_out_4_3_7, B1=>nx9888);
   ix7822 : aoi22 port map ( Y=>nx7821, A0=>que_out_0_3_7, A1=>nx9836, B0=>
      que_out_2_3_7, B1=>nx9862);
   ix2689 : nand03 port map ( Y=>nx2688, A0=>nx7825, A1=>nx7827, A2=>nx7829
   );
   ix7826 : aoi222 port map ( Y=>nx7825, A0=>que_out_26_3_7, A1=>nx9810, B0
      =>que_out_14_3_7, B1=>nx9784, C0=>que_out_11_3_7, C1=>nx9758);
   ix7828 : aoi22 port map ( Y=>nx7827, A0=>que_out_13_3_7, A1=>nx9732, B0=>
      que_out_7_3_7, B1=>nx9706);
   ix7830 : aoi22 port map ( Y=>nx7829, A0=>que_out_12_3_7, A1=>nx9680, B0=>
      que_out_1_3_7, B1=>nx9654);
   ix2883 : or04 port map ( Y=>out_column_3_8, A0=>nx2878, A1=>nx2852, A2=>
      nx2824, A3=>nx2798);
   ix2879 : nand03 port map ( Y=>nx2878, A0=>nx7835, A1=>nx7837, A2=>nx7839
   );
   ix7836 : aoi222 port map ( Y=>nx7835, A0=>que_out_10_3_8, A1=>nx10304, B0
      =>que_out_6_3_8, B1=>nx10356, C0=>que_out_9_3_8, C1=>nx10330);
   ix7838 : aoi22 port map ( Y=>nx7837, A0=>que_out_5_3_8, A1=>nx10252, B0=>
      que_out_18_3_8, B1=>nx10278);
   ix7840 : aoi22 port map ( Y=>nx7839, A0=>que_out_17_3_8, A1=>nx10226, B0
      =>que_out_20_3_8, B1=>nx10200);
   ix2853 : nand03 port map ( Y=>nx2852, A0=>nx7843, A1=>nx7845, A2=>nx7847
   );
   ix7844 : aoi222 port map ( Y=>nx7843, A0=>que_out_19_3_8, A1=>nx10174, B0
      =>que_out_21_3_8, B1=>nx10148, C0=>que_out_8_3_8, C1=>nx10122);
   ix7846 : aoi22 port map ( Y=>nx7845, A0=>que_out_25_3_8, A1=>nx10070, B0
      =>que_out_16_3_8, B1=>nx10096);
   ix7848 : aoi22 port map ( Y=>nx7847, A0=>que_out_24_3_8, A1=>nx10044, B0
      =>que_out_22_3_8, B1=>nx10018);
   ix2825 : nand03 port map ( Y=>nx2824, A0=>nx7851, A1=>nx7853, A2=>nx7855
   );
   ix7852 : aoi222 port map ( Y=>nx7851, A0=>que_out_15_3_8, A1=>nx9966, B0
      =>que_out_3_3_8, B1=>nx9992, C0=>que_out_23_3_8, C1=>nx9940);
   ix7854 : aoi22 port map ( Y=>nx7853, A0=>que_out_27_3_8, A1=>nx9914, B0=>
      que_out_4_3_8, B1=>nx9888);
   ix7856 : aoi22 port map ( Y=>nx7855, A0=>que_out_0_3_8, A1=>nx9836, B0=>
      que_out_2_3_8, B1=>nx9862);
   ix2799 : nand03 port map ( Y=>nx2798, A0=>nx7859, A1=>nx7861, A2=>nx7863
   );
   ix7860 : aoi222 port map ( Y=>nx7859, A0=>que_out_26_3_8, A1=>nx9810, B0
      =>que_out_14_3_8, B1=>nx9784, C0=>que_out_11_3_8, C1=>nx9758);
   ix7862 : aoi22 port map ( Y=>nx7861, A0=>que_out_13_3_8, A1=>nx9732, B0=>
      que_out_7_3_8, B1=>nx9706);
   ix7864 : aoi22 port map ( Y=>nx7863, A0=>que_out_12_3_8, A1=>nx9680, B0=>
      que_out_1_3_8, B1=>nx9654);
   ix2993 : or04 port map ( Y=>out_column_3_9, A0=>nx2988, A1=>nx2962, A2=>
      nx2934, A3=>nx2908);
   ix2989 : nand03 port map ( Y=>nx2988, A0=>nx7869, A1=>nx7871, A2=>nx7873
   );
   ix7870 : aoi222 port map ( Y=>nx7869, A0=>que_out_10_3_9, A1=>nx10304, B0
      =>que_out_6_3_9, B1=>nx10356, C0=>que_out_9_3_9, C1=>nx10330);
   ix7872 : aoi22 port map ( Y=>nx7871, A0=>que_out_5_3_9, A1=>nx10252, B0=>
      que_out_18_3_9, B1=>nx10278);
   ix7874 : aoi22 port map ( Y=>nx7873, A0=>que_out_17_3_9, A1=>nx10226, B0
      =>que_out_20_3_9, B1=>nx10200);
   ix2963 : nand03 port map ( Y=>nx2962, A0=>nx7877, A1=>nx7879, A2=>nx7881
   );
   ix7878 : aoi222 port map ( Y=>nx7877, A0=>que_out_19_3_9, A1=>nx10174, B0
      =>que_out_21_3_9, B1=>nx10148, C0=>que_out_8_3_9, C1=>nx10122);
   ix7880 : aoi22 port map ( Y=>nx7879, A0=>que_out_25_3_9, A1=>nx10070, B0
      =>que_out_16_3_9, B1=>nx10096);
   ix7882 : aoi22 port map ( Y=>nx7881, A0=>que_out_24_3_9, A1=>nx10044, B0
      =>que_out_22_3_9, B1=>nx10018);
   ix2935 : nand03 port map ( Y=>nx2934, A0=>nx7885, A1=>nx7887, A2=>nx7889
   );
   ix7886 : aoi222 port map ( Y=>nx7885, A0=>que_out_15_3_9, A1=>nx9966, B0
      =>que_out_3_3_9, B1=>nx9992, C0=>que_out_23_3_9, C1=>nx9940);
   ix7888 : aoi22 port map ( Y=>nx7887, A0=>que_out_27_3_9, A1=>nx9914, B0=>
      que_out_4_3_9, B1=>nx9888);
   ix7890 : aoi22 port map ( Y=>nx7889, A0=>que_out_0_3_9, A1=>nx9836, B0=>
      que_out_2_3_9, B1=>nx9862);
   ix2909 : nand03 port map ( Y=>nx2908, A0=>nx7893, A1=>nx7895, A2=>nx7897
   );
   ix7894 : aoi222 port map ( Y=>nx7893, A0=>que_out_26_3_9, A1=>nx9810, B0
      =>que_out_14_3_9, B1=>nx9784, C0=>que_out_11_3_9, C1=>nx9758);
   ix7896 : aoi22 port map ( Y=>nx7895, A0=>que_out_13_3_9, A1=>nx9732, B0=>
      que_out_7_3_9, B1=>nx9706);
   ix7898 : aoi22 port map ( Y=>nx7897, A0=>que_out_12_3_9, A1=>nx9680, B0=>
      que_out_1_3_9, B1=>nx9654);
   ix3103 : or04 port map ( Y=>out_column_3_10, A0=>nx3098, A1=>nx3072, A2=>
      nx3044, A3=>nx3018);
   ix3099 : nand03 port map ( Y=>nx3098, A0=>nx7903, A1=>nx7905, A2=>nx7907
   );
   ix7904 : aoi222 port map ( Y=>nx7903, A0=>que_out_10_3_10, A1=>nx10304, 
      B0=>que_out_6_3_10, B1=>nx10356, C0=>que_out_9_3_10, C1=>nx10330);
   ix7906 : aoi22 port map ( Y=>nx7905, A0=>que_out_5_3_10, A1=>nx10252, B0
      =>que_out_18_3_10, B1=>nx10278);
   ix7908 : aoi22 port map ( Y=>nx7907, A0=>que_out_17_3_10, A1=>nx10226, B0
      =>que_out_20_3_10, B1=>nx10200);
   ix3073 : nand03 port map ( Y=>nx3072, A0=>nx7911, A1=>nx7913, A2=>nx7915
   );
   ix7912 : aoi222 port map ( Y=>nx7911, A0=>que_out_19_3_10, A1=>nx10174, 
      B0=>que_out_21_3_10, B1=>nx10148, C0=>que_out_8_3_10, C1=>nx10122);
   ix7914 : aoi22 port map ( Y=>nx7913, A0=>que_out_25_3_10, A1=>nx10070, B0
      =>que_out_16_3_10, B1=>nx10096);
   ix7916 : aoi22 port map ( Y=>nx7915, A0=>que_out_24_3_10, A1=>nx10044, B0
      =>que_out_22_3_10, B1=>nx10018);
   ix3045 : nand03 port map ( Y=>nx3044, A0=>nx7919, A1=>nx7921, A2=>nx7923
   );
   ix7920 : aoi222 port map ( Y=>nx7919, A0=>que_out_15_3_10, A1=>nx9966, B0
      =>que_out_3_3_10, B1=>nx9992, C0=>que_out_23_3_10, C1=>nx9940);
   ix7922 : aoi22 port map ( Y=>nx7921, A0=>que_out_27_3_10, A1=>nx9914, B0
      =>que_out_4_3_10, B1=>nx9888);
   ix7924 : aoi22 port map ( Y=>nx7923, A0=>que_out_0_3_10, A1=>nx9836, B0=>
      que_out_2_3_10, B1=>nx9862);
   ix3019 : nand03 port map ( Y=>nx3018, A0=>nx7927, A1=>nx7929, A2=>nx7931
   );
   ix7928 : aoi222 port map ( Y=>nx7927, A0=>que_out_26_3_10, A1=>nx9810, B0
      =>que_out_14_3_10, B1=>nx9784, C0=>que_out_11_3_10, C1=>nx9758);
   ix7930 : aoi22 port map ( Y=>nx7929, A0=>que_out_13_3_10, A1=>nx9732, B0
      =>que_out_7_3_10, B1=>nx9706);
   ix7932 : aoi22 port map ( Y=>nx7931, A0=>que_out_12_3_10, A1=>nx9680, B0
      =>que_out_1_3_10, B1=>nx9654);
   ix3213 : or04 port map ( Y=>out_column_3_11, A0=>nx3208, A1=>nx3182, A2=>
      nx3154, A3=>nx3128);
   ix3209 : nand03 port map ( Y=>nx3208, A0=>nx7937, A1=>nx7939, A2=>nx7941
   );
   ix7938 : aoi222 port map ( Y=>nx7937, A0=>que_out_10_3_11, A1=>nx10304, 
      B0=>que_out_6_3_11, B1=>nx10356, C0=>que_out_9_3_11, C1=>nx10330);
   ix7940 : aoi22 port map ( Y=>nx7939, A0=>que_out_5_3_11, A1=>nx10252, B0
      =>que_out_18_3_11, B1=>nx10278);
   ix7942 : aoi22 port map ( Y=>nx7941, A0=>que_out_17_3_11, A1=>nx10226, B0
      =>que_out_20_3_11, B1=>nx10200);
   ix3183 : nand03 port map ( Y=>nx3182, A0=>nx7945, A1=>nx7947, A2=>nx7949
   );
   ix7946 : aoi222 port map ( Y=>nx7945, A0=>que_out_19_3_11, A1=>nx10174, 
      B0=>que_out_21_3_11, B1=>nx10148, C0=>que_out_8_3_11, C1=>nx10122);
   ix7948 : aoi22 port map ( Y=>nx7947, A0=>que_out_25_3_11, A1=>nx10070, B0
      =>que_out_16_3_11, B1=>nx10096);
   ix7950 : aoi22 port map ( Y=>nx7949, A0=>que_out_24_3_11, A1=>nx10044, B0
      =>que_out_22_3_11, B1=>nx10018);
   ix3155 : nand03 port map ( Y=>nx3154, A0=>nx7953, A1=>nx7955, A2=>nx7957
   );
   ix7954 : aoi222 port map ( Y=>nx7953, A0=>que_out_15_3_11, A1=>nx9966, B0
      =>que_out_3_3_11, B1=>nx9992, C0=>que_out_23_3_11, C1=>nx9940);
   ix7956 : aoi22 port map ( Y=>nx7955, A0=>que_out_27_3_11, A1=>nx9914, B0
      =>que_out_4_3_11, B1=>nx9888);
   ix7958 : aoi22 port map ( Y=>nx7957, A0=>que_out_0_3_11, A1=>nx9836, B0=>
      que_out_2_3_11, B1=>nx9862);
   ix3129 : nand03 port map ( Y=>nx3128, A0=>nx7961, A1=>nx7963, A2=>nx7965
   );
   ix7962 : aoi222 port map ( Y=>nx7961, A0=>que_out_26_3_11, A1=>nx9810, B0
      =>que_out_14_3_11, B1=>nx9784, C0=>que_out_11_3_11, C1=>nx9758);
   ix7964 : aoi22 port map ( Y=>nx7963, A0=>que_out_13_3_11, A1=>nx9732, B0
      =>que_out_7_3_11, B1=>nx9706);
   ix7966 : aoi22 port map ( Y=>nx7965, A0=>que_out_12_3_11, A1=>nx9680, B0
      =>que_out_1_3_11, B1=>nx9654);
   ix3323 : or04 port map ( Y=>out_column_3_12, A0=>nx3318, A1=>nx3292, A2=>
      nx3264, A3=>nx3238);
   ix3319 : nand03 port map ( Y=>nx3318, A0=>nx7971, A1=>nx7973, A2=>nx7975
   );
   ix7972 : aoi222 port map ( Y=>nx7971, A0=>que_out_10_3_12, A1=>nx10306, 
      B0=>que_out_6_3_12, B1=>nx10358, C0=>que_out_9_3_12, C1=>nx10332);
   ix7974 : aoi22 port map ( Y=>nx7973, A0=>que_out_5_3_12, A1=>nx10254, B0
      =>que_out_18_3_12, B1=>nx10280);
   ix7976 : aoi22 port map ( Y=>nx7975, A0=>que_out_17_3_12, A1=>nx10228, B0
      =>que_out_20_3_12, B1=>nx10202);
   ix3293 : nand03 port map ( Y=>nx3292, A0=>nx7979, A1=>nx7981, A2=>nx7983
   );
   ix7980 : aoi222 port map ( Y=>nx7979, A0=>que_out_19_3_12, A1=>nx10176, 
      B0=>que_out_21_3_12, B1=>nx10150, C0=>que_out_8_3_12, C1=>nx10124);
   ix7982 : aoi22 port map ( Y=>nx7981, A0=>que_out_25_3_12, A1=>nx10072, B0
      =>que_out_16_3_12, B1=>nx10098);
   ix7984 : aoi22 port map ( Y=>nx7983, A0=>que_out_24_3_12, A1=>nx10046, B0
      =>que_out_22_3_12, B1=>nx10020);
   ix3265 : nand03 port map ( Y=>nx3264, A0=>nx7987, A1=>nx7989, A2=>nx7991
   );
   ix7988 : aoi222 port map ( Y=>nx7987, A0=>que_out_15_3_12, A1=>nx9968, B0
      =>que_out_3_3_12, B1=>nx9994, C0=>que_out_23_3_12, C1=>nx9942);
   ix7990 : aoi22 port map ( Y=>nx7989, A0=>que_out_27_3_12, A1=>nx9916, B0
      =>que_out_4_3_12, B1=>nx9890);
   ix7992 : aoi22 port map ( Y=>nx7991, A0=>que_out_0_3_12, A1=>nx9838, B0=>
      que_out_2_3_12, B1=>nx9864);
   ix3239 : nand03 port map ( Y=>nx3238, A0=>nx7995, A1=>nx7997, A2=>nx7999
   );
   ix7996 : aoi222 port map ( Y=>nx7995, A0=>que_out_26_3_12, A1=>nx9812, B0
      =>que_out_14_3_12, B1=>nx9786, C0=>que_out_11_3_12, C1=>nx9760);
   ix7998 : aoi22 port map ( Y=>nx7997, A0=>que_out_13_3_12, A1=>nx9734, B0
      =>que_out_7_3_12, B1=>nx9708);
   ix8000 : aoi22 port map ( Y=>nx7999, A0=>que_out_12_3_12, A1=>nx9682, B0
      =>que_out_1_3_12, B1=>nx9656);
   ix3433 : or04 port map ( Y=>out_column_3_13, A0=>nx3428, A1=>nx3402, A2=>
      nx3374, A3=>nx3348);
   ix3429 : nand03 port map ( Y=>nx3428, A0=>nx8005, A1=>nx8007, A2=>nx8009
   );
   ix8006 : aoi222 port map ( Y=>nx8005, A0=>que_out_10_3_13, A1=>nx10306, 
      B0=>que_out_6_3_13, B1=>nx10358, C0=>que_out_9_3_13, C1=>nx10332);
   ix8008 : aoi22 port map ( Y=>nx8007, A0=>que_out_5_3_13, A1=>nx10254, B0
      =>que_out_18_3_13, B1=>nx10280);
   ix8010 : aoi22 port map ( Y=>nx8009, A0=>que_out_17_3_13, A1=>nx10228, B0
      =>que_out_20_3_13, B1=>nx10202);
   ix3403 : nand03 port map ( Y=>nx3402, A0=>nx8013, A1=>nx8015, A2=>nx8017
   );
   ix8014 : aoi222 port map ( Y=>nx8013, A0=>que_out_19_3_13, A1=>nx10176, 
      B0=>que_out_21_3_13, B1=>nx10150, C0=>que_out_8_3_13, C1=>nx10124);
   ix8016 : aoi22 port map ( Y=>nx8015, A0=>que_out_25_3_13, A1=>nx10072, B0
      =>que_out_16_3_13, B1=>nx10098);
   ix8018 : aoi22 port map ( Y=>nx8017, A0=>que_out_24_3_13, A1=>nx10046, B0
      =>que_out_22_3_13, B1=>nx10020);
   ix3375 : nand03 port map ( Y=>nx3374, A0=>nx8021, A1=>nx8023, A2=>nx8025
   );
   ix8022 : aoi222 port map ( Y=>nx8021, A0=>que_out_15_3_13, A1=>nx9968, B0
      =>que_out_3_3_13, B1=>nx9994, C0=>que_out_23_3_13, C1=>nx9942);
   ix8024 : aoi22 port map ( Y=>nx8023, A0=>que_out_27_3_13, A1=>nx9916, B0
      =>que_out_4_3_13, B1=>nx9890);
   ix8026 : aoi22 port map ( Y=>nx8025, A0=>que_out_0_3_13, A1=>nx9838, B0=>
      que_out_2_3_13, B1=>nx9864);
   ix3349 : nand03 port map ( Y=>nx3348, A0=>nx8029, A1=>nx8031, A2=>nx8033
   );
   ix8030 : aoi222 port map ( Y=>nx8029, A0=>que_out_26_3_13, A1=>nx9812, B0
      =>que_out_14_3_13, B1=>nx9786, C0=>que_out_11_3_13, C1=>nx9760);
   ix8032 : aoi22 port map ( Y=>nx8031, A0=>que_out_13_3_13, A1=>nx9734, B0
      =>que_out_7_3_13, B1=>nx9708);
   ix8034 : aoi22 port map ( Y=>nx8033, A0=>que_out_12_3_13, A1=>nx9682, B0
      =>que_out_1_3_13, B1=>nx9656);
   ix3543 : or04 port map ( Y=>out_column_3_14, A0=>nx3538, A1=>nx3512, A2=>
      nx3484, A3=>nx3458);
   ix3539 : nand03 port map ( Y=>nx3538, A0=>nx8039, A1=>nx8041, A2=>nx8043
   );
   ix8040 : aoi222 port map ( Y=>nx8039, A0=>que_out_10_3_14, A1=>nx10306, 
      B0=>que_out_6_3_14, B1=>nx10358, C0=>que_out_9_3_14, C1=>nx10332);
   ix8042 : aoi22 port map ( Y=>nx8041, A0=>que_out_5_3_14, A1=>nx10254, B0
      =>que_out_18_3_14, B1=>nx10280);
   ix8044 : aoi22 port map ( Y=>nx8043, A0=>que_out_17_3_14, A1=>nx10228, B0
      =>que_out_20_3_14, B1=>nx10202);
   ix3513 : nand03 port map ( Y=>nx3512, A0=>nx8047, A1=>nx8049, A2=>nx8051
   );
   ix8048 : aoi222 port map ( Y=>nx8047, A0=>que_out_19_3_14, A1=>nx10176, 
      B0=>que_out_21_3_14, B1=>nx10150, C0=>que_out_8_3_14, C1=>nx10124);
   ix8050 : aoi22 port map ( Y=>nx8049, A0=>que_out_25_3_14, A1=>nx10072, B0
      =>que_out_16_3_14, B1=>nx10098);
   ix8052 : aoi22 port map ( Y=>nx8051, A0=>que_out_24_3_14, A1=>nx10046, B0
      =>que_out_22_3_14, B1=>nx10020);
   ix3485 : nand03 port map ( Y=>nx3484, A0=>nx8055, A1=>nx8057, A2=>nx8059
   );
   ix8056 : aoi222 port map ( Y=>nx8055, A0=>que_out_15_3_14, A1=>nx9968, B0
      =>que_out_3_3_14, B1=>nx9994, C0=>que_out_23_3_14, C1=>nx9942);
   ix8058 : aoi22 port map ( Y=>nx8057, A0=>que_out_27_3_14, A1=>nx9916, B0
      =>que_out_4_3_14, B1=>nx9890);
   ix8060 : aoi22 port map ( Y=>nx8059, A0=>que_out_0_3_14, A1=>nx9838, B0=>
      que_out_2_3_14, B1=>nx9864);
   ix3459 : nand03 port map ( Y=>nx3458, A0=>nx8063, A1=>nx8065, A2=>nx8067
   );
   ix8064 : aoi222 port map ( Y=>nx8063, A0=>que_out_26_3_14, A1=>nx9812, B0
      =>que_out_14_3_14, B1=>nx9786, C0=>que_out_11_3_14, C1=>nx9760);
   ix8066 : aoi22 port map ( Y=>nx8065, A0=>que_out_13_3_14, A1=>nx9734, B0
      =>que_out_7_3_14, B1=>nx9708);
   ix8068 : aoi22 port map ( Y=>nx8067, A0=>que_out_12_3_14, A1=>nx9682, B0
      =>que_out_1_3_14, B1=>nx9656);
   ix3653 : or04 port map ( Y=>out_column_3_15, A0=>nx3648, A1=>nx3622, A2=>
      nx3594, A3=>nx3568);
   ix3649 : nand03 port map ( Y=>nx3648, A0=>nx8073, A1=>nx8075, A2=>nx8077
   );
   ix8074 : aoi222 port map ( Y=>nx8073, A0=>que_out_10_3_15, A1=>nx10306, 
      B0=>que_out_6_3_15, B1=>nx10358, C0=>que_out_9_3_15, C1=>nx10332);
   ix8076 : aoi22 port map ( Y=>nx8075, A0=>que_out_5_3_15, A1=>nx10254, B0
      =>que_out_18_3_15, B1=>nx10280);
   ix8078 : aoi22 port map ( Y=>nx8077, A0=>que_out_17_3_15, A1=>nx10228, B0
      =>que_out_20_3_15, B1=>nx10202);
   ix3623 : nand03 port map ( Y=>nx3622, A0=>nx8081, A1=>nx8083, A2=>nx8085
   );
   ix8082 : aoi222 port map ( Y=>nx8081, A0=>que_out_19_3_15, A1=>nx10176, 
      B0=>que_out_21_3_15, B1=>nx10150, C0=>que_out_8_3_15, C1=>nx10124);
   ix8084 : aoi22 port map ( Y=>nx8083, A0=>que_out_25_3_15, A1=>nx10072, B0
      =>que_out_16_3_15, B1=>nx10098);
   ix8086 : aoi22 port map ( Y=>nx8085, A0=>que_out_24_3_15, A1=>nx10046, B0
      =>que_out_22_3_15, B1=>nx10020);
   ix3595 : nand03 port map ( Y=>nx3594, A0=>nx8089, A1=>nx8091, A2=>nx8093
   );
   ix8090 : aoi222 port map ( Y=>nx8089, A0=>que_out_15_3_15, A1=>nx9968, B0
      =>que_out_3_3_15, B1=>nx9994, C0=>que_out_23_3_15, C1=>nx9942);
   ix8092 : aoi22 port map ( Y=>nx8091, A0=>que_out_27_3_15, A1=>nx9916, B0
      =>que_out_4_3_15, B1=>nx9890);
   ix8094 : aoi22 port map ( Y=>nx8093, A0=>que_out_0_3_15, A1=>nx9838, B0=>
      que_out_2_3_15, B1=>nx9864);
   ix3569 : nand03 port map ( Y=>nx3568, A0=>nx8097, A1=>nx8099, A2=>nx8101
   );
   ix8098 : aoi222 port map ( Y=>nx8097, A0=>que_out_26_3_15, A1=>nx9812, B0
      =>que_out_14_3_15, B1=>nx9786, C0=>que_out_11_3_15, C1=>nx9760);
   ix8100 : aoi22 port map ( Y=>nx8099, A0=>que_out_13_3_15, A1=>nx9734, B0
      =>que_out_7_3_15, B1=>nx9708);
   ix8102 : aoi22 port map ( Y=>nx8101, A0=>que_out_12_3_15, A1=>nx9682, B0
      =>que_out_1_3_15, B1=>nx9656);
   ix3763 : or04 port map ( Y=>out_column_2_0, A0=>nx3758, A1=>nx3732, A2=>
      nx3704, A3=>nx3678);
   ix3759 : nand03 port map ( Y=>nx3758, A0=>nx8107, A1=>nx8109, A2=>nx8111
   );
   ix8108 : aoi222 port map ( Y=>nx8107, A0=>que_out_10_2_0, A1=>nx10306, B0
      =>que_out_6_2_0, B1=>nx10358, C0=>que_out_9_2_0, C1=>nx10332);
   ix8110 : aoi22 port map ( Y=>nx8109, A0=>que_out_5_2_0, A1=>nx10254, B0=>
      que_out_18_2_0, B1=>nx10280);
   ix8112 : aoi22 port map ( Y=>nx8111, A0=>que_out_17_2_0, A1=>nx10228, B0
      =>que_out_20_2_0, B1=>nx10202);
   ix3733 : nand03 port map ( Y=>nx3732, A0=>nx8115, A1=>nx8117, A2=>nx8119
   );
   ix8116 : aoi222 port map ( Y=>nx8115, A0=>que_out_19_2_0, A1=>nx10176, B0
      =>que_out_21_2_0, B1=>nx10150, C0=>que_out_8_2_0, C1=>nx10124);
   ix8118 : aoi22 port map ( Y=>nx8117, A0=>que_out_25_2_0, A1=>nx10072, B0
      =>que_out_16_2_0, B1=>nx10098);
   ix8120 : aoi22 port map ( Y=>nx8119, A0=>que_out_24_2_0, A1=>nx10046, B0
      =>que_out_22_2_0, B1=>nx10020);
   ix3705 : nand03 port map ( Y=>nx3704, A0=>nx8123, A1=>nx8125, A2=>nx8127
   );
   ix8124 : aoi222 port map ( Y=>nx8123, A0=>que_out_15_2_0, A1=>nx9968, B0
      =>que_out_3_2_0, B1=>nx9994, C0=>que_out_23_2_0, C1=>nx9942);
   ix8126 : aoi22 port map ( Y=>nx8125, A0=>que_out_27_2_0, A1=>nx9916, B0=>
      que_out_4_2_0, B1=>nx9890);
   ix8128 : aoi22 port map ( Y=>nx8127, A0=>que_out_0_2_0, A1=>nx9838, B0=>
      que_out_2_2_0, B1=>nx9864);
   ix3679 : nand03 port map ( Y=>nx3678, A0=>nx8131, A1=>nx8133, A2=>nx8135
   );
   ix8132 : aoi222 port map ( Y=>nx8131, A0=>que_out_26_2_0, A1=>nx9812, B0
      =>que_out_14_2_0, B1=>nx9786, C0=>que_out_11_2_0, C1=>nx9760);
   ix8134 : aoi22 port map ( Y=>nx8133, A0=>que_out_13_2_0, A1=>nx9734, B0=>
      que_out_7_2_0, B1=>nx9708);
   ix8136 : aoi22 port map ( Y=>nx8135, A0=>que_out_12_2_0, A1=>nx9682, B0=>
      que_out_1_2_0, B1=>nx9656);
   ix3873 : or04 port map ( Y=>out_column_2_1, A0=>nx3868, A1=>nx3842, A2=>
      nx3814, A3=>nx3788);
   ix3869 : nand03 port map ( Y=>nx3868, A0=>nx8141, A1=>nx8143, A2=>nx8145
   );
   ix8142 : aoi222 port map ( Y=>nx8141, A0=>que_out_10_2_1, A1=>nx10306, B0
      =>que_out_6_2_1, B1=>nx10358, C0=>que_out_9_2_1, C1=>nx10332);
   ix8144 : aoi22 port map ( Y=>nx8143, A0=>que_out_5_2_1, A1=>nx10254, B0=>
      que_out_18_2_1, B1=>nx10280);
   ix8146 : aoi22 port map ( Y=>nx8145, A0=>que_out_17_2_1, A1=>nx10228, B0
      =>que_out_20_2_1, B1=>nx10202);
   ix3843 : nand03 port map ( Y=>nx3842, A0=>nx8149, A1=>nx8151, A2=>nx8153
   );
   ix8150 : aoi222 port map ( Y=>nx8149, A0=>que_out_19_2_1, A1=>nx10176, B0
      =>que_out_21_2_1, B1=>nx10150, C0=>que_out_8_2_1, C1=>nx10124);
   ix8152 : aoi22 port map ( Y=>nx8151, A0=>que_out_25_2_1, A1=>nx10072, B0
      =>que_out_16_2_1, B1=>nx10098);
   ix8154 : aoi22 port map ( Y=>nx8153, A0=>que_out_24_2_1, A1=>nx10046, B0
      =>que_out_22_2_1, B1=>nx10020);
   ix3815 : nand03 port map ( Y=>nx3814, A0=>nx8157, A1=>nx8159, A2=>nx8161
   );
   ix8158 : aoi222 port map ( Y=>nx8157, A0=>que_out_15_2_1, A1=>nx9968, B0
      =>que_out_3_2_1, B1=>nx9994, C0=>que_out_23_2_1, C1=>nx9942);
   ix8160 : aoi22 port map ( Y=>nx8159, A0=>que_out_27_2_1, A1=>nx9916, B0=>
      que_out_4_2_1, B1=>nx9890);
   ix8162 : aoi22 port map ( Y=>nx8161, A0=>que_out_0_2_1, A1=>nx9838, B0=>
      que_out_2_2_1, B1=>nx9864);
   ix3789 : nand03 port map ( Y=>nx3788, A0=>nx8165, A1=>nx8167, A2=>nx8169
   );
   ix8166 : aoi222 port map ( Y=>nx8165, A0=>que_out_26_2_1, A1=>nx9812, B0
      =>que_out_14_2_1, B1=>nx9786, C0=>que_out_11_2_1, C1=>nx9760);
   ix8168 : aoi22 port map ( Y=>nx8167, A0=>que_out_13_2_1, A1=>nx9734, B0=>
      que_out_7_2_1, B1=>nx9708);
   ix8170 : aoi22 port map ( Y=>nx8169, A0=>que_out_12_2_1, A1=>nx9682, B0=>
      que_out_1_2_1, B1=>nx9656);
   ix3983 : or04 port map ( Y=>out_column_2_2, A0=>nx3978, A1=>nx3952, A2=>
      nx3924, A3=>nx3898);
   ix3979 : nand03 port map ( Y=>nx3978, A0=>nx8175, A1=>nx8177, A2=>nx8179
   );
   ix8176 : aoi222 port map ( Y=>nx8175, A0=>que_out_10_2_2, A1=>nx10306, B0
      =>que_out_6_2_2, B1=>nx10358, C0=>que_out_9_2_2, C1=>nx10332);
   ix8178 : aoi22 port map ( Y=>nx8177, A0=>que_out_5_2_2, A1=>nx10254, B0=>
      que_out_18_2_2, B1=>nx10280);
   ix8180 : aoi22 port map ( Y=>nx8179, A0=>que_out_17_2_2, A1=>nx10228, B0
      =>que_out_20_2_2, B1=>nx10202);
   ix3953 : nand03 port map ( Y=>nx3952, A0=>nx8183, A1=>nx8185, A2=>nx8187
   );
   ix8184 : aoi222 port map ( Y=>nx8183, A0=>que_out_19_2_2, A1=>nx10176, B0
      =>que_out_21_2_2, B1=>nx10150, C0=>que_out_8_2_2, C1=>nx10124);
   ix8186 : aoi22 port map ( Y=>nx8185, A0=>que_out_25_2_2, A1=>nx10072, B0
      =>que_out_16_2_2, B1=>nx10098);
   ix8188 : aoi22 port map ( Y=>nx8187, A0=>que_out_24_2_2, A1=>nx10046, B0
      =>que_out_22_2_2, B1=>nx10020);
   ix3925 : nand03 port map ( Y=>nx3924, A0=>nx8191, A1=>nx8193, A2=>nx8195
   );
   ix8192 : aoi222 port map ( Y=>nx8191, A0=>que_out_15_2_2, A1=>nx9968, B0
      =>que_out_3_2_2, B1=>nx9994, C0=>que_out_23_2_2, C1=>nx9942);
   ix8194 : aoi22 port map ( Y=>nx8193, A0=>que_out_27_2_2, A1=>nx9916, B0=>
      que_out_4_2_2, B1=>nx9890);
   ix8196 : aoi22 port map ( Y=>nx8195, A0=>que_out_0_2_2, A1=>nx9838, B0=>
      que_out_2_2_2, B1=>nx9864);
   ix3899 : nand03 port map ( Y=>nx3898, A0=>nx8199, A1=>nx8201, A2=>nx8203
   );
   ix8200 : aoi222 port map ( Y=>nx8199, A0=>que_out_26_2_2, A1=>nx9812, B0
      =>que_out_14_2_2, B1=>nx9786, C0=>que_out_11_2_2, C1=>nx9760);
   ix8202 : aoi22 port map ( Y=>nx8201, A0=>que_out_13_2_2, A1=>nx9734, B0=>
      que_out_7_2_2, B1=>nx9708);
   ix8204 : aoi22 port map ( Y=>nx8203, A0=>que_out_12_2_2, A1=>nx9682, B0=>
      que_out_1_2_2, B1=>nx9656);
   ix4093 : or04 port map ( Y=>out_column_2_3, A0=>nx4088, A1=>nx4062, A2=>
      nx4034, A3=>nx4008);
   ix4089 : nand03 port map ( Y=>nx4088, A0=>nx8209, A1=>nx8211, A2=>nx8213
   );
   ix8210 : aoi222 port map ( Y=>nx8209, A0=>que_out_10_2_3, A1=>nx10308, B0
      =>que_out_6_2_3, B1=>nx10360, C0=>que_out_9_2_3, C1=>nx10334);
   ix8212 : aoi22 port map ( Y=>nx8211, A0=>que_out_5_2_3, A1=>nx10256, B0=>
      que_out_18_2_3, B1=>nx10282);
   ix8214 : aoi22 port map ( Y=>nx8213, A0=>que_out_17_2_3, A1=>nx10230, B0
      =>que_out_20_2_3, B1=>nx10204);
   ix4063 : nand03 port map ( Y=>nx4062, A0=>nx8217, A1=>nx8219, A2=>nx8221
   );
   ix8218 : aoi222 port map ( Y=>nx8217, A0=>que_out_19_2_3, A1=>nx10178, B0
      =>que_out_21_2_3, B1=>nx10152, C0=>que_out_8_2_3, C1=>nx10126);
   ix8220 : aoi22 port map ( Y=>nx8219, A0=>que_out_25_2_3, A1=>nx10074, B0
      =>que_out_16_2_3, B1=>nx10100);
   ix8222 : aoi22 port map ( Y=>nx8221, A0=>que_out_24_2_3, A1=>nx10048, B0
      =>que_out_22_2_3, B1=>nx10022);
   ix4035 : nand03 port map ( Y=>nx4034, A0=>nx8225, A1=>nx8227, A2=>nx8229
   );
   ix8226 : aoi222 port map ( Y=>nx8225, A0=>que_out_15_2_3, A1=>nx9970, B0
      =>que_out_3_2_3, B1=>nx9996, C0=>que_out_23_2_3, C1=>nx9944);
   ix8228 : aoi22 port map ( Y=>nx8227, A0=>que_out_27_2_3, A1=>nx9918, B0=>
      que_out_4_2_3, B1=>nx9892);
   ix8230 : aoi22 port map ( Y=>nx8229, A0=>que_out_0_2_3, A1=>nx9840, B0=>
      que_out_2_2_3, B1=>nx9866);
   ix4009 : nand03 port map ( Y=>nx4008, A0=>nx8233, A1=>nx8235, A2=>nx8237
   );
   ix8234 : aoi222 port map ( Y=>nx8233, A0=>que_out_26_2_3, A1=>nx9814, B0
      =>que_out_14_2_3, B1=>nx9788, C0=>que_out_11_2_3, C1=>nx9762);
   ix8236 : aoi22 port map ( Y=>nx8235, A0=>que_out_13_2_3, A1=>nx9736, B0=>
      que_out_7_2_3, B1=>nx9710);
   ix8238 : aoi22 port map ( Y=>nx8237, A0=>que_out_12_2_3, A1=>nx9684, B0=>
      que_out_1_2_3, B1=>nx9658);
   ix4203 : or04 port map ( Y=>out_column_2_4, A0=>nx4198, A1=>nx4172, A2=>
      nx4144, A3=>nx4118);
   ix4199 : nand03 port map ( Y=>nx4198, A0=>nx8243, A1=>nx8245, A2=>nx8247
   );
   ix8244 : aoi222 port map ( Y=>nx8243, A0=>que_out_10_2_4, A1=>nx10308, B0
      =>que_out_6_2_4, B1=>nx10360, C0=>que_out_9_2_4, C1=>nx10334);
   ix8246 : aoi22 port map ( Y=>nx8245, A0=>que_out_5_2_4, A1=>nx10256, B0=>
      que_out_18_2_4, B1=>nx10282);
   ix8248 : aoi22 port map ( Y=>nx8247, A0=>que_out_17_2_4, A1=>nx10230, B0
      =>que_out_20_2_4, B1=>nx10204);
   ix4173 : nand03 port map ( Y=>nx4172, A0=>nx8251, A1=>nx8253, A2=>nx8255
   );
   ix8252 : aoi222 port map ( Y=>nx8251, A0=>que_out_19_2_4, A1=>nx10178, B0
      =>que_out_21_2_4, B1=>nx10152, C0=>que_out_8_2_4, C1=>nx10126);
   ix8254 : aoi22 port map ( Y=>nx8253, A0=>que_out_25_2_4, A1=>nx10074, B0
      =>que_out_16_2_4, B1=>nx10100);
   ix8256 : aoi22 port map ( Y=>nx8255, A0=>que_out_24_2_4, A1=>nx10048, B0
      =>que_out_22_2_4, B1=>nx10022);
   ix4145 : nand03 port map ( Y=>nx4144, A0=>nx8259, A1=>nx8261, A2=>nx8263
   );
   ix8260 : aoi222 port map ( Y=>nx8259, A0=>que_out_15_2_4, A1=>nx9970, B0
      =>que_out_3_2_4, B1=>nx9996, C0=>que_out_23_2_4, C1=>nx9944);
   ix8262 : aoi22 port map ( Y=>nx8261, A0=>que_out_27_2_4, A1=>nx9918, B0=>
      que_out_4_2_4, B1=>nx9892);
   ix8264 : aoi22 port map ( Y=>nx8263, A0=>que_out_0_2_4, A1=>nx9840, B0=>
      que_out_2_2_4, B1=>nx9866);
   ix4119 : nand03 port map ( Y=>nx4118, A0=>nx8267, A1=>nx8269, A2=>nx8271
   );
   ix8268 : aoi222 port map ( Y=>nx8267, A0=>que_out_26_2_4, A1=>nx9814, B0
      =>que_out_14_2_4, B1=>nx9788, C0=>que_out_11_2_4, C1=>nx9762);
   ix8270 : aoi22 port map ( Y=>nx8269, A0=>que_out_13_2_4, A1=>nx9736, B0=>
      que_out_7_2_4, B1=>nx9710);
   ix8272 : aoi22 port map ( Y=>nx8271, A0=>que_out_12_2_4, A1=>nx9684, B0=>
      que_out_1_2_4, B1=>nx9658);
   ix4313 : or04 port map ( Y=>out_column_2_5, A0=>nx4308, A1=>nx4282, A2=>
      nx4254, A3=>nx4228);
   ix4309 : nand03 port map ( Y=>nx4308, A0=>nx8277, A1=>nx8279, A2=>nx8281
   );
   ix8278 : aoi222 port map ( Y=>nx8277, A0=>que_out_10_2_5, A1=>nx10308, B0
      =>que_out_6_2_5, B1=>nx10360, C0=>que_out_9_2_5, C1=>nx10334);
   ix8280 : aoi22 port map ( Y=>nx8279, A0=>que_out_5_2_5, A1=>nx10256, B0=>
      que_out_18_2_5, B1=>nx10282);
   ix8282 : aoi22 port map ( Y=>nx8281, A0=>que_out_17_2_5, A1=>nx10230, B0
      =>que_out_20_2_5, B1=>nx10204);
   ix4283 : nand03 port map ( Y=>nx4282, A0=>nx8285, A1=>nx8287, A2=>nx8289
   );
   ix8286 : aoi222 port map ( Y=>nx8285, A0=>que_out_19_2_5, A1=>nx10178, B0
      =>que_out_21_2_5, B1=>nx10152, C0=>que_out_8_2_5, C1=>nx10126);
   ix8288 : aoi22 port map ( Y=>nx8287, A0=>que_out_25_2_5, A1=>nx10074, B0
      =>que_out_16_2_5, B1=>nx10100);
   ix8290 : aoi22 port map ( Y=>nx8289, A0=>que_out_24_2_5, A1=>nx10048, B0
      =>que_out_22_2_5, B1=>nx10022);
   ix4255 : nand03 port map ( Y=>nx4254, A0=>nx8293, A1=>nx8295, A2=>nx8297
   );
   ix8294 : aoi222 port map ( Y=>nx8293, A0=>que_out_15_2_5, A1=>nx9970, B0
      =>que_out_3_2_5, B1=>nx9996, C0=>que_out_23_2_5, C1=>nx9944);
   ix8296 : aoi22 port map ( Y=>nx8295, A0=>que_out_27_2_5, A1=>nx9918, B0=>
      que_out_4_2_5, B1=>nx9892);
   ix8298 : aoi22 port map ( Y=>nx8297, A0=>que_out_0_2_5, A1=>nx9840, B0=>
      que_out_2_2_5, B1=>nx9866);
   ix4229 : nand03 port map ( Y=>nx4228, A0=>nx8301, A1=>nx8303, A2=>nx8305
   );
   ix8302 : aoi222 port map ( Y=>nx8301, A0=>que_out_26_2_5, A1=>nx9814, B0
      =>que_out_14_2_5, B1=>nx9788, C0=>que_out_11_2_5, C1=>nx9762);
   ix8304 : aoi22 port map ( Y=>nx8303, A0=>que_out_13_2_5, A1=>nx9736, B0=>
      que_out_7_2_5, B1=>nx9710);
   ix8306 : aoi22 port map ( Y=>nx8305, A0=>que_out_12_2_5, A1=>nx9684, B0=>
      que_out_1_2_5, B1=>nx9658);
   ix4423 : or04 port map ( Y=>out_column_2_6, A0=>nx4418, A1=>nx4392, A2=>
      nx4364, A3=>nx4338);
   ix4419 : nand03 port map ( Y=>nx4418, A0=>nx8311, A1=>nx8313, A2=>nx8315
   );
   ix8312 : aoi222 port map ( Y=>nx8311, A0=>que_out_10_2_6, A1=>nx10308, B0
      =>que_out_6_2_6, B1=>nx10360, C0=>que_out_9_2_6, C1=>nx10334);
   ix8314 : aoi22 port map ( Y=>nx8313, A0=>que_out_5_2_6, A1=>nx10256, B0=>
      que_out_18_2_6, B1=>nx10282);
   ix8316 : aoi22 port map ( Y=>nx8315, A0=>que_out_17_2_6, A1=>nx10230, B0
      =>que_out_20_2_6, B1=>nx10204);
   ix4393 : nand03 port map ( Y=>nx4392, A0=>nx8319, A1=>nx8321, A2=>nx8323
   );
   ix8320 : aoi222 port map ( Y=>nx8319, A0=>que_out_19_2_6, A1=>nx10178, B0
      =>que_out_21_2_6, B1=>nx10152, C0=>que_out_8_2_6, C1=>nx10126);
   ix8322 : aoi22 port map ( Y=>nx8321, A0=>que_out_25_2_6, A1=>nx10074, B0
      =>que_out_16_2_6, B1=>nx10100);
   ix8324 : aoi22 port map ( Y=>nx8323, A0=>que_out_24_2_6, A1=>nx10048, B0
      =>que_out_22_2_6, B1=>nx10022);
   ix4365 : nand03 port map ( Y=>nx4364, A0=>nx8327, A1=>nx8329, A2=>nx8331
   );
   ix8328 : aoi222 port map ( Y=>nx8327, A0=>que_out_15_2_6, A1=>nx9970, B0
      =>que_out_3_2_6, B1=>nx9996, C0=>que_out_23_2_6, C1=>nx9944);
   ix8330 : aoi22 port map ( Y=>nx8329, A0=>que_out_27_2_6, A1=>nx9918, B0=>
      que_out_4_2_6, B1=>nx9892);
   ix8332 : aoi22 port map ( Y=>nx8331, A0=>que_out_0_2_6, A1=>nx9840, B0=>
      que_out_2_2_6, B1=>nx9866);
   ix4339 : nand03 port map ( Y=>nx4338, A0=>nx8335, A1=>nx8337, A2=>nx8339
   );
   ix8336 : aoi222 port map ( Y=>nx8335, A0=>que_out_26_2_6, A1=>nx9814, B0
      =>que_out_14_2_6, B1=>nx9788, C0=>que_out_11_2_6, C1=>nx9762);
   ix8338 : aoi22 port map ( Y=>nx8337, A0=>que_out_13_2_6, A1=>nx9736, B0=>
      que_out_7_2_6, B1=>nx9710);
   ix8340 : aoi22 port map ( Y=>nx8339, A0=>que_out_12_2_6, A1=>nx9684, B0=>
      que_out_1_2_6, B1=>nx9658);
   ix4533 : or04 port map ( Y=>out_column_2_7, A0=>nx4528, A1=>nx4502, A2=>
      nx4474, A3=>nx4448);
   ix4529 : nand03 port map ( Y=>nx4528, A0=>nx8345, A1=>nx8347, A2=>nx8349
   );
   ix8346 : aoi222 port map ( Y=>nx8345, A0=>que_out_10_2_7, A1=>nx10308, B0
      =>que_out_6_2_7, B1=>nx10360, C0=>que_out_9_2_7, C1=>nx10334);
   ix8348 : aoi22 port map ( Y=>nx8347, A0=>que_out_5_2_7, A1=>nx10256, B0=>
      que_out_18_2_7, B1=>nx10282);
   ix8350 : aoi22 port map ( Y=>nx8349, A0=>que_out_17_2_7, A1=>nx10230, B0
      =>que_out_20_2_7, B1=>nx10204);
   ix4503 : nand03 port map ( Y=>nx4502, A0=>nx8353, A1=>nx8355, A2=>nx8357
   );
   ix8354 : aoi222 port map ( Y=>nx8353, A0=>que_out_19_2_7, A1=>nx10178, B0
      =>que_out_21_2_7, B1=>nx10152, C0=>que_out_8_2_7, C1=>nx10126);
   ix8356 : aoi22 port map ( Y=>nx8355, A0=>que_out_25_2_7, A1=>nx10074, B0
      =>que_out_16_2_7, B1=>nx10100);
   ix8358 : aoi22 port map ( Y=>nx8357, A0=>que_out_24_2_7, A1=>nx10048, B0
      =>que_out_22_2_7, B1=>nx10022);
   ix4475 : nand03 port map ( Y=>nx4474, A0=>nx8361, A1=>nx8363, A2=>nx8365
   );
   ix8362 : aoi222 port map ( Y=>nx8361, A0=>que_out_15_2_7, A1=>nx9970, B0
      =>que_out_3_2_7, B1=>nx9996, C0=>que_out_23_2_7, C1=>nx9944);
   ix8364 : aoi22 port map ( Y=>nx8363, A0=>que_out_27_2_7, A1=>nx9918, B0=>
      que_out_4_2_7, B1=>nx9892);
   ix8366 : aoi22 port map ( Y=>nx8365, A0=>que_out_0_2_7, A1=>nx9840, B0=>
      que_out_2_2_7, B1=>nx9866);
   ix4449 : nand03 port map ( Y=>nx4448, A0=>nx8369, A1=>nx8371, A2=>nx8373
   );
   ix8370 : aoi222 port map ( Y=>nx8369, A0=>que_out_26_2_7, A1=>nx9814, B0
      =>que_out_14_2_7, B1=>nx9788, C0=>que_out_11_2_7, C1=>nx9762);
   ix8372 : aoi22 port map ( Y=>nx8371, A0=>que_out_13_2_7, A1=>nx9736, B0=>
      que_out_7_2_7, B1=>nx9710);
   ix8374 : aoi22 port map ( Y=>nx8373, A0=>que_out_12_2_7, A1=>nx9684, B0=>
      que_out_1_2_7, B1=>nx9658);
   ix4643 : or04 port map ( Y=>out_column_2_8, A0=>nx4638, A1=>nx4612, A2=>
      nx4584, A3=>nx4558);
   ix4639 : nand03 port map ( Y=>nx4638, A0=>nx8379, A1=>nx8381, A2=>nx8383
   );
   ix8380 : aoi222 port map ( Y=>nx8379, A0=>que_out_10_2_8, A1=>nx10308, B0
      =>que_out_6_2_8, B1=>nx10360, C0=>que_out_9_2_8, C1=>nx10334);
   ix8382 : aoi22 port map ( Y=>nx8381, A0=>que_out_5_2_8, A1=>nx10256, B0=>
      que_out_18_2_8, B1=>nx10282);
   ix8384 : aoi22 port map ( Y=>nx8383, A0=>que_out_17_2_8, A1=>nx10230, B0
      =>que_out_20_2_8, B1=>nx10204);
   ix4613 : nand03 port map ( Y=>nx4612, A0=>nx8387, A1=>nx8389, A2=>nx8391
   );
   ix8388 : aoi222 port map ( Y=>nx8387, A0=>que_out_19_2_8, A1=>nx10178, B0
      =>que_out_21_2_8, B1=>nx10152, C0=>que_out_8_2_8, C1=>nx10126);
   ix8390 : aoi22 port map ( Y=>nx8389, A0=>que_out_25_2_8, A1=>nx10074, B0
      =>que_out_16_2_8, B1=>nx10100);
   ix8392 : aoi22 port map ( Y=>nx8391, A0=>que_out_24_2_8, A1=>nx10048, B0
      =>que_out_22_2_8, B1=>nx10022);
   ix4585 : nand03 port map ( Y=>nx4584, A0=>nx8395, A1=>nx8397, A2=>nx8399
   );
   ix8396 : aoi222 port map ( Y=>nx8395, A0=>que_out_15_2_8, A1=>nx9970, B0
      =>que_out_3_2_8, B1=>nx9996, C0=>que_out_23_2_8, C1=>nx9944);
   ix8398 : aoi22 port map ( Y=>nx8397, A0=>que_out_27_2_8, A1=>nx9918, B0=>
      que_out_4_2_8, B1=>nx9892);
   ix8400 : aoi22 port map ( Y=>nx8399, A0=>que_out_0_2_8, A1=>nx9840, B0=>
      que_out_2_2_8, B1=>nx9866);
   ix4559 : nand03 port map ( Y=>nx4558, A0=>nx8403, A1=>nx8405, A2=>nx8407
   );
   ix8404 : aoi222 port map ( Y=>nx8403, A0=>que_out_26_2_8, A1=>nx9814, B0
      =>que_out_14_2_8, B1=>nx9788, C0=>que_out_11_2_8, C1=>nx9762);
   ix8406 : aoi22 port map ( Y=>nx8405, A0=>que_out_13_2_8, A1=>nx9736, B0=>
      que_out_7_2_8, B1=>nx9710);
   ix8408 : aoi22 port map ( Y=>nx8407, A0=>que_out_12_2_8, A1=>nx9684, B0=>
      que_out_1_2_8, B1=>nx9658);
   ix4753 : or04 port map ( Y=>out_column_2_9, A0=>nx4748, A1=>nx4722, A2=>
      nx4694, A3=>nx4668);
   ix4749 : nand03 port map ( Y=>nx4748, A0=>nx8413, A1=>nx8415, A2=>nx8417
   );
   ix8414 : aoi222 port map ( Y=>nx8413, A0=>que_out_10_2_9, A1=>nx10308, B0
      =>que_out_6_2_9, B1=>nx10360, C0=>que_out_9_2_9, C1=>nx10334);
   ix8416 : aoi22 port map ( Y=>nx8415, A0=>que_out_5_2_9, A1=>nx10256, B0=>
      que_out_18_2_9, B1=>nx10282);
   ix8418 : aoi22 port map ( Y=>nx8417, A0=>que_out_17_2_9, A1=>nx10230, B0
      =>que_out_20_2_9, B1=>nx10204);
   ix4723 : nand03 port map ( Y=>nx4722, A0=>nx8421, A1=>nx8423, A2=>nx8425
   );
   ix8422 : aoi222 port map ( Y=>nx8421, A0=>que_out_19_2_9, A1=>nx10178, B0
      =>que_out_21_2_9, B1=>nx10152, C0=>que_out_8_2_9, C1=>nx10126);
   ix8424 : aoi22 port map ( Y=>nx8423, A0=>que_out_25_2_9, A1=>nx10074, B0
      =>que_out_16_2_9, B1=>nx10100);
   ix8426 : aoi22 port map ( Y=>nx8425, A0=>que_out_24_2_9, A1=>nx10048, B0
      =>que_out_22_2_9, B1=>nx10022);
   ix4695 : nand03 port map ( Y=>nx4694, A0=>nx8429, A1=>nx8431, A2=>nx8433
   );
   ix8430 : aoi222 port map ( Y=>nx8429, A0=>que_out_15_2_9, A1=>nx9970, B0
      =>que_out_3_2_9, B1=>nx9996, C0=>que_out_23_2_9, C1=>nx9944);
   ix8432 : aoi22 port map ( Y=>nx8431, A0=>que_out_27_2_9, A1=>nx9918, B0=>
      que_out_4_2_9, B1=>nx9892);
   ix8434 : aoi22 port map ( Y=>nx8433, A0=>que_out_0_2_9, A1=>nx9840, B0=>
      que_out_2_2_9, B1=>nx9866);
   ix4669 : nand03 port map ( Y=>nx4668, A0=>nx8437, A1=>nx8439, A2=>nx8441
   );
   ix8438 : aoi222 port map ( Y=>nx8437, A0=>que_out_26_2_9, A1=>nx9814, B0
      =>que_out_14_2_9, B1=>nx9788, C0=>que_out_11_2_9, C1=>nx9762);
   ix8440 : aoi22 port map ( Y=>nx8439, A0=>que_out_13_2_9, A1=>nx9736, B0=>
      que_out_7_2_9, B1=>nx9710);
   ix8442 : aoi22 port map ( Y=>nx8441, A0=>que_out_12_2_9, A1=>nx9684, B0=>
      que_out_1_2_9, B1=>nx9658);
   ix4863 : or04 port map ( Y=>out_column_2_10, A0=>nx4858, A1=>nx4832, A2=>
      nx4804, A3=>nx4778);
   ix4859 : nand03 port map ( Y=>nx4858, A0=>nx8447, A1=>nx8449, A2=>nx8451
   );
   ix8448 : aoi222 port map ( Y=>nx8447, A0=>que_out_10_2_10, A1=>nx10310, 
      B0=>que_out_6_2_10, B1=>nx10362, C0=>que_out_9_2_10, C1=>nx10336);
   ix8450 : aoi22 port map ( Y=>nx8449, A0=>que_out_5_2_10, A1=>nx10258, B0
      =>que_out_18_2_10, B1=>nx10284);
   ix8452 : aoi22 port map ( Y=>nx8451, A0=>que_out_17_2_10, A1=>nx10232, B0
      =>que_out_20_2_10, B1=>nx10206);
   ix4833 : nand03 port map ( Y=>nx4832, A0=>nx8455, A1=>nx8457, A2=>nx8459
   );
   ix8456 : aoi222 port map ( Y=>nx8455, A0=>que_out_19_2_10, A1=>nx10180, 
      B0=>que_out_21_2_10, B1=>nx10154, C0=>que_out_8_2_10, C1=>nx10128);
   ix8458 : aoi22 port map ( Y=>nx8457, A0=>que_out_25_2_10, A1=>nx10076, B0
      =>que_out_16_2_10, B1=>nx10102);
   ix8460 : aoi22 port map ( Y=>nx8459, A0=>que_out_24_2_10, A1=>nx10050, B0
      =>que_out_22_2_10, B1=>nx10024);
   ix4805 : nand03 port map ( Y=>nx4804, A0=>nx8463, A1=>nx8465, A2=>nx8467
   );
   ix8464 : aoi222 port map ( Y=>nx8463, A0=>que_out_15_2_10, A1=>nx9972, B0
      =>que_out_3_2_10, B1=>nx9998, C0=>que_out_23_2_10, C1=>nx9946);
   ix8466 : aoi22 port map ( Y=>nx8465, A0=>que_out_27_2_10, A1=>nx9920, B0
      =>que_out_4_2_10, B1=>nx9894);
   ix8468 : aoi22 port map ( Y=>nx8467, A0=>que_out_0_2_10, A1=>nx9842, B0=>
      que_out_2_2_10, B1=>nx9868);
   ix4779 : nand03 port map ( Y=>nx4778, A0=>nx8471, A1=>nx8473, A2=>nx8475
   );
   ix8472 : aoi222 port map ( Y=>nx8471, A0=>que_out_26_2_10, A1=>nx9816, B0
      =>que_out_14_2_10, B1=>nx9790, C0=>que_out_11_2_10, C1=>nx9764);
   ix8474 : aoi22 port map ( Y=>nx8473, A0=>que_out_13_2_10, A1=>nx9738, B0
      =>que_out_7_2_10, B1=>nx9712);
   ix8476 : aoi22 port map ( Y=>nx8475, A0=>que_out_12_2_10, A1=>nx9686, B0
      =>que_out_1_2_10, B1=>nx9660);
   ix4973 : or04 port map ( Y=>out_column_2_11, A0=>nx4968, A1=>nx4942, A2=>
      nx4914, A3=>nx4888);
   ix4969 : nand03 port map ( Y=>nx4968, A0=>nx8481, A1=>nx8483, A2=>nx8485
   );
   ix8482 : aoi222 port map ( Y=>nx8481, A0=>que_out_10_2_11, A1=>nx10310, 
      B0=>que_out_6_2_11, B1=>nx10362, C0=>que_out_9_2_11, C1=>nx10336);
   ix8484 : aoi22 port map ( Y=>nx8483, A0=>que_out_5_2_11, A1=>nx10258, B0
      =>que_out_18_2_11, B1=>nx10284);
   ix8486 : aoi22 port map ( Y=>nx8485, A0=>que_out_17_2_11, A1=>nx10232, B0
      =>que_out_20_2_11, B1=>nx10206);
   ix4943 : nand03 port map ( Y=>nx4942, A0=>nx8489, A1=>nx8491, A2=>nx8493
   );
   ix8490 : aoi222 port map ( Y=>nx8489, A0=>que_out_19_2_11, A1=>nx10180, 
      B0=>que_out_21_2_11, B1=>nx10154, C0=>que_out_8_2_11, C1=>nx10128);
   ix8492 : aoi22 port map ( Y=>nx8491, A0=>que_out_25_2_11, A1=>nx10076, B0
      =>que_out_16_2_11, B1=>nx10102);
   ix8494 : aoi22 port map ( Y=>nx8493, A0=>que_out_24_2_11, A1=>nx10050, B0
      =>que_out_22_2_11, B1=>nx10024);
   ix4915 : nand03 port map ( Y=>nx4914, A0=>nx8497, A1=>nx8499, A2=>nx8501
   );
   ix8498 : aoi222 port map ( Y=>nx8497, A0=>que_out_15_2_11, A1=>nx9972, B0
      =>que_out_3_2_11, B1=>nx9998, C0=>que_out_23_2_11, C1=>nx9946);
   ix8500 : aoi22 port map ( Y=>nx8499, A0=>que_out_27_2_11, A1=>nx9920, B0
      =>que_out_4_2_11, B1=>nx9894);
   ix8502 : aoi22 port map ( Y=>nx8501, A0=>que_out_0_2_11, A1=>nx9842, B0=>
      que_out_2_2_11, B1=>nx9868);
   ix4889 : nand03 port map ( Y=>nx4888, A0=>nx8505, A1=>nx8507, A2=>nx8509
   );
   ix8506 : aoi222 port map ( Y=>nx8505, A0=>que_out_26_2_11, A1=>nx9816, B0
      =>que_out_14_2_11, B1=>nx9790, C0=>que_out_11_2_11, C1=>nx9764);
   ix8508 : aoi22 port map ( Y=>nx8507, A0=>que_out_13_2_11, A1=>nx9738, B0
      =>que_out_7_2_11, B1=>nx9712);
   ix8510 : aoi22 port map ( Y=>nx8509, A0=>que_out_12_2_11, A1=>nx9686, B0
      =>que_out_1_2_11, B1=>nx9660);
   ix5083 : or04 port map ( Y=>out_column_2_12, A0=>nx5078, A1=>nx5052, A2=>
      nx5024, A3=>nx4998);
   ix5079 : nand03 port map ( Y=>nx5078, A0=>nx8515, A1=>nx8517, A2=>nx8519
   );
   ix8516 : aoi222 port map ( Y=>nx8515, A0=>que_out_10_2_12, A1=>nx10310, 
      B0=>que_out_6_2_12, B1=>nx10362, C0=>que_out_9_2_12, C1=>nx10336);
   ix8518 : aoi22 port map ( Y=>nx8517, A0=>que_out_5_2_12, A1=>nx10258, B0
      =>que_out_18_2_12, B1=>nx10284);
   ix8520 : aoi22 port map ( Y=>nx8519, A0=>que_out_17_2_12, A1=>nx10232, B0
      =>que_out_20_2_12, B1=>nx10206);
   ix5053 : nand03 port map ( Y=>nx5052, A0=>nx8523, A1=>nx8525, A2=>nx8527
   );
   ix8524 : aoi222 port map ( Y=>nx8523, A0=>que_out_19_2_12, A1=>nx10180, 
      B0=>que_out_21_2_12, B1=>nx10154, C0=>que_out_8_2_12, C1=>nx10128);
   ix8526 : aoi22 port map ( Y=>nx8525, A0=>que_out_25_2_12, A1=>nx10076, B0
      =>que_out_16_2_12, B1=>nx10102);
   ix8528 : aoi22 port map ( Y=>nx8527, A0=>que_out_24_2_12, A1=>nx10050, B0
      =>que_out_22_2_12, B1=>nx10024);
   ix5025 : nand03 port map ( Y=>nx5024, A0=>nx8531, A1=>nx8533, A2=>nx8535
   );
   ix8532 : aoi222 port map ( Y=>nx8531, A0=>que_out_15_2_12, A1=>nx9972, B0
      =>que_out_3_2_12, B1=>nx9998, C0=>que_out_23_2_12, C1=>nx9946);
   ix8534 : aoi22 port map ( Y=>nx8533, A0=>que_out_27_2_12, A1=>nx9920, B0
      =>que_out_4_2_12, B1=>nx9894);
   ix8536 : aoi22 port map ( Y=>nx8535, A0=>que_out_0_2_12, A1=>nx9842, B0=>
      que_out_2_2_12, B1=>nx9868);
   ix4999 : nand03 port map ( Y=>nx4998, A0=>nx8539, A1=>nx8541, A2=>nx8543
   );
   ix8540 : aoi222 port map ( Y=>nx8539, A0=>que_out_26_2_12, A1=>nx9816, B0
      =>que_out_14_2_12, B1=>nx9790, C0=>que_out_11_2_12, C1=>nx9764);
   ix8542 : aoi22 port map ( Y=>nx8541, A0=>que_out_13_2_12, A1=>nx9738, B0
      =>que_out_7_2_12, B1=>nx9712);
   ix8544 : aoi22 port map ( Y=>nx8543, A0=>que_out_12_2_12, A1=>nx9686, B0
      =>que_out_1_2_12, B1=>nx9660);
   ix5193 : or04 port map ( Y=>out_column_2_13, A0=>nx5188, A1=>nx5162, A2=>
      nx5134, A3=>nx5108);
   ix5189 : nand03 port map ( Y=>nx5188, A0=>nx8549, A1=>nx8551, A2=>nx8553
   );
   ix8550 : aoi222 port map ( Y=>nx8549, A0=>que_out_10_2_13, A1=>nx10310, 
      B0=>que_out_6_2_13, B1=>nx10362, C0=>que_out_9_2_13, C1=>nx10336);
   ix8552 : aoi22 port map ( Y=>nx8551, A0=>que_out_5_2_13, A1=>nx10258, B0
      =>que_out_18_2_13, B1=>nx10284);
   ix8554 : aoi22 port map ( Y=>nx8553, A0=>que_out_17_2_13, A1=>nx10232, B0
      =>que_out_20_2_13, B1=>nx10206);
   ix5163 : nand03 port map ( Y=>nx5162, A0=>nx8557, A1=>nx8559, A2=>nx8561
   );
   ix8558 : aoi222 port map ( Y=>nx8557, A0=>que_out_19_2_13, A1=>nx10180, 
      B0=>que_out_21_2_13, B1=>nx10154, C0=>que_out_8_2_13, C1=>nx10128);
   ix8560 : aoi22 port map ( Y=>nx8559, A0=>que_out_25_2_13, A1=>nx10076, B0
      =>que_out_16_2_13, B1=>nx10102);
   ix8562 : aoi22 port map ( Y=>nx8561, A0=>que_out_24_2_13, A1=>nx10050, B0
      =>que_out_22_2_13, B1=>nx10024);
   ix5135 : nand03 port map ( Y=>nx5134, A0=>nx8565, A1=>nx8567, A2=>nx8569
   );
   ix8566 : aoi222 port map ( Y=>nx8565, A0=>que_out_15_2_13, A1=>nx9972, B0
      =>que_out_3_2_13, B1=>nx9998, C0=>que_out_23_2_13, C1=>nx9946);
   ix8568 : aoi22 port map ( Y=>nx8567, A0=>que_out_27_2_13, A1=>nx9920, B0
      =>que_out_4_2_13, B1=>nx9894);
   ix8570 : aoi22 port map ( Y=>nx8569, A0=>que_out_0_2_13, A1=>nx9842, B0=>
      que_out_2_2_13, B1=>nx9868);
   ix5109 : nand03 port map ( Y=>nx5108, A0=>nx8573, A1=>nx8575, A2=>nx8577
   );
   ix8574 : aoi222 port map ( Y=>nx8573, A0=>que_out_26_2_13, A1=>nx9816, B0
      =>que_out_14_2_13, B1=>nx9790, C0=>que_out_11_2_13, C1=>nx9764);
   ix8576 : aoi22 port map ( Y=>nx8575, A0=>que_out_13_2_13, A1=>nx9738, B0
      =>que_out_7_2_13, B1=>nx9712);
   ix8578 : aoi22 port map ( Y=>nx8577, A0=>que_out_12_2_13, A1=>nx9686, B0
      =>que_out_1_2_13, B1=>nx9660);
   ix5303 : or04 port map ( Y=>out_column_2_14, A0=>nx5298, A1=>nx5272, A2=>
      nx5244, A3=>nx5218);
   ix5299 : nand03 port map ( Y=>nx5298, A0=>nx8583, A1=>nx8585, A2=>nx8587
   );
   ix8584 : aoi222 port map ( Y=>nx8583, A0=>que_out_10_2_14, A1=>nx10310, 
      B0=>que_out_6_2_14, B1=>nx10362, C0=>que_out_9_2_14, C1=>nx10336);
   ix8586 : aoi22 port map ( Y=>nx8585, A0=>que_out_5_2_14, A1=>nx10258, B0
      =>que_out_18_2_14, B1=>nx10284);
   ix8588 : aoi22 port map ( Y=>nx8587, A0=>que_out_17_2_14, A1=>nx10232, B0
      =>que_out_20_2_14, B1=>nx10206);
   ix5273 : nand03 port map ( Y=>nx5272, A0=>nx8591, A1=>nx8593, A2=>nx8595
   );
   ix8592 : aoi222 port map ( Y=>nx8591, A0=>que_out_19_2_14, A1=>nx10180, 
      B0=>que_out_21_2_14, B1=>nx10154, C0=>que_out_8_2_14, C1=>nx10128);
   ix8594 : aoi22 port map ( Y=>nx8593, A0=>que_out_25_2_14, A1=>nx10076, B0
      =>que_out_16_2_14, B1=>nx10102);
   ix8596 : aoi22 port map ( Y=>nx8595, A0=>que_out_24_2_14, A1=>nx10050, B0
      =>que_out_22_2_14, B1=>nx10024);
   ix5245 : nand03 port map ( Y=>nx5244, A0=>nx8599, A1=>nx8601, A2=>nx8603
   );
   ix8600 : aoi222 port map ( Y=>nx8599, A0=>que_out_15_2_14, A1=>nx9972, B0
      =>que_out_3_2_14, B1=>nx9998, C0=>que_out_23_2_14, C1=>nx9946);
   ix8602 : aoi22 port map ( Y=>nx8601, A0=>que_out_27_2_14, A1=>nx9920, B0
      =>que_out_4_2_14, B1=>nx9894);
   ix8604 : aoi22 port map ( Y=>nx8603, A0=>que_out_0_2_14, A1=>nx9842, B0=>
      que_out_2_2_14, B1=>nx9868);
   ix5219 : nand03 port map ( Y=>nx5218, A0=>nx8607, A1=>nx8609, A2=>nx8611
   );
   ix8608 : aoi222 port map ( Y=>nx8607, A0=>que_out_26_2_14, A1=>nx9816, B0
      =>que_out_14_2_14, B1=>nx9790, C0=>que_out_11_2_14, C1=>nx9764);
   ix8610 : aoi22 port map ( Y=>nx8609, A0=>que_out_13_2_14, A1=>nx9738, B0
      =>que_out_7_2_14, B1=>nx9712);
   ix8612 : aoi22 port map ( Y=>nx8611, A0=>que_out_12_2_14, A1=>nx9686, B0
      =>que_out_1_2_14, B1=>nx9660);
   ix5413 : or04 port map ( Y=>out_column_2_15, A0=>nx5408, A1=>nx5382, A2=>
      nx5354, A3=>nx5328);
   ix5409 : nand03 port map ( Y=>nx5408, A0=>nx8617, A1=>nx8619, A2=>nx8621
   );
   ix8618 : aoi222 port map ( Y=>nx8617, A0=>que_out_10_2_15, A1=>nx10310, 
      B0=>que_out_6_2_15, B1=>nx10362, C0=>que_out_9_2_15, C1=>nx10336);
   ix8620 : aoi22 port map ( Y=>nx8619, A0=>que_out_5_2_15, A1=>nx10258, B0
      =>que_out_18_2_15, B1=>nx10284);
   ix8622 : aoi22 port map ( Y=>nx8621, A0=>que_out_17_2_15, A1=>nx10232, B0
      =>que_out_20_2_15, B1=>nx10206);
   ix5383 : nand03 port map ( Y=>nx5382, A0=>nx8625, A1=>nx8627, A2=>nx8629
   );
   ix8626 : aoi222 port map ( Y=>nx8625, A0=>que_out_19_2_15, A1=>nx10180, 
      B0=>que_out_21_2_15, B1=>nx10154, C0=>que_out_8_2_15, C1=>nx10128);
   ix8628 : aoi22 port map ( Y=>nx8627, A0=>que_out_25_2_15, A1=>nx10076, B0
      =>que_out_16_2_15, B1=>nx10102);
   ix8630 : aoi22 port map ( Y=>nx8629, A0=>que_out_24_2_15, A1=>nx10050, B0
      =>que_out_22_2_15, B1=>nx10024);
   ix5355 : nand03 port map ( Y=>nx5354, A0=>nx8633, A1=>nx8635, A2=>nx8637
   );
   ix8634 : aoi222 port map ( Y=>nx8633, A0=>que_out_15_2_15, A1=>nx9972, B0
      =>que_out_3_2_15, B1=>nx9998, C0=>que_out_23_2_15, C1=>nx9946);
   ix8636 : aoi22 port map ( Y=>nx8635, A0=>que_out_27_2_15, A1=>nx9920, B0
      =>que_out_4_2_15, B1=>nx9894);
   ix8638 : aoi22 port map ( Y=>nx8637, A0=>que_out_0_2_15, A1=>nx9842, B0=>
      que_out_2_2_15, B1=>nx9868);
   ix5329 : nand03 port map ( Y=>nx5328, A0=>nx8641, A1=>nx8643, A2=>nx8645
   );
   ix8642 : aoi222 port map ( Y=>nx8641, A0=>que_out_26_2_15, A1=>nx9816, B0
      =>que_out_14_2_15, B1=>nx9790, C0=>que_out_11_2_15, C1=>nx9764);
   ix8644 : aoi22 port map ( Y=>nx8643, A0=>que_out_13_2_15, A1=>nx9738, B0
      =>que_out_7_2_15, B1=>nx9712);
   ix8646 : aoi22 port map ( Y=>nx8645, A0=>que_out_12_2_15, A1=>nx9686, B0
      =>que_out_1_2_15, B1=>nx9660);
   ix5523 : or04 port map ( Y=>out_column_1_0, A0=>nx5518, A1=>nx5492, A2=>
      nx5464, A3=>nx5438);
   ix5519 : nand03 port map ( Y=>nx5518, A0=>nx8651, A1=>nx8653, A2=>nx8655
   );
   ix8652 : aoi222 port map ( Y=>nx8651, A0=>que_out_10_1_0, A1=>nx10310, B0
      =>que_out_6_1_0, B1=>nx10362, C0=>que_out_9_1_0, C1=>nx10336);
   ix8654 : aoi22 port map ( Y=>nx8653, A0=>que_out_5_1_0, A1=>nx10258, B0=>
      que_out_18_1_0, B1=>nx10284);
   ix8656 : aoi22 port map ( Y=>nx8655, A0=>que_out_17_1_0, A1=>nx10232, B0
      =>que_out_20_1_0, B1=>nx10206);
   ix5493 : nand03 port map ( Y=>nx5492, A0=>nx8659, A1=>nx8661, A2=>nx8663
   );
   ix8660 : aoi222 port map ( Y=>nx8659, A0=>que_out_19_1_0, A1=>nx10180, B0
      =>que_out_21_1_0, B1=>nx10154, C0=>que_out_8_1_0, C1=>nx10128);
   ix8662 : aoi22 port map ( Y=>nx8661, A0=>que_out_25_1_0, A1=>nx10076, B0
      =>que_out_16_1_0, B1=>nx10102);
   ix8664 : aoi22 port map ( Y=>nx8663, A0=>que_out_24_1_0, A1=>nx10050, B0
      =>que_out_22_1_0, B1=>nx10024);
   ix5465 : nand03 port map ( Y=>nx5464, A0=>nx8667, A1=>nx8669, A2=>nx8671
   );
   ix8668 : aoi222 port map ( Y=>nx8667, A0=>que_out_15_1_0, A1=>nx9972, B0
      =>que_out_3_1_0, B1=>nx9998, C0=>que_out_23_1_0, C1=>nx9946);
   ix8670 : aoi22 port map ( Y=>nx8669, A0=>que_out_27_1_0, A1=>nx9920, B0=>
      que_out_4_1_0, B1=>nx9894);
   ix8672 : aoi22 port map ( Y=>nx8671, A0=>que_out_0_1_0, A1=>nx9842, B0=>
      que_out_2_1_0, B1=>nx9868);
   ix5439 : nand03 port map ( Y=>nx5438, A0=>nx8675, A1=>nx8677, A2=>nx8679
   );
   ix8676 : aoi222 port map ( Y=>nx8675, A0=>que_out_26_1_0, A1=>nx9816, B0
      =>que_out_14_1_0, B1=>nx9790, C0=>que_out_11_1_0, C1=>nx9764);
   ix8678 : aoi22 port map ( Y=>nx8677, A0=>que_out_13_1_0, A1=>nx9738, B0=>
      que_out_7_1_0, B1=>nx9712);
   ix8680 : aoi22 port map ( Y=>nx8679, A0=>que_out_12_1_0, A1=>nx9686, B0=>
      que_out_1_1_0, B1=>nx9660);
   ix5633 : or04 port map ( Y=>out_column_1_1, A0=>nx5628, A1=>nx5602, A2=>
      nx5574, A3=>nx5548);
   ix5629 : nand03 port map ( Y=>nx5628, A0=>nx8685, A1=>nx8687, A2=>nx8689
   );
   ix8686 : aoi222 port map ( Y=>nx8685, A0=>que_out_10_1_1, A1=>nx10312, B0
      =>que_out_6_1_1, B1=>nx10364, C0=>que_out_9_1_1, C1=>nx10338);
   ix8688 : aoi22 port map ( Y=>nx8687, A0=>que_out_5_1_1, A1=>nx10260, B0=>
      que_out_18_1_1, B1=>nx10286);
   ix8690 : aoi22 port map ( Y=>nx8689, A0=>que_out_17_1_1, A1=>nx10234, B0
      =>que_out_20_1_1, B1=>nx10208);
   ix5603 : nand03 port map ( Y=>nx5602, A0=>nx8693, A1=>nx8695, A2=>nx8697
   );
   ix8694 : aoi222 port map ( Y=>nx8693, A0=>que_out_19_1_1, A1=>nx10182, B0
      =>que_out_21_1_1, B1=>nx10156, C0=>que_out_8_1_1, C1=>nx10130);
   ix8696 : aoi22 port map ( Y=>nx8695, A0=>que_out_25_1_1, A1=>nx10078, B0
      =>que_out_16_1_1, B1=>nx10104);
   ix8698 : aoi22 port map ( Y=>nx8697, A0=>que_out_24_1_1, A1=>nx10052, B0
      =>que_out_22_1_1, B1=>nx10026);
   ix5575 : nand03 port map ( Y=>nx5574, A0=>nx8701, A1=>nx8703, A2=>nx8705
   );
   ix8702 : aoi222 port map ( Y=>nx8701, A0=>que_out_15_1_1, A1=>nx9974, B0
      =>que_out_3_1_1, B1=>nx10000, C0=>que_out_23_1_1, C1=>nx9948);
   ix8704 : aoi22 port map ( Y=>nx8703, A0=>que_out_27_1_1, A1=>nx9922, B0=>
      que_out_4_1_1, B1=>nx9896);
   ix8706 : aoi22 port map ( Y=>nx8705, A0=>que_out_0_1_1, A1=>nx9844, B0=>
      que_out_2_1_1, B1=>nx9870);
   ix5549 : nand03 port map ( Y=>nx5548, A0=>nx8709, A1=>nx8711, A2=>nx8713
   );
   ix8710 : aoi222 port map ( Y=>nx8709, A0=>que_out_26_1_1, A1=>nx9818, B0
      =>que_out_14_1_1, B1=>nx9792, C0=>que_out_11_1_1, C1=>nx9766);
   ix8712 : aoi22 port map ( Y=>nx8711, A0=>que_out_13_1_1, A1=>nx9740, B0=>
      que_out_7_1_1, B1=>nx9714);
   ix8714 : aoi22 port map ( Y=>nx8713, A0=>que_out_12_1_1, A1=>nx9688, B0=>
      que_out_1_1_1, B1=>nx9662);
   ix5743 : or04 port map ( Y=>out_column_1_2, A0=>nx5738, A1=>nx5712, A2=>
      nx5684, A3=>nx5658);
   ix5739 : nand03 port map ( Y=>nx5738, A0=>nx8719, A1=>nx8721, A2=>nx8723
   );
   ix8720 : aoi222 port map ( Y=>nx8719, A0=>que_out_10_1_2, A1=>nx10312, B0
      =>que_out_6_1_2, B1=>nx10364, C0=>que_out_9_1_2, C1=>nx10338);
   ix8722 : aoi22 port map ( Y=>nx8721, A0=>que_out_5_1_2, A1=>nx10260, B0=>
      que_out_18_1_2, B1=>nx10286);
   ix8724 : aoi22 port map ( Y=>nx8723, A0=>que_out_17_1_2, A1=>nx10234, B0
      =>que_out_20_1_2, B1=>nx10208);
   ix5713 : nand03 port map ( Y=>nx5712, A0=>nx8727, A1=>nx8729, A2=>nx8731
   );
   ix8728 : aoi222 port map ( Y=>nx8727, A0=>que_out_19_1_2, A1=>nx10182, B0
      =>que_out_21_1_2, B1=>nx10156, C0=>que_out_8_1_2, C1=>nx10130);
   ix8730 : aoi22 port map ( Y=>nx8729, A0=>que_out_25_1_2, A1=>nx10078, B0
      =>que_out_16_1_2, B1=>nx10104);
   ix8732 : aoi22 port map ( Y=>nx8731, A0=>que_out_24_1_2, A1=>nx10052, B0
      =>que_out_22_1_2, B1=>nx10026);
   ix5685 : nand03 port map ( Y=>nx5684, A0=>nx8735, A1=>nx8737, A2=>nx8739
   );
   ix8736 : aoi222 port map ( Y=>nx8735, A0=>que_out_15_1_2, A1=>nx9974, B0
      =>que_out_3_1_2, B1=>nx10000, C0=>que_out_23_1_2, C1=>nx9948);
   ix8738 : aoi22 port map ( Y=>nx8737, A0=>que_out_27_1_2, A1=>nx9922, B0=>
      que_out_4_1_2, B1=>nx9896);
   ix8740 : aoi22 port map ( Y=>nx8739, A0=>que_out_0_1_2, A1=>nx9844, B0=>
      que_out_2_1_2, B1=>nx9870);
   ix5659 : nand03 port map ( Y=>nx5658, A0=>nx8743, A1=>nx8745, A2=>nx8747
   );
   ix8744 : aoi222 port map ( Y=>nx8743, A0=>que_out_26_1_2, A1=>nx9818, B0
      =>que_out_14_1_2, B1=>nx9792, C0=>que_out_11_1_2, C1=>nx9766);
   ix8746 : aoi22 port map ( Y=>nx8745, A0=>que_out_13_1_2, A1=>nx9740, B0=>
      que_out_7_1_2, B1=>nx9714);
   ix8748 : aoi22 port map ( Y=>nx8747, A0=>que_out_12_1_2, A1=>nx9688, B0=>
      que_out_1_1_2, B1=>nx9662);
   ix5853 : or04 port map ( Y=>out_column_1_3, A0=>nx5848, A1=>nx5822, A2=>
      nx5794, A3=>nx5768);
   ix5849 : nand03 port map ( Y=>nx5848, A0=>nx8753, A1=>nx8755, A2=>nx8757
   );
   ix8754 : aoi222 port map ( Y=>nx8753, A0=>que_out_10_1_3, A1=>nx10312, B0
      =>que_out_6_1_3, B1=>nx10364, C0=>que_out_9_1_3, C1=>nx10338);
   ix8756 : aoi22 port map ( Y=>nx8755, A0=>que_out_5_1_3, A1=>nx10260, B0=>
      que_out_18_1_3, B1=>nx10286);
   ix8758 : aoi22 port map ( Y=>nx8757, A0=>que_out_17_1_3, A1=>nx10234, B0
      =>que_out_20_1_3, B1=>nx10208);
   ix5823 : nand03 port map ( Y=>nx5822, A0=>nx8761, A1=>nx8763, A2=>nx8765
   );
   ix8762 : aoi222 port map ( Y=>nx8761, A0=>que_out_19_1_3, A1=>nx10182, B0
      =>que_out_21_1_3, B1=>nx10156, C0=>que_out_8_1_3, C1=>nx10130);
   ix8764 : aoi22 port map ( Y=>nx8763, A0=>que_out_25_1_3, A1=>nx10078, B0
      =>que_out_16_1_3, B1=>nx10104);
   ix8766 : aoi22 port map ( Y=>nx8765, A0=>que_out_24_1_3, A1=>nx10052, B0
      =>que_out_22_1_3, B1=>nx10026);
   ix5795 : nand03 port map ( Y=>nx5794, A0=>nx8769, A1=>nx8771, A2=>nx8773
   );
   ix8770 : aoi222 port map ( Y=>nx8769, A0=>que_out_15_1_3, A1=>nx9974, B0
      =>que_out_3_1_3, B1=>nx10000, C0=>que_out_23_1_3, C1=>nx9948);
   ix8772 : aoi22 port map ( Y=>nx8771, A0=>que_out_27_1_3, A1=>nx9922, B0=>
      que_out_4_1_3, B1=>nx9896);
   ix8774 : aoi22 port map ( Y=>nx8773, A0=>que_out_0_1_3, A1=>nx9844, B0=>
      que_out_2_1_3, B1=>nx9870);
   ix5769 : nand03 port map ( Y=>nx5768, A0=>nx8777, A1=>nx8779, A2=>nx8781
   );
   ix8778 : aoi222 port map ( Y=>nx8777, A0=>que_out_26_1_3, A1=>nx9818, B0
      =>que_out_14_1_3, B1=>nx9792, C0=>que_out_11_1_3, C1=>nx9766);
   ix8780 : aoi22 port map ( Y=>nx8779, A0=>que_out_13_1_3, A1=>nx9740, B0=>
      que_out_7_1_3, B1=>nx9714);
   ix8782 : aoi22 port map ( Y=>nx8781, A0=>que_out_12_1_3, A1=>nx9688, B0=>
      que_out_1_1_3, B1=>nx9662);
   ix5963 : or04 port map ( Y=>out_column_1_4, A0=>nx5958, A1=>nx5932, A2=>
      nx5904, A3=>nx5878);
   ix5959 : nand03 port map ( Y=>nx5958, A0=>nx8787, A1=>nx8789, A2=>nx8791
   );
   ix8788 : aoi222 port map ( Y=>nx8787, A0=>que_out_10_1_4, A1=>nx10312, B0
      =>que_out_6_1_4, B1=>nx10364, C0=>que_out_9_1_4, C1=>nx10338);
   ix8790 : aoi22 port map ( Y=>nx8789, A0=>que_out_5_1_4, A1=>nx10260, B0=>
      que_out_18_1_4, B1=>nx10286);
   ix8792 : aoi22 port map ( Y=>nx8791, A0=>que_out_17_1_4, A1=>nx10234, B0
      =>que_out_20_1_4, B1=>nx10208);
   ix5933 : nand03 port map ( Y=>nx5932, A0=>nx8795, A1=>nx8797, A2=>nx8799
   );
   ix8796 : aoi222 port map ( Y=>nx8795, A0=>que_out_19_1_4, A1=>nx10182, B0
      =>que_out_21_1_4, B1=>nx10156, C0=>que_out_8_1_4, C1=>nx10130);
   ix8798 : aoi22 port map ( Y=>nx8797, A0=>que_out_25_1_4, A1=>nx10078, B0
      =>que_out_16_1_4, B1=>nx10104);
   ix8800 : aoi22 port map ( Y=>nx8799, A0=>que_out_24_1_4, A1=>nx10052, B0
      =>que_out_22_1_4, B1=>nx10026);
   ix5905 : nand03 port map ( Y=>nx5904, A0=>nx8803, A1=>nx8805, A2=>nx8807
   );
   ix8804 : aoi222 port map ( Y=>nx8803, A0=>que_out_15_1_4, A1=>nx9974, B0
      =>que_out_3_1_4, B1=>nx10000, C0=>que_out_23_1_4, C1=>nx9948);
   ix8806 : aoi22 port map ( Y=>nx8805, A0=>que_out_27_1_4, A1=>nx9922, B0=>
      que_out_4_1_4, B1=>nx9896);
   ix8808 : aoi22 port map ( Y=>nx8807, A0=>que_out_0_1_4, A1=>nx9844, B0=>
      que_out_2_1_4, B1=>nx9870);
   ix5879 : nand03 port map ( Y=>nx5878, A0=>nx8811, A1=>nx8813, A2=>nx8815
   );
   ix8812 : aoi222 port map ( Y=>nx8811, A0=>que_out_26_1_4, A1=>nx9818, B0
      =>que_out_14_1_4, B1=>nx9792, C0=>que_out_11_1_4, C1=>nx9766);
   ix8814 : aoi22 port map ( Y=>nx8813, A0=>que_out_13_1_4, A1=>nx9740, B0=>
      que_out_7_1_4, B1=>nx9714);
   ix8816 : aoi22 port map ( Y=>nx8815, A0=>que_out_12_1_4, A1=>nx9688, B0=>
      que_out_1_1_4, B1=>nx9662);
   ix6073 : or04 port map ( Y=>out_column_1_5, A0=>nx6068, A1=>nx6042, A2=>
      nx6014, A3=>nx5988);
   ix6069 : nand03 port map ( Y=>nx6068, A0=>nx8821, A1=>nx8823, A2=>nx8825
   );
   ix8822 : aoi222 port map ( Y=>nx8821, A0=>que_out_10_1_5, A1=>nx10312, B0
      =>que_out_6_1_5, B1=>nx10364, C0=>que_out_9_1_5, C1=>nx10338);
   ix8824 : aoi22 port map ( Y=>nx8823, A0=>que_out_5_1_5, A1=>nx10260, B0=>
      que_out_18_1_5, B1=>nx10286);
   ix8826 : aoi22 port map ( Y=>nx8825, A0=>que_out_17_1_5, A1=>nx10234, B0
      =>que_out_20_1_5, B1=>nx10208);
   ix6043 : nand03 port map ( Y=>nx6042, A0=>nx8829, A1=>nx8831, A2=>nx8833
   );
   ix8830 : aoi222 port map ( Y=>nx8829, A0=>que_out_19_1_5, A1=>nx10182, B0
      =>que_out_21_1_5, B1=>nx10156, C0=>que_out_8_1_5, C1=>nx10130);
   ix8832 : aoi22 port map ( Y=>nx8831, A0=>que_out_25_1_5, A1=>nx10078, B0
      =>que_out_16_1_5, B1=>nx10104);
   ix8834 : aoi22 port map ( Y=>nx8833, A0=>que_out_24_1_5, A1=>nx10052, B0
      =>que_out_22_1_5, B1=>nx10026);
   ix6015 : nand03 port map ( Y=>nx6014, A0=>nx8837, A1=>nx8839, A2=>nx8841
   );
   ix8838 : aoi222 port map ( Y=>nx8837, A0=>que_out_15_1_5, A1=>nx9974, B0
      =>que_out_3_1_5, B1=>nx10000, C0=>que_out_23_1_5, C1=>nx9948);
   ix8840 : aoi22 port map ( Y=>nx8839, A0=>que_out_27_1_5, A1=>nx9922, B0=>
      que_out_4_1_5, B1=>nx9896);
   ix8842 : aoi22 port map ( Y=>nx8841, A0=>que_out_0_1_5, A1=>nx9844, B0=>
      que_out_2_1_5, B1=>nx9870);
   ix5989 : nand03 port map ( Y=>nx5988, A0=>nx8845, A1=>nx8847, A2=>nx8849
   );
   ix8846 : aoi222 port map ( Y=>nx8845, A0=>que_out_26_1_5, A1=>nx9818, B0
      =>que_out_14_1_5, B1=>nx9792, C0=>que_out_11_1_5, C1=>nx9766);
   ix8848 : aoi22 port map ( Y=>nx8847, A0=>que_out_13_1_5, A1=>nx9740, B0=>
      que_out_7_1_5, B1=>nx9714);
   ix8850 : aoi22 port map ( Y=>nx8849, A0=>que_out_12_1_5, A1=>nx9688, B0=>
      que_out_1_1_5, B1=>nx9662);
   ix6183 : or04 port map ( Y=>out_column_1_6, A0=>nx6178, A1=>nx6152, A2=>
      nx6124, A3=>nx6098);
   ix6179 : nand03 port map ( Y=>nx6178, A0=>nx8855, A1=>nx8857, A2=>nx8859
   );
   ix8856 : aoi222 port map ( Y=>nx8855, A0=>que_out_10_1_6, A1=>nx10312, B0
      =>que_out_6_1_6, B1=>nx10364, C0=>que_out_9_1_6, C1=>nx10338);
   ix8858 : aoi22 port map ( Y=>nx8857, A0=>que_out_5_1_6, A1=>nx10260, B0=>
      que_out_18_1_6, B1=>nx10286);
   ix8860 : aoi22 port map ( Y=>nx8859, A0=>que_out_17_1_6, A1=>nx10234, B0
      =>que_out_20_1_6, B1=>nx10208);
   ix6153 : nand03 port map ( Y=>nx6152, A0=>nx8863, A1=>nx8865, A2=>nx8867
   );
   ix8864 : aoi222 port map ( Y=>nx8863, A0=>que_out_19_1_6, A1=>nx10182, B0
      =>que_out_21_1_6, B1=>nx10156, C0=>que_out_8_1_6, C1=>nx10130);
   ix8866 : aoi22 port map ( Y=>nx8865, A0=>que_out_25_1_6, A1=>nx10078, B0
      =>que_out_16_1_6, B1=>nx10104);
   ix8868 : aoi22 port map ( Y=>nx8867, A0=>que_out_24_1_6, A1=>nx10052, B0
      =>que_out_22_1_6, B1=>nx10026);
   ix6125 : nand03 port map ( Y=>nx6124, A0=>nx8871, A1=>nx8873, A2=>nx8875
   );
   ix8872 : aoi222 port map ( Y=>nx8871, A0=>que_out_15_1_6, A1=>nx9974, B0
      =>que_out_3_1_6, B1=>nx10000, C0=>que_out_23_1_6, C1=>nx9948);
   ix8874 : aoi22 port map ( Y=>nx8873, A0=>que_out_27_1_6, A1=>nx9922, B0=>
      que_out_4_1_6, B1=>nx9896);
   ix8876 : aoi22 port map ( Y=>nx8875, A0=>que_out_0_1_6, A1=>nx9844, B0=>
      que_out_2_1_6, B1=>nx9870);
   ix6099 : nand03 port map ( Y=>nx6098, A0=>nx8879, A1=>nx8881, A2=>nx8883
   );
   ix8880 : aoi222 port map ( Y=>nx8879, A0=>que_out_26_1_6, A1=>nx9818, B0
      =>que_out_14_1_6, B1=>nx9792, C0=>que_out_11_1_6, C1=>nx9766);
   ix8882 : aoi22 port map ( Y=>nx8881, A0=>que_out_13_1_6, A1=>nx9740, B0=>
      que_out_7_1_6, B1=>nx9714);
   ix8884 : aoi22 port map ( Y=>nx8883, A0=>que_out_12_1_6, A1=>nx9688, B0=>
      que_out_1_1_6, B1=>nx9662);
   ix6293 : or04 port map ( Y=>out_column_1_7, A0=>nx6288, A1=>nx6262, A2=>
      nx6234, A3=>nx6208);
   ix6289 : nand03 port map ( Y=>nx6288, A0=>nx8889, A1=>nx8891, A2=>nx8893
   );
   ix8890 : aoi222 port map ( Y=>nx8889, A0=>que_out_10_1_7, A1=>nx10312, B0
      =>que_out_6_1_7, B1=>nx10364, C0=>que_out_9_1_7, C1=>nx10338);
   ix8892 : aoi22 port map ( Y=>nx8891, A0=>que_out_5_1_7, A1=>nx10260, B0=>
      que_out_18_1_7, B1=>nx10286);
   ix8894 : aoi22 port map ( Y=>nx8893, A0=>que_out_17_1_7, A1=>nx10234, B0
      =>que_out_20_1_7, B1=>nx10208);
   ix6263 : nand03 port map ( Y=>nx6262, A0=>nx8897, A1=>nx8899, A2=>nx8901
   );
   ix8898 : aoi222 port map ( Y=>nx8897, A0=>que_out_19_1_7, A1=>nx10182, B0
      =>que_out_21_1_7, B1=>nx10156, C0=>que_out_8_1_7, C1=>nx10130);
   ix8900 : aoi22 port map ( Y=>nx8899, A0=>que_out_25_1_7, A1=>nx10078, B0
      =>que_out_16_1_7, B1=>nx10104);
   ix8902 : aoi22 port map ( Y=>nx8901, A0=>que_out_24_1_7, A1=>nx10052, B0
      =>que_out_22_1_7, B1=>nx10026);
   ix6235 : nand03 port map ( Y=>nx6234, A0=>nx8905, A1=>nx8907, A2=>nx8909
   );
   ix8906 : aoi222 port map ( Y=>nx8905, A0=>que_out_15_1_7, A1=>nx9974, B0
      =>que_out_3_1_7, B1=>nx10000, C0=>que_out_23_1_7, C1=>nx9948);
   ix8908 : aoi22 port map ( Y=>nx8907, A0=>que_out_27_1_7, A1=>nx9922, B0=>
      que_out_4_1_7, B1=>nx9896);
   ix8910 : aoi22 port map ( Y=>nx8909, A0=>que_out_0_1_7, A1=>nx9844, B0=>
      que_out_2_1_7, B1=>nx9870);
   ix6209 : nand03 port map ( Y=>nx6208, A0=>nx8913, A1=>nx8915, A2=>nx8917
   );
   ix8914 : aoi222 port map ( Y=>nx8913, A0=>que_out_26_1_7, A1=>nx9818, B0
      =>que_out_14_1_7, B1=>nx9792, C0=>que_out_11_1_7, C1=>nx9766);
   ix8916 : aoi22 port map ( Y=>nx8915, A0=>que_out_13_1_7, A1=>nx9740, B0=>
      que_out_7_1_7, B1=>nx9714);
   ix8918 : aoi22 port map ( Y=>nx8917, A0=>que_out_12_1_7, A1=>nx9688, B0=>
      que_out_1_1_7, B1=>nx9662);
   ix6403 : or04 port map ( Y=>out_column_1_8, A0=>nx6398, A1=>nx6372, A2=>
      nx6344, A3=>nx6318);
   ix6399 : nand03 port map ( Y=>nx6398, A0=>nx8923, A1=>nx8925, A2=>nx8927
   );
   ix8924 : aoi222 port map ( Y=>nx8923, A0=>que_out_10_1_8, A1=>nx10314, B0
      =>que_out_6_1_8, B1=>nx10366, C0=>que_out_9_1_8, C1=>nx10340);
   ix8926 : aoi22 port map ( Y=>nx8925, A0=>que_out_5_1_8, A1=>nx10262, B0=>
      que_out_18_1_8, B1=>nx10288);
   ix8928 : aoi22 port map ( Y=>nx8927, A0=>que_out_17_1_8, A1=>nx10236, B0
      =>que_out_20_1_8, B1=>nx10210);
   ix6373 : nand03 port map ( Y=>nx6372, A0=>nx8931, A1=>nx8933, A2=>nx8935
   );
   ix8932 : aoi222 port map ( Y=>nx8931, A0=>que_out_19_1_8, A1=>nx10184, B0
      =>que_out_21_1_8, B1=>nx10158, C0=>que_out_8_1_8, C1=>nx10132);
   ix8934 : aoi22 port map ( Y=>nx8933, A0=>que_out_25_1_8, A1=>nx10080, B0
      =>que_out_16_1_8, B1=>nx10106);
   ix8936 : aoi22 port map ( Y=>nx8935, A0=>que_out_24_1_8, A1=>nx10054, B0
      =>que_out_22_1_8, B1=>nx10028);
   ix6345 : nand03 port map ( Y=>nx6344, A0=>nx8939, A1=>nx8941, A2=>nx8943
   );
   ix8940 : aoi222 port map ( Y=>nx8939, A0=>que_out_15_1_8, A1=>nx9976, B0
      =>que_out_3_1_8, B1=>nx10002, C0=>que_out_23_1_8, C1=>nx9950);
   ix8942 : aoi22 port map ( Y=>nx8941, A0=>que_out_27_1_8, A1=>nx9924, B0=>
      que_out_4_1_8, B1=>nx9898);
   ix8944 : aoi22 port map ( Y=>nx8943, A0=>que_out_0_1_8, A1=>nx9846, B0=>
      que_out_2_1_8, B1=>nx9872);
   ix6319 : nand03 port map ( Y=>nx6318, A0=>nx8947, A1=>nx8949, A2=>nx8951
   );
   ix8948 : aoi222 port map ( Y=>nx8947, A0=>que_out_26_1_8, A1=>nx9820, B0
      =>que_out_14_1_8, B1=>nx9794, C0=>que_out_11_1_8, C1=>nx9768);
   ix8950 : aoi22 port map ( Y=>nx8949, A0=>que_out_13_1_8, A1=>nx9742, B0=>
      que_out_7_1_8, B1=>nx9716);
   ix8952 : aoi22 port map ( Y=>nx8951, A0=>que_out_12_1_8, A1=>nx9690, B0=>
      que_out_1_1_8, B1=>nx9664);
   ix6513 : or04 port map ( Y=>out_column_1_9, A0=>nx6508, A1=>nx6482, A2=>
      nx6454, A3=>nx6428);
   ix6509 : nand03 port map ( Y=>nx6508, A0=>nx8955, A1=>nx8957, A2=>nx8959
   );
   ix8956 : aoi222 port map ( Y=>nx8955, A0=>que_out_10_1_9, A1=>nx10314, B0
      =>que_out_6_1_9, B1=>nx10366, C0=>que_out_9_1_9, C1=>nx10340);
   ix8958 : aoi22 port map ( Y=>nx8957, A0=>que_out_5_1_9, A1=>nx10262, B0=>
      que_out_18_1_9, B1=>nx10288);
   ix8960 : aoi22 port map ( Y=>nx8959, A0=>que_out_17_1_9, A1=>nx10236, B0
      =>que_out_20_1_9, B1=>nx10210);
   ix6483 : nand03 port map ( Y=>nx6482, A0=>nx8963, A1=>nx8965, A2=>nx8967
   );
   ix8964 : aoi222 port map ( Y=>nx8963, A0=>que_out_19_1_9, A1=>nx10184, B0
      =>que_out_21_1_9, B1=>nx10158, C0=>que_out_8_1_9, C1=>nx10132);
   ix8966 : aoi22 port map ( Y=>nx8965, A0=>que_out_25_1_9, A1=>nx10080, B0
      =>que_out_16_1_9, B1=>nx10106);
   ix8968 : aoi22 port map ( Y=>nx8967, A0=>que_out_24_1_9, A1=>nx10054, B0
      =>que_out_22_1_9, B1=>nx10028);
   ix6455 : nand03 port map ( Y=>nx6454, A0=>nx8970, A1=>nx8973, A2=>nx8975
   );
   ix8972 : aoi222 port map ( Y=>nx8970, A0=>que_out_15_1_9, A1=>nx9976, B0
      =>que_out_3_1_9, B1=>nx10002, C0=>que_out_23_1_9, C1=>nx9950);
   ix8974 : aoi22 port map ( Y=>nx8973, A0=>que_out_27_1_9, A1=>nx9924, B0=>
      que_out_4_1_9, B1=>nx9898);
   ix8976 : aoi22 port map ( Y=>nx8975, A0=>que_out_0_1_9, A1=>nx9846, B0=>
      que_out_2_1_9, B1=>nx9872);
   ix6429 : nand03 port map ( Y=>nx6428, A0=>nx8978, A1=>nx8981, A2=>nx8983
   );
   ix8980 : aoi222 port map ( Y=>nx8978, A0=>que_out_26_1_9, A1=>nx9820, B0
      =>que_out_14_1_9, B1=>nx9794, C0=>que_out_11_1_9, C1=>nx9768);
   ix8982 : aoi22 port map ( Y=>nx8981, A0=>que_out_13_1_9, A1=>nx9742, B0=>
      que_out_7_1_9, B1=>nx9716);
   ix8984 : aoi22 port map ( Y=>nx8983, A0=>que_out_12_1_9, A1=>nx9690, B0=>
      que_out_1_1_9, B1=>nx9664);
   ix6623 : or04 port map ( Y=>out_column_1_10, A0=>nx6618, A1=>nx6592, A2=>
      nx6564, A3=>nx6538);
   ix6619 : nand03 port map ( Y=>nx6618, A0=>nx8989, A1=>nx8991, A2=>nx8993
   );
   ix8990 : aoi222 port map ( Y=>nx8989, A0=>que_out_10_1_10, A1=>nx10314, 
      B0=>que_out_6_1_10, B1=>nx10366, C0=>que_out_9_1_10, C1=>nx10340);
   ix8992 : aoi22 port map ( Y=>nx8991, A0=>que_out_5_1_10, A1=>nx10262, B0
      =>que_out_18_1_10, B1=>nx10288);
   ix8994 : aoi22 port map ( Y=>nx8993, A0=>que_out_17_1_10, A1=>nx10236, B0
      =>que_out_20_1_10, B1=>nx10210);
   ix6593 : nand03 port map ( Y=>nx6592, A0=>nx8997, A1=>nx8999, A2=>nx9001
   );
   ix8998 : aoi222 port map ( Y=>nx8997, A0=>que_out_19_1_10, A1=>nx10184, 
      B0=>que_out_21_1_10, B1=>nx10158, C0=>que_out_8_1_10, C1=>nx10132);
   ix9000 : aoi22 port map ( Y=>nx8999, A0=>que_out_25_1_10, A1=>nx10080, B0
      =>que_out_16_1_10, B1=>nx10106);
   ix9002 : aoi22 port map ( Y=>nx9001, A0=>que_out_24_1_10, A1=>nx10054, B0
      =>que_out_22_1_10, B1=>nx10028);
   ix6565 : nand03 port map ( Y=>nx6564, A0=>nx9005, A1=>nx9007, A2=>nx9009
   );
   ix9006 : aoi222 port map ( Y=>nx9005, A0=>que_out_15_1_10, A1=>nx9976, B0
      =>que_out_3_1_10, B1=>nx10002, C0=>que_out_23_1_10, C1=>nx9950);
   ix9008 : aoi22 port map ( Y=>nx9007, A0=>que_out_27_1_10, A1=>nx9924, B0
      =>que_out_4_1_10, B1=>nx9898);
   ix9010 : aoi22 port map ( Y=>nx9009, A0=>que_out_0_1_10, A1=>nx9846, B0=>
      que_out_2_1_10, B1=>nx9872);
   ix6539 : nand03 port map ( Y=>nx6538, A0=>nx9013, A1=>nx9015, A2=>nx9017
   );
   ix9014 : aoi222 port map ( Y=>nx9013, A0=>que_out_26_1_10, A1=>nx9820, B0
      =>que_out_14_1_10, B1=>nx9794, C0=>que_out_11_1_10, C1=>nx9768);
   ix9016 : aoi22 port map ( Y=>nx9015, A0=>que_out_13_1_10, A1=>nx9742, B0
      =>que_out_7_1_10, B1=>nx9716);
   ix9018 : aoi22 port map ( Y=>nx9017, A0=>que_out_12_1_10, A1=>nx9690, B0
      =>que_out_1_1_10, B1=>nx9664);
   ix6733 : or04 port map ( Y=>out_column_1_11, A0=>nx6728, A1=>nx6702, A2=>
      nx6674, A3=>nx6648);
   ix6729 : nand03 port map ( Y=>nx6728, A0=>nx9023, A1=>nx9025, A2=>nx9027
   );
   ix9024 : aoi222 port map ( Y=>nx9023, A0=>que_out_10_1_11, A1=>nx10314, 
      B0=>que_out_6_1_11, B1=>nx10366, C0=>que_out_9_1_11, C1=>nx10340);
   ix9026 : aoi22 port map ( Y=>nx9025, A0=>que_out_5_1_11, A1=>nx10262, B0
      =>que_out_18_1_11, B1=>nx10288);
   ix9028 : aoi22 port map ( Y=>nx9027, A0=>que_out_17_1_11, A1=>nx10236, B0
      =>que_out_20_1_11, B1=>nx10210);
   ix6703 : nand03 port map ( Y=>nx6702, A0=>nx9031, A1=>nx9033, A2=>nx9035
   );
   ix9032 : aoi222 port map ( Y=>nx9031, A0=>que_out_19_1_11, A1=>nx10184, 
      B0=>que_out_21_1_11, B1=>nx10158, C0=>que_out_8_1_11, C1=>nx10132);
   ix9034 : aoi22 port map ( Y=>nx9033, A0=>que_out_25_1_11, A1=>nx10080, B0
      =>que_out_16_1_11, B1=>nx10106);
   ix9036 : aoi22 port map ( Y=>nx9035, A0=>que_out_24_1_11, A1=>nx10054, B0
      =>que_out_22_1_11, B1=>nx10028);
   ix6675 : nand03 port map ( Y=>nx6674, A0=>nx9039, A1=>nx9041, A2=>nx9043
   );
   ix9040 : aoi222 port map ( Y=>nx9039, A0=>que_out_15_1_11, A1=>nx9976, B0
      =>que_out_3_1_11, B1=>nx10002, C0=>que_out_23_1_11, C1=>nx9950);
   ix9042 : aoi22 port map ( Y=>nx9041, A0=>que_out_27_1_11, A1=>nx9924, B0
      =>que_out_4_1_11, B1=>nx9898);
   ix9044 : aoi22 port map ( Y=>nx9043, A0=>que_out_0_1_11, A1=>nx9846, B0=>
      que_out_2_1_11, B1=>nx9872);
   ix6649 : nand03 port map ( Y=>nx6648, A0=>nx9047, A1=>nx9049, A2=>nx9051
   );
   ix9048 : aoi222 port map ( Y=>nx9047, A0=>que_out_26_1_11, A1=>nx9820, B0
      =>que_out_14_1_11, B1=>nx9794, C0=>que_out_11_1_11, C1=>nx9768);
   ix9050 : aoi22 port map ( Y=>nx9049, A0=>que_out_13_1_11, A1=>nx9742, B0
      =>que_out_7_1_11, B1=>nx9716);
   ix9052 : aoi22 port map ( Y=>nx9051, A0=>que_out_12_1_11, A1=>nx9690, B0
      =>que_out_1_1_11, B1=>nx9664);
   ix6843 : or04 port map ( Y=>out_column_1_12, A0=>nx6838, A1=>nx6812, A2=>
      nx6784, A3=>nx6758);
   ix6839 : nand03 port map ( Y=>nx6838, A0=>nx9057, A1=>nx9059, A2=>nx9061
   );
   ix9058 : aoi222 port map ( Y=>nx9057, A0=>que_out_10_1_12, A1=>nx10314, 
      B0=>que_out_6_1_12, B1=>nx10366, C0=>que_out_9_1_12, C1=>nx10340);
   ix9060 : aoi22 port map ( Y=>nx9059, A0=>que_out_5_1_12, A1=>nx10262, B0
      =>que_out_18_1_12, B1=>nx10288);
   ix9062 : aoi22 port map ( Y=>nx9061, A0=>que_out_17_1_12, A1=>nx10236, B0
      =>que_out_20_1_12, B1=>nx10210);
   ix6813 : nand03 port map ( Y=>nx6812, A0=>nx9065, A1=>nx9067, A2=>nx9069
   );
   ix9066 : aoi222 port map ( Y=>nx9065, A0=>que_out_19_1_12, A1=>nx10184, 
      B0=>que_out_21_1_12, B1=>nx10158, C0=>que_out_8_1_12, C1=>nx10132);
   ix9068 : aoi22 port map ( Y=>nx9067, A0=>que_out_25_1_12, A1=>nx10080, B0
      =>que_out_16_1_12, B1=>nx10106);
   ix9070 : aoi22 port map ( Y=>nx9069, A0=>que_out_24_1_12, A1=>nx10054, B0
      =>que_out_22_1_12, B1=>nx10028);
   ix6785 : nand03 port map ( Y=>nx6784, A0=>nx9073, A1=>nx9075, A2=>nx9077
   );
   ix9074 : aoi222 port map ( Y=>nx9073, A0=>que_out_15_1_12, A1=>nx9976, B0
      =>que_out_3_1_12, B1=>nx10002, C0=>que_out_23_1_12, C1=>nx9950);
   ix9076 : aoi22 port map ( Y=>nx9075, A0=>que_out_27_1_12, A1=>nx9924, B0
      =>que_out_4_1_12, B1=>nx9898);
   ix9078 : aoi22 port map ( Y=>nx9077, A0=>que_out_0_1_12, A1=>nx9846, B0=>
      que_out_2_1_12, B1=>nx9872);
   ix6759 : nand03 port map ( Y=>nx6758, A0=>nx9081, A1=>nx9083, A2=>nx9085
   );
   ix9082 : aoi222 port map ( Y=>nx9081, A0=>que_out_26_1_12, A1=>nx9820, B0
      =>que_out_14_1_12, B1=>nx9794, C0=>que_out_11_1_12, C1=>nx9768);
   ix9084 : aoi22 port map ( Y=>nx9083, A0=>que_out_13_1_12, A1=>nx9742, B0
      =>que_out_7_1_12, B1=>nx9716);
   ix9086 : aoi22 port map ( Y=>nx9085, A0=>que_out_12_1_12, A1=>nx9690, B0
      =>que_out_1_1_12, B1=>nx9664);
   ix6953 : or04 port map ( Y=>out_column_1_13, A0=>nx6948, A1=>nx6922, A2=>
      nx6894, A3=>nx6868);
   ix6949 : nand03 port map ( Y=>nx6948, A0=>nx9090, A1=>nx9093, A2=>nx9095
   );
   ix9092 : aoi222 port map ( Y=>nx9090, A0=>que_out_10_1_13, A1=>nx10314, 
      B0=>que_out_6_1_13, B1=>nx10366, C0=>que_out_9_1_13, C1=>nx10340);
   ix9094 : aoi22 port map ( Y=>nx9093, A0=>que_out_5_1_13, A1=>nx10262, B0
      =>que_out_18_1_13, B1=>nx10288);
   ix9096 : aoi22 port map ( Y=>nx9095, A0=>que_out_17_1_13, A1=>nx10236, B0
      =>que_out_20_1_13, B1=>nx10210);
   ix6923 : nand03 port map ( Y=>nx6922, A0=>nx9098, A1=>nx9101, A2=>nx9103
   );
   ix9100 : aoi222 port map ( Y=>nx9098, A0=>que_out_19_1_13, A1=>nx10184, 
      B0=>que_out_21_1_13, B1=>nx10158, C0=>que_out_8_1_13, C1=>nx10132);
   ix9102 : aoi22 port map ( Y=>nx9101, A0=>que_out_25_1_13, A1=>nx10080, B0
      =>que_out_16_1_13, B1=>nx10106);
   ix9104 : aoi22 port map ( Y=>nx9103, A0=>que_out_24_1_13, A1=>nx10054, B0
      =>que_out_22_1_13, B1=>nx10028);
   ix6895 : nand03 port map ( Y=>nx6894, A0=>nx9106, A1=>nx9108, A2=>nx9110
   );
   ix9107 : aoi222 port map ( Y=>nx9106, A0=>que_out_15_1_13, A1=>nx9976, B0
      =>que_out_3_1_13, B1=>nx10002, C0=>que_out_23_1_13, C1=>nx9950);
   ix9109 : aoi22 port map ( Y=>nx9108, A0=>que_out_27_1_13, A1=>nx9924, B0
      =>que_out_4_1_13, B1=>nx9898);
   ix9111 : aoi22 port map ( Y=>nx9110, A0=>que_out_0_1_13, A1=>nx9846, B0=>
      que_out_2_1_13, B1=>nx9872);
   ix6869 : nand03 port map ( Y=>nx6868, A0=>nx9113, A1=>nx9115, A2=>nx9117
   );
   ix9114 : aoi222 port map ( Y=>nx9113, A0=>que_out_26_1_13, A1=>nx9820, B0
      =>que_out_14_1_13, B1=>nx9794, C0=>que_out_11_1_13, C1=>nx9768);
   ix9116 : aoi22 port map ( Y=>nx9115, A0=>que_out_13_1_13, A1=>nx9742, B0
      =>que_out_7_1_13, B1=>nx9716);
   ix9118 : aoi22 port map ( Y=>nx9117, A0=>que_out_12_1_13, A1=>nx9690, B0
      =>que_out_1_1_13, B1=>nx9664);
   ix7063 : or04 port map ( Y=>out_column_1_14, A0=>nx7058, A1=>nx7032, A2=>
      nx7004, A3=>nx6978);
   ix7059 : nand03 port map ( Y=>nx7058, A0=>nx9121, A1=>nx9123, A2=>nx9125
   );
   ix9122 : aoi222 port map ( Y=>nx9121, A0=>que_out_10_1_14, A1=>nx10314, 
      B0=>que_out_6_1_14, B1=>nx10366, C0=>que_out_9_1_14, C1=>nx10340);
   ix9124 : aoi22 port map ( Y=>nx9123, A0=>que_out_5_1_14, A1=>nx10262, B0
      =>que_out_18_1_14, B1=>nx10288);
   ix9126 : aoi22 port map ( Y=>nx9125, A0=>que_out_17_1_14, A1=>nx10236, B0
      =>que_out_20_1_14, B1=>nx10210);
   ix7033 : nand03 port map ( Y=>nx7032, A0=>nx9128, A1=>nx9130, A2=>nx9132
   );
   ix9129 : aoi222 port map ( Y=>nx9128, A0=>que_out_19_1_14, A1=>nx10184, 
      B0=>que_out_21_1_14, B1=>nx10158, C0=>que_out_8_1_14, C1=>nx10132);
   ix9131 : aoi22 port map ( Y=>nx9130, A0=>que_out_25_1_14, A1=>nx10080, B0
      =>que_out_16_1_14, B1=>nx10106);
   ix9133 : aoi22 port map ( Y=>nx9132, A0=>que_out_24_1_14, A1=>nx10054, B0
      =>que_out_22_1_14, B1=>nx10028);
   ix7005 : nand03 port map ( Y=>nx7004, A0=>nx9135, A1=>nx9137, A2=>nx9139
   );
   ix9136 : aoi222 port map ( Y=>nx9135, A0=>que_out_15_1_14, A1=>nx9976, B0
      =>que_out_3_1_14, B1=>nx10002, C0=>que_out_23_1_14, C1=>nx9950);
   ix9138 : aoi22 port map ( Y=>nx9137, A0=>que_out_27_1_14, A1=>nx9924, B0
      =>que_out_4_1_14, B1=>nx9898);
   ix9140 : aoi22 port map ( Y=>nx9139, A0=>que_out_0_1_14, A1=>nx9846, B0=>
      que_out_2_1_14, B1=>nx9872);
   ix6979 : nand03 port map ( Y=>nx6978, A0=>nx9142, A1=>nx9144, A2=>nx9146
   );
   ix9143 : aoi222 port map ( Y=>nx9142, A0=>que_out_26_1_14, A1=>nx9820, B0
      =>que_out_14_1_14, B1=>nx9794, C0=>que_out_11_1_14, C1=>nx9768);
   ix9145 : aoi22 port map ( Y=>nx9144, A0=>que_out_13_1_14, A1=>nx9742, B0
      =>que_out_7_1_14, B1=>nx9716);
   ix9147 : aoi22 port map ( Y=>nx9146, A0=>que_out_12_1_14, A1=>nx9690, B0
      =>que_out_1_1_14, B1=>nx9664);
   ix7173 : or04 port map ( Y=>out_column_1_15, A0=>nx7168, A1=>nx7142, A2=>
      nx7114, A3=>nx7088);
   ix7169 : nand03 port map ( Y=>nx7168, A0=>nx9150, A1=>nx9152, A2=>nx9154
   );
   ix9151 : aoi222 port map ( Y=>nx9150, A0=>que_out_10_1_15, A1=>nx10316, 
      B0=>que_out_6_1_15, B1=>nx10368, C0=>que_out_9_1_15, C1=>nx10342);
   ix9153 : aoi22 port map ( Y=>nx9152, A0=>que_out_5_1_15, A1=>nx10264, B0
      =>que_out_18_1_15, B1=>nx10290);
   ix9155 : aoi22 port map ( Y=>nx9154, A0=>que_out_17_1_15, A1=>nx10238, B0
      =>que_out_20_1_15, B1=>nx10212);
   ix7143 : nand03 port map ( Y=>nx7142, A0=>nx9157, A1=>nx9159, A2=>nx9161
   );
   ix9158 : aoi222 port map ( Y=>nx9157, A0=>que_out_19_1_15, A1=>nx10186, 
      B0=>que_out_21_1_15, B1=>nx10160, C0=>que_out_8_1_15, C1=>nx10134);
   ix9160 : aoi22 port map ( Y=>nx9159, A0=>que_out_25_1_15, A1=>nx10082, B0
      =>que_out_16_1_15, B1=>nx10108);
   ix9162 : aoi22 port map ( Y=>nx9161, A0=>que_out_24_1_15, A1=>nx10056, B0
      =>que_out_22_1_15, B1=>nx10030);
   ix7115 : nand03 port map ( Y=>nx7114, A0=>nx9164, A1=>nx9166, A2=>nx9168
   );
   ix9165 : aoi222 port map ( Y=>nx9164, A0=>que_out_15_1_15, A1=>nx9978, B0
      =>que_out_3_1_15, B1=>nx10004, C0=>que_out_23_1_15, C1=>nx9952);
   ix9167 : aoi22 port map ( Y=>nx9166, A0=>que_out_27_1_15, A1=>nx9926, B0
      =>que_out_4_1_15, B1=>nx9900);
   ix9169 : aoi22 port map ( Y=>nx9168, A0=>que_out_0_1_15, A1=>nx9848, B0=>
      que_out_2_1_15, B1=>nx9874);
   ix7089 : nand03 port map ( Y=>nx7088, A0=>nx9171, A1=>nx9173, A2=>nx9175
   );
   ix9172 : aoi222 port map ( Y=>nx9171, A0=>que_out_26_1_15, A1=>nx9822, B0
      =>que_out_14_1_15, B1=>nx9796, C0=>que_out_11_1_15, C1=>nx9770);
   ix9174 : aoi22 port map ( Y=>nx9173, A0=>que_out_13_1_15, A1=>nx9744, B0
      =>que_out_7_1_15, B1=>nx9718);
   ix9176 : aoi22 port map ( Y=>nx9175, A0=>que_out_12_1_15, A1=>nx9692, B0
      =>que_out_1_1_15, B1=>nx9666);
   ix7283 : or04 port map ( Y=>out_column_0_0, A0=>nx7278, A1=>nx7252, A2=>
      nx7224, A3=>nx7198);
   ix7279 : nand03 port map ( Y=>nx7278, A0=>nx9179, A1=>nx9181, A2=>nx9183
   );
   ix9180 : aoi222 port map ( Y=>nx9179, A0=>que_out_10_0_0, A1=>nx10316, B0
      =>que_out_6_0_0, B1=>nx10368, C0=>que_out_9_0_0, C1=>nx10342);
   ix9182 : aoi22 port map ( Y=>nx9181, A0=>que_out_5_0_0, A1=>nx10264, B0=>
      que_out_18_0_0, B1=>nx10290);
   ix9184 : aoi22 port map ( Y=>nx9183, A0=>que_out_17_0_0, A1=>nx10238, B0
      =>que_out_20_0_0, B1=>nx10212);
   ix7253 : nand03 port map ( Y=>nx7252, A0=>nx9186, A1=>nx9188, A2=>nx9190
   );
   ix9187 : aoi222 port map ( Y=>nx9186, A0=>que_out_19_0_0, A1=>nx10186, B0
      =>que_out_21_0_0, B1=>nx10160, C0=>que_out_8_0_0, C1=>nx10134);
   ix9189 : aoi22 port map ( Y=>nx9188, A0=>que_out_25_0_0, A1=>nx10082, B0
      =>que_out_16_0_0, B1=>nx10108);
   ix9191 : aoi22 port map ( Y=>nx9190, A0=>que_out_24_0_0, A1=>nx10056, B0
      =>que_out_22_0_0, B1=>nx10030);
   ix7225 : nand03 port map ( Y=>nx7224, A0=>nx9193, A1=>nx9195, A2=>nx9197
   );
   ix9194 : aoi222 port map ( Y=>nx9193, A0=>que_out_15_0_0, A1=>nx9978, B0
      =>que_out_3_0_0, B1=>nx10004, C0=>que_out_23_0_0, C1=>nx9952);
   ix9196 : aoi22 port map ( Y=>nx9195, A0=>que_out_27_0_0, A1=>nx9926, B0=>
      que_out_4_0_0, B1=>nx9900);
   ix9198 : aoi22 port map ( Y=>nx9197, A0=>que_out_0_0_0, A1=>nx9848, B0=>
      que_out_2_0_0, B1=>nx9874);
   ix7199 : nand03 port map ( Y=>nx7198, A0=>nx9200, A1=>nx9202, A2=>nx9204
   );
   ix9201 : aoi222 port map ( Y=>nx9200, A0=>que_out_26_0_0, A1=>nx9822, B0
      =>que_out_14_0_0, B1=>nx9796, C0=>que_out_11_0_0, C1=>nx9770);
   ix9203 : aoi22 port map ( Y=>nx9202, A0=>que_out_13_0_0, A1=>nx9744, B0=>
      que_out_7_0_0, B1=>nx9718);
   ix9205 : aoi22 port map ( Y=>nx9204, A0=>que_out_12_0_0, A1=>nx9692, B0=>
      que_out_1_0_0, B1=>nx9666);
   ix7393 : or04 port map ( Y=>out_column_0_1, A0=>nx7388, A1=>nx7362, A2=>
      nx7334, A3=>nx7308);
   ix7389 : nand03 port map ( Y=>nx7388, A0=>nx9208, A1=>nx9210, A2=>nx9212
   );
   ix9209 : aoi222 port map ( Y=>nx9208, A0=>que_out_10_0_1, A1=>nx10316, B0
      =>que_out_6_0_1, B1=>nx10368, C0=>que_out_9_0_1, C1=>nx10342);
   ix9211 : aoi22 port map ( Y=>nx9210, A0=>que_out_5_0_1, A1=>nx10264, B0=>
      que_out_18_0_1, B1=>nx10290);
   ix9213 : aoi22 port map ( Y=>nx9212, A0=>que_out_17_0_1, A1=>nx10238, B0
      =>que_out_20_0_1, B1=>nx10212);
   ix7363 : nand03 port map ( Y=>nx7362, A0=>nx9215, A1=>nx9217, A2=>nx9219
   );
   ix9216 : aoi222 port map ( Y=>nx9215, A0=>que_out_19_0_1, A1=>nx10186, B0
      =>que_out_21_0_1, B1=>nx10160, C0=>que_out_8_0_1, C1=>nx10134);
   ix9218 : aoi22 port map ( Y=>nx9217, A0=>que_out_25_0_1, A1=>nx10082, B0
      =>que_out_16_0_1, B1=>nx10108);
   ix9220 : aoi22 port map ( Y=>nx9219, A0=>que_out_24_0_1, A1=>nx10056, B0
      =>que_out_22_0_1, B1=>nx10030);
   ix7335 : nand03 port map ( Y=>nx7334, A0=>nx9222, A1=>nx9224, A2=>nx9226
   );
   ix9223 : aoi222 port map ( Y=>nx9222, A0=>que_out_15_0_1, A1=>nx9978, B0
      =>que_out_3_0_1, B1=>nx10004, C0=>que_out_23_0_1, C1=>nx9952);
   ix9225 : aoi22 port map ( Y=>nx9224, A0=>que_out_27_0_1, A1=>nx9926, B0=>
      que_out_4_0_1, B1=>nx9900);
   ix9227 : aoi22 port map ( Y=>nx9226, A0=>que_out_0_0_1, A1=>nx9848, B0=>
      que_out_2_0_1, B1=>nx9874);
   ix7309 : nand03 port map ( Y=>nx7308, A0=>nx9229, A1=>nx9231, A2=>nx9233
   );
   ix9230 : aoi222 port map ( Y=>nx9229, A0=>que_out_26_0_1, A1=>nx9822, B0
      =>que_out_14_0_1, B1=>nx9796, C0=>que_out_11_0_1, C1=>nx9770);
   ix9232 : aoi22 port map ( Y=>nx9231, A0=>que_out_13_0_1, A1=>nx9744, B0=>
      que_out_7_0_1, B1=>nx9718);
   ix9234 : aoi22 port map ( Y=>nx9233, A0=>que_out_12_0_1, A1=>nx9692, B0=>
      que_out_1_0_1, B1=>nx9666);
   ix7503 : or04 port map ( Y=>out_column_0_2, A0=>nx7498, A1=>nx7472, A2=>
      nx7444, A3=>nx7418);
   ix7499 : nand03 port map ( Y=>nx7498, A0=>nx9237, A1=>nx9239, A2=>nx9241
   );
   ix9238 : aoi222 port map ( Y=>nx9237, A0=>que_out_10_0_2, A1=>nx10316, B0
      =>que_out_6_0_2, B1=>nx10368, C0=>que_out_9_0_2, C1=>nx10342);
   ix9240 : aoi22 port map ( Y=>nx9239, A0=>que_out_5_0_2, A1=>nx10264, B0=>
      que_out_18_0_2, B1=>nx10290);
   ix9242 : aoi22 port map ( Y=>nx9241, A0=>que_out_17_0_2, A1=>nx10238, B0
      =>que_out_20_0_2, B1=>nx10212);
   ix7473 : nand03 port map ( Y=>nx7472, A0=>nx9244, A1=>nx9246, A2=>nx9248
   );
   ix9245 : aoi222 port map ( Y=>nx9244, A0=>que_out_19_0_2, A1=>nx10186, B0
      =>que_out_21_0_2, B1=>nx10160, C0=>que_out_8_0_2, C1=>nx10134);
   ix9247 : aoi22 port map ( Y=>nx9246, A0=>que_out_25_0_2, A1=>nx10082, B0
      =>que_out_16_0_2, B1=>nx10108);
   ix9249 : aoi22 port map ( Y=>nx9248, A0=>que_out_24_0_2, A1=>nx10056, B0
      =>que_out_22_0_2, B1=>nx10030);
   ix7445 : nand03 port map ( Y=>nx7444, A0=>nx9251, A1=>nx9253, A2=>nx9255
   );
   ix9252 : aoi222 port map ( Y=>nx9251, A0=>que_out_15_0_2, A1=>nx9978, B0
      =>que_out_3_0_2, B1=>nx10004, C0=>que_out_23_0_2, C1=>nx9952);
   ix9254 : aoi22 port map ( Y=>nx9253, A0=>que_out_27_0_2, A1=>nx9926, B0=>
      que_out_4_0_2, B1=>nx9900);
   ix9256 : aoi22 port map ( Y=>nx9255, A0=>que_out_0_0_2, A1=>nx9848, B0=>
      que_out_2_0_2, B1=>nx9874);
   ix7419 : nand03 port map ( Y=>nx7418, A0=>nx9258, A1=>nx9260, A2=>nx9262
   );
   ix9259 : aoi222 port map ( Y=>nx9258, A0=>que_out_26_0_2, A1=>nx9822, B0
      =>que_out_14_0_2, B1=>nx9796, C0=>que_out_11_0_2, C1=>nx9770);
   ix9261 : aoi22 port map ( Y=>nx9260, A0=>que_out_13_0_2, A1=>nx9744, B0=>
      que_out_7_0_2, B1=>nx9718);
   ix9263 : aoi22 port map ( Y=>nx9262, A0=>que_out_12_0_2, A1=>nx9692, B0=>
      que_out_1_0_2, B1=>nx9666);
   ix7613 : or04 port map ( Y=>out_column_0_3, A0=>nx7608, A1=>nx7582, A2=>
      nx7554, A3=>nx7528);
   ix7609 : nand03 port map ( Y=>nx7608, A0=>nx9266, A1=>nx9268, A2=>nx9270
   );
   ix9267 : aoi222 port map ( Y=>nx9266, A0=>que_out_10_0_3, A1=>nx10316, B0
      =>que_out_6_0_3, B1=>nx10368, C0=>que_out_9_0_3, C1=>nx10342);
   ix9269 : aoi22 port map ( Y=>nx9268, A0=>que_out_5_0_3, A1=>nx10264, B0=>
      que_out_18_0_3, B1=>nx10290);
   ix9271 : aoi22 port map ( Y=>nx9270, A0=>que_out_17_0_3, A1=>nx10238, B0
      =>que_out_20_0_3, B1=>nx10212);
   ix7583 : nand03 port map ( Y=>nx7582, A0=>nx9273, A1=>nx9275, A2=>nx9277
   );
   ix9274 : aoi222 port map ( Y=>nx9273, A0=>que_out_19_0_3, A1=>nx10186, B0
      =>que_out_21_0_3, B1=>nx10160, C0=>que_out_8_0_3, C1=>nx10134);
   ix9276 : aoi22 port map ( Y=>nx9275, A0=>que_out_25_0_3, A1=>nx10082, B0
      =>que_out_16_0_3, B1=>nx10108);
   ix9278 : aoi22 port map ( Y=>nx9277, A0=>que_out_24_0_3, A1=>nx10056, B0
      =>que_out_22_0_3, B1=>nx10030);
   ix7555 : nand03 port map ( Y=>nx7554, A0=>nx9280, A1=>nx9282, A2=>nx9284
   );
   ix9281 : aoi222 port map ( Y=>nx9280, A0=>que_out_15_0_3, A1=>nx9978, B0
      =>que_out_3_0_3, B1=>nx10004, C0=>que_out_23_0_3, C1=>nx9952);
   ix9283 : aoi22 port map ( Y=>nx9282, A0=>que_out_27_0_3, A1=>nx9926, B0=>
      que_out_4_0_3, B1=>nx9900);
   ix9285 : aoi22 port map ( Y=>nx9284, A0=>que_out_0_0_3, A1=>nx9848, B0=>
      que_out_2_0_3, B1=>nx9874);
   ix7529 : nand03 port map ( Y=>nx7528, A0=>nx9287, A1=>nx9289, A2=>nx9291
   );
   ix9288 : aoi222 port map ( Y=>nx9287, A0=>que_out_26_0_3, A1=>nx9822, B0
      =>que_out_14_0_3, B1=>nx9796, C0=>que_out_11_0_3, C1=>nx9770);
   ix9290 : aoi22 port map ( Y=>nx9289, A0=>que_out_13_0_3, A1=>nx9744, B0=>
      que_out_7_0_3, B1=>nx9718);
   ix9292 : aoi22 port map ( Y=>nx9291, A0=>que_out_12_0_3, A1=>nx9692, B0=>
      que_out_1_0_3, B1=>nx9666);
   ix7723 : or04 port map ( Y=>out_column_0_4, A0=>nx7718, A1=>nx7692, A2=>
      nx7664, A3=>nx7638);
   ix7719 : nand03 port map ( Y=>nx7718, A0=>nx9295, A1=>nx9297, A2=>nx9299
   );
   ix9296 : aoi222 port map ( Y=>nx9295, A0=>que_out_10_0_4, A1=>nx10316, B0
      =>que_out_6_0_4, B1=>nx10368, C0=>que_out_9_0_4, C1=>nx10342);
   ix9298 : aoi22 port map ( Y=>nx9297, A0=>que_out_5_0_4, A1=>nx10264, B0=>
      que_out_18_0_4, B1=>nx10290);
   ix9300 : aoi22 port map ( Y=>nx9299, A0=>que_out_17_0_4, A1=>nx10238, B0
      =>que_out_20_0_4, B1=>nx10212);
   ix7693 : nand03 port map ( Y=>nx7692, A0=>nx9302, A1=>nx9304, A2=>nx9306
   );
   ix9303 : aoi222 port map ( Y=>nx9302, A0=>que_out_19_0_4, A1=>nx10186, B0
      =>que_out_21_0_4, B1=>nx10160, C0=>que_out_8_0_4, C1=>nx10134);
   ix9305 : aoi22 port map ( Y=>nx9304, A0=>que_out_25_0_4, A1=>nx10082, B0
      =>que_out_16_0_4, B1=>nx10108);
   ix9307 : aoi22 port map ( Y=>nx9306, A0=>que_out_24_0_4, A1=>nx10056, B0
      =>que_out_22_0_4, B1=>nx10030);
   ix7665 : nand03 port map ( Y=>nx7664, A0=>nx9309, A1=>nx9311, A2=>nx9313
   );
   ix9310 : aoi222 port map ( Y=>nx9309, A0=>que_out_15_0_4, A1=>nx9978, B0
      =>que_out_3_0_4, B1=>nx10004, C0=>que_out_23_0_4, C1=>nx9952);
   ix9312 : aoi22 port map ( Y=>nx9311, A0=>que_out_27_0_4, A1=>nx9926, B0=>
      que_out_4_0_4, B1=>nx9900);
   ix9314 : aoi22 port map ( Y=>nx9313, A0=>que_out_0_0_4, A1=>nx9848, B0=>
      que_out_2_0_4, B1=>nx9874);
   ix7639 : nand03 port map ( Y=>nx7638, A0=>nx9316, A1=>nx9318, A2=>nx9320
   );
   ix9317 : aoi222 port map ( Y=>nx9316, A0=>que_out_26_0_4, A1=>nx9822, B0
      =>que_out_14_0_4, B1=>nx9796, C0=>que_out_11_0_4, C1=>nx9770);
   ix9319 : aoi22 port map ( Y=>nx9318, A0=>que_out_13_0_4, A1=>nx9744, B0=>
      que_out_7_0_4, B1=>nx9718);
   ix9321 : aoi22 port map ( Y=>nx9320, A0=>que_out_12_0_4, A1=>nx9692, B0=>
      que_out_1_0_4, B1=>nx9666);
   ix7833 : or04 port map ( Y=>out_column_0_5, A0=>nx7828, A1=>nx7802, A2=>
      nx7774, A3=>nx7748);
   ix7829 : nand03 port map ( Y=>nx7828, A0=>nx9324, A1=>nx9326, A2=>nx9328
   );
   ix9325 : aoi222 port map ( Y=>nx9324, A0=>que_out_10_0_5, A1=>nx10316, B0
      =>que_out_6_0_5, B1=>nx10368, C0=>que_out_9_0_5, C1=>nx10342);
   ix9327 : aoi22 port map ( Y=>nx9326, A0=>que_out_5_0_5, A1=>nx10264, B0=>
      que_out_18_0_5, B1=>nx10290);
   ix9329 : aoi22 port map ( Y=>nx9328, A0=>que_out_17_0_5, A1=>nx10238, B0
      =>que_out_20_0_5, B1=>nx10212);
   ix7803 : nand03 port map ( Y=>nx7802, A0=>nx9331, A1=>nx9333, A2=>nx9335
   );
   ix9332 : aoi222 port map ( Y=>nx9331, A0=>que_out_19_0_5, A1=>nx10186, B0
      =>que_out_21_0_5, B1=>nx10160, C0=>que_out_8_0_5, C1=>nx10134);
   ix9334 : aoi22 port map ( Y=>nx9333, A0=>que_out_25_0_5, A1=>nx10082, B0
      =>que_out_16_0_5, B1=>nx10108);
   ix9336 : aoi22 port map ( Y=>nx9335, A0=>que_out_24_0_5, A1=>nx10056, B0
      =>que_out_22_0_5, B1=>nx10030);
   ix7775 : nand03 port map ( Y=>nx7774, A0=>nx9338, A1=>nx9340, A2=>nx9342
   );
   ix9339 : aoi222 port map ( Y=>nx9338, A0=>que_out_15_0_5, A1=>nx9978, B0
      =>que_out_3_0_5, B1=>nx10004, C0=>que_out_23_0_5, C1=>nx9952);
   ix9341 : aoi22 port map ( Y=>nx9340, A0=>que_out_27_0_5, A1=>nx9926, B0=>
      que_out_4_0_5, B1=>nx9900);
   ix9343 : aoi22 port map ( Y=>nx9342, A0=>que_out_0_0_5, A1=>nx9848, B0=>
      que_out_2_0_5, B1=>nx9874);
   ix7749 : nand03 port map ( Y=>nx7748, A0=>nx9345, A1=>nx9347, A2=>nx9349
   );
   ix9346 : aoi222 port map ( Y=>nx9345, A0=>que_out_26_0_5, A1=>nx9822, B0
      =>que_out_14_0_5, B1=>nx9796, C0=>que_out_11_0_5, C1=>nx9770);
   ix9348 : aoi22 port map ( Y=>nx9347, A0=>que_out_13_0_5, A1=>nx9744, B0=>
      que_out_7_0_5, B1=>nx9718);
   ix9350 : aoi22 port map ( Y=>nx9349, A0=>que_out_12_0_5, A1=>nx9692, B0=>
      que_out_1_0_5, B1=>nx9666);
   ix7943 : or04 port map ( Y=>out_column_0_6, A0=>nx7938, A1=>nx7912, A2=>
      nx7884, A3=>nx7858);
   ix7939 : nand03 port map ( Y=>nx7938, A0=>nx9353, A1=>nx9355, A2=>nx9357
   );
   ix9354 : aoi222 port map ( Y=>nx9353, A0=>que_out_10_0_6, A1=>nx10318, B0
      =>que_out_6_0_6, B1=>nx10370, C0=>que_out_9_0_6, C1=>nx10344);
   ix9356 : aoi22 port map ( Y=>nx9355, A0=>que_out_5_0_6, A1=>nx10266, B0=>
      que_out_18_0_6, B1=>nx10292);
   ix9358 : aoi22 port map ( Y=>nx9357, A0=>que_out_17_0_6, A1=>nx10240, B0
      =>que_out_20_0_6, B1=>nx10214);
   ix7913 : nand03 port map ( Y=>nx7912, A0=>nx9360, A1=>nx9362, A2=>nx9364
   );
   ix9361 : aoi222 port map ( Y=>nx9360, A0=>que_out_19_0_6, A1=>nx10188, B0
      =>que_out_21_0_6, B1=>nx10162, C0=>que_out_8_0_6, C1=>nx10136);
   ix9363 : aoi22 port map ( Y=>nx9362, A0=>que_out_25_0_6, A1=>nx10084, B0
      =>que_out_16_0_6, B1=>nx10110);
   ix9365 : aoi22 port map ( Y=>nx9364, A0=>que_out_24_0_6, A1=>nx10058, B0
      =>que_out_22_0_6, B1=>nx10032);
   ix7885 : nand03 port map ( Y=>nx7884, A0=>nx9367, A1=>nx9369, A2=>nx9371
   );
   ix9368 : aoi222 port map ( Y=>nx9367, A0=>que_out_15_0_6, A1=>nx9980, B0
      =>que_out_3_0_6, B1=>nx10006, C0=>que_out_23_0_6, C1=>nx9954);
   ix9370 : aoi22 port map ( Y=>nx9369, A0=>que_out_27_0_6, A1=>nx9928, B0=>
      que_out_4_0_6, B1=>nx9902);
   ix9372 : aoi22 port map ( Y=>nx9371, A0=>que_out_0_0_6, A1=>nx9850, B0=>
      que_out_2_0_6, B1=>nx9876);
   ix7859 : nand03 port map ( Y=>nx7858, A0=>nx9374, A1=>nx9376, A2=>nx9378
   );
   ix9375 : aoi222 port map ( Y=>nx9374, A0=>que_out_26_0_6, A1=>nx9824, B0
      =>que_out_14_0_6, B1=>nx9798, C0=>que_out_11_0_6, C1=>nx9772);
   ix9377 : aoi22 port map ( Y=>nx9376, A0=>que_out_13_0_6, A1=>nx9746, B0=>
      que_out_7_0_6, B1=>nx9720);
   ix9379 : aoi22 port map ( Y=>nx9378, A0=>que_out_12_0_6, A1=>nx9694, B0=>
      que_out_1_0_6, B1=>nx9668);
   ix8053 : or04 port map ( Y=>out_column_0_7, A0=>nx8048, A1=>nx8022, A2=>
      nx7994, A3=>nx7968);
   ix8049 : nand03 port map ( Y=>nx8048, A0=>nx9382, A1=>nx9384, A2=>nx9386
   );
   ix9383 : aoi222 port map ( Y=>nx9382, A0=>que_out_10_0_7, A1=>nx10318, B0
      =>que_out_6_0_7, B1=>nx10370, C0=>que_out_9_0_7, C1=>nx10344);
   ix9385 : aoi22 port map ( Y=>nx9384, A0=>que_out_5_0_7, A1=>nx10266, B0=>
      que_out_18_0_7, B1=>nx10292);
   ix9387 : aoi22 port map ( Y=>nx9386, A0=>que_out_17_0_7, A1=>nx10240, B0
      =>que_out_20_0_7, B1=>nx10214);
   ix8023 : nand03 port map ( Y=>nx8022, A0=>nx9389, A1=>nx9391, A2=>nx9393
   );
   ix9390 : aoi222 port map ( Y=>nx9389, A0=>que_out_19_0_7, A1=>nx10188, B0
      =>que_out_21_0_7, B1=>nx10162, C0=>que_out_8_0_7, C1=>nx10136);
   ix9392 : aoi22 port map ( Y=>nx9391, A0=>que_out_25_0_7, A1=>nx10084, B0
      =>que_out_16_0_7, B1=>nx10110);
   ix9394 : aoi22 port map ( Y=>nx9393, A0=>que_out_24_0_7, A1=>nx10058, B0
      =>que_out_22_0_7, B1=>nx10032);
   ix7995 : nand03 port map ( Y=>nx7994, A0=>nx9396, A1=>nx9398, A2=>nx9400
   );
   ix9397 : aoi222 port map ( Y=>nx9396, A0=>que_out_15_0_7, A1=>nx9980, B0
      =>que_out_3_0_7, B1=>nx10006, C0=>que_out_23_0_7, C1=>nx9954);
   ix9399 : aoi22 port map ( Y=>nx9398, A0=>que_out_27_0_7, A1=>nx9928, B0=>
      que_out_4_0_7, B1=>nx9902);
   ix9401 : aoi22 port map ( Y=>nx9400, A0=>que_out_0_0_7, A1=>nx9850, B0=>
      que_out_2_0_7, B1=>nx9876);
   ix7969 : nand03 port map ( Y=>nx7968, A0=>nx9403, A1=>nx9405, A2=>nx9407
   );
   ix9404 : aoi222 port map ( Y=>nx9403, A0=>que_out_26_0_7, A1=>nx9824, B0
      =>que_out_14_0_7, B1=>nx9798, C0=>que_out_11_0_7, C1=>nx9772);
   ix9406 : aoi22 port map ( Y=>nx9405, A0=>que_out_13_0_7, A1=>nx9746, B0=>
      que_out_7_0_7, B1=>nx9720);
   ix9408 : aoi22 port map ( Y=>nx9407, A0=>que_out_12_0_7, A1=>nx9694, B0=>
      que_out_1_0_7, B1=>nx9668);
   ix8163 : or04 port map ( Y=>out_column_0_8, A0=>nx8158, A1=>nx8132, A2=>
      nx8104, A3=>nx8078);
   ix8159 : nand03 port map ( Y=>nx8158, A0=>nx9411, A1=>nx9413, A2=>nx9415
   );
   ix9412 : aoi222 port map ( Y=>nx9411, A0=>que_out_10_0_8, A1=>nx10318, B0
      =>que_out_6_0_8, B1=>nx10370, C0=>que_out_9_0_8, C1=>nx10344);
   ix9414 : aoi22 port map ( Y=>nx9413, A0=>que_out_5_0_8, A1=>nx10266, B0=>
      que_out_18_0_8, B1=>nx10292);
   ix9416 : aoi22 port map ( Y=>nx9415, A0=>que_out_17_0_8, A1=>nx10240, B0
      =>que_out_20_0_8, B1=>nx10214);
   ix8133 : nand03 port map ( Y=>nx8132, A0=>nx9418, A1=>nx9420, A2=>nx9422
   );
   ix9419 : aoi222 port map ( Y=>nx9418, A0=>que_out_19_0_8, A1=>nx10188, B0
      =>que_out_21_0_8, B1=>nx10162, C0=>que_out_8_0_8, C1=>nx10136);
   ix9421 : aoi22 port map ( Y=>nx9420, A0=>que_out_25_0_8, A1=>nx10084, B0
      =>que_out_16_0_8, B1=>nx10110);
   ix9423 : aoi22 port map ( Y=>nx9422, A0=>que_out_24_0_8, A1=>nx10058, B0
      =>que_out_22_0_8, B1=>nx10032);
   ix8105 : nand03 port map ( Y=>nx8104, A0=>nx9425, A1=>nx9427, A2=>nx9429
   );
   ix9426 : aoi222 port map ( Y=>nx9425, A0=>que_out_15_0_8, A1=>nx9980, B0
      =>que_out_3_0_8, B1=>nx10006, C0=>que_out_23_0_8, C1=>nx9954);
   ix9428 : aoi22 port map ( Y=>nx9427, A0=>que_out_27_0_8, A1=>nx9928, B0=>
      que_out_4_0_8, B1=>nx9902);
   ix9430 : aoi22 port map ( Y=>nx9429, A0=>que_out_0_0_8, A1=>nx9850, B0=>
      que_out_2_0_8, B1=>nx9876);
   ix8079 : nand03 port map ( Y=>nx8078, A0=>nx9432, A1=>nx9434, A2=>nx9436
   );
   ix9433 : aoi222 port map ( Y=>nx9432, A0=>que_out_26_0_8, A1=>nx9824, B0
      =>que_out_14_0_8, B1=>nx9798, C0=>que_out_11_0_8, C1=>nx9772);
   ix9435 : aoi22 port map ( Y=>nx9434, A0=>que_out_13_0_8, A1=>nx9746, B0=>
      que_out_7_0_8, B1=>nx9720);
   ix9437 : aoi22 port map ( Y=>nx9436, A0=>que_out_12_0_8, A1=>nx9694, B0=>
      que_out_1_0_8, B1=>nx9668);
   ix8273 : or04 port map ( Y=>out_column_0_9, A0=>nx8268, A1=>nx8242, A2=>
      nx8214, A3=>nx8188);
   ix8269 : nand03 port map ( Y=>nx8268, A0=>nx9440, A1=>nx9442, A2=>nx9444
   );
   ix9441 : aoi222 port map ( Y=>nx9440, A0=>que_out_10_0_9, A1=>nx10318, B0
      =>que_out_6_0_9, B1=>nx10370, C0=>que_out_9_0_9, C1=>nx10344);
   ix9443 : aoi22 port map ( Y=>nx9442, A0=>que_out_5_0_9, A1=>nx10266, B0=>
      que_out_18_0_9, B1=>nx10292);
   ix9445 : aoi22 port map ( Y=>nx9444, A0=>que_out_17_0_9, A1=>nx10240, B0
      =>que_out_20_0_9, B1=>nx10214);
   ix8243 : nand03 port map ( Y=>nx8242, A0=>nx9447, A1=>nx9449, A2=>nx9451
   );
   ix9448 : aoi222 port map ( Y=>nx9447, A0=>que_out_19_0_9, A1=>nx10188, B0
      =>que_out_21_0_9, B1=>nx10162, C0=>que_out_8_0_9, C1=>nx10136);
   ix9450 : aoi22 port map ( Y=>nx9449, A0=>que_out_25_0_9, A1=>nx10084, B0
      =>que_out_16_0_9, B1=>nx10110);
   ix9452 : aoi22 port map ( Y=>nx9451, A0=>que_out_24_0_9, A1=>nx10058, B0
      =>que_out_22_0_9, B1=>nx10032);
   ix8215 : nand03 port map ( Y=>nx8214, A0=>nx9454, A1=>nx9456, A2=>nx9458
   );
   ix9455 : aoi222 port map ( Y=>nx9454, A0=>que_out_15_0_9, A1=>nx9980, B0
      =>que_out_3_0_9, B1=>nx10006, C0=>que_out_23_0_9, C1=>nx9954);
   ix9457 : aoi22 port map ( Y=>nx9456, A0=>que_out_27_0_9, A1=>nx9928, B0=>
      que_out_4_0_9, B1=>nx9902);
   ix9459 : aoi22 port map ( Y=>nx9458, A0=>que_out_0_0_9, A1=>nx9850, B0=>
      que_out_2_0_9, B1=>nx9876);
   ix8189 : nand03 port map ( Y=>nx8188, A0=>nx9461, A1=>nx9463, A2=>nx9465
   );
   ix9462 : aoi222 port map ( Y=>nx9461, A0=>que_out_26_0_9, A1=>nx9824, B0
      =>que_out_14_0_9, B1=>nx9798, C0=>que_out_11_0_9, C1=>nx9772);
   ix9464 : aoi22 port map ( Y=>nx9463, A0=>que_out_13_0_9, A1=>nx9746, B0=>
      que_out_7_0_9, B1=>nx9720);
   ix9466 : aoi22 port map ( Y=>nx9465, A0=>que_out_12_0_9, A1=>nx9694, B0=>
      que_out_1_0_9, B1=>nx9668);
   ix8383 : or04 port map ( Y=>out_column_0_10, A0=>nx8378, A1=>nx8352, A2=>
      nx8324, A3=>nx8298);
   ix8379 : nand03 port map ( Y=>nx8378, A0=>nx9469, A1=>nx9471, A2=>nx9473
   );
   ix9470 : aoi222 port map ( Y=>nx9469, A0=>que_out_10_0_10, A1=>nx10318, 
      B0=>que_out_6_0_10, B1=>nx10370, C0=>que_out_9_0_10, C1=>nx10344);
   ix9472 : aoi22 port map ( Y=>nx9471, A0=>que_out_5_0_10, A1=>nx10266, B0
      =>que_out_18_0_10, B1=>nx10292);
   ix9474 : aoi22 port map ( Y=>nx9473, A0=>que_out_17_0_10, A1=>nx10240, B0
      =>que_out_20_0_10, B1=>nx10214);
   ix8353 : nand03 port map ( Y=>nx8352, A0=>nx9476, A1=>nx9478, A2=>nx9480
   );
   ix9477 : aoi222 port map ( Y=>nx9476, A0=>que_out_19_0_10, A1=>nx10188, 
      B0=>que_out_21_0_10, B1=>nx10162, C0=>que_out_8_0_10, C1=>nx10136);
   ix9479 : aoi22 port map ( Y=>nx9478, A0=>que_out_25_0_10, A1=>nx10084, B0
      =>que_out_16_0_10, B1=>nx10110);
   ix9481 : aoi22 port map ( Y=>nx9480, A0=>que_out_24_0_10, A1=>nx10058, B0
      =>que_out_22_0_10, B1=>nx10032);
   ix8325 : nand03 port map ( Y=>nx8324, A0=>nx9483, A1=>nx9485, A2=>nx9487
   );
   ix9484 : aoi222 port map ( Y=>nx9483, A0=>que_out_15_0_10, A1=>nx9980, B0
      =>que_out_3_0_10, B1=>nx10006, C0=>que_out_23_0_10, C1=>nx9954);
   ix9486 : aoi22 port map ( Y=>nx9485, A0=>que_out_27_0_10, A1=>nx9928, B0
      =>que_out_4_0_10, B1=>nx9902);
   ix9488 : aoi22 port map ( Y=>nx9487, A0=>que_out_0_0_10, A1=>nx9850, B0=>
      que_out_2_0_10, B1=>nx9876);
   ix8299 : nand03 port map ( Y=>nx8298, A0=>nx9490, A1=>nx9492, A2=>nx9494
   );
   ix9491 : aoi222 port map ( Y=>nx9490, A0=>que_out_26_0_10, A1=>nx9824, B0
      =>que_out_14_0_10, B1=>nx9798, C0=>que_out_11_0_10, C1=>nx9772);
   ix9493 : aoi22 port map ( Y=>nx9492, A0=>que_out_13_0_10, A1=>nx9746, B0
      =>que_out_7_0_10, B1=>nx9720);
   ix9495 : aoi22 port map ( Y=>nx9494, A0=>que_out_12_0_10, A1=>nx9694, B0
      =>que_out_1_0_10, B1=>nx9668);
   ix8493 : or04 port map ( Y=>out_column_0_11, A0=>nx8488, A1=>nx8462, A2=>
      nx8434, A3=>nx8408);
   ix8489 : nand03 port map ( Y=>nx8488, A0=>nx9498, A1=>nx9500, A2=>nx9502
   );
   ix9499 : aoi222 port map ( Y=>nx9498, A0=>que_out_10_0_11, A1=>nx10318, 
      B0=>que_out_6_0_11, B1=>nx10370, C0=>que_out_9_0_11, C1=>nx10344);
   ix9501 : aoi22 port map ( Y=>nx9500, A0=>que_out_5_0_11, A1=>nx10266, B0
      =>que_out_18_0_11, B1=>nx10292);
   ix9503 : aoi22 port map ( Y=>nx9502, A0=>que_out_17_0_11, A1=>nx10240, B0
      =>que_out_20_0_11, B1=>nx10214);
   ix8463 : nand03 port map ( Y=>nx8462, A0=>nx9505, A1=>nx9507, A2=>nx9509
   );
   ix9506 : aoi222 port map ( Y=>nx9505, A0=>que_out_19_0_11, A1=>nx10188, 
      B0=>que_out_21_0_11, B1=>nx10162, C0=>que_out_8_0_11, C1=>nx10136);
   ix9508 : aoi22 port map ( Y=>nx9507, A0=>que_out_25_0_11, A1=>nx10084, B0
      =>que_out_16_0_11, B1=>nx10110);
   ix9510 : aoi22 port map ( Y=>nx9509, A0=>que_out_24_0_11, A1=>nx10058, B0
      =>que_out_22_0_11, B1=>nx10032);
   ix8435 : nand03 port map ( Y=>nx8434, A0=>nx9512, A1=>nx9514, A2=>nx9516
   );
   ix9513 : aoi222 port map ( Y=>nx9512, A0=>que_out_15_0_11, A1=>nx9980, B0
      =>que_out_3_0_11, B1=>nx10006, C0=>que_out_23_0_11, C1=>nx9954);
   ix9515 : aoi22 port map ( Y=>nx9514, A0=>que_out_27_0_11, A1=>nx9928, B0
      =>que_out_4_0_11, B1=>nx9902);
   ix9517 : aoi22 port map ( Y=>nx9516, A0=>que_out_0_0_11, A1=>nx9850, B0=>
      que_out_2_0_11, B1=>nx9876);
   ix8409 : nand03 port map ( Y=>nx8408, A0=>nx9519, A1=>nx9521, A2=>nx9523
   );
   ix9520 : aoi222 port map ( Y=>nx9519, A0=>que_out_26_0_11, A1=>nx9824, B0
      =>que_out_14_0_11, B1=>nx9798, C0=>que_out_11_0_11, C1=>nx9772);
   ix9522 : aoi22 port map ( Y=>nx9521, A0=>que_out_13_0_11, A1=>nx9746, B0
      =>que_out_7_0_11, B1=>nx9720);
   ix9524 : aoi22 port map ( Y=>nx9523, A0=>que_out_12_0_11, A1=>nx9694, B0
      =>que_out_1_0_11, B1=>nx9668);
   ix8603 : or04 port map ( Y=>out_column_0_12, A0=>nx8598, A1=>nx8572, A2=>
      nx8544, A3=>nx8518);
   ix8599 : nand03 port map ( Y=>nx8598, A0=>nx9527, A1=>nx9529, A2=>nx9531
   );
   ix9528 : aoi222 port map ( Y=>nx9527, A0=>que_out_10_0_12, A1=>nx10318, 
      B0=>que_out_6_0_12, B1=>nx10370, C0=>que_out_9_0_12, C1=>nx10344);
   ix9530 : aoi22 port map ( Y=>nx9529, A0=>que_out_5_0_12, A1=>nx10266, B0
      =>que_out_18_0_12, B1=>nx10292);
   ix9532 : aoi22 port map ( Y=>nx9531, A0=>que_out_17_0_12, A1=>nx10240, B0
      =>que_out_20_0_12, B1=>nx10214);
   ix8573 : nand03 port map ( Y=>nx8572, A0=>nx9534, A1=>nx9536, A2=>nx9538
   );
   ix9535 : aoi222 port map ( Y=>nx9534, A0=>que_out_19_0_12, A1=>nx10188, 
      B0=>que_out_21_0_12, B1=>nx10162, C0=>que_out_8_0_12, C1=>nx10136);
   ix9537 : aoi22 port map ( Y=>nx9536, A0=>que_out_25_0_12, A1=>nx10084, B0
      =>que_out_16_0_12, B1=>nx10110);
   ix9539 : aoi22 port map ( Y=>nx9538, A0=>que_out_24_0_12, A1=>nx10058, B0
      =>que_out_22_0_12, B1=>nx10032);
   ix8545 : nand03 port map ( Y=>nx8544, A0=>nx9541, A1=>nx9543, A2=>nx9545
   );
   ix9542 : aoi222 port map ( Y=>nx9541, A0=>que_out_15_0_12, A1=>nx9980, B0
      =>que_out_3_0_12, B1=>nx10006, C0=>que_out_23_0_12, C1=>nx9954);
   ix9544 : aoi22 port map ( Y=>nx9543, A0=>que_out_27_0_12, A1=>nx9928, B0
      =>que_out_4_0_12, B1=>nx9902);
   ix9546 : aoi22 port map ( Y=>nx9545, A0=>que_out_0_0_12, A1=>nx9850, B0=>
      que_out_2_0_12, B1=>nx9876);
   ix8519 : nand03 port map ( Y=>nx8518, A0=>nx9548, A1=>nx9550, A2=>nx9552
   );
   ix9549 : aoi222 port map ( Y=>nx9548, A0=>que_out_26_0_12, A1=>nx9824, B0
      =>que_out_14_0_12, B1=>nx9798, C0=>que_out_11_0_12, C1=>nx9772);
   ix9551 : aoi22 port map ( Y=>nx9550, A0=>que_out_13_0_12, A1=>nx9746, B0
      =>que_out_7_0_12, B1=>nx9720);
   ix9553 : aoi22 port map ( Y=>nx9552, A0=>que_out_12_0_12, A1=>nx9694, B0
      =>que_out_1_0_12, B1=>nx9668);
   ix8713 : or04 port map ( Y=>out_column_0_13, A0=>nx8708, A1=>nx8682, A2=>
      nx8654, A3=>nx8628);
   ix8709 : nand03 port map ( Y=>nx8708, A0=>nx9556, A1=>nx9558, A2=>nx9560
   );
   ix9557 : aoi222 port map ( Y=>nx9556, A0=>que_out_10_0_13, A1=>nx10320, 
      B0=>que_out_6_0_13, B1=>nx10372, C0=>que_out_9_0_13, C1=>nx10346);
   ix9559 : aoi22 port map ( Y=>nx9558, A0=>que_out_5_0_13, A1=>nx10268, B0
      =>que_out_18_0_13, B1=>nx10294);
   ix9561 : aoi22 port map ( Y=>nx9560, A0=>que_out_17_0_13, A1=>nx10242, B0
      =>que_out_20_0_13, B1=>nx10216);
   ix8683 : nand03 port map ( Y=>nx8682, A0=>nx9563, A1=>nx9565, A2=>nx9567
   );
   ix9564 : aoi222 port map ( Y=>nx9563, A0=>que_out_19_0_13, A1=>nx10190, 
      B0=>que_out_21_0_13, B1=>nx10164, C0=>que_out_8_0_13, C1=>nx10138);
   ix9566 : aoi22 port map ( Y=>nx9565, A0=>que_out_25_0_13, A1=>nx10086, B0
      =>que_out_16_0_13, B1=>nx10112);
   ix9568 : aoi22 port map ( Y=>nx9567, A0=>que_out_24_0_13, A1=>nx10060, B0
      =>que_out_22_0_13, B1=>nx10034);
   ix8655 : nand03 port map ( Y=>nx8654, A0=>nx9570, A1=>nx9572, A2=>nx9574
   );
   ix9571 : aoi222 port map ( Y=>nx9570, A0=>que_out_15_0_13, A1=>nx9982, B0
      =>que_out_3_0_13, B1=>nx10008, C0=>que_out_23_0_13, C1=>nx9956);
   ix9573 : aoi22 port map ( Y=>nx9572, A0=>que_out_27_0_13, A1=>nx9930, B0
      =>que_out_4_0_13, B1=>nx9904);
   ix9575 : aoi22 port map ( Y=>nx9574, A0=>que_out_0_0_13, A1=>nx9852, B0=>
      que_out_2_0_13, B1=>nx9878);
   ix8629 : nand03 port map ( Y=>nx8628, A0=>nx9577, A1=>nx9579, A2=>nx9581
   );
   ix9578 : aoi222 port map ( Y=>nx9577, A0=>que_out_26_0_13, A1=>nx9826, B0
      =>que_out_14_0_13, B1=>nx9800, C0=>que_out_11_0_13, C1=>nx9774);
   ix9580 : aoi22 port map ( Y=>nx9579, A0=>que_out_13_0_13, A1=>nx9748, B0
      =>que_out_7_0_13, B1=>nx9722);
   ix9582 : aoi22 port map ( Y=>nx9581, A0=>que_out_12_0_13, A1=>nx9696, B0
      =>que_out_1_0_13, B1=>nx9670);
   ix8823 : or04 port map ( Y=>out_column_0_14, A0=>nx8818, A1=>nx8792, A2=>
      nx8764, A3=>nx8738);
   ix8819 : nand03 port map ( Y=>nx8818, A0=>nx9585, A1=>nx9587, A2=>nx9589
   );
   ix9586 : aoi222 port map ( Y=>nx9585, A0=>que_out_10_0_14, A1=>nx10320, 
      B0=>que_out_6_0_14, B1=>nx10372, C0=>que_out_9_0_14, C1=>nx10346);
   ix9588 : aoi22 port map ( Y=>nx9587, A0=>que_out_5_0_14, A1=>nx10268, B0
      =>que_out_18_0_14, B1=>nx10294);
   ix9590 : aoi22 port map ( Y=>nx9589, A0=>que_out_17_0_14, A1=>nx10242, B0
      =>que_out_20_0_14, B1=>nx10216);
   ix8793 : nand03 port map ( Y=>nx8792, A0=>nx9592, A1=>nx9594, A2=>nx9596
   );
   ix9593 : aoi222 port map ( Y=>nx9592, A0=>que_out_19_0_14, A1=>nx10190, 
      B0=>que_out_21_0_14, B1=>nx10164, C0=>que_out_8_0_14, C1=>nx10138);
   ix9595 : aoi22 port map ( Y=>nx9594, A0=>que_out_25_0_14, A1=>nx10086, B0
      =>que_out_16_0_14, B1=>nx10112);
   ix9597 : aoi22 port map ( Y=>nx9596, A0=>que_out_24_0_14, A1=>nx10060, B0
      =>que_out_22_0_14, B1=>nx10034);
   ix8765 : nand03 port map ( Y=>nx8764, A0=>nx9599, A1=>nx9601, A2=>nx9603
   );
   ix9600 : aoi222 port map ( Y=>nx9599, A0=>que_out_15_0_14, A1=>nx9982, B0
      =>que_out_3_0_14, B1=>nx10008, C0=>que_out_23_0_14, C1=>nx9956);
   ix9602 : aoi22 port map ( Y=>nx9601, A0=>que_out_27_0_14, A1=>nx9930, B0
      =>que_out_4_0_14, B1=>nx9904);
   ix9604 : aoi22 port map ( Y=>nx9603, A0=>que_out_0_0_14, A1=>nx9852, B0=>
      que_out_2_0_14, B1=>nx9878);
   ix8739 : nand03 port map ( Y=>nx8738, A0=>nx9606, A1=>nx9608, A2=>nx9610
   );
   ix9607 : aoi222 port map ( Y=>nx9606, A0=>que_out_26_0_14, A1=>nx9826, B0
      =>que_out_14_0_14, B1=>nx9800, C0=>que_out_11_0_14, C1=>nx9774);
   ix9609 : aoi22 port map ( Y=>nx9608, A0=>que_out_13_0_14, A1=>nx9748, B0
      =>que_out_7_0_14, B1=>nx9722);
   ix9611 : aoi22 port map ( Y=>nx9610, A0=>que_out_12_0_14, A1=>nx9696, B0
      =>que_out_1_0_14, B1=>nx9670);
   ix8933 : or04 port map ( Y=>out_column_0_15, A0=>nx8928, A1=>nx8902, A2=>
      nx8874, A3=>nx8848);
   ix8929 : nand03 port map ( Y=>nx8928, A0=>nx9614, A1=>nx9616, A2=>nx9618
   );
   ix9615 : aoi222 port map ( Y=>nx9614, A0=>que_out_10_0_15, A1=>nx10320, 
      B0=>que_out_6_0_15, B1=>nx10372, C0=>que_out_9_0_15, C1=>nx10346);
   ix9617 : aoi22 port map ( Y=>nx9616, A0=>que_out_5_0_15, A1=>nx10268, B0
      =>que_out_18_0_15, B1=>nx10294);
   ix9619 : aoi22 port map ( Y=>nx9618, A0=>que_out_17_0_15, A1=>nx10242, B0
      =>que_out_20_0_15, B1=>nx10216);
   ix8903 : nand03 port map ( Y=>nx8902, A0=>nx9621, A1=>nx9623, A2=>nx9625
   );
   ix9622 : aoi222 port map ( Y=>nx9621, A0=>que_out_19_0_15, A1=>nx10190, 
      B0=>que_out_21_0_15, B1=>nx10164, C0=>que_out_8_0_15, C1=>nx10138);
   ix9624 : aoi22 port map ( Y=>nx9623, A0=>que_out_25_0_15, A1=>nx10086, B0
      =>que_out_16_0_15, B1=>nx10112);
   ix9626 : aoi22 port map ( Y=>nx9625, A0=>que_out_24_0_15, A1=>nx10060, B0
      =>que_out_22_0_15, B1=>nx10034);
   ix8875 : nand03 port map ( Y=>nx8874, A0=>nx9628, A1=>nx9630, A2=>nx9632
   );
   ix9629 : aoi222 port map ( Y=>nx9628, A0=>que_out_15_0_15, A1=>nx9982, B0
      =>que_out_3_0_15, B1=>nx10008, C0=>que_out_23_0_15, C1=>nx9956);
   ix9631 : aoi22 port map ( Y=>nx9630, A0=>que_out_27_0_15, A1=>nx9930, B0
      =>que_out_4_0_15, B1=>nx9904);
   ix9633 : aoi22 port map ( Y=>nx9632, A0=>que_out_0_0_15, A1=>nx9852, B0=>
      que_out_2_0_15, B1=>nx9878);
   ix8849 : nand03 port map ( Y=>nx8848, A0=>nx9635, A1=>nx9637, A2=>nx9639
   );
   ix9636 : aoi222 port map ( Y=>nx9635, A0=>que_out_26_0_15, A1=>nx9826, B0
      =>que_out_14_0_15, B1=>nx9800, C0=>que_out_11_0_15, C1=>nx9774);
   ix9638 : aoi22 port map ( Y=>nx9637, A0=>que_out_13_0_15, A1=>nx9748, B0
      =>que_out_7_0_15, B1=>nx9722);
   ix9640 : aoi22 port map ( Y=>nx9639, A0=>que_out_12_0_15, A1=>nx9696, B0
      =>que_out_1_0_15, B1=>nx9670);
   ix6944 : inv02 port map ( Y=>nx6943, A=>nx88);
   ix9647 : inv02 port map ( Y=>nx9648, A=>nx10378);
   ix9649 : inv02 port map ( Y=>nx9650, A=>nx10378);
   ix9651 : inv02 port map ( Y=>nx9652, A=>nx10378);
   ix9653 : inv02 port map ( Y=>nx9654, A=>nx10378);
   ix9655 : inv02 port map ( Y=>nx9656, A=>nx10378);
   ix9657 : inv02 port map ( Y=>nx9658, A=>nx10378);
   ix9659 : inv02 port map ( Y=>nx9660, A=>nx10378);
   ix9661 : inv02 port map ( Y=>nx9662, A=>nx10380);
   ix9663 : inv02 port map ( Y=>nx9664, A=>nx10380);
   ix9665 : inv02 port map ( Y=>nx9666, A=>nx10380);
   ix9667 : inv02 port map ( Y=>nx9668, A=>nx10380);
   ix9669 : inv02 port map ( Y=>nx9670, A=>nx10380);
   ix9673 : inv02 port map ( Y=>nx9674, A=>nx10382);
   ix9675 : inv02 port map ( Y=>nx9676, A=>nx10382);
   ix9677 : inv02 port map ( Y=>nx9678, A=>nx10382);
   ix9679 : inv02 port map ( Y=>nx9680, A=>nx10382);
   ix9681 : inv02 port map ( Y=>nx9682, A=>nx10382);
   ix9683 : inv02 port map ( Y=>nx9684, A=>nx10382);
   ix9685 : inv02 port map ( Y=>nx9686, A=>nx10382);
   ix9687 : inv02 port map ( Y=>nx9688, A=>nx10384);
   ix9689 : inv02 port map ( Y=>nx9690, A=>nx10384);
   ix9691 : inv02 port map ( Y=>nx9692, A=>nx10384);
   ix9693 : inv02 port map ( Y=>nx9694, A=>nx10384);
   ix9695 : inv02 port map ( Y=>nx9696, A=>nx10384);
   ix9699 : inv02 port map ( Y=>nx9700, A=>nx10386);
   ix9701 : inv02 port map ( Y=>nx9702, A=>nx10386);
   ix9703 : inv02 port map ( Y=>nx9704, A=>nx10386);
   ix9705 : inv02 port map ( Y=>nx9706, A=>nx10386);
   ix9707 : inv02 port map ( Y=>nx9708, A=>nx10386);
   ix9709 : inv02 port map ( Y=>nx9710, A=>nx10386);
   ix9711 : inv02 port map ( Y=>nx9712, A=>nx10386);
   ix9713 : inv02 port map ( Y=>nx9714, A=>nx10388);
   ix9715 : inv02 port map ( Y=>nx9716, A=>nx10388);
   ix9717 : inv02 port map ( Y=>nx9718, A=>nx10388);
   ix9719 : inv02 port map ( Y=>nx9720, A=>nx10388);
   ix9721 : inv02 port map ( Y=>nx9722, A=>nx10388);
   ix9725 : inv02 port map ( Y=>nx9726, A=>nx10390);
   ix9727 : inv02 port map ( Y=>nx9728, A=>nx10390);
   ix9729 : inv02 port map ( Y=>nx9730, A=>nx10390);
   ix9731 : inv02 port map ( Y=>nx9732, A=>nx10390);
   ix9733 : inv02 port map ( Y=>nx9734, A=>nx10390);
   ix9735 : inv02 port map ( Y=>nx9736, A=>nx10390);
   ix9737 : inv02 port map ( Y=>nx9738, A=>nx10390);
   ix9739 : inv02 port map ( Y=>nx9740, A=>nx10392);
   ix9741 : inv02 port map ( Y=>nx9742, A=>nx10392);
   ix9743 : inv02 port map ( Y=>nx9744, A=>nx10392);
   ix9745 : inv02 port map ( Y=>nx9746, A=>nx10392);
   ix9747 : inv02 port map ( Y=>nx9748, A=>nx10392);
   ix9751 : inv02 port map ( Y=>nx9752, A=>nx10394);
   ix9753 : inv02 port map ( Y=>nx9754, A=>nx10394);
   ix9755 : inv02 port map ( Y=>nx9756, A=>nx10394);
   ix9757 : inv02 port map ( Y=>nx9758, A=>nx10394);
   ix9759 : inv02 port map ( Y=>nx9760, A=>nx10394);
   ix9761 : inv02 port map ( Y=>nx9762, A=>nx10394);
   ix9763 : inv02 port map ( Y=>nx9764, A=>nx10394);
   ix9765 : inv02 port map ( Y=>nx9766, A=>nx10396);
   ix9767 : inv02 port map ( Y=>nx9768, A=>nx10396);
   ix9769 : inv02 port map ( Y=>nx9770, A=>nx10396);
   ix9771 : inv02 port map ( Y=>nx9772, A=>nx10396);
   ix9773 : inv02 port map ( Y=>nx9774, A=>nx10396);
   ix9777 : inv02 port map ( Y=>nx9778, A=>nx10398);
   ix9779 : inv02 port map ( Y=>nx9780, A=>nx10398);
   ix9781 : inv02 port map ( Y=>nx9782, A=>nx10398);
   ix9783 : inv02 port map ( Y=>nx9784, A=>nx10398);
   ix9785 : inv02 port map ( Y=>nx9786, A=>nx10398);
   ix9787 : inv02 port map ( Y=>nx9788, A=>nx10398);
   ix9789 : inv02 port map ( Y=>nx9790, A=>nx10398);
   ix9791 : inv02 port map ( Y=>nx9792, A=>nx10400);
   ix9793 : inv02 port map ( Y=>nx9794, A=>nx10400);
   ix9795 : inv02 port map ( Y=>nx9796, A=>nx10400);
   ix9797 : inv02 port map ( Y=>nx9798, A=>nx10400);
   ix9799 : inv02 port map ( Y=>nx9800, A=>nx10400);
   ix9803 : inv02 port map ( Y=>nx9804, A=>nx10402);
   ix9805 : inv02 port map ( Y=>nx9806, A=>nx10402);
   ix9807 : inv02 port map ( Y=>nx9808, A=>nx10402);
   ix9809 : inv02 port map ( Y=>nx9810, A=>nx10402);
   ix9811 : inv02 port map ( Y=>nx9812, A=>nx10402);
   ix9813 : inv02 port map ( Y=>nx9814, A=>nx10402);
   ix9815 : inv02 port map ( Y=>nx9816, A=>nx10402);
   ix9817 : inv02 port map ( Y=>nx9818, A=>nx10404);
   ix9819 : inv02 port map ( Y=>nx9820, A=>nx10404);
   ix9821 : inv02 port map ( Y=>nx9822, A=>nx10404);
   ix9823 : inv02 port map ( Y=>nx9824, A=>nx10404);
   ix9825 : inv02 port map ( Y=>nx9826, A=>nx10404);
   ix9829 : inv02 port map ( Y=>nx9830, A=>nx10406);
   ix9831 : inv02 port map ( Y=>nx9832, A=>nx10406);
   ix9833 : inv02 port map ( Y=>nx9834, A=>nx10406);
   ix9835 : inv02 port map ( Y=>nx9836, A=>nx10406);
   ix9837 : inv02 port map ( Y=>nx9838, A=>nx10406);
   ix9839 : inv02 port map ( Y=>nx9840, A=>nx10406);
   ix9841 : inv02 port map ( Y=>nx9842, A=>nx10406);
   ix9843 : inv02 port map ( Y=>nx9844, A=>nx10408);
   ix9845 : inv02 port map ( Y=>nx9846, A=>nx10408);
   ix9847 : inv02 port map ( Y=>nx9848, A=>nx10408);
   ix9849 : inv02 port map ( Y=>nx9850, A=>nx10408);
   ix9851 : inv02 port map ( Y=>nx9852, A=>nx10408);
   ix9855 : inv02 port map ( Y=>nx9856, A=>nx10410);
   ix9857 : inv02 port map ( Y=>nx9858, A=>nx10410);
   ix9859 : inv02 port map ( Y=>nx9860, A=>nx10410);
   ix9861 : inv02 port map ( Y=>nx9862, A=>nx10410);
   ix9863 : inv02 port map ( Y=>nx9864, A=>nx10410);
   ix9865 : inv02 port map ( Y=>nx9866, A=>nx10410);
   ix9867 : inv02 port map ( Y=>nx9868, A=>nx10410);
   ix9869 : inv02 port map ( Y=>nx9870, A=>nx10412);
   ix9871 : inv02 port map ( Y=>nx9872, A=>nx10412);
   ix9873 : inv02 port map ( Y=>nx9874, A=>nx10412);
   ix9875 : inv02 port map ( Y=>nx9876, A=>nx10412);
   ix9877 : inv02 port map ( Y=>nx9878, A=>nx10412);
   ix9881 : inv02 port map ( Y=>nx9882, A=>nx10414);
   ix9883 : inv02 port map ( Y=>nx9884, A=>nx10414);
   ix9885 : inv02 port map ( Y=>nx9886, A=>nx10414);
   ix9887 : inv02 port map ( Y=>nx9888, A=>nx10414);
   ix9889 : inv02 port map ( Y=>nx9890, A=>nx10414);
   ix9891 : inv02 port map ( Y=>nx9892, A=>nx10414);
   ix9893 : inv02 port map ( Y=>nx9894, A=>nx10414);
   ix9895 : inv02 port map ( Y=>nx9896, A=>nx10416);
   ix9897 : inv02 port map ( Y=>nx9898, A=>nx10416);
   ix9899 : inv02 port map ( Y=>nx9900, A=>nx10416);
   ix9901 : inv02 port map ( Y=>nx9902, A=>nx10416);
   ix9903 : inv02 port map ( Y=>nx9904, A=>nx10416);
   ix9907 : inv02 port map ( Y=>nx9908, A=>nx10418);
   ix9909 : inv02 port map ( Y=>nx9910, A=>nx10418);
   ix9911 : inv02 port map ( Y=>nx9912, A=>nx10418);
   ix9913 : inv02 port map ( Y=>nx9914, A=>nx10418);
   ix9915 : inv02 port map ( Y=>nx9916, A=>nx10418);
   ix9917 : inv02 port map ( Y=>nx9918, A=>nx10418);
   ix9919 : inv02 port map ( Y=>nx9920, A=>nx10418);
   ix9921 : inv02 port map ( Y=>nx9922, A=>nx10420);
   ix9923 : inv02 port map ( Y=>nx9924, A=>nx10420);
   ix9925 : inv02 port map ( Y=>nx9926, A=>nx10420);
   ix9927 : inv02 port map ( Y=>nx9928, A=>nx10420);
   ix9929 : inv02 port map ( Y=>nx9930, A=>nx10420);
   ix9933 : inv02 port map ( Y=>nx9934, A=>nx10422);
   ix9935 : inv02 port map ( Y=>nx9936, A=>nx10422);
   ix9937 : inv02 port map ( Y=>nx9938, A=>nx10422);
   ix9939 : inv02 port map ( Y=>nx9940, A=>nx10422);
   ix9941 : inv02 port map ( Y=>nx9942, A=>nx10422);
   ix9943 : inv02 port map ( Y=>nx9944, A=>nx10422);
   ix9945 : inv02 port map ( Y=>nx9946, A=>nx10422);
   ix9947 : inv02 port map ( Y=>nx9948, A=>nx10424);
   ix9949 : inv02 port map ( Y=>nx9950, A=>nx10424);
   ix9951 : inv02 port map ( Y=>nx9952, A=>nx10424);
   ix9953 : inv02 port map ( Y=>nx9954, A=>nx10424);
   ix9955 : inv02 port map ( Y=>nx9956, A=>nx10424);
   ix9959 : inv02 port map ( Y=>nx9960, A=>nx10426);
   ix9961 : inv02 port map ( Y=>nx9962, A=>nx10426);
   ix9963 : inv02 port map ( Y=>nx9964, A=>nx10426);
   ix9965 : inv02 port map ( Y=>nx9966, A=>nx10426);
   ix9967 : inv02 port map ( Y=>nx9968, A=>nx10426);
   ix9969 : inv02 port map ( Y=>nx9970, A=>nx10426);
   ix9971 : inv02 port map ( Y=>nx9972, A=>nx10426);
   ix9973 : inv02 port map ( Y=>nx9974, A=>nx10428);
   ix9975 : inv02 port map ( Y=>nx9976, A=>nx10428);
   ix9977 : inv02 port map ( Y=>nx9978, A=>nx10428);
   ix9979 : inv02 port map ( Y=>nx9980, A=>nx10428);
   ix9981 : inv02 port map ( Y=>nx9982, A=>nx10428);
   ix9985 : inv02 port map ( Y=>nx9986, A=>nx10430);
   ix9987 : inv02 port map ( Y=>nx9988, A=>nx10430);
   ix9989 : inv02 port map ( Y=>nx9990, A=>nx10430);
   ix9991 : inv02 port map ( Y=>nx9992, A=>nx10430);
   ix9993 : inv02 port map ( Y=>nx9994, A=>nx10430);
   ix9995 : inv02 port map ( Y=>nx9996, A=>nx10430);
   ix9997 : inv02 port map ( Y=>nx9998, A=>nx10430);
   ix9999 : inv02 port map ( Y=>nx10000, A=>nx10432);
   ix10001 : inv02 port map ( Y=>nx10002, A=>nx10432);
   ix10003 : inv02 port map ( Y=>nx10004, A=>nx10432);
   ix10005 : inv02 port map ( Y=>nx10006, A=>nx10432);
   ix10007 : inv02 port map ( Y=>nx10008, A=>nx10432);
   ix10011 : inv02 port map ( Y=>nx10012, A=>nx10434);
   ix10013 : inv02 port map ( Y=>nx10014, A=>nx10434);
   ix10015 : inv02 port map ( Y=>nx10016, A=>nx10434);
   ix10017 : inv02 port map ( Y=>nx10018, A=>nx10434);
   ix10019 : inv02 port map ( Y=>nx10020, A=>nx10434);
   ix10021 : inv02 port map ( Y=>nx10022, A=>nx10434);
   ix10023 : inv02 port map ( Y=>nx10024, A=>nx10434);
   ix10025 : inv02 port map ( Y=>nx10026, A=>nx10436);
   ix10027 : inv02 port map ( Y=>nx10028, A=>nx10436);
   ix10029 : inv02 port map ( Y=>nx10030, A=>nx10436);
   ix10031 : inv02 port map ( Y=>nx10032, A=>nx10436);
   ix10033 : inv02 port map ( Y=>nx10034, A=>nx10436);
   ix10037 : inv02 port map ( Y=>nx10038, A=>nx10438);
   ix10039 : inv02 port map ( Y=>nx10040, A=>nx10438);
   ix10041 : inv02 port map ( Y=>nx10042, A=>nx10438);
   ix10043 : inv02 port map ( Y=>nx10044, A=>nx10438);
   ix10045 : inv02 port map ( Y=>nx10046, A=>nx10438);
   ix10047 : inv02 port map ( Y=>nx10048, A=>nx10438);
   ix10049 : inv02 port map ( Y=>nx10050, A=>nx10438);
   ix10051 : inv02 port map ( Y=>nx10052, A=>nx10440);
   ix10053 : inv02 port map ( Y=>nx10054, A=>nx10440);
   ix10055 : inv02 port map ( Y=>nx10056, A=>nx10440);
   ix10057 : inv02 port map ( Y=>nx10058, A=>nx10440);
   ix10059 : inv02 port map ( Y=>nx10060, A=>nx10440);
   ix10063 : inv02 port map ( Y=>nx10064, A=>nx10442);
   ix10065 : inv02 port map ( Y=>nx10066, A=>nx10442);
   ix10067 : inv02 port map ( Y=>nx10068, A=>nx10442);
   ix10069 : inv02 port map ( Y=>nx10070, A=>nx10442);
   ix10071 : inv02 port map ( Y=>nx10072, A=>nx10442);
   ix10073 : inv02 port map ( Y=>nx10074, A=>nx10442);
   ix10075 : inv02 port map ( Y=>nx10076, A=>nx10442);
   ix10077 : inv02 port map ( Y=>nx10078, A=>nx10444);
   ix10079 : inv02 port map ( Y=>nx10080, A=>nx10444);
   ix10081 : inv02 port map ( Y=>nx10082, A=>nx10444);
   ix10083 : inv02 port map ( Y=>nx10084, A=>nx10444);
   ix10085 : inv02 port map ( Y=>nx10086, A=>nx10444);
   ix10089 : inv02 port map ( Y=>nx10090, A=>nx10446);
   ix10091 : inv02 port map ( Y=>nx10092, A=>nx10446);
   ix10093 : inv02 port map ( Y=>nx10094, A=>nx10446);
   ix10095 : inv02 port map ( Y=>nx10096, A=>nx10446);
   ix10097 : inv02 port map ( Y=>nx10098, A=>nx10446);
   ix10099 : inv02 port map ( Y=>nx10100, A=>nx10446);
   ix10101 : inv02 port map ( Y=>nx10102, A=>nx10446);
   ix10103 : inv02 port map ( Y=>nx10104, A=>nx10448);
   ix10105 : inv02 port map ( Y=>nx10106, A=>nx10448);
   ix10107 : inv02 port map ( Y=>nx10108, A=>nx10448);
   ix10109 : inv02 port map ( Y=>nx10110, A=>nx10448);
   ix10111 : inv02 port map ( Y=>nx10112, A=>nx10448);
   ix10115 : inv02 port map ( Y=>nx10116, A=>nx10450);
   ix10117 : inv02 port map ( Y=>nx10118, A=>nx10450);
   ix10119 : inv02 port map ( Y=>nx10120, A=>nx10450);
   ix10121 : inv02 port map ( Y=>nx10122, A=>nx10450);
   ix10123 : inv02 port map ( Y=>nx10124, A=>nx10450);
   ix10125 : inv02 port map ( Y=>nx10126, A=>nx10450);
   ix10127 : inv02 port map ( Y=>nx10128, A=>nx10450);
   ix10129 : inv02 port map ( Y=>nx10130, A=>nx10452);
   ix10131 : inv02 port map ( Y=>nx10132, A=>nx10452);
   ix10133 : inv02 port map ( Y=>nx10134, A=>nx10452);
   ix10135 : inv02 port map ( Y=>nx10136, A=>nx10452);
   ix10137 : inv02 port map ( Y=>nx10138, A=>nx10452);
   ix10141 : inv02 port map ( Y=>nx10142, A=>nx10454);
   ix10143 : inv02 port map ( Y=>nx10144, A=>nx10454);
   ix10145 : inv02 port map ( Y=>nx10146, A=>nx10454);
   ix10147 : inv02 port map ( Y=>nx10148, A=>nx10454);
   ix10149 : inv02 port map ( Y=>nx10150, A=>nx10454);
   ix10151 : inv02 port map ( Y=>nx10152, A=>nx10454);
   ix10153 : inv02 port map ( Y=>nx10154, A=>nx10454);
   ix10155 : inv02 port map ( Y=>nx10156, A=>nx10456);
   ix10157 : inv02 port map ( Y=>nx10158, A=>nx10456);
   ix10159 : inv02 port map ( Y=>nx10160, A=>nx10456);
   ix10161 : inv02 port map ( Y=>nx10162, A=>nx10456);
   ix10163 : inv02 port map ( Y=>nx10164, A=>nx10456);
   ix10167 : inv02 port map ( Y=>nx10168, A=>nx10458);
   ix10169 : inv02 port map ( Y=>nx10170, A=>nx10458);
   ix10171 : inv02 port map ( Y=>nx10172, A=>nx10458);
   ix10173 : inv02 port map ( Y=>nx10174, A=>nx10458);
   ix10175 : inv02 port map ( Y=>nx10176, A=>nx10458);
   ix10177 : inv02 port map ( Y=>nx10178, A=>nx10458);
   ix10179 : inv02 port map ( Y=>nx10180, A=>nx10458);
   ix10181 : inv02 port map ( Y=>nx10182, A=>nx10460);
   ix10183 : inv02 port map ( Y=>nx10184, A=>nx10460);
   ix10185 : inv02 port map ( Y=>nx10186, A=>nx10460);
   ix10187 : inv02 port map ( Y=>nx10188, A=>nx10460);
   ix10189 : inv02 port map ( Y=>nx10190, A=>nx10460);
   ix10193 : inv02 port map ( Y=>nx10194, A=>nx10462);
   ix10195 : inv02 port map ( Y=>nx10196, A=>nx10462);
   ix10197 : inv02 port map ( Y=>nx10198, A=>nx10462);
   ix10199 : inv02 port map ( Y=>nx10200, A=>nx10462);
   ix10201 : inv02 port map ( Y=>nx10202, A=>nx10462);
   ix10203 : inv02 port map ( Y=>nx10204, A=>nx10462);
   ix10205 : inv02 port map ( Y=>nx10206, A=>nx10462);
   ix10207 : inv02 port map ( Y=>nx10208, A=>nx10464);
   ix10209 : inv02 port map ( Y=>nx10210, A=>nx10464);
   ix10211 : inv02 port map ( Y=>nx10212, A=>nx10464);
   ix10213 : inv02 port map ( Y=>nx10214, A=>nx10464);
   ix10215 : inv02 port map ( Y=>nx10216, A=>nx10464);
   ix10219 : inv02 port map ( Y=>nx10220, A=>nx10466);
   ix10221 : inv02 port map ( Y=>nx10222, A=>nx10466);
   ix10223 : inv02 port map ( Y=>nx10224, A=>nx10466);
   ix10225 : inv02 port map ( Y=>nx10226, A=>nx10466);
   ix10227 : inv02 port map ( Y=>nx10228, A=>nx10466);
   ix10229 : inv02 port map ( Y=>nx10230, A=>nx10466);
   ix10231 : inv02 port map ( Y=>nx10232, A=>nx10466);
   ix10233 : inv02 port map ( Y=>nx10234, A=>nx10468);
   ix10235 : inv02 port map ( Y=>nx10236, A=>nx10468);
   ix10237 : inv02 port map ( Y=>nx10238, A=>nx10468);
   ix10239 : inv02 port map ( Y=>nx10240, A=>nx10468);
   ix10241 : inv02 port map ( Y=>nx10242, A=>nx10468);
   ix10245 : inv02 port map ( Y=>nx10246, A=>nx10470);
   ix10247 : inv02 port map ( Y=>nx10248, A=>nx10470);
   ix10249 : inv02 port map ( Y=>nx10250, A=>nx10470);
   ix10251 : inv02 port map ( Y=>nx10252, A=>nx10470);
   ix10253 : inv02 port map ( Y=>nx10254, A=>nx10470);
   ix10255 : inv02 port map ( Y=>nx10256, A=>nx10470);
   ix10257 : inv02 port map ( Y=>nx10258, A=>nx10470);
   ix10259 : inv02 port map ( Y=>nx10260, A=>nx10472);
   ix10261 : inv02 port map ( Y=>nx10262, A=>nx10472);
   ix10263 : inv02 port map ( Y=>nx10264, A=>nx10472);
   ix10265 : inv02 port map ( Y=>nx10266, A=>nx10472);
   ix10267 : inv02 port map ( Y=>nx10268, A=>nx10472);
   ix10271 : inv02 port map ( Y=>nx10272, A=>nx10474);
   ix10273 : inv02 port map ( Y=>nx10274, A=>nx10474);
   ix10275 : inv02 port map ( Y=>nx10276, A=>nx10474);
   ix10277 : inv02 port map ( Y=>nx10278, A=>nx10474);
   ix10279 : inv02 port map ( Y=>nx10280, A=>nx10474);
   ix10281 : inv02 port map ( Y=>nx10282, A=>nx10474);
   ix10283 : inv02 port map ( Y=>nx10284, A=>nx10474);
   ix10285 : inv02 port map ( Y=>nx10286, A=>nx10476);
   ix10287 : inv02 port map ( Y=>nx10288, A=>nx10476);
   ix10289 : inv02 port map ( Y=>nx10290, A=>nx10476);
   ix10291 : inv02 port map ( Y=>nx10292, A=>nx10476);
   ix10293 : inv02 port map ( Y=>nx10294, A=>nx10476);
   ix10297 : inv02 port map ( Y=>nx10298, A=>nx10478);
   ix10299 : inv02 port map ( Y=>nx10300, A=>nx10478);
   ix10301 : inv02 port map ( Y=>nx10302, A=>nx10478);
   ix10303 : inv02 port map ( Y=>nx10304, A=>nx10478);
   ix10305 : inv02 port map ( Y=>nx10306, A=>nx10478);
   ix10307 : inv02 port map ( Y=>nx10308, A=>nx10478);
   ix10309 : inv02 port map ( Y=>nx10310, A=>nx10478);
   ix10311 : inv02 port map ( Y=>nx10312, A=>nx10480);
   ix10313 : inv02 port map ( Y=>nx10314, A=>nx10480);
   ix10315 : inv02 port map ( Y=>nx10316, A=>nx10480);
   ix10317 : inv02 port map ( Y=>nx10318, A=>nx10480);
   ix10319 : inv02 port map ( Y=>nx10320, A=>nx10480);
   ix10323 : inv02 port map ( Y=>nx10324, A=>nx10482);
   ix10325 : inv02 port map ( Y=>nx10326, A=>nx10482);
   ix10327 : inv02 port map ( Y=>nx10328, A=>nx10482);
   ix10329 : inv02 port map ( Y=>nx10330, A=>nx10482);
   ix10331 : inv02 port map ( Y=>nx10332, A=>nx10482);
   ix10333 : inv02 port map ( Y=>nx10334, A=>nx10482);
   ix10335 : inv02 port map ( Y=>nx10336, A=>nx10482);
   ix10337 : inv02 port map ( Y=>nx10338, A=>nx10484);
   ix10339 : inv02 port map ( Y=>nx10340, A=>nx10484);
   ix10341 : inv02 port map ( Y=>nx10342, A=>nx10484);
   ix10343 : inv02 port map ( Y=>nx10344, A=>nx10484);
   ix10345 : inv02 port map ( Y=>nx10346, A=>nx10484);
   ix10349 : inv02 port map ( Y=>nx10350, A=>nx10486);
   ix10351 : inv02 port map ( Y=>nx10352, A=>nx10486);
   ix10353 : inv02 port map ( Y=>nx10354, A=>nx10486);
   ix10355 : inv02 port map ( Y=>nx10356, A=>nx10486);
   ix10357 : inv02 port map ( Y=>nx10358, A=>nx10486);
   ix10359 : inv02 port map ( Y=>nx10360, A=>nx10486);
   ix10361 : inv02 port map ( Y=>nx10362, A=>nx10486);
   ix10363 : inv02 port map ( Y=>nx10364, A=>nx10488);
   ix10365 : inv02 port map ( Y=>nx10366, A=>nx10488);
   ix10367 : inv02 port map ( Y=>nx10368, A=>nx10488);
   ix10369 : inv02 port map ( Y=>nx10370, A=>nx10488);
   ix10371 : inv02 port map ( Y=>nx10372, A=>nx10488);
   ix10373 : buf02 port map ( Y=>nx10374, A=>nx6955);
   ix10375 : buf02 port map ( Y=>nx10376, A=>nx6955);
   ix10377 : inv02 port map ( Y=>nx10378, A=>nx14);
   ix10379 : inv02 port map ( Y=>nx10380, A=>nx14);
   ix10381 : inv02 port map ( Y=>nx10382, A=>nx30);
   ix10383 : inv02 port map ( Y=>nx10384, A=>nx30);
   ix10385 : inv02 port map ( Y=>nx10386, A=>nx42);
   ix10387 : inv02 port map ( Y=>nx10388, A=>nx42);
   ix10389 : inv02 port map ( Y=>nx10390, A=>nx48);
   ix10391 : inv02 port map ( Y=>nx10392, A=>nx48);
   ix10393 : inv02 port map ( Y=>nx10394, A=>nx64);
   ix10395 : inv02 port map ( Y=>nx10396, A=>nx64);
   ix10397 : inv02 port map ( Y=>nx10398, A=>nx68);
   ix10399 : inv02 port map ( Y=>nx10400, A=>nx68);
   ix10401 : inv02 port map ( Y=>nx10402, A=>nx74);
   ix10403 : inv02 port map ( Y=>nx10404, A=>nx74);
   ix10405 : inv02 port map ( Y=>nx10406, A=>nx90);
   ix10407 : inv02 port map ( Y=>nx10408, A=>nx90);
   ix10409 : inv02 port map ( Y=>nx10410, A=>nx94);
   ix10411 : inv02 port map ( Y=>nx10412, A=>nx94);
   ix10413 : inv02 port map ( Y=>nx10414, A=>nx100);
   ix10415 : inv02 port map ( Y=>nx10416, A=>nx100);
   ix10417 : inv02 port map ( Y=>nx10418, A=>nx104);
   ix10419 : inv02 port map ( Y=>nx10420, A=>nx104);
   ix10421 : inv02 port map ( Y=>nx10422, A=>nx114);
   ix10423 : inv02 port map ( Y=>nx10424, A=>nx114);
   ix10425 : inv02 port map ( Y=>nx10426, A=>nx118);
   ix10427 : inv02 port map ( Y=>nx10428, A=>nx118);
   ix10429 : inv02 port map ( Y=>nx10430, A=>nx122);
   ix10431 : inv02 port map ( Y=>nx10432, A=>nx122);
   ix10433 : inv02 port map ( Y=>nx10434, A=>nx136);
   ix10435 : inv02 port map ( Y=>nx10436, A=>nx136);
   ix10437 : inv02 port map ( Y=>nx10438, A=>nx144);
   ix10439 : inv02 port map ( Y=>nx10440, A=>nx144);
   ix10441 : inv02 port map ( Y=>nx10442, A=>nx150);
   ix10443 : inv02 port map ( Y=>nx10444, A=>nx150);
   ix10445 : inv02 port map ( Y=>nx10446, A=>nx158);
   ix10447 : inv02 port map ( Y=>nx10448, A=>nx158);
   ix10449 : inv02 port map ( Y=>nx10450, A=>nx166);
   ix10451 : inv02 port map ( Y=>nx10452, A=>nx166);
   ix10453 : inv02 port map ( Y=>nx10454, A=>nx172);
   ix10455 : inv02 port map ( Y=>nx10456, A=>nx172);
   ix10457 : inv02 port map ( Y=>nx10458, A=>nx180);
   ix10459 : inv02 port map ( Y=>nx10460, A=>nx180);
   ix10461 : inv02 port map ( Y=>nx10462, A=>nx192);
   ix10463 : inv02 port map ( Y=>nx10464, A=>nx192);
   ix10465 : inv02 port map ( Y=>nx10466, A=>nx200);
   ix10467 : inv02 port map ( Y=>nx10468, A=>nx200);
   ix10469 : inv02 port map ( Y=>nx10470, A=>nx206);
   ix10471 : inv02 port map ( Y=>nx10472, A=>nx206);
   ix10473 : inv02 port map ( Y=>nx10474, A=>nx214);
   ix10475 : inv02 port map ( Y=>nx10476, A=>nx214);
   ix10477 : inv02 port map ( Y=>nx10478, A=>nx222);
   ix10479 : inv02 port map ( Y=>nx10480, A=>nx222);
   ix10481 : inv02 port map ( Y=>nx10482, A=>nx226);
   ix10483 : inv02 port map ( Y=>nx10484, A=>nx226);
   ix10485 : inv02 port map ( Y=>nx10486, A=>nx230);
   ix10487 : inv02 port map ( Y=>nx10488, A=>nx230);
   ix8951 : nor02ii port map ( Y=>sel_que_0, A0=>nx6829, A1=>nx6885);
   ix8961 : nor02ii port map ( Y=>sel_que_1, A0=>nx6839, A1=>nx6885);
   ix8971 : nor02ii port map ( Y=>sel_que_2, A0=>nx6843, A1=>nx6885);
   ix8979 : nor02ii port map ( Y=>sel_que_3, A0=>nx6847, A1=>nx6885);
   ix8987 : nor02ii port map ( Y=>sel_que_4, A0=>nx6829, A1=>nx6905);
   ix8991 : nor02ii port map ( Y=>sel_que_5, A0=>nx6839, A1=>nx6905);
   ix8995 : nor02ii port map ( Y=>sel_que_6, A0=>nx6843, A1=>nx6905);
   ix8999 : nor02ii port map ( Y=>sel_que_7, A0=>nx6847, A1=>nx6905);
   ix9007 : nor02ii port map ( Y=>sel_que_8, A0=>nx6829, A1=>nx6915);
   ix9011 : nor02ii port map ( Y=>sel_que_9, A0=>nx6839, A1=>nx6915);
   ix9015 : nor02ii port map ( Y=>sel_que_10, A0=>nx6843, A1=>nx6915);
   ix9019 : nor02ii port map ( Y=>sel_que_11, A0=>nx6847, A1=>nx6915);
   ix9053 : nor02ii port map ( Y=>sel_que_17, A0=>nx6893, A1=>nx6885);
   ix9063 : nor02ii port map ( Y=>sel_que_18, A0=>nx6897, A1=>nx6885);
   ix9071 : nor02ii port map ( Y=>sel_que_19, A0=>nx6901, A1=>nx6885);
   ix6906 : nor02ii port map ( Y=>nx6905, A0=>cache_in_sel(3), A1=>
      cache_in_sel(2));
   ix9079 : nor02ii port map ( Y=>sel_que_21, A0=>nx6893, A1=>nx6905);
   ix9083 : nor02ii port map ( Y=>sel_que_22, A0=>nx6897, A1=>nx6905);
   ix9087 : nor02ii port map ( Y=>sel_que_23, A0=>nx6901, A1=>nx6905);
   ix6916 : nor02ii port map ( Y=>nx6915, A0=>cache_in_sel(2), A1=>
      cache_in_sel(3));
   ix9095 : nor02ii port map ( Y=>sel_que_25, A0=>nx6893, A1=>nx6915);
   ix9099 : nor02ii port map ( Y=>sel_que_26, A0=>nx6897, A1=>nx6915);
   ix9103 : nor02ii port map ( Y=>sel_que_27, A0=>nx6901, A1=>nx6915);
   ix223 : nor02ii port map ( Y=>nx222, A0=>nx6931, A1=>nx62);
   ix231 : nor02ii port map ( Y=>nx230, A0=>nx6945, A1=>nx88);
   ix207 : nor02ii port map ( Y=>nx206, A0=>nx10374, A1=>nx28);
   ix123 : nor02ii port map ( Y=>nx122, A0=>nx10374, A1=>nx62);
   ix65 : nor02ii port map ( Y=>nx64, A0=>nx6949, A1=>nx62);
   ix49 : nor02ii port map ( Y=>nx48, A0=>nx6949, A1=>nx28);
   ix31 : nor02ii port map ( Y=>nx30, A0=>nx6931, A1=>nx28);
   ix10493 : inv02 port map ( Y=>nx10494, A=>nx6937);
   ix10495 : inv02 port map ( Y=>nx10496, A=>nx6937);
   ix10497 : inv02 port map ( Y=>nx10498, A=>nx6939);
   ix10499 : inv02 port map ( Y=>nx10500, A=>nx6939);
   ix10501 : inv01 port map ( Y=>nx10502, A=>nx6961);
   ix10503 : inv01 port map ( Y=>nx10504, A=>nx6961);
   ix10505 : inv02 port map ( Y=>nx10506, A=>nx6833);
   ix10507 : inv02 port map ( Y=>nx10508, A=>nx6835);
   ix10509 : inv01 port map ( Y=>nx10510, A=>in_word(15));
   ix10511 : inv01 port map ( Y=>nx10512, A=>nx10510);
   ix10513 : inv01 port map ( Y=>nx10514, A=>nx10510);
   ix10515 : inv01 port map ( Y=>nx10516, A=>nx10510);
   ix10517 : inv01 port map ( Y=>nx10518, A=>nx10510);
   ix10519 : inv01 port map ( Y=>nx10520, A=>in_word(14));
   ix10521 : inv01 port map ( Y=>nx10522, A=>nx10520);
   ix10523 : inv01 port map ( Y=>nx10524, A=>nx10520);
   ix10525 : inv01 port map ( Y=>nx10526, A=>nx10520);
   ix10527 : inv01 port map ( Y=>nx10528, A=>nx10520);
   ix10529 : inv01 port map ( Y=>nx10530, A=>in_word(13));
   ix10531 : inv01 port map ( Y=>nx10532, A=>nx10530);
   ix10533 : inv01 port map ( Y=>nx10534, A=>nx10530);
   ix10535 : inv01 port map ( Y=>nx10536, A=>nx10530);
   ix10537 : inv01 port map ( Y=>nx10538, A=>nx10530);
   ix10539 : inv01 port map ( Y=>nx10540, A=>in_word(12));
   ix10541 : inv01 port map ( Y=>nx10542, A=>nx10540);
   ix10543 : inv01 port map ( Y=>nx10544, A=>nx10540);
   ix10545 : inv01 port map ( Y=>nx10546, A=>nx10540);
   ix10547 : inv01 port map ( Y=>nx10548, A=>nx10540);
   ix10549 : inv01 port map ( Y=>nx10550, A=>in_word(11));
   ix10551 : inv01 port map ( Y=>nx10552, A=>nx10550);
   ix10553 : inv01 port map ( Y=>nx10554, A=>nx10550);
   ix10555 : inv01 port map ( Y=>nx10556, A=>nx10550);
   ix10557 : inv01 port map ( Y=>nx10558, A=>nx10550);
   ix10559 : inv01 port map ( Y=>nx10560, A=>in_word(10));
   ix10561 : inv01 port map ( Y=>nx10562, A=>nx10560);
   ix10563 : inv01 port map ( Y=>nx10564, A=>nx10560);
   ix10565 : inv01 port map ( Y=>nx10566, A=>nx10560);
   ix10567 : inv01 port map ( Y=>nx10568, A=>nx10560);
   ix10569 : inv01 port map ( Y=>nx10570, A=>in_word(9));
   ix10571 : inv01 port map ( Y=>nx10572, A=>nx10570);
   ix10573 : inv01 port map ( Y=>nx10574, A=>nx10570);
   ix10575 : inv01 port map ( Y=>nx10576, A=>nx10570);
   ix10577 : inv01 port map ( Y=>nx10578, A=>nx10570);
   ix10579 : inv01 port map ( Y=>nx10580, A=>in_word(8));
   ix10581 : inv01 port map ( Y=>nx10582, A=>nx10580);
   ix10583 : inv01 port map ( Y=>nx10584, A=>nx10580);
   ix10585 : inv01 port map ( Y=>nx10586, A=>nx10580);
   ix10587 : inv01 port map ( Y=>nx10588, A=>nx10580);
   ix10589 : inv01 port map ( Y=>nx10590, A=>in_word(7));
   ix10591 : inv01 port map ( Y=>nx10592, A=>nx10590);
   ix10593 : inv01 port map ( Y=>nx10594, A=>nx10590);
   ix10595 : inv01 port map ( Y=>nx10596, A=>nx10590);
   ix10597 : inv01 port map ( Y=>nx10598, A=>nx10590);
   ix10599 : inv01 port map ( Y=>nx10600, A=>in_word(6));
   ix10601 : inv01 port map ( Y=>nx10602, A=>nx10600);
   ix10603 : inv01 port map ( Y=>nx10604, A=>nx10600);
   ix10605 : inv01 port map ( Y=>nx10606, A=>nx10600);
   ix10607 : inv01 port map ( Y=>nx10608, A=>nx10600);
   ix10609 : inv01 port map ( Y=>nx10610, A=>in_word(5));
   ix10611 : inv01 port map ( Y=>nx10612, A=>nx10610);
   ix10613 : inv01 port map ( Y=>nx10614, A=>nx10610);
   ix10615 : inv01 port map ( Y=>nx10616, A=>nx10610);
   ix10617 : inv01 port map ( Y=>nx10618, A=>nx10610);
   ix10619 : inv01 port map ( Y=>nx10620, A=>in_word(4));
   ix10621 : inv01 port map ( Y=>nx10622, A=>nx10620);
   ix10623 : inv01 port map ( Y=>nx10624, A=>nx10620);
   ix10625 : inv01 port map ( Y=>nx10626, A=>nx10620);
   ix10627 : inv01 port map ( Y=>nx10628, A=>nx10620);
   ix10629 : inv01 port map ( Y=>nx10630, A=>in_word(3));
   ix10631 : inv01 port map ( Y=>nx10632, A=>nx10630);
   ix10633 : inv01 port map ( Y=>nx10634, A=>nx10630);
   ix10635 : inv01 port map ( Y=>nx10636, A=>nx10630);
   ix10637 : inv01 port map ( Y=>nx10638, A=>nx10630);
   ix10639 : inv01 port map ( Y=>nx10640, A=>in_word(2));
   ix10641 : inv01 port map ( Y=>nx10642, A=>nx10640);
   ix10643 : inv01 port map ( Y=>nx10644, A=>nx10640);
   ix10645 : inv01 port map ( Y=>nx10646, A=>nx10640);
   ix10647 : inv01 port map ( Y=>nx10648, A=>nx10640);
   ix10649 : inv01 port map ( Y=>nx10650, A=>in_word(1));
   ix10651 : inv01 port map ( Y=>nx10652, A=>nx10650);
   ix10653 : inv01 port map ( Y=>nx10654, A=>nx10650);
   ix10655 : inv01 port map ( Y=>nx10656, A=>nx10650);
   ix10657 : inv01 port map ( Y=>nx10658, A=>nx10650);
   ix10659 : inv01 port map ( Y=>nx10660, A=>in_word(0));
   ix10661 : inv01 port map ( Y=>nx10662, A=>nx10660);
   ix10663 : inv01 port map ( Y=>nx10664, A=>nx10660);
   ix10665 : inv01 port map ( Y=>nx10666, A=>nx10660);
   ix10667 : inv01 port map ( Y=>nx10668, A=>nx10660);
   ix10689 : inv02 port map ( Y=>nx10690, A=>nx10742);
   ix10691 : inv02 port map ( Y=>nx10692, A=>nx10742);
   ix10693 : inv02 port map ( Y=>nx10694, A=>nx10742);
   ix10695 : inv02 port map ( Y=>nx10696, A=>nx10742);
   ix10697 : inv02 port map ( Y=>nx10698, A=>nx10742);
   ix10699 : inv02 port map ( Y=>nx10700, A=>nx10742);
   ix10701 : inv02 port map ( Y=>nx10702, A=>nx10742);
   ix10703 : inv02 port map ( Y=>nx10704, A=>nx10744);
   ix10705 : inv02 port map ( Y=>nx10706, A=>nx10744);
   ix10707 : inv02 port map ( Y=>nx10708, A=>nx10744);
   ix10709 : inv02 port map ( Y=>nx10710, A=>nx10744);
   ix10711 : inv02 port map ( Y=>nx10712, A=>nx10744);
   ix10713 : inv02 port map ( Y=>nx10714, A=>nx10746);
   ix10715 : inv02 port map ( Y=>nx10716, A=>nx10746);
   ix10717 : inv02 port map ( Y=>nx10718, A=>nx10746);
   ix10719 : inv02 port map ( Y=>nx10720, A=>nx10746);
   ix10721 : inv02 port map ( Y=>nx10722, A=>nx10746);
   ix10723 : inv02 port map ( Y=>nx10724, A=>nx10746);
   ix10725 : inv02 port map ( Y=>nx10726, A=>nx10746);
   ix10727 : inv02 port map ( Y=>nx10728, A=>nx10748);
   ix10729 : inv02 port map ( Y=>nx10730, A=>nx10748);
   ix10731 : inv02 port map ( Y=>nx10732, A=>nx10748);
   ix10733 : inv02 port map ( Y=>nx10734, A=>nx10748);
   ix10735 : inv02 port map ( Y=>nx10736, A=>nx10748);
   ix10741 : inv02 port map ( Y=>nx10742, A=>reset);
   ix10743 : inv02 port map ( Y=>nx10744, A=>reset);
   ix10745 : inv02 port map ( Y=>nx10746, A=>clk);
   ix10747 : inv02 port map ( Y=>nx10748, A=>clk);
end Dataflow ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity AdvancedCounter_16 is
   port (
      clk : IN std_logic ;
      reset : IN std_logic ;
      enable : IN std_logic ;
      mode_in : IN std_logic_vector (1 DOWNTO 0) ;
      max_val_in : IN std_logic_vector (15 DOWNTO 0) ;
      max_reached_out : OUT std_logic ;
      counter_out : OUT std_logic_vector (15 DOWNTO 0)) ;
end AdvancedCounter_16 ;

architecture behavioural_unfold_2902 of AdvancedCounter_16 is
   signal counter_out_0_EXMPLR, counter_out_15_EXMPLR, counter_out_14_EXMPLR, 
      nx149, counter_out_13_EXMPLR, counter_out_12_EXMPLR, nx152, 
      counter_out_11_EXMPLR, counter_out_10_EXMPLR, nx155, 
      counter_out_9_EXMPLR, counter_out_8_EXMPLR, nx157, 
      counter_out_7_EXMPLR, counter_out_6_EXMPLR, nx159, 
      counter_out_5_EXMPLR, counter_out_4_EXMPLR, nx161, 
      counter_out_3_EXMPLR, counter_out_2_EXMPLR, counter_out_1_EXMPLR, 
      counter_out_dup0_0, nx22, nx34, nx46, nx70, nx94, nx118, nx142, nx166, 
      nx174, nx192, nx206, nx224, nx246, nx173, nx183, nx193, nx203, nx213, 
      nx223, nx233, nx243, nx253, nx263, nx273, nx283, nx293, nx303, nx313, 
      nx323, nx339, nx344, nx348, nx350, nx353, nx358, nx362, nx364, nx367, 
      nx372, nx376, nx378, nx381, nx386, nx390, nx392, nx395, nx400, nx404, 
      nx406, nx409, nx414, nx419, nx424, nx428, nx430, nx436, nx439, nx445, 
      nx447, nx449, nx451, nx458, nx460, nx462, nx464, nx466, nx468, nx470, 
      nx472, nx474: std_logic ;

begin
   counter_out(15) <= counter_out_0_EXMPLR ;
   counter_out(14) <= counter_out_0_EXMPLR ;
   counter_out(13) <= counter_out_0_EXMPLR ;
   counter_out(12) <= counter_out_0_EXMPLR ;
   counter_out(11) <= counter_out_0_EXMPLR ;
   counter_out(10) <= counter_out_0_EXMPLR ;
   counter_out(9) <= counter_out_0_EXMPLR ;
   counter_out(8) <= counter_out_0_EXMPLR ;
   counter_out(7) <= counter_out_0_EXMPLR ;
   counter_out(6) <= counter_out_0_EXMPLR ;
   counter_out(5) <= counter_out_0_EXMPLR ;
   counter_out(4) <= counter_out_0_EXMPLR ;
   counter_out(3) <= counter_out_0_EXMPLR ;
   counter_out(2) <= counter_out_0_EXMPLR ;
   counter_out(1) <= counter_out_0_EXMPLR ;
   counter_out(0) <= counter_out_0_EXMPLR ;
   ix140 : fake_gnd port map ( Y=>counter_out_0_EXMPLR);
   ix251 : and04 port map ( Y=>max_reached_out, A0=>nx192, A1=>nx206, A2=>
      nx224, A3=>nx246);
   ix324 : mux21_ni port map ( Y=>nx323, A0=>counter_out_15_EXMPLR, A1=>
      nx174, S0=>nx474);
   ix314 : mux21_ni port map ( Y=>nx313, A0=>counter_out_14_EXMPLR, A1=>
      nx166, S0=>nx472);
   reg_counter_data_14 : dffr port map ( Q=>counter_out_14_EXMPLR, QB=>nx339, 
      D=>nx313, CLK=>clk, R=>nx462);
   ix345 : nand02 port map ( Y=>nx344, A0=>counter_out_13_EXMPLR, A1=>nx152
   );
   ix304 : mux21 port map ( Y=>nx303, A0=>nx348, A1=>nx350, S0=>nx472);
   reg_counter_data_13 : dffr port map ( Q=>counter_out_13_EXMPLR, QB=>nx348, 
      D=>nx303, CLK=>clk, R=>nx462);
   ix351 : oai21 port map ( Y=>nx350, A0=>nx152, A1=>counter_out_13_EXMPLR, 
      B0=>nx344);
   ix294 : mux21_ni port map ( Y=>nx293, A0=>counter_out_12_EXMPLR, A1=>
      nx142, S0=>nx472);
   reg_counter_data_12 : dffr port map ( Q=>counter_out_12_EXMPLR, QB=>nx353, 
      D=>nx293, CLK=>clk, R=>nx462);
   ix359 : nand02 port map ( Y=>nx358, A0=>counter_out_11_EXMPLR, A1=>nx155
   );
   ix284 : mux21 port map ( Y=>nx283, A0=>nx362, A1=>nx364, S0=>nx472);
   reg_counter_data_11 : dffr port map ( Q=>counter_out_11_EXMPLR, QB=>nx362, 
      D=>nx283, CLK=>clk, R=>nx462);
   ix365 : oai21 port map ( Y=>nx364, A0=>nx155, A1=>counter_out_11_EXMPLR, 
      B0=>nx358);
   ix274 : mux21_ni port map ( Y=>nx273, A0=>counter_out_10_EXMPLR, A1=>
      nx118, S0=>nx472);
   reg_counter_data_10 : dffr port map ( Q=>counter_out_10_EXMPLR, QB=>nx367, 
      D=>nx273, CLK=>clk, R=>nx462);
   ix373 : nand02 port map ( Y=>nx372, A0=>counter_out_9_EXMPLR, A1=>nx157);
   ix264 : mux21 port map ( Y=>nx263, A0=>nx376, A1=>nx378, S0=>nx472);
   reg_counter_data_9 : dffr port map ( Q=>counter_out_9_EXMPLR, QB=>nx376, 
      D=>nx263, CLK=>clk, R=>nx462);
   ix379 : oai21 port map ( Y=>nx378, A0=>nx157, A1=>counter_out_9_EXMPLR, 
      B0=>nx372);
   ix254 : mux21_ni port map ( Y=>nx253, A0=>counter_out_8_EXMPLR, A1=>nx94, 
      S0=>nx472);
   reg_counter_data_8 : dffr port map ( Q=>counter_out_8_EXMPLR, QB=>nx381, 
      D=>nx253, CLK=>clk, R=>nx462);
   ix387 : nand02 port map ( Y=>nx386, A0=>counter_out_7_EXMPLR, A1=>nx159);
   ix244 : mux21 port map ( Y=>nx243, A0=>nx390, A1=>nx392, S0=>nx470);
   reg_counter_data_7 : dffr port map ( Q=>counter_out_7_EXMPLR, QB=>nx390, 
      D=>nx243, CLK=>clk, R=>nx464);
   ix393 : oai21 port map ( Y=>nx392, A0=>nx159, A1=>counter_out_7_EXMPLR, 
      B0=>nx386);
   ix234 : mux21_ni port map ( Y=>nx233, A0=>counter_out_6_EXMPLR, A1=>nx70, 
      S0=>nx470);
   reg_counter_data_6 : dffr port map ( Q=>counter_out_6_EXMPLR, QB=>nx395, 
      D=>nx233, CLK=>clk, R=>nx464);
   ix401 : nand02 port map ( Y=>nx400, A0=>counter_out_5_EXMPLR, A1=>nx161);
   ix224 : mux21 port map ( Y=>nx223, A0=>nx404, A1=>nx406, S0=>nx470);
   reg_counter_data_5 : dffr port map ( Q=>counter_out_5_EXMPLR, QB=>nx404, 
      D=>nx223, CLK=>clk, R=>nx464);
   ix407 : oai21 port map ( Y=>nx406, A0=>nx161, A1=>counter_out_5_EXMPLR, 
      B0=>nx400);
   ix214 : mux21_ni port map ( Y=>nx213, A0=>counter_out_4_EXMPLR, A1=>nx46, 
      S0=>nx470);
   reg_counter_data_4 : dffr port map ( Q=>counter_out_4_EXMPLR, QB=>nx409, 
      D=>nx213, CLK=>clk, R=>nx464);
   ix47 : aoi21 port map ( Y=>nx46, A0=>nx414, A1=>nx409, B0=>nx161);
   ix415 : nand04 port map ( Y=>nx414, A0=>counter_out_3_EXMPLR, A1=>
      counter_out_2_EXMPLR, A2=>counter_out_1_EXMPLR, A3=>counter_out_dup0_0
   );
   reg_counter_data_3 : dffr port map ( Q=>counter_out_3_EXMPLR, QB=>OPEN, D
      =>nx203, CLK=>clk, R=>nx466);
   ix204 : mux21_ni port map ( Y=>nx203, A0=>counter_out_3_EXMPLR, A1=>nx34, 
      S0=>nx470);
   ix35 : xnor2 port map ( Y=>nx34, A0=>counter_out_3_EXMPLR, A1=>nx419);
   ix420 : nand03 port map ( Y=>nx419, A0=>counter_out_2_EXMPLR, A1=>
      counter_out_1_EXMPLR, A2=>counter_out_dup0_0);
   reg_counter_data_2 : dffr port map ( Q=>counter_out_2_EXMPLR, QB=>OPEN, D
      =>nx193, CLK=>clk, R=>nx464);
   ix194 : mux21_ni port map ( Y=>nx193, A0=>counter_out_2_EXMPLR, A1=>nx22, 
      S0=>nx470);
   ix23 : xnor2 port map ( Y=>nx22, A0=>counter_out_2_EXMPLR, A1=>nx424);
   ix184 : mux21 port map ( Y=>nx183, A0=>nx428, A1=>nx430, S0=>nx470);
   reg_counter_data_1 : dffr port map ( Q=>counter_out_1_EXMPLR, QB=>nx428, 
      D=>nx183, CLK=>clk, R=>nx464);
   ix431 : oai21 port map ( Y=>nx430, A0=>counter_out_dup0_0, A1=>
      counter_out_1_EXMPLR, B0=>nx424);
   reg_counter_data_0 : dffr port map ( Q=>counter_out_dup0_0, QB=>nx436, D
      =>nx173, CLK=>clk, R=>nx464);
   reg_counter_data_15 : dffr port map ( Q=>counter_out_15_EXMPLR, QB=>nx439, 
      D=>nx323, CLK=>clk, R=>nx466);
   ix247 : and04 port map ( Y=>nx246, A0=>nx445, A1=>nx447, A2=>nx449, A3=>
      nx451);
   ix448 : xnor2 port map ( Y=>nx447, A0=>counter_out_2_EXMPLR, A1=>
      max_val_in(2));
   ix450 : xnor2 port map ( Y=>nx449, A0=>counter_out_3_EXMPLR, A1=>
      max_val_in(3));
   ix193 : and04 port map ( Y=>nx192, A0=>nx439, A1=>nx339, A2=>nx348, A3=>
      nx353);
   ix175 : xor2 port map ( Y=>nx174, A0=>nx149, A1=>counter_out_15_EXMPLR);
   ix173 : nor02ii port map ( Y=>nx149, A0=>nx344, A1=>counter_out_14_EXMPLR
   );
   ix167 : xor2 port map ( Y=>nx166, A0=>nx339, A1=>nx344);
   ix149 : nor02ii port map ( Y=>nx152, A0=>nx358, A1=>counter_out_12_EXMPLR
   );
   ix143 : xor2 port map ( Y=>nx142, A0=>nx353, A1=>nx358);
   ix125 : nor02ii port map ( Y=>nx155, A0=>nx372, A1=>counter_out_10_EXMPLR
   );
   ix119 : xor2 port map ( Y=>nx118, A0=>nx367, A1=>nx372);
   ix101 : nor02ii port map ( Y=>nx157, A0=>nx386, A1=>counter_out_8_EXMPLR
   );
   ix95 : xor2 port map ( Y=>nx94, A0=>nx381, A1=>nx386);
   ix77 : nor02ii port map ( Y=>nx159, A0=>nx400, A1=>counter_out_6_EXMPLR);
   ix71 : xor2 port map ( Y=>nx70, A0=>nx395, A1=>nx400);
   ix53 : nor02ii port map ( Y=>nx161, A0=>nx414, A1=>counter_out_4_EXMPLR);
   ix425 : or02 port map ( Y=>nx424, A0=>nx428, A1=>nx436);
   ix174 : xnor2 port map ( Y=>nx173, A0=>nx436, A1=>nx474);
   ix207 : and04 port map ( Y=>nx206, A0=>nx362, A1=>nx367, A2=>nx376, A3=>
      nx381);
   ix225 : and04 port map ( Y=>nx224, A0=>nx390, A1=>nx395, A2=>nx404, A3=>
      nx458);
   ix217 : xnor2 port map ( Y=>nx458, A0=>max_val_in(0), A1=>
      counter_out_dup0_0);
   ix446 : xor2 port map ( Y=>nx445, A0=>nx428, A1=>max_val_in(1));
   ix452 : xor2 port map ( Y=>nx451, A0=>nx409, A1=>max_val_in(4));
   ix459 : inv01 port map ( Y=>nx460, A=>reset);
   ix461 : inv02 port map ( Y=>nx462, A=>nx460);
   ix463 : inv02 port map ( Y=>nx464, A=>nx460);
   ix465 : inv02 port map ( Y=>nx466, A=>nx460);
   ix467 : inv01 port map ( Y=>nx468, A=>enable);
   ix469 : inv02 port map ( Y=>nx470, A=>nx468);
   ix471 : inv02 port map ( Y=>nx472, A=>nx468);
   ix473 : inv02 port map ( Y=>nx474, A=>nx468);
end behavioural_unfold_2902 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Controller is
   port (
      clk : IN std_logic ;
      reset : IN std_logic ;
      io_ready_in : IN std_logic ;
      io_done_out : OUT std_logic ;
      mem_data_in : IN std_logic_vector (15 DOWNTO 0) ;
      mem_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
      mem_addr_out : OUT std_logic_vector (15 DOWNTO 0) ;
      mem_write_out : OUT std_logic ;
      mem_read_out : OUT std_logic ;
      wind_en : OUT std_logic ;
      wind_rst : OUT std_logic ;
      wind_col_in_4_15 : OUT std_logic ;
      wind_col_in_4_14 : OUT std_logic ;
      wind_col_in_4_13 : OUT std_logic ;
      wind_col_in_4_12 : OUT std_logic ;
      wind_col_in_4_11 : OUT std_logic ;
      wind_col_in_4_10 : OUT std_logic ;
      wind_col_in_4_9 : OUT std_logic ;
      wind_col_in_4_8 : OUT std_logic ;
      wind_col_in_4_7 : OUT std_logic ;
      wind_col_in_4_6 : OUT std_logic ;
      wind_col_in_4_5 : OUT std_logic ;
      wind_col_in_4_4 : OUT std_logic ;
      wind_col_in_4_3 : OUT std_logic ;
      wind_col_in_4_2 : OUT std_logic ;
      wind_col_in_4_1 : OUT std_logic ;
      wind_col_in_4_0 : OUT std_logic ;
      wind_col_in_3_15 : OUT std_logic ;
      wind_col_in_3_14 : OUT std_logic ;
      wind_col_in_3_13 : OUT std_logic ;
      wind_col_in_3_12 : OUT std_logic ;
      wind_col_in_3_11 : OUT std_logic ;
      wind_col_in_3_10 : OUT std_logic ;
      wind_col_in_3_9 : OUT std_logic ;
      wind_col_in_3_8 : OUT std_logic ;
      wind_col_in_3_7 : OUT std_logic ;
      wind_col_in_3_6 : OUT std_logic ;
      wind_col_in_3_5 : OUT std_logic ;
      wind_col_in_3_4 : OUT std_logic ;
      wind_col_in_3_3 : OUT std_logic ;
      wind_col_in_3_2 : OUT std_logic ;
      wind_col_in_3_1 : OUT std_logic ;
      wind_col_in_3_0 : OUT std_logic ;
      wind_col_in_2_15 : OUT std_logic ;
      wind_col_in_2_14 : OUT std_logic ;
      wind_col_in_2_13 : OUT std_logic ;
      wind_col_in_2_12 : OUT std_logic ;
      wind_col_in_2_11 : OUT std_logic ;
      wind_col_in_2_10 : OUT std_logic ;
      wind_col_in_2_9 : OUT std_logic ;
      wind_col_in_2_8 : OUT std_logic ;
      wind_col_in_2_7 : OUT std_logic ;
      wind_col_in_2_6 : OUT std_logic ;
      wind_col_in_2_5 : OUT std_logic ;
      wind_col_in_2_4 : OUT std_logic ;
      wind_col_in_2_3 : OUT std_logic ;
      wind_col_in_2_2 : OUT std_logic ;
      wind_col_in_2_1 : OUT std_logic ;
      wind_col_in_2_0 : OUT std_logic ;
      wind_col_in_1_15 : OUT std_logic ;
      wind_col_in_1_14 : OUT std_logic ;
      wind_col_in_1_13 : OUT std_logic ;
      wind_col_in_1_12 : OUT std_logic ;
      wind_col_in_1_11 : OUT std_logic ;
      wind_col_in_1_10 : OUT std_logic ;
      wind_col_in_1_9 : OUT std_logic ;
      wind_col_in_1_8 : OUT std_logic ;
      wind_col_in_1_7 : OUT std_logic ;
      wind_col_in_1_6 : OUT std_logic ;
      wind_col_in_1_5 : OUT std_logic ;
      wind_col_in_1_4 : OUT std_logic ;
      wind_col_in_1_3 : OUT std_logic ;
      wind_col_in_1_2 : OUT std_logic ;
      wind_col_in_1_1 : OUT std_logic ;
      wind_col_in_1_0 : OUT std_logic ;
      wind_col_in_0_15 : OUT std_logic ;
      wind_col_in_0_14 : OUT std_logic ;
      wind_col_in_0_13 : OUT std_logic ;
      wind_col_in_0_12 : OUT std_logic ;
      wind_col_in_0_11 : OUT std_logic ;
      wind_col_in_0_10 : OUT std_logic ;
      wind_col_in_0_9 : OUT std_logic ;
      wind_col_in_0_8 : OUT std_logic ;
      wind_col_in_0_7 : OUT std_logic ;
      wind_col_in_0_6 : OUT std_logic ;
      wind_col_in_0_5 : OUT std_logic ;
      wind_col_in_0_4 : OUT std_logic ;
      wind_col_in_0_3 : OUT std_logic ;
      wind_col_in_0_2 : OUT std_logic ;
      wind_col_in_0_1 : OUT std_logic ;
      wind_col_in_0_0 : OUT std_logic ;
      filter_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
      filter_ready_out : OUT std_logic ;
      filter_reset : OUT std_logic ;
      comp_unit_ready : OUT std_logic ;
      comp_unit_operation : OUT std_logic ;
      comp_unit_flt_size : OUT std_logic ;
      comp_unit_relu : OUT std_logic ;
      comp_unit_data1_out : OUT std_logic_vector (15 DOWNTO 0) ;
      comp_unit_data2_out : OUT std_logic_vector (15 DOWNTO 0) ;
      comp_unit_buffer_finished : IN std_logic ;
      comp_unit_finished : IN std_logic ;
      comp_unit_data1_in : IN std_logic_vector (15 DOWNTO 0) ;
      comp_unit_data2_in : IN std_logic_vector (15 DOWNTO 0) ;
      argmax_ready : OUT std_logic ;
      argmax_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
      argmax_data_in : IN std_logic_vector (15 DOWNTO 0)) ;
end Controller ;

architecture Mixed of Controller is
   component Cache_5_16_28_5
      port (
         in_word : IN std_logic_vector (15 DOWNTO 0) ;
         cache_in_sel : IN std_logic_vector (4 DOWNTO 0) ;
         cache_out_sel : IN std_logic_vector (4 DOWNTO 0) ;
         decoder_enable : IN std_logic ;
         out_column_0_15 : OUT std_logic ;
         out_column_0_14 : OUT std_logic ;
         out_column_0_13 : OUT std_logic ;
         out_column_0_12 : OUT std_logic ;
         out_column_0_11 : OUT std_logic ;
         out_column_0_10 : OUT std_logic ;
         out_column_0_9 : OUT std_logic ;
         out_column_0_8 : OUT std_logic ;
         out_column_0_7 : OUT std_logic ;
         out_column_0_6 : OUT std_logic ;
         out_column_0_5 : OUT std_logic ;
         out_column_0_4 : OUT std_logic ;
         out_column_0_3 : OUT std_logic ;
         out_column_0_2 : OUT std_logic ;
         out_column_0_1 : OUT std_logic ;
         out_column_0_0 : OUT std_logic ;
         out_column_1_15 : OUT std_logic ;
         out_column_1_14 : OUT std_logic ;
         out_column_1_13 : OUT std_logic ;
         out_column_1_12 : OUT std_logic ;
         out_column_1_11 : OUT std_logic ;
         out_column_1_10 : OUT std_logic ;
         out_column_1_9 : OUT std_logic ;
         out_column_1_8 : OUT std_logic ;
         out_column_1_7 : OUT std_logic ;
         out_column_1_6 : OUT std_logic ;
         out_column_1_5 : OUT std_logic ;
         out_column_1_4 : OUT std_logic ;
         out_column_1_3 : OUT std_logic ;
         out_column_1_2 : OUT std_logic ;
         out_column_1_1 : OUT std_logic ;
         out_column_1_0 : OUT std_logic ;
         out_column_2_15 : OUT std_logic ;
         out_column_2_14 : OUT std_logic ;
         out_column_2_13 : OUT std_logic ;
         out_column_2_12 : OUT std_logic ;
         out_column_2_11 : OUT std_logic ;
         out_column_2_10 : OUT std_logic ;
         out_column_2_9 : OUT std_logic ;
         out_column_2_8 : OUT std_logic ;
         out_column_2_7 : OUT std_logic ;
         out_column_2_6 : OUT std_logic ;
         out_column_2_5 : OUT std_logic ;
         out_column_2_4 : OUT std_logic ;
         out_column_2_3 : OUT std_logic ;
         out_column_2_2 : OUT std_logic ;
         out_column_2_1 : OUT std_logic ;
         out_column_2_0 : OUT std_logic ;
         out_column_3_15 : OUT std_logic ;
         out_column_3_14 : OUT std_logic ;
         out_column_3_13 : OUT std_logic ;
         out_column_3_12 : OUT std_logic ;
         out_column_3_11 : OUT std_logic ;
         out_column_3_10 : OUT std_logic ;
         out_column_3_9 : OUT std_logic ;
         out_column_3_8 : OUT std_logic ;
         out_column_3_7 : OUT std_logic ;
         out_column_3_6 : OUT std_logic ;
         out_column_3_5 : OUT std_logic ;
         out_column_3_4 : OUT std_logic ;
         out_column_3_3 : OUT std_logic ;
         out_column_3_2 : OUT std_logic ;
         out_column_3_1 : OUT std_logic ;
         out_column_3_0 : OUT std_logic ;
         out_column_4_15 : OUT std_logic ;
         out_column_4_14 : OUT std_logic ;
         out_column_4_13 : OUT std_logic ;
         out_column_4_12 : OUT std_logic ;
         out_column_4_11 : OUT std_logic ;
         out_column_4_10 : OUT std_logic ;
         out_column_4_9 : OUT std_logic ;
         out_column_4_8 : OUT std_logic ;
         out_column_4_7 : OUT std_logic ;
         out_column_4_6 : OUT std_logic ;
         out_column_4_5 : OUT std_logic ;
         out_column_4_4 : OUT std_logic ;
         out_column_4_3 : OUT std_logic ;
         out_column_4_2 : OUT std_logic ;
         out_column_4_1 : OUT std_logic ;
         out_column_4_0 : OUT std_logic ;
         clk : IN std_logic ;
         reset : IN std_logic) ;
   end component ;
   component AdvancedCounter_16
      port (
         clk : IN std_logic ;
         reset : IN std_logic ;
         enable : IN std_logic ;
         mode_in : IN std_logic_vector (1 DOWNTO 0) ;
         max_val_in : IN std_logic_vector (15 DOWNTO 0) ;
         max_reached_out : OUT std_logic ;
         counter_out : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   signal current_state_12, wind_width_count_4, wind_width_count_3, 
      wind_width_count_2, wind_width_count_1, wind_width_count_0, 
      cache_height_count_en, cache_height_ended, max_height_4, max_height_3, 
      max_height_2, max_height_0, cache_width_count_4, cache_width_count_3, 
      cache_width_count_2, cache_width_count_1, cache_width_count_0, 
      cache_data_in_15, cache_data_in_14, cache_data_in_13, cache_data_in_12, 
      cache_data_in_11, cache_data_in_10, cache_data_in_9, cache_data_in_8, 
      cache_data_in_7, cache_data_in_6, cache_data_in_5, cache_data_in_4, 
      cache_data_in_3, cache_data_in_2, cache_data_in_1, cache_data_in_0, 
      cache_data_out_4_15, cache_data_out_4_14, cache_data_out_4_13, 
      cache_data_out_4_12, cache_data_out_4_11, cache_data_out_4_10, 
      cache_data_out_4_9, cache_data_out_4_8, cache_data_out_4_7, 
      cache_data_out_4_6, cache_data_out_4_5, cache_data_out_4_4, 
      cache_data_out_4_3, cache_data_out_4_2, cache_data_out_4_1, 
      cache_data_out_4_0, cache_data_out_3_15, cache_data_out_3_14, 
      cache_data_out_3_13, cache_data_out_3_12, cache_data_out_3_11, 
      cache_data_out_3_10, cache_data_out_3_9, cache_data_out_3_8, 
      cache_data_out_3_7, cache_data_out_3_6, cache_data_out_3_5, 
      cache_data_out_3_4, cache_data_out_3_3, cache_data_out_3_2, 
      cache_data_out_3_1, cache_data_out_3_0, cache_data_out_2_15, 
      cache_data_out_2_14, cache_data_out_2_13, cache_data_out_2_12, 
      cache_data_out_2_11, cache_data_out_2_10, cache_data_out_2_9, 
      cache_data_out_2_8, cache_data_out_2_7, cache_data_out_2_6, 
      cache_data_out_2_5, cache_data_out_2_4, cache_data_out_2_3, 
      cache_data_out_2_2, cache_data_out_2_1, cache_data_out_2_0, 
      cache_data_out_1_15, cache_data_out_1_14, cache_data_out_1_13, 
      cache_data_out_1_12, cache_data_out_1_11, cache_data_out_1_10, 
      cache_data_out_1_9, cache_data_out_1_8, cache_data_out_1_7, 
      cache_data_out_1_6, cache_data_out_1_5, cache_data_out_1_4, 
      cache_data_out_1_3, cache_data_out_1_2, cache_data_out_1_1, 
      cache_data_out_1_0, cache_data_out_0_15, cache_data_out_0_14, 
      cache_data_out_0_13, cache_data_out_0_12, cache_data_out_0_11, 
      cache_data_out_0_10, cache_data_out_0_9, cache_data_out_0_8, 
      cache_data_out_0_7, cache_data_out_0_6, cache_data_out_0_5, 
      cache_data_out_0_4, cache_data_out_0_3, cache_data_out_0_2, 
      cache_data_out_0_1, cache_data_out_0_0, cache_load, cache_rst_actual, 
      max_height_1, comp_unit_operation_EXMPLR, argmax_ready_EXMPLR, 
      filter_ready_out_EXMPLR, wind_rst_EXMPLR, current_state_20, 
      ftc_cntrl_reg_out_8, current_state_15, current_state_14, 
      current_state_23, ftc_cntrl_reg_out_12, ftc_cntrl_reg_out_10, 
      current_state_9, current_state_8, current_state_6, current_state_5, 
      current_state_4, current_state_2, current_state_24, 
      num_channels_counter_out_2, nx12230, nx4, nx12231, 
      write_offset_data_out_0, nx8, new_size_squared_out_0, 
      write_offset_data_out_1, nx26, new_size_squared_out_1, 
      write_offset_data_out_2, new_size_squared_out_2, 
      write_offset_data_out_3, nx78, new_size_squared_out_3, nx96, 
      write_offset_data_out_4, nx98, nx104, new_size_squared_out_4, 
      write_offset_data_out_5, new_size_squared_out_5, 
      write_offset_data_out_6, nx144, nx150, new_size_squared_out_6, 
      write_offset_data_out_7, new_size_squared_out_7, nx190, 
      write_offset_data_out_8, nx194, nx200, new_size_squared_out_8, 
      write_offset_data_out_9, new_size_squared_out_9, 
      write_offset_data_out_10, nx240, nx246, new_size_squared_out_10, 
      write_offset_data_out_11, new_size_squared_out_11, nx286, 
      write_offset_data_out_12, nx288, nx294, new_size_squared_out_12, 
      write_offset_data_out_13, new_size_squared_out_13, 
      write_offset_data_out_14, nx334, nx340, new_size_squared_out_14, 
      new_size_squared_out_15, nx374, nx386, num_channels_counter_out_1, 
      num_channels_counter_out_0, nflt_layer_temp_0, current_state_1, 
      current_state_0, nx426, nflt_layer_temp_1, nx454, nx466, 
      nflt_layer_temp_2, nx492, nflt_layer_cntr_counter_out_3, nx496, 
      nflt_layer_cntr_counter_out_2, nflt_layer_cntr_counter_out_1, 
      nflt_layer_cntr_counter_out_0, nx506, nx524, nx544, nx560, 
      nlayers_counter_out_0, nlayers_counter_out_2, nlayers_counter_out_1, 
      nx600, layer_type_out_1, nx646, nx650, nx662, nx670, nx680, 
      cntr1_inst_counter_out_1, cntr1_inst_counter_out_0, nx684, nx702, 
      cntr1_inst_counter_out_3, cntr1_inst_counter_out_2, nx708, nx722, 
      nx728, cntr1_inst_counter_out_5, cntr1_inst_counter_out_4, nx12238, 
      nx740, flt_size_out_0, flt_size_out_2, flt_size_out_1, nx786, nx794, 
      nx808, nx12239, nx814, ftc_cntrl_reg_out_13, nx830, nx856, nx862, 
      cache_width_cntr_counter_out_14, nx12241, 
      cache_width_cntr_counter_out_13, cache_width_cntr_counter_out_12, 
      nx12243, cache_width_cntr_counter_out_11, 
      cache_width_cntr_counter_out_10, nx12245, 
      cache_width_cntr_counter_out_9, cache_width_cntr_counter_out_8, 
      nx12247, cache_width_cntr_counter_out_7, 
      cache_width_cntr_counter_out_6, nx12249, nx866, nx874, nx880, nx888, 
      nx896, nx904, cache_width_cntr_counter_out_5, nx910, nx930, nx954, 
      nx978, nx1002, nx1026, nx1052, nx1066, img_width_out_0, 
      new_width_out_0, nx1098, img_width_out_1, new_width_out_1, nx1112, 
      nx1120, img_width_out_2, new_width_out_2, nx1144, img_width_out_3, 
      new_width_out_3, nx1172, img_width_out_4, new_width_out_4, nx1188, 
      nx1196, nx1200, ftc_cntrl_reg_out_14, nx12251, nx1226, nx1240, nx1246, 
      nx1256, nx1266, ftc_cntrl_reg_out_9, ftc_cntrl_reg_out_11, nx12253, 
      window_width_cntr_counter_out_14, nx12254, 
      window_width_cntr_counter_out_13, window_width_cntr_counter_out_12, 
      nx12256, window_width_cntr_counter_out_11, 
      window_width_cntr_counter_out_10, nx12258, 
      window_width_cntr_counter_out_9, window_width_cntr_counter_out_8, 
      nx12260, window_width_cntr_counter_out_7, 
      window_width_cntr_counter_out_6, nx12262, 
      window_width_cntr_counter_out_5, nx1278, nx1284, nx1292, nx1300, 
      nx1308, nx1328, nx1352, nx1376, nx1400, nx1424, nx1450, nx1464, 
      nx12265, nx1478, nx1486, nx1488, nx1494, nx1504, nx1508, nx1518, 
      nx1534, nx1542, nx1556, nx12266, nx1576, nx1584, nx12267, 
      current_state_18, current_state_17, nx1622, nx1628, nx1644, nx1654, 
      nx1692, current_state_25, class_cntr_counter_out_3, 
      class_cntr_counter_out_2, class_cntr_counter_out_1, 
      class_cntr_counter_out_0, nx1720, nx1728, nx1742, nx1754, nx1762, 
      flt_bias_out_0, nx1960, nx1966, flt_bias_out_1, nx1994, flt_bias_out_2, 
      nx2020, flt_bias_out_3, nx2046, flt_bias_out_4, nx2072, flt_bias_out_5, 
      nx2098, flt_bias_out_6, nx2124, flt_bias_out_7, nx2150, flt_bias_out_8, 
      nx2176, flt_bias_out_9, nx2202, flt_bias_out_10, nx2228, 
      flt_bias_out_11, nx2254, flt_bias_out_12, nx2280, flt_bias_out_13, 
      nx2306, flt_bias_out_14, nx2332, flt_bias_out_15, nx2358, nx2372, 
      ftc_cntrl_reg_out_15, nx2392, nx2406, nx2478, layer_mem_size_out_0, 
      nx2494, nx2502, nx2520, nx2526, nx2532, bias_offset_data_out_0, 
      addr1_data_0, nx2568, nx2572, img_addr_offset_0, nx2610, 
      img_addr_offset_1, write_base_data_out_1, layer_mem_size_out_1, nx2658, 
      bias_offset_data_out_1, nx2670, addr1_data_1, write_base_data_out_2, 
      layer_mem_size_out_2, nx2758, img_addr_offset_2, nx2768, nx2774, 
      nx2780, nx2794, addr1_data_2, nx2822, bias_offset_data_out_3, 
      write_base_data_out_3, layer_mem_size_out_3, nx2890, img_addr_offset_3, 
      nx2900, nx2906, nx2908, nx2926, addr1_data_3, nx2954, 
      write_base_data_out_4, layer_mem_size_out_4, nx3016, img_addr_offset_4, 
      nx3038, nx3044, nx3060, bias_offset_data_out_4, addr1_data_4, nx3084, 
      nx3090, write_base_data_out_5, layer_mem_size_out_5, nx3152, 
      img_addr_offset_5, nx3170, nx3188, bias_offset_data_out_5, 
      addr1_data_5, write_base_data_out_6, layer_mem_size_out_6, nx3280, 
      nx3286, img_addr_offset_6, nx3294, nx3300, nx3316, 
      bias_offset_data_out_6, addr1_data_6, nx3340, nx3346, 
      write_base_data_out_7, layer_mem_size_out_7, nx3408, img_addr_offset_7, 
      nx3426, nx3444, bias_offset_data_out_7, addr1_data_7, nx3492, 
      write_base_data_out_8, layer_mem_size_out_8, nx3534, nx3536, 
      img_addr_offset_8, nx3540, nx3546, nx3554, nx3564, nx3572, 
      bias_offset_data_out_8, addr1_data_8, nx3596, nx3602, 
      write_base_data_out_9, layer_mem_size_out_9, nx3664, img_addr_offset_9, 
      nx3682, nx3692, nx3700, bias_offset_data_out_9, addr1_data_9, nx3748, 
      write_base_data_out_10, layer_mem_size_out_10, nx3792, 
      img_addr_offset_10, nx3796, nx3802, nx3810, nx3820, nx3828, 
      bias_offset_data_out_10, addr1_data_10, nx3852, nx3858, 
      write_base_data_out_11, layer_mem_size_out_11, nx3920, 
      img_addr_offset_11, nx3946, nx3956, bias_offset_data_out_11, 
      addr1_data_11, write_base_data_out_12, layer_mem_size_out_12, nx4048, 
      nx4054, img_addr_offset_12, nx4062, nx4068, nx4084, 
      bias_offset_data_out_12, addr1_data_12, nx4108, nx4114, 
      write_base_data_out_13, layer_mem_size_out_13, img_addr_offset_13, 
      nx4194, bias_offset_data_out_13, addr1_data_13, write_base_data_out_14, 
      layer_mem_size_out_14, nx4304, img_addr_offset_14, nx4308, nx4314, 
      nx4320, nx4330, bias_offset_data_out_14, addr1_data_14, nx4364, nx4370, 
      write_base_data_out_15, nx4406, layer_mem_size_out_15, nx4428, 
      addr1_data_15, nx12277, nx12287, nx12297, nx12307, nx12317, nx12327, 
      nx12337, nx12347, nx12357, nx12367, nx12377, nx12387, nx12397, nx12407, 
      nx12417, nx12427, nx12437, nx12447, nx12457, nx12467, nx12477, nx12487, 
      nx12497, nx12507, nx12517, nx12527, nx12537, nx12547, nx12557, nx12567, 
      nx12577, nx12587, nx12597, nx12607, nx12617, nx12627, nx12637, nx12647, 
      nx12657, nx12667, nx12677, nx12687, nx12697, nx12707, nx12717, nx12727, 
      nx12737, nx12747, nx12757, nx12767, nx12777, nx12787, nx12797, nx12807, 
      nx12817, nx12827, nx12837, nx12847, nx12857, nx12867, nx12877, nx12887, 
      nx12897, nx12907, nx12917, nx12927, nx12937, nx12947, nx12957, nx12967, 
      nx12977, nx12987, nx12997, nx13007, nx13017, nx13027, nx13037, nx13047, 
      nx13057, nx13067, nx13077, nx13087, nx13097, nx13107, nx13117, nx13127, 
      nx13137, nx13147, nx13157, nx13167, nx13177, nx13187, nx13197, nx13207, 
      nx13217, nx13227, nx13237, nx13247, nx13257, nx13267, nx13277, nx13287, 
      nx13297, nx13307, nx13317, nx13327, nx13337, nx13347, nx13357, nx13367, 
      nx13377, nx13387, nx13397, nx13407, nx13417, nx13427, nx13437, nx13447, 
      nx13457, nx13467, nx13477, nx13487, nx13497, nx13507, nx13517, nx13527, 
      nx13537, nx13547, nx13557, nx13567, nx13577, nx13587, nx13597, nx13607, 
      nx13617, nx13627, nx13637, nx13647, nx13657, nx13667, nx13677, nx13687, 
      nx13697, nx13707, nx13717, nx13727, nx13737, nx13747, nx13757, nx13767, 
      nx13777, nx13787, nx13797, nx13807, nx13817, nx13827, nx13837, nx13847, 
      nx13857, nx13867, nx13877, nx13887, nx13897, nx13907, nx13917, nx13927, 
      nx13937, nx13947, nx13957, nx13967, nx13977, nx13987, nx13997, nx14007, 
      nx14017, nx14027, nx14037, nx14047, nx14057, nx14067, nx14077, nx14087, 
      nx14097, nx14107, nx14117, nx14127, nx14137, nx14147, nx14157, nx14167, 
      nx14177, nx14187, nx14197, nx14207, nx14217, nx14227, nx14237, nx14247, 
      nx14257, nx14277, nx14287, nx14297, nx14307, nx14317, nx14327, nx14337, 
      nx14347, nx14357, nx14367, nx14377, nx14387, nx14397, nx14407, nx14427, 
      nx14437, nx14447, nx14457, nx14467, nx14487, nx14497, nx14508, nx14512, 
      nx14515, nx14520, nx14525, nx14530, nx14534, nx14540, nx14542, nx14544, 
      nx14546, nx14549, nx14553, nx14555, nx14561, nx14564, nx14567, nx14571, 
      nx14573, nx14577, nx14585, nx14597, nx14604, nx14606, nx14615, nx14620, 
      nx14627, nx14632, nx14635, nx14640, nx14644, nx14647, nx14651, nx14653, 
      nx14656, nx14660, nx14663, nx14669, nx14673, nx14676, nx14682, nx14686, 
      nx14689, nx14695, nx14699, nx14702, nx14708, nx14712, nx14715, nx14717, 
      nx14722, nx14723, nx14726, nx14732, nx14736, nx14738, nx14741, nx14747, 
      nx14751, nx14756, nx14759, nx14762, nx14765, nx14769, nx14771, nx14774, 
      nx14776, nx14778, nx14780, nx14782, nx14787, nx14791, nx14792, nx14797, 
      nx14801, nx14803, nx14808, nx14812, nx14813, nx14818, nx14822, nx14824, 
      nx14829, nx14833, nx14834, nx14839, nx14843, nx14845, nx14850, nx14854, 
      nx14855, nx14860, nx14865, nx14867, nx14871, nx14873, nx14875, nx14878, 
      nx14882, nx14884, nx14887, nx14892, nx14895, nx14897, nx14899, nx14902, 
      nx14905, nx14910, nx14914, nx14916, nx14919, nx14924, nx14928, nx14930, 
      nx14933, nx14938, nx14942, nx14944, nx14947, nx14952, nx14956, nx14958, 
      nx14961, nx14966, nx14971, nx14983, nx14985, nx14988, nx14990, nx15000, 
      nx15006, nx15012, nx15014, nx15027, nx15029, nx15032, nx15040, nx15043, 
      nx15052, nx15055, nx15064, nx15072, nx15075, nx15077, nx15080, nx15082, 
      nx15087, nx15089, nx15092, nx15094, nx15097, nx15102, nx15106, nx15108, 
      nx15111, nx15116, nx15120, nx15122, nx15125, nx15130, nx15134, nx15136, 
      nx15139, nx15144, nx15148, nx15150, nx15153, nx15158, nx15163, nx15180, 
      nx15186, nx15192, nx15194, nx15201, nx15204, nx15207, nx15210, nx15213, 
      nx15216, nx15219, nx15223, nx15226, nx15231, nx15240, nx15242, nx15247, 
      nx15249, nx15251, nx15257, nx15259, nx15265, nx15267, nx15269, nx15272, 
      nx15274, nx15293, nx15297, nx15304, nx15309, nx15311, nx15313, nx15320, 
      nx15322, nx15329, nx15332, nx15336, nx15339, nx15344, nx15347, nx15350, 
      nx15353, nx15358, nx15360, nx15362, nx15364, nx15372, nx15374, nx15399, 
      nx15480, nx15483, nx15489, nx15531, nx15538, nx15541, nx15547, nx15550, 
      nx15553, nx15556, nx15559, nx15562, nx15565, nx15568, nx15571, nx15574, 
      nx15577, nx15580, nx15583, nx15586, nx15589, nx15592, nx15595, nx15598, 
      nx15601, nx15604, nx15607, nx15610, nx15613, nx15616, nx15619, nx15622, 
      nx15625, nx15628, nx15631, nx15634, nx15637, nx15656, nx15739, nx15742, 
      nx15747, nx15750, nx15753, nx15755, nx15758, nx15762, nx15777, nx15781, 
      nx15785, nx15791, nx15793, nx15795, nx15803, nx15805, nx15811, nx15815, 
      nx15818, nx15821, nx15823, nx15829, nx15832, nx15834, nx15838, nx15840, 
      nx15849, nx15851, nx15855, nx15857, nx15860, nx15864, nx15870, nx15875, 
      nx15878, nx15884, nx15891, nx15900, nx15901, nx15905, nx15908, nx15913, 
      nx15924, nx15927, nx15932, nx15934, nx15943, nx15948, nx15951, nx15956, 
      nx15958, nx15961, nx15963, nx15968, nx15970, nx15974, nx15987, nx15991, 
      nx15995, nx16005, nx16010, nx16017, nx16026, nx16027, nx16029, nx16033, 
      nx16036, nx16040, nx16045, nx16047, nx16051, nx16054, nx16057, nx16061, 
      nx16065, nx16068, nx16070, nx16073, nx16078, nx16080, nx16083, nx16086, 
      nx16088, nx16097, nx16102, nx16106, nx16108, nx16110, nx16114, nx16124, 
      nx16127, nx16134, nx16143, nx16146, nx16151, nx16155, nx16158, nx16161, 
      nx16166, nx16169, nx16172, nx16175, nx16179, nx16183, nx16186, nx16188, 
      nx16191, nx16196, nx16198, nx16201, nx16205, nx16207, nx16213, nx16216, 
      nx16221, nx16225, nx16227, nx16229, nx16233, nx16243, nx16246, nx16253, 
      nx16262, nx16265, nx16270, nx16274, nx16277, nx16280, nx16285, nx16290, 
      nx16293, nx16297, nx16301, nx16304, nx16306, nx16309, nx16314, nx16316, 
      nx16319, nx16323, nx16325, nx16328, nx16331, nx16334, nx16339, nx16343, 
      nx16345, nx16347, nx16349, nx16353, nx16363, nx16366, nx16373, nx16382, 
      nx16385, nx16390, nx16394, nx16397, nx16400, nx16405, nx16410, nx16413, 
      nx16417, nx16434, nx16436, nx16439, nx16443, nx16445, nx16454, nx16459, 
      nx16463, nx16465, nx16467, nx16469, nx16472, nx16482, nx16485, nx16492, 
      nx16501, nx16504, nx16509, nx16513, nx16516, nx16519, nx16524, nx16528, 
      nx16538, nx16547, nx16550, nx16555, nx16557, nx16560, nx16564, nx16580, 
      nx16584, nx16586, nx16588, nx16592, nx16602, nx16621, nx16622, nx16624, 
      nx16629, nx16635, nx16636, nx16642, nx16647, nx16650, nx16661, nx16663, 
      nx16677, nx16686, nx16689, nx16693, nx16696, nx16699, nx16702, nx16705, 
      nx16708, nx16711, nx16714, nx16717, nx16720, nx16723, nx16726, nx16729, 
      nx16732, nx16735, nx16738, nx16741, nx16744, nx16751, nx16753, nx16755, 
      nx16757, nx16759, nx16761, nx16763, nx16765, nx16767, nx16769, nx16771, 
      nx16773, nx16775, nx16777, nx16779, nx16781, nx16783, nx16795, nx16797, 
      nx16803, nx16805, nx16809, nx16811, nx16815, nx16817, nx16819, nx16821, 
      nx16835, nx16837, nx16839, nx16841, nx16843, nx16847, nx16849, nx16851, 
      nx16857, nx16865, nx16867, nx16869, nx16871, nx16879, nx16881, nx16883, 
      nx16885, nx16891, nx16893, nx16895, nx16897, nx16905, nx16913, nx16915, 
      nx16917, nx16923, nx16925, nx16927, nx16935, nx16937, nx16939, nx16941, 
      nx16945, nx16947, nx16949, nx16951, nx16953, nx16955, nx16957, nx16959, 
      nx16961, nx16963, nx16967, nx16969, nx16971, nx16977, nx16979, nx16981, 
      nx16983, nx16985, nx17009, nx17011, nx17013, nx17015, nx17017, nx17019, 
      nx17021, nx17023, nx17027, nx17029, nx17035, nx17037, nx17039, nx17045, 
      nx17047, nx17049, nx17051, nx17053, nx17055, nx17057, nx17059, nx17061, 
      nx17063, nx17065, nx17067, nx17069, nx17071, nx17073, nx17075, nx17077, 
      nx17079, nx17081, nx17083, nx17085, nx17087, nx17089, nx17091, nx17093, 
      nx17095, nx17097, nx17099, nx17101, nx17103, nx17105, nx17107, nx17109, 
      nx17111, nx17113, nx17115, nx17117, nx17119, nx17121, nx17123, nx17125, 
      nx17127, nx17129, nx17131, nx17133, nx17135, nx17137, nx17139, nx17141, 
      nx17143, nx17145, nx17147, nx17149, nx17151, nx17153, nx17155, nx17159, 
      nx17161, nx17163, nx17165, nx17167, nx17171, nx17175, nx17179, nx17183, 
      nx17187, nx17191, nx17193, nx17195, nx17197, nx17199, nx17201, nx17203, 
      nx17205, nx17207, nx17209, nx17211, nx17213, nx17217, nx17219, nx17221, 
      nx17223, nx17225, nx17227, nx17229, nx17231, nx17233, nx17235, nx17237, 
      nx17239, nx17245, nx17247, nx17390, nx15886, nx15889, nx17391, nx17392, 
      nx17393, nx17394, nx17395, nx17396, nx17397, nx17398, nx17399, nx17400, 
      nx17401, nx4420, nx17402, nx17403, nx17404, nx16494, nx16497, nx17405, 
      nx16378, nx17406, nx16614, nx17407, nx17408, nx17409, nx17410, nx17411, 
      nx17412, nx17413, nx17414, nx17415, nx17416, nx17417, nx17418, nx17419, 
      nx17420, nx17421, nx17422, nx14417, nx16610, nx16490, nx17423, nx17424, 
      nx17425, nx17426, nx17427, nx17428, nx17429, nx17430, nx17431, nx16371, 
      nx17432, nx17433, nx17434, nx17435, nx17436, nx17437, nx17438, nx15893, 
      nx17439, nx15896, nx15842, nx17440, nx17441, nx17442, nx17443, nx17444, 
      nx17445, nx17446, nx17447, nx17448, nx17449, nx17450, nx17451, nx17452, 
      nx17453, nx17454, nx17455, nx17456, nx17457, nx17458, nx17459, nx17460, 
      nx17461, nx17462, nx17463, nx17464, nx2472, nx17465, nx16597, nx4260, 
      nx17466, nx17467, nx17468, nx17469, nx17470, nx17471, nx17472, nx17473, 
      nx15981, nx17474, nx2790, nx15800, nx15867, nx16919, nx17475, nx17476, 
      nx16487, nx17477, nx17478, nx17479, nx17480, nx17481, nx17482, nx17483, 
      nx17484, nx16542, nx16545, nx17485, nx17486, nx17487, nx17488, nx17489, 
      nx17490, nx17491, nx17492, nx17493, nx17494, nx17495, nx17496, nx16594, 
      nx17497, nx16474, nx17189, nx16477, nx17498, nx17499, nx17500, nx17501, 
      nx17502, nx17503, nx17504, nx17505, nx17506, nx17507, nx17508, nx17509, 
      nx17510, nx15946, nx15836, nx17511, nx17512, nx15917, nx17513, nx17514, 
      nx17515, nx17169, nx17516, nx17517, nx17518, nx17519, nx17520, nx15997, 
      nx17521, nx16000, nx17522, nx15920, nx17523, nx17524, nx17525, nx17526, 
      nx17527, nx17528, nx16019, nx17529, nx17530, nx17531, nx17532, nx17533, 
      nx17534, nx17535, nx17536, nx17537, nx17538, nx17539, nx17540, nx17541, 
      nx17542, nx17543, nx17544, nx17545, nx4004, nx17546, nx16448, nx16451, 
      nx17547, nx17548, nx17549, nx17550, nx17551, nx17552, nx17553, nx17554, 
      nx17555, nx17556, nx17557, nx17558, nx4154, nx17559, nx17560, nx17561, 
      nx16375, nx17562, nx17563, nx16255, nx16258, nx17564, nx17565, nx17566, 
      nx17567, nx17568, nx17569, nx17570, nx17571, nx17185, nx17572, nx17573, 
      nx17574, nx17575, nx17576, nx17577, nx17578, nx17579, nx17580, nx17581, 
      nx3966, nx17582, nx17583, nx17584, nx17585, nx17586, nx16355, nx16358, 
      nx17587, nx16235, nx16238, nx17588, nx17589, nx17590, nx17591, nx4336, 
      nx17592, nx17593, nx17594, nx3926, nx16456, nx17595, nx17596, nx17597, 
      nx17598, nx16605, nx17599, nx17600, nx17601, nx17602, nx2854, nx17603, 
      nx17604, nx17605, nx17606, nx16129, nx17607, nx3116, nx17608, nx16012, 
      nx16015, nx17025, nx17609, nx17610, nx4222, nx17611, nx17612, nx17613, 
      nx17614, nx17615, nx17616, nx17617, nx16572, nx17618, nx17619, nx17620, 
      nx17621, nx17622, nx17623, nx17624, nx17625, nx17626, nx17627, nx17628, 
      nx17629, nx17630, nx17631, nx17632, nx16534, nx17633, nx4204, 
      NOT_nx16569, nx16577, nx17634, nx17635, nx17636, nx17637, nx17638, 
      nx17639, nx17640, nx3236, nx17641, nx17642, nx17643, nx17644, nx16091, 
      nx17645, nx17646, nx16094, nx2972, nx15984, nx17647, nx17648, nx17649, 
      nx17650, nx17651, nx17652, nx17653, nx17654, nx17655, nx17656, nx17657, 
      nx17658, nx17659, nx3180, nx17660, nx17661, nx17662, nx3026, nx17663, 
      nx16099, nx17664, nx17665, nx17666, nx17667, nx15936, nx15939, nx2808, 
      nx17668, nx17669, nx15825, nx17670, nx17671, nx17672, nx17673, nx17674, 
      nx17675, nx17676, nx17677, nx17678, nx17679, nx16210, nx17680, nx17681, 
      nx17682, nx17683, nx17684, nx17685, nx17686, nx17687, nx17688, nx17689, 
      nx17690, nx17691, nx3710, nx17692, nx17693, nx17694, nx16116, nx17695, 
      nx16119, nx17696, nx17697, nx17698, nx17699, nx17700, nx17701, nx17702, 
      nx17703, nx17704, nx17705, nx17706, nx17707, nx17708, nx17709, nx17710, 
      nx17711, nx17712, nx17713, nx17714, nx17715, nx3198, nx17716, nx3454, 
      nx17717, nx17718, nx17719, nx16336, nx3436, nx16218, nx17720, nx17721, 
      nx17722, nx17723, nx17724, nx17725, nx17726, nx17727, nx17728, nx17729, 
      nx17181, nx17730, nx17731, nx3628, nx17732, nx17733, nx17734, nx17735, 
      NOT_nx16607, nx17736, nx17737, nx17738, nx16368, nx17739, nx17740, 
      nx16248, nx16251, nx3372, nx16132, nx17741, nx17173, nx17742, nx17743, 
      nx17744, nx17745, nx17746, nx17747, nx17177, nx17748, nx17749, nx17750, 
      nx3642, nx17751, nx17752, nx17753, nx17754, nx17755, nx17756, nx17757, 
      nx16136, nx16139, nx3130, nx17758, nx16022, nx17759, nx17760, nx17761, 
      nx17762, nx17763, NOT_nx3386, nx17764, nx17765, nx17766, nx17767, 
      nx17768, nx17769, nx17770, nx17771, nx17772, nx17215, nx17773, nx17774, 
      nx17775, nx17776, nx17777, nx17778, nx14477, nx17779, nx17780, nx17781, 
      nx17782, nx17783, nx17784, nx17785, nx17786, nx17787, nx17788, nx17789, 
      nx17790, nx16943, nx17791, nx17792, nx17793, nx17794, nx17795, nx17796, 
      nx17797, nx14267, nx16424, nx16429, nx17798, nx17799, nx17800, nx17801, 
      nx17802, nx2868, nx17803, nx17804, nx17805, nx17806, nx17807, nx17808, 
      nx17809, nx17810, nx17811, nx17812, nx17813, nx17814, nx17815, nx17816, 
      nx17817, nx17818, nx17819, nx17820, nx17821, nx17822, nx17823, nx17824, 
      nx17825, nx17826, nx17827, nx17828, nx17829, nx17830, nx17831, nx17832, 
      nx17833, nx17834, nx17835, nx17836, nx17837, nx17838, nx17839, nx17840, 
      nx18293, nx18295, nx18297, nx18299, nx18301, nx18303, nx18305, nx18307
   : std_logic ;
   
   signal DANGLING : std_logic_vector (15 downto 0 );

begin
   io_done_out <= wind_rst_EXMPLR ;
   wind_rst <= wind_rst_EXMPLR ;
   filter_ready_out <= filter_ready_out_EXMPLR ;
   filter_reset <= reset ;
   comp_unit_operation <= comp_unit_operation_EXMPLR ;
   argmax_ready <= argmax_ready_EXMPLR ;
   img_cache : Cache_5_16_28_5 port map ( in_word(15)=>cache_data_in_15, 
      in_word(14)=>cache_data_in_14, in_word(13)=>cache_data_in_13, 
      in_word(12)=>cache_data_in_12, in_word(11)=>cache_data_in_11, 
      in_word(10)=>cache_data_in_10, in_word(9)=>cache_data_in_9, in_word(8)
      =>cache_data_in_8, in_word(7)=>cache_data_in_7, in_word(6)=>
      cache_data_in_6, in_word(5)=>cache_data_in_5, in_word(4)=>
      cache_data_in_4, in_word(3)=>cache_data_in_3, in_word(2)=>
      cache_data_in_2, in_word(1)=>cache_data_in_1, in_word(0)=>
      cache_data_in_0, cache_in_sel(4)=>nx16759, cache_in_sel(3)=>
      cache_width_count_3, cache_in_sel(2)=>nx16763, cache_in_sel(1)=>
      cache_width_count_1, cache_in_sel(0)=>cache_width_count_0, 
      cache_out_sel(4)=>wind_width_count_4, cache_out_sel(3)=>
      wind_width_count_3, cache_out_sel(2)=>wind_width_count_2, 
      cache_out_sel(1)=>wind_width_count_1, cache_out_sel(0)=>nx16755, 
      decoder_enable=>cache_load, out_column_0_15=>cache_data_out_4_15, 
      out_column_0_14=>cache_data_out_4_14, out_column_0_13=>
      cache_data_out_4_13, out_column_0_12=>cache_data_out_4_12, 
      out_column_0_11=>cache_data_out_4_11, out_column_0_10=>
      cache_data_out_4_10, out_column_0_9=>cache_data_out_4_9, 
      out_column_0_8=>cache_data_out_4_8, out_column_0_7=>cache_data_out_4_7, 
      out_column_0_6=>cache_data_out_4_6, out_column_0_5=>cache_data_out_4_5, 
      out_column_0_4=>cache_data_out_4_4, out_column_0_3=>cache_data_out_4_3, 
      out_column_0_2=>cache_data_out_4_2, out_column_0_1=>cache_data_out_4_1, 
      out_column_0_0=>cache_data_out_4_0, out_column_1_15=>
      cache_data_out_3_15, out_column_1_14=>cache_data_out_3_14, 
      out_column_1_13=>cache_data_out_3_13, out_column_1_12=>
      cache_data_out_3_12, out_column_1_11=>cache_data_out_3_11, 
      out_column_1_10=>cache_data_out_3_10, out_column_1_9=>
      cache_data_out_3_9, out_column_1_8=>cache_data_out_3_8, out_column_1_7
      =>cache_data_out_3_7, out_column_1_6=>cache_data_out_3_6, 
      out_column_1_5=>cache_data_out_3_5, out_column_1_4=>cache_data_out_3_4, 
      out_column_1_3=>cache_data_out_3_3, out_column_1_2=>cache_data_out_3_2, 
      out_column_1_1=>cache_data_out_3_1, out_column_1_0=>cache_data_out_3_0, 
      out_column_2_15=>cache_data_out_2_15, out_column_2_14=>
      cache_data_out_2_14, out_column_2_13=>cache_data_out_2_13, 
      out_column_2_12=>cache_data_out_2_12, out_column_2_11=>
      cache_data_out_2_11, out_column_2_10=>cache_data_out_2_10, 
      out_column_2_9=>cache_data_out_2_9, out_column_2_8=>cache_data_out_2_8, 
      out_column_2_7=>cache_data_out_2_7, out_column_2_6=>cache_data_out_2_6, 
      out_column_2_5=>cache_data_out_2_5, out_column_2_4=>cache_data_out_2_4, 
      out_column_2_3=>cache_data_out_2_3, out_column_2_2=>cache_data_out_2_2, 
      out_column_2_1=>cache_data_out_2_1, out_column_2_0=>cache_data_out_2_0, 
      out_column_3_15=>cache_data_out_1_15, out_column_3_14=>
      cache_data_out_1_14, out_column_3_13=>cache_data_out_1_13, 
      out_column_3_12=>cache_data_out_1_12, out_column_3_11=>
      cache_data_out_1_11, out_column_3_10=>cache_data_out_1_10, 
      out_column_3_9=>cache_data_out_1_9, out_column_3_8=>cache_data_out_1_8, 
      out_column_3_7=>cache_data_out_1_7, out_column_3_6=>cache_data_out_1_6, 
      out_column_3_5=>cache_data_out_1_5, out_column_3_4=>cache_data_out_1_4, 
      out_column_3_3=>cache_data_out_1_3, out_column_3_2=>cache_data_out_1_2, 
      out_column_3_1=>cache_data_out_1_1, out_column_3_0=>cache_data_out_1_0, 
      out_column_4_15=>cache_data_out_0_15, out_column_4_14=>
      cache_data_out_0_14, out_column_4_13=>cache_data_out_0_13, 
      out_column_4_12=>cache_data_out_0_12, out_column_4_11=>
      cache_data_out_0_11, out_column_4_10=>cache_data_out_0_10, 
      out_column_4_9=>cache_data_out_0_9, out_column_4_8=>cache_data_out_0_8, 
      out_column_4_7=>cache_data_out_0_7, out_column_4_6=>cache_data_out_0_6, 
      out_column_4_5=>cache_data_out_0_5, out_column_4_4=>cache_data_out_0_4, 
      out_column_4_3=>cache_data_out_0_3, out_column_4_2=>cache_data_out_0_2, 
      out_column_4_1=>cache_data_out_0_1, out_column_4_0=>cache_data_out_0_0, 
      clk=>nx16767, reset=>cache_rst_actual);
   cache_height_cntr : AdvancedCounter_16 port map ( clk=>clk, reset=>
      nx16751, enable=>cache_height_count_en, mode_in(1)=>wind_rst_EXMPLR, 
      mode_in(0)=>wind_rst_EXMPLR, max_val_in(15)=>wind_rst_EXMPLR, 
      max_val_in(14)=>wind_rst_EXMPLR, max_val_in(13)=>wind_rst_EXMPLR, 
      max_val_in(12)=>wind_rst_EXMPLR, max_val_in(11)=>wind_rst_EXMPLR, 
      max_val_in(10)=>wind_rst_EXMPLR, max_val_in(9)=>wind_rst_EXMPLR, 
      max_val_in(8)=>wind_rst_EXMPLR, max_val_in(7)=>wind_rst_EXMPLR, 
      max_val_in(6)=>wind_rst_EXMPLR, max_val_in(5)=>wind_rst_EXMPLR, 
      max_val_in(4)=>max_height_4, max_val_in(3)=>max_height_3, 
      max_val_in(2)=>max_height_2, max_val_in(1)=>max_height_1, 
      max_val_in(0)=>max_height_0, max_reached_out=>cache_height_ended, 
      counter_out(15)=>DANGLING(0), counter_out(14)=>DANGLING(1), 
      counter_out(13)=>DANGLING(2), counter_out(12)=>DANGLING(3), 
      counter_out(11)=>DANGLING(4), counter_out(10)=>DANGLING(5), 
      counter_out(9)=>DANGLING(6), counter_out(8)=>DANGLING(7), 
      counter_out(7)=>DANGLING(8), counter_out(6)=>DANGLING(9), 
      counter_out(5)=>DANGLING(10), counter_out(4)=>DANGLING(11), 
      counter_out(3)=>DANGLING(12), counter_out(2)=>DANGLING(13), 
      counter_out(1)=>DANGLING(14), counter_out(0)=>DANGLING(15));
   ix12069 : fake_gnd port map ( Y=>wind_rst_EXMPLR);
   ix799 : oai21 port map ( Y=>filter_ready_out_EXMPLR, A0=>nx17097, A1=>
      nx14512, B0=>nx15339);
   reg_current_state_10 : dffr port map ( Q=>OPEN, QB=>nx14508, D=>nx16797, 
      CLK=>nx16767, R=>reset);
   ix14521 : nand04 port map ( Y=>nx14520, A0=>cntr1_inst_counter_out_3, A1
      =>cntr1_inst_counter_out_2, A2=>cntr1_inst_counter_out_1, A3=>
      cntr1_inst_counter_out_0);
   ix14526 : nand03 port map ( Y=>nx14525, A0=>cntr1_inst_counter_out_2, A1
      =>cntr1_inst_counter_out_1, A2=>cntr1_inst_counter_out_0);
   ix14531 : nand02 port map ( Y=>nx14530, A0=>cntr1_inst_counter_out_1, A1
      =>cntr1_inst_counter_out_0);
   reg_cntr1_inst_counter_out_1 : dffr port map ( Q=>
      cntr1_inst_counter_out_1, QB=>nx14534, D=>nx12757, CLK=>clk, R=>
      nx16857);
   ix685 : or02 port map ( Y=>nx684, A0=>nx16753, A1=>nx680);
   reg_current_state_12 : dffr port map ( Q=>current_state_12, QB=>OPEN, D=>
      nx808, CLK=>nx16779, R=>reset);
   ix809 : oai22 port map ( Y=>nx808, A0=>nx17097, A1=>nx794, B0=>nx14564, 
      B1=>nx646);
   ix795 : nand04 port map ( Y=>nx794, A0=>nx14515, A1=>nx14540, A2=>nx14544, 
      A3=>nx14555);
   reg_cntr1_inst_counter_out_2 : dffr port map ( Q=>
      cntr1_inst_counter_out_2, QB=>nx14542, D=>nx12767, CLK=>clk, R=>
      nx16857);
   reg_cntr1_inst_counter_out_5 : dffr port map ( Q=>
      cntr1_inst_counter_out_5, QB=>nx14546, D=>nx12797, CLK=>clk, R=>
      nx16857);
   reg_cntr1_inst_counter_out_4 : dffr port map ( Q=>
      cntr1_inst_counter_out_4, QB=>nx14553, D=>nx12787, CLK=>clk, R=>
      nx16857);
   ix14556 : nor03_2x port map ( Y=>nx14555, A0=>nx728, A1=>nx14561, A2=>
      nx702);
   reg_cntr1_inst_counter_out_0 : dffr port map ( Q=>
      cntr1_inst_counter_out_0, QB=>OPEN, D=>nx12747, CLK=>clk, R=>nx16857);
   ix12748 : xnor2 port map ( Y=>nx12747, A0=>cntr1_inst_counter_out_0, A1=>
      nx17097);
   reg_cntr1_inst_counter_out_3 : dffr port map ( Q=>
      cntr1_inst_counter_out_3, QB=>nx14561, D=>nx12777, CLK=>clk, R=>
      nx16857);
   reg_current_state_9 : dffr port map ( Q=>current_state_9, QB=>nx14564, D
      =>nx670, CLK=>nx16779, R=>reset);
   ix671 : oai21 port map ( Y=>nx670, A0=>nx14567, A1=>nx14715, B0=>nx15329
   );
   ix14568 : nor03_2x port map ( Y=>nx14567, A0=>num_channels_counter_out_0, 
      A1=>num_channels_counter_out_1, A2=>num_channels_counter_out_2);
   ix12608 : mux21 port map ( Y=>nx12607, A0=>nx14571, A1=>nx14573, S0=>
      nx386);
   reg_num_channels_counter_out_0 : dffr port map ( Q=>
      num_channels_counter_out_0, QB=>nx14571, D=>nx12607, CLK=>clk, R=>
      reset);
   ix14574 : aoi221 port map ( Y=>nx14573, A0=>mem_data_in(0), A1=>
      current_state_8, B0=>nflt_layer_temp_0, B1=>nx16841, C0=>nx426);
   reg_current_state_8 : dffr port map ( Q=>current_state_8, QB=>nx15297, D
      =>nx650, CLK=>nx16779, R=>reset);
   ix651 : nor02_2x port map ( Y=>nx650, A0=>nx17103, A1=>nx646);
   reg_current_state_7 : dffr port map ( Q=>OPEN, QB=>nx14577, D=>nx16835, 
      CLK=>nx16779, R=>reset);
   reg_current_state_6 : dffr port map ( Q=>current_state_6, QB=>OPEN, D=>
      current_state_5, CLK=>nx16779, R=>reset);
   reg_current_state_5 : dffr port map ( Q=>current_state_5, QB=>OPEN, D=>
      current_state_4, CLK=>nx16779, R=>reset);
   reg_current_state_4 : dffr port map ( Q=>current_state_4, QB=>OPEN, D=>
      nx16837, CLK=>nx16777, R=>reset);
   reg_current_state_2 : dffr port map ( Q=>current_state_2, QB=>OPEN, D=>
      nx12230, CLK=>nx16777, R=>reset);
   reg_current_state_1 : dffr port map ( Q=>current_state_1, QB=>nx14585, D
      =>current_state_0, CLK=>nx16767, R=>reset);
   reg_current_state_0 : dffs_ni port map ( Q=>current_state_0, QB=>OPEN, D
      =>wind_rst_EXMPLR, CLK=>nx16767, S=>reset);
   ix1257 : oai21 port map ( Y=>nx1256, A0=>nx14597, A1=>nx16783, B0=>
      nx14722);
   ix13128 : mux21_ni port map ( Y=>nx13127, A0=>nx1226, A1=>
      ftc_cntrl_reg_out_14, S0=>nx16953);
   ix1227 : oai22 port map ( Y=>nx1226, A0=>nx14604, A1=>nx14620, B0=>
      nx14606, B1=>nx15231);
   ftc_cntrl_reg_reg_q_14 : dffr port map ( Q=>ftc_cntrl_reg_out_14, QB=>
      nx14606, D=>nx13127, CLK=>nx16767, R=>nx16751);
   ix12808 : mux21_ni port map ( Y=>nx12807, A0=>flt_size_out_0, A1=>
      mem_data_in(0), S0=>current_state_4);
   flt_size_reg_q_0 : dffr port map ( Q=>flt_size_out_0, QB=>OPEN, D=>
      nx12807, CLK=>clk, R=>reset);
   flt_size_reg_q_2 : dffr port map ( Q=>flt_size_out_2, QB=>nx14615, D=>
      nx12817, CLK=>clk, R=>reset);
   ix12818 : mux21_ni port map ( Y=>nx12817, A0=>flt_size_out_2, A1=>
      mem_data_in(2), S0=>current_state_4);
   ix12828 : mux21_ni port map ( Y=>nx12827, A0=>flt_size_out_1, A1=>
      mem_data_in(1), S0=>current_state_4);
   flt_size_reg_q_1 : dffr port map ( Q=>flt_size_out_1, QB=>OPEN, D=>
      nx12827, CLK=>clk, R=>reset);
   ix14621 : aoi21 port map ( Y=>nx14620, A0=>nx16805, A1=>nx14884, B0=>
      current_state_20);
   ix1655 : oai221 port map ( Y=>nx1654, A0=>nx12251, A1=>nx1584, B0=>
      nx14875, B1=>nx15216, C0=>nx15219);
   ix13288 : mux21 port map ( Y=>nx13287, A0=>nx14627, A1=>nx14871, S0=>
      nx16953);
   ix14628 : nand04 port map ( Y=>nx14627, A0=>nx1450, A1=>nx1464, A2=>
      nx1486, A3=>nx1518);
   window_width_cntr_counter_out_15 : dffr port map ( Q=>OPEN, QB=>nx14632, 
      D=>nx13277, CLK=>clk, R=>nx16881);
   ix1279 : nand02 port map ( Y=>nx1278, A0=>nx14635, A1=>nx14873);
   ix14636 : aoi22 port map ( Y=>nx14635, A0=>nx16819, A1=>
      ftc_cntrl_reg_out_13, B0=>nx16805, B1=>ftc_cntrl_reg_out_12);
   ix815 : or02 port map ( Y=>nx814, A0=>nx12239, A1=>nx16753);
   reg_current_state_13 : dffr port map ( Q=>OPEN, QB=>nx14640, D=>nx814, 
      CLK=>nx16767, R=>reset);
   ix12838 : mux21_ni port map ( Y=>nx12837, A0=>cache_height_ended, A1=>
      ftc_cntrl_reg_out_13, S0=>nx16953);
   reg_current_state_19 : dffr port map ( Q=>OPEN, QB=>nx14647, D=>nx1654, 
      CLK=>nx16767, R=>reset);
   reg_current_state_14 : dffr port map ( Q=>current_state_14, QB=>nx14867, 
      D=>nx1266, CLK=>nx16773, R=>reset);
   ix1267 : oai22 port map ( Y=>nx1266, A0=>nx14651, A1=>nx14653, B0=>
      nx17109, B1=>nx14865);
   reg_current_state_23 : dffr port map ( Q=>current_state_23, QB=>nx14651, 
      D=>nx1256, CLK=>nx16769, R=>reset);
   ix14654 : nor04 port map ( Y=>nx14653, A0=>nx374, A1=>nx286, A2=>nx190, 
      A3=>nx96);
   ix375 : nand04 port map ( Y=>nx374, A0=>nx14656, A1=>nx14787, A2=>nx14792, 
      A3=>nx14797);
   ix12578 : oai22 port map ( Y=>nx12577, A0=>nx14660, A1=>nx14717, B0=>
      nx14782, B1=>nx16851);
   reg_write_offset_reg_q_14 : dffr port map ( Q=>write_offset_data_out_14, 
      QB=>nx14663, D=>nx12557, CLK=>nx16769, R=>reset);
   ix14670 : nand02 port map ( Y=>nx14669, A0=>write_offset_data_out_13, A1
      =>nx288);
   ix12538 : oai22 port map ( Y=>nx12537, A0=>nx14673, A1=>nx14717, B0=>
      nx14780, B1=>nx16849);
   ix14674 : oai21 port map ( Y=>nx14673, A0=>nx288, A1=>
      write_offset_data_out_13, B0=>nx14669);
   reg_write_offset_reg_q_12 : dffr port map ( Q=>write_offset_data_out_12, 
      QB=>nx14676, D=>nx12517, CLK=>nx16769, R=>reset);
   ix14683 : nand02 port map ( Y=>nx14682, A0=>write_offset_data_out_11, A1
      =>nx240);
   ix12498 : oai22 port map ( Y=>nx12497, A0=>nx14686, A1=>nx16959, B0=>
      nx14778, B1=>nx16849);
   ix14687 : oai21 port map ( Y=>nx14686, A0=>nx240, A1=>
      write_offset_data_out_11, B0=>nx14682);
   reg_write_offset_reg_q_10 : dffr port map ( Q=>write_offset_data_out_10, 
      QB=>nx14689, D=>nx12477, CLK=>nx16769, R=>reset);
   ix14696 : nand02 port map ( Y=>nx14695, A0=>write_offset_data_out_9, A1=>
      nx194);
   ix12458 : oai22 port map ( Y=>nx12457, A0=>nx14699, A1=>nx16959, B0=>
      nx14776, B1=>nx16849);
   ix14700 : oai21 port map ( Y=>nx14699, A0=>nx194, A1=>
      write_offset_data_out_9, B0=>nx14695);
   reg_write_offset_reg_q_8 : dffr port map ( Q=>write_offset_data_out_8, QB
      =>nx14702, D=>nx12437, CLK=>nx16769, R=>reset);
   ix14709 : nand02 port map ( Y=>nx14708, A0=>write_offset_data_out_7, A1=>
      nx144);
   ix12418 : oai22 port map ( Y=>nx12417, A0=>nx14712, A1=>nx16847, B0=>
      nx14723, B1=>nx16959);
   reg_write_offset_reg_q_7 : dffr port map ( Q=>write_offset_data_out_7, QB
      =>nx14712, D=>nx12417, CLK=>nx16769, R=>reset);
   ix9 : nand02 port map ( Y=>nx8, A0=>nx14715, A1=>nx16957);
   ix14716 : nand02 port map ( Y=>nx14715, A0=>current_state_23, A1=>nx14653
   );
   reg_current_state_21 : dffr port map ( Q=>OPEN, QB=>nx14597, D=>nx1240, 
      CLK=>nx16769, R=>reset);
   reg_current_state_22 : dffr port map ( Q=>OPEN, QB=>nx14722, D=>nx1246, 
      CLK=>nx16771, R=>reset);
   ix14724 : oai21 port map ( Y=>nx14723, A0=>nx144, A1=>
      write_offset_data_out_7, B0=>nx14708);
   reg_write_offset_reg_q_6 : dffr port map ( Q=>write_offset_data_out_6, QB
      =>nx14726, D=>nx12397, CLK=>nx16771, R=>reset);
   ix14733 : nand02 port map ( Y=>nx14732, A0=>write_offset_data_out_5, A1=>
      nx98);
   ix12378 : oai22 port map ( Y=>nx12377, A0=>nx14736, A1=>nx16847, B0=>
      nx14738, B1=>nx16957);
   reg_write_offset_reg_q_5 : dffr port map ( Q=>write_offset_data_out_5, QB
      =>nx14736, D=>nx12377, CLK=>nx16771, R=>reset);
   ix14739 : oai21 port map ( Y=>nx14738, A0=>nx98, A1=>
      write_offset_data_out_5, B0=>nx14732);
   reg_write_offset_reg_q_4 : dffr port map ( Q=>write_offset_data_out_4, QB
      =>nx14741, D=>nx12357, CLK=>nx16771, R=>reset);
   reg_write_offset_reg_q_3 : dffr port map ( Q=>write_offset_data_out_3, QB
      =>nx14751, D=>nx12337, CLK=>nx16771, R=>reset);
   ix12318 : oai22 port map ( Y=>nx12317, A0=>nx14756, A1=>nx16847, B0=>
      nx14759, B1=>nx16957);
   ix14760 : oai21 port map ( Y=>nx14759, A0=>nx26, A1=>
      write_offset_data_out_2, B0=>nx14774);
   ix12298 : oai22 port map ( Y=>nx12297, A0=>nx17803, A1=>nx16847, B0=>
      nx14765, B1=>nx16957);
   ix14766 : oai21 port map ( Y=>nx14765, A0=>write_offset_data_out_0, A1=>
      write_offset_data_out_1, B0=>nx14771);
   reg_write_offset_reg_q_0 : dffr port map ( Q=>write_offset_data_out_0, QB
      =>nx14769, D=>nx12277, CLK=>nx16771, R=>reset);
   reg_write_offset_reg_q_1 : dffr port map ( Q=>write_offset_data_out_1, QB
      =>nx14762, D=>nx12297, CLK=>nx16771, R=>reset);
   reg_write_offset_reg_q_2 : dffr port map ( Q=>write_offset_data_out_2, QB
      =>nx14756, D=>nx12317, CLK=>nx16773, R=>reset);
   reg_write_offset_reg_q_9 : dffr port map ( Q=>write_offset_data_out_9, QB
      =>nx14776, D=>nx12457, CLK=>nx16773, R=>reset);
   reg_write_offset_reg_q_11 : dffr port map ( Q=>write_offset_data_out_11, 
      QB=>nx14778, D=>nx12497, CLK=>nx16773, R=>reset);
   reg_write_offset_reg_q_13 : dffr port map ( Q=>write_offset_data_out_13, 
      QB=>nx14780, D=>nx12537, CLK=>nx16773, R=>reset);
   reg_write_offset_reg_q_15 : dffr port map ( Q=>OPEN, QB=>nx14782, D=>
      nx12577, CLK=>nx16773, R=>reset);
   new_size_squared_reg_q_15 : dffr port map ( Q=>new_size_squared_out_15, 
      QB=>OPEN, D=>nx12587, CLK=>clk, R=>reset);
   new_size_squared_reg_q_14 : dffr port map ( Q=>new_size_squared_out_14, 
      QB=>nx14791, D=>nx12567, CLK=>clk, R=>reset);
   new_size_squared_reg_q_13 : dffr port map ( Q=>new_size_squared_out_13, 
      QB=>OPEN, D=>nx12547, CLK=>clk, R=>reset);
   new_size_squared_reg_q_12 : dffr port map ( Q=>new_size_squared_out_12, 
      QB=>nx14801, D=>nx12527, CLK=>clk, R=>reset);
   ix287 : nand04 port map ( Y=>nx286, A0=>nx14803, A1=>nx14808, A2=>nx14813, 
      A3=>nx14818);
   new_size_squared_reg_q_11 : dffr port map ( Q=>new_size_squared_out_11, 
      QB=>OPEN, D=>nx12507, CLK=>clk, R=>reset);
   new_size_squared_reg_q_10 : dffr port map ( Q=>new_size_squared_out_10, 
      QB=>nx14812, D=>nx12487, CLK=>clk, R=>reset);
   new_size_squared_reg_q_9 : dffr port map ( Q=>new_size_squared_out_9, QB
      =>OPEN, D=>nx12467, CLK=>clk, R=>reset);
   new_size_squared_reg_q_8 : dffr port map ( Q=>new_size_squared_out_8, QB
      =>nx14822, D=>nx12447, CLK=>clk, R=>reset);
   ix191 : nand04 port map ( Y=>nx190, A0=>nx14824, A1=>nx14829, A2=>nx14834, 
      A3=>nx14839);
   new_size_squared_reg_q_7 : dffr port map ( Q=>new_size_squared_out_7, QB
      =>OPEN, D=>nx12427, CLK=>clk, R=>reset);
   new_size_squared_reg_q_6 : dffr port map ( Q=>new_size_squared_out_6, QB
      =>nx14833, D=>nx12407, CLK=>clk, R=>reset);
   new_size_squared_reg_q_5 : dffr port map ( Q=>new_size_squared_out_5, QB
      =>OPEN, D=>nx12387, CLK=>clk, R=>reset);
   new_size_squared_reg_q_4 : dffr port map ( Q=>new_size_squared_out_4, QB
      =>nx14843, D=>nx12367, CLK=>clk, R=>reset);
   ix97 : nand04 port map ( Y=>nx96, A0=>nx14845, A1=>nx14850, A2=>nx14855, 
      A3=>nx14860);
   new_size_squared_reg_q_3 : dffr port map ( Q=>new_size_squared_out_3, QB
      =>OPEN, D=>nx12347, CLK=>clk, R=>reset);
   new_size_squared_reg_q_2 : dffr port map ( Q=>new_size_squared_out_2, QB
      =>nx14854, D=>nx12327, CLK=>clk, R=>reset);
   new_size_squared_reg_q_1 : dffr port map ( Q=>new_size_squared_out_1, QB
      =>OPEN, D=>nx12307, CLK=>clk, R=>reset);
   new_size_squared_reg_q_0 : dffr port map ( Q=>new_size_squared_out_0, QB
      =>OPEN, D=>nx12287, CLK=>clk, R=>reset);
   ftc_cntrl_reg_reg_q_13 : dffr port map ( Q=>ftc_cntrl_reg_out_13, QB=>
      nx14865, D=>nx12837, CLK=>nx16773, R=>nx16751);
   ix1557 : nand02 port map ( Y=>nx1556, A0=>nx17071, A1=>nx14873);
   ftc_cntrl_reg_reg_q_11 : dffr port map ( Q=>ftc_cntrl_reg_out_11, QB=>
      nx14871, D=>nx13287, CLK=>nx16775, R=>nx16751);
   ix13308 : mux21 port map ( Y=>nx13307, A0=>nx14878, A1=>nx14875, S0=>
      nx16953);
   ix14879 : aoi32 port map ( Y=>nx14878, A0=>nx14604, A1=>
      ftc_cntrl_reg_out_11, A2=>current_state_20, B0=>ftc_cntrl_reg_out_8, 
      B1=>nx1576);
   ix13118 : mux21 port map ( Y=>nx13117, A0=>nx14887, A1=>nx14884, S0=>
      nx16953);
   ix14888 : nand04 port map ( Y=>nx14887, A0=>nx1052, A1=>nx1066, A2=>
      nx1098, A3=>nx1196);
   cache_width_cntr_counter_out_15 : dffr port map ( Q=>OPEN, QB=>nx14892, D
      =>nx13007, CLK=>clk, R=>nx16867);
   ix875 : nand02 port map ( Y=>nx874, A0=>nx14895, A1=>nx14899);
   ix14896 : aoi21 port map ( Y=>nx14895, A0=>nx14897, A1=>nx16819, B0=>
      nx16751);
   ftc_cntrl_reg_reg_q_12 : dffr port map ( Q=>ftc_cntrl_reg_out_12, QB=>
      nx14884, D=>nx13117, CLK=>nx16775, R=>nx16751);
   reg_cache_width_cntr_counter_out_14 : dffr port map ( Q=>
      cache_width_cntr_counter_out_14, QB=>nx14905, D=>nx12997, CLK=>clk, R
      =>nx16867);
   ix14911 : nand02 port map ( Y=>nx14910, A0=>
      cache_width_cntr_counter_out_13, A1=>nx12243);
   reg_cache_width_cntr_counter_out_13 : dffr port map ( Q=>
      cache_width_cntr_counter_out_13, QB=>nx14914, D=>nx12987, CLK=>clk, R
      =>nx16867);
   ix14917 : oai21 port map ( Y=>nx14916, A0=>nx12243, A1=>
      cache_width_cntr_counter_out_13, B0=>nx14910);
   reg_cache_width_cntr_counter_out_12 : dffr port map ( Q=>
      cache_width_cntr_counter_out_12, QB=>nx14919, D=>nx12977, CLK=>clk, R
      =>nx16867);
   ix14925 : nand02 port map ( Y=>nx14924, A0=>
      cache_width_cntr_counter_out_11, A1=>nx12245);
   reg_cache_width_cntr_counter_out_11 : dffr port map ( Q=>
      cache_width_cntr_counter_out_11, QB=>nx14928, D=>nx12967, CLK=>clk, R
      =>nx16867);
   ix14931 : oai21 port map ( Y=>nx14930, A0=>nx12245, A1=>
      cache_width_cntr_counter_out_11, B0=>nx14924);
   reg_cache_width_cntr_counter_out_10 : dffr port map ( Q=>
      cache_width_cntr_counter_out_10, QB=>nx14933, D=>nx12957, CLK=>clk, R
      =>nx16867);
   ix14939 : nand02 port map ( Y=>nx14938, A0=>
      cache_width_cntr_counter_out_9, A1=>nx12247);
   reg_cache_width_cntr_counter_out_9 : dffr port map ( Q=>
      cache_width_cntr_counter_out_9, QB=>nx14942, D=>nx12947, CLK=>clk, R=>
      nx16867);
   ix14945 : oai21 port map ( Y=>nx14944, A0=>nx12247, A1=>
      cache_width_cntr_counter_out_9, B0=>nx14938);
   reg_cache_width_cntr_counter_out_8 : dffr port map ( Q=>
      cache_width_cntr_counter_out_8, QB=>nx14947, D=>nx12937, CLK=>clk, R=>
      nx16869);
   ix14953 : nand02 port map ( Y=>nx14952, A0=>
      cache_width_cntr_counter_out_7, A1=>nx12249);
   reg_cache_width_cntr_counter_out_7 : dffr port map ( Q=>
      cache_width_cntr_counter_out_7, QB=>nx14956, D=>nx12927, CLK=>clk, R=>
      nx16869);
   ix14959 : oai21 port map ( Y=>nx14958, A0=>nx12249, A1=>
      cache_width_cntr_counter_out_7, B0=>nx14952);
   reg_cache_width_cntr_counter_out_6 : dffr port map ( Q=>
      cache_width_cntr_counter_out_6, QB=>nx14961, D=>nx12917, CLK=>clk, R=>
      nx16869);
   reg_cache_width_count_4 : dffr port map ( Q=>cache_width_count_4, QB=>
      OPEN, D=>nx12897, CLK=>clk, R=>nx16871);
   ix905 : xnor2 port map ( Y=>nx904, A0=>nx16759, A1=>nx14971);
   ix14972 : nand04 port map ( Y=>nx14971, A0=>cache_width_count_1, A1=>
      cache_width_count_0, A2=>nx16763, A3=>cache_width_count_3);
   reg_cache_width_count_1 : dffr port map ( Q=>cache_width_count_1, QB=>
      OPEN, D=>nx12867, CLK=>clk, R=>nx16869);
   ix881 : xor2 port map ( Y=>nx880, A0=>cache_width_count_1, A1=>
      cache_width_count_0);
   reg_cache_width_count_0 : dffr port map ( Q=>cache_width_count_0, QB=>
      OPEN, D=>nx12857, CLK=>clk, R=>nx16869);
   ix12848 : mux21_ni port map ( Y=>nx12847, A0=>nx856, A1=>
      ftc_cntrl_reg_out_10, S0=>nx16953);
   ix857 : oai21 port map ( Y=>nx856, A0=>nx14983, A1=>nx14985, B0=>nx14990
   );
   ftc_cntrl_reg_reg_q_10 : dffr port map ( Q=>ftc_cntrl_reg_out_10, QB=>
      nx14983, D=>nx12847, CLK=>nx16775, R=>nx16751);
   ix845 : nor03_2x port map ( Y=>cache_height_count_en, A0=>nx14988, A1=>
      ftc_cntrl_reg_out_13, A2=>nx14884);
   ix14991 : aoi21 port map ( Y=>nx14990, A0=>nx16803, A1=>nx14884, B0=>
      nx830);
   ix831 : nor03_2x port map ( Y=>nx830, A0=>ftc_cntrl_reg_out_12, A1=>
      nx17109, A2=>ftc_cntrl_reg_out_13);
   reg_cache_width_count_2 : dffr port map ( Q=>cache_width_count_2, QB=>
      OPEN, D=>nx12877, CLK=>clk, R=>nx16869);
   ix889 : xnor2 port map ( Y=>nx888, A0=>nx16763, A1=>nx15000);
   ix15001 : nand02 port map ( Y=>nx15000, A0=>cache_width_count_1, A1=>
      cache_width_count_0);
   reg_cache_width_count_3 : dffr port map ( Q=>cache_width_count_3, QB=>
      OPEN, D=>nx12887, CLK=>clk, R=>nx16869);
   ix897 : xnor2 port map ( Y=>nx896, A0=>cache_width_count_3, A1=>nx15006);
   ix15007 : nand03 port map ( Y=>nx15006, A0=>cache_width_count_1, A1=>
      cache_width_count_0, A2=>nx16765);
   reg_cache_width_cntr_counter_out_5 : dffr port map ( Q=>
      cache_width_cntr_counter_out_5, QB=>nx15012, D=>nx12907, CLK=>clk, R=>
      nx16871);
   ix15015 : oai21 port map ( Y=>nx15014, A0=>nx910, A1=>
      cache_width_cntr_counter_out_5, B0=>nx14966);
   ix911 : nor02ii port map ( Y=>nx910, A0=>nx14971, A1=>nx16761);
   img_width_reg_q_0 : dffr port map ( Q=>img_width_out_0, QB=>nx15029, D=>
      nx13027, CLK=>clk, R=>reset);
   reg_current_state_24 : dffr port map ( Q=>current_state_24, QB=>OPEN, D=>
      nx600, CLK=>nx16775, R=>reset);
   new_width_reg_q_0 : dffr port map ( Q=>new_width_out_0, QB=>OPEN, D=>
      nx13017, CLK=>clk, R=>reset);
   ix13018 : mux21_ni port map ( Y=>nx13017, A0=>new_width_out_0, A1=>
      mem_data_in(0), S0=>current_state_5);
   ix1197 : nor04 port map ( Y=>nx1196, A0=>nx1120, A1=>nx1144, A2=>nx1172, 
      A3=>nx1188);
   ix1121 : xnor2 port map ( Y=>nx1120, A0=>cache_width_count_1, A1=>nx16961
   );
   ix15033 : aoi21 port map ( Y=>nx15032, A0=>img_width_out_1, A1=>
      img_width_out_0, B0=>nx15040);
   img_width_reg_q_1 : dffr port map ( Q=>img_width_out_1, QB=>OPEN, D=>
      nx13047, CLK=>clk, R=>reset);
   ix13048 : ao22 port map ( Y=>nx13047, A0=>nx16841, A1=>new_width_out_1, 
      B0=>img_width_out_1, B1=>nx15027);
   new_width_reg_q_1 : dffr port map ( Q=>new_width_out_1, QB=>OPEN, D=>
      nx13037, CLK=>clk, R=>reset);
   ix13038 : mux21_ni port map ( Y=>nx13037, A0=>new_width_out_1, A1=>
      mem_data_in(1), S0=>current_state_5);
   ix1145 : xnor2 port map ( Y=>nx1144, A0=>nx16765, A1=>nx15043);
   ix15044 : aoi21 port map ( Y=>nx15043, A0=>img_width_out_2, A1=>nx1112, 
      B0=>nx15052);
   img_width_reg_q_2 : dffs_ni port map ( Q=>img_width_out_2, QB=>OPEN, D=>
      nx13067, CLK=>clk, S=>reset);
   ix13068 : ao221 port map ( Y=>nx13067, A0=>nx16841, A1=>new_width_out_2, 
      B0=>img_width_out_2, B1=>nx15027, C0=>current_state_8);
   new_width_reg_q_2 : dffr port map ( Q=>new_width_out_2, QB=>OPEN, D=>
      nx13057, CLK=>clk, R=>reset);
   ix13058 : mux21_ni port map ( Y=>nx13057, A0=>new_width_out_2, A1=>
      mem_data_in(2), S0=>current_state_5);
   ix15053 : nor03_2x port map ( Y=>nx15052, A0=>img_width_out_0, A1=>
      img_width_out_1, A2=>img_width_out_2);
   ix1173 : xnor2 port map ( Y=>nx1172, A0=>cache_width_count_3, A1=>nx15055
   );
   ix15056 : xnor2 port map ( Y=>nx15055, A0=>img_width_out_3, A1=>nx15052);
   img_width_reg_q_3 : dffs_ni port map ( Q=>img_width_out_3, QB=>OPEN, D=>
      nx13087, CLK=>clk, S=>reset);
   ix13088 : ao22 port map ( Y=>nx13087, A0=>nx16841, A1=>new_width_out_3, 
      B0=>img_width_out_3, B1=>nx15027);
   new_width_reg_q_3 : dffr port map ( Q=>new_width_out_3, QB=>OPEN, D=>
      nx13077, CLK=>clk, R=>reset);
   ix13078 : mux21_ni port map ( Y=>nx13077, A0=>new_width_out_3, A1=>
      mem_data_in(3), S0=>current_state_5);
   ix1189 : xnor2 port map ( Y=>nx1188, A0=>nx16761, A1=>nx15064);
   ix15065 : xnor2 port map ( Y=>nx15064, A0=>img_width_out_4, A1=>nx15072);
   img_width_reg_q_4 : dffs_ni port map ( Q=>img_width_out_4, QB=>OPEN, D=>
      nx13107, CLK=>clk, S=>reset);
   ix13108 : ao22 port map ( Y=>nx13107, A0=>nx16841, A1=>new_width_out_4, 
      B0=>img_width_out_4, B1=>nx15027);
   new_width_reg_q_4 : dffr port map ( Q=>new_width_out_4, QB=>OPEN, D=>
      nx13097, CLK=>clk, R=>reset);
   ix13098 : mux21_ni port map ( Y=>nx13097, A0=>new_width_out_4, A1=>
      mem_data_in(4), S0=>current_state_5);
   ix15073 : nor04 port map ( Y=>nx15072, A0=>img_width_out_0, A1=>
      img_width_out_1, A2=>img_width_out_2, A3=>img_width_out_3);
   ftc_cntrl_reg_reg_q_8 : dffr port map ( Q=>ftc_cntrl_reg_out_8, QB=>
      nx14875, D=>nx13307, CLK=>nx16775, R=>nx16753);
   reg_current_state_20 : dffr port map ( Q=>current_state_20, QB=>nx15075, 
      D=>nx12266, CLK=>nx16775, R=>reset);
   ix15078 : nand03 port map ( Y=>nx15077, A0=>flt_size_out_0, A1=>nx14615, 
      A2=>flt_size_out_1);
   ix1577 : nand02 port map ( Y=>nx1576, A0=>nx15080, A1=>nx15082);
   ix15081 : oai21 port map ( Y=>nx15080, A0=>nx16803, A1=>nx15075, B0=>
      nx14899);
   ix15083 : aoi43 port map ( Y=>nx15082, A0=>nx16803, A1=>nx14884, A2=>
      nx14875, A3=>nx14604, B0=>current_state_20, B1=>nx14606, B2=>nx16783);
   ix13298 : mux21_ni port map ( Y=>nx13297, A0=>nx1542, A1=>
      ftc_cntrl_reg_out_9, S0=>nx16953);
   ix1543 : oai21 port map ( Y=>nx1542, A0=>nx15087, A1=>nx15089, B0=>
      nx14635);
   ftc_cntrl_reg_reg_q_9 : dffr port map ( Q=>ftc_cntrl_reg_out_9, QB=>
      nx15087, D=>nx13297, CLK=>nx16775, R=>nx16753);
   ix15090 : aoi21 port map ( Y=>nx15089, A0=>nx17071, A1=>nx1534, B0=>
      nx16819);
   reg_current_state_15 : dffr port map ( Q=>current_state_15, QB=>nx15092, 
      D=>nx1556, CLK=>nx16777, R=>reset);
   reg_window_width_cntr_counter_out_14 : dffr port map ( Q=>
      window_width_cntr_counter_out_14, QB=>nx15097, D=>nx13267, CLK=>clk, R
      =>nx16881);
   ix15103 : nand02 port map ( Y=>nx15102, A0=>
      window_width_cntr_counter_out_13, A1=>nx12256);
   reg_window_width_cntr_counter_out_13 : dffr port map ( Q=>
      window_width_cntr_counter_out_13, QB=>nx15106, D=>nx13257, CLK=>clk, R
      =>nx16881);
   ix15109 : oai21 port map ( Y=>nx15108, A0=>nx12256, A1=>
      window_width_cntr_counter_out_13, B0=>nx15102);
   reg_window_width_cntr_counter_out_12 : dffr port map ( Q=>
      window_width_cntr_counter_out_12, QB=>nx15111, D=>nx13247, CLK=>clk, R
      =>nx16881);
   ix15117 : nand02 port map ( Y=>nx15116, A0=>
      window_width_cntr_counter_out_11, A1=>nx12258);
   reg_window_width_cntr_counter_out_11 : dffr port map ( Q=>
      window_width_cntr_counter_out_11, QB=>nx15120, D=>nx13237, CLK=>clk, R
      =>nx16881);
   ix15123 : oai21 port map ( Y=>nx15122, A0=>nx12258, A1=>
      window_width_cntr_counter_out_11, B0=>nx15116);
   reg_window_width_cntr_counter_out_10 : dffr port map ( Q=>
      window_width_cntr_counter_out_10, QB=>nx15125, D=>nx13227, CLK=>clk, R
      =>nx16881);
   ix15131 : nand02 port map ( Y=>nx15130, A0=>
      window_width_cntr_counter_out_9, A1=>nx12260);
   reg_window_width_cntr_counter_out_9 : dffr port map ( Q=>
      window_width_cntr_counter_out_9, QB=>nx15134, D=>nx13217, CLK=>clk, R
      =>nx16881);
   ix15137 : oai21 port map ( Y=>nx15136, A0=>nx12260, A1=>
      window_width_cntr_counter_out_9, B0=>nx15130);
   reg_window_width_cntr_counter_out_8 : dffr port map ( Q=>
      window_width_cntr_counter_out_8, QB=>nx15139, D=>nx13207, CLK=>clk, R
      =>nx16883);
   ix15145 : nand02 port map ( Y=>nx15144, A0=>
      window_width_cntr_counter_out_7, A1=>nx12262);
   reg_window_width_cntr_counter_out_7 : dffr port map ( Q=>
      window_width_cntr_counter_out_7, QB=>nx15148, D=>nx13197, CLK=>clk, R
      =>nx16883);
   ix15151 : oai21 port map ( Y=>nx15150, A0=>nx12262, A1=>
      window_width_cntr_counter_out_7, B0=>nx15144);
   reg_window_width_cntr_counter_out_6 : dffr port map ( Q=>
      window_width_cntr_counter_out_6, QB=>nx15153, D=>nx13187, CLK=>clk, R
      =>nx16883);
   reg_wind_width_count_4 : dffr port map ( Q=>wind_width_count_4, QB=>OPEN, 
      D=>nx13317, CLK=>clk, R=>nx16885);
   ix1693 : xnor2 port map ( Y=>nx1692, A0=>wind_width_count_4, A1=>nx15163
   );
   ix15164 : nand04 port map ( Y=>nx15163, A0=>wind_width_count_1, A1=>
      nx16755, A2=>wind_width_count_2, A3=>wind_width_count_3);
   reg_wind_width_count_1 : dffr port map ( Q=>wind_width_count_1, QB=>OPEN, 
      D=>nx13147, CLK=>clk, R=>nx16883);
   ix1285 : xor2 port map ( Y=>nx1284, A0=>wind_width_count_1, A1=>nx16755);
   reg_wind_width_count_0 : dffr port map ( Q=>wind_width_count_0, QB=>OPEN, 
      D=>nx13137, CLK=>clk, R=>nx16883);
   ix1691 : oai22 port map ( Y=>nx12253, A0=>ftc_cntrl_reg_out_9, A1=>
      nx17071, B0=>nx15075, B1=>ftc_cntrl_reg_out_11);
   reg_wind_width_count_2 : dffr port map ( Q=>wind_width_count_2, QB=>OPEN, 
      D=>nx13157, CLK=>clk, R=>nx16883);
   ix1293 : xnor2 port map ( Y=>nx1292, A0=>wind_width_count_2, A1=>nx15180
   );
   ix15181 : nand02 port map ( Y=>nx15180, A0=>wind_width_count_1, A1=>
      nx16757);
   reg_wind_width_count_3 : dffr port map ( Q=>wind_width_count_3, QB=>OPEN, 
      D=>nx13167, CLK=>clk, R=>nx16883);
   ix1301 : xnor2 port map ( Y=>nx1300, A0=>wind_width_count_3, A1=>nx15186
   );
   ix15187 : nand03 port map ( Y=>nx15186, A0=>wind_width_count_1, A1=>
      nx16757, A2=>wind_width_count_2);
   reg_window_width_cntr_counter_out_5 : dffr port map ( Q=>
      window_width_cntr_counter_out_5, QB=>nx15192, D=>nx13177, CLK=>clk, R
      =>nx16885);
   ix15195 : oai21 port map ( Y=>nx15194, A0=>nx1308, A1=>
      window_width_cntr_counter_out_5, B0=>nx15158);
   ix1309 : nor02ii port map ( Y=>nx1308, A0=>nx15163, A1=>
      wind_width_count_4);
   ix1479 : xnor2 port map ( Y=>nx1478, A0=>nx15201, A1=>nx16757);
   ix15202 : nand02 port map ( Y=>nx15201, A0=>nx15029, A1=>nx17071);
   ix1519 : and04 port map ( Y=>nx1518, A0=>nx15204, A1=>nx15207, A2=>
      nx15210, A3=>nx15213);
   ix15205 : xnor2 port map ( Y=>nx15204, A0=>wind_width_count_1, A1=>nx1488
   );
   ix15208 : xnor2 port map ( Y=>nx15207, A0=>wind_width_count_2, A1=>nx1494
   );
   ix1495 : nand02 port map ( Y=>nx1494, A0=>nx17071, A1=>nx15043);
   ix15211 : xnor2 port map ( Y=>nx15210, A0=>wind_width_count_3, A1=>nx1504
   );
   ix15214 : xnor2 port map ( Y=>nx15213, A0=>wind_width_count_4, A1=>nx1508
   );
   ix15220 : aoi22 port map ( Y=>nx15219, A0=>comp_unit_finished, A1=>
      current_state_18, B0=>nx12251, B1=>nx12267);
   ix1645 : oai221 port map ( Y=>nx1644, A0=>nx17129, A1=>nx16783, B0=>
      comp_unit_finished, B1=>nx15226, C0=>nx16963);
   reg_current_state_16 : dffr port map ( Q=>OPEN, QB=>nx15223, D=>nx1622, 
      CLK=>nx16777, R=>reset);
   reg_current_state_18 : dffr port map ( Q=>current_state_18, QB=>nx15226, 
      D=>nx1644, CLK=>nx16777, R=>reset);
   reg_current_state_17 : dffr port map ( Q=>current_state_17, QB=>OPEN, D=>
      nx1628, CLK=>nx16777, R=>reset);
   ix15232 : aoi22 port map ( Y=>nx15231, A0=>nx16819, A1=>nx14865, B0=>
      nx15075, B1=>nx14988);
   ix12658 : mux21_ni port map ( Y=>nx12657, A0=>
      nflt_layer_cntr_counter_out_0, A1=>nx506, S0=>nx496);
   ix497 : oai21 port map ( Y=>nx496, A0=>nx15240, A1=>nx16947, B0=>nx17135
   );
   ix15241 : nor04 port map ( Y=>nx15240, A0=>nx15242, A1=>
      nflt_layer_cntr_counter_out_1, A2=>nflt_layer_cntr_counter_out_2, A3=>
      nflt_layer_cntr_counter_out_3);
   reg_nflt_layer_cntr_counter_out_0 : dffr port map ( Q=>
      nflt_layer_cntr_counter_out_0, QB=>nx15242, D=>nx12657, CLK=>clk, R=>
      reset);
   reg_nflt_layer_cntr_counter_out_1 : dffr port map ( Q=>
      nflt_layer_cntr_counter_out_1, QB=>OPEN, D=>nx12667, CLK=>clk, R=>
      reset);
   ix12668 : mux21_ni port map ( Y=>nx12667, A0=>
      nflt_layer_cntr_counter_out_1, A1=>nx524, S0=>nx496);
   ix15248 : aoi21 port map ( Y=>nx15247, A0=>nflt_layer_cntr_counter_out_1, 
      A1=>nflt_layer_cntr_counter_out_0, B0=>nx15249);
   ix15252 : inv01 port map ( Y=>nx15251, A=>mem_data_in(1));
   reg_nflt_layer_cntr_counter_out_2 : dffr port map ( Q=>
      nflt_layer_cntr_counter_out_2, QB=>OPEN, D=>nx12677, CLK=>clk, R=>
      reset);
   ix12678 : mux21_ni port map ( Y=>nx12677, A0=>
      nflt_layer_cntr_counter_out_2, A1=>nx544, S0=>nx496);
   ix15258 : xnor2 port map ( Y=>nx15257, A0=>nflt_layer_cntr_counter_out_2, 
      A1=>nx15249);
   ix15260 : inv01 port map ( Y=>nx15259, A=>mem_data_in(2));
   reg_nflt_layer_cntr_counter_out_3 : dffr port map ( Q=>
      nflt_layer_cntr_counter_out_3, QB=>OPEN, D=>nx12687, CLK=>clk, R=>
      reset);
   ix12688 : mux21_ni port map ( Y=>nx12687, A0=>
      nflt_layer_cntr_counter_out_3, A1=>nx560, S0=>nx496);
   ix15266 : xnor2 port map ( Y=>nx15265, A0=>nflt_layer_cntr_counter_out_3, 
      A1=>nx15267);
   ix15268 : nor03_2x port map ( Y=>nx15267, A0=>
      nflt_layer_cntr_counter_out_0, A1=>nflt_layer_cntr_counter_out_1, A2=>
      nflt_layer_cntr_counter_out_2);
   ix15270 : inv01 port map ( Y=>nx15269, A=>mem_data_in(3));
   reg_current_state_3 : dffr port map ( Q=>OPEN, QB=>nx15272, D=>
      current_state_2, CLK=>nx16777, R=>reset);
   ix15275 : nor03_2x port map ( Y=>nx15274, A0=>nlayers_counter_out_1, A1=>
      nlayers_counter_out_2, A2=>nlayers_counter_out_0);
   nlayers_reg_counter_data_1 : dffr port map ( Q=>nlayers_counter_out_1, QB
      =>OPEN, D=>nx12717, CLK=>clk, R=>reset);
   nlayers_reg_counter_data_2 : dffr port map ( Q=>nlayers_counter_out_2, QB
      =>OPEN, D=>nx12707, CLK=>clk, R=>reset);
   nlayers_reg_counter_data_0 : dffr port map ( Q=>nlayers_counter_out_0, QB
      =>OPEN, D=>nx12697, CLK=>clk, R=>reset);
   ix647 : nand02 port map ( Y=>nx646, A0=>comp_unit_operation_EXMPLR, A1=>
      nx15293);
   layer_type_reg_q_0 : dffr port map ( Q=>comp_unit_operation_EXMPLR, QB=>
      OPEN, D=>nx12737, CLK=>clk, R=>reset);
   ix12738 : mux21_ni port map ( Y=>nx12737, A0=>comp_unit_operation_EXMPLR, 
      A1=>mem_data_in(0), S0=>current_state_2);
   ix12728 : mux21_ni port map ( Y=>nx12727, A0=>layer_type_out_1, A1=>
      mem_data_in(1), S0=>current_state_2);
   layer_type_reg_q_1 : dffr port map ( Q=>layer_type_out_1, QB=>nx15293, D
      =>nx12727, CLK=>clk, R=>reset);
   nflt_layer_total_reg_q_0 : dffr port map ( Q=>nflt_layer_temp_0, QB=>OPEN, 
      D=>nx12597, CLK=>clk, R=>reset);
   ix387 : oai21 port map ( Y=>nx386, A0=>nx14567, A1=>nx14715, B0=>nx15304
   );
   reg_num_channels_counter_out_1 : dffr port map ( Q=>
      num_channels_counter_out_1, QB=>OPEN, D=>nx12627, CLK=>clk, R=>reset);
   ix12628 : mux21_ni port map ( Y=>nx12627, A0=>num_channels_counter_out_1, 
      A1=>nx454, S0=>nx386);
   ix455 : oai222 port map ( Y=>nx454, A0=>nx4, A1=>nx15309, B0=>nx15313, B1
      =>nx16941, C0=>nx15251, C1=>nx15297);
   ix15310 : aoi21 port map ( Y=>nx15309, A0=>num_channels_counter_out_1, A1
      =>num_channels_counter_out_0, B0=>nx15311);
   nflt_layer_total_reg_q_1 : dffr port map ( Q=>nflt_layer_temp_1, QB=>
      nx15313, D=>nx12617, CLK=>clk, R=>reset);
   ix12648 : mux21 port map ( Y=>nx12647, A0=>nx15320, A1=>nx15322, S0=>
      nx386);
   reg_num_channels_counter_out_2 : dffr port map ( Q=>
      num_channels_counter_out_2, QB=>nx15320, D=>nx12647, CLK=>clk, R=>
      reset);
   ix15323 : aoi222 port map ( Y=>nx15322, A0=>nflt_layer_temp_2, A1=>
      nx16843, B0=>mem_data_in(2), B1=>current_state_8, C0=>nx15304, C1=>
      nx466);
   nflt_layer_total_reg_q_2 : dffr port map ( Q=>nflt_layer_temp_2, QB=>OPEN, 
      D=>nx12637, CLK=>clk, R=>reset);
   ix467 : oai21 port map ( Y=>nx466, A0=>nx15320, A1=>nx15311, B0=>nx12231
   );
   reg_current_state_11 : dffr port map ( Q=>OPEN, QB=>nx15329, D=>nx662, 
      CLK=>nx16779, R=>reset);
   ix663 : oai221 port map ( Y=>nx662, A0=>nx15240, A1=>nx16947, B0=>nx17103, 
      B1=>nx15332, C0=>nx15297);
   ix15337 : oai21 port map ( Y=>nx15336, A0=>cntr1_inst_counter_out_0, A1=>
      cntr1_inst_counter_out_1, B0=>nx14530);
   ix15340 : nand02 port map ( Y=>nx15339, A0=>current_state_9, A1=>nx646);
   ix1755 : nand02 port map ( Y=>nx1754, A0=>nx15344, A1=>nx17139);
   ix15345 : nand03 port map ( Y=>nx15344, A0=>nx17069, A1=>nx15240, A2=>
      nx15274);
   ix15348 : nand02 port map ( Y=>nx15347, A0=>current_state_25, A1=>nx1742
   );
   reg_current_state_25 : dffr port map ( Q=>current_state_25, QB=>nx15353, 
      D=>nx1754, CLK=>nx16781, R=>reset);
   reg_class_cntr_counter_out_0 : dffr port map ( Q=>
      class_cntr_counter_out_0, QB=>nx15350, D=>nx13327, CLK=>clk, R=>reset
   );
   reg_class_cntr_counter_out_1 : dffr port map ( Q=>
      class_cntr_counter_out_1, QB=>nx15358, D=>nx13337, CLK=>clk, R=>reset
   );
   ix15361 : oai21 port map ( Y=>nx15360, A0=>class_cntr_counter_out_0, A1=>
      class_cntr_counter_out_1, B0=>nx15362);
   reg_class_cntr_counter_out_2 : dffr port map ( Q=>
      class_cntr_counter_out_2, QB=>nx15364, D=>nx13347, CLK=>clk, R=>reset
   );
   reg_class_cntr_counter_out_3 : dffr port map ( Q=>
      class_cntr_counter_out_3, QB=>nx15374, D=>nx13357, CLK=>clk, R=>reset
   );
   reg_flt_bias1_reg_q_0 : dff port map ( Q=>flt_bias_out_0, QB=>OPEN, D=>
      nx13377, CLK=>clk);
   ix13368 : nand02 port map ( Y=>nx13367, A0=>nx17149, A1=>nx15329);
   channel_zero_reg_q_0 : dffr port map ( Q=>OPEN, QB=>nx15399, D=>nx13367, 
      CLK=>clk, R=>reset);
   reg_flt_bias1_reg_q_1 : dff port map ( Q=>flt_bias_out_1, QB=>OPEN, D=>
      nx13397, CLK=>clk);
   reg_flt_bias1_reg_q_2 : dff port map ( Q=>flt_bias_out_2, QB=>OPEN, D=>
      nx13417, CLK=>clk);
   reg_flt_bias1_reg_q_3 : dff port map ( Q=>flt_bias_out_3, QB=>OPEN, D=>
      nx13437, CLK=>clk);
   reg_flt_bias1_reg_q_4 : dff port map ( Q=>flt_bias_out_4, QB=>OPEN, D=>
      nx13457, CLK=>clk);
   reg_flt_bias1_reg_q_5 : dff port map ( Q=>flt_bias_out_5, QB=>OPEN, D=>
      nx13477, CLK=>clk);
   reg_flt_bias1_reg_q_6 : dff port map ( Q=>flt_bias_out_6, QB=>OPEN, D=>
      nx13497, CLK=>clk);
   reg_flt_bias1_reg_q_7 : dff port map ( Q=>flt_bias_out_7, QB=>OPEN, D=>
      nx13517, CLK=>clk);
   reg_flt_bias1_reg_q_8 : dff port map ( Q=>flt_bias_out_8, QB=>OPEN, D=>
      nx13537, CLK=>clk);
   reg_flt_bias1_reg_q_9 : dff port map ( Q=>flt_bias_out_9, QB=>OPEN, D=>
      nx13557, CLK=>clk);
   reg_flt_bias1_reg_q_10 : dff port map ( Q=>flt_bias_out_10, QB=>OPEN, D=>
      nx13577, CLK=>clk);
   reg_flt_bias1_reg_q_11 : dff port map ( Q=>flt_bias_out_11, QB=>OPEN, D=>
      nx13597, CLK=>clk);
   reg_flt_bias1_reg_q_12 : dff port map ( Q=>flt_bias_out_12, QB=>OPEN, D=>
      nx13617, CLK=>clk);
   reg_flt_bias1_reg_q_13 : dff port map ( Q=>flt_bias_out_13, QB=>OPEN, D=>
      nx13637, CLK=>clk);
   reg_flt_bias1_reg_q_14 : dff port map ( Q=>flt_bias_out_14, QB=>OPEN, D=>
      nx13657, CLK=>clk);
   reg_flt_bias1_reg_q_15 : dff port map ( Q=>flt_bias_out_15, QB=>OPEN, D=>
      nx13677, CLK=>clk);
   ix4611 : aoi21 port map ( Y=>comp_unit_relu, A0=>nx17129, A1=>nx16967, B0
      =>nx12231);
   ix4773 : nor02_2x port map ( Y=>max_height_1, A0=>nx17113, A1=>nx16961);
   ix4487 : or02 port map ( Y=>cache_rst_actual, A0=>nx16753, A1=>reset);
   ix2445 : oai321 port map ( Y=>cache_load, A0=>ftc_cntrl_reg_out_12, A1=>
      nx17109, A2=>ftc_cntrl_reg_out_13, B0=>nx17113, B1=>nx15480, C0=>
      nx14882);
   ix13698 : mux21 port map ( Y=>nx13697, A0=>nx15483, A1=>nx15480, S0=>
      nx16955);
   ix15484 : aoi32 port map ( Y=>nx15483, A0=>nx1200, A1=>cache_height_ended, 
      A2=>nx16805, B0=>ftc_cntrl_reg_out_15, B1=>nx2392);
   ftc_cntrl_reg_reg_q_15 : dffr port map ( Q=>ftc_cntrl_reg_out_15, QB=>
      nx15480, D=>nx13697, CLK=>nx16781, R=>nx16753);
   ix2393 : nand03 port map ( Y=>nx2392, A0=>ftc_cntrl_reg_out_13, A1=>
      nx17113, A2=>nx16821);
   ix15490 : aoi21 port map ( Y=>nx15489, A0=>nx15480, A1=>nx12267, B0=>
      nx830);
   ix2451 : oai21 port map ( Y=>max_height_0, A0=>nx17113, A1=>
      img_width_out_0, B0=>nx15531);
   ix4777 : nand02 port map ( Y=>max_height_2, A0=>nx15043, A1=>nx16805);
   ix1979 : oai21 port map ( Y=>comp_unit_data1_out(0), A0=>nx16967, A1=>
      nx15538, B0=>nx15541);
   bias1_reg_reg_q_0 : dffr port map ( Q=>OPEN, QB=>nx15538, D=>nx13387, CLK
      =>clk, R=>reset);
   ix15542 : nand02 port map ( Y=>nx15541, A0=>nx1960, A1=>nx16913);
   ix2005 : oai21 port map ( Y=>comp_unit_data1_out(1), A0=>nx16967, A1=>
      nx15547, B0=>nx15550);
   bias1_reg_reg_q_1 : dffr port map ( Q=>OPEN, QB=>nx15547, D=>nx13407, CLK
      =>clk, R=>reset);
   ix15551 : nand02 port map ( Y=>nx15550, A0=>nx1994, A1=>nx16913);
   ix2031 : oai21 port map ( Y=>comp_unit_data1_out(2), A0=>nx16967, A1=>
      nx15553, B0=>nx15556);
   bias1_reg_reg_q_2 : dffr port map ( Q=>OPEN, QB=>nx15553, D=>nx13427, CLK
      =>clk, R=>reset);
   ix15557 : nand02 port map ( Y=>nx15556, A0=>nx2020, A1=>nx16913);
   ix2057 : oai21 port map ( Y=>comp_unit_data1_out(3), A0=>nx16969, A1=>
      nx15559, B0=>nx15562);
   bias1_reg_reg_q_3 : dffr port map ( Q=>OPEN, QB=>nx15559, D=>nx13447, CLK
      =>clk, R=>reset);
   ix15563 : nand02 port map ( Y=>nx15562, A0=>nx2046, A1=>nx16913);
   ix2083 : oai21 port map ( Y=>comp_unit_data1_out(4), A0=>nx16969, A1=>
      nx15565, B0=>nx15568);
   bias1_reg_reg_q_4 : dffr port map ( Q=>OPEN, QB=>nx15565, D=>nx13467, CLK
      =>clk, R=>reset);
   ix15569 : nand02 port map ( Y=>nx15568, A0=>nx2072, A1=>nx16913);
   ix2109 : oai21 port map ( Y=>comp_unit_data1_out(5), A0=>nx16969, A1=>
      nx15571, B0=>nx15574);
   bias1_reg_reg_q_5 : dffr port map ( Q=>OPEN, QB=>nx15571, D=>nx13487, CLK
      =>clk, R=>reset);
   ix15575 : nand02 port map ( Y=>nx15574, A0=>nx2098, A1=>nx16913);
   ix2135 : oai21 port map ( Y=>comp_unit_data1_out(6), A0=>nx16969, A1=>
      nx15577, B0=>nx15580);
   bias1_reg_reg_q_6 : dffr port map ( Q=>OPEN, QB=>nx15577, D=>nx13507, CLK
      =>clk, R=>reset);
   ix15581 : nand02 port map ( Y=>nx15580, A0=>nx2124, A1=>nx16913);
   ix2161 : oai21 port map ( Y=>comp_unit_data1_out(7), A0=>nx16969, A1=>
      nx15583, B0=>nx15586);
   bias1_reg_reg_q_7 : dffr port map ( Q=>OPEN, QB=>nx15583, D=>nx13527, CLK
      =>clk, R=>reset);
   ix15587 : nand02 port map ( Y=>nx15586, A0=>nx2150, A1=>nx16915);
   ix2187 : oai21 port map ( Y=>comp_unit_data1_out(8), A0=>nx16969, A1=>
      nx15589, B0=>nx15592);
   bias1_reg_reg_q_8 : dffr port map ( Q=>OPEN, QB=>nx15589, D=>nx13547, CLK
      =>clk, R=>reset);
   ix15593 : nand02 port map ( Y=>nx15592, A0=>nx2176, A1=>nx16915);
   ix2213 : oai21 port map ( Y=>comp_unit_data1_out(9), A0=>nx16969, A1=>
      nx15595, B0=>nx15598);
   bias1_reg_reg_q_9 : dffr port map ( Q=>OPEN, QB=>nx15595, D=>nx13567, CLK
      =>clk, R=>reset);
   ix15599 : nand02 port map ( Y=>nx15598, A0=>nx2202, A1=>nx16915);
   ix2239 : oai21 port map ( Y=>comp_unit_data1_out(10), A0=>nx16971, A1=>
      nx15601, B0=>nx15604);
   bias1_reg_reg_q_10 : dffr port map ( Q=>OPEN, QB=>nx15601, D=>nx13587, 
      CLK=>clk, R=>reset);
   ix15605 : nand02 port map ( Y=>nx15604, A0=>nx2228, A1=>nx16915);
   ix2265 : oai21 port map ( Y=>comp_unit_data1_out(11), A0=>nx16971, A1=>
      nx15607, B0=>nx15610);
   bias1_reg_reg_q_11 : dffr port map ( Q=>OPEN, QB=>nx15607, D=>nx13607, 
      CLK=>clk, R=>reset);
   ix15611 : nand02 port map ( Y=>nx15610, A0=>nx2254, A1=>nx16915);
   ix2291 : oai21 port map ( Y=>comp_unit_data1_out(12), A0=>nx16971, A1=>
      nx15613, B0=>nx15616);
   bias1_reg_reg_q_12 : dffr port map ( Q=>OPEN, QB=>nx15613, D=>nx13627, 
      CLK=>clk, R=>reset);
   ix15617 : nand02 port map ( Y=>nx15616, A0=>nx2280, A1=>nx16915);
   ix2317 : oai21 port map ( Y=>comp_unit_data1_out(13), A0=>nx16971, A1=>
      nx15619, B0=>nx15622);
   bias1_reg_reg_q_13 : dffr port map ( Q=>OPEN, QB=>nx15619, D=>nx13647, 
      CLK=>clk, R=>reset);
   ix15623 : nand02 port map ( Y=>nx15622, A0=>nx2306, A1=>nx16915);
   ix2343 : oai21 port map ( Y=>comp_unit_data1_out(14), A0=>nx16971, A1=>
      nx15625, B0=>nx15628);
   bias1_reg_reg_q_14 : dffr port map ( Q=>OPEN, QB=>nx15625, D=>nx13667, 
      CLK=>clk, R=>reset);
   ix15629 : nand02 port map ( Y=>nx15628, A0=>nx2332, A1=>nx16917);
   ix2369 : oai21 port map ( Y=>comp_unit_data1_out(15), A0=>nx16971, A1=>
      nx15631, B0=>nx15634);
   bias1_reg_reg_q_15 : dffr port map ( Q=>OPEN, QB=>nx15631, D=>nx13687, 
      CLK=>clk, R=>reset);
   ix15635 : nand02 port map ( Y=>nx15634, A0=>nx2358, A1=>nx16917);
   ix1933 : oai21 port map ( Y=>comp_unit_ready, A0=>nx17129, A1=>nx646, B0
      =>nx15637);
   ix15638 : aoi21 port map ( Y=>nx15637, A0=>nx16891, A1=>nx15077, B0=>
      nx17075);
   ix2381 : nand03 port map ( Y=>wind_en, A0=>nx17071, A1=>nx17217, A2=>
      nx15739);
   ix4509 : aoi21 port map ( Y=>mem_read_out, A0=>nx15742, A1=>nx15750, B0=>
      reset);
   ix15748 : oai21 port map ( Y=>nx15747, A0=>comp_unit_operation_EXMPLR, A1
      =>nx15293, B0=>nx1966);
   ix2569 : nand02 port map ( Y=>nx2568, A0=>nx15753, A1=>nx15755);
   ix15754 : nor04 port map ( Y=>nx15753, A0=>current_state_1, A1=>
      current_state_2, A2=>nx16839, A3=>current_state_4);
   ix4493 : aoi21 port map ( Y=>mem_write_out, A0=>nx14717, A1=>nx15758, B0
      =>reset);
   reg_current_state_26 : dffr port map ( Q=>OPEN, QB=>nx15758, D=>nx1762, 
      CLK=>nx16781, R=>reset);
   ix2615 : nand02 port map ( Y=>mem_addr_out(0), A0=>nx15762, A1=>nx15811);
   ix15763 : aoi21 port map ( Y=>nx15762, A0=>addr1_data_0, A1=>nx17089, B0
      =>nx2610);
   reg_addr1_data_0 : dffr port map ( Q=>addr1_data_0, QB=>OPEN, D=>nx13737, 
      CLK=>clk, R=>reset);
   ix2611 : oai22 port map ( Y=>nx2610, A0=>nx17805, A1=>nx15793, B0=>
      img_addr_offset_0, B1=>nx16977);
   ix13718 : mux21_ni port map ( Y=>nx13717, A0=>nx2502, A1=>nx16919, S0=>
      nx15791);
   ix2503 : oai33 port map ( Y=>nx2502, A0=>nx15781, A1=>nx2478, A2=>nx16947, 
      B0=>nx15785, B1=>nx16941, B2=>nx2494);
   reg_write_base_reg_q_0 : dffr port map ( Q=>OPEN, QB=>nx15777, D=>nx13717, 
      CLK=>clk, R=>reset);
   layer_mem_size_reg_q_0 : dffr port map ( Q=>layer_mem_size_out_0, QB=>
      OPEN, D=>nx13707, CLK=>clk, R=>reset);
   ix15794 : aoi222 port map ( Y=>nx15793, A0=>nx15795, A1=>nx2532, B0=>
      nx15800, B1=>nx16935, C0=>nx18293, C1=>nx2472);
   ix15796 : nand02 port map ( Y=>nx15795, A0=>bias_offset_data_out_0, A1=>
      nx16919);
   reg_bias_offset_reg_q_0 : dffr port map ( Q=>bias_offset_data_out_0, QB=>
      OPEN, D=>nx13727, CLK=>clk, R=>reset);
   ix2521 : nand02 port map ( Y=>nx2520, A0=>nx17163, A1=>nx14717);
   reg_img_addr_offset_0 : dffr port map ( Q=>img_addr_offset_0, QB=>OPEN, D
      =>nx13747, CLK=>clk, R=>reset);
   ix15812 : aoi332 port map ( Y=>nx15811, A0=>nx2532, A1=>
      bias_offset_data_out_0, A2=>nx17805, B0=>nx2472, B1=>
      class_cntr_counter_out_0, B2=>nx18293, C0=>nx16935, C1=>nx2526);
   ix2701 : oai221 port map ( Y=>mem_addr_out(1), A0=>nx15815, A1=>nx17009, 
      B0=>nx15823, B1=>nx17019, C0=>nx15849);
   ix15819 : oai21 port map ( Y=>nx15818, A0=>addr1_data_0, A1=>addr1_data_1, 
      B0=>nx15821);
   reg_addr1_data_1 : dffr port map ( Q=>addr1_data_1, QB=>nx15815, D=>
      nx13797, CLK=>clk, R=>reset);
   ix15822 : nand02 port map ( Y=>nx15821, A0=>addr1_data_1, A1=>
      addr1_data_0);
   ix15824 : xnor2 port map ( Y=>nx15823, A0=>nx18293, A1=>nx15825);
   ix13778 : oai222 port map ( Y=>nx13777, A0=>nx17811, A1=>nx16923, B0=>
      nx15832, B1=>nx16947, C0=>nx16941, C1=>nx15838);
   reg_write_base_reg_q_1 : dffr port map ( Q=>write_base_data_out_1, QB=>
      nx15829, D=>nx13777, CLK=>clk, R=>reset);
   ix15833 : xnor2 port map ( Y=>nx15832, A0=>nx15834, A1=>nx15836);
   ix15835 : nand02 port map ( Y=>nx15834, A0=>new_size_squared_out_0, A1=>
      nx16919);
   ix15839 : xnor2 port map ( Y=>nx15838, A0=>nx15840, A1=>nx15842);
   ix15841 : nand02 port map ( Y=>nx15840, A0=>layer_mem_size_out_0, A1=>
      nx16919);
   layer_mem_size_reg_q_1 : dffr port map ( Q=>layer_mem_size_out_1, QB=>
      OPEN, D=>nx13767, CLK=>clk, R=>reset);
   ix15850 : aoi222 port map ( Y=>nx15849, A0=>nx15851, A1=>nx17237, B0=>
      nx2670, B1=>nx2532, C0=>nx2658, C1=>nx16935);
   ix15852 : oai21 port map ( Y=>nx15851, A0=>img_addr_offset_0, A1=>
      img_addr_offset_1, B0=>nx15857);
   reg_img_addr_offset_1 : dffr port map ( Q=>img_addr_offset_1, QB=>nx15855, 
      D=>nx13757, CLK=>clk, R=>reset);
   ix15858 : nand02 port map ( Y=>nx15857, A0=>img_addr_offset_1, A1=>
      img_addr_offset_0);
   ix2671 : xor2 port map ( Y=>nx2670, A0=>nx15795, A1=>nx15860);
   reg_bias_offset_reg_q_1 : dffr port map ( Q=>bias_offset_data_out_1, QB=>
      nx15864, D=>nx13787, CLK=>clk, R=>reset);
   ix2659 : xor2 port map ( Y=>nx2658, A0=>nx15800, A1=>nx15867);
   ix2833 : oai221 port map ( Y=>mem_addr_out(2), A0=>nx15870, A1=>nx17009, 
      B0=>nx15875, B1=>nx17019, C0=>nx15901);
   reg_addr1_data_2 : dffr port map ( Q=>addr1_data_2, QB=>nx15870, D=>
      nx13847, CLK=>clk, R=>reset);
   ix15876 : xor2 port map ( Y=>nx15875, A0=>nx2808, A1=>nx15878);
   ix13828 : oai222 port map ( Y=>nx13827, A0=>nx17169, A1=>nx16923, B0=>
      nx15884, B1=>nx16947, C0=>nx16941, C1=>nx15891);
   reg_write_base_reg_q_2 : dffr port map ( Q=>write_base_data_out_2, QB=>
      OPEN, D=>nx13827, CLK=>clk, R=>reset);
   ix15885 : xnor2 port map ( Y=>nx15884, A0=>nx15886, A1=>nx15889);
   ix15892 : xnor2 port map ( Y=>nx15891, A0=>nx15893, A1=>nx15896);
   layer_mem_size_reg_q_2 : dffr port map ( Q=>layer_mem_size_out_2, QB=>
      nx15900, D=>nx13817, CLK=>clk, R=>reset);
   ix15902 : aoi222 port map ( Y=>nx15901, A0=>nx2794, A1=>nx16935, B0=>
      nx17237, B1=>nx2780, C0=>nx2758, C1=>nx2532);
   ix2795 : xnor2 port map ( Y=>nx2794, A0=>nx2790, A1=>nx15905);
   ix2781 : oai21 port map ( Y=>nx2780, A0=>nx15908, A1=>nx15913, B0=>nx2774
   );
   reg_img_addr_offset_2 : dffr port map ( Q=>img_addr_offset_2, QB=>nx15908, 
      D=>nx13837, CLK=>clk, R=>reset);
   ix2759 : xor2 port map ( Y=>nx2758, A0=>nx15917, A1=>nx15920);
   reg_bias_offset_reg_q_2 : dffr port map ( Q=>OPEN, QB=>nx15924, D=>
      nx13807, CLK=>clk, R=>reset);
   ix2965 : oai221 port map ( Y=>mem_addr_out(3), A0=>nx15927, A1=>nx17009, 
      B0=>nx15934, B1=>nx17019, C0=>nx15958);
   reg_addr1_data_3 : dffr port map ( Q=>addr1_data_3, QB=>nx15927, D=>
      nx13897, CLK=>clk, R=>reset);
   ix15933 : nand03 port map ( Y=>nx15932, A0=>addr1_data_2, A1=>
      addr1_data_1, A2=>addr1_data_0);
   ix15935 : xnor2 port map ( Y=>nx15934, A0=>nx15936, A1=>nx15939);
   ix13878 : oai222 port map ( Y=>nx13877, A0=>nx15943, A1=>nx16947, B0=>
      nx16941, B1=>nx15948, C0=>nx17816, C1=>nx16923);
   ix15944 : xor2 port map ( Y=>nx15943, A0=>nx2854, A1=>nx15946);
   ix15949 : xor2 port map ( Y=>nx15948, A0=>nx2868, A1=>nx15951);
   layer_mem_size_reg_q_3 : dffr port map ( Q=>layer_mem_size_out_3, QB=>
      OPEN, D=>nx13867, CLK=>clk, R=>reset);
   reg_write_base_reg_q_3 : dffs_ni port map ( Q=>write_base_data_out_3, QB
      =>nx15956, D=>nx13877, CLK=>clk, S=>reset);
   ix15959 : aoi332 port map ( Y=>nx15958, A0=>nx2906, A1=>nx15970, A2=>
      nx17237, B0=>nx2890, B1=>nx17075, B2=>nx17149, C0=>nx2926, C1=>nx16935
   );
   ix2907 : nand02 port map ( Y=>nx2906, A0=>nx15961, A1=>nx15963);
   ix15962 : nor03_2x port map ( Y=>nx15961, A0=>img_addr_offset_0, A1=>
      img_addr_offset_1, A2=>img_addr_offset_2);
   reg_img_addr_offset_3 : dffr port map ( Q=>img_addr_offset_3, QB=>nx15963, 
      D=>nx13887, CLK=>clk, R=>reset);
   ix15969 : nand03 port map ( Y=>nx15968, A0=>img_addr_offset_2, A1=>
      img_addr_offset_1, A2=>img_addr_offset_0);
   ix2891 : xnor2 port map ( Y=>nx2890, A0=>nx17522, A1=>nx18295);
   reg_bias_offset_reg_q_3 : dffr port map ( Q=>bias_offset_data_out_3, QB=>
      OPEN, D=>nx13857, CLK=>clk, R=>reset);
   ix2927 : xor2 port map ( Y=>nx2926, A0=>nx15981, A1=>nx15984);
   ix3101 : oai221 port map ( Y=>mem_addr_out(4), A0=>nx15987, A1=>nx17011, 
      B0=>nx15995, B1=>nx17023, C0=>nx16029);
   ix3091 : aoi21 port map ( Y=>nx3090, A0=>nx15991, A1=>nx15987, B0=>nx3084
   );
   ix15992 : nand04 port map ( Y=>nx15991, A0=>addr1_data_3, A1=>
      addr1_data_2, A2=>addr1_data_1, A3=>addr1_data_0);
   reg_addr1_data_4 : dffr port map ( Q=>addr1_data_4, QB=>nx15987, D=>
      nx13947, CLK=>clk, R=>reset);
   ix15996 : xnor2 port map ( Y=>nx15995, A0=>nx15997, A1=>nx16000);
   reg_bias_offset_reg_q_4 : dffr port map ( Q=>bias_offset_data_out_4, QB=>
      nx16005, D=>nx13937, CLK=>clk, R=>reset);
   ix105 : aoi21 port map ( Y=>nx104, A0=>nx14747, A1=>nx14741, B0=>nx98);
   ix13918 : oai222 port map ( Y=>nx13917, A0=>nx17173, A1=>nx16923, B0=>
      nx16010, B1=>nx16949, C0=>nx16941, C1=>nx16017);
   reg_write_base_reg_q_4 : dffr port map ( Q=>write_base_data_out_4, QB=>
      OPEN, D=>nx13917, CLK=>clk, R=>reset);
   ix16011 : xnor2 port map ( Y=>nx16010, A0=>nx16012, A1=>nx16015);
   ix16018 : xnor2 port map ( Y=>nx16017, A0=>nx16019, A1=>nx16022);
   layer_mem_size_reg_q_4 : dffr port map ( Q=>layer_mem_size_out_4, QB=>
      nx16026, D=>nx13907, CLK=>clk, R=>reset);
   ix16028 : nand02 port map ( Y=>nx16027, A0=>nx17075, A1=>nx17149);
   ix16030 : aoi21 port map ( Y=>nx16029, A0=>nx3016, A1=>nx16935, B0=>
      nx3060);
   ix3017 : xnor2 port map ( Y=>nx3016, A0=>nx2972, A1=>nx16033);
   ix3061 : oai32 port map ( Y=>nx3060, A0=>nx16036, A1=>nx16099, A2=>
      nx17019, B0=>nx16979, B1=>nx16040);
   ix16041 : aoi21 port map ( Y=>nx16040, A0=>img_addr_offset_4, A1=>nx2908, 
      B0=>nx16051);
   ix3045 : aoi21 port map ( Y=>nx3044, A0=>nx16045, A1=>nx16047, B0=>nx3038
   );
   ix16046 : nand04 port map ( Y=>nx16045, A0=>img_addr_offset_3, A1=>
      img_addr_offset_2, A2=>img_addr_offset_1, A3=>img_addr_offset_0);
   reg_img_addr_offset_4 : dffr port map ( Q=>img_addr_offset_4, QB=>nx16047, 
      D=>nx13927, CLK=>clk, R=>reset);
   ix3229 : oai221 port map ( Y=>mem_addr_out(5), A0=>nx16054, A1=>nx17023, 
      B0=>nx16080, B1=>nx17011, C0=>nx16088);
   ix16055 : xor2 port map ( Y=>nx16054, A0=>nx3198, A1=>nx16057);
   reg_bias_offset_reg_q_5 : dffr port map ( Q=>bias_offset_data_out_5, QB=>
      nx16061, D=>nx13987, CLK=>clk, R=>reset);
   ix13968 : oai222 port map ( Y=>nx13967, A0=>nx16065, A1=>nx16949, B0=>
      nx16943, B1=>nx16070, C0=>nx17820, C1=>nx16923);
   ix16066 : xor2 port map ( Y=>nx16065, A0=>nx3116, A1=>nx16068);
   ix16071 : xor2 port map ( Y=>nx16070, A0=>nx3130, A1=>nx16073);
   layer_mem_size_reg_q_5 : dffr port map ( Q=>layer_mem_size_out_5, QB=>
      OPEN, D=>nx13957, CLK=>clk, R=>reset);
   reg_write_base_reg_q_5 : dffs_ni port map ( Q=>write_base_data_out_5, QB
      =>nx16078, D=>nx13967, CLK=>clk, S=>reset);
   ix16084 : oai21 port map ( Y=>nx16083, A0=>nx3084, A1=>addr1_data_5, B0=>
      nx16086);
   reg_addr1_data_5 : dffr port map ( Q=>addr1_data_5, QB=>nx16080, D=>
      nx13997, CLK=>clk, R=>reset);
   ix16087 : nand02 port map ( Y=>nx16086, A0=>addr1_data_5, A1=>nx3084);
   ix16089 : aoi21 port map ( Y=>nx16088, A0=>nx3152, A1=>nx16935, B0=>
      nx3188);
   ix3153 : xor2 port map ( Y=>nx3152, A0=>nx16091, A1=>nx16094);
   ix3189 : oai33 port map ( Y=>nx3188, A0=>nx16097, A1=>nx3180, A2=>nx17019, 
      B0=>nx16102, B1=>nx3170, B2=>nx16979);
   ix16107 : oai21 port map ( Y=>nx16106, A0=>nx3038, A1=>img_addr_offset_5, 
      B0=>nx16108);
   ix16109 : nand02 port map ( Y=>nx16108, A0=>img_addr_offset_5, A1=>nx3038
   );
   reg_img_addr_offset_5 : dffr port map ( Q=>img_addr_offset_5, QB=>nx16110, 
      D=>nx13977, CLK=>clk, R=>reset);
   ix3357 : oai221 port map ( Y=>mem_addr_out(6), A0=>nx16114, A1=>nx17023, 
      B0=>nx16146, B1=>nx17011, C0=>nx16151);
   ix16115 : xnor2 port map ( Y=>nx16114, A0=>nx16116, A1=>nx16119);
   reg_bias_offset_reg_q_6 : dffr port map ( Q=>bias_offset_data_out_6, QB=>
      nx16124, D=>nx14037, CLK=>clk, R=>reset);
   ix151 : aoi21 port map ( Y=>nx150, A0=>nx14732, A1=>nx14726, B0=>nx144);
   ix14018 : oai222 port map ( Y=>nx14017, A0=>nx16127, A1=>nx16949, B0=>
      nx16943, B1=>nx16134, C0=>nx17177, C1=>nx16923);
   ix16128 : xnor2 port map ( Y=>nx16127, A0=>nx16129, A1=>nx16132);
   ix16135 : xnor2 port map ( Y=>nx16134, A0=>nx16136, A1=>nx16139);
   layer_mem_size_reg_q_6 : dffr port map ( Q=>layer_mem_size_out_6, QB=>
      nx16143, D=>nx14007, CLK=>clk, R=>reset);
   reg_write_base_reg_q_6 : dffs_ni port map ( Q=>write_base_data_out_6, QB
      =>OPEN, D=>nx14017, CLK=>clk, S=>reset);
   reg_addr1_data_6 : dffr port map ( Q=>addr1_data_6, QB=>nx16146, D=>
      nx14047, CLK=>clk, R=>reset);
   ix16152 : aoi21 port map ( Y=>nx16151, A0=>nx3280, A1=>nx16937, B0=>
      nx3316);
   ix3281 : xnor2 port map ( Y=>nx3280, A0=>nx3236, A1=>nx16155);
   ix3317 : oai32 port map ( Y=>nx3316, A0=>nx16158, A1=>nx3286, A2=>nx17019, 
      B0=>nx16979, B1=>nx16161);
   ix16162 : aoi21 port map ( Y=>nx16161, A0=>img_addr_offset_6, A1=>nx3170, 
      B0=>nx16169);
   ix3301 : aoi21 port map ( Y=>nx3300, A0=>nx16108, A1=>nx16166, B0=>nx3294
   );
   reg_img_addr_offset_6 : dffr port map ( Q=>img_addr_offset_6, QB=>nx16166, 
      D=>nx14027, CLK=>clk, R=>reset);
   ix3485 : oai221 port map ( Y=>mem_addr_out(7), A0=>nx16172, A1=>nx17023, 
      B0=>nx16198, B1=>nx17013, C0=>nx16207);
   ix16173 : xor2 port map ( Y=>nx16172, A0=>nx3454, A1=>nx16175);
   reg_bias_offset_reg_q_7 : dffr port map ( Q=>bias_offset_data_out_7, QB=>
      nx16179, D=>nx14087, CLK=>clk, R=>reset);
   ix14068 : oai222 port map ( Y=>nx14067, A0=>nx16183, A1=>nx16949, B0=>
      nx16943, B1=>nx16188, C0=>nx16196, C1=>nx16923);
   ix16184 : xor2 port map ( Y=>nx16183, A0=>nx3372, A1=>nx16186);
   ix16189 : xor2 port map ( Y=>nx16188, A0=>nx17753, A1=>nx16191);
   layer_mem_size_reg_q_7 : dffr port map ( Q=>layer_mem_size_out_7, QB=>
      OPEN, D=>nx14057, CLK=>clk, R=>reset);
   reg_write_base_reg_q_7 : dffr port map ( Q=>write_base_data_out_7, QB=>
      nx16196, D=>nx14067, CLK=>clk, R=>reset);
   ix16202 : oai21 port map ( Y=>nx16201, A0=>nx3340, A1=>addr1_data_7, B0=>
      nx16205);
   reg_addr1_data_7 : dffr port map ( Q=>addr1_data_7, QB=>nx16198, D=>
      nx14097, CLK=>clk, R=>reset);
   ix16206 : nand02 port map ( Y=>nx16205, A0=>addr1_data_7, A1=>nx3340);
   ix16208 : aoi21 port map ( Y=>nx16207, A0=>nx3408, A1=>nx16937, B0=>
      nx3444);
   ix3409 : xor2 port map ( Y=>nx3408, A0=>nx16210, A1=>nx16213);
   ix3445 : oai33 port map ( Y=>nx3444, A0=>nx16216, A1=>nx3436, A2=>nx17019, 
      B0=>nx16221, B1=>nx3426, B2=>nx16981);
   ix16226 : oai21 port map ( Y=>nx16225, A0=>nx3294, A1=>img_addr_offset_7, 
      B0=>nx16227);
   ix16228 : nand02 port map ( Y=>nx16227, A0=>img_addr_offset_7, A1=>nx3294
   );
   reg_img_addr_offset_7 : dffr port map ( Q=>img_addr_offset_7, QB=>nx16229, 
      D=>nx14077, CLK=>clk, R=>reset);
   ix3613 : oai221 port map ( Y=>mem_addr_out(8), A0=>nx16233, A1=>nx17023, 
      B0=>nx16265, B1=>nx17013, C0=>nx16270);
   ix16234 : xnor2 port map ( Y=>nx16233, A0=>nx16235, A1=>nx16238);
   reg_bias_offset_reg_q_8 : dffr port map ( Q=>bias_offset_data_out_8, QB=>
      nx16243, D=>nx14137, CLK=>clk, R=>reset);
   ix201 : aoi21 port map ( Y=>nx200, A0=>nx14708, A1=>nx14702, B0=>nx194);
   ix14118 : oai222 port map ( Y=>nx14117, A0=>nx16246, A1=>nx16949, B0=>
      nx16943, B1=>nx16253, C0=>nx17181, C1=>nx16925);
   ix16247 : xnor2 port map ( Y=>nx16246, A0=>nx16248, A1=>nx16251);
   ix16254 : xnor2 port map ( Y=>nx16253, A0=>nx16255, A1=>nx16258);
   layer_mem_size_reg_q_8 : dffr port map ( Q=>layer_mem_size_out_8, QB=>
      nx16262, D=>nx14107, CLK=>clk, R=>reset);
   reg_write_base_reg_q_8 : dffs_ni port map ( Q=>write_base_data_out_8, QB
      =>OPEN, D=>nx14117, CLK=>clk, S=>reset);
   reg_addr1_data_8 : dffr port map ( Q=>addr1_data_8, QB=>nx16265, D=>
      nx14147, CLK=>clk, R=>reset);
   ix16271 : aoi21 port map ( Y=>nx16270, A0=>nx3536, A1=>nx16937, B0=>
      nx3572);
   ix3537 : xnor2 port map ( Y=>nx3536, A0=>nx3492, A1=>nx16274);
   ix3493 : oai22 port map ( Y=>nx3492, A0=>nx17680, A1=>nx16213, B0=>
      nx14712, B1=>nx16196);
   ix3573 : oai33 port map ( Y=>nx3572, A0=>nx16277, A1=>nx3564, A2=>nx17826, 
      B0=>nx16280, B1=>nx3554, B2=>nx16981);
   ix3547 : aoi21 port map ( Y=>nx3546, A0=>nx16227, A1=>nx16285, B0=>nx3540
   );
   reg_img_addr_offset_8 : dffr port map ( Q=>img_addr_offset_8, QB=>nx16285, 
      D=>nx14127, CLK=>clk, R=>reset);
   ix3741 : oai221 port map ( Y=>mem_addr_out(9), A0=>nx16290, A1=>nx17023, 
      B0=>nx16316, B1=>nx17013, C0=>nx16325);
   ix16291 : xor2 port map ( Y=>nx16290, A0=>nx3710, A1=>nx16293);
   reg_bias_offset_reg_q_9 : dffr port map ( Q=>bias_offset_data_out_9, QB=>
      nx16297, D=>nx14187, CLK=>clk, R=>reset);
   ix14168 : oai222 port map ( Y=>nx14167, A0=>nx16301, A1=>nx16949, B0=>
      nx16943, B1=>nx16306, C0=>nx16314, C1=>nx16925);
   ix16302 : xor2 port map ( Y=>nx16301, A0=>nx17739, A1=>nx16304);
   ix16307 : xor2 port map ( Y=>nx16306, A0=>nx3642, A1=>nx16309);
   layer_mem_size_reg_q_9 : dffr port map ( Q=>layer_mem_size_out_9, QB=>
      OPEN, D=>nx14157, CLK=>clk, R=>reset);
   reg_write_base_reg_q_9 : dffs_ni port map ( Q=>write_base_data_out_9, QB
      =>nx16314, D=>nx14167, CLK=>clk, S=>reset);
   ix16320 : oai21 port map ( Y=>nx16319, A0=>nx3596, A1=>addr1_data_9, B0=>
      nx16323);
   reg_addr1_data_9 : dffr port map ( Q=>addr1_data_9, QB=>nx16316, D=>
      nx14197, CLK=>clk, R=>reset);
   ix16324 : nand02 port map ( Y=>nx16323, A0=>addr1_data_9, A1=>nx3596);
   ix16326 : aoi21 port map ( Y=>nx16325, A0=>nx3664, A1=>nx16937, B0=>
      nx3700);
   ix3665 : xor2 port map ( Y=>nx3664, A0=>nx16328, A1=>nx16331);
   ix16329 : aoi22 port map ( Y=>nx16328, A0=>write_offset_data_out_8, A1=>
      nx17824, B0=>nx3492, B1=>nx3534);
   ix3701 : oai33 port map ( Y=>nx3700, A0=>nx16334, A1=>nx17828, A2=>
      nx17826, B0=>nx16339, B1=>nx3682, B2=>nx16981);
   ix16344 : oai21 port map ( Y=>nx16343, A0=>nx3540, A1=>img_addr_offset_9, 
      B0=>nx16345);
   ix16346 : nand02 port map ( Y=>nx16345, A0=>img_addr_offset_9, A1=>nx3540
   );
   reg_img_addr_offset_9 : dffr port map ( Q=>img_addr_offset_9, QB=>nx16347, 
      D=>nx14177, CLK=>clk, R=>reset);
   ix16350 : nand02 port map ( Y=>nx16349, A0=>img_addr_offset_8, A1=>nx3426
   );
   ix3869 : oai221 port map ( Y=>mem_addr_out(10), A0=>nx16353, A1=>nx17023, 
      B0=>nx16385, B1=>nx17013, C0=>nx16390);
   ix16354 : xnor2 port map ( Y=>nx16353, A0=>nx16355, A1=>nx16358);
   reg_bias_offset_reg_q_10 : dffr port map ( Q=>bias_offset_data_out_10, QB
      =>nx16363, D=>nx14237, CLK=>clk, R=>reset);
   ix247 : aoi21 port map ( Y=>nx246, A0=>nx14695, A1=>nx14689, B0=>nx240);
   ix14218 : oai222 port map ( Y=>nx14217, A0=>nx16366, A1=>nx16949, B0=>
      nx16943, B1=>nx16373, C0=>nx17185, C1=>nx16925);
   ix16367 : xnor2 port map ( Y=>nx16366, A0=>nx16368, A1=>nx16371);
   ix16374 : xnor2 port map ( Y=>nx16373, A0=>nx16375, A1=>nx16378);
   layer_mem_size_reg_q_10 : dffr port map ( Q=>layer_mem_size_out_10, QB=>
      nx16382, D=>nx14207, CLK=>clk, R=>reset);
   reg_write_base_reg_q_10 : dffr port map ( Q=>write_base_data_out_10, QB=>
      OPEN, D=>nx14217, CLK=>clk, R=>reset);
   reg_addr1_data_10 : dffr port map ( Q=>addr1_data_10, QB=>nx16385, D=>
      nx14247, CLK=>clk, R=>reset);
   ix16391 : aoi21 port map ( Y=>nx16390, A0=>nx3792, A1=>nx16937, B0=>
      nx3828);
   ix3793 : xnor2 port map ( Y=>nx3792, A0=>nx3748, A1=>nx16394);
   ix3749 : oai22 port map ( Y=>nx3748, A0=>nx16328, A1=>nx16331, B0=>
      nx14776, B1=>nx16314);
   ix3829 : oai33 port map ( Y=>nx3828, A0=>nx16397, A1=>nx3820, A2=>nx17826, 
      B0=>nx16400, B1=>nx3810, B2=>nx16981);
   ix3803 : aoi21 port map ( Y=>nx3802, A0=>nx16345, A1=>nx16405, B0=>nx3796
   );
   reg_img_addr_offset_10 : dffr port map ( Q=>img_addr_offset_10, QB=>
      nx16405, D=>nx14227, CLK=>clk, R=>reset);
   ix3997 : oai221 port map ( Y=>mem_addr_out(11), A0=>nx16410, A1=>nx17025, 
      B0=>nx16436, B1=>nx17015, C0=>nx16445);
   ix16411 : xor2 port map ( Y=>nx16410, A0=>nx3966, A1=>nx16413);
   reg_bias_offset_reg_q_11 : dffr port map ( Q=>bias_offset_data_out_11, QB
      =>nx16417, D=>nx14287, CLK=>clk, R=>reset);
   layer_mem_size_reg_q_11 : dffr port map ( Q=>layer_mem_size_out_11, QB=>
      OPEN, D=>nx14257, CLK=>clk, R=>reset);
   reg_write_base_reg_q_11 : dffs_ni port map ( Q=>write_base_data_out_11, 
      QB=>nx16434, D=>nx14267, CLK=>clk, S=>reset);
   ix16440 : oai21 port map ( Y=>nx16439, A0=>nx3852, A1=>addr1_data_11, B0
      =>nx16443);
   reg_addr1_data_11 : dffr port map ( Q=>addr1_data_11, QB=>nx16436, D=>
      nx14297, CLK=>clk, R=>reset);
   ix16444 : nand02 port map ( Y=>nx16443, A0=>addr1_data_11, A1=>nx3852);
   ix16446 : aoi21 port map ( Y=>nx16445, A0=>nx3920, A1=>nx16937, B0=>
      nx3956);
   ix3921 : xor2 port map ( Y=>nx3920, A0=>nx16448, A1=>nx16451);
   ix3957 : oai32 port map ( Y=>nx3956, A0=>nx16454, A1=>nx3926, A2=>nx17826, 
      B0=>nx16983, B1=>nx16459);
   ix16464 : oai21 port map ( Y=>nx16463, A0=>nx3796, A1=>img_addr_offset_11, 
      B0=>nx16465);
   ix16466 : nand02 port map ( Y=>nx16465, A0=>img_addr_offset_11, A1=>
      nx3796);
   reg_img_addr_offset_11 : dffr port map ( Q=>img_addr_offset_11, QB=>
      nx16467, D=>nx14277, CLK=>clk, R=>reset);
   ix16470 : nand02 port map ( Y=>nx16469, A0=>img_addr_offset_10, A1=>
      nx3682);
   ix4125 : oai221 port map ( Y=>mem_addr_out(12), A0=>nx16472, A1=>nx17025, 
      B0=>nx16504, B1=>nx17015, C0=>nx16509);
   ix16473 : xnor2 port map ( Y=>nx16472, A0=>nx16474, A1=>nx16477);
   reg_bias_offset_reg_q_12 : dffr port map ( Q=>bias_offset_data_out_12, QB
      =>nx16482, D=>nx14337, CLK=>clk, R=>reset);
   ix295 : aoi21 port map ( Y=>nx294, A0=>nx14682, A1=>nx14676, B0=>nx288);
   ix14318 : oai222 port map ( Y=>nx14317, A0=>nx16485, A1=>nx16951, B0=>
      nx17215, B1=>nx16492, C0=>nx17189, C1=>nx16925);
   ix16486 : xnor2 port map ( Y=>nx16485, A0=>nx18303, A1=>nx16490);
   ix16493 : xnor2 port map ( Y=>nx16492, A0=>nx16494, A1=>nx16497);
   layer_mem_size_reg_q_12 : dffr port map ( Q=>layer_mem_size_out_12, QB=>
      nx16501, D=>nx14307, CLK=>clk, R=>reset);
   reg_write_base_reg_q_12 : dffs_ni port map ( Q=>write_base_data_out_12, 
      QB=>OPEN, D=>nx14317, CLK=>clk, S=>reset);
   reg_addr1_data_12 : dffr port map ( Q=>addr1_data_12, QB=>nx16504, D=>
      nx14347, CLK=>clk, R=>reset);
   ix16510 : aoi21 port map ( Y=>nx16509, A0=>nx4048, A1=>nx16937, B0=>
      nx4084);
   ix4049 : xnor2 port map ( Y=>nx4048, A0=>nx4004, A1=>nx16513);
   ix4085 : oai32 port map ( Y=>nx4084, A0=>nx16516, A1=>nx4054, A2=>nx17826, 
      B0=>nx16983, B1=>nx16519);
   ix16520 : aoi21 port map ( Y=>nx16519, A0=>img_addr_offset_12, A1=>nx3946, 
      B0=>nx16528);
   ix4069 : aoi21 port map ( Y=>nx4068, A0=>nx16465, A1=>nx16524, B0=>nx4062
   );
   reg_img_addr_offset_12 : dffr port map ( Q=>img_addr_offset_12, QB=>
      nx16524, D=>nx14327, CLK=>clk, R=>reset);
   ix3947 : nand02 port map ( Y=>nx3946, A0=>nx16469, A1=>nx16467);
   reg_bias_offset_reg_q_13 : dffr port map ( Q=>bias_offset_data_out_13, QB
      =>nx16538, D=>nx14387, CLK=>clk, R=>reset);
   ix14368 : oai222 port map ( Y=>nx14367, A0=>nx16542, A1=>nx16951, B0=>
      nx17215, B1=>nx16547, C0=>nx17836, C1=>nx16925);
   ix16548 : xor2 port map ( Y=>nx16547, A0=>nx4154, A1=>nx16550);
   layer_mem_size_reg_q_13 : dffr port map ( Q=>layer_mem_size_out_13, QB=>
      OPEN, D=>nx14357, CLK=>clk, R=>reset);
   reg_write_base_reg_q_13 : dffr port map ( Q=>write_base_data_out_13, QB=>
      nx16555, D=>nx14367, CLK=>clk, R=>reset);
   ix16561 : oai21 port map ( Y=>nx16560, A0=>nx4108, A1=>addr1_data_13, B0
      =>nx16564);
   reg_addr1_data_13 : dffr port map ( Q=>addr1_data_13, QB=>nx16557, D=>
      nx14397, CLK=>clk, R=>reset);
   ix16565 : nand02 port map ( Y=>nx16564, A0=>addr1_data_13, A1=>nx4108);
   ix16585 : oai21 port map ( Y=>nx16584, A0=>nx4062, A1=>img_addr_offset_13, 
      B0=>nx16586);
   ix16587 : nand02 port map ( Y=>nx16586, A0=>img_addr_offset_13, A1=>
      nx4062);
   reg_img_addr_offset_13 : dffr port map ( Q=>img_addr_offset_13, QB=>
      nx16588, D=>nx14377, CLK=>clk, R=>reset);
   ix4381 : oai221 port map ( Y=>mem_addr_out(14), A0=>nx16592, A1=>nx17025, 
      B0=>nx16624, B1=>nx17017, C0=>nx16629);
   ix16593 : xnor2 port map ( Y=>nx16592, A0=>nx16594, A1=>nx16597);
   reg_bias_offset_reg_q_14 : dffr port map ( Q=>bias_offset_data_out_14, QB
      =>nx16602, D=>nx14437, CLK=>clk, R=>reset);
   layer_mem_size_reg_q_14 : dffr port map ( Q=>layer_mem_size_out_14, QB=>
      nx16621, D=>nx14407, CLK=>clk, R=>reset);
   reg_write_base_reg_q_14 : dffr port map ( Q=>write_base_data_out_14, QB=>
      nx16622, D=>nx14417, CLK=>clk, R=>reset);
   reg_addr1_data_14 : dffr port map ( Q=>addr1_data_14, QB=>nx16624, D=>
      nx14447, CLK=>clk, R=>reset);
   ix16630 : aoi322 port map ( Y=>nx16629, A0=>nx4320, A1=>nx16636, A2=>
      nx17237, B0=>nx4330, B1=>nx4336, C0=>nx4304, C1=>nx16939);
   ix4321 : or02 port map ( Y=>nx4320, A0=>nx4194, A1=>img_addr_offset_14);
   reg_img_addr_offset_14 : dffr port map ( Q=>img_addr_offset_14, QB=>
      nx16635, D=>nx14427, CLK=>clk, R=>reset);
   ix16637 : nand02 port map ( Y=>nx16636, A0=>img_addr_offset_14, A1=>
      nx4194);
   ix4331 : or02 port map ( Y=>nx4330, A0=>nx4204, A1=>
      write_base_data_out_14);
   ix4305 : xnor2 port map ( Y=>nx4304, A0=>nx4260, A1=>nx16642);
   reg_addr1_data_15 : dffr port map ( Q=>addr1_data_15, QB=>nx16650, D=>
      nx14497, CLK=>clk, R=>reset);
   ix4407 : oai22 port map ( Y=>nx4406, A0=>NOT_nx16607, A1=>nx16610, B0=>
      nx17838, B1=>nx14791);
   reg_write_base_reg_q_15 : dffs_ni port map ( Q=>write_base_data_out_15, 
      QB=>nx16661, D=>nx14477, CLK=>clk, S=>reset);
   ix16664 : xnor2 port map ( Y=>nx16663, A0=>nx18299, A1=>nx4428);
   layer_mem_size_reg_q_15 : dffr port map ( Q=>layer_mem_size_out_15, QB=>
      OPEN, D=>nx14467, CLK=>clk, R=>reset);
   reg_bias_offset_reg_q_15 : dffr port map ( Q=>OPEN, QB=>nx16677, D=>
      nx14487, CLK=>clk, R=>reset);
   img_addr_offset_15 : dffr port map ( Q=>OPEN, QB=>nx16696, D=>nx14457, 
      CLK=>clk, R=>reset);
   ix1777 : inv01 port map ( Y=>mem_data_out(0), A=>nx16699);
   ix16700 : aoi222 port map ( Y=>nx16699, A0=>comp_unit_data2_in(0), A1=>
      nx17027, B0=>comp_unit_data1_in(0), B1=>nx17029, C0=>argmax_data_in(0), 
      C1=>nx16893);
   ix1787 : inv01 port map ( Y=>mem_data_out(1), A=>nx16702);
   ix16703 : aoi222 port map ( Y=>nx16702, A0=>comp_unit_data2_in(1), A1=>
      nx17027, B0=>comp_unit_data1_in(1), B1=>nx17029, C0=>argmax_data_in(1), 
      C1=>nx16893);
   ix1797 : inv01 port map ( Y=>mem_data_out(2), A=>nx16705);
   ix16706 : aoi222 port map ( Y=>nx16705, A0=>comp_unit_data2_in(2), A1=>
      nx17027, B0=>comp_unit_data1_in(2), B1=>nx17029, C0=>argmax_data_in(2), 
      C1=>nx16893);
   ix1807 : inv01 port map ( Y=>mem_data_out(3), A=>nx16708);
   ix16709 : aoi222 port map ( Y=>nx16708, A0=>comp_unit_data2_in(3), A1=>
      nx17027, B0=>comp_unit_data1_in(3), B1=>nx17029, C0=>argmax_data_in(3), 
      C1=>nx16893);
   ix1817 : inv01 port map ( Y=>mem_data_out(4), A=>nx16711);
   ix16712 : aoi222 port map ( Y=>nx16711, A0=>comp_unit_data2_in(4), A1=>
      nx17027, B0=>comp_unit_data1_in(4), B1=>nx17029, C0=>argmax_data_in(4), 
      C1=>nx16893);
   ix1827 : inv01 port map ( Y=>mem_data_out(5), A=>nx16714);
   ix16715 : aoi222 port map ( Y=>nx16714, A0=>comp_unit_data2_in(5), A1=>
      nx17027, B0=>comp_unit_data1_in(5), B1=>nx16815, C0=>argmax_data_in(5), 
      C1=>nx16893);
   ix1837 : inv01 port map ( Y=>mem_data_out(6), A=>nx16717);
   ix16718 : aoi222 port map ( Y=>nx16717, A0=>comp_unit_data2_in(6), A1=>
      nx16809, B0=>comp_unit_data1_in(6), B1=>nx16815, C0=>argmax_data_in(6), 
      C1=>nx16895);
   ix1847 : inv01 port map ( Y=>mem_data_out(7), A=>nx16720);
   ix16721 : aoi222 port map ( Y=>nx16720, A0=>comp_unit_data2_in(7), A1=>
      nx16809, B0=>comp_unit_data1_in(7), B1=>nx16815, C0=>argmax_data_in(7), 
      C1=>nx16895);
   ix1857 : inv01 port map ( Y=>mem_data_out(8), A=>nx16723);
   ix16724 : aoi222 port map ( Y=>nx16723, A0=>comp_unit_data2_in(8), A1=>
      nx16809, B0=>comp_unit_data1_in(8), B1=>nx16815, C0=>argmax_data_in(8), 
      C1=>nx16895);
   ix1867 : inv01 port map ( Y=>mem_data_out(9), A=>nx16726);
   ix16727 : aoi222 port map ( Y=>nx16726, A0=>comp_unit_data2_in(9), A1=>
      nx16809, B0=>comp_unit_data1_in(9), B1=>nx16815, C0=>argmax_data_in(9), 
      C1=>nx16895);
   ix1877 : inv01 port map ( Y=>mem_data_out(10), A=>nx16729);
   ix16730 : aoi222 port map ( Y=>nx16729, A0=>comp_unit_data2_in(10), A1=>
      nx16809, B0=>comp_unit_data1_in(10), B1=>nx16815, C0=>
      argmax_data_in(10), C1=>nx16895);
   ix1887 : inv01 port map ( Y=>mem_data_out(11), A=>nx16732);
   ix16733 : aoi222 port map ( Y=>nx16732, A0=>comp_unit_data2_in(11), A1=>
      nx16809, B0=>comp_unit_data1_in(11), B1=>nx16815, C0=>
      argmax_data_in(11), C1=>nx16895);
   ix1897 : inv01 port map ( Y=>mem_data_out(12), A=>nx16735);
   ix16736 : aoi222 port map ( Y=>nx16735, A0=>comp_unit_data2_in(12), A1=>
      nx16809, B0=>comp_unit_data1_in(12), B1=>nx16817, C0=>
      argmax_data_in(12), C1=>nx16895);
   ix1907 : inv01 port map ( Y=>mem_data_out(13), A=>nx16738);
   ix16739 : aoi222 port map ( Y=>nx16738, A0=>comp_unit_data2_in(13), A1=>
      nx16811, B0=>comp_unit_data1_in(13), B1=>nx16817, C0=>
      argmax_data_in(13), C1=>nx16897);
   ix1917 : inv01 port map ( Y=>mem_data_out(14), A=>nx16741);
   ix16742 : aoi222 port map ( Y=>nx16741, A0=>comp_unit_data2_in(14), A1=>
      nx16811, B0=>comp_unit_data1_in(14), B1=>nx16817, C0=>
      argmax_data_in(14), C1=>nx16897);
   ix1927 : inv01 port map ( Y=>mem_data_out(15), A=>nx16744);
   ix16745 : aoi222 port map ( Y=>nx16744, A0=>comp_unit_data2_in(15), A1=>
      nx16811, B0=>comp_unit_data1_in(15), B1=>nx16817, C0=>
      argmax_data_in(15), C1=>nx16897);
   ix4055 : inv01 port map ( Y=>nx4054, A=>nx16577);
   ix3821 : inv01 port map ( Y=>nx3820, A=>nx16456);
   ix3811 : inv01 port map ( Y=>nx3810, A=>nx16469);
   ix3565 : inv01 port map ( Y=>nx3564, A=>nx16336);
   ix3555 : inv01 port map ( Y=>nx3554, A=>nx16349);
   ix3535 : inv01 port map ( Y=>nx3534, A=>nx16274);
   ix3287 : inv01 port map ( Y=>nx3286, A=>nx16218);
   ix15971 : inv01 port map ( Y=>nx15970, A=>nx2908);
   ix2775 : inv01 port map ( Y=>nx2774, A=>nx15961);
   ix2533 : inv02 port map ( Y=>nx2532, A=>nx16027);
   ix16687 : inv01 port map ( Y=>nx16686, A=>nx2520);
   ix2495 : inv01 port map ( Y=>nx2494, A=>nx15840);
   ix2479 : inv01 port map ( Y=>nx2478, A=>nx15834);
   ix2407 : inv02 port map ( Y=>nx2406, A=>nx15489);
   ix15657 : inv01 port map ( Y=>nx15656, A=>nx2372);
   ix14883 : inv01 port map ( Y=>nx14882, A=>nx12267);
   ix1675 : inv01 port map ( Y=>nx12266, A=>nx15082);
   ix1235 : inv01 port map ( Y=>nx12251, A=>nx14604);
   ix1201 : inv01 port map ( Y=>nx1200, A=>nx14887);
   ix1113 : inv01 port map ( Y=>nx1112, A=>nx15040);
   ix867 : inv01 port map ( Y=>nx866, A=>nx15531);
   ix14898 : inv01 port map ( Y=>nx14897, A=>nx830);
   ix14513 : inv01 port map ( Y=>nx14512, A=>nx794);
   ix681 : inv01 port map ( Y=>nx680, A=>nx15339);
   ix15333 : inv01 port map ( Y=>nx15332, A=>nx646);
   ix27 : inv01 port map ( Y=>nx26, A=>nx14771);
   ix489 : inv01 port map ( Y=>nx12231, A=>nx14567);
   ix5 : inv01 port map ( Y=>nx4, A=>nx15304);
   ix1745 : inv01 port map ( Y=>argmax_ready_EXMPLR, A=>nx15347);
   ix781 : inv01 port map ( Y=>comp_unit_flt_size, A=>nx15077);
   ix16750 : buf02 port map ( Y=>nx16751, A=>current_state_12);
   ix16752 : buf02 port map ( Y=>nx16753, A=>current_state_12);
   ix16754 : buf02 port map ( Y=>nx16755, A=>wind_width_count_0);
   ix16756 : buf02 port map ( Y=>nx16757, A=>wind_width_count_0);
   ix16758 : buf02 port map ( Y=>nx16759, A=>cache_width_count_4);
   ix16760 : buf02 port map ( Y=>nx16761, A=>cache_width_count_4);
   ix16762 : buf02 port map ( Y=>nx16763, A=>cache_width_count_2);
   ix16764 : buf02 port map ( Y=>nx16765, A=>cache_width_count_2);
   ix16766 : inv02 port map ( Y=>nx16767, A=>clk);
   ix16768 : inv02 port map ( Y=>nx16769, A=>clk);
   ix16770 : inv02 port map ( Y=>nx16771, A=>clk);
   ix16772 : inv02 port map ( Y=>nx16773, A=>clk);
   ix16774 : inv02 port map ( Y=>nx16775, A=>clk);
   ix16776 : inv02 port map ( Y=>nx16777, A=>clk);
   ix16778 : inv02 port map ( Y=>nx16779, A=>clk);
   ix16780 : inv02 port map ( Y=>nx16781, A=>clk);
   ix16782 : inv01 port map ( Y=>nx16783, A=>nx15077);
   ix16794 : inv01 port map ( Y=>nx16795, A=>filter_ready_out_EXMPLR);
   ix16796 : inv02 port map ( Y=>nx16797, A=>nx17193);
   ix16802 : inv02 port map ( Y=>nx16803, A=>nx14647);
   ix16804 : inv02 port map ( Y=>nx16805, A=>nx17113);
   ix16808 : inv02 port map ( Y=>nx16809, A=>nx14722);
   ix16810 : inv02 port map ( Y=>nx16811, A=>nx14722);
   ix16814 : inv02 port map ( Y=>nx16815, A=>nx14597);
   ix16816 : inv02 port map ( Y=>nx16817, A=>nx14597);
   ix16818 : inv02 port map ( Y=>nx16819, A=>nx14640);
   ix16820 : inv02 port map ( Y=>nx16821, A=>nx17109);
   ix16834 : inv02 port map ( Y=>nx16835, A=>nx17197);
   ix16836 : inv02 port map ( Y=>nx16837, A=>nx15272);
   ix16838 : inv02 port map ( Y=>nx16839, A=>nx17135);
   ix16840 : inv02 port map ( Y=>nx16841, A=>nx17215);
   ix16842 : inv02 port map ( Y=>nx16843, A=>nx17215);
   ix16846 : inv02 port map ( Y=>nx16847, A=>nx17203);
   ix16848 : inv02 port map ( Y=>nx16849, A=>nx17203);
   ix16850 : inv02 port map ( Y=>nx16851, A=>nx17203);
   ix16856 : buf02 port map ( Y=>nx16857, A=>nx684);
   ix16864 : inv01 port map ( Y=>nx16865, A=>nx874);
   ix16866 : inv02 port map ( Y=>nx16867, A=>nx16865);
   ix16868 : inv02 port map ( Y=>nx16869, A=>nx16865);
   ix16870 : inv02 port map ( Y=>nx16871, A=>nx16865);
   ix16878 : inv01 port map ( Y=>nx16879, A=>nx1278);
   ix16880 : inv02 port map ( Y=>nx16881, A=>nx16879);
   ix16882 : inv02 port map ( Y=>nx16883, A=>nx16879);
   ix16884 : inv02 port map ( Y=>nx16885, A=>nx16879);
   ix16890 : inv02 port map ( Y=>nx16891, A=>nx15223);
   ix16892 : inv02 port map ( Y=>nx16893, A=>nx15758);
   ix16894 : inv02 port map ( Y=>nx16895, A=>nx15758);
   ix16896 : inv02 port map ( Y=>nx16897, A=>nx15758);
   ix16912 : inv02 port map ( Y=>nx16913, A=>nx15747);
   ix16914 : inv02 port map ( Y=>nx16915, A=>nx15747);
   ix16916 : inv02 port map ( Y=>nx16917, A=>nx15747);
   ix16922 : inv02 port map ( Y=>nx16923, A=>nx15791);
   ix16924 : inv02 port map ( Y=>nx16925, A=>nx15791);
   ix16926 : inv02 port map ( Y=>nx16927, A=>nx15791);
   ix16934 : inv02 port map ( Y=>nx16935, A=>nx16686);
   ix16936 : inv02 port map ( Y=>nx16937, A=>nx16686);
   ix16938 : inv02 port map ( Y=>nx16939, A=>nx16686);
   ix16940 : inv02 port map ( Y=>nx16941, A=>current_state_24);
   ix16944 : inv02 port map ( Y=>nx16945, A=>current_state_24);
   ix16946 : inv02 port map ( Y=>nx16947, A=>nx492);
   ix16948 : inv02 port map ( Y=>nx16949, A=>nx17069);
   ix16950 : inv02 port map ( Y=>nx16951, A=>nx17069);
   ix16952 : buf02 port map ( Y=>nx16953, A=>nx14644);
   ix16954 : buf02 port map ( Y=>nx16955, A=>nx14644);
   ix16960 : buf02 port map ( Y=>nx16961, A=>nx15032);
   ix16962 : inv02 port map ( Y=>nx16963, A=>current_state_17);
   ix16966 : inv02 port map ( Y=>nx16967, A=>nx17075);
   ix16968 : inv02 port map ( Y=>nx16969, A=>nx17075);
   ix16970 : inv02 port map ( Y=>nx16971, A=>nx17075);
   ix16976 : inv02 port map ( Y=>nx16977, A=>nx17083);
   ix16978 : inv02 port map ( Y=>nx16979, A=>nx17083);
   ix16980 : inv02 port map ( Y=>nx16981, A=>nx17083);
   ix16982 : inv02 port map ( Y=>nx16983, A=>nx17083);
   ix16984 : inv02 port map ( Y=>nx16985, A=>nx17083);
   ix17008 : inv02 port map ( Y=>nx17009, A=>nx2572);
   ix17010 : inv02 port map ( Y=>nx17011, A=>nx17089);
   ix17012 : inv02 port map ( Y=>nx17013, A=>nx17089);
   ix17014 : inv02 port map ( Y=>nx17015, A=>nx17089);
   ix17016 : inv02 port map ( Y=>nx17017, A=>nx17089);
   ix17018 : inv02 port map ( Y=>nx17019, A=>nx2472);
   ix17020 : inv02 port map ( Y=>nx17021, A=>nx2472);
   ix17022 : inv02 port map ( Y=>nx17023, A=>nx2532);
   ix17026 : inv02 port map ( Y=>nx17027, A=>nx14722);
   ix17028 : inv02 port map ( Y=>nx17029, A=>nx14597);
   ix17034 : inv01 port map ( Y=>nx17035, A=>nx17247);
   ix17036 : inv01 port map ( Y=>nx17037, A=>nx17247);
   ix17038 : inv02 port map ( Y=>nx17039, A=>nx17155);
   ix14516 : xor2 port map ( Y=>nx14515, A0=>nx14553, A1=>nx786);
   ix12788 : mux21_ni port map ( Y=>nx12787, A0=>nx740, A1=>
      cntr1_inst_counter_out_4, S0=>nx17097);
   ix741 : xor2 port map ( Y=>nx740, A0=>nx14553, A1=>nx14520);
   ix12778 : mux21_ni port map ( Y=>nx12777, A0=>nx722, A1=>
      cntr1_inst_counter_out_3, S0=>nx17097);
   ix723 : xor2 port map ( Y=>nx722, A0=>nx14561, A1=>nx14525);
   ix12768 : mux21_ni port map ( Y=>nx12767, A0=>nx708, A1=>
      cntr1_inst_counter_out_2, S0=>nx17097);
   ix709 : xor2 port map ( Y=>nx708, A0=>nx14542, A1=>nx14530);
   ix12758 : mux21 port map ( Y=>nx12757, A0=>nx15336, A1=>nx14534, S0=>
      nx17097);
   ix14541 : xnor2 port map ( Y=>nx14540, A0=>nx17099, A1=>
      cntr1_inst_counter_out_2);
   ix14545 : xnor2 port map ( Y=>nx14544, A0=>nx17099, A1=>
      cntr1_inst_counter_out_5);
   ix12798 : mux21 port map ( Y=>nx12797, A0=>nx14549, A1=>nx14546, S0=>
      nx17099);
   ix14550 : xor2 port map ( Y=>nx14549, A0=>nx14546, A1=>nx12238);
   ix747 : nor02ii port map ( Y=>nx12238, A0=>nx14520, A1=>
      cntr1_inst_counter_out_4);
   ix729 : xor2 port map ( Y=>nx728, A0=>nx17099, A1=>
      cntr1_inst_counter_out_0);
   ix703 : xnor2 port map ( Y=>nx702, A0=>nx17099, A1=>nx14534);
   ix607 : or02 port map ( Y=>nx12230, A0=>current_state_1, A1=>
      current_state_24);
   ix601 : and03 port map ( Y=>nx600, A0=>nx17069, A1=>nx15240, A2=>nx17045
   );
   ix17044 : inv01 port map ( Y=>nx17045, A=>nx15274);
   ix1241 : ao32 port map ( Y=>nx1240, A0=>nx14604, A1=>current_state_20, A2
      =>nx14871, B0=>nx16803, B1=>ftc_cntrl_reg_out_12);
   ix14605 : or02 port map ( Y=>nx14604, A0=>ftc_cntrl_reg_out_14, A1=>
      nx15077);
   ix1585 : or02 port map ( Y=>nx1584, A0=>nx14871, A1=>nx15075);
   ix1451 : and04 port map ( Y=>nx1450, A0=>nx14632, A1=>nx15097, A2=>
      nx15106, A3=>nx15111);
   ix13278 : mux21 port map ( Y=>nx13277, A0=>nx15094, A1=>nx14632, S0=>
      nx17123);
   ix827 : nor02ii port map ( Y=>nx12239, A0=>nx17109, A1=>nx14865);
   ix14645 : and04 port map ( Y=>nx14644, A0=>nx14988, A1=>nx14867, A2=>
      nx15092, A3=>nx15075);
   ix14657 : xor2 port map ( Y=>nx14656, A0=>nx14782, A1=>
      new_size_squared_out_15);
   ix14661 : xor2 port map ( Y=>nx14660, A0=>nx14782, A1=>nx334);
   ix335 : nor02ii port map ( Y=>nx334, A0=>nx14669, A1=>
      write_offset_data_out_14);
   ix12558 : ao22 port map ( Y=>nx12557, A0=>write_offset_data_out_14, A1=>
      nx17203, B0=>nx340, B1=>nx17047);
   ix17046 : inv01 port map ( Y=>nx17047, A=>nx14717);
   ix289 : nor02ii port map ( Y=>nx288, A0=>nx14682, A1=>
      write_offset_data_out_12);
   ix12518 : ao22 port map ( Y=>nx12517, A0=>write_offset_data_out_12, A1=>
      nx17203, B0=>nx294, B1=>nx17049);
   ix17048 : inv01 port map ( Y=>nx17049, A=>nx16959);
   ix241 : nor02ii port map ( Y=>nx240, A0=>nx14695, A1=>
      write_offset_data_out_10);
   ix12478 : ao22 port map ( Y=>nx12477, A0=>write_offset_data_out_10, A1=>
      nx17203, B0=>nx246, B1=>nx17049);
   ix195 : nor02ii port map ( Y=>nx194, A0=>nx14708, A1=>
      write_offset_data_out_8);
   ix12438 : ao22 port map ( Y=>nx12437, A0=>write_offset_data_out_8, A1=>
      nx17203, B0=>nx200, B1=>nx17049);
   ix14718 : and02 port map ( Y=>nx14717, A0=>nx14597, A1=>nx14722);
   ix1247 : nor02_2x port map ( Y=>nx1246, A0=>nx14597, A1=>nx15077);
   ix145 : nor02ii port map ( Y=>nx144, A0=>nx14732, A1=>
      write_offset_data_out_6);
   ix12398 : ao22 port map ( Y=>nx12397, A0=>write_offset_data_out_6, A1=>
      nx17205, B0=>nx150, B1=>nx17049);
   ix99 : nor02ii port map ( Y=>nx98, A0=>nx14747, A1=>
      write_offset_data_out_4);
   ix12358 : ao22 port map ( Y=>nx12357, A0=>write_offset_data_out_4, A1=>
      nx17205, B0=>nx104, B1=>nx17051);
   ix17050 : inv01 port map ( Y=>nx17051, A=>nx16957);
   ix14748 : or04 port map ( Y=>nx14747, A0=>nx14751, A1=>nx14756, A2=>
      nx17803, A3=>nx17807);
   ix12338 : ao22 port map ( Y=>nx12337, A0=>write_offset_data_out_3, A1=>
      nx17205, B0=>nx78, B1=>nx17051);
   ix12278 : mux21 port map ( Y=>nx12277, A0=>nx16847, A1=>nx16957, S0=>
      nx17807);
   ix14772 : or02 port map ( Y=>nx14771, A0=>nx17803, A1=>nx17807);
   ix14775 : or03 port map ( Y=>nx14774, A0=>nx14756, A1=>nx17803, A2=>
      nx17807);
   ix12588 : mux21_ni port map ( Y=>nx12587, A0=>mem_data_in(15), A1=>
      new_size_squared_out_15, S0=>nx17197);
   ix14788 : xnor2 port map ( Y=>nx14787, A0=>nx14663, A1=>nx14791);
   ix12568 : mux21_ni port map ( Y=>nx12567, A0=>mem_data_in(14), A1=>
      new_size_squared_out_14, S0=>nx17197);
   ix14793 : xor2 port map ( Y=>nx14792, A0=>nx14780, A1=>
      new_size_squared_out_13);
   ix12548 : mux21_ni port map ( Y=>nx12547, A0=>mem_data_in(13), A1=>
      new_size_squared_out_13, S0=>nx17197);
   ix14798 : xnor2 port map ( Y=>nx14797, A0=>nx14676, A1=>nx14801);
   ix12528 : mux21_ni port map ( Y=>nx12527, A0=>mem_data_in(12), A1=>
      new_size_squared_out_12, S0=>nx17197);
   ix14804 : xor2 port map ( Y=>nx14803, A0=>nx14778, A1=>
      new_size_squared_out_11);
   ix12508 : mux21_ni port map ( Y=>nx12507, A0=>mem_data_in(11), A1=>
      new_size_squared_out_11, S0=>nx17197);
   ix14809 : xnor2 port map ( Y=>nx14808, A0=>nx14689, A1=>nx14812);
   ix12488 : mux21_ni port map ( Y=>nx12487, A0=>mem_data_in(10), A1=>
      new_size_squared_out_10, S0=>nx17197);
   ix14814 : xor2 port map ( Y=>nx14813, A0=>nx14776, A1=>
      new_size_squared_out_9);
   ix12468 : mux21_ni port map ( Y=>nx12467, A0=>mem_data_in(9), A1=>
      new_size_squared_out_9, S0=>nx17199);
   ix14819 : xnor2 port map ( Y=>nx14818, A0=>nx14702, A1=>nx14822);
   ix12448 : mux21_ni port map ( Y=>nx12447, A0=>mem_data_in(8), A1=>
      new_size_squared_out_8, S0=>nx17199);
   ix14825 : xor2 port map ( Y=>nx14824, A0=>nx14712, A1=>
      new_size_squared_out_7);
   ix12428 : mux21_ni port map ( Y=>nx12427, A0=>mem_data_in(7), A1=>
      new_size_squared_out_7, S0=>nx17199);
   ix14830 : xnor2 port map ( Y=>nx14829, A0=>nx14726, A1=>nx14833);
   ix12408 : mux21_ni port map ( Y=>nx12407, A0=>mem_data_in(6), A1=>
      new_size_squared_out_6, S0=>nx17199);
   ix14835 : xor2 port map ( Y=>nx14834, A0=>nx14736, A1=>
      new_size_squared_out_5);
   ix12388 : mux21_ni port map ( Y=>nx12387, A0=>mem_data_in(5), A1=>
      new_size_squared_out_5, S0=>nx17199);
   ix14840 : xnor2 port map ( Y=>nx14839, A0=>nx14741, A1=>nx14843);
   ix12368 : mux21_ni port map ( Y=>nx12367, A0=>mem_data_in(4), A1=>
      new_size_squared_out_4, S0=>nx17199);
   ix14846 : xor2 port map ( Y=>nx14845, A0=>nx14751, A1=>
      new_size_squared_out_3);
   ix12348 : mux21_ni port map ( Y=>nx12347, A0=>mem_data_in(3), A1=>
      new_size_squared_out_3, S0=>nx17199);
   ix14851 : xnor2 port map ( Y=>nx14850, A0=>nx14756, A1=>nx14854);
   ix12328 : mux21_ni port map ( Y=>nx12327, A0=>mem_data_in(2), A1=>
      new_size_squared_out_2, S0=>nx17201);
   ix14856 : xor2 port map ( Y=>nx14855, A0=>nx17803, A1=>
      new_size_squared_out_1);
   ix12308 : mux21_ni port map ( Y=>nx12307, A0=>mem_data_in(1), A1=>
      new_size_squared_out_1, S0=>nx17201);
   ix14861 : xor2 port map ( Y=>nx14860, A0=>nx17808, A1=>
      new_size_squared_out_0);
   ix12288 : mux21_ni port map ( Y=>nx12287, A0=>mem_data_in(0), A1=>
      new_size_squared_out_0, S0=>nx17201);
   ix1531 : or02 port map ( Y=>nx12265, A0=>ftc_cntrl_reg_out_11, A1=>
      nx15092);
   ix14874 : or03 port map ( Y=>nx14873, A0=>ftc_cntrl_reg_out_8, A1=>
      nx14867, A2=>nx15087);
   ix1053 : and04 port map ( Y=>nx1052, A0=>nx14892, A1=>nx14905, A2=>
      nx14914, A3=>nx14919);
   ix13008 : mux21 port map ( Y=>nx13007, A0=>nx14902, A1=>nx14892, S0=>
      nx17117);
   ix14900 : or02 port map ( Y=>nx14899, A0=>nx17113, A1=>nx14884);
   ix14903 : xor2 port map ( Y=>nx14902, A0=>nx14892, A1=>nx12241);
   ix1033 : nor02ii port map ( Y=>nx12241, A0=>nx14910, A1=>
      cache_width_cntr_counter_out_14);
   ix12998 : mux21_ni port map ( Y=>nx12997, A0=>nx1026, A1=>
      cache_width_cntr_counter_out_14, S0=>nx17117);
   ix1027 : xor2 port map ( Y=>nx1026, A0=>nx14905, A1=>nx14910);
   ix12988 : mux21 port map ( Y=>nx12987, A0=>nx14916, A1=>nx14914, S0=>
      nx17117);
   ix1009 : nor02ii port map ( Y=>nx12243, A0=>nx14924, A1=>
      cache_width_cntr_counter_out_12);
   ix12978 : mux21_ni port map ( Y=>nx12977, A0=>nx1002, A1=>
      cache_width_cntr_counter_out_12, S0=>nx17117);
   ix1003 : xor2 port map ( Y=>nx1002, A0=>nx14919, A1=>nx14924);
   ix12968 : mux21 port map ( Y=>nx12967, A0=>nx14930, A1=>nx14928, S0=>
      nx17117);
   ix985 : nor02ii port map ( Y=>nx12245, A0=>nx14938, A1=>
      cache_width_cntr_counter_out_10);
   ix12958 : mux21_ni port map ( Y=>nx12957, A0=>nx978, A1=>
      cache_width_cntr_counter_out_10, S0=>nx17117);
   ix979 : xor2 port map ( Y=>nx978, A0=>nx14933, A1=>nx14938);
   ix12948 : mux21 port map ( Y=>nx12947, A0=>nx14944, A1=>nx14942, S0=>
      nx17117);
   ix961 : nor02ii port map ( Y=>nx12247, A0=>nx14952, A1=>
      cache_width_cntr_counter_out_8);
   ix12938 : mux21_ni port map ( Y=>nx12937, A0=>nx954, A1=>
      cache_width_cntr_counter_out_8, S0=>nx17119);
   ix955 : xor2 port map ( Y=>nx954, A0=>nx14947, A1=>nx14952);
   ix12928 : mux21 port map ( Y=>nx12927, A0=>nx14958, A1=>nx14956, S0=>
      nx17119);
   ix937 : nor02ii port map ( Y=>nx12249, A0=>nx14966, A1=>
      cache_width_cntr_counter_out_6);
   ix12918 : mux21_ni port map ( Y=>nx12917, A0=>nx930, A1=>
      cache_width_cntr_counter_out_6, S0=>nx17119);
   ix931 : xor2 port map ( Y=>nx930, A0=>nx14961, A1=>nx14966);
   ix14967 : or03 port map ( Y=>nx14966, A0=>nx17053, A1=>nx15012, A2=>
      nx14971);
   ix17052 : inv01 port map ( Y=>nx17053, A=>nx16761);
   ix12898 : mux21_ni port map ( Y=>nx12897, A0=>nx904, A1=>nx16759, S0=>
      nx17119);
   ix12868 : mux21_ni port map ( Y=>nx12867, A0=>nx880, A1=>
      cache_width_count_1, S0=>nx17119);
   ix12858 : xor2 port map ( Y=>nx12857, A0=>cache_width_count_0, A1=>
      nx17245);
   ix14986 : mux21_ni port map ( Y=>nx14985, A0=>cache_height_count_en, A1=>
      nx16803, S0=>nx17109);
   ix14989 : and02 port map ( Y=>nx14988, A0=>nx17109, A1=>nx17113);
   ix863 : nor02ii port map ( Y=>nx862, A0=>nx14990, A1=>
      ftc_cntrl_reg_out_10);
   ix12878 : mux21_ni port map ( Y=>nx12877, A0=>nx888, A1=>nx16763, S0=>
      nx17119);
   ix12888 : mux21_ni port map ( Y=>nx12887, A0=>nx896, A1=>
      cache_width_count_3, S0=>nx17119);
   ix12908 : mux21 port map ( Y=>nx12907, A0=>nx15014, A1=>nx15012, S0=>
      nx17121);
   ix1067 : and04 port map ( Y=>nx1066, A0=>nx14928, A1=>nx14933, A2=>
      nx14942, A3=>nx14947);
   ix1099 : and04 port map ( Y=>nx1098, A0=>nx14956, A1=>nx14961, A2=>
      nx15012, A3=>nx17055);
   ix1091 : xnor2 port map ( Y=>nx17055, A0=>nx15029, A1=>
      cache_width_count_0);
   ix13028 : oai221 port map ( Y=>nx13027, A0=>nx17215, A1=>nx17057, B0=>
      nx15029, B1=>nx17059, C0=>nx15297);
   ix17056 : inv01 port map ( Y=>nx17057, A=>new_width_out_0);
   ix17058 : inv01 port map ( Y=>nx17059, A=>nx15027);
   ix15028 : and02 port map ( Y=>nx15027, A0=>nx15297, A1=>nx16945);
   ix15041 : nor02ii port map ( Y=>nx15040, A0=>img_width_out_1, A1=>nx15029
   );
   ix1535 : ao21 port map ( Y=>nx1534, A0=>nx17111, A1=>nx17115, B0=>
      current_state_15);
   ix15095 : xor2 port map ( Y=>nx15094, A0=>nx14632, A1=>nx12254);
   ix1431 : nor02ii port map ( Y=>nx12254, A0=>nx15102, A1=>
      window_width_cntr_counter_out_14);
   ix13268 : mux21_ni port map ( Y=>nx13267, A0=>nx1424, A1=>
      window_width_cntr_counter_out_14, S0=>nx17123);
   ix1425 : xor2 port map ( Y=>nx1424, A0=>nx15097, A1=>nx15102);
   ix13258 : mux21 port map ( Y=>nx13257, A0=>nx15108, A1=>nx15106, S0=>
      nx17123);
   ix1407 : nor02ii port map ( Y=>nx12256, A0=>nx15116, A1=>
      window_width_cntr_counter_out_12);
   ix13248 : mux21_ni port map ( Y=>nx13247, A0=>nx1400, A1=>
      window_width_cntr_counter_out_12, S0=>nx17123);
   ix1401 : xor2 port map ( Y=>nx1400, A0=>nx15111, A1=>nx15116);
   ix13238 : mux21 port map ( Y=>nx13237, A0=>nx15122, A1=>nx15120, S0=>
      nx17123);
   ix1383 : nor02ii port map ( Y=>nx12258, A0=>nx15130, A1=>
      window_width_cntr_counter_out_10);
   ix13228 : mux21_ni port map ( Y=>nx13227, A0=>nx1376, A1=>
      window_width_cntr_counter_out_10, S0=>nx17123);
   ix1377 : xor2 port map ( Y=>nx1376, A0=>nx15125, A1=>nx15130);
   ix13218 : mux21 port map ( Y=>nx13217, A0=>nx15136, A1=>nx15134, S0=>
      nx17123);
   ix1359 : nor02ii port map ( Y=>nx12260, A0=>nx15144, A1=>
      window_width_cntr_counter_out_8);
   ix13208 : mux21_ni port map ( Y=>nx13207, A0=>nx1352, A1=>
      window_width_cntr_counter_out_8, S0=>nx17125);
   ix1353 : xor2 port map ( Y=>nx1352, A0=>nx15139, A1=>nx15144);
   ix13198 : mux21 port map ( Y=>nx13197, A0=>nx15150, A1=>nx15148, S0=>
      nx17125);
   ix1335 : nor02ii port map ( Y=>nx12262, A0=>nx15158, A1=>
      window_width_cntr_counter_out_6);
   ix13188 : mux21_ni port map ( Y=>nx13187, A0=>nx1328, A1=>
      window_width_cntr_counter_out_6, S0=>nx17125);
   ix1329 : xor2 port map ( Y=>nx1328, A0=>nx15153, A1=>nx15158);
   ix15159 : or03 port map ( Y=>nx15158, A0=>nx17061, A1=>nx15192, A2=>
      nx15163);
   ix17060 : inv01 port map ( Y=>nx17061, A=>wind_width_count_4);
   ix13318 : mux21_ni port map ( Y=>nx13317, A0=>nx1692, A1=>
      wind_width_count_4, S0=>nx17125);
   ix13148 : mux21_ni port map ( Y=>nx13147, A0=>nx1284, A1=>
      wind_width_count_1, S0=>nx17125);
   ix13138 : xor2 port map ( Y=>nx13137, A0=>nx16755, A1=>nx12253);
   ix13158 : mux21_ni port map ( Y=>nx13157, A0=>nx1292, A1=>
      wind_width_count_2, S0=>nx17125);
   ix13168 : mux21_ni port map ( Y=>nx13167, A0=>nx1300, A1=>
      wind_width_count_3, S0=>nx17125);
   ix13178 : mux21 port map ( Y=>nx13177, A0=>nx15194, A1=>nx15192, S0=>
      nx17127);
   ix1465 : and04 port map ( Y=>nx1464, A0=>nx15120, A1=>nx15125, A2=>
      nx15134, A3=>nx15139);
   ix1487 : and04 port map ( Y=>nx1486, A0=>nx15148, A1=>nx15153, A2=>
      nx15192, A3=>nx17063);
   ix17062 : inv01 port map ( Y=>nx17063, A=>nx1478);
   ix1489 : nor02ii port map ( Y=>nx1488, A0=>nx16961, A1=>nx17071);
   ix1505 : nor02ii port map ( Y=>nx1504, A0=>nx15055, A1=>nx17073);
   ix1509 : nor02ii port map ( Y=>nx1508, A0=>nx15064, A1=>nx17073);
   ix15217 : nor02ii port map ( Y=>nx15216, A0=>nx12267, A1=>nx14867);
   ix1663 : nor02ii port map ( Y=>nx12267, A0=>nx17115, A1=>nx14884);
   ix1623 : ao32 port map ( Y=>nx1622, A0=>nx14875, A1=>current_state_14, A2
      =>nx15087, B0=>current_state_15, B1=>ftc_cntrl_reg_out_11);
   ix1629 : nor02_2x port map ( Y=>nx1628, A0=>nx17129, A1=>nx15077);
   ix507 : mux21_ni port map ( Y=>nx506, A0=>mem_data_in(0), A1=>nx15242, S0
      =>nx17135);
   ix525 : mux21 port map ( Y=>nx524, A0=>nx15251, A1=>nx15247, S0=>nx17135
   );
   ix15250 : nor02ii port map ( Y=>nx15249, A0=>
      nflt_layer_cntr_counter_out_1, A1=>nx15242);
   ix545 : mux21 port map ( Y=>nx544, A0=>nx15259, A1=>nx15257, S0=>nx17135
   );
   ix561 : mux21 port map ( Y=>nx560, A0=>nx15269, A1=>nx15265, S0=>nx17135
   );
   ix12718 : mux21_ni port map ( Y=>nx12717, A0=>mem_data_in(1), A1=>
      nlayers_counter_out_1, S0=>nx14585);
   ix12708 : mux21_ni port map ( Y=>nx12707, A0=>mem_data_in(2), A1=>
      nlayers_counter_out_2, S0=>nx14585);
   ix12698 : mux21_ni port map ( Y=>nx12697, A0=>mem_data_in(0), A1=>
      nlayers_counter_out_0, S0=>nx14585);
   ix12598 : mux21_ni port map ( Y=>nx12597, A0=>mem_data_in(0), A1=>
      nflt_layer_temp_0, S0=>nx17135);
   ix427 : ao21 port map ( Y=>nx426, A0=>nx14571, A1=>nx15304, B0=>
      current_state_1);
   ix15305 : and03 port map ( Y=>nx15304, A0=>nx15297, A1=>nx16945, A2=>
      nx14585);
   ix15312 : nor02ii port map ( Y=>nx15311, A0=>num_channels_counter_out_1, 
      A1=>nx14571);
   ix12618 : mux21_ni port map ( Y=>nx12617, A0=>mem_data_in(1), A1=>
      nflt_layer_temp_1, S0=>nx17137);
   ix12638 : mux21_ni port map ( Y=>nx12637, A0=>mem_data_in(2), A1=>
      nflt_layer_temp_2, S0=>nx17137);
   ix787 : or02 port map ( Y=>nx786, A0=>nx15077, A1=>nx17099);
   ix493 : nor02ii port map ( Y=>nx492, A0=>nx14715, A1=>nx14567);
   ix1743 : or04 port map ( Y=>nx1742, A0=>class_cntr_counter_out_0, A1=>
      nx17809, A2=>class_cntr_counter_out_2, A3=>nx15374);
   ix13328 : mux21 port map ( Y=>nx13327, A0=>current_state_25, A1=>nx17139, 
      S0=>nx15350);
   ix13338 : mux21 port map ( Y=>nx13337, A0=>nx15360, A1=>nx17809, S0=>
      nx17139);
   ix15363 : or02 port map ( Y=>nx15362, A0=>nx17809, A1=>nx15350);
   ix13348 : mux21_ni port map ( Y=>nx13347, A0=>nx1720, A1=>
      class_cntr_counter_out_2, S0=>nx17139);
   ix1721 : xor2 port map ( Y=>nx1720, A0=>nx15364, A1=>nx15362);
   ix13358 : mux21_ni port map ( Y=>nx13357, A0=>nx1728, A1=>
      class_cntr_counter_out_3, S0=>nx17139);
   ix1729 : xor2 port map ( Y=>nx1728, A0=>nx15374, A1=>nx15372);
   ix15373 : or03 port map ( Y=>nx15372, A0=>nx15364, A1=>nx17809, A2=>
      nx15350);
   ix4543 : nor02ii port map ( Y=>argmax_data_out(0), A0=>nx17139, A1=>
      mem_data_in(0));
   ix4545 : nor02ii port map ( Y=>argmax_data_out(1), A0=>nx17139, A1=>
      mem_data_in(1));
   ix4547 : nor02ii port map ( Y=>argmax_data_out(2), A0=>nx17141, A1=>
      mem_data_in(2));
   ix4549 : nor02ii port map ( Y=>argmax_data_out(3), A0=>nx17141, A1=>
      mem_data_in(3));
   ix4551 : nor02ii port map ( Y=>argmax_data_out(4), A0=>nx17141, A1=>
      mem_data_in(4));
   ix4553 : nor02ii port map ( Y=>argmax_data_out(5), A0=>nx17141, A1=>
      mem_data_in(5));
   ix4555 : nor02ii port map ( Y=>argmax_data_out(6), A0=>nx17141, A1=>
      mem_data_in(6));
   ix4557 : nor02ii port map ( Y=>argmax_data_out(7), A0=>nx17141, A1=>
      mem_data_in(7));
   ix4559 : nor02ii port map ( Y=>argmax_data_out(8), A0=>nx17141, A1=>
      mem_data_in(8));
   ix4561 : nor02ii port map ( Y=>argmax_data_out(9), A0=>nx17143, A1=>
      mem_data_in(9));
   ix4563 : nor02ii port map ( Y=>argmax_data_out(10), A0=>nx17143, A1=>
      mem_data_in(10));
   ix4565 : nor02ii port map ( Y=>argmax_data_out(11), A0=>nx17143, A1=>
      mem_data_in(11));
   ix4567 : nor02ii port map ( Y=>argmax_data_out(12), A0=>nx17143, A1=>
      mem_data_in(12));
   ix4569 : nor02ii port map ( Y=>argmax_data_out(13), A0=>nx17143, A1=>
      mem_data_in(13));
   ix4571 : nor02ii port map ( Y=>argmax_data_out(14), A0=>nx17143, A1=>
      mem_data_in(14));
   ix4573 : nor02ii port map ( Y=>argmax_data_out(15), A0=>nx17143, A1=>
      mem_data_in(15));
   ix4575 : and02 port map ( Y=>comp_unit_data2_out(0), A0=>nx17075, A1=>
      nx1960);
   ix1961 : mux21_ni port map ( Y=>nx1960, A0=>flt_bias_out_0, A1=>
      mem_data_in(0), S0=>nx17149);
   ix13378 : mux21_ni port map ( Y=>nx13377, A0=>mem_data_in(0), A1=>
      flt_bias_out_0, S0=>nx17209);
   ix1949 : or03 port map ( Y=>nx16905, A0=>comp_unit_operation_EXMPLR, A1=>
      nx15329, A2=>layer_type_out_1);
   ix4577 : and02 port map ( Y=>comp_unit_data2_out(1), A0=>nx17077, A1=>
      nx1994);
   ix1995 : mux21_ni port map ( Y=>nx1994, A0=>flt_bias_out_1, A1=>
      mem_data_in(1), S0=>nx17149);
   ix13398 : mux21_ni port map ( Y=>nx13397, A0=>mem_data_in(1), A1=>
      flt_bias_out_1, S0=>nx17209);
   ix4579 : and02 port map ( Y=>comp_unit_data2_out(2), A0=>nx17077, A1=>
      nx2020);
   ix2021 : mux21_ni port map ( Y=>nx2020, A0=>flt_bias_out_2, A1=>
      mem_data_in(2), S0=>nx17149);
   ix13418 : mux21_ni port map ( Y=>nx13417, A0=>mem_data_in(2), A1=>
      flt_bias_out_2, S0=>nx17209);
   ix4581 : and02 port map ( Y=>comp_unit_data2_out(3), A0=>nx17077, A1=>
      nx2046);
   ix2047 : mux21_ni port map ( Y=>nx2046, A0=>flt_bias_out_3, A1=>
      mem_data_in(3), S0=>nx17149);
   ix13438 : mux21_ni port map ( Y=>nx13437, A0=>mem_data_in(3), A1=>
      flt_bias_out_3, S0=>nx17209);
   ix4583 : and02 port map ( Y=>comp_unit_data2_out(4), A0=>nx17077, A1=>
      nx2072);
   ix2073 : mux21_ni port map ( Y=>nx2072, A0=>flt_bias_out_4, A1=>
      mem_data_in(4), S0=>nx17151);
   ix13458 : mux21_ni port map ( Y=>nx13457, A0=>mem_data_in(4), A1=>
      flt_bias_out_4, S0=>nx17209);
   ix4585 : and02 port map ( Y=>comp_unit_data2_out(5), A0=>nx17077, A1=>
      nx2098);
   ix2099 : mux21_ni port map ( Y=>nx2098, A0=>flt_bias_out_5, A1=>
      mem_data_in(5), S0=>nx17151);
   ix13478 : mux21_ni port map ( Y=>nx13477, A0=>mem_data_in(5), A1=>
      flt_bias_out_5, S0=>nx17209);
   ix4587 : and02 port map ( Y=>comp_unit_data2_out(6), A0=>nx17077, A1=>
      nx2124);
   ix2125 : mux21_ni port map ( Y=>nx2124, A0=>flt_bias_out_6, A1=>
      mem_data_in(6), S0=>nx17151);
   ix13498 : mux21_ni port map ( Y=>nx13497, A0=>mem_data_in(6), A1=>
      flt_bias_out_6, S0=>nx17209);
   ix4589 : and02 port map ( Y=>comp_unit_data2_out(7), A0=>nx17077, A1=>
      nx2150);
   ix2151 : mux21_ni port map ( Y=>nx2150, A0=>flt_bias_out_7, A1=>
      mem_data_in(7), S0=>nx17151);
   ix13518 : mux21_ni port map ( Y=>nx13517, A0=>mem_data_in(7), A1=>
      flt_bias_out_7, S0=>nx17211);
   ix4591 : and02 port map ( Y=>comp_unit_data2_out(8), A0=>nx17079, A1=>
      nx2176);
   ix2177 : mux21_ni port map ( Y=>nx2176, A0=>flt_bias_out_8, A1=>
      mem_data_in(8), S0=>nx17151);
   ix13538 : mux21_ni port map ( Y=>nx13537, A0=>mem_data_in(8), A1=>
      flt_bias_out_8, S0=>nx17211);
   ix4593 : and02 port map ( Y=>comp_unit_data2_out(9), A0=>nx17079, A1=>
      nx2202);
   ix2203 : mux21_ni port map ( Y=>nx2202, A0=>flt_bias_out_9, A1=>
      mem_data_in(9), S0=>nx17151);
   ix13558 : mux21_ni port map ( Y=>nx13557, A0=>mem_data_in(9), A1=>
      flt_bias_out_9, S0=>nx17211);
   ix4595 : and02 port map ( Y=>comp_unit_data2_out(10), A0=>nx17079, A1=>
      nx2228);
   ix2229 : mux21_ni port map ( Y=>nx2228, A0=>flt_bias_out_10, A1=>
      mem_data_in(10), S0=>nx17151);
   ix13578 : mux21_ni port map ( Y=>nx13577, A0=>mem_data_in(10), A1=>
      flt_bias_out_10, S0=>nx17211);
   ix4597 : and02 port map ( Y=>comp_unit_data2_out(11), A0=>nx17079, A1=>
      nx2254);
   ix2255 : mux21_ni port map ( Y=>nx2254, A0=>flt_bias_out_11, A1=>
      mem_data_in(11), S0=>nx17153);
   ix13598 : mux21_ni port map ( Y=>nx13597, A0=>mem_data_in(11), A1=>
      flt_bias_out_11, S0=>nx17211);
   ix4599 : and02 port map ( Y=>comp_unit_data2_out(12), A0=>nx17079, A1=>
      nx2280);
   ix2281 : mux21_ni port map ( Y=>nx2280, A0=>flt_bias_out_12, A1=>
      mem_data_in(12), S0=>nx17153);
   ix13618 : mux21_ni port map ( Y=>nx13617, A0=>mem_data_in(12), A1=>
      flt_bias_out_12, S0=>nx17211);
   ix4601 : and02 port map ( Y=>comp_unit_data2_out(13), A0=>nx17079, A1=>
      nx2306);
   ix2307 : mux21_ni port map ( Y=>nx2306, A0=>flt_bias_out_13, A1=>
      mem_data_in(13), S0=>nx17153);
   ix13638 : mux21_ni port map ( Y=>nx13637, A0=>mem_data_in(13), A1=>
      flt_bias_out_13, S0=>nx17211);
   ix4603 : and02 port map ( Y=>comp_unit_data2_out(14), A0=>nx17079, A1=>
      nx2332);
   ix2333 : mux21_ni port map ( Y=>nx2332, A0=>flt_bias_out_14, A1=>
      mem_data_in(14), S0=>nx17153);
   ix13658 : mux21_ni port map ( Y=>nx13657, A0=>mem_data_in(14), A1=>
      flt_bias_out_14, S0=>nx17213);
   ix4605 : and02 port map ( Y=>comp_unit_data2_out(15), A0=>nx17081, A1=>
      nx2358);
   ix2359 : mux21_ni port map ( Y=>nx2358, A0=>flt_bias_out_15, A1=>
      mem_data_in(15), S0=>nx17153);
   ix13678 : mux21_ni port map ( Y=>nx13677, A0=>mem_data_in(15), A1=>
      flt_bias_out_15, S0=>nx17213);
   ix2409 : and02 port map ( Y=>cache_data_in_0, A0=>mem_data_in(0), A1=>
      nx17237);
   ix2411 : and02 port map ( Y=>cache_data_in_1, A0=>mem_data_in(1), A1=>
      nx17237);
   ix2413 : and02 port map ( Y=>cache_data_in_2, A0=>mem_data_in(2), A1=>
      nx17237);
   ix2415 : and02 port map ( Y=>cache_data_in_3, A0=>mem_data_in(3), A1=>
      nx17239);
   ix2417 : and02 port map ( Y=>cache_data_in_4, A0=>mem_data_in(4), A1=>
      nx17239);
   ix2419 : and02 port map ( Y=>cache_data_in_5, A0=>mem_data_in(5), A1=>
      nx17239);
   ix2421 : and02 port map ( Y=>cache_data_in_6, A0=>mem_data_in(6), A1=>
      nx17239);
   ix2423 : and02 port map ( Y=>cache_data_in_7, A0=>mem_data_in(7), A1=>
      nx17239);
   ix2425 : and02 port map ( Y=>cache_data_in_8, A0=>mem_data_in(8), A1=>
      nx17239);
   ix2427 : and02 port map ( Y=>cache_data_in_9, A0=>mem_data_in(9), A1=>
      nx17239);
   ix2429 : and02 port map ( Y=>cache_data_in_10, A0=>mem_data_in(10), A1=>
      nx17039);
   ix2431 : and02 port map ( Y=>cache_data_in_11, A0=>mem_data_in(11), A1=>
      nx17039);
   ix2433 : and02 port map ( Y=>cache_data_in_12, A0=>mem_data_in(12), A1=>
      nx17039);
   ix2435 : and02 port map ( Y=>cache_data_in_13, A0=>mem_data_in(13), A1=>
      nx17039);
   ix2437 : and02 port map ( Y=>cache_data_in_14, A0=>mem_data_in(14), A1=>
      nx17083);
   ix2439 : and02 port map ( Y=>cache_data_in_15, A0=>mem_data_in(15), A1=>
      nx17083);
   ix15532 : nor02ii port map ( Y=>nx15531, A0=>nx16753, A1=>nx17111);
   ix2461 : mux21 port map ( Y=>max_height_3, A0=>nx15055, A1=>nx866, S0=>
      nx17115);
   ix2471 : mux21 port map ( Y=>max_height_4, A0=>nx15064, A1=>nx866, S0=>
      nx17115);
   ix13388 : mux21 port map ( Y=>nx13387, A0=>nx15541, A1=>nx15538, S0=>
      nx17129);
   ix13408 : mux21 port map ( Y=>nx13407, A0=>nx15550, A1=>nx15547, S0=>
      nx17129);
   ix13428 : mux21 port map ( Y=>nx13427, A0=>nx15556, A1=>nx15553, S0=>
      nx17129);
   ix13448 : mux21 port map ( Y=>nx13447, A0=>nx15562, A1=>nx15559, S0=>
      nx17131);
   ix13468 : mux21 port map ( Y=>nx13467, A0=>nx15568, A1=>nx15565, S0=>
      nx17131);
   ix13488 : mux21 port map ( Y=>nx13487, A0=>nx15574, A1=>nx15571, S0=>
      nx17131);
   ix13508 : mux21 port map ( Y=>nx13507, A0=>nx15580, A1=>nx15577, S0=>
      nx17131);
   ix13528 : mux21 port map ( Y=>nx13527, A0=>nx15586, A1=>nx15583, S0=>
      nx17131);
   ix13548 : mux21 port map ( Y=>nx13547, A0=>nx15592, A1=>nx15589, S0=>
      nx17131);
   ix13568 : mux21 port map ( Y=>nx13567, A0=>nx15598, A1=>nx15595, S0=>
      nx17131);
   ix13588 : mux21 port map ( Y=>nx13587, A0=>nx15604, A1=>nx15601, S0=>
      nx17133);
   ix13608 : mux21 port map ( Y=>nx13607, A0=>nx15610, A1=>nx15607, S0=>
      nx17133);
   ix13628 : mux21 port map ( Y=>nx13627, A0=>nx15616, A1=>nx15613, S0=>
      nx17133);
   ix13648 : mux21 port map ( Y=>nx13647, A0=>nx15622, A1=>nx15619, S0=>
      nx17133);
   ix13668 : mux21 port map ( Y=>nx13667, A0=>nx15628, A1=>nx15625, S0=>
      nx17133);
   ix13688 : mux21 port map ( Y=>nx13687, A0=>nx15634, A1=>nx15631, S0=>
      nx17133);
   ix4511 : nor02ii port map ( Y=>filter_data_out(0), A0=>nx17193, A1=>
      mem_data_in(0));
   ix4513 : nor02ii port map ( Y=>filter_data_out(1), A0=>nx17193, A1=>
      mem_data_in(1));
   ix4515 : nor02ii port map ( Y=>filter_data_out(2), A0=>nx17193, A1=>
      mem_data_in(2));
   ix4517 : nor02ii port map ( Y=>filter_data_out(3), A0=>nx17193, A1=>
      mem_data_in(3));
   ix4519 : nor02ii port map ( Y=>filter_data_out(4), A0=>nx17193, A1=>
      mem_data_in(4));
   ix4521 : nor02ii port map ( Y=>filter_data_out(5), A0=>nx17193, A1=>
      mem_data_in(5));
   ix4523 : nor02ii port map ( Y=>filter_data_out(6), A0=>nx17195, A1=>
      mem_data_in(6));
   ix4525 : nor02ii port map ( Y=>filter_data_out(7), A0=>nx17195, A1=>
      mem_data_in(7));
   ix4527 : nor02ii port map ( Y=>filter_data_out(8), A0=>nx17195, A1=>
      mem_data_in(8));
   ix4529 : nor02ii port map ( Y=>filter_data_out(9), A0=>nx17195, A1=>
      mem_data_in(9));
   ix4531 : nor02ii port map ( Y=>filter_data_out(10), A0=>nx17195, A1=>
      mem_data_in(10));
   ix4533 : nor02ii port map ( Y=>filter_data_out(11), A0=>nx17195, A1=>
      mem_data_in(11));
   ix4535 : nor02ii port map ( Y=>filter_data_out(12), A0=>nx17195, A1=>
      mem_data_in(12));
   ix4537 : nor02ii port map ( Y=>filter_data_out(13), A0=>nx16795, A1=>
      mem_data_in(13));
   ix4539 : nor02ii port map ( Y=>filter_data_out(14), A0=>nx16795, A1=>
      mem_data_in(14));
   ix4541 : nor02ii port map ( Y=>filter_data_out(15), A0=>nx16795, A1=>
      mem_data_in(15));
   ix4613 : and02 port map ( Y=>wind_col_in_0_0, A0=>nx17217, A1=>
      cache_data_out_0_0);
   ix4615 : and02 port map ( Y=>wind_col_in_0_1, A0=>nx17217, A1=>
      cache_data_out_0_1);
   ix4617 : and02 port map ( Y=>wind_col_in_0_2, A0=>nx17217, A1=>
      cache_data_out_0_2);
   ix4619 : and02 port map ( Y=>wind_col_in_0_3, A0=>nx17217, A1=>
      cache_data_out_0_3);
   ix4621 : and02 port map ( Y=>wind_col_in_0_4, A0=>nx17217, A1=>
      cache_data_out_0_4);
   ix4623 : and02 port map ( Y=>wind_col_in_0_5, A0=>nx17217, A1=>
      cache_data_out_0_5);
   ix4625 : and02 port map ( Y=>wind_col_in_0_6, A0=>nx17219, A1=>
      cache_data_out_0_6);
   ix4627 : and02 port map ( Y=>wind_col_in_0_7, A0=>nx17219, A1=>
      cache_data_out_0_7);
   ix4629 : and02 port map ( Y=>wind_col_in_0_8, A0=>nx17219, A1=>
      cache_data_out_0_8);
   ix4631 : and02 port map ( Y=>wind_col_in_0_9, A0=>nx17219, A1=>
      cache_data_out_0_9);
   ix4633 : and02 port map ( Y=>wind_col_in_0_10, A0=>nx17219, A1=>
      cache_data_out_0_10);
   ix4635 : and02 port map ( Y=>wind_col_in_0_11, A0=>nx17219, A1=>
      cache_data_out_0_11);
   ix4637 : and02 port map ( Y=>wind_col_in_0_12, A0=>nx17219, A1=>
      cache_data_out_0_12);
   ix4639 : and02 port map ( Y=>wind_col_in_0_13, A0=>nx17221, A1=>
      cache_data_out_0_13);
   ix4641 : and02 port map ( Y=>wind_col_in_0_14, A0=>nx17221, A1=>
      cache_data_out_0_14);
   ix4643 : and02 port map ( Y=>wind_col_in_0_15, A0=>nx17221, A1=>
      cache_data_out_0_15);
   ix4645 : and02 port map ( Y=>wind_col_in_1_0, A0=>nx17221, A1=>
      cache_data_out_1_0);
   ix4647 : and02 port map ( Y=>wind_col_in_1_1, A0=>nx17221, A1=>
      cache_data_out_1_1);
   ix4649 : and02 port map ( Y=>wind_col_in_1_2, A0=>nx17221, A1=>
      cache_data_out_1_2);
   ix4651 : and02 port map ( Y=>wind_col_in_1_3, A0=>nx17221, A1=>
      cache_data_out_1_3);
   ix4653 : and02 port map ( Y=>wind_col_in_1_4, A0=>nx17223, A1=>
      cache_data_out_1_4);
   ix4655 : and02 port map ( Y=>wind_col_in_1_5, A0=>nx17223, A1=>
      cache_data_out_1_5);
   ix4657 : and02 port map ( Y=>wind_col_in_1_6, A0=>nx17223, A1=>
      cache_data_out_1_6);
   ix4659 : and02 port map ( Y=>wind_col_in_1_7, A0=>nx17223, A1=>
      cache_data_out_1_7);
   ix4661 : and02 port map ( Y=>wind_col_in_1_8, A0=>nx17223, A1=>
      cache_data_out_1_8);
   ix4663 : and02 port map ( Y=>wind_col_in_1_9, A0=>nx17223, A1=>
      cache_data_out_1_9);
   ix4665 : and02 port map ( Y=>wind_col_in_1_10, A0=>nx17223, A1=>
      cache_data_out_1_10);
   ix4667 : and02 port map ( Y=>wind_col_in_1_11, A0=>nx17225, A1=>
      cache_data_out_1_11);
   ix4669 : and02 port map ( Y=>wind_col_in_1_12, A0=>nx17225, A1=>
      cache_data_out_1_12);
   ix4671 : and02 port map ( Y=>wind_col_in_1_13, A0=>nx17225, A1=>
      cache_data_out_1_13);
   ix4673 : and02 port map ( Y=>wind_col_in_1_14, A0=>nx17225, A1=>
      cache_data_out_1_14);
   ix4675 : and02 port map ( Y=>wind_col_in_1_15, A0=>nx17225, A1=>
      cache_data_out_1_15);
   ix4677 : and02 port map ( Y=>wind_col_in_2_0, A0=>nx17225, A1=>
      cache_data_out_2_0);
   ix4679 : and02 port map ( Y=>wind_col_in_2_1, A0=>nx17225, A1=>
      cache_data_out_2_1);
   ix4681 : and02 port map ( Y=>wind_col_in_2_2, A0=>nx17227, A1=>
      cache_data_out_2_2);
   ix4683 : and02 port map ( Y=>wind_col_in_2_3, A0=>nx17227, A1=>
      cache_data_out_2_3);
   ix4685 : and02 port map ( Y=>wind_col_in_2_4, A0=>nx17227, A1=>
      cache_data_out_2_4);
   ix4687 : and02 port map ( Y=>wind_col_in_2_5, A0=>nx17227, A1=>
      cache_data_out_2_5);
   ix4689 : and02 port map ( Y=>wind_col_in_2_6, A0=>nx17227, A1=>
      cache_data_out_2_6);
   ix4691 : and02 port map ( Y=>wind_col_in_2_7, A0=>nx17227, A1=>
      cache_data_out_2_7);
   ix4693 : and02 port map ( Y=>wind_col_in_2_8, A0=>nx17227, A1=>
      cache_data_out_2_8);
   ix4695 : and02 port map ( Y=>wind_col_in_2_9, A0=>nx17035, A1=>
      cache_data_out_2_9);
   ix4697 : and02 port map ( Y=>wind_col_in_2_10, A0=>nx17229, A1=>
      cache_data_out_2_10);
   ix4699 : and02 port map ( Y=>wind_col_in_2_11, A0=>nx17229, A1=>
      cache_data_out_2_11);
   ix4701 : and02 port map ( Y=>wind_col_in_2_12, A0=>nx17229, A1=>
      cache_data_out_2_12);
   ix4703 : and02 port map ( Y=>wind_col_in_2_13, A0=>nx17229, A1=>
      cache_data_out_2_13);
   ix4705 : and02 port map ( Y=>wind_col_in_2_14, A0=>nx17229, A1=>
      cache_data_out_2_14);
   ix4707 : and02 port map ( Y=>wind_col_in_2_15, A0=>nx17229, A1=>
      cache_data_out_2_15);
   ix4709 : and02 port map ( Y=>wind_col_in_3_0, A0=>nx17229, A1=>
      cache_data_out_3_0);
   ix4711 : and02 port map ( Y=>wind_col_in_3_1, A0=>nx17231, A1=>
      cache_data_out_3_1);
   ix4713 : and02 port map ( Y=>wind_col_in_3_2, A0=>nx17231, A1=>
      cache_data_out_3_2);
   ix4715 : and02 port map ( Y=>wind_col_in_3_3, A0=>nx17231, A1=>
      cache_data_out_3_3);
   ix4717 : and02 port map ( Y=>wind_col_in_3_4, A0=>nx17231, A1=>
      cache_data_out_3_4);
   ix4719 : and02 port map ( Y=>wind_col_in_3_5, A0=>nx17231, A1=>
      cache_data_out_3_5);
   ix4721 : and02 port map ( Y=>wind_col_in_3_6, A0=>nx17231, A1=>
      cache_data_out_3_6);
   ix4723 : and02 port map ( Y=>wind_col_in_3_7, A0=>nx17231, A1=>
      cache_data_out_3_7);
   ix4725 : and02 port map ( Y=>wind_col_in_3_8, A0=>nx17233, A1=>
      cache_data_out_3_8);
   ix4727 : and02 port map ( Y=>wind_col_in_3_9, A0=>nx17233, A1=>
      cache_data_out_3_9);
   ix4729 : and02 port map ( Y=>wind_col_in_3_10, A0=>nx17233, A1=>
      cache_data_out_3_10);
   ix4731 : and02 port map ( Y=>wind_col_in_3_11, A0=>nx17233, A1=>
      cache_data_out_3_11);
   ix4733 : and02 port map ( Y=>wind_col_in_3_12, A0=>nx17233, A1=>
      cache_data_out_3_12);
   ix4735 : and02 port map ( Y=>wind_col_in_3_13, A0=>nx17233, A1=>
      cache_data_out_3_13);
   ix4737 : and02 port map ( Y=>wind_col_in_3_14, A0=>nx17233, A1=>
      cache_data_out_3_14);
   ix4739 : and02 port map ( Y=>wind_col_in_3_15, A0=>nx17235, A1=>
      cache_data_out_3_15);
   ix4741 : and02 port map ( Y=>wind_col_in_4_0, A0=>nx17235, A1=>
      cache_data_out_4_0);
   ix4743 : and02 port map ( Y=>wind_col_in_4_1, A0=>nx17235, A1=>
      cache_data_out_4_1);
   ix4745 : and02 port map ( Y=>wind_col_in_4_2, A0=>nx17235, A1=>
      cache_data_out_4_2);
   ix4747 : and02 port map ( Y=>wind_col_in_4_3, A0=>nx17235, A1=>
      cache_data_out_4_3);
   ix4749 : and02 port map ( Y=>wind_col_in_4_4, A0=>nx17235, A1=>
      cache_data_out_4_4);
   ix4751 : and02 port map ( Y=>wind_col_in_4_5, A0=>nx17235, A1=>
      cache_data_out_4_5);
   ix4753 : and02 port map ( Y=>wind_col_in_4_6, A0=>nx17037, A1=>
      cache_data_out_4_6);
   ix4755 : and02 port map ( Y=>wind_col_in_4_7, A0=>nx17037, A1=>
      cache_data_out_4_7);
   ix4757 : and02 port map ( Y=>wind_col_in_4_8, A0=>nx17037, A1=>
      cache_data_out_4_8);
   ix4759 : and02 port map ( Y=>wind_col_in_4_9, A0=>nx17037, A1=>
      cache_data_out_4_9);
   ix4761 : and02 port map ( Y=>wind_col_in_4_10, A0=>nx17037, A1=>
      cache_data_out_4_10);
   ix4763 : and02 port map ( Y=>wind_col_in_4_11, A0=>nx17037, A1=>
      cache_data_out_4_11);
   ix4765 : and02 port map ( Y=>wind_col_in_4_12, A0=>nx17037, A1=>
      cache_data_out_4_12);
   ix4767 : and02 port map ( Y=>wind_col_in_4_13, A0=>nx2372, A1=>
      cache_data_out_4_13);
   ix4769 : and02 port map ( Y=>wind_col_in_4_14, A0=>nx2372, A1=>
      cache_data_out_4_14);
   ix4771 : and02 port map ( Y=>wind_col_in_4_15, A0=>nx2372, A1=>
      cache_data_out_4_15);
   ix2373 : or03 port map ( Y=>nx2372, A0=>nx14871, A1=>nx15075, A2=>nx15077
   );
   ix15740 : or02 port map ( Y=>nx15739, A0=>nx15075, A1=>
      ftc_cntrl_reg_out_11);
   ix15743 : and03 port map ( Y=>nx15742, A0=>nx16027, A1=>nx17155, A2=>
      nx17163);
   ix2519 : nand02 port map ( Y=>nx15803, A0=>nx17153, A1=>nx16913);
   ix1967 : nor02ii port map ( Y=>nx1966, A0=>nx17133, A1=>nx646);
   ix15751 : and04 port map ( Y=>nx15750, A0=>nx16795, A1=>nx17145, A2=>
      nx17065, A3=>nx17213);
   ix17064 : inv01 port map ( Y=>nx17065, A=>nx2568);
   ix15756 : and04 port map ( Y=>nx15755, A0=>nx17067, A1=>nx17201, A2=>
      nx17103, A3=>nx15297);
   ix17066 : inv01 port map ( Y=>nx17067, A=>current_state_5);
   ix1763 : nor02_2x port map ( Y=>nx1762, A0=>nx1742, A1=>nx15353);
   ix13738 : xor2 port map ( Y=>nx13737, A0=>addr1_data_0, A1=>nx17089);
   ix15767 : nand04 port map ( Y=>nx2572, A0=>nx17065, A1=>nx17213, A2=>
      nx15339, A3=>nx17099);
   ix15782 : nor02ii port map ( Y=>nx15781, A0=>new_size_squared_out_0, A1=>
      nx17805);
   ix15786 : nor02ii port map ( Y=>nx15785, A0=>layer_mem_size_out_0, A1=>
      nx17805);
   ix13708 : mux21_ni port map ( Y=>nx13707, A0=>mem_data_in(0), A1=>
      layer_mem_size_out_0, S0=>nx17103);
   ix15792 : nor02ii port map ( Y=>nx15791, A0=>nx17069, A1=>nx16945);
   ix13728 : mux21_ni port map ( Y=>nx13727, A0=>nx17808, A1=>
      bias_offset_data_out_0, S0=>nx17163);
   ix15806 : or02 port map ( Y=>nx15805, A0=>nx17159, A1=>nx15350);
   ix13748 : xor2 port map ( Y=>nx13747, A0=>img_addr_offset_0, A1=>nx17085
   );
   ix2527 : and02 port map ( Y=>nx2526, A0=>write_offset_data_out_0, A1=>
      nx17159);
   ix13798 : mux21 port map ( Y=>nx13797, A0=>nx15815, A1=>nx15818, S0=>
      nx17091);
   ix13768 : mux21_ni port map ( Y=>nx13767, A0=>mem_data_in(1), A1=>
      layer_mem_size_out_1, S0=>nx17103);
   ix13758 : mux21 port map ( Y=>nx13757, A0=>nx15855, A1=>nx15851, S0=>
      nx17085);
   ix15861 : xnor2 port map ( Y=>nx15860, A0=>nx15864, A1=>nx17811);
   ix13788 : mux21 port map ( Y=>nx13787, A0=>nx14765, A1=>nx15864, S0=>
      nx17163);
   ix13848 : mux21_ni port map ( Y=>nx13847, A0=>addr1_data_2, A1=>nx2822, 
      S0=>nx17091);
   ix2823 : xor2 port map ( Y=>nx2822, A0=>nx15870, A1=>nx15821);
   ix15879 : xnor2 port map ( Y=>nx15878, A0=>nx17169, A1=>nx15364);
   ix13818 : mux21_ni port map ( Y=>nx13817, A0=>mem_data_in(2), A1=>
      layer_mem_size_out_2, S0=>nx17103);
   ix15906 : xnor2 port map ( Y=>nx15905, A0=>nx17171, A1=>nx14756);
   ix13838 : mux21_ni port map ( Y=>nx13837, A0=>img_addr_offset_2, A1=>
      nx2768, S0=>nx17085);
   ix2769 : xor2 port map ( Y=>nx2768, A0=>nx15908, A1=>nx15857);
   ix15914 : nor02ii port map ( Y=>nx15913, A0=>img_addr_offset_0, A1=>
      nx15855);
   ix13808 : mux21 port map ( Y=>nx13807, A0=>nx14759, A1=>nx15924, S0=>
      nx17163);
   ix13898 : mux21_ni port map ( Y=>nx13897, A0=>addr1_data_3, A1=>nx2954, 
      S0=>nx17091);
   ix2955 : xor2 port map ( Y=>nx2954, A0=>nx15927, A1=>nx15932);
   ix15952 : xor2 port map ( Y=>nx15951, A0=>layer_mem_size_out_3, A1=>
      nx17816);
   ix13868 : mux21_ni port map ( Y=>nx13867, A0=>mem_data_in(3), A1=>
      layer_mem_size_out_3, S0=>nx17103);
   ix13888 : mux21_ni port map ( Y=>nx13887, A0=>img_addr_offset_3, A1=>
      nx2900, S0=>nx17085);
   ix2901 : xor2 port map ( Y=>nx2900, A0=>nx15963, A1=>nx15968);
   ix15975 : xor2 port map ( Y=>nx15974, A0=>bias_offset_data_out_3, A1=>
      nx17816);
   ix13858 : mux21_ni port map ( Y=>nx13857, A0=>nx78, A1=>
      bias_offset_data_out_3, S0=>nx17163);
   ix79 : xor2 port map ( Y=>nx78, A0=>nx14751, A1=>nx14774);
   ix13948 : mux21_ni port map ( Y=>nx13947, A0=>addr1_data_4, A1=>nx3090, 
      S0=>nx17091);
   ix3085 : nor02ii port map ( Y=>nx3084, A0=>nx15991, A1=>addr1_data_4);
   ix13938 : mux21_ni port map ( Y=>nx13937, A0=>nx104, A1=>
      bias_offset_data_out_4, S0=>nx17163);
   ix13908 : mux21_ni port map ( Y=>nx13907, A0=>mem_data_in(4), A1=>
      layer_mem_size_out_4, S0=>nx17105);
   ix16034 : xnor2 port map ( Y=>nx16033, A0=>nx17175, A1=>nx14741);
   ix16037 : nor02ii port map ( Y=>nx16036, A0=>nx17665, A1=>nx17175);
   ix13928 : mux21_ni port map ( Y=>nx13927, A0=>img_addr_offset_4, A1=>
      nx3044, S0=>nx17085);
   ix3039 : nor02ii port map ( Y=>nx3038, A0=>nx16045, A1=>img_addr_offset_4
   );
   ix2909 : nor02ii port map ( Y=>nx2908, A0=>nx15961, A1=>img_addr_offset_3
   );
   ix16052 : nor02ii port map ( Y=>nx16051, A0=>nx2908, A1=>nx16047);
   ix16058 : xnor2 port map ( Y=>nx16057, A0=>nx16061, A1=>nx17820);
   ix13988 : mux21 port map ( Y=>nx13987, A0=>nx14738, A1=>nx16061, S0=>
      nx17165);
   ix16069 : xor2 port map ( Y=>nx16068, A0=>new_size_squared_out_5, A1=>
      nx17820);
   ix16074 : xor2 port map ( Y=>nx16073, A0=>layer_mem_size_out_5, A1=>
      nx17820);
   ix13958 : mux21_ni port map ( Y=>nx13957, A0=>mem_data_in(5), A1=>
      layer_mem_size_out_5, S0=>nx17105);
   ix13998 : mux21 port map ( Y=>nx13997, A0=>nx16080, A1=>nx16083, S0=>
      nx17091);
   ix16098 : and02 port map ( Y=>nx16097, A0=>nx17821, A1=>nx17664);
   ix16103 : and02 port map ( Y=>nx16102, A0=>nx16110, A1=>nx16051);
   ix13978 : mux21 port map ( Y=>nx13977, A0=>nx16110, A1=>nx16106, S0=>
      nx17085);
   ix3171 : nor02ii port map ( Y=>nx3170, A0=>nx16051, A1=>img_addr_offset_5
   );
   ix14038 : mux21_ni port map ( Y=>nx14037, A0=>nx150, A1=>
      bias_offset_data_out_6, S0=>nx17165);
   ix14008 : mux21_ni port map ( Y=>nx14007, A0=>mem_data_in(6), A1=>
      layer_mem_size_out_6, S0=>nx17105);
   ix14048 : mux21_ni port map ( Y=>nx14047, A0=>addr1_data_6, A1=>nx3346, 
      S0=>nx17091);
   ix3347 : xor2 port map ( Y=>nx3346, A0=>nx16146, A1=>nx16086);
   ix16156 : xnor2 port map ( Y=>nx16155, A0=>nx17179, A1=>nx14726);
   ix16159 : nor02ii port map ( Y=>nx16158, A0=>nx17660, A1=>nx17179);
   ix14028 : mux21_ni port map ( Y=>nx14027, A0=>img_addr_offset_6, A1=>
      nx3300, S0=>nx17085);
   ix3295 : nor02ii port map ( Y=>nx3294, A0=>nx16108, A1=>img_addr_offset_6
   );
   ix16170 : nor02ii port map ( Y=>nx16169, A0=>nx3170, A1=>nx16166);
   ix16176 : xnor2 port map ( Y=>nx16175, A0=>nx16179, A1=>nx16196);
   ix14088 : mux21 port map ( Y=>nx14087, A0=>nx14723, A1=>nx16179, S0=>
      nx17165);
   ix16187 : xor2 port map ( Y=>nx16186, A0=>new_size_squared_out_7, A1=>
      nx16196);
   ix16192 : xor2 port map ( Y=>nx16191, A0=>layer_mem_size_out_7, A1=>
      nx16196);
   ix14058 : mux21_ni port map ( Y=>nx14057, A0=>mem_data_in(7), A1=>
      layer_mem_size_out_7, S0=>nx17105);
   ix14098 : mux21 port map ( Y=>nx14097, A0=>nx16198, A1=>nx16201, S0=>
      nx17091);
   ix3341 : nor02ii port map ( Y=>nx3340, A0=>nx16086, A1=>addr1_data_6);
   ix16214 : xnor2 port map ( Y=>nx16213, A0=>nx16196, A1=>nx14712);
   ix16217 : and02 port map ( Y=>nx16216, A0=>nx16196, A1=>nx16218);
   ix16222 : and02 port map ( Y=>nx16221, A0=>nx16229, A1=>nx16169);
   ix14078 : mux21 port map ( Y=>nx14077, A0=>nx16229, A1=>nx16225, S0=>
      nx17087);
   ix3427 : nor02ii port map ( Y=>nx3426, A0=>nx16169, A1=>img_addr_offset_7
   );
   ix14138 : mux21_ni port map ( Y=>nx14137, A0=>nx200, A1=>
      bias_offset_data_out_8, S0=>nx17165);
   ix14108 : mux21_ni port map ( Y=>nx14107, A0=>mem_data_in(8), A1=>
      layer_mem_size_out_8, S0=>nx17105);
   ix14148 : mux21_ni port map ( Y=>nx14147, A0=>addr1_data_8, A1=>nx3602, 
      S0=>nx17093);
   ix3603 : xor2 port map ( Y=>nx3602, A0=>nx16265, A1=>nx16205);
   ix16275 : xnor2 port map ( Y=>nx16274, A0=>nx17183, A1=>nx14702);
   ix16278 : nor02ii port map ( Y=>nx16277, A0=>nx3436, A1=>nx17183);
   ix16281 : nor02ii port map ( Y=>nx16280, A0=>nx3426, A1=>nx16285);
   ix14128 : mux21_ni port map ( Y=>nx14127, A0=>img_addr_offset_8, A1=>
      nx3546, S0=>nx17087);
   ix3541 : nor02ii port map ( Y=>nx3540, A0=>nx16227, A1=>img_addr_offset_8
   );
   ix16294 : xnor2 port map ( Y=>nx16293, A0=>nx16297, A1=>nx16314);
   ix14188 : mux21 port map ( Y=>nx14187, A0=>nx14699, A1=>nx16297, S0=>
      nx17165);
   ix16305 : xor2 port map ( Y=>nx16304, A0=>new_size_squared_out_9, A1=>
      nx16314);
   ix16310 : xor2 port map ( Y=>nx16309, A0=>layer_mem_size_out_9, A1=>
      nx16314);
   ix14158 : mux21_ni port map ( Y=>nx14157, A0=>mem_data_in(9), A1=>
      layer_mem_size_out_9, S0=>nx17105);
   ix14198 : mux21 port map ( Y=>nx14197, A0=>nx16316, A1=>nx16319, S0=>
      nx17093);
   ix3597 : nor02ii port map ( Y=>nx3596, A0=>nx16205, A1=>addr1_data_8);
   ix16332 : xnor2 port map ( Y=>nx16331, A0=>nx16314, A1=>nx14776);
   ix16335 : and02 port map ( Y=>nx16334, A0=>nx16314, A1=>nx16336);
   ix3693 : nor02ii port map ( Y=>nx3692, A0=>nx16336, A1=>
      write_base_data_out_9);
   ix16340 : and02 port map ( Y=>nx16339, A0=>nx16347, A1=>nx16349);
   ix14178 : mux21 port map ( Y=>nx14177, A0=>nx16347, A1=>nx16343, S0=>
      nx17087);
   ix3683 : nor02ii port map ( Y=>nx3682, A0=>nx16349, A1=>img_addr_offset_9
   );
   ix14238 : mux21_ni port map ( Y=>nx14237, A0=>nx246, A1=>
      bias_offset_data_out_10, S0=>nx17165);
   ix14208 : mux21_ni port map ( Y=>nx14207, A0=>mem_data_in(10), A1=>
      layer_mem_size_out_10, S0=>nx17105);
   ix14248 : mux21_ni port map ( Y=>nx14247, A0=>addr1_data_10, A1=>nx3858, 
      S0=>nx17093);
   ix3859 : xor2 port map ( Y=>nx3858, A0=>nx16385, A1=>nx16323);
   ix16395 : xnor2 port map ( Y=>nx16394, A0=>nx17187, A1=>nx14689);
   ix16398 : nor02ii port map ( Y=>nx16397, A0=>nx17828, A1=>nx17187);
   ix16401 : nor02ii port map ( Y=>nx16400, A0=>nx3682, A1=>nx16405);
   ix14228 : mux21_ni port map ( Y=>nx14227, A0=>img_addr_offset_10, A1=>
      nx3802, S0=>nx17087);
   ix3797 : nor02ii port map ( Y=>nx3796, A0=>nx16345, A1=>
      img_addr_offset_10);
   ix16414 : xnor2 port map ( Y=>nx16413, A0=>nx16417, A1=>nx17832);
   ix14288 : mux21 port map ( Y=>nx14287, A0=>nx14686, A1=>nx16417, S0=>
      nx17165);
   ix14258 : mux21_ni port map ( Y=>nx14257, A0=>mem_data_in(11), A1=>
      layer_mem_size_out_11, S0=>nx17107);
   ix14298 : mux21 port map ( Y=>nx14297, A0=>nx16436, A1=>nx16439, S0=>
      nx17093);
   ix3853 : nor02ii port map ( Y=>nx3852, A0=>nx16323, A1=>addr1_data_10);
   ix16455 : and02 port map ( Y=>nx16454, A0=>nx17832, A1=>nx16456);
   ix16460 : xor2 port map ( Y=>nx16459, A0=>nx16467, A1=>nx16469);
   ix14278 : mux21 port map ( Y=>nx14277, A0=>nx16467, A1=>nx16463, S0=>
      nx17087);
   ix14338 : mux21_ni port map ( Y=>nx14337, A0=>nx294, A1=>
      bias_offset_data_out_12, S0=>nx17167);
   ix14308 : mux21_ni port map ( Y=>nx14307, A0=>mem_data_in(12), A1=>
      layer_mem_size_out_12, S0=>nx17107);
   ix14348 : mux21_ni port map ( Y=>nx14347, A0=>addr1_data_12, A1=>nx4114, 
      S0=>nx17093);
   ix4115 : xor2 port map ( Y=>nx4114, A0=>nx16504, A1=>nx16443);
   ix16514 : xnor2 port map ( Y=>nx16513, A0=>nx17191, A1=>nx14676);
   ix16517 : nor02ii port map ( Y=>nx16516, A0=>nx3926, A1=>nx17191);
   ix14328 : mux21_ni port map ( Y=>nx14327, A0=>img_addr_offset_12, A1=>
      nx4068, S0=>nx17087);
   ix4063 : nor02ii port map ( Y=>nx4062, A0=>nx16465, A1=>
      img_addr_offset_12);
   ix16529 : nor02ii port map ( Y=>nx16528, A0=>nx3946, A1=>nx16524);
   ix14388 : mux21 port map ( Y=>nx14387, A0=>nx14673, A1=>nx16538, S0=>
      nx17167);
   ix16551 : xor2 port map ( Y=>nx16550, A0=>layer_mem_size_out_13, A1=>
      nx17836);
   ix14358 : mux21_ni port map ( Y=>nx14357, A0=>mem_data_in(13), A1=>
      layer_mem_size_out_13, S0=>nx17107);
   ix14398 : mux21 port map ( Y=>nx14397, A0=>nx16557, A1=>nx16560, S0=>
      nx17093);
   ix4109 : nor02ii port map ( Y=>nx4108, A0=>nx16443, A1=>addr1_data_12);
   ix16581 : and02 port map ( Y=>nx16580, A0=>nx16588, A1=>nx16528);
   ix14378 : mux21 port map ( Y=>nx14377, A0=>nx16588, A1=>nx16584, S0=>
      nx17087);
   ix4195 : nor02ii port map ( Y=>nx4194, A0=>nx16528, A1=>
      img_addr_offset_13);
   ix14438 : mux21_ni port map ( Y=>nx14437, A0=>nx340, A1=>
      bias_offset_data_out_14, S0=>nx17167);
   ix341 : xor2 port map ( Y=>nx340, A0=>nx14663, A1=>nx14669);
   ix14408 : mux21_ni port map ( Y=>nx14407, A0=>mem_data_in(14), A1=>
      layer_mem_size_out_14, S0=>nx17107);
   ix14448 : mux21_ni port map ( Y=>nx14447, A0=>addr1_data_14, A1=>nx4370, 
      S0=>nx17093);
   ix4371 : xor2 port map ( Y=>nx4370, A0=>nx16624, A1=>nx16564);
   ix14428 : mux21_ni port map ( Y=>nx14427, A0=>img_addr_offset_14, A1=>
      nx4314, S0=>nx2406);
   ix4315 : xor2 port map ( Y=>nx4314, A0=>nx16635, A1=>nx16586);
   ix16643 : xnor2 port map ( Y=>nx16642, A0=>nx17838, A1=>nx14663);
   ix14498 : mux21 port map ( Y=>nx14497, A0=>nx16650, A1=>nx16647, S0=>
      nx17095);
   ix16648 : xor2 port map ( Y=>nx16647, A0=>nx16650, A1=>nx4364);
   ix4365 : nor02ii port map ( Y=>nx4364, A0=>nx16564, A1=>addr1_data_14);
   ix4429 : xor2 port map ( Y=>nx4428, A0=>layer_mem_size_out_15, A1=>
      write_base_data_out_15);
   ix14468 : mux21_ni port map ( Y=>nx14467, A0=>mem_data_in(15), A1=>
      layer_mem_size_out_15, S0=>nx17107);
   ix14488 : mux21 port map ( Y=>nx14487, A0=>nx14660, A1=>nx16677, S0=>
      nx17167);
   ix16690 : xor2 port map ( Y=>nx16689, A0=>nx16696, A1=>nx16636);
   ix14458 : mux21 port map ( Y=>nx14457, A0=>nx16696, A1=>nx16693, S0=>
      nx2406);
   ix16694 : xor2 port map ( Y=>nx16693, A0=>nx16696, A1=>nx4308);
   ix4309 : nor02ii port map ( Y=>nx4308, A0=>nx16586, A1=>
      img_addr_offset_14);
   ix16956 : and02 port map ( Y=>nx16957, A0=>nx14597, A1=>nx14722);
   ix16958 : and02 port map ( Y=>nx16959, A0=>nx14597, A1=>nx14722);
   ix17068 : inv01 port map ( Y=>nx17069, A=>nx16947);
   ix17070 : buf02 port map ( Y=>nx17071, A=>nx12265);
   ix17072 : buf02 port map ( Y=>nx17073, A=>nx12265);
   ix17074 : inv02 port map ( Y=>nx17075, A=>nx16963);
   ix17076 : inv02 port map ( Y=>nx17077, A=>nx16963);
   ix17078 : inv02 port map ( Y=>nx17079, A=>nx16963);
   ix17080 : inv02 port map ( Y=>nx17081, A=>nx16963);
   ix17082 : inv02 port map ( Y=>nx17083, A=>nx17155);
   ix17084 : inv02 port map ( Y=>nx17085, A=>nx17155);
   ix17086 : inv02 port map ( Y=>nx17087, A=>nx17155);
   ix17088 : inv02 port map ( Y=>nx17089, A=>nx17009);
   ix17090 : inv02 port map ( Y=>nx17091, A=>nx17009);
   ix17092 : inv02 port map ( Y=>nx17093, A=>nx17009);
   ix17094 : inv02 port map ( Y=>nx17095, A=>nx17009);
   ix17096 : buf02 port map ( Y=>nx17097, A=>nx14508);
   ix17098 : buf02 port map ( Y=>nx17099, A=>nx14508);
   ix17100 : inv01 port map ( Y=>nx17101, A=>nx14577);
   ix17102 : inv02 port map ( Y=>nx17103, A=>nx17101);
   ix17104 : inv02 port map ( Y=>nx17105, A=>nx17101);
   ix17106 : inv02 port map ( Y=>nx17107, A=>nx17101);
   ix17108 : inv02 port map ( Y=>nx17109, A=>nx16819);
   ix17110 : inv02 port map ( Y=>nx17111, A=>nx16819);
   ix17112 : inv02 port map ( Y=>nx17113, A=>nx16803);
   ix17114 : inv02 port map ( Y=>nx17115, A=>nx16803);
   ix17116 : inv02 port map ( Y=>nx17117, A=>nx862);
   ix17118 : inv02 port map ( Y=>nx17119, A=>nx17245);
   ix17120 : inv02 port map ( Y=>nx17121, A=>nx17245);
   ix17122 : inv02 port map ( Y=>nx17123, A=>nx12253);
   ix17124 : inv02 port map ( Y=>nx17125, A=>nx12253);
   ix17126 : inv02 port map ( Y=>nx17127, A=>nx12253);
   ix17128 : inv02 port map ( Y=>nx17129, A=>nx16891);
   ix17130 : inv02 port map ( Y=>nx17131, A=>nx16891);
   ix17132 : inv02 port map ( Y=>nx17133, A=>nx16891);
   ix17134 : inv02 port map ( Y=>nx17135, A=>nx16837);
   ix17136 : inv02 port map ( Y=>nx17137, A=>nx16837);
   ix17138 : inv02 port map ( Y=>nx17139, A=>argmax_ready_EXMPLR);
   ix17140 : inv02 port map ( Y=>nx17141, A=>argmax_ready_EXMPLR);
   ix17142 : inv02 port map ( Y=>nx17143, A=>argmax_ready_EXMPLR);
   ix17144 : inv02 port map ( Y=>nx17145, A=>argmax_ready_EXMPLR);
   ix17146 : inv01 port map ( Y=>nx17147, A=>nx15399);
   ix17148 : inv02 port map ( Y=>nx17149, A=>nx17147);
   ix17150 : inv02 port map ( Y=>nx17151, A=>nx17147);
   ix17152 : inv02 port map ( Y=>nx17153, A=>nx17147);
   ix17154 : inv02 port map ( Y=>nx17155, A=>nx2406);
   ix17158 : inv01 port map ( Y=>nx17159, A=>nx16919);
   ix17160 : inv01 port map ( Y=>nx17161, A=>nx15803);
   ix17162 : inv02 port map ( Y=>nx17163, A=>nx17161);
   ix17164 : inv02 port map ( Y=>nx17165, A=>nx17161);
   ix17166 : inv02 port map ( Y=>nx17167, A=>nx17161);
   ix17170 : inv02 port map ( Y=>nx17171, A=>nx17814);
   ix17174 : inv02 port map ( Y=>nx17175, A=>nx17818);
   ix17178 : inv02 port map ( Y=>nx17179, A=>nx17822);
   ix17182 : inv02 port map ( Y=>nx17183, A=>nx17824);
   ix17186 : inv02 port map ( Y=>nx17187, A=>nx17830);
   ix17190 : inv02 port map ( Y=>nx17191, A=>nx17834);
   ix17192 : inv01 port map ( Y=>nx17193, A=>filter_ready_out_EXMPLR);
   ix17194 : inv01 port map ( Y=>nx17195, A=>filter_ready_out_EXMPLR);
   ix17196 : inv02 port map ( Y=>nx17197, A=>current_state_6);
   ix17198 : inv02 port map ( Y=>nx17199, A=>current_state_6);
   ix17200 : inv02 port map ( Y=>nx17201, A=>current_state_6);
   ix17202 : inv02 port map ( Y=>nx17203, A=>nx8);
   ix17204 : inv02 port map ( Y=>nx17205, A=>nx8);
   ix17206 : inv01 port map ( Y=>nx17207, A=>nx16905);
   ix17208 : inv02 port map ( Y=>nx17209, A=>nx17207);
   ix17210 : inv02 port map ( Y=>nx17211, A=>nx17207);
   ix17212 : inv02 port map ( Y=>nx17213, A=>nx17207);
   ix17216 : inv01 port map ( Y=>nx17217, A=>nx17247);
   ix17218 : inv01 port map ( Y=>nx17219, A=>nx17247);
   ix17220 : inv01 port map ( Y=>nx17221, A=>nx17247);
   ix17222 : inv01 port map ( Y=>nx17223, A=>nx17247);
   ix17224 : inv01 port map ( Y=>nx17225, A=>nx17247);
   ix17226 : inv01 port map ( Y=>nx17227, A=>nx15656);
   ix17228 : inv01 port map ( Y=>nx17229, A=>nx15656);
   ix17230 : inv01 port map ( Y=>nx17231, A=>nx15656);
   ix17232 : inv01 port map ( Y=>nx17233, A=>nx15656);
   ix17234 : inv01 port map ( Y=>nx17235, A=>nx15656);
   ix17236 : inv02 port map ( Y=>nx17237, A=>nx17155);
   ix17238 : inv02 port map ( Y=>nx17239, A=>nx17155);
   ix17244 : inv01 port map ( Y=>nx17245, A=>nx17117);
   ix17246 : inv01 port map ( Y=>nx17247, A=>nx2372);
   ix17841 : nor03_2x port map ( Y=>nx17390, A0=>nx15836, A1=>nx17511, A2=>
      nx17805);
   reg_nx15886 : aoi21 port map ( Y=>nx15886, A0=>write_base_data_out_1, A1
      =>new_size_squared_out_1, B0=>nx17390);
   reg_nx15889 : oai22 port map ( Y=>nx15889, A0=>nx17510, A1=>nx17814, B0=>
      nx17169, B1=>nx14854);
   ix17842 : nor02ii port map ( Y=>nx17391, A0=>nx16382, A1=>nx17830);
   ix17843 : nor02ii port map ( Y=>nx17392, A0=>nx17830, A1=>nx16382);
   ix17844 : inv02 port map ( Y=>nx17393, A=>nx16501);
   ix17845 : nor02_2x port map ( Y=>nx17394, A0=>nx17393, A1=>nx17834);
   ix17846 : inv02 port map ( Y=>nx17395, A=>write_base_data_out_11);
   ix17847 : inv02 port map ( Y=>nx17396, A=>layer_mem_size_out_11);
   ix17848 : and02 port map ( Y=>nx17397, A0=>write_base_data_out_11, A1=>
      layer_mem_size_out_11);
   ix17849 : nor02_2x port map ( Y=>nx17398, A0=>nx17393, A1=>nx17397);
   ix17850 : and02 port map ( Y=>nx17399, A0=>nx17838, A1=>nx16621);
   ix17851 : inv02 port map ( Y=>nx17400, A=>write_base_data_out_13);
   ix17852 : inv02 port map ( Y=>nx17401, A=>layer_mem_size_out_13);
   reg_nx4420 : oai332 port map ( Y=>nx4420, A0=>nx17559, A1=>nx17399, A2=>
      nx16550, B0=>nx17399, B1=>nx17400, B2=>nx17401, C0=>nx17838, C1=>
      nx16621);
   ix17853 : oai21 port map ( Y=>nx17402, A0=>nx17400, A1=>nx17401, B0=>
      nx16550);
   ix17854 : nor02_2x port map ( Y=>nx17403, A0=>nx17838, A1=>nx16621);
   ix17855 : inv02 port map ( Y=>nx17404, A=>nx16429);
   reg_nx16494 : oai32 port map ( Y=>nx16494, A0=>nx17397, A1=>nx17391, A2=>
      nx17501, B0=>nx17404, B1=>nx17397);
   reg_nx16497 : oai22 port map ( Y=>nx16497, A0=>nx17189, A1=>nx16501, B0=>
      nx17393, B1=>nx17834);
   ix17856 : inv02 port map ( Y=>nx17405, A=>nx16382);
   reg_nx16378 : oai22 port map ( Y=>nx16378, A0=>nx17405, A1=>nx17830, B0=>
      nx17185, B1=>nx16382);
   ix17857 : nor02_2x port map ( Y=>nx17406, A0=>nx17400, A1=>nx17401);
   reg_nx16614 : oai21 port map ( Y=>nx16614, A0=>nx4154, A1=>nx17406, B0=>
      nx17402);
   ix17858 : aoi21 port map ( Y=>nx17407, A0=>nx17839, A1=>nx16621, B0=>
      nx17403);
   ix17859 : ao21 port map ( Y=>nx17408, A0=>nx17839, A1=>nx16621, B0=>
      nx17403);
   ix17860 : inv01 port map ( Y=>nx17409, A=>nx17400);
   ix17861 : inv01 port map ( Y=>nx17410, A=>nx17401);
   ix17862 : aoi21 port map ( Y=>nx17411, A0=>nx17409, A1=>nx17410, B0=>
      nx4154);
   ix17863 : nor02ii port map ( Y=>nx17412, A0=>nx17411, A1=>nx17402);
   ix17864 : aoi22 port map ( Y=>nx17413, A0=>nx16614, A1=>nx17407, B0=>
      nx17408, B1=>nx17412);
   ix17865 : inv02 port map ( Y=>nx17414, A=>write_base_data_out_13);
   ix17866 : inv02 port map ( Y=>nx17415, A=>new_size_squared_out_13);
   ix17867 : oai21 port map ( Y=>nx17416, A0=>nx17414, A1=>nx17415, B0=>
      nx16545);
   ix17868 : inv02 port map ( Y=>nx17417, A=>nx14801);
   ix17869 : nor02_2x port map ( Y=>nx17418, A0=>nx17417, A1=>nx17834);
   ix17870 : inv01 port map ( Y=>nx17419, A=>nx17839);
   ix17871 : inv02 port map ( Y=>nx17420, A=>nx14791);
   ix17872 : aoi22 port map ( Y=>nx17421, A0=>nx17839, A1=>nx14791, B0=>
      nx17419, B1=>nx17420);
   ix17873 : oai22 port map ( Y=>nx17422, A0=>nx17420, A1=>nx17839, B0=>
      nx17419, B1=>nx14791);
   reg_nx14417 : oai222 port map ( Y=>nx14417, A0=>nx17215, A1=>nx17413, B0
      =>nx17840, B1=>nx16925, C0=>nx16951, C1=>nx16605);
   reg_nx16610 : oai22 port map ( Y=>nx16610, A0=>nx17419, A1=>nx17420, B0=>
      nx17840, B1=>nx14791);
   reg_nx16490 : oai22 port map ( Y=>nx16490, A0=>nx17417, A1=>nx17834, B0=>
      nx17189, B1=>nx14801);
   ix17874 : inv02 port map ( Y=>nx17423, A=>nx14812);
   ix17875 : nor02_2x port map ( Y=>nx17424, A0=>nx17423, A1=>nx17830);
   ix17876 : nor02_2x port map ( Y=>nx17425, A0=>nx17424, A1=>nx16424);
   ix17877 : nor02ii port map ( Y=>nx17426, A0=>nx17418, A1=>nx17416);
   ix17878 : oai22 port map ( Y=>nx17427, A0=>nx17189, A1=>nx14801, B0=>
      nx17414, B1=>nx17415);
   ix17879 : inv02 port map ( Y=>nx17428, A=>write_base_data_out_11);
   ix17880 : inv02 port map ( Y=>nx17429, A=>new_size_squared_out_11);
   ix17881 : oai32 port map ( Y=>nx17430, A0=>nx16424, A1=>nx17185, A2=>
      nx14812, B0=>nx17428, B1=>nx17429);
   ix17882 : oai21 port map ( Y=>nx17431, A0=>nx17428, A1=>nx17429, B0=>
      nx16424);
   reg_nx16371 : oai22 port map ( Y=>nx16371, A0=>nx17423, A1=>nx17830, B0=>
      nx17185, B1=>nx14812);
   ix17883 : nand02_2x port map ( Y=>nx17432, A0=>nx15900, A1=>nx17169);
   ix17884 : inv01 port map ( Y=>nx17433, A=>nx17811);
   ix17885 : nand02_2x port map ( Y=>nx17434, A0=>layer_mem_size_out_1, A1=>
      nx17433);
   ix17886 : inv02 port map ( Y=>nx17435, A=>write_base_data_out_1);
   ix17887 : nand03_2x port map ( Y=>nx17436, A0=>layer_mem_size_out_0, A1=>
      nx16919, A2=>nx17433);
   ix17888 : inv02 port map ( Y=>nx17437, A=>layer_mem_size_out_1);
   ix17889 : nor02ii port map ( Y=>nx17438, A0=>nx15900, A1=>nx17814);
   reg_nx15893 : inv01 port map ( Y=>nx15893, A=>nx17529);
   ix17890 : inv02 port map ( Y=>nx17439, A=>nx15900);
   reg_nx15896 : oai22 port map ( Y=>nx15896, A0=>nx17439, A1=>nx17814, B0=>
      nx17169, B1=>nx15900);
   reg_nx15842 : oai22 port map ( Y=>nx15842, A0=>nx17433, A1=>
      layer_mem_size_out_1, B0=>nx17437, B1=>nx17811);
   ix17891 : or02 port map ( Y=>nx17440, A0=>nx17840, A1=>nx16602);
   ix17892 : inv02 port map ( Y=>nx17441, A=>nx16677);
   ix17893 : inv02 port map ( Y=>nx17442, A=>write_base_data_out_15);
   ix17894 : aoi22 port map ( Y=>nx17443, A0=>nx16677, A1=>
      write_base_data_out_15, B0=>nx17441, B1=>nx17442);
   ix17895 : and02 port map ( Y=>nx17444, A0=>nx17840, A1=>nx16602);
   ix17896 : nor02_2x port map ( Y=>nx17445, A0=>nx18301, A1=>nx17444);
   ix17897 : nor03_2x port map ( Y=>nx17446, A0=>nx18301, A1=>nx17840, A2=>
      nx16602);
   ix17898 : ao21 port map ( Y=>nx17447, A0=>nx18301, A1=>nx17444, B0=>
      nx17446);
   ix17899 : inv02 port map ( Y=>nx17448, A=>nx16686);
   ix17900 : inv02 port map ( Y=>nx17449, A=>nx14782);
   ix17901 : inv02 port map ( Y=>nx17450, A=>nx16661);
   ix17902 : oai22 port map ( Y=>nx17451, A0=>nx17449, A1=>nx16661, B0=>
      nx17450, B1=>nx14782);
   ix17903 : inv02 port map ( Y=>nx17452, A=>write_base_data_out_14);
   ix17904 : inv02 port map ( Y=>nx17453, A=>write_offset_data_out_14);
   ix17905 : oai21 port map ( Y=>nx17454, A0=>nx17452, A1=>nx17453, B0=>
      nx16642);
   ix17906 : and02 port map ( Y=>nx17455, A0=>nx14780, A1=>nx17836);
   ix17907 : aoi22 port map ( Y=>nx17456, A0=>nx16661, A1=>nx14782, B0=>
      nx17450, B1=>nx17449);
   ix17908 : nor02_2x port map ( Y=>nx17457, A0=>nx17542, A1=>nx17456);
   ix17909 : inv02 port map ( Y=>nx17458, A=>addr1_data_15);
   ix17910 : inv02 port map ( Y=>nx17459, A=>nx17089);
   ix17911 : and02 port map ( Y=>nx17460, A0=>nx17145, A1=>nx15758);
   ix17912 : inv02 port map ( Y=>nx17461, A=>write_base_data_out_13);
   ix17913 : nor03_2x port map ( Y=>nx17462, A0=>nx16577, A1=>nx17452, A2=>
      nx17461);
   ix17914 : nor02_2x port map ( Y=>nx17463, A0=>nx17462, A1=>nx16661);
   ix17915 : aoi21 port map ( Y=>nx17464, A0=>nx16661, A1=>nx17462, B0=>
      nx17463);
   reg_nx2472 : nand02_2x port map ( Y=>nx2472, A0=>nx17145, A1=>nx15758);
   ix17916 : nor02_2x port map ( Y=>nx17465, A0=>nx17840, A1=>nx16602);
   reg_nx16597 : ao21 port map ( Y=>nx16597, A0=>nx17840, A1=>nx16602, B0=>
      nx17465);
   reg_nx4260 : oai22 port map ( Y=>nx4260, A0=>nx14780, A1=>nx17836, B0=>
      nx17455, B1=>nx17545);
   ix17917 : inv02 port map ( Y=>nx17466, A=>nx14780);
   ix17918 : inv02 port map ( Y=>nx17467, A=>nx17836);
   ix17919 : nand02_2x port map ( Y=>nx17468, A0=>write_offset_data_out_2, 
      A1=>nx17814);
   ix17920 : inv01 port map ( Y=>nx17469, A=>nx17804);
   ix17921 : inv01 port map ( Y=>nx17470, A=>nx17811);
   ix17922 : nand02_2x port map ( Y=>nx17471, A0=>nx17804, A1=>nx17812);
   ix17923 : nor02_2x port map ( Y=>nx17472, A0=>nx17806, A1=>nx17808);
   ix17924 : aoi22 port map ( Y=>nx17473, A0=>nx17469, A1=>nx17470, B0=>
      nx17471, B1=>nx17472);
   reg_nx15981 : inv02 port map ( Y=>nx15981, A=>nx17637);
   ix17925 : and02 port map ( Y=>nx17474, A0=>nx17804, A1=>nx17812);
   reg_nx2790 : oai32 port map ( Y=>nx2790, A0=>nx17474, A1=>nx17806, A2=>
      nx17808, B0=>nx17804, B1=>nx17812);
   reg_nx15800 : or02 port map ( Y=>nx15800, A0=>nx17806, A1=>nx17808);
   reg_nx15867 : oai22 port map ( Y=>nx15867, A0=>nx17469, A1=>nx17470, B0=>
      nx17804, B1=>nx17812);
   reg_nx16919 : inv02 port map ( Y=>nx16919, A=>nx17806);
   ix17926 : inv01 port map ( Y=>nx17475, A=>nx17424);
   ix17927 : oai22 port map ( Y=>nx17476, A0=>nx17185, A1=>nx14812, B0=>
      nx17428, B1=>nx17429);
   reg_nx16487 : aoi32 port map ( Y=>nx16487, A0=>nx17798, A1=>nx17431, A2=>
      nx17475, B0=>nx17431, B1=>nx17476);
   ix17928 : inv01 port map ( Y=>nx17477, A=>nx17418);
   ix17929 : inv02 port map ( Y=>nx17478, A=>new_size_squared_out_13);
   ix17930 : inv02 port map ( Y=>nx17479, A=>nx17836);
   ix17931 : aoi22 port map ( Y=>nx17480, A0=>nx17836, A1=>nx17478, B0=>
      new_size_squared_out_13, B1=>nx17479);
   ix17932 : nand02_2x port map ( Y=>nx17481, A0=>nx17477, A1=>nx17480);
   ix17933 : nor02_2x port map ( Y=>nx17482, A0=>nx17189, A1=>nx14801);
   ix17934 : nor02_2x port map ( Y=>nx17483, A0=>nx17480, A1=>nx17482);
   ix17935 : aoi222 port map ( Y=>nx17484, A0=>nx17418, A1=>nx17483, B0=>
      nx17480, B1=>nx17482, C0=>nx18303, C1=>nx17483);
   reg_nx16542 : oai21 port map ( Y=>nx16542, A0=>nx18303, A1=>nx17481, B0=>
      nx17484);
   reg_nx16545 : oai22 port map ( Y=>nx16545, A0=>nx17479, A1=>
      new_size_squared_out_13, B0=>nx17478, B1=>nx17837);
   ix17936 : nand02_2x port map ( Y=>nx17485, A0=>write_base_data_out_13, A1
      =>bias_offset_data_out_13);
   ix17937 : nand02_2x port map ( Y=>nx17486, A0=>write_base_data_out_11, A1
      =>bias_offset_data_out_11);
   ix17938 : nand02_2x port map ( Y=>nx17487, A0=>nx16482, A1=>nx17486);
   ix17939 : inv02 port map ( Y=>nx17488, A=>nx16482);
   ix17940 : and02 port map ( Y=>nx17489, A0=>write_base_data_out_11, A1=>
      bias_offset_data_out_11);
   ix17941 : nor02_2x port map ( Y=>nx17490, A0=>nx17488, A1=>nx17834);
   ix17942 : nor02_2x port map ( Y=>nx17491, A0=>nx17490, A1=>nx16413);
   ix17943 : aoi22 port map ( Y=>nx17492, A0=>nx17485, A1=>nx4222, B0=>
      nx16534, B1=>nx17485);
   ix17944 : nor02_2x port map ( Y=>nx17493, A0=>nx17447, A1=>nx17445);
   ix17945 : nand02_2x port map ( Y=>nx17494, A0=>nx17440, A1=>nx18301);
   ix17946 : and02 port map ( Y=>nx17495, A0=>nx17440, A1=>nx18301);
   ix17947 : nor03_2x port map ( Y=>nx17496, A0=>nx17492, A1=>nx17495, A2=>
      nx17447);
   reg_nx16594 : inv02 port map ( Y=>nx16594, A=>nx17492);
   ix17948 : inv02 port map ( Y=>nx17497, A=>nx16413);
   reg_nx16474 : oai22 port map ( Y=>nx16474, A0=>nx17489, A1=>nx17582, B0=>
      nx17497, B1=>nx17489);
   reg_nx17189 : inv02 port map ( Y=>nx17189, A=>nx17834);
   reg_nx16477 : oai22 port map ( Y=>nx16477, A0=>nx17189, A1=>nx16482, B0=>
      nx17488, B1=>nx17835);
   ix17949 : inv01 port map ( Y=>nx17498, A=>nx17392);
   ix17950 : nor02_2x port map ( Y=>nx17499, A0=>nx17394, A1=>nx16429);
   ix17951 : oai32 port map ( Y=>nx17500, A0=>nx17395, A1=>nx16501, A2=>
      nx17396, B0=>nx17189, B1=>nx17398);
   ix17952 : nor02_2x port map ( Y=>nx17501, A0=>nx17562, A1=>nx17392);
   ix17953 : inv02 port map ( Y=>nx17502, A=>new_size_squared_out_3);
   ix17954 : inv02 port map ( Y=>nx17503, A=>nx17816);
   ix17955 : oai22 port map ( Y=>nx17504, A0=>nx17502, A1=>nx17503, B0=>
      new_size_squared_out_3, B1=>nx17816);
   ix17956 : and02 port map ( Y=>nx17505, A0=>nx14854, A1=>nx17169);
   ix17957 : inv01 port map ( Y=>nx17506, A=>new_size_squared_out_1);
   ix17958 : inv01 port map ( Y=>nx17507, A=>nx17812);
   ix17959 : oai22 port map ( Y=>nx17508, A0=>nx17506, A1=>nx17507, B0=>
      new_size_squared_out_1, B1=>nx17813);
   ix17960 : inv02 port map ( Y=>nx17509, A=>nx17806);
   ix17961 : inv02 port map ( Y=>nx17510, A=>nx14854);
   reg_nx15946 : oai22 port map ( Y=>nx15946, A0=>nx17503, A1=>
      new_size_squared_out_3, B0=>nx17502, B1=>nx17816);
   reg_nx15836 : oai22 port map ( Y=>nx15836, A0=>nx17507, A1=>
      new_size_squared_out_1, B0=>nx17506, B1=>nx17813);
   ix17962 : inv02 port map ( Y=>nx17511, A=>new_size_squared_out_0);
   ix17963 : inv02 port map ( Y=>nx17512, A=>nx15860);
   reg_nx15917 : aoi32 port map ( Y=>nx15917, A0=>nx17512, A1=>
      bias_offset_data_out_0, A2=>nx16919, B0=>write_base_data_out_1, B1=>
      bias_offset_data_out_1);
   ix17964 : inv02 port map ( Y=>nx17513, A=>nx15924);
   ix17965 : inv02 port map ( Y=>nx17514, A=>nx17171);
   ix17966 : aoi22 port map ( Y=>nx17515, A0=>nx17171, A1=>nx17513, B0=>
      nx15924, B1=>nx17514);
   reg_nx17169 : inv02 port map ( Y=>nx17169, A=>nx17815);
   ix17967 : nor02ii port map ( Y=>nx17516, A0=>nx17818, A1=>nx16005);
   ix17968 : inv02 port map ( Y=>nx17517, A=>write_base_data_out_3);
   ix17969 : inv02 port map ( Y=>nx17518, A=>bias_offset_data_out_3);
   ix17970 : oai21 port map ( Y=>nx17519, A0=>nx17517, A1=>nx17518, B0=>
      nx18295);
   ix17971 : oai21 port map ( Y=>nx17520, A0=>nx17517, A1=>nx17518, B0=>
      nx17568);
   reg_nx15997 : nand02_2x port map ( Y=>nx15997, A0=>nx17519, A1=>nx17520);
   ix17972 : inv02 port map ( Y=>nx17521, A=>nx16005);
   reg_nx16000 : oai22 port map ( Y=>nx16000, A0=>nx17521, A1=>nx17818, B0=>
      nx17173, B1=>nx16005);
   ix17973 : inv01 port map ( Y=>nx17522, A=>nx17568);
   reg_nx15920 : oai22 port map ( Y=>nx15920, A0=>nx17513, A1=>nx17514, B0=>
      nx15924, B1=>nx17171);
   ix17974 : and02 port map ( Y=>nx17523, A0=>write_base_data_out_3, A1=>
      layer_mem_size_out_3);
   ix17975 : nor02ii port map ( Y=>nx17524, A0=>nx17523, A1=>nx15951);
   ix17976 : nand03_2x port map ( Y=>nx17525, A0=>nx17434, A1=>
      layer_mem_size_out_0, A2=>nx16919);
   ix17977 : inv02 port map ( Y=>nx17526, A=>nx17438);
   ix17978 : nand02_2x port map ( Y=>nx17527, A0=>nx17436, A1=>nx17437);
   ix17979 : nand02_2x port map ( Y=>nx17528, A0=>nx17432, A1=>nx17527);
   reg_nx16019 : inv02 port map ( Y=>nx16019, A=>nx17766);
   ix17980 : aoi22 port map ( Y=>nx17529, A0=>nx17435, A1=>nx17525, B0=>
      nx17436, B1=>nx17437);
   ix17981 : nor02ii port map ( Y=>nx17530, A0=>nx17455, A1=>nx17454);
   ix17982 : oai22 port map ( Y=>nx17531, A0=>nx14780, A1=>nx17837, B0=>
      nx17452, B1=>nx17453);
   ix17983 : inv02 port map ( Y=>nx17532, A=>nx14778);
   ix17984 : inv02 port map ( Y=>nx17533, A=>nx17832);
   ix17985 : nand02_2x port map ( Y=>nx17534, A0=>nx14778, A1=>nx17832);
   ix17986 : and02 port map ( Y=>nx17535, A0=>write_offset_data_out_10, A1=>
      nx17830);
   ix17987 : and02 port map ( Y=>nx17536, A0=>nx14778, A1=>nx17832);
   ix17988 : nor02_2x port map ( Y=>nx17537, A0=>nx17536, A1=>nx16394);
   ix17989 : aoi222 port map ( Y=>nx17538, A0=>nx17532, A1=>nx17533, B0=>
      nx17534, B1=>nx17535, C0=>nx3748, C1=>nx17537);
   ix17990 : inv02 port map ( Y=>nx17539, A=>nx17454);
   ix17991 : nor04_2x port map ( Y=>nx17540, A0=>nx17538, A1=>nx16513, A2=>
      nx17539, A3=>nx17455);
   ix17992 : aoi321 port map ( Y=>nx17541, A0=>nx17530, A1=>
      write_offset_data_out_12, A2=>nx17835, B0=>nx17454, B1=>nx17531, C0=>
      nx17540);
   ix17993 : inv01 port map ( Y=>nx17542, A=>nx17541);
   ix17994 : inv01 port map ( Y=>nx17543, A=>nx17541);
   ix17995 : nand02_2x port map ( Y=>nx17544, A0=>write_offset_data_out_12, 
      A1=>nx17835);
   ix17996 : inv02 port map ( Y=>nx17545, A=>NOT_nx16569);
   reg_nx4004 : inv01 port map ( Y=>nx4004, A=>nx17538);
   ix17997 : inv02 port map ( Y=>nx17546, A=>nx16394);
   reg_nx16448 : oai22 port map ( Y=>nx16448, A0=>nx17535, A1=>nx3748, B0=>
      nx17546, B1=>nx17535);
   reg_nx16451 : oai22 port map ( Y=>nx16451, A0=>nx17532, A1=>nx17533, B0=>
      nx14778, B1=>nx17832);
   ix17998 : nand02_2x port map ( Y=>nx17547, A0=>write_base_data_out_7, A1
      =>layer_mem_size_out_7);
   ix17999 : nand02_2x port map ( Y=>nx17548, A0=>nx16262, A1=>nx17547);
   ix18000 : inv02 port map ( Y=>nx17549, A=>nx16262);
   ix18001 : and02 port map ( Y=>nx17550, A0=>write_base_data_out_7, A1=>
      layer_mem_size_out_7);
   ix18002 : nor02_2x port map ( Y=>nx17551, A0=>nx17549, A1=>nx17824);
   ix18003 : nor02_2x port map ( Y=>nx17552, A0=>nx17551, A1=>nx16191);
   ix18004 : and02 port map ( Y=>nx17553, A0=>write_base_data_out_9, A1=>
      layer_mem_size_out_9);
   ix18005 : nor03_2x port map ( Y=>nx17554, A0=>nx17500, A1=>nx17553, A2=>
      nx17391);
   ix18006 : nor02ii port map ( Y=>nx17555, A0=>nx17553, A1=>nx16309);
   ix18007 : nor02ii port map ( Y=>nx17556, A0=>nx17555, A1=>nx17498);
   ix18008 : oai21 port map ( Y=>nx17557, A0=>nx17556, A1=>nx17391, B0=>
      nx17499);
   ix18009 : inv02 port map ( Y=>nx17558, A=>nx17500);
   reg_nx4154 : aoi22 port map ( Y=>nx4154, A0=>nx17751, A1=>nx17554, B0=>
      nx17557, B1=>nx17558);
   ix18010 : inv01 port map ( Y=>nx17559, A=>nx4154);
   ix18011 : nand02_2x port map ( Y=>nx17560, A0=>write_base_data_out_9, A1
      =>layer_mem_size_out_9);
   ix18012 : aoi21 port map ( Y=>nx17561, A0=>nx17560, A1=>nx17752, B0=>
      nx17555);
   reg_nx16375 : inv01 port map ( Y=>nx16375, A=>nx17561);
   ix18013 : inv01 port map ( Y=>nx17562, A=>nx17561);
   ix18014 : inv02 port map ( Y=>nx17563, A=>nx16191);
   reg_nx16255 : oai22 port map ( Y=>nx16255, A0=>nx17550, A1=>nx17754, B0=>
      nx17563, B1=>nx17550);
   reg_nx16258 : oai22 port map ( Y=>nx16258, A0=>nx17181, A1=>nx16262, B0=>
      nx17549, B1=>nx17824);
   ix18015 : inv01 port map ( Y=>nx17564, A=>nx17517);
   ix18016 : inv01 port map ( Y=>nx17565, A=>nx17516);
   ix18017 : inv01 port map ( Y=>nx17566, A=>nx17518);
   ix18018 : oai22 port map ( Y=>nx17567, A0=>nx15917, A1=>nx17515, B0=>
      nx17169, B1=>nx15924);
   ix18019 : inv02 port map ( Y=>nx17568, A=>nx17567);
   ix18020 : inv01 port map ( Y=>nx17569, A=>nx17173);
   ix18021 : inv02 port map ( Y=>nx17570, A=>nx16005);
   ix18022 : aoi22 port map ( Y=>nx17571, A0=>nx17835, A1=>nx17487, B0=>
      nx17488, B1=>nx17489);
   reg_nx17185 : inv02 port map ( Y=>nx17185, A=>nx17831);
   ix18023 : nand02_2x port map ( Y=>nx17572, A0=>nx16363, A1=>nx17185);
   ix18024 : inv02 port map ( Y=>nx17573, A=>nx16363);
   ix18025 : nand02_2x port map ( Y=>nx17574, A0=>write_base_data_out_7, A1
      =>bias_offset_data_out_7);
   ix18026 : nand02_2x port map ( Y=>nx17575, A0=>nx16243, A1=>nx17574);
   ix18027 : inv02 port map ( Y=>nx17576, A=>nx16243);
   ix18028 : and02 port map ( Y=>nx17577, A0=>write_base_data_out_7, A1=>
      bias_offset_data_out_7);
   ix18029 : nor02_2x port map ( Y=>nx17578, A0=>nx17576, A1=>nx17824);
   ix18030 : nor02_2x port map ( Y=>nx17579, A0=>nx17578, A1=>nx16175);
   ix18031 : nor02ii port map ( Y=>nx17580, A0=>nx17831, A1=>nx16363);
   ix18032 : inv02 port map ( Y=>nx17581, A=>nx17491);
   reg_nx3966 : inv01 port map ( Y=>nx3966, A=>nx17633);
   ix18033 : inv01 port map ( Y=>nx17582, A=>nx17633);
   ix18034 : nand02_2x port map ( Y=>nx17583, A0=>write_base_data_out_9, A1
      =>bias_offset_data_out_9);
   ix18035 : inv02 port map ( Y=>nx17584, A=>nx16293);
   ix18036 : and02 port map ( Y=>nx17585, A0=>write_base_data_out_9, A1=>
      bias_offset_data_out_9);
   ix18037 : nor02_2x port map ( Y=>nx17586, A0=>nx17584, A1=>nx17585);
   reg_nx16355 : ao21 port map ( Y=>nx16355, A0=>nx17583, A1=>nx17692, B0=>
      nx17586);
   reg_nx16358 : oai22 port map ( Y=>nx16358, A0=>nx17573, A1=>nx17831, B0=>
      nx17185, B1=>nx16363);
   ix18038 : inv02 port map ( Y=>nx17587, A=>nx16175);
   reg_nx16235 : oai22 port map ( Y=>nx16235, A0=>nx17577, A1=>nx3454, B0=>
      nx17587, B1=>nx17577);
   reg_nx16238 : oai22 port map ( Y=>nx16238, A0=>nx17181, A1=>nx16243, B0=>
      nx17576, B1=>nx17824);
   ix18039 : inv02 port map ( Y=>nx17588, A=>write_base_data_out_11);
   ix18040 : inv02 port map ( Y=>nx17589, A=>nx17835);
   ix18041 : nand02_2x port map ( Y=>nx17590, A0=>write_base_data_out_14, A1
      =>nx17831);
   ix18042 : nor04_2x port map ( Y=>nx17591, A0=>nx17588, A1=>nx17461, A2=>
      nx17589, A3=>nx17590);
   reg_nx4336 : oai22 port map ( Y=>nx4336, A0=>nx17591, A1=>nx17827, B0=>
      nx17827, B1=>nx17828);
   ix18043 : inv02 port map ( Y=>nx17592, A=>nx17831);
   ix18044 : nor04_2x port map ( Y=>nx17593, A0=>nx17589, A1=>nx17588, A2=>
      nx17592, A3=>nx17461);
   ix18045 : and02 port map ( Y=>nx17594, A0=>write_base_data_out_11, A1=>
      nx17831);
   reg_nx3926 : and02 port map ( Y=>nx3926, A0=>nx17828, A1=>nx17594);
   reg_nx16456 : nand02_2x port map ( Y=>nx16456, A0=>nx17831, A1=>nx17829);
   ix18046 : nand02_2x port map ( Y=>nx17595, A0=>nx17416, A1=>nx17427);
   ix18047 : inv02 port map ( Y=>nx17596, A=>nx17430);
   ix18048 : oai21 port map ( Y=>nx17597, A0=>nx17430, A1=>nx17425, B0=>
      nx17426);
   ix18049 : nand02_2x port map ( Y=>nx17598, A0=>nx17422, A1=>nx17736);
   reg_nx16605 : oai21 port map ( Y=>nx16605, A0=>nx17737, A1=>nx17421, B0=>
      nx17598);
   ix18050 : nand02_2x port map ( Y=>nx17599, A0=>write_base_data_out_5, A1
      =>new_size_squared_out_5);
   ix18051 : nand02_2x port map ( Y=>nx17600, A0=>nx14843, A1=>nx17173);
   ix18052 : inv02 port map ( Y=>nx17601, A=>nx14843);
   ix18053 : aoi322 port map ( Y=>nx17602, A0=>nx17508, A1=>
      new_size_squared_out_0, A2=>nx17509, B0=>nx17815, B1=>nx17510, C0=>
      new_size_squared_out_1, C1=>write_base_data_out_1);
   reg_nx2854 : nor02_2x port map ( Y=>nx2854, A0=>nx17602, A1=>nx17505);
   ix18054 : nor02_2x port map ( Y=>nx17603, A0=>nx17601, A1=>nx17818);
   ix18055 : nor02ii port map ( Y=>nx17604, A0=>nx17603, A1=>nx17504);
   ix18056 : aoi322 port map ( Y=>nx17605, A0=>nx17600, A1=>
      write_base_data_out_3, A2=>new_size_squared_out_3, B0=>nx17818, B1=>
      nx17601, C0=>nx2854, C1=>nx17604);
   ix18057 : aoi22 port map ( Y=>nx17606, A0=>nx17599, A1=>nx17605, B0=>
      nx16068, B1=>nx17599);
   reg_nx16129 : inv01 port map ( Y=>nx16129, A=>nx17606);
   ix18058 : inv01 port map ( Y=>nx17607, A=>nx17606);
   reg_nx3116 : inv02 port map ( Y=>nx3116, A=>nx17605);
   ix18059 : and02 port map ( Y=>nx17608, A0=>write_base_data_out_3, A1=>
      new_size_squared_out_3);
   reg_nx16012 : oai22 port map ( Y=>nx16012, A0=>nx17608, A1=>nx17504, B0=>
      nx2854, B1=>nx17608);
   reg_nx16015 : oai22 port map ( Y=>nx16015, A0=>nx17601, A1=>nx17818, B0=>
      nx17173, B1=>nx14843);
   reg_nx17025 : inv02 port map ( Y=>nx17025, A=>nx2532);
   ix18060 : aoi32 port map ( Y=>nx17609, A0=>nx17572, A1=>
      write_base_data_out_9, A2=>bias_offset_data_out_9, B0=>nx17831, B1=>
      nx17573);
   ix18061 : or02 port map ( Y=>nx17610, A0=>nx17609, A1=>nx17581);
   reg_nx4222 : and03 port map ( Y=>nx4222, A0=>nx17610, A1=>nx17571, A2=>
      nx17690);
   ix18062 : inv02 port map ( Y=>nx17611, A=>nx16538);
   ix18063 : inv02 port map ( Y=>nx17612, A=>nx17837);
   ix18064 : aoi22 port map ( Y=>nx17613, A0=>nx16538, A1=>nx17837, B0=>
      nx17611, B1=>nx17612);
   ix18065 : and02 port map ( Y=>nx17614, A0=>nx4222, A1=>nx17613);
   ix18066 : nor02_2x port map ( Y=>nx17615, A0=>nx4222, A1=>nx17613);
   ix18067 : nor02_2x port map ( Y=>nx17616, A0=>nx17614, A1=>nx17615);
   ix18068 : inv02 port map ( Y=>nx17617, A=>nx16939);
   reg_nx16572 : oai22 port map ( Y=>nx16572, A0=>nx17466, A1=>nx17467, B0=>
      nx17837, B1=>nx14780);
   ix18069 : inv02 port map ( Y=>nx17618, A=>nx16572);
   ix18070 : nor02_2x port map ( Y=>nx17619, A0=>nx17538, A1=>nx16513);
   ix18071 : nor02ii port map ( Y=>nx17620, A0=>nx17619, A1=>nx17544);
   ix18072 : nor02_2x port map ( Y=>nx17621, A0=>nx17618, A1=>nx17620);
   ix18073 : aoi21 port map ( Y=>nx17622, A0=>nx17618, A1=>nx17620, B0=>
      nx17621);
   ix18074 : nor02_2x port map ( Y=>nx17623, A0=>nx16557, A1=>nx17015);
   ix18075 : inv02 port map ( Y=>nx17624, A=>nx17829);
   ix18076 : inv01 port map ( Y=>nx17625, A=>nx17827);
   ix18077 : inv01 port map ( Y=>nx17626, A=>nx17593);
   ix18078 : nand02_2x port map ( Y=>nx17627, A0=>nx17625, A1=>nx17626);
   ix18079 : inv02 port map ( Y=>nx17628, A=>nx17835);
   ix18080 : inv02 port map ( Y=>nx17629, A=>nx17594);
   ix18081 : oai43 port map ( Y=>nx17630, A0=>nx17624, A1=>nx17627, A2=>
      nx17628, A3=>nx17629, B0=>nx16580, B1=>nx4194, B2=>nx16983);
   ix18082 : oai33 port map ( Y=>nx17631, A0=>nx17827, A1=>nx17837, A2=>
      nx17593, B0=>nx17829, B1=>nx17837, B2=>nx17827);
   ix18083 : nor03_2x port map ( Y=>nx17632, A0=>nx17623, A1=>nx17630, A2=>
      nx17631);
   reg_mem_addr_out_13 : oai221 port map ( Y=>mem_addr_out(13), A0=>nx17025, 
      A1=>nx17616, B0=>nx17617, B1=>nx17622, C0=>nx17632);
   reg_nx16534 : oai22 port map ( Y=>nx16534, A0=>nx17611, A1=>nx17612, B0=>
      nx16538, B1=>nx17837);
   ix18084 : nor02ii port map ( Y=>nx17633, A0=>nx17691, A1=>nx17609);
   reg_nx4204 : and02 port map ( Y=>nx4204, A0=>nx17829, A1=>nx17593);
   reg_NOT_nx16569 : oai21 port map ( Y=>NOT_nx16569, A0=>nx17538, A1=>
      nx16513, B0=>nx17544);
   reg_nx16577 : nand03_2x port map ( Y=>nx16577, A0=>nx17829, A1=>nx17835, 
      A2=>nx17594);
   ix18085 : inv02 port map ( Y=>nx17634, A=>nx14751);
   ix18086 : inv02 port map ( Y=>nx17635, A=>nx17816);
   ix18087 : nand02_2x port map ( Y=>nx17636, A0=>nx14751, A1=>nx17817);
   ix18088 : oai21 port map ( Y=>nx17637, A0=>nx17473, A1=>nx15905, B0=>
      nx17468);
   ix18089 : and02 port map ( Y=>nx17638, A0=>nx14736, A1=>nx17821);
   ix18090 : inv02 port map ( Y=>nx17639, A=>write_offset_data_out_4);
   ix18091 : inv02 port map ( Y=>nx17640, A=>nx17818);
   reg_nx3236 : inv02 port map ( Y=>nx3236, A=>nx17678);
   ix18092 : nand02_2x port map ( Y=>nx17641, A0=>write_offset_data_out_4, 
      A1=>nx17819);
   ix18093 : inv02 port map ( Y=>nx17642, A=>nx16033);
   ix18094 : and02 port map ( Y=>nx17643, A0=>write_offset_data_out_4, A1=>
      nx17819);
   ix18095 : nor02_2x port map ( Y=>nx17644, A0=>nx17642, A1=>nx17643);
   reg_nx16091 : ao21 port map ( Y=>nx16091, A0=>nx17641, A1=>nx17681, B0=>
      nx17644);
   ix18096 : inv02 port map ( Y=>nx17645, A=>nx14736);
   ix18097 : inv02 port map ( Y=>nx17646, A=>nx17821);
   reg_nx16094 : oai22 port map ( Y=>nx16094, A0=>nx17645, A1=>nx17646, B0=>
      nx14736, B1=>nx17821);
   reg_nx2972 : inv01 port map ( Y=>nx2972, A=>nx17681);
   reg_nx15984 : oai22 port map ( Y=>nx15984, A0=>nx17634, A1=>nx17635, B0=>
      nx14751, B1=>nx17817);
   ix18098 : and02 port map ( Y=>nx17647, A0=>nx17810, A1=>nx17813);
   ix18099 : nor02_2x port map ( Y=>nx17648, A0=>nx17647, A1=>nx18293);
   ix18100 : nor02_2x port map ( Y=>nx17649, A0=>nx17810, A1=>nx17813);
   ix18101 : nor02_2x port map ( Y=>nx17650, A0=>nx17648, A1=>nx17649);
   ix18102 : nand02_2x port map ( Y=>nx17651, A0=>write_base_data_out_5, A1
      =>nx17819);
   ix18103 : and02 port map ( Y=>nx17652, A0=>nx15374, A1=>nx17817);
   ix18104 : nand02_2x port map ( Y=>nx17653, A0=>nx15374, A1=>nx17817);
   ix18105 : inv02 port map ( Y=>nx17654, A=>nx15374);
   ix18106 : inv02 port map ( Y=>nx17655, A=>nx17817);
   ix18107 : aoi32 port map ( Y=>nx17656, A0=>nx17653, A1=>
      class_cntr_counter_out_2, A2=>nx17815, B0=>nx17654, B1=>nx17655);
   ix18108 : inv02 port map ( Y=>nx17657, A=>write_base_data_out_5);
   ix18109 : inv02 port map ( Y=>nx17658, A=>nx17819);
   ix18110 : oai43 port map ( Y=>nx17659, A0=>nx17650, A1=>nx17651, A2=>
      nx17652, A3=>nx15878, B0=>nx17656, B1=>nx17657, B2=>nx17658);
   reg_nx3180 : inv02 port map ( Y=>nx3180, A=>nx17720);
   ix18111 : inv02 port map ( Y=>nx17660, A=>nx17720);
   ix18112 : inv02 port map ( Y=>nx17661, A=>class_cntr_counter_out_2);
   ix18113 : inv02 port map ( Y=>nx17662, A=>nx17815);
   reg_nx3026 : oai332 port map ( Y=>nx3026, A0=>nx17650, A1=>nx17652, A2=>
      nx15878, B0=>nx17652, B1=>nx17661, B2=>nx17662, C0=>nx15374, C1=>
      nx17817);
   ix18114 : inv02 port map ( Y=>nx17663, A=>nx3026);
   reg_nx16099 : nor02_2x port map ( Y=>nx16099, A0=>nx17658, A1=>nx17663);
   ix18115 : inv02 port map ( Y=>nx17664, A=>nx16099);
   ix18116 : inv01 port map ( Y=>nx17665, A=>nx17663);
   ix18117 : and02 port map ( Y=>nx17666, A0=>class_cntr_counter_out_2, A1=>
      nx17815);
   ix18118 : inv02 port map ( Y=>nx17667, A=>nx15878);
   reg_nx15936 : oai32 port map ( Y=>nx15936, A0=>nx17666, A1=>nx17648, A2=>
      nx17649, B0=>nx17667, B1=>nx17666);
   reg_nx15939 : oai22 port map ( Y=>nx15939, A0=>nx17654, A1=>nx17655, B0=>
      nx15374, B1=>nx17817);
   reg_nx2808 : oai22 port map ( Y=>nx2808, A0=>nx17810, A1=>nx17813, B0=>
      nx17647, B1=>nx18293);
   ix18119 : inv01 port map ( Y=>nx17668, A=>nx17810);
   ix18120 : inv01 port map ( Y=>nx17669, A=>nx17813);
   reg_nx15825 : oai22 port map ( Y=>nx15825, A0=>nx17668, A1=>nx17669, B0=>
      nx17810, B1=>nx17813);
   ix18121 : nand02_2x port map ( Y=>nx17670, A0=>write_offset_data_out_6, 
      A1=>nx17822);
   ix18122 : inv02 port map ( Y=>nx17671, A=>nx17638);
   ix18123 : inv02 port map ( Y=>nx17672, A=>nx16033);
   ix18124 : inv02 port map ( Y=>nx17673, A=>nx14736);
   ix18125 : inv02 port map ( Y=>nx17674, A=>nx17821);
   ix18126 : inv02 port map ( Y=>nx17675, A=>nx17635);
   ix18127 : inv02 port map ( Y=>nx17676, A=>nx17634);
   ix18128 : oai32 port map ( Y=>nx17677, A0=>nx17675, A1=>nx17676, A2=>
      nx16033, B0=>nx17639, B1=>nx17640);
   ix18129 : aoi422 port map ( Y=>nx17678, A0=>nx17671, A1=>nx17637, A2=>
      nx17636, A3=>nx17672, B0=>nx17673, B1=>nx17674, C0=>nx17677, C1=>
      nx17671);
   ix18130 : aoi22 port map ( Y=>nx17679, A0=>nx16155, A1=>nx17670, B0=>
      nx17670, B1=>nx17678);
   reg_nx16210 : inv02 port map ( Y=>nx16210, A=>nx17679);
   ix18131 : inv02 port map ( Y=>nx17680, A=>nx17679);
   ix18132 : aoi22 port map ( Y=>nx17681, A0=>nx17634, A1=>nx17635, B0=>
      nx17636, B1=>nx17637);
   ix18133 : aoi22 port map ( Y=>nx17682, A0=>nx17825, A1=>nx17575, B0=>
      nx17576, B1=>nx17577);
   ix18134 : nor03_2x port map ( Y=>nx17683, A0=>nx17682, A1=>nx17580, A2=>
      nx16293);
   ix18135 : nand02_2x port map ( Y=>nx17684, A0=>nx16124, A1=>nx17177);
   ix18136 : nor02ii port map ( Y=>nx17685, A0=>nx17822, A1=>nx16124);
   ix18137 : nor02_2x port map ( Y=>nx17686, A0=>nx17685, A1=>nx16057);
   ix18138 : nor02ii port map ( Y=>nx17687, A0=>nx16124, A1=>nx17822);
   ix18139 : inv02 port map ( Y=>nx17688, A=>nx17579);
   ix18140 : nor02_2x port map ( Y=>nx17689, A0=>nx17683, A1=>nx17704);
   ix18141 : or02 port map ( Y=>nx17690, A0=>nx17581, A1=>nx17689);
   ix18142 : inv01 port map ( Y=>nx17691, A=>nx17689);
   reg_nx3710 : aoi22 port map ( Y=>nx3710, A0=>nx17682, A1=>nx17717, B0=>
      nx17682, B1=>nx17688);
   ix18143 : inv02 port map ( Y=>nx17692, A=>nx3710);
   ix18144 : and02 port map ( Y=>nx17693, A0=>write_base_data_out_5, A1=>
      bias_offset_data_out_5);
   ix18145 : inv02 port map ( Y=>nx17694, A=>nx16057);
   reg_nx16116 : oai22 port map ( Y=>nx16116, A0=>nx17693, A1=>nx18305, B0=>
      nx17694, B1=>nx17693);
   ix18146 : inv02 port map ( Y=>nx17695, A=>nx16124);
   reg_nx16119 : oai22 port map ( Y=>nx16119, A0=>nx17695, A1=>nx17822, B0=>
      nx17177, B1=>nx16124);
   ix18147 : inv02 port map ( Y=>nx17696, A=>nx17564);
   ix18148 : inv02 port map ( Y=>nx17697, A=>nx17566);
   ix18149 : oai22 port map ( Y=>nx17698, A0=>nx17696, A1=>nx17697, B0=>
      nx18295, B1=>nx17568);
   ix18150 : nand03_2x port map ( Y=>nx17699, A0=>nx17698, A1=>nx17686, A2=>
      nx17565);
   ix18151 : nand03_2x port map ( Y=>nx17700, A0=>nx17569, A1=>nx17686, A2=>
      nx17570);
   ix18152 : and03 port map ( Y=>nx17701, A0=>nx17684, A1=>
      write_base_data_out_5, A2=>bias_offset_data_out_5);
   ix18153 : nor02_2x port map ( Y=>nx17702, A0=>nx17701, A1=>nx17687);
   ix18154 : and03 port map ( Y=>nx17703, A0=>nx17699, A1=>nx17700, A2=>
      nx17702);
   ix18155 : nor04_2x port map ( Y=>nx17704, A0=>nx17703, A1=>nx17688, A2=>
      nx17580, A3=>nx16293);
   ix18156 : inv02 port map ( Y=>nx17705, A=>nx17569);
   ix18157 : nor02_2x port map ( Y=>nx17706, A0=>nx17566, A1=>nx17570);
   ix18158 : aoi322 port map ( Y=>nx17707, A0=>nx17568, A1=>nx17697, A2=>
      nx17705, B0=>nx17568, B1=>nx17706, C0=>nx18295, C1=>nx17706);
   ix18159 : nor02_2x port map ( Y=>nx17708, A0=>nx17564, A1=>nx17569);
   ix18160 : nor02_2x port map ( Y=>nx17709, A0=>nx17566, A1=>nx17569);
   ix18161 : aoi22 port map ( Y=>nx17710, A0=>nx17568, A1=>nx17708, B0=>
      nx18295, B1=>nx17709);
   ix18162 : nor02_2x port map ( Y=>nx17711, A0=>nx17564, A1=>nx17570);
   ix18163 : aoi22 port map ( Y=>nx17712, A0=>nx18295, A1=>nx17711, B0=>
      nx17568, B1=>nx17711);
   ix18164 : inv02 port map ( Y=>nx17713, A=>nx17565);
   ix18165 : inv02 port map ( Y=>nx17714, A=>nx17570);
   ix18166 : aoi222 port map ( Y=>nx17715, A0=>nx17713, A1=>nx17705, B0=>
      nx17713, B1=>nx17714, C0=>nx18295, C1=>nx17708);
   reg_nx3198 : and04 port map ( Y=>nx3198, A0=>nx17707, A1=>nx17710, A2=>
      nx17712, A3=>nx17715);
   ix18167 : oai33 port map ( Y=>nx17716, A0=>nx3198, A1=>nx17701, A2=>
      nx17687, B0=>nx17701, B1=>nx17686, B2=>nx17687);
   reg_nx3454 : inv01 port map ( Y=>nx3454, A=>nx17716);
   ix18168 : inv02 port map ( Y=>nx17717, A=>nx3454);
   ix18169 : oai332 port map ( Y=>nx17718, A0=>nx17713, A1=>nx18297, A2=>
      nx17568, B0=>nx17713, B1=>nx17696, B2=>nx17697, C0=>nx17705, C1=>
      nx17714);
   ix18170 : and02 port map ( Y=>nx17719, A0=>write_base_data_out_7, A1=>
      nx17822);
   reg_nx16336 : nand03_2x port map ( Y=>nx16336, A0=>nx17659, A1=>nx17825, 
      A2=>nx17719);
   reg_nx3436 : and02 port map ( Y=>nx3436, A0=>nx17659, A1=>nx17719);
   reg_nx16218 : nand02_2x port map ( Y=>nx16218, A0=>nx17823, A1=>nx17659);
   ix18171 : inv02 port map ( Y=>nx17720, A=>nx17659);
   ix18172 : nor02ii port map ( Y=>nx17721, A0=>nx14833, A1=>nx17823);
   ix18173 : inv02 port map ( Y=>nx17722, A=>nx14833);
   ix18174 : nor02_2x port map ( Y=>nx17723, A0=>nx17722, A1=>nx17823);
   ix18175 : nor02_2x port map ( Y=>nx17724, A0=>nx17723, A1=>nx17607);
   ix18176 : nor02_2x port map ( Y=>nx17725, A0=>nx17721, A1=>nx17724);
   ix18177 : inv02 port map ( Y=>nx17726, A=>nx14822);
   ix18178 : nor02_2x port map ( Y=>nx17727, A0=>nx17726, A1=>nx17825);
   ix18179 : inv02 port map ( Y=>nx17728, A=>write_base_data_out_7);
   ix18180 : inv02 port map ( Y=>nx17729, A=>new_size_squared_out_7);
   reg_nx17181 : inv02 port map ( Y=>nx17181, A=>nx17825);
   ix18181 : and02 port map ( Y=>nx17730, A0=>write_base_data_out_7, A1=>
      new_size_squared_out_7);
   ix18182 : nor02_2x port map ( Y=>nx17731, A0=>nx17726, A1=>nx17730);
   reg_nx3628 : oai332 port map ( Y=>nx3628, A0=>nx17725, A1=>nx17727, A2=>
      nx16186, B0=>nx14822, B1=>nx17728, B2=>nx17729, C0=>nx17181, C1=>
      nx17731);
   ix18183 : inv01 port map ( Y=>nx17732, A=>nx3628);
   ix18184 : and02 port map ( Y=>nx17733, A0=>write_base_data_out_9, A1=>
      new_size_squared_out_9);
   ix18185 : nor02ii port map ( Y=>nx17734, A0=>nx17733, A1=>nx17596);
   ix18186 : oai321 port map ( Y=>nx17735, A0=>nx17732, A1=>nx17597, A2=>
      nx16304, B0=>nx17734, B1=>nx17597, C0=>nx17595);
   reg_NOT_nx16607 : inv01 port map ( Y=>NOT_nx16607, A=>nx17735);
   ix18187 : inv01 port map ( Y=>nx17736, A=>NOT_nx16607);
   ix18188 : inv01 port map ( Y=>nx17737, A=>NOT_nx16607);
   ix18189 : nand02_2x port map ( Y=>nx17738, A0=>write_base_data_out_9, A1
      =>new_size_squared_out_9);
   reg_nx16368 : inv02 port map ( Y=>nx16368, A=>nx17798);
   ix18190 : inv02 port map ( Y=>nx17739, A=>nx17732);
   ix18191 : inv02 port map ( Y=>nx17740, A=>nx16186);
   reg_nx16248 : oai32 port map ( Y=>nx16248, A0=>nx17730, A1=>nx17721, A2=>
      nx17724, B0=>nx17740, B1=>nx17730);
   reg_nx16251 : oai22 port map ( Y=>nx16251, A0=>nx17181, A1=>nx14822, B0=>
      nx17726, B1=>nx17825);
   reg_nx3372 : oai22 port map ( Y=>nx3372, A0=>nx17723, A1=>nx17607, B0=>
      nx17177, B1=>nx14833);
   reg_nx16132 : oai22 port map ( Y=>nx16132, A0=>nx17722, A1=>nx17823, B0=>
      nx17177, B1=>nx14833);
   ix18192 : aoi22 port map ( Y=>nx17741, A0=>nx17825, A1=>nx17548, B0=>
      nx17549, B1=>nx17550);
   reg_nx17173 : inv02 port map ( Y=>nx17173, A=>nx17819);
   ix18193 : nand02_2x port map ( Y=>nx17742, A0=>nx16026, A1=>nx17173);
   ix18194 : nor02ii port map ( Y=>nx17743, A0=>nx16026, A1=>nx17819);
   ix18195 : inv02 port map ( Y=>nx17744, A=>nx16143);
   ix18196 : nor02_2x port map ( Y=>nx17745, A0=>nx17744, A1=>nx17823);
   ix18197 : inv02 port map ( Y=>nx17746, A=>write_base_data_out_5);
   ix18198 : inv02 port map ( Y=>nx17747, A=>layer_mem_size_out_5);
   reg_nx17177 : inv02 port map ( Y=>nx17177, A=>nx17823);
   ix18199 : and02 port map ( Y=>nx17748, A0=>write_base_data_out_5, A1=>
      layer_mem_size_out_5);
   ix18200 : nor02_2x port map ( Y=>nx17749, A0=>nx17744, A1=>nx17748);
   ix18201 : inv02 port map ( Y=>nx17750, A=>nx17552);
   reg_nx3642 : aoi22 port map ( Y=>nx3642, A0=>nx17741, A1=>NOT_nx3386, B0
      =>nx17750, B1=>nx17741);
   ix18202 : inv01 port map ( Y=>nx17751, A=>nx3642);
   ix18203 : inv01 port map ( Y=>nx17752, A=>nx3642);
   ix18204 : inv02 port map ( Y=>nx17753, A=>NOT_nx3386);
   ix18205 : inv02 port map ( Y=>nx17754, A=>NOT_nx3386);
   ix18206 : nor02ii port map ( Y=>nx17755, A0=>nx17819, A1=>nx16026);
   ix18207 : nor02ii port map ( Y=>nx17756, A0=>nx17755, A1=>nx17766);
   ix18208 : inv02 port map ( Y=>nx17757, A=>nx16073);
   reg_nx16136 : oai32 port map ( Y=>nx16136, A0=>nx17748, A1=>nx17743, A2=>
      nx17756, B0=>nx17757, B1=>nx17748);
   reg_nx16139 : oai22 port map ( Y=>nx16139, A0=>nx17177, A1=>nx16143, B0=>
      nx17744, B1=>nx17823);
   reg_nx3130 : inv02 port map ( Y=>nx3130, A=>nx17765);
   ix18209 : inv02 port map ( Y=>nx17758, A=>nx16026);
   reg_nx16022 : oai22 port map ( Y=>nx16022, A0=>nx17758, A1=>nx17819, B0=>
      nx17173, B1=>nx16026);
   ix18210 : inv02 port map ( Y=>nx17759, A=>nx17742);
   ix18211 : or02 port map ( Y=>nx17760, A0=>nx17745, A1=>nx16073);
   ix18212 : nor04_2x port map ( Y=>nx17761, A0=>nx17759, A1=>nx17524, A2=>
      nx17801, A3=>nx17760);
   ix18213 : inv02 port map ( Y=>nx17762, A=>nx17743);
   ix18214 : oai332 port map ( Y=>nx17763, A0=>nx17762, A1=>nx17745, A2=>
      nx16073, B0=>nx17746, B1=>nx16143, B2=>nx17747, C0=>nx17177, C1=>
      nx17749);
   reg_NOT_nx3386 : nor02_2x port map ( Y=>NOT_nx3386, A0=>nx17761, A1=>
      nx18307);
   ix18215 : oai21 port map ( Y=>nx17764, A0=>nx2868, A1=>nx17523, B0=>
      nx17742);
   ix18216 : ao22 port map ( Y=>nx17765, A0=>nx17764, A1=>nx17762, B0=>
      nx17524, B1=>nx17762);
   ix18217 : nor02_2x port map ( Y=>nx17766, A0=>nx17801, A1=>nx17524);
   ix18218 : oai222 port map ( Y=>nx17767, A0=>nx17458, A1=>nx17459, B0=>
      nx17460, B1=>nx17464, C0=>nx16689, C1=>nx16985);
   ix18219 : inv02 port map ( Y=>nx17768, A=>nx17767);
   ix18220 : or02 port map ( Y=>nx17769, A0=>nx17492, A1=>nx17494);
   ix18221 : nand02_2x port map ( Y=>nx17770, A0=>nx17451, A1=>nx17543);
   ix18222 : nor02ii port map ( Y=>nx17771, A0=>nx17457, A1=>nx17448);
   ix18223 : aoi322 port map ( Y=>nx17772, A0=>nx17769, A1=>nx2532, A2=>
      nx17493, B0=>nx2532, B1=>nx17496, C0=>nx17770, C1=>nx17771);
   reg_mem_addr_out_15 : nand02_2x port map ( Y=>mem_addr_out(15), A0=>
      nx17768, A1=>nx17772);
   reg_nx17215 : inv02 port map ( Y=>nx17215, A=>current_state_24);
   ix18224 : inv02 port map ( Y=>nx17773, A=>new_size_squared_out_15);
   ix18225 : inv02 port map ( Y=>nx17774, A=>write_base_data_out_15);
   ix18226 : oai22 port map ( Y=>nx17775, A0=>nx17773, A1=>nx17774, B0=>
      new_size_squared_out_15, B1=>write_base_data_out_15);
   ix18227 : oai22 port map ( Y=>nx17776, A0=>nx17774, A1=>
      new_size_squared_out_15, B0=>nx17773, B1=>write_base_data_out_15);
   ix18228 : inv01 port map ( Y=>nx17777, A=>nx4406);
   ix18229 : aoi22 port map ( Y=>nx17778, A0=>nx4406, A1=>nx17775, B0=>
      nx17776, B1=>nx17777);
   reg_nx14477 : oai222 port map ( Y=>nx14477, A0=>nx17215, A1=>nx16663, B0
      =>nx16661, B1=>nx16927, C0=>nx17778, C1=>nx16951);
   ix18230 : inv02 port map ( Y=>nx17779, A=>nx17732);
   ix18231 : inv01 port map ( Y=>nx17780, A=>nx17424);
   ix18232 : inv02 port map ( Y=>nx17781, A=>nx16304);
   ix18233 : inv01 port map ( Y=>nx17782, A=>nx17185);
   ix18234 : inv02 port map ( Y=>nx17783, A=>nx14812);
   ix18235 : inv02 port map ( Y=>nx17784, A=>nx17738);
   ix18236 : aoi322 port map ( Y=>nx17785, A0=>nx17779, A1=>nx17780, A2=>
      nx17781, B0=>nx17782, B1=>nx17783, C0=>nx17780, C1=>nx17784);
   ix18237 : inv02 port map ( Y=>nx17786, A=>new_size_squared_out_11);
   ix18238 : inv02 port map ( Y=>nx17787, A=>nx17833);
   ix18239 : aoi22 port map ( Y=>nx17788, A0=>nx17833, A1=>nx17786, B0=>
      new_size_squared_out_11, B1=>nx17787);
   ix18240 : nor02_2x port map ( Y=>nx17789, A0=>nx17785, A1=>nx17788);
   ix18241 : aoi21 port map ( Y=>nx17790, A0=>nx17785, A1=>nx17788, B0=>
      nx17789);
   reg_nx16943 : inv02 port map ( Y=>nx16943, A=>current_state_24);
   ix18242 : inv02 port map ( Y=>nx17791, A=>nx16382);
   ix18243 : inv01 port map ( Y=>nx17792, A=>nx17392);
   ix18244 : aoi22 port map ( Y=>nx17793, A0=>nx17782, A1=>nx17791, B0=>
      nx17561, B1=>nx17792);
   ix18245 : inv02 port map ( Y=>nx17794, A=>layer_mem_size_out_11);
   ix18246 : aoi22 port map ( Y=>nx17795, A0=>nx17833, A1=>nx17794, B0=>
      layer_mem_size_out_11, B1=>nx17787);
   ix18247 : nor02_2x port map ( Y=>nx17796, A0=>nx17793, A1=>nx17795);
   ix18248 : aoi21 port map ( Y=>nx17797, A0=>nx17793, A1=>nx17795, B0=>
      nx17796);
   reg_nx14267 : oai222 port map ( Y=>nx14267, A0=>nx17790, A1=>nx16951, B0
      =>nx17833, B1=>nx16925, C0=>nx16943, C1=>nx17797);
   reg_nx16424 : oai22 port map ( Y=>nx16424, A0=>nx17787, A1=>
      new_size_squared_out_11, B0=>nx17786, B1=>nx17833);
   reg_nx16429 : oai22 port map ( Y=>nx16429, A0=>nx17787, A1=>
      layer_mem_size_out_11, B0=>nx17794, B1=>nx17833);
   ix18249 : oai21 port map ( Y=>nx17798, A0=>nx17732, A1=>nx16304, B0=>
      nx17738);
   ix18250 : aoi21 port map ( Y=>nx17799, A0=>nx17525, A1=>nx17435, B0=>
      nx17528);
   ix18251 : inv01 port map ( Y=>nx17800, A=>nx17526);
   ix18252 : nor03_2x port map ( Y=>nx17801, A0=>nx17799, A1=>nx17800, A2=>
      nx17523);
   ix18253 : ao21 port map ( Y=>nx17802, A0=>nx17525, A1=>nx17435, B0=>
      nx17528);
   reg_nx2868 : nand02_2x port map ( Y=>nx2868, A0=>nx17526, A1=>nx17802);
   ix18254 : buf16 port map ( Y=>nx17803, A=>nx14762);
   ix18255 : buf16 port map ( Y=>nx17804, A=>nx14762);
   ix18256 : buf16 port map ( Y=>nx17805, A=>nx15777);
   ix18257 : buf16 port map ( Y=>nx17806, A=>nx15777);
   ix18258 : buf16 port map ( Y=>nx17807, A=>nx14769);
   ix18259 : buf16 port map ( Y=>nx17808, A=>nx14769);
   ix18260 : buf16 port map ( Y=>nx17809, A=>nx15358);
   ix18261 : buf16 port map ( Y=>nx17810, A=>nx15358);
   ix18262 : buf16 port map ( Y=>nx17811, A=>nx15829);
   ix18263 : buf16 port map ( Y=>nx17812, A=>nx15829);
   ix18264 : buf16 port map ( Y=>nx17813, A=>nx15829);
   ix18265 : buf16 port map ( Y=>nx17814, A=>write_base_data_out_2);
   ix18266 : buf16 port map ( Y=>nx17815, A=>write_base_data_out_2);
   ix18267 : buf16 port map ( Y=>nx17816, A=>nx15956);
   ix18268 : buf16 port map ( Y=>nx17817, A=>nx15956);
   ix18269 : buf16 port map ( Y=>nx17818, A=>write_base_data_out_4);
   ix18270 : buf16 port map ( Y=>nx17819, A=>write_base_data_out_4);
   ix18271 : buf16 port map ( Y=>nx17820, A=>nx16078);
   ix18272 : buf16 port map ( Y=>nx17821, A=>nx16078);
   ix18273 : buf16 port map ( Y=>nx17822, A=>write_base_data_out_6);
   ix18274 : buf16 port map ( Y=>nx17823, A=>write_base_data_out_6);
   ix18275 : buf16 port map ( Y=>nx17824, A=>write_base_data_out_8);
   ix18276 : buf16 port map ( Y=>nx17825, A=>write_base_data_out_8);
   ix18277 : buf16 port map ( Y=>nx17826, A=>nx17021);
   ix18278 : buf16 port map ( Y=>nx17827, A=>nx17021);
   ix18279 : buf16 port map ( Y=>nx17828, A=>nx3692);
   ix18280 : buf16 port map ( Y=>nx17829, A=>nx3692);
   ix18281 : buf16 port map ( Y=>nx17830, A=>write_base_data_out_10);
   ix18282 : buf16 port map ( Y=>nx17831, A=>write_base_data_out_10);
   ix18283 : buf16 port map ( Y=>nx17832, A=>nx16434);
   ix18284 : buf16 port map ( Y=>nx17833, A=>nx16434);
   ix18285 : buf16 port map ( Y=>nx17834, A=>write_base_data_out_12);
   ix18286 : buf16 port map ( Y=>nx17835, A=>write_base_data_out_12);
   ix18287 : buf16 port map ( Y=>nx17836, A=>nx16555);
   ix18288 : buf16 port map ( Y=>nx17837, A=>nx16555);
   ix18289 : buf16 port map ( Y=>nx17838, A=>nx16622);
   ix18290 : buf16 port map ( Y=>nx17839, A=>nx16622);
   ix18291 : buf16 port map ( Y=>nx17840, A=>nx16622);
   ix18292 : buf02 port map ( Y=>nx18293, A=>nx15805);
   ix18294 : buf02 port map ( Y=>nx18295, A=>nx15974);
   ix18296 : buf02 port map ( Y=>nx18297, A=>nx15974);
   ix18298 : buf02 port map ( Y=>nx18299, A=>nx4420);
   ix18300 : buf02 port map ( Y=>nx18301, A=>nx17443);
   ix18302 : buf02 port map ( Y=>nx18303, A=>nx16487);
   ix18304 : buf02 port map ( Y=>nx18305, A=>nx17718);
   ix18306 : buf02 port map ( Y=>nx18307, A=>nx17763);
end Mixed ;

