
-- 
-- Definition of  Ram
-- 
--      Fri Mar 22 20:16:45 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use dcnn.adk_components.all;

entity Ram is
   port (
      clk : IN std_logic ;
      read_in : IN std_logic ;
      write_out : IN std_logic ;
      address : IN std_logic_vector (7 DOWNTO 0) ;
      data_in : IN std_logic_vector (15 DOWNTO 0) ;
      data_out : OUT std_logic_vector (15 DOWNTO 0)) ;
end Ram ;

architecture Behavioral of Ram is
   signal nx2, nx8, nx14, nx18, nx42, nx44, nx48, nx52, nx72, nx90, nx96, 
      nx98, nx116, nx122, nx126, nx128, nx150, nx158, nx174, nx178, nx192, 
      nx210, nx218, nx226, nx260, nx264, nx278, nx296, nx338, nx358, nx378, 
      nx404, nx424, nx426, nx444, nx450, nx452, nx456, nx470, nx476, 
      modgen_ram_ix74_a_28_dup_1191, nx560, modgen_ram_ix74_a_12_dup_1207, 
      nx598, nx612, nx630, nx634, nx656, nx672, nx694, nx698, nx714, nx726, 
      nx778, nx780, nx806, nx860, nx888, nx922, nx942, nx968, nx1002, nx1004, 
      nx1026, nx1086, nx1088, nx1092, nx1106, nx1124, nx1166, nx1184, nx1188, 
      nx1202, nx1248, nx1286, nx1292, nx1310, nx1330, nx1364, nx1392, nx1400, 
      nx1408, nx1430, nx1438, nx1446, nx1470, nx1478, nx1486, nx1508, nx1526, 
      nx1550, nx1558, nx1566, modgen_ram_ix74_a_28_dup_1126, 
      modgen_ram_ix74_a_12_dup_1142, nx1636, nx1644, nx1648, nx1666, nx1684, 
      nx1718, nx1788, nx1826, nx1868, nx1876, nx1884, nx1906, nx1914, nx1922, 
      nx1946, nx1964, nx2002, nx2030, nx2038, nx2046, nx2068, nx2076, nx2084, 
      nx2108, nx2116, nx2124, nx2146, nx2164, nx2188, nx2196, nx2204, 
      modgen_ram_ix74_a_28_dup_1060, modgen_ram_ix74_a_12_dup_1076, nx2274, 
      nx2282, nx2286, nx2304, nx2322, nx2356, nx2426, nx2464, nx2506, nx2514, 
      nx2522, nx2544, nx2552, nx2560, nx2584, nx2602, nx2640, nx2668, nx2676, 
      nx2684, nx2706, nx2714, nx2722, nx2746, nx2754, nx2762, nx2784, nx2802, 
      nx2826, nx2834, nx2842, nx2864, nx2872, nx2880, 
      modgen_ram_ix74_a_28_dup_995, modgen_ram_ix74_a_12_dup_1011, nx2912, 
      nx2920, nx2924, nx2942, nx2960, nx2986, nx2994, nx3024, nx3064, nx3102, 
      nx3144, nx3152, nx3160, nx3182, nx3190, nx3198, nx3222, nx3240, nx3260, 
      nx3278, nx3306, nx3314, nx3322, nx3344, nx3352, nx3360, nx3384, nx3392, 
      nx3400, nx3422, nx3440, nx3464, nx3472, nx3480, nx3502, nx3510, nx3518, 
      modgen_ram_ix74_a_28_dup_930, modgen_ram_ix74_a_12_dup_946, nx3550, 
      nx3558, nx3562, nx3580, nx3598, nx3624, nx3632, nx3662, nx3702, nx3740, 
      nx3782, nx3790, nx3798, nx3820, nx3828, nx3836, nx3860, nx3878, nx3898, 
      nx3916, nx3944, nx3952, nx3960, nx3982, nx3990, nx3998, nx4022, nx4030, 
      nx4038, nx4060, nx4078, nx4102, nx4110, nx4118, nx4140, nx4148, nx4156, 
      modgen_ram_ix74_a_28_dup_865, modgen_ram_ix74_a_12_dup_881, nx4188, 
      nx4196, nx4200, nx4218, nx4236, nx4262, nx4270, nx4300, nx4340, nx4378, 
      nx4420, nx4428, nx4436, nx4458, nx4466, nx4474, nx4498, nx4516, nx4536, 
      nx4554, nx4582, nx4590, nx4598, nx4620, nx4628, nx4636, nx4660, nx4668, 
      nx4676, nx4698, nx4716, nx4748, nx4756, nx4778, nx4786, nx4794, 
      modgen_ram_ix74_a_28_dup_799, modgen_ram_ix74_a_12_dup_815, nx4826, 
      nx4834, nx4838, nx4856, nx4874, nx4900, nx4908, nx4938, nx4978, nx5016, 
      nx5058, nx5066, nx5074, nx5096, nx5104, nx5112, nx5136, nx5154, nx5174, 
      nx5192, nx5220, nx5228, nx5236, nx5258, nx5266, nx5274, nx5298, nx5306, 
      nx5314, nx5336, nx5354, nx5378, nx5386, nx5394, nx5416, nx5424, nx5432, 
      modgen_ram_ix74_a_28_dup_734, modgen_ram_ix74_a_12_dup_750, nx5464, 
      nx5472, nx5476, nx5494, nx5512, nx5538, nx5546, nx5576, nx5616, nx5654, 
      nx5696, nx5704, nx5712, nx5734, nx5742, nx5750, nx5774, nx5792, nx5812, 
      nx5830, nx5858, nx5866, nx5874, nx5896, nx5904, nx5912, nx5936, nx5944, 
      nx5952, nx5974, nx5992, nx6016, nx6024, nx6032, nx6054, nx6062, nx6070, 
      modgen_ram_ix74_a_28_dup_669, modgen_ram_ix74_a_12_dup_685, nx6102, 
      nx6110, nx6114, nx6132, nx6150, nx6176, nx6184, nx6214, nx6254, nx6292, 
      nx6334, nx6342, nx6350, nx6372, nx6380, nx6388, nx6412, nx6430, nx6450, 
      nx6468, nx6496, nx6504, nx6512, nx6534, nx6542, nx6550, nx6574, nx6582, 
      nx6590, nx6612, nx6630, nx6654, nx6662, nx6670, nx6692, nx6700, nx6708, 
      modgen_ram_ix74_a_28_dup_604, modgen_ram_ix74_a_12_dup_620, nx6740, 
      nx6748, nx6752, nx6770, nx6788, nx6814, nx6822, nx6852, nx6892, nx6930, 
      nx6972, nx6980, nx6988, nx7010, nx7018, nx7026, nx7050, nx7068, nx7088, 
      nx7106, nx7134, nx7142, nx7150, nx7172, nx7180, nx7188, nx7212, nx7220, 
      nx7228, nx7250, nx7268, nx7292, nx7300, nx7308, nx7330, nx7338, nx7346, 
      modgen_ram_ix74_a_28_dup_538, modgen_ram_ix74_a_12_dup_554, nx7378, 
      nx7386, nx7390, nx7408, nx7426, nx7452, nx7460, nx7490, nx7530, nx7568, 
      nx7610, nx7618, nx7626, nx7648, nx7656, nx7664, nx7688, nx7706, nx7726, 
      nx7744, nx7772, nx7780, nx7788, nx7810, nx7818, nx7826, nx7850, nx7858, 
      nx7866, nx7888, nx7906, nx7930, nx7938, nx7946, nx7968, nx7976, nx7984, 
      modgen_ram_ix74_a_28_dup_473, modgen_ram_ix74_a_12_dup_489, nx8016, 
      nx8024, nx8028, nx8046, nx8064, nx8090, nx8098, nx8128, nx8168, nx8206, 
      nx8248, nx8256, nx8264, nx8286, nx8294, nx8302, nx8326, nx8344, nx8364, 
      nx8382, nx8410, nx8418, nx8426, nx8448, nx8456, nx8464, nx8488, nx8496, 
      nx8504, nx8526, nx8544, nx8568, nx8576, nx8584, nx8606, nx8614, nx8622, 
      modgen_ram_ix74_a_28_dup_408, modgen_ram_ix74_a_12_dup_424, nx8654, 
      nx8662, nx8666, nx8684, nx8702, nx8728, nx8736, nx8766, nx8806, nx8844, 
      nx8886, nx8894, nx8902, nx8924, nx8932, nx8940, nx8964, nx8982, nx9002, 
      nx9020, nx9048, nx9056, nx9064, nx9086, nx9094, nx9102, nx9126, nx9134, 
      nx9142, nx9164, nx9182, nx9206, nx9214, nx9222, 
      modgen_ram_ix74_a_28_dup_342, modgen_ram_ix74_a_12_dup_358, nx9292, 
      nx9300, nx9304, nx9322, nx9340, nx9374, nx9444, nx9482, nx9524, nx9532, 
      nx9540, nx9562, nx9570, nx9578, nx9602, nx9620, nx9658, nx9686, nx9694, 
      nx9702, nx9724, nx9732, nx9740, nx9764, nx9772, nx9780, nx9802, nx9820, 
      nx9844, nx9852, nx9860, nx9882, nx9890, nx9898, 
      modgen_ram_ix74_a_28_dup_277, modgen_ram_ix74_a_12_dup_293, nx9930, 
      nx9938, nx9942, nx9960, nx9978, nx10004, nx10012, nx10042, nx10082, 
      nx10120, nx10162, nx10170, nx10178, nx10200, nx10208, nx10216, nx10240, 
      nx10258, nx10278, nx10296, nx10324, nx10332, nx10340, nx10362, nx10370, 
      nx10378, nx10402, nx10410, nx10418, nx10440, nx10458, nx10482, nx10490, 
      nx10498, nx10520, nx10528, nx10536, modgen_ram_ix74_a_28, 
      modgen_ram_ix74_a_12, nx10568, nx10576, nx10580, nx10598, nx10616, 
      nx10642, nx10650, nx10680, nx10720, nx10758, nx10800, nx10808, nx10816, 
      nx10838, nx10846, nx10854, nx10878, nx10896, nx10916, nx10934, nx249, 
      nx259, nx269, nx279, nx289, nx299, nx309, nx319, nx329, nx339, nx349, 
      nx359, nx369, nx379, nx389, nx399, nx409, nx419, nx429, nx439, nx449, 
      nx459, nx469, nx479, nx489, nx499, nx509, nx519, nx529, nx539, nx549, 
      nx559, nx569, nx579, nx589, nx599, nx609, nx619, nx629, nx639, nx649, 
      nx659, nx669, nx679, nx689, nx699, nx709, nx719, nx729, nx739, nx749, 
      nx759, nx769, nx779, nx789, nx799, nx809, nx819, nx829, nx839, nx849, 
      nx859, nx869, nx879, nx889, nx899, nx909, nx919, nx929, nx939, nx949, 
      nx959, nx969, nx979, nx989, nx999, nx1009, nx1019, nx1029, nx1039, 
      nx1049, nx1059, nx1069, nx1079, nx1089, nx1099, nx1109, nx1119, nx1129, 
      nx1139, nx1149, nx1159, nx1169, nx1179, nx1189, nx1199, nx1209, nx1219, 
      nx1229, nx1239, nx1249, nx1259, nx1269, nx1279, nx1289, nx1299, nx1309, 
      nx1319, nx1329, nx1339, nx1349, nx1359, nx1369, nx1379, nx1389, nx1399, 
      nx1409, nx1419, nx1429, nx1439, nx1449, nx1459, nx1469, nx1479, nx1489, 
      nx1499, nx1509, nx1519, nx1529, nx1539, nx1549, nx1559, nx1569, nx1579, 
      nx1589, nx1599, nx1609, nx1619, nx1629, nx1639, nx1649, nx1659, nx1669, 
      nx1679, nx1689, nx1699, nx1709, nx1719, nx1729, nx1739, nx1749, nx1759, 
      nx1769, nx1779, nx1789, nx1799, nx1809, nx1819, nx1829, nx1839, nx1849, 
      nx1859, nx1869, nx1879, nx1889, nx1899, nx1909, nx1919, nx1929, nx1939, 
      nx1949, nx1959, nx1969, nx1979, nx1989, nx1999, nx2009, nx2019, nx2029, 
      nx2039, nx2049, nx2059, nx2069, nx2079, nx2089, nx2099, nx2109, nx2119, 
      nx2129, nx2139, nx2149, nx2159, nx2169, nx2179, nx2189, nx2199, nx2209, 
      nx2219, nx2229, nx2239, nx2249, nx2259, nx2269, nx2279, nx2289, nx2299, 
      nx2309, nx2319, nx2329, nx2339, nx2349, nx2359, nx2369, nx2379, nx2389, 
      nx2399, nx2409, nx2419, nx2429, nx2439, nx2449, nx2459, nx2469, nx2479, 
      nx2489, nx2499, nx2509, nx2519, nx2529, nx2539, nx2549, nx2559, nx2569, 
      nx2579, nx2589, nx2599, nx2609, nx2619, nx2629, nx2639, nx2649, nx2659, 
      nx2669, nx2679, nx2689, nx2699, nx2709, nx2719, nx2729, nx2739, nx2749, 
      nx2759, nx2769, nx2779, nx2789, nx2799, nx2809, nx2819, nx2829, nx2839, 
      nx2849, nx2859, nx2869, nx2879, nx2889, nx2899, nx2909, nx2919, nx2929, 
      nx2939, nx2949, nx2959, nx2969, nx2979, nx2989, nx2999, nx3009, nx3019, 
      nx3029, nx3039, nx3049, nx3059, nx3069, nx3079, nx3089, nx3099, nx3109, 
      nx3119, nx3129, nx3139, nx3149, nx3159, nx3169, nx3179, nx3189, nx3199, 
      nx3209, nx3219, nx3229, nx3239, nx3249, nx3259, nx3269, nx3279, nx3289, 
      nx3299, nx3309, nx3319, nx3329, nx3339, nx3349, nx3359, nx3369, nx3379, 
      nx3389, nx3399, nx3409, nx3419, nx3429, nx3439, nx3449, nx3459, nx3469, 
      nx3479, nx3489, nx3499, nx3509, nx3519, nx3529, nx3539, nx3549, nx3559, 
      nx3569, nx3579, nx3589, nx3599, nx3609, nx3619, nx3629, nx3639, nx3649, 
      nx3659, nx3669, nx3679, nx3689, nx3699, nx3709, nx3719, nx3729, nx3739, 
      nx3749, nx3759, nx3769, nx3779, nx3789, nx3799, nx3809, nx3819, nx3829, 
      nx3839, nx3849, nx3859, nx3869, nx3879, nx3889, nx3899, nx3909, nx3919, 
      nx3929, nx3939, nx3949, nx3959, nx3969, nx3979, nx3989, nx3999, nx4009, 
      nx4019, nx4029, nx4039, nx4049, nx4059, nx4069, nx4079, nx4089, nx4099, 
      nx4109, nx4119, nx4129, nx4139, nx4149, nx4159, nx4169, nx4179, nx4189, 
      nx4199, nx4209, nx4219, nx4229, nx4239, nx4249, nx4259, nx4269, nx4279, 
      nx4289, nx4299, nx4309, nx4319, nx4329, nx4339, nx4349, nx4359, nx4369, 
      nx4379, nx4389, nx4399, nx4409, nx4419, nx4429, nx4439, nx4449, nx4459, 
      nx4469, nx4479, nx4489, nx4499, nx4509, nx4519, nx4529, nx4539, nx4549, 
      nx4559, nx4569, nx4579, nx4589, nx4599, nx4609, nx4619, nx4629, nx4639, 
      nx4649, nx4659, nx4669, nx4679, nx4689, nx4699, nx4709, nx4719, nx4729, 
      nx4739, nx4749, nx4759, nx4769, nx4779, nx4789, nx4799, nx4809, nx4819, 
      nx4829, nx4839, nx4849, nx4859, nx4869, nx4879, nx4889, nx4899, nx4909, 
      nx4919, nx4929, nx4939, nx4949, nx4959, nx4969, nx4979, nx4989, nx4999, 
      nx5009, nx5019, nx5029, nx5039, nx5049, nx5059, nx5069, nx5079, nx5089, 
      nx5099, nx5109, nx5119, nx5129, nx5139, nx5149, nx5159, nx5169, nx5179, 
      nx5189, nx5199, nx5209, nx5219, nx5229, nx5239, nx5249, nx5259, nx5269, 
      nx5279, nx5289, nx5299, nx5309, nx5319, nx5329, nx5339, nx5349, nx5359, 
      nx5369, nx5379, nx5389, nx5399, nx5409, nx5419, nx5429, nx5439, nx5449, 
      nx5459, nx5469, nx5479, nx5489, nx5499, nx5509, nx5519, nx5529, nx5539, 
      nx5549, nx5559, nx5569, nx5579, nx5589, nx5599, nx5609, nx5619, nx5629, 
      nx5639, nx5649, nx5659, nx5669, nx5679, nx5689, nx5699, nx5709, nx5719, 
      nx5729, nx5739, nx5749, nx5759, nx5769, nx5779, nx5789, nx5799, nx5809, 
      nx5819, nx5829, nx5839, nx5849, nx5859, nx5869, nx5879, nx5889, nx5899, 
      nx5909, nx5919, nx5929, nx5939, nx5949, nx5959, nx5969, nx5979, nx5989, 
      nx5999, nx6009, nx6019, nx6029, nx6039, nx6049, nx6059, nx6069, nx6079, 
      nx6089, nx6099, nx6109, nx6119, nx6129, nx6139, nx6149, nx6159, nx6169, 
      nx6179, nx6189, nx6199, nx6209, nx6219, nx6229, nx6239, nx6249, nx6259, 
      nx6269, nx6279, nx6289, nx6299, nx6309, nx6319, nx6329, nx6339, nx6349, 
      nx6359, nx6369, nx6379, nx6389, nx6399, nx6409, nx6419, nx6429, nx6439, 
      nx6449, nx6459, nx6469, nx6479, nx6489, nx6499, nx6509, nx6519, nx6529, 
      nx6539, nx6549, nx6559, nx6569, nx6579, nx6589, nx6599, nx6609, nx6619, 
      nx6629, nx6639, nx6649, nx6659, nx6669, nx6679, nx6689, nx6699, nx6709, 
      nx6719, nx6729, nx6739, nx6749, nx6759, nx6769, nx6779, nx6789, nx6799, 
      nx6809, nx6819, nx6829, nx6839, nx6849, nx6859, nx6869, nx6879, nx6889, 
      nx6899, nx6909, nx6919, nx6929, nx6939, nx6949, nx6959, nx6969, nx6979, 
      nx6989, nx6999, nx7009, nx7019, nx7029, nx7039, nx7049, nx7059, nx7069, 
      nx7079, nx7089, nx7099, nx7109, nx7119, nx7129, nx7139, nx7149, nx7159, 
      nx7169, nx7179, nx7189, nx7199, nx7209, nx7219, nx7229, nx7239, nx7249, 
      nx7259, nx7269, nx7279, nx7289, nx7299, nx7309, nx7319, nx7329, nx7339, 
      nx7349, nx7359, nx7369, nx7379, nx7389, nx7399, nx7409, nx7419, nx7429, 
      nx7439, nx7449, nx7459, nx7469, nx7479, nx7489, nx7499, nx7509, nx7519, 
      nx7529, nx7539, nx7549, nx7559, nx7569, nx7579, nx7589, nx7599, nx7609, 
      nx7619, nx7629, nx7639, nx7649, nx7659, nx7669, nx7679, nx7689, nx7699, 
      nx7709, nx7719, nx7729, nx7739, nx7749, nx7759, nx7769, nx7779, nx7789, 
      nx7799, nx7809, nx7819, nx7829, nx7839, nx7849, nx7859, nx7869, nx7879, 
      nx7889, nx7899, nx7909, nx7919, nx7929, nx7939, nx7949, nx7959, nx7969, 
      nx7979, nx7989, nx7999, nx8009, nx8019, nx8029, nx8039, nx8049, nx8059, 
      nx8069, nx8079, nx8089, nx8099, nx8109, nx8119, nx8129, nx8139, nx8149, 
      nx8159, nx8169, nx8179, nx8189, nx8199, nx8209, nx8219, nx8229, nx8239, 
      nx8249, nx8259, nx8269, nx8279, nx8289, nx8299, nx8309, nx8319, nx8329, 
      nx8339, nx8349, nx8359, nx8369, nx8379, nx8389, nx8399, nx8409, nx8419, 
      nx8429, nx8439, nx8449, nx8459, nx8469, nx8479, nx8489, nx8499, nx8509, 
      nx8519, nx8529, nx8539, nx8549, nx8559, nx8569, nx8579, nx8589, nx8599, 
      nx8609, nx8619, nx8629, nx8639, nx8649, nx8659, nx8669, nx8679, nx8689, 
      nx8699, nx8709, nx8719, nx8729, nx8739, nx8749, nx8759, nx8769, nx8779, 
      nx8789, nx8799, nx8809, nx8819, nx8829, nx8839, nx8849, nx8859, nx8869, 
      nx8879, nx8889, nx8899, nx8909, nx8919, nx8929, nx8939, nx8949, nx8959, 
      nx8969, nx8979, nx8989, nx8999, nx9009, nx9019, nx9029, nx9039, nx9049, 
      nx9059, nx9069, nx9079, nx9089, nx9099, nx9109, nx9119, nx9129, nx9139, 
      nx9149, nx9159, nx9169, nx9179, nx9189, nx9199, nx9209, nx9219, nx9229, 
      nx9239, nx9249, nx9259, nx9269, nx9279, nx9289, nx9299, nx9309, nx9319, 
      nx9329, nx9339, nx9349, nx9359, nx9369, nx9379, nx9389, nx9399, nx9409, 
      nx9419, nx9429, nx9439, nx9449, nx9459, nx9469, nx9479, nx9489, nx9499, 
      nx9509, nx9519, nx9529, nx9539, nx9549, nx9559, nx9569, nx9579, nx9589, 
      nx9599, nx9609, nx9619, nx9629, nx9639, nx9649, nx9659, nx9669, nx9679, 
      nx9689, nx9699, nx9709, nx9719, nx9729, nx9739, nx9749, nx9759, nx9769, 
      nx9779, nx9789, nx9799, nx9809, nx9819, nx9829, nx9839, nx9849, nx9859, 
      nx9869, nx9879, nx9889, nx9899, nx9909, nx9919, nx9929, nx9939, nx9949, 
      nx9959, nx9969, nx9979, nx9989, nx9999, nx10009, nx10019, nx10029, 
      nx10039, nx10049, nx10059, nx10069, nx10079, nx10089, nx10099, nx10109, 
      nx10119, nx10129, nx10139, nx10149, nx10159, nx10169, nx10179, nx10189, 
      nx10199, nx10209, nx10219, nx10229, nx10239, nx10249, nx10259, nx10269, 
      nx10279, nx10289, nx10299, nx10309, nx10319, nx10329, nx10339, nx10349, 
      nx10359, nx10369, nx10379, nx10389, nx10399, nx10409, nx10419, nx10429, 
      nx10439, nx10449, nx10459, nx10469, nx10479, nx10497, nx10503, nx10505, 
      nx10507, nx10514, nx10519, nx10521, nx10527, nx10529, nx10534, nx10537, 
      nx10541, nx10543, nx10548, nx10555, nx10557, nx10559, nx10567, nx10571, 
      nx10574, nx10577, nx10579, nx10584, nx10587, nx10589, nx10592, nx10595, 
      nx10599, nx10603, nx10607, nx10611, nx10613, nx10615, nx10619, nx10625, 
      nx10629, nx10633, nx10637, nx10641, nx10643, nx10645, nx10648, nx10651, 
      nx10654, nx10657, nx10659, nx10663, nx10666, nx10671, nx10674, nx10677, 
      nx10679, nx10681, nx10684, nx10686, nx10692, nx10699, nx10703, nx10706, 
      nx10711, nx10713, nx10716, nx10719, nx10724, nx10727, nx10731, nx10734, 
      nx10737, nx10744, nx10749, nx10751, nx10754, nx10757, nx10762, nx10765, 
      nx10769, nx10772, nx10775, nx10783, nx10787, nx10789, nx10793, nx10795, 
      nx10801, nx10804, nx10807, nx10811, nx10813, nx10817, nx10823, nx10825, 
      nx10829, nx10831, nx10841, nx10844, nx10847, nx10850, nx10852, nx10857, 
      nx10861, nx10866, nx10869, nx10872, nx10874, nx10877, nx10881, nx10884, 
      nx10887, nx10889, nx10893, nx10899, nx10903, nx10907, nx10909, nx10913, 
      nx10922, nx10928, nx10931, nx10935, nx10939, nx10941, nx10943, nx10951, 
      nx10954, nx10959, nx10962, nx10965, nx10968, nx10970, nx10972, nx10975, 
      nx10977, nx10983, nx10986, nx10988, nx10990, nx10992, nx10995, nx10997, 
      nx11000, nx11003, nx11007, nx11010, nx11012, nx11016, nx11019, nx11022, 
      nx11026, nx11032, nx11035, nx11037, nx11039, nx11041, nx11048, nx11051, 
      nx11054, nx11056, nx11059, nx11064, nx11070, nx11073, nx11075, nx11077, 
      nx11080, nx11083, nx11086, nx11089, nx11092, nx11095, nx11097, nx11099, 
      nx11102, nx11104, nx11113, nx11118, nx11122, nx11125, nx11128, nx11131, 
      nx11134, nx11138, nx11141, nx11144, nx11147, nx11151, nx11155, nx11158, 
      nx11161, nx11164, nx11168, nx11172, nx11175, nx11182, nx11186, nx11190, 
      nx11193, nx11199, nx11203, nx11207, nx11210, nx11216, nx11220, nx11224, 
      nx11227, nx11233, nx11237, nx11241, nx11244, nx11254, nx11257, nx11261, 
      nx11264, nx11268, nx11271, nx11275, nx11278, nx11282, nx11284, nx11288, 
      nx11293, nx11297, nx11301, nx11304, nx11307, nx11310, nx11314, nx11318, 
      nx11321, nx11328, nx11331, nx11335, nx11338, nx11341, nx11344, nx11348, 
      nx11352, nx11355, nx11358, nx11361, nx11365, nx11369, nx11372, nx11375, 
      nx11378, nx11382, nx11386, nx11389, nx11399, nx11404, nx11408, nx11411, 
      nx11414, nx11417, nx11420, nx11424, nx11427, nx11430, nx11433, nx11437, 
      nx11441, nx11444, nx11447, nx11450, nx11454, nx11458, nx11461, nx11468, 
      nx11472, nx11476, nx11479, nx11485, nx11489, nx11493, nx11496, nx11502, 
      nx11506, nx11510, nx11513, nx11519, nx11523, nx11527, nx11530, nx11540, 
      nx11543, nx11547, nx11550, nx11554, nx11557, nx11561, nx11564, nx11568, 
      nx11570, nx11574, nx11579, nx11583, nx11587, nx11590, nx11593, nx11596, 
      nx11600, nx11604, nx11607, nx11614, nx11617, nx11621, nx11624, nx11627, 
      nx11630, nx11634, nx11638, nx11641, nx11644, nx11647, nx11651, nx11655, 
      nx11658, nx11661, nx11664, nx11668, nx11672, nx11675, nx11685, nx11690, 
      nx11694, nx11697, nx11700, nx11703, nx11706, nx11710, nx11713, nx11716, 
      nx11719, nx11723, nx11727, nx11730, nx11733, nx11736, nx11740, nx11744, 
      nx11747, nx11754, nx11758, nx11762, nx11765, nx11771, nx11775, nx11779, 
      nx11782, nx11788, nx11792, nx11796, nx11799, nx11805, nx11809, nx11813, 
      nx11816, nx11826, nx11829, nx11833, nx11836, nx11840, nx11843, nx11847, 
      nx11850, nx11854, nx11856, nx11860, nx11862, nx11865, nx11869, nx11873, 
      nx11876, nx11879, nx11882, nx11886, nx11890, nx11893, nx11900, nx11903, 
      nx11907, nx11910, nx11913, nx11916, nx11920, nx11924, nx11927, nx11930, 
      nx11933, nx11937, nx11941, nx11944, nx11947, nx11950, nx11954, nx11958, 
      nx11961, nx11971, nx11976, nx11980, nx11983, nx11986, nx11989, nx11992, 
      nx11996, nx11999, nx12002, nx12005, nx12009, nx12013, nx12016, nx12019, 
      nx12022, nx12026, nx12030, nx12033, nx12040, nx12044, nx12048, nx12051, 
      nx12057, nx12061, nx12065, nx12068, nx12074, nx12078, nx12082, nx12085, 
      nx12091, nx12095, nx12099, nx12102, nx12112, nx12115, nx12119, nx12122, 
      nx12126, nx12129, nx12133, nx12136, nx12140, nx12142, nx12146, nx12148, 
      nx12151, nx12155, nx12159, nx12162, nx12165, nx12168, nx12172, nx12176, 
      nx12179, nx12186, nx12189, nx12193, nx12196, nx12199, nx12202, nx12206, 
      nx12210, nx12213, nx12216, nx12219, nx12223, nx12227, nx12230, nx12233, 
      nx12236, nx12240, nx12244, nx12247, nx12257, nx12262, nx12266, nx12269, 
      nx12272, nx12275, nx12278, nx12282, nx12285, nx12288, nx12291, nx12295, 
      nx12299, nx12302, nx12305, nx12308, nx12312, nx12316, nx12319, nx12326, 
      nx12330, nx12334, nx12337, nx12343, nx12347, nx12351, nx12354, nx12360, 
      nx12364, nx12368, nx12371, nx12377, nx12381, nx12385, nx12388, nx12398, 
      nx12401, nx12405, nx12408, nx12412, nx12415, nx12419, nx12422, nx12426, 
      nx12428, nx12432, nx12434, nx12437, nx12441, nx12445, nx12448, nx12451, 
      nx12454, nx12458, nx12462, nx12465, nx12472, nx12475, nx12479, nx12482, 
      nx12485, nx12488, nx12492, nx12496, nx12499, nx12502, nx12505, nx12509, 
      nx12513, nx12516, nx12519, nx12522, nx12526, nx12530, nx12533, nx12543, 
      nx12548, nx12552, nx12555, nx12558, nx12561, nx12564, nx12568, nx12571, 
      nx12574, nx12577, nx12581, nx12585, nx12588, nx12591, nx12594, nx12598, 
      nx12602, nx12605, nx12612, nx12616, nx12620, nx12623, nx12629, nx12633, 
      nx12637, nx12640, nx12646, nx12650, nx12654, nx12657, nx12663, nx12667, 
      nx12671, nx12674, nx12684, nx12687, nx12691, nx12694, nx12698, nx12701, 
      nx12705, nx12708, nx12712, nx12714, nx12718, nx12720, nx12723, nx12727, 
      nx12731, nx12734, nx12740, nx12744, nx12748, nx12751, nx12758, nx12761, 
      nx12765, nx12768, nx12771, nx12774, nx12778, nx12782, nx12785, nx12788, 
      nx12791, nx12795, nx12799, nx12802, nx12805, nx12808, nx12812, nx12816, 
      nx12819, nx12829, nx12834, nx12838, nx12841, nx12844, nx12847, nx12850, 
      nx12854, nx12857, nx12860, nx12863, nx12867, nx12871, nx12874, nx12877, 
      nx12880, nx12884, nx12888, nx12891, nx12898, nx12902, nx12906, nx12909, 
      nx12915, nx12919, nx12923, nx12926, nx12932, nx12936, nx12940, nx12943, 
      nx12949, nx12953, nx12957, nx12960, nx12970, nx12973, nx12977, nx12980, 
      nx12984, nx12987, nx12991, nx12994, nx12998, nx13000, nx13004, nx13006, 
      nx13009, nx13013, nx13017, nx13020, nx13023, nx13026, nx13030, nx13034, 
      nx13037, nx13044, nx13047, nx13051, nx13054, nx13057, nx13060, nx13064, 
      nx13068, nx13071, nx13074, nx13077, nx13081, nx13085, nx13088, nx13091, 
      nx13094, nx13098, nx13102, nx13105, nx13115, nx13120, nx13124, nx13127, 
      nx13130, nx13133, nx13136, nx13140, nx13143, nx13146, nx13149, nx13153, 
      nx13157, nx13160, nx13163, nx13166, nx13170, nx13174, nx13177, nx13184, 
      nx13188, nx13192, nx13195, nx13201, nx13205, nx13209, nx13212, nx13218, 
      nx13222, nx13226, nx13229, nx13235, nx13239, nx13243, nx13246, nx13256, 
      nx13259, nx13263, nx13266, nx13270, nx13273, nx13277, nx13280, nx13284, 
      nx13286, nx13290, nx13292, nx13295, nx13299, nx13303, nx13306, nx13309, 
      nx13312, nx13316, nx13320, nx13323, nx13330, nx13333, nx13337, nx13340, 
      nx13343, nx13346, nx13350, nx13354, nx13357, nx13360, nx13363, nx13367, 
      nx13371, nx13374, nx13377, nx13380, nx13384, nx13388, nx13391, nx13401, 
      nx13406, nx13410, nx13413, nx13416, nx13419, nx13422, nx13426, nx13429, 
      nx13432, nx13435, nx13439, nx13443, nx13446, nx13449, nx13452, nx13456, 
      nx13460, nx13463, nx13470, nx13474, nx13478, nx13481, nx13487, nx13491, 
      nx13495, nx13498, nx13504, nx13508, nx13512, nx13515, nx13521, nx13525, 
      nx13529, nx13532, nx13542, nx13545, nx13549, nx13552, nx13556, nx13559, 
      nx13563, nx13566, nx13570, nx13572, nx13576, nx13578, nx13581, nx13585, 
      nx13589, nx13592, nx13595, nx13598, nx13602, nx13606, nx13609, nx13616, 
      nx13619, nx13623, nx13626, nx13629, nx13632, nx13636, nx13640, nx13643, 
      nx13646, nx13649, nx13653, nx13657, nx13660, nx13663, nx13666, nx13670, 
      nx13674, nx13677, nx13687, nx13692, nx13696, nx13699, nx13702, nx13705, 
      nx13708, nx13712, nx13715, nx13718, nx13721, nx13725, nx13729, nx13732, 
      nx13735, nx13738, nx13742, nx13746, nx13749, nx13756, nx13760, nx13764, 
      nx13767, nx13773, nx13777, nx13781, nx13784, nx13790, nx13794, nx13798, 
      nx13801, nx13807, nx13811, nx13815, nx13818, nx13828, nx13831, nx13835, 
      nx13838, nx13842, nx13845, nx13849, nx13852, nx13856, nx13858, nx13862, 
      nx13864, nx13867, nx13871, nx13875, nx13878, nx13881, nx13884, nx13888, 
      nx13892, nx13895, nx13902, nx13905, nx13909, nx13912, nx13915, nx13918, 
      nx13922, nx13926, nx13929, nx13932, nx13935, nx13939, nx13943, nx13946, 
      nx13949, nx13952, nx13956, nx13960, nx13963, nx13973, nx13978, nx13982, 
      nx13985, nx13988, nx13991, nx13994, nx13998, nx14001, nx14004, nx14007, 
      nx14011, nx14015, nx14018, nx14021, nx14024, nx14028, nx14032, nx14035, 
      nx14042, nx14046, nx14050, nx14053, nx14059, nx14063, nx14067, nx14070, 
      nx14076, nx14080, nx14084, nx14087, nx14093, nx14097, nx14101, nx14104, 
      nx14114, nx14117, nx14121, nx14124, nx14128, nx14131, nx14135, nx14138, 
      nx14142, nx14144, nx14148, nx14150, nx14153, nx14157, nx14161, nx14164, 
      nx14167, nx14170, nx14174, nx14178, nx14181, nx14188, nx14191, nx14195, 
      nx14198, nx14201, nx14204, nx14208, nx14212, nx14215, nx14218, nx14221, 
      nx14225, nx14229, nx14232, nx14235, nx14238, nx14242, nx14246, nx14249, 
      nx14259, nx14264, nx14268, nx14271, nx14274, nx14277, nx14280, nx14284, 
      nx14287, nx14290, nx14293, nx14297, nx14301, nx14304, nx14307, nx14310, 
      nx14314, nx14318, nx14321, nx14328, nx14332, nx14336, nx14339, nx14345, 
      nx14349, nx14353, nx14356, nx14362, nx14366, nx14370, nx14373, nx14379, 
      nx14383, nx14387, nx14390, nx14400, nx14403, nx14407, nx14410, nx14414, 
      nx14417, nx14421, nx14424, nx14428, nx14430, nx14434, nx14436, nx14439, 
      nx14443, nx14447, nx14450, nx14453, nx14456, nx14460, nx14464, nx14467, 
      nx14474, nx14477, nx14481, nx14484, nx14487, nx14490, nx14494, nx14498, 
      nx14501, nx14504, nx14507, nx14511, nx14515, nx14518, nx14521, nx14524, 
      nx14528, nx14532, nx14535, nx14545, nx14550, nx14554, nx14557, nx14560, 
      nx14563, nx14566, nx14570, nx14573, nx14576, nx14579, nx14583, nx14587, 
      nx14590, nx14593, nx14596, nx14600, nx14604, nx14607, nx14614, nx14618, 
      nx14622, nx14625, nx14631, nx14635, nx14639, nx14642, nx14648, nx14652, 
      nx14656, nx14659, nx14665, nx14669, nx14673, nx14676, nx14686, nx14689, 
      nx14693, nx14696, nx14700, nx14703, nx14707, nx14710, nx14714, nx14716, 
      nx14720, nx14725, nx14729, nx14733, nx14736, nx14739, nx14742, nx14746, 
      nx14750, nx14753, nx14760, nx14763, nx14767, nx14770, nx14773, nx14776, 
      nx14780, nx14784, nx14787, nx14790, nx14793, nx14797, nx14801, nx14804, 
      nx14807, nx14810, nx14814, nx14818, nx14821, nx14831, nx14836, nx14840, 
      nx14843, nx14846, nx14849, nx14852, nx14856, nx14859, nx14862, nx14865, 
      nx14869, nx14873, nx14876, nx14879, nx14882, nx14886, nx14890, nx14893, 
      nx14900, nx14904, nx14908, nx14911, nx14917, nx14921, nx14925, nx14928, 
      nx14934, nx14938, nx14942, nx14945, nx14951, nx14955, nx14959, nx14962, 
      nx14972, nx14975, nx14979, nx14982, nx14986, nx14989, nx14993, nx14996, 
      nx15000, nx15002, nx15006, nx15008, nx15011, nx15015, nx15019, nx15022, 
      nx15025, nx15028, nx15032, nx15036, nx15039, nx15046, nx15049, nx15053, 
      nx15056, nx15059, nx15062, nx15066, nx15070, nx15073, nx15076, nx15079, 
      nx15083, nx15087, nx15090, nx15093, nx15096, nx15100, nx15104, nx15107, 
      nx15117, nx15122, nx15126, nx15129, nx15132, nx15135, nx15138, nx15142, 
      nx15145, nx15148, nx15151, nx15155, nx15159, nx15162, nx15165, nx15168, 
      nx15172, nx15176, nx15179, nx15186, nx15190, nx15194, nx15197, nx15203, 
      nx15207, nx15211, nx15214, nx15220, nx15224, nx15228, nx15231, nx15237, 
      nx15241, nx15245, nx15248, nx15258, nx15261, nx15265, nx15268, nx15272, 
      nx15275, nx15279, nx15282, nx15286, nx15288, nx15292, nx15294, nx15297, 
      nx15301, nx15305, nx15308, nx15311, nx15314, nx15318, nx15322, nx15325, 
      nx15332, nx15335, nx15339, nx15342, nx15345, nx15348, nx15352, nx15356, 
      nx15359, nx15362, nx15365, nx15369, nx15373, nx15376, nx15379, nx15382, 
      nx15386, nx15390, nx15393, nx15401, nx15403, nx15405, nx15407, nx15409, 
      nx15411, nx15413, nx15415, nx15417, nx15419, nx15421, nx15423, nx15425, 
      nx15427, nx15429, nx15431, nx15433, nx15435, nx15437, nx15439, nx15441, 
      nx15443, nx15445, nx15447, nx15449, nx15451, nx15453, nx15455, nx15457, 
      nx15459, nx15461, nx15463, nx15465, nx15467, nx15469, nx15471, nx15473, 
      nx15475, nx15477, nx15479, nx15481, nx15483, nx15485, nx15487, nx15489, 
      nx15491, nx15493, nx15495, nx15497, nx15499, nx15501, nx15503, nx15505, 
      nx15507, nx15509, nx15511, nx15513, nx15515, nx15517, nx15519, nx15521, 
      nx15523, nx15525, nx15527, nx15529, nx15531, nx15533, nx15535, nx15537, 
      nx15539, nx15541, nx15543, nx15545, nx15547, nx15549, nx15551, nx15553, 
      nx15555, nx15557, nx15559, nx15561, nx15563, nx15565, nx15567, nx15569, 
      nx15571, nx15573, nx15575, nx15577, nx15579, nx15581, nx15583, nx15585, 
      nx15587, nx15589, nx15591, nx15593, nx15595, nx15597, nx15599, nx15601, 
      nx15603, nx15605, nx15607, nx15609, nx15611, nx15613, nx15615, nx15617, 
      nx15619, nx15621, nx15623, nx15625, nx15627, nx15629, nx15631, nx15633, 
      nx15635, nx15637, nx15639, nx15641, nx15643, nx15645, nx15647, nx15649, 
      nx15651, nx15653, nx15655, nx15657, nx15659, nx15661, nx15663, nx15665, 
      nx15667, nx15669, nx15671, nx15673, nx15675, nx15677, nx15679, nx15681, 
      nx15683, nx15685, nx15687, nx15689, nx15691, nx15693, nx15695, nx15697, 
      nx15699, nx15701, nx15703, nx15705, nx15707, nx15709, nx15711, nx15713, 
      nx15715, nx15717, nx15719, nx15721, nx15723, nx15725, nx15727, nx15729, 
      nx15731, nx15733, nx15735, nx15737, nx15739, nx15741, nx15743, nx15745, 
      nx15747, nx15749, nx15751, nx15753, nx15755, nx15757, nx15759, nx15761, 
      nx15763, nx15765, nx15767, nx15769, nx15771, nx15773, nx15775, nx15777, 
      nx15779, nx15781, nx15783, nx15785, nx15787, nx15789, nx15791, nx15793, 
      nx15797, nx15799, nx15801, nx15803, nx15805, nx15807, nx15809, nx15813, 
      nx15815, nx15817, nx15819, nx15821, nx15823, nx15825, nx15827, nx15829, 
      nx15831, nx15849, nx15851, nx15853, nx15855, nx15857, nx15859, nx15861, 
      nx15863, nx15865, nx15867, nx15869, nx15871, nx15889, nx15891, nx15893, 
      nx15895, nx15897, nx15899, nx15901, nx15903, nx15905, nx15907, nx15909, 
      nx15911, nx15913, nx15915, nx15917, nx15919, nx15929, nx15931, nx15933, 
      nx15959, nx15961, nx15963, nx15981, nx15983, nx15985, nx15987, nx15989, 
      nx15991, nx16001, nx16003, nx16005, nx16007, nx16009, nx16019, nx16021, 
      nx16023, nx16025, nx16027, nx16029, nx16039, nx16041, nx16043, nx16045, 
      nx16047, nx16049, nx16051, nx16061, nx16063, nx16065, nx16067, nx16069, 
      nx16071, nx16073, nx16091, nx16093, nx16095, nx16097, nx16123, nx16125, 
      nx16127, nx16129, nx16131, nx16133, nx16135, nx16137, nx16139, nx16141, 
      nx16155, nx16157, nx16159, nx16161, nx16163, nx16165, nx16167, nx16169, 
      nx16171, nx16173, nx16175, nx16177, nx16179, nx16181, nx16183, nx16185, 
      nx16187, nx16191, nx16195, nx16197, nx16199, nx16213, nx16215, nx16225, 
      nx16227, nx16229, nx16231, nx16233, nx16235, nx16237, nx16247, nx16257, 
      nx16259, nx16261, nx16263, nx16273, nx16275, nx16277, nx16279, nx16281, 
      nx16325, nx16327, nx16329, nx16331, nx16341, nx16343, nx16345, nx16347, 
      nx16357, nx16359, nx16361, nx16363, nx16373, nx16375, nx16377, nx16379, 
      nx16397, nx16399, nx16401, nx16403, nx16413, nx16415, nx16417, nx16419, 
      nx16437, nx16443, nx16453, nx16459, nx16477, nx16483, nx16493, nx16499, 
      nx16509, nx16511, nx16513, nx16515, nx16517, nx16519, nx16521, nx16523, 
      nx16525, nx16527, nx16529, nx16531, nx16541, nx16543, nx16545, nx16547, 
      nx16557, nx16567, nx16569, nx16571, nx16573, nx16575, nx16577, nx16601, 
      nx16607, nx16609, nx16617, nx16619, nx16621, nx16623, nx16641, nx16643, 
      nx16645, nx16647, nx16657, nx16659, nx16661, nx16663, nx16673, nx16675, 
      nx16677, nx16679, nx16689, nx16691, nx16693, nx16695, nx16705, nx16707, 
      nx16709, nx16711, nx16721, nx16723, nx16725, nx16727, nx16745, nx16747, 
      nx16749, nx16751, nx16753, nx16755, nx16757, nx16759, nx16769, nx16771, 
      nx16773, nx16775, nx16785, nx16787, nx16789, nx16791, nx16817, nx16819, 
      nx16821, nx16823, nx16833, nx16835, nx16837, nx16839, nx16841, nx16843, 
      nx16845, nx16847, nx16849, nx16851, nx16853, nx16855, nx16857, nx16859, 
      nx16861, nx16863, nx16865, nx16867, nx16869, nx16871, nx16873, nx16875, 
      nx16877, nx16879, nx16881, nx16883, nx16885, nx16887, nx16889, nx16891, 
      nx16893, nx16895, nx16897, nx16899, nx16901, nx16903, nx16905, nx16907, 
      nx16909, nx16911, nx16913, nx16915, nx16917, nx16919, nx16921, nx16923, 
      nx16925, nx16927, nx16929, nx16931, nx16933, nx16935, nx16937, nx16939, 
      nx16941, nx16943, nx16945, nx16947, nx16949, nx16951, nx16953, nx16955, 
      nx16957, nx16959, nx16961, nx16963, nx16965, nx16967, nx16969, nx16971, 
      nx16973, nx16975, nx16977, nx16979, nx16981, nx16983, nx16985, nx16987, 
      nx16989, nx16991, nx16993, nx16995, nx16997, nx16999, nx17001, nx17003, 
      nx17005, nx17007, nx17009, nx17011, nx17013, nx17015, nx17017, nx17019, 
      nx17021, nx17023, nx17025, nx17027, nx17029, nx17031, nx17033, nx17035, 
      nx17037, nx17039, nx17041, nx17043, nx17045, nx17047, nx17049, nx17051, 
      nx17053, nx17055, nx17057, nx17059, nx17061, nx17063, nx17065, nx17067, 
      nx17069, nx17071, nx17073, nx17075, nx17077, nx17079, nx17081, nx17083, 
      nx17085, nx17087, nx17089, nx17091, nx17093, nx17095, nx17097, nx17099, 
      nx17101, nx17103, nx17105, nx17107, nx17109, nx17111, nx17113, nx17115, 
      nx17117, nx17119, nx17121, nx17123, nx17125, nx17127, nx17129, nx17131, 
      nx17133, nx17135, nx17137, nx17139, nx17141, nx17143, nx17147, nx17153, 
      nx17155, nx17157, nx17159, nx17165, nx17167, nx17169, nx17171, nx17173, 
      nx17175, nx17179, nx17181, nx17183, nx17185, nx17187, nx17189, nx17191, 
      nx17193, nx17195, nx17197, nx17199, nx17201, nx17203, nx17205, nx17207, 
      nx17209, nx17211, nx17213, nx17215, nx17217, nx17219, nx17221, nx17223, 
      nx17225, nx17227, nx17229, nx17231, nx17233, nx17235, nx17237, nx17239, 
      nx17241, nx17243, nx17245, nx17247, nx17249, nx17251, nx17253, nx17255, 
      nx17257, nx17259, nx17261, nx17263, nx17265, nx17267, nx17269, nx17271, 
      nx17273, nx17275, nx17277, nx17279, nx17281, nx17283, nx17285, nx17287, 
      nx17289, nx17291, nx17293, nx17295, nx17297, nx17299, nx17303, nx17305, 
      nx17307, nx17309, nx17311, nx17313, nx17315, nx17317, nx17319, nx17321, 
      nx17323, nx17325, nx17327, nx17329, nx17331, nx17333, nx17335, nx17337, 
      nx17339, nx17341, nx17343, nx17345, nx17347, nx17349, nx17351, nx17353, 
      nx17355, nx17357, nx17359, nx17361, nx17363, nx17365, nx17367, nx17369, 
      nx17371, nx17373, nx17375, nx17377, nx17379, nx17381, nx17383, nx17385, 
      nx17387, nx17389, nx17391, nx17393, nx17395, nx17397, nx17399, nx17401, 
      nx17403, nx17405, nx17407, nx17409, nx17411, nx17413, nx17415, nx17417, 
      nx17419, nx17421, nx17423, nx17425, nx17427, nx17429, nx17431, nx17433, 
      nx17435, nx17437, nx17439, nx17441, nx17443, nx17445, nx17447, nx17449, 
      nx17451, nx17453, nx17455, nx17457, nx17459, nx17461, nx17463, nx17465, 
      nx17467, nx17469, nx17471, nx17473, nx17475, nx17477, nx17479, nx17481, 
      nx17483, nx17485, nx17487, nx17489, nx17491, nx17493, nx17495, nx17497, 
      nx17499, nx17501, nx17503, nx17505, nx17507, nx17509, nx17511, nx17513, 
      nx17515, nx17517, nx17519, nx17521, nx17523, nx17525, nx17527, nx17529, 
      nx17531, nx17533, nx17535, nx17537, nx17539, nx17541, nx17543, nx17545, 
      nx17547, nx17549, nx17551, nx17553, nx17555, nx17557, nx17559, nx17561, 
      nx17563, nx17565, nx17567, nx17569, nx17571, nx17573, nx17575, nx17577, 
      nx18578, nx18579, nx7274, nx18580, nx18581, nx18582, nx18583, nx18584, 
      nx18585, nx18586, nx18587, NOT_nx7538, nx18588, nx18589, nx18590, 
      nx18591, NOT_nx7576, nx18592, nx18593, nx18594, nx18595, nx18596, 
      nx18597, nx18598, nx18599, nx18600, nx18601, nx13681, nx18602, nx18603, 
      nx3446, nx18604, nx18605, nx18606, nx18607, nx18608, nx18609, nx18610, 
      nx18611, NOT_nx3710, nx18612, nx18613, nx18614, nx18615, NOT_nx3748, 
      nx18616, nx18617, nx18618, nx18619, nx18620, nx18621, nx18622, nx18623, 
      nx18624, nx18625, nx11965, nx18626, nx18627, nx8550, nx18628, nx18629, 
      nx18630, nx18631, nx18632, nx18633, nx18634, nx18635, NOT_nx8814, 
      nx18636, nx18637, nx18638, nx18639, NOT_nx8852, nx18640, nx18641, 
      nx18642, nx18643, nx18644, nx18645, nx18646, nx18647, nx18648, nx18649, 
      nx14253, nx18650, nx18651, nx2808, nx18652, nx18653, nx18654, nx18655, 
      nx18656, nx18657, nx18658, nx18659, NOT_nx3072, nx18660, nx18661, 
      nx18662, nx18663, NOT_nx3110, nx18664, nx18665, nx18666, nx18667, 
      nx18668, nx18669, nx18670, nx18671, nx18672, nx18673, nx11679, nx18674, 
      nx18675, nx6636, nx18676, nx18677, nx18678, nx18679, nx18680, nx18681, 
      nx18682, nx18683, NOT_nx6900, nx18684, nx18685, nx18686, nx18687, 
      NOT_nx6938, nx18688, nx18689, nx18690, nx18691, nx18692, nx18693, 
      nx18694, nx18695, nx18696, nx18697, nx13395, nx18698, nx18699, nx7912, 
      nx18700, nx18701, nx18702, nx18703, nx18704, nx18705, nx18706, nx18707, 
      NOT_nx8176, nx18708, nx18709, nx18710, nx18711, NOT_nx8214, nx18712, 
      nx18713, nx18714, nx18715, nx18716, nx18717, nx18718, nx18719, nx18720, 
      nx18721, nx13967, nx18722, nx18723, nx4084, nx18724, nx18725, nx18726, 
      nx18727, nx18728, nx18729, nx18730, nx18731, NOT_nx4348, nx18732, 
      nx18733, nx18734, nx18735, NOT_nx4386, nx18736, nx18737, nx18738, 
      nx18739, nx18740, nx18741, nx18742, nx18743, nx18744, nx18745, nx12251, 
      nx18746, nx18747, nx2170, nx18748, nx18749, nx18750, nx18751, nx18752, 
      nx18753, nx18754, nx18755, NOT_nx2434, nx18756, nx18757, nx18758, 
      NOT_nx2364, nx18759, nx18760, nx18761, NOT_nx2472, NOT_nx2442, nx18762, 
      nx18763, nx18764, nx18765, nx11393, nx18766, nx18767, nx5360, nx18768, 
      nx18769, nx18770, nx18771, nx18772, nx18773, nx18774, nx18775, 
      NOT_nx5624, nx18776, nx18777, nx18778, nx18779, NOT_nx5662, nx18780, 
      nx18781, nx18782, nx18783, nx18784, nx18785, nx18786, nx18787, nx18788, 
      nx18789, nx12823, nx18790, nx18791, nx5998, nx18792, nx18793, nx18794, 
      nx18795, nx18796, nx18797, nx18798, nx18799, NOT_nx6262, nx18800, 
      nx18801, nx18802, nx18803, NOT_nx6300, nx18804, nx18805, nx18806, 
      nx18807, nx18808, nx18809, nx18810, nx18811, nx18812, nx18813, nx13109, 
      nx18814, nx18815, nx4722, nx18816, nx18817, nx18818, nx18819, 
      NOT_nx4986, nx18820, nx18821, nx18822, nx18823, NOT_nx5024, nx18824, 
      nx18825, nx18826, nx18827, NOT_nx4954, nx18828, nx18829, nx18830, 
      nx12537, nx18831, nx18832, nx384, nx18833, nx18834, nx18835, nx18836, 
      nx18837, nx18838, nx18839, nx18840, NOT_nx940, nx18841, nx18842, 
      nx18843, NOT_nx798, nx18844, nx18845, nx18846, NOT_nx1022, NOT_nx960, 
      nx18847, nx18848, nx18849, nx18850, nx10491, nx18851, nx18852, nx1532, 
      nx18853, nx18854, nx18855, nx18856, nx18857, nx18858, nx18859, nx18860, 
      NOT_nx1796, nx18861, nx18862, nx18863, NOT_nx1726, nx18864, nx18865, 
      nx18866, NOT_nx1834, NOT_nx1804, nx18867, nx18868, nx18869, nx18870, 
      nx11107, nx18871, nx18872, nx9188, nx18873, nx18874, NOT_nx9452, 
      nx18875, nx18876, nx18877, NOT_nx9420, nx18878, nx18879, nx18880, 
      nx18881, nx18882, nx18883, nx18884, nx18885, nx18886, nx14539, nx18887, 
      nx18888, nx10464, nx18889, nx18890, nx18891, NOT_nx10688, nx18892, 
      nx18893, nx18894, nx18895, nx18896, nx18897, nx18898, nx18899, nx18900, 
      nx18901, nx18902, nx18903, nx18904, nx15111, nx18905, nx18906, nx9826, 
      nx18907, nx18908, nx18909, nx18910, NOT_nx10090, nx18911, nx18912, 
      nx18913, nx18914, nx18915, nx18916, nx18917, nx18918, nx18919, nx18920, 
      nx18921, nx18922, nx18923, nx14825, nx10545, nx18924, nx17301, nx10523, 
      nx10511, nx16283, nx10949, nx10525, nx17177, nx16151, nx18925, nx18926, 
      nx18927, nx18928, nx18929, nx2622, nx18930, nx2226, nx18931, nx18932, 
      nx18933, nx18934, nx18935, nx18936, nx18937, nx1984, nx18938, nx1588, 
      nx18939, nx18940, nx18941, nx18942, nx18943, nx18944, nx18945, nx1326, 
      nx16495, nx16479, nx18946, nx16603, nx514, nx16455, nx16439, nx18947, 
      nx18948, nx16201, nx10565, nx18949, nx18950, nx9640, nx16497, nx16481, 
      nx18951, nx16605, nx9244, nx16457, nx16441, nx18952, nx18953, nx16203, 
      nx18954, nx12737, nx18955, nx18956, nx18957, nx18958, nx19341, nx19343
   : std_logic ;

begin
   tri_data_out_0 : tri01 port map ( Y=>data_out(0), A=>nx10491, E=>
      write_out);
   ix1365 : oai22 port map ( Y=>nx1364, A0=>nx10497, A1=>nx16157, B0=>
      nx10529, B1=>nx16183);
   modgen_ram_ix74_ix4012 : dff port map ( Q=>OPEN, QB=>nx10497, D=>nx879, 
      CLK=>nx15457);
   ix10504 : nand02 port map ( Y=>nx10503, A0=>nx10505, A1=>nx15453);
   ix10506 : nor03_2x port map ( Y=>nx10505, A0=>nx10507, A1=>address(3), A2
      =>nx17177);
   ix10508 : inv02 port map ( Y=>nx10507, A=>address(2));
   ix123 : inv02 port map ( Y=>nx122, A=>nx18955);
   ix19 : nor02_2x port map ( Y=>nx18, A0=>nx10514, A1=>nx17141);
   ix10515 : inv02 port map ( Y=>nx10514, A=>read_in);
   ix15 : nand02 port map ( Y=>nx14, A0=>address(4), A1=>address(5));
   ix10520 : nand03 port map ( Y=>nx10519, A0=>nx10521, A1=>nx16163, A2=>
      nx18955);
   ix10522 : nor02_2x port map ( Y=>nx10521, A0=>nx10523, A1=>nx10525);
   ix10528 : nor02_2x port map ( Y=>nx10527, A0=>nx10507, A1=>address(3));
   modgen_ram_ix74_ix4120 : dff port map ( Q=>OPEN, QB=>nx10529, D=>nx869, 
      CLK=>nx15457);
   ix1331 : nor02_2x port map ( Y=>nx1330, A0=>nx15889, A1=>nx16177);
   ix405 : nand03 port map ( Y=>nx404, A0=>nx16167, A1=>address(0), A2=>
      nx16171);
   ix10535 : nor02_2x port map ( Y=>nx10534, A0=>address(2), A1=>nx10537);
   ix10538 : inv02 port map ( Y=>nx10537, A=>address(3));
   ix10542 : nand03 port map ( Y=>nx10541, A0=>read_in, A1=>address(4), A2=>
      nx10525);
   ix10544 : nand04 port map ( Y=>nx10543, A0=>nx17147, A1=>nx16167, A2=>
      address(0), A3=>nx16171);
   modgen_ram_ix74_ix4096 : dff port map ( Q=>OPEN, QB=>nx10548, D=>nx849, 
      CLK=>nx15457);
   ix1293 : nor03_2x port map ( Y=>nx1292, A0=>nx96, A1=>nx450, A2=>nx16177
   );
   ix97 : nand02_2x port map ( Y=>nx96, A0=>address(0), A1=>address(1));
   ix451 : nand02_2x port map ( Y=>nx450, A0=>address(2), A1=>address(3));
   ix10556 : nand02 port map ( Y=>nx10555, A0=>nx17147, A1=>nx10557);
   ix10558 : nor02_2x port map ( Y=>nx10557, A0=>nx96, A1=>nx450);
   modgen_ram_ix74_ix4104 : dff port map ( Q=>OPEN, QB=>nx10559, D=>nx859, 
      CLK=>nx15457);
   ix1311 : nor02_2x port map ( Y=>nx1310, A0=>nx15911, A1=>nx16177);
   ix453 : nand04 port map ( Y=>nx452, A0=>address(0), A1=>nx16171, A2=>
      address(2), A3=>address(3));
   ix10568 : nor02_2x port map ( Y=>nx10567, A0=>nx16213, A1=>address(1));
   ix10572 : nor02_2x port map ( Y=>nx10571, A0=>nx1286, A1=>nx1248);
   ix1287 : oai33 port map ( Y=>nx1286, A0=>nx10574, A1=>nx15849, A2=>
      nx16093, B0=>nx10584, B1=>nx17141, B2=>nx16021);
   modgen_ram_ix74_ix4204 : dff port map ( Q=>OPEN, QB=>nx10574, D=>nx829, 
      CLK=>nx15457);
   ix10578 : nand04 port map ( Y=>nx10577, A0=>nx16163, A1=>nx18955, A2=>
      read_in, A3=>nx16225);
   ix10580 : nor02_2x port map ( Y=>nx10579, A0=>address(4), A1=>address(5)
   );
   ix219 : inv04 port map ( Y=>nx218, A=>nx10579);
   modgen_ram_ix74_ix4016 : dff port map ( Q=>OPEN, QB=>nx10584, D=>nx839, 
      CLK=>nx15457);
   ix10588 : nand02 port map ( Y=>nx10587, A0=>nx10589, A1=>nx15453);
   ix10590 : nor03_2x port map ( Y=>nx10589, A0=>address(2), A1=>address(3), 
      A2=>nx96);
   ix943 : nand03 port map ( Y=>nx942, A0=>nx16247, A1=>address(0), A2=>
      address(1));
   ix10593 : nor02_2x port map ( Y=>nx10592, A0=>address(2), A1=>address(3)
   );
   ix1249 : oai22 port map ( Y=>nx1248, A0=>nx10595, A1=>nx16259, B0=>
      nx10603, B1=>nx16275);
   modgen_ram_ix74_ix4140 : dff port map ( Q=>OPEN, QB=>nx10595, D=>nx819, 
      CLK=>nx15457);
   ix10600 : nand03 port map ( Y=>nx10599, A0=>nx10505, A1=>read_in, A2=>
      nx17147);
   modgen_ram_ix74_ix4076 : dff port map ( Q=>OPEN, QB=>nx10603, D=>nx809, 
      CLK=>nx15459);
   ix10608 : nand02 port map ( Y=>nx10607, A0=>nx10505, A1=>nx15793);
   ix53 : nor02_2x port map ( Y=>nx52, A0=>nx10514, A1=>nx15759);
   ix49 : nand02 port map ( Y=>nx48, A0=>nx10523, A1=>address(5));
   ix10612 : nand03 port map ( Y=>nx10611, A0=>nx16281, A1=>nx16163, A2=>
      nx18955);
   ix10614 : nor02_2x port map ( Y=>nx10613, A0=>address(4), A1=>nx10525);
   ix10616 : nor03_2x port map ( Y=>nx10615, A0=>nx1202, A1=>nx1184, A2=>
      nx1166);
   ix1203 : nor03_2x port map ( Y=>nx1202, A0=>nx10619, A1=>nx15759, A2=>
      nx16061);
   modgen_ram_ix74_ix4032 : dff port map ( Q=>OPEN, QB=>nx10619, D=>nx799, 
      CLK=>nx15459);
   ix1189 : nor03_2x port map ( Y=>nx1188, A0=>nx96, A1=>nx450, A2=>nx10625
   );
   ix10626 : nand03 port map ( Y=>nx10625, A0=>read_in, A1=>nx10523, A2=>
      address(5));
   ix1089 : nand04 port map ( Y=>nx1088, A0=>address(0), A1=>address(1), A2
      =>address(2), A3=>address(3));
   ix1185 : nor03_2x port map ( Y=>nx1184, A0=>nx10629, A1=>nx15849, A2=>
      nx15403);
   modgen_ram_ix74_ix4200 : dff port map ( Q=>OPEN, QB=>nx10629, D=>nx789, 
      CLK=>nx15459);
   ix10634 : nand04 port map ( Y=>nx10633, A0=>nx16163, A1=>nx10567, A2=>
      read_in, A3=>nx16225);
   ix9 : nand03 port map ( Y=>nx8, A0=>nx16163, A1=>address(0), A2=>nx16171
   );
   ix1167 : oai33 port map ( Y=>nx1166, A0=>nx10637, A1=>nx15759, A2=>
      nx15911, B0=>nx10645, B1=>nx17141, B2=>nx16061);
   modgen_ram_ix74_ix4040 : dff port map ( Q=>OPEN, QB=>nx10637, D=>nx769, 
      CLK=>nx15459);
   ix10642 : nand02 port map ( Y=>nx10641, A0=>nx10643, A1=>nx15793);
   ix10644 : nor03_2x port map ( Y=>nx10643, A0=>nx16213, A1=>address(1), A2
      =>nx450);
   modgen_ram_ix74_ix3968 : dff port map ( Q=>OPEN, QB=>nx10645, D=>nx779, 
      CLK=>nx15459);
   ix10649 : nand02 port map ( Y=>nx10648, A0=>nx10557, A1=>nx15453);
   ix10652 : nor03_2x port map ( Y=>nx10651, A0=>nx1124, A1=>nx1106, A2=>
      nx1086);
   ix1125 : nor03_2x port map ( Y=>nx1124, A0=>nx10654, A1=>nx15759, A2=>
      nx16039);
   modgen_ram_ix74_ix4036 : dff port map ( Q=>OPEN, QB=>nx10654, D=>nx759, 
      CLK=>nx15459);
   ix10658 : nand03 port map ( Y=>nx10657, A0=>nx10659, A1=>read_in, A2=>
      nx16281);
   ix10660 : nor03_2x port map ( Y=>nx10659, A0=>address(0), A1=>nx16171, A2
      =>nx450);
   ix1005 : nand03 port map ( Y=>nx1004, A0=>nx10663, A1=>address(2), A2=>
      address(3));
   ix10664 : nor02_2x port map ( Y=>nx10663, A0=>address(0), A1=>nx16171);
   ix1107 : nor04 port map ( Y=>nx1106, A0=>nx10666, A1=>address(4), A2=>
      address(5), A3=>nx16061);
   modgen_ram_ix74_ix4160 : dff port map ( Q=>OPEN, QB=>nx10666, D=>nx749, 
      CLK=>nx15459);
   ix1093 : nor03_2x port map ( Y=>nx1092, A0=>nx96, A1=>nx450, A2=>nx10671
   );
   ix10672 : nand02 port map ( Y=>nx10671, A0=>read_in, A1=>nx16225);
   ix1087 : oai22 port map ( Y=>nx1086, A0=>nx10674, A1=>nx16327, B0=>
      nx10681, B1=>nx16343);
   modgen_ram_ix74_ix3976 : dff port map ( Q=>OPEN, QB=>nx10674, D=>nx729, 
      CLK=>nx15461);
   ix10678 : nand02 port map ( Y=>nx10677, A0=>nx10643, A1=>nx15453);
   ix10680 : nand04 port map ( Y=>nx10679, A0=>nx10521, A1=>nx10567, A2=>
      address(2), A3=>address(3));
   modgen_ram_ix74_ix3972 : dff port map ( Q=>OPEN, QB=>nx10681, D=>nx739, 
      CLK=>nx15461);
   ix10685 : nand02 port map ( Y=>nx10684, A0=>nx10659, A1=>nx15453);
   ix10687 : nand04 port map ( Y=>nx10686, A0=>nx10521, A1=>nx10663, A2=>
      address(2), A3=>address(3));
   modgen_ram_ix74_ix4100 : dff port map ( Q=>OPEN, QB=>nx10692, D=>nx719, 
      CLK=>nx15461);
   ix1027 : nor02_2x port map ( Y=>nx1026, A0=>nx16039, A1=>nx16177);
   ix151 : nand02 port map ( Y=>nx150, A0=>address(4), A1=>nx10525);
   modgen_ram_ix74_ix4164 : dff port map ( Q=>OPEN, QB=>nx10699, D=>nx709, 
      CLK=>nx15461);
   ix10704 : nand03 port map ( Y=>nx10703, A0=>nx10659, A1=>read_in, A2=>
      nx16225);
   ix1003 : oai22 port map ( Y=>nx1002, A0=>nx10706, A1=>nx16359, B0=>
      nx10713, B1=>nx16375);
   modgen_ram_ix74_ix4144 : dff port map ( Q=>OPEN, QB=>nx10706, D=>nx689, 
      CLK=>nx15461);
   ix969 : nor02_2x port map ( Y=>nx968, A0=>nx16021, A1=>nx16177);
   ix10712 : nand04 port map ( Y=>nx10711, A0=>nx17147, A1=>nx16247, A2=>
      address(0), A3=>address(1));
   modgen_ram_ix74_ix4080 : dff port map ( Q=>OPEN, QB=>nx10713, D=>nx699, 
      CLK=>nx15461);
   ix10717 : nand03 port map ( Y=>nx10716, A0=>nx10589, A1=>read_in, A2=>
      nx16281);
   ix10720 : nand04 port map ( Y=>nx10719, A0=>nx16281, A1=>nx16247, A2=>
      address(0), A3=>address(1));
   modgen_ram_ix74_ix4208 : dff port map ( Q=>OPEN, QB=>nx10724, D=>nx679, 
      CLK=>nx15461);
   ix10728 : nand03 port map ( Y=>nx10727, A0=>nx10589, A1=>read_in, A2=>
      nx16225);
   modgen_ram_ix74_ix4020 : dff port map ( Q=>OPEN, QB=>nx10731, D=>nx669, 
      CLK=>nx15463);
   ix10735 : nand02 port map ( Y=>nx10734, A0=>nx10737, A1=>nx15453);
   ix10738 : nor03_2x port map ( Y=>nx10737, A0=>address(2), A1=>address(3), 
      A2=>nx42);
   ix43 : nand02 port map ( Y=>nx42, A0=>nx16213, A1=>address(1));
   ix861 : nand03 port map ( Y=>nx860, A0=>nx16247, A1=>nx16213, A2=>
      address(1));
   ix923 : oai22 port map ( Y=>nx922, A0=>nx10744, A1=>nx16399, B0=>nx10751, 
      B1=>nx16415);
   modgen_ram_ix74_ix4148 : dff port map ( Q=>OPEN, QB=>nx10744, D=>nx649, 
      CLK=>nx15463);
   ix889 : nor02_2x port map ( Y=>nx888, A0=>nx16001, A1=>nx16177);
   ix10750 : nand04 port map ( Y=>nx10749, A0=>nx17147, A1=>nx16247, A2=>
      nx16213, A3=>address(1));
   modgen_ram_ix74_ix4084 : dff port map ( Q=>OPEN, QB=>nx10751, D=>nx659, 
      CLK=>nx15463);
   ix10755 : nand03 port map ( Y=>nx10754, A0=>nx10737, A1=>read_in, A2=>
      nx16281);
   ix10758 : nand04 port map ( Y=>nx10757, A0=>nx16281, A1=>nx16247, A2=>
      nx16213, A3=>address(1));
   modgen_ram_ix74_ix4212 : dff port map ( Q=>OPEN, QB=>nx10762, D=>nx639, 
      CLK=>nx15463);
   ix10766 : nand03 port map ( Y=>nx10765, A0=>nx10737, A1=>read_in, A2=>
      nx16225);
   modgen_ram_ix74_ix4024 : dff port map ( Q=>OPEN, QB=>nx10769, D=>nx629, 
      CLK=>nx15463);
   ix10773 : nand02 port map ( Y=>nx10772, A0=>nx10775, A1=>nx15453);
   ix10776 : nor03_2x port map ( Y=>nx10775, A0=>address(2), A1=>address(3), 
      A2=>nx2);
   ix3 : nand02 port map ( Y=>nx2, A0=>address(0), A1=>nx16171);
   ix781 : nand03 port map ( Y=>nx780, A0=>nx16247, A1=>address(0), A2=>
      nx16173);
   modgen_ram_ix74_ix4152 : dff port map ( Q=>OPEN, QB=>nx10783, D=>nx609, 
      CLK=>nx15463);
   ix807 : nor02_2x port map ( Y=>nx806, A0=>nx15983, A1=>nx16177);
   ix10788 : nand04 port map ( Y=>nx10787, A0=>nx19341, A1=>nx10592, A2=>
      address(0), A3=>nx16173);
   modgen_ram_ix74_ix4088 : dff port map ( Q=>OPEN, QB=>nx10789, D=>nx619, 
      CLK=>nx15463);
   ix10794 : nand02 port map ( Y=>nx10793, A0=>nx10775, A1=>nx15793);
   ix10796 : nand04 port map ( Y=>nx10795, A0=>nx16281, A1=>nx10592, A2=>
      address(0), A3=>nx16173);
   modgen_ram_ix74_ix4216 : dff port map ( Q=>OPEN, QB=>nx10801, D=>nx599, 
      CLK=>nx15465);
   ix10805 : nand04 port map ( Y=>nx10804, A0=>nx10592, A1=>nx10567, A2=>
      read_in, A3=>nx16225);
   ix779 : nor03_2x port map ( Y=>nx778, A0=>nx10807, A1=>nx17141, A2=>
      nx15959);
   modgen_ram_ix74_ix4028 : dff port map ( Q=>OPEN, QB=>nx10807, D=>nx589, 
      CLK=>nx15465);
   ix10812 : nand02 port map ( Y=>nx10811, A0=>nx10813, A1=>nx15455);
   ix10814 : nor03_2x port map ( Y=>nx10813, A0=>address(2), A1=>address(3), 
      A2=>nx16151);
   ix695 : nand02 port map ( Y=>nx694, A0=>nx10592, A1=>nx18955);
   modgen_ram_ix74_ix4156 : dff port map ( Q=>OPEN, QB=>nx10817, D=>nx569, 
      CLK=>nx15465);
   ix727 : nor02_2x port map ( Y=>nx726, A0=>nx15959, A1=>nx16179);
   ix10824 : nand04 port map ( Y=>nx10823, A0=>nx19341, A1=>nx10592, A2=>
      nx16213, A3=>nx16173);
   modgen_ram_ix74_ix4092 : dff port map ( Q=>OPEN, QB=>nx10825, D=>nx579, 
      CLK=>nx15465);
   ix10830 : nand02 port map ( Y=>nx10829, A0=>nx10813, A1=>nx15793);
   ix10832 : nand04 port map ( Y=>nx10831, A0=>nx19343, A1=>nx10592, A2=>
      nx16215, A3=>nx16173);
   ix715 : oai22 port map ( Y=>nx714, A0=>nx10841, A1=>nx16511, B0=>nx10852, 
      B1=>nx16519);
   modgen_ram_ix74_ix4184 : dff port map ( Q=>OPEN, QB=>nx10841, D=>nx549, 
      CLK=>nx15465);
   ix10845 : nand03 port map ( Y=>nx10844, A0=>nx10847, A1=>read_in, A2=>
      nx16227);
   ix10848 : nor02_2x port map ( Y=>nx10847, A0=>nx126, A1=>nx2);
   ix127 : nand02 port map ( Y=>nx126, A0=>nx10507, A1=>address(3));
   ix10851 : nand04 port map ( Y=>nx10850, A0=>nx16227, A1=>nx16167, A2=>
      address(0), A3=>nx16173);
   modgen_ram_ix74_ix4220 : dff port map ( Q=>OPEN, QB=>nx10852, D=>nx559, 
      CLK=>nx15465);
   ix699 : nor02_2x port map ( Y=>nx698, A0=>nx15959, A1=>nx10671);
   ix10858 : nand04 port map ( Y=>nx10857, A0=>nx16227, A1=>nx10592, A2=>
      nx16215, A3=>nx16173);
   ix673 : oai22 port map ( Y=>nx672, A0=>nx10861, A1=>nx16527, B0=>nx10869, 
      B1=>nx16543);
   modgen_ram_ix74_ix4116 : dff port map ( Q=>OPEN, QB=>nx10861, D=>nx539, 
      CLK=>nx15465);
   ix657 : nor02_2x port map ( Y=>nx656, A0=>nx358, A1=>nx16179);
   ix359 : nand03 port map ( Y=>nx358, A0=>nx16167, A1=>nx16215, A2=>
      address(1));
   ix10867 : nand04 port map ( Y=>nx10866, A0=>nx19341, A1=>nx16167, A2=>
      nx16215, A3=>address(1));
   modgen_ram_ix74_ix4052 : dff port map ( Q=>OPEN, QB=>nx10869, D=>nx529, 
      CLK=>nx15467);
   ix10873 : nand03 port map ( Y=>nx10872, A0=>nx10874, A1=>read_in, A2=>
      nx19343);
   ix10875 : nor03_2x port map ( Y=>nx10874, A0=>address(2), A1=>nx10537, A2
      =>nx42);
   ix10878 : nand04 port map ( Y=>nx10877, A0=>nx19343, A1=>nx16167, A2=>
      nx16215, A3=>address(1));
   ix635 : nand03 port map ( Y=>nx634, A0=>nx10881, A1=>nx10899, A2=>nx10909
   );
   ix10882 : nor02_2x port map ( Y=>nx10881, A0=>nx630, A1=>nx612);
   ix631 : nor04 port map ( Y=>nx630, A0=>nx10884, A1=>address(4), A2=>
      address(5), A3=>nx15895);
   modgen_ram_ix74_ix4176 : dff port map ( Q=>OPEN, QB=>nx10884, D=>nx519, 
      CLK=>nx15467);
   ix10888 : nand03 port map ( Y=>nx10887, A0=>nx10889, A1=>read_in, A2=>
      nx16227);
   ix10890 : nor03_2x port map ( Y=>nx10889, A0=>address(2), A1=>nx10537, A2
      =>nx96);
   ix427 : nand03 port map ( Y=>nx426, A0=>nx16167, A1=>address(0), A2=>
      address(1));
   ix613 : nor03_2x port map ( Y=>nx612, A0=>nx10893, A1=>nx15819, A2=>
      nx15895);
   modgen_ram_ix74_ix4112 : dff port map ( Q=>OPEN, QB=>nx10893, D=>nx509, 
      CLK=>nx15467);
   ix599 : nor02_2x port map ( Y=>nx598, A0=>nx15895, A1=>nx16179);
   ix10900 : nand03 port map ( Y=>nx10899, A0=>modgen_ram_ix74_a_12_dup_1207, 
      A1=>nx16227, A2=>nx16567);
   modgen_ram_ix74_ix4172 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_1207, 
      QB=>nx10903, D=>nx499, CLK=>nx15467);
   ix10908 : nor03_2x port map ( Y=>nx10907, A0=>address(0), A1=>address(1), 
      A2=>nx450);
   ix10910 : nand03 port map ( Y=>nx10909, A0=>modgen_ram_ix74_a_28_dup_1191, 
      A1=>nx19341, A2=>nx16567);
   modgen_ram_ix74_ix4108 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_1191, 
      QB=>nx10913, D=>nx489, CLK=>nx15467);
   ix561 : nor02_2x port map ( Y=>nx560, A0=>nx15929, A1=>nx16179);
   ix477 : nand03 port map ( Y=>nx476, A0=>nx18955, A1=>address(2), A2=>
      address(3));
   modgen_ram_ix74_ix3980 : dff port map ( Q=>OPEN, QB=>nx10922, D=>nx479, 
      CLK=>nx15467);
   modgen_ram_ix74_ix4056 : dff port map ( Q=>OPEN, QB=>nx10928, D=>nx469, 
      CLK=>nx15467);
   ix10932 : nand02 port map ( Y=>nx10931, A0=>nx10847, A1=>nx15793);
   modgen_ram_ix74_ix4048 : dff port map ( Q=>OPEN, QB=>nx10935, D=>nx459, 
      CLK=>nx15469);
   ix10940 : nand03 port map ( Y=>nx10939, A0=>nx10889, A1=>read_in, A2=>
      nx19343);
   ix10942 : nand04 port map ( Y=>nx10941, A0=>nx19343, A1=>nx16169, A2=>
      address(0), A3=>address(1));
   modgen_ram_ix74_ix4044 : dff port map ( Q=>OPEN, QB=>nx10943, D=>nx449, 
      CLK=>nx15469);
   ix10952 : nor03_2x port map ( Y=>nx10951, A0=>nx470, A1=>nx444, A2=>nx424
   );
   ix471 : nor03_2x port map ( Y=>nx470, A0=>nx10954, A1=>nx15849, A2=>
      nx15911);
   modgen_ram_ix74_ix4168 : dff port map ( Q=>OPEN, QB=>nx10954, D=>nx439, 
      CLK=>nx15469);
   ix457 : nor02_2x port map ( Y=>nx456, A0=>nx15911, A1=>nx10671);
   ix445 : nor03_2x port map ( Y=>nx444, A0=>nx10959, A1=>nx15417, A2=>
      nx15895);
   modgen_ram_ix74_ix3984 : dff port map ( Q=>OPEN, QB=>nx10959, D=>nx429, 
      CLK=>nx15469);
   ix10963 : nand02 port map ( Y=>nx10962, A0=>nx10889, A1=>nx15455);
   ix425 : oai22 port map ( Y=>nx424, A0=>nx10965, A1=>nx16643, B0=>nx10972, 
      B1=>nx16659);
   modgen_ram_ix74_ix3992 : dff port map ( Q=>OPEN, QB=>nx10965, D=>nx419, 
      CLK=>nx15469);
   ix10969 : nand02 port map ( Y=>nx10968, A0=>nx10847, A1=>nx15455);
   ix10971 : nand04 port map ( Y=>nx10970, A0=>nx10521, A1=>nx16169, A2=>
      address(0), A3=>nx16175);
   modgen_ram_ix74_ix3988 : dff port map ( Q=>OPEN, QB=>nx10972, D=>nx409, 
      CLK=>nx15469);
   ix10976 : nand02 port map ( Y=>nx10975, A0=>nx10874, A1=>nx15455);
   ix10978 : nand04 port map ( Y=>nx10977, A0=>nx10521, A1=>nx16169, A2=>
      nx16215, A3=>address(1));
   ix379 : oai22 port map ( Y=>nx378, A0=>nx10983, A1=>nx16675, B0=>nx10992, 
      B1=>nx16691);
   modgen_ram_ix74_ix4136 : dff port map ( Q=>OPEN, QB=>nx10983, D=>nx389, 
      CLK=>nx15469);
   ix10987 : nand03 port map ( Y=>nx10986, A0=>nx10988, A1=>read_in, A2=>
      nx19341);
   ix10989 : nor03_2x port map ( Y=>nx10988, A0=>nx10507, A1=>address(3), A2
      =>nx2);
   ix10991 : nand04 port map ( Y=>nx10990, A0=>nx19341, A1=>nx16165, A2=>
      address(0), A3=>nx16175);
   modgen_ram_ix74_ix4180 : dff port map ( Q=>OPEN, QB=>nx10992, D=>nx399, 
      CLK=>nx15471);
   ix10996 : nand03 port map ( Y=>nx10995, A0=>nx10874, A1=>read_in, A2=>
      nx16227);
   ix10998 : nand04 port map ( Y=>nx10997, A0=>nx16229, A1=>nx16169, A2=>
      nx16215, A3=>address(1));
   ix339 : oai22 port map ( Y=>nx338, A0=>nx11000, A1=>nx16707, B0=>nx11007, 
      B1=>nx16723);
   modgen_ram_ix74_ix4196 : dff port map ( Q=>OPEN, QB=>nx11000, D=>nx379, 
      CLK=>nx15471);
   ix11004 : nand04 port map ( Y=>nx11003, A0=>nx16165, A1=>nx10663, A2=>
      read_in, A3=>nx16229);
   modgen_ram_ix74_ix4132 : dff port map ( Q=>OPEN, QB=>nx11007, D=>nx369, 
      CLK=>nx15471);
   ix11011 : nand03 port map ( Y=>nx11010, A0=>nx11012, A1=>read_in, A2=>
      nx19341);
   ix11013 : nor03_2x port map ( Y=>nx11012, A0=>nx10507, A1=>address(3), A2
      =>nx42);
   ix11017 : nor03_2x port map ( Y=>nx11016, A0=>nx296, A1=>nx278, A2=>nx260
   );
   ix297 : nor03_2x port map ( Y=>nx296, A0=>nx11019, A1=>nx15417, A2=>
      nx15753);
   modgen_ram_ix74_ix4004 : dff port map ( Q=>OPEN, QB=>nx11019, D=>nx359, 
      CLK=>nx15471);
   ix11023 : nand02 port map ( Y=>nx11022, A0=>nx11012, A1=>nx15455);
   ix45 : nand02 port map ( Y=>nx44, A0=>nx16165, A1=>nx10663);
   ix279 : nor03_2x port map ( Y=>nx278, A0=>nx11026, A1=>nx15849, A2=>
      nx15797);
   modgen_ram_ix74_ix4192 : dff port map ( Q=>OPEN, QB=>nx11026, D=>nx349, 
      CLK=>nx15471);
   ix265 : nor02_2x port map ( Y=>nx264, A0=>nx15797, A1=>nx10671);
   ix99 : nand04 port map ( Y=>nx98, A0=>address(2), A1=>nx10537, A2=>
      address(0), A3=>address(1));
   ix261 : oai22 port map ( Y=>nx260, A0=>nx11032, A1=>nx16747, B0=>nx11041, 
      B1=>nx16755);
   modgen_ram_ix74_ix4000 : dff port map ( Q=>OPEN, QB=>nx11032, D=>nx339, 
      CLK=>nx15471);
   ix11036 : nand02 port map ( Y=>nx11035, A0=>nx11037, A1=>nx15455);
   ix11038 : nor03_2x port map ( Y=>nx11037, A0=>nx10507, A1=>address(3), A2
      =>nx96);
   ix11040 : nand04 port map ( Y=>nx11039, A0=>nx10521, A1=>nx16165, A2=>
      address(0), A3=>address(1));
   modgen_ram_ix74_ix4188 : dff port map ( Q=>OPEN, QB=>nx11041, D=>nx329, 
      CLK=>nx15471);
   ix227 : nor02_2x port map ( Y=>nx226, A0=>nx15813, A1=>nx10671);
   ix129 : nand02 port map ( Y=>nx128, A0=>nx16169, A1=>nx18955);
   ix11049 : nor03_2x port map ( Y=>nx11048, A0=>nx210, A1=>nx192, A2=>nx174
   );
   ix211 : nor03_2x port map ( Y=>nx210, A0=>nx11051, A1=>nx15759, A2=>
      nx15813);
   modgen_ram_ix74_ix4060 : dff port map ( Q=>OPEN, QB=>nx11051, D=>nx319, 
      CLK=>nx15473);
   ix11055 : nand02 port map ( Y=>nx11054, A0=>nx11056, A1=>nx15793);
   ix11057 : nor03_2x port map ( Y=>nx11056, A0=>address(2), A1=>nx10537, A2
      =>nx18925);
   ix193 : nor03_2x port map ( Y=>nx192, A0=>nx11059, A1=>nx15819, A2=>
      nx15797);
   modgen_ram_ix74_ix4128 : dff port map ( Q=>OPEN, QB=>nx11059, D=>nx309, 
      CLK=>nx15473);
   ix179 : nor02_2x port map ( Y=>nx178, A0=>nx15797, A1=>nx16179);
   ix175 : oai22 port map ( Y=>nx174, A0=>nx11064, A1=>nx16771, B0=>nx11070, 
      B1=>nx16787);
   modgen_ram_ix74_ix4124 : dff port map ( Q=>OPEN, QB=>nx11064, D=>nx299, 
      CLK=>nx15473);
   ix159 : nor02_2x port map ( Y=>nx158, A0=>nx15813, A1=>nx16179);
   modgen_ram_ix74_ix3996 : dff port map ( Q=>OPEN, QB=>nx11070, D=>nx289, 
      CLK=>nx15473);
   ix11074 : nand02 port map ( Y=>nx11073, A0=>nx11056, A1=>nx18);
   ix11076 : nand03 port map ( Y=>nx11075, A0=>nx10521, A1=>nx10534, A2=>
      nx18956);
   ix11078 : nor03_2x port map ( Y=>nx11077, A0=>nx116, A1=>nx90, A2=>nx72);
   ix117 : nor03_2x port map ( Y=>nx116, A0=>nx11080, A1=>nx15759, A2=>
      nx15797);
   modgen_ram_ix74_ix4064 : dff port map ( Q=>OPEN, QB=>nx11080, D=>nx279, 
      CLK=>nx15473);
   ix11084 : nand02 port map ( Y=>nx11083, A0=>nx11037, A1=>nx15793);
   ix91 : nor03_2x port map ( Y=>nx90, A0=>nx11086, A1=>nx15761, A2=>nx15403
   );
   modgen_ram_ix74_ix4072 : dff port map ( Q=>OPEN, QB=>nx11086, D=>nx269, 
      CLK=>nx15473);
   ix11090 : nand02 port map ( Y=>nx11089, A0=>nx10988, A1=>nx52);
   ix73 : oai22 port map ( Y=>nx72, A0=>nx11092, A1=>nx16819, B0=>nx11099, 
      B1=>nx16835);
   modgen_ram_ix74_ix4008 : dff port map ( Q=>OPEN, QB=>nx11092, D=>nx249, 
      CLK=>nx15473);
   ix11096 : nand02 port map ( Y=>nx11095, A0=>nx10988, A1=>nx18);
   ix11098 : nand04 port map ( Y=>nx11097, A0=>nx10521, A1=>nx16165, A2=>
      address(0), A3=>nx16175);
   modgen_ram_ix74_ix4068 : dff port map ( Q=>OPEN, QB=>nx11099, D=>nx259, 
      CLK=>nx15475);
   ix11103 : nand02 port map ( Y=>nx11102, A0=>nx11012, A1=>nx52);
   ix11105 : nand03 port map ( Y=>nx11104, A0=>nx10613, A1=>nx10527, A2=>
      nx10663);
   tri_data_out_1 : tri01 port map ( Y=>data_out(1), A=>nx11107, E=>
      write_out);
   ix2003 : oai22 port map ( Y=>nx2002, A0=>nx11113, A1=>nx16157, B0=>
      nx11118, B1=>nx16183);
   modgen_ram_ix74_ix3755 : dff port map ( Q=>OPEN, QB=>nx11113, D=>nx1519, 
      CLK=>nx15475);
   modgen_ram_ix74_ix3863 : dff port map ( Q=>OPEN, QB=>nx11118, D=>nx1509, 
      CLK=>nx15475);
   modgen_ram_ix74_ix3839 : dff port map ( Q=>OPEN, QB=>nx11122, D=>nx1489, 
      CLK=>nx15475);
   modgen_ram_ix74_ix3847 : dff port map ( Q=>OPEN, QB=>nx11125, D=>nx1499, 
      CLK=>nx15475);
   ix11129 : nor02_2x port map ( Y=>nx11128, A0=>nx1964, A1=>nx1946);
   ix1965 : oai33 port map ( Y=>nx1964, A0=>nx11131, A1=>nx15849, A2=>
      nx16093, B0=>nx11134, B1=>nx15417, B2=>nx16021);
   modgen_ram_ix74_ix3947 : dff port map ( Q=>OPEN, QB=>nx11131, D=>nx1469, 
      CLK=>nx15475);
   modgen_ram_ix74_ix3759 : dff port map ( Q=>OPEN, QB=>nx11134, D=>nx1479, 
      CLK=>nx15475);
   ix1947 : oai22 port map ( Y=>nx1946, A0=>nx11138, A1=>nx16259, B0=>
      nx11141, B1=>nx16275);
   modgen_ram_ix74_ix3883 : dff port map ( Q=>OPEN, QB=>nx11138, D=>nx1459, 
      CLK=>nx15477);
   modgen_ram_ix74_ix3819 : dff port map ( Q=>OPEN, QB=>nx11141, D=>nx1449, 
      CLK=>nx15477);
   ix11145 : nor03_2x port map ( Y=>nx11144, A0=>nx1922, A1=>nx1914, A2=>
      nx1906);
   ix1923 : nor03_2x port map ( Y=>nx1922, A0=>nx11147, A1=>nx15761, A2=>
      nx16061);
   modgen_ram_ix74_ix3775 : dff port map ( Q=>OPEN, QB=>nx11147, D=>nx1439, 
      CLK=>nx15477);
   ix1915 : nor03_2x port map ( Y=>nx1914, A0=>nx11151, A1=>nx15849, A2=>
      nx15403);
   modgen_ram_ix74_ix3943 : dff port map ( Q=>OPEN, QB=>nx11151, D=>nx1429, 
      CLK=>nx15477);
   ix1907 : oai33 port map ( Y=>nx1906, A0=>nx11155, A1=>nx15761, A2=>
      nx15911, B0=>nx11158, B1=>nx15417, B2=>nx16061);
   modgen_ram_ix74_ix3783 : dff port map ( Q=>OPEN, QB=>nx11155, D=>nx1409, 
      CLK=>nx15477);
   modgen_ram_ix74_ix3711 : dff port map ( Q=>OPEN, QB=>nx11158, D=>nx1419, 
      CLK=>nx15477);
   ix11162 : nor03_2x port map ( Y=>nx11161, A0=>nx1884, A1=>nx1876, A2=>
      nx1868);
   ix1885 : nor03_2x port map ( Y=>nx1884, A0=>nx11164, A1=>nx15761, A2=>
      nx16039);
   modgen_ram_ix74_ix3779 : dff port map ( Q=>OPEN, QB=>nx11164, D=>nx1399, 
      CLK=>nx15477);
   ix1877 : nor04 port map ( Y=>nx1876, A0=>nx11168, A1=>address(4), A2=>
      address(5), A3=>nx16061);
   modgen_ram_ix74_ix3903 : dff port map ( Q=>OPEN, QB=>nx11168, D=>nx1389, 
      CLK=>nx15479);
   ix1869 : oai22 port map ( Y=>nx1868, A0=>nx11172, A1=>nx16327, B0=>
      nx11175, B1=>nx16343);
   modgen_ram_ix74_ix3719 : dff port map ( Q=>OPEN, QB=>nx11172, D=>nx1369, 
      CLK=>nx15479);
   modgen_ram_ix74_ix3715 : dff port map ( Q=>OPEN, QB=>nx11175, D=>nx1379, 
      CLK=>nx15479);
   modgen_ram_ix74_ix3843 : dff port map ( Q=>OPEN, QB=>nx11182, D=>nx1359, 
      CLK=>nx15479);
   modgen_ram_ix74_ix3907 : dff port map ( Q=>OPEN, QB=>nx11186, D=>nx1349, 
      CLK=>nx15479);
   ix1827 : oai22 port map ( Y=>nx1826, A0=>nx11190, A1=>nx16359, B0=>
      nx11193, B1=>nx16375);
   modgen_ram_ix74_ix3887 : dff port map ( Q=>OPEN, QB=>nx11190, D=>nx1329, 
      CLK=>nx15479);
   modgen_ram_ix74_ix3823 : dff port map ( Q=>OPEN, QB=>nx11193, D=>nx1339, 
      CLK=>nx15479);
   modgen_ram_ix74_ix3951 : dff port map ( Q=>OPEN, QB=>nx11199, D=>nx1319, 
      CLK=>nx15481);
   modgen_ram_ix74_ix3763 : dff port map ( Q=>OPEN, QB=>nx11203, D=>nx1309, 
      CLK=>nx15481);
   ix1789 : oai22 port map ( Y=>nx1788, A0=>nx11207, A1=>nx16399, B0=>
      nx11210, B1=>nx16415);
   modgen_ram_ix74_ix3891 : dff port map ( Q=>OPEN, QB=>nx11207, D=>nx1289, 
      CLK=>nx15481);
   modgen_ram_ix74_ix3827 : dff port map ( Q=>OPEN, QB=>nx11210, D=>nx1299, 
      CLK=>nx15481);
   modgen_ram_ix74_ix3955 : dff port map ( Q=>OPEN, QB=>nx11216, D=>nx1279, 
      CLK=>nx15481);
   modgen_ram_ix74_ix3767 : dff port map ( Q=>OPEN, QB=>nx11220, D=>nx1269, 
      CLK=>nx15481);
   modgen_ram_ix74_ix3895 : dff port map ( Q=>OPEN, QB=>nx11224, D=>nx1249, 
      CLK=>nx15481);
   modgen_ram_ix74_ix3831 : dff port map ( Q=>OPEN, QB=>nx11227, D=>nx1259, 
      CLK=>nx15483);
   modgen_ram_ix74_ix3959 : dff port map ( Q=>OPEN, QB=>nx11233, D=>nx1239, 
      CLK=>nx15483);
   ix1719 : nor03_2x port map ( Y=>nx1718, A0=>nx11237, A1=>nx15417, A2=>
      nx15959);
   modgen_ram_ix74_ix3771 : dff port map ( Q=>OPEN, QB=>nx11237, D=>nx1229, 
      CLK=>nx15483);
   modgen_ram_ix74_ix3899 : dff port map ( Q=>OPEN, QB=>nx11241, D=>nx1209, 
      CLK=>nx15483);
   modgen_ram_ix74_ix3835 : dff port map ( Q=>OPEN, QB=>nx11244, D=>nx1219, 
      CLK=>nx15483);
   ix1685 : oai22 port map ( Y=>nx1684, A0=>nx11254, A1=>nx16511, B0=>
      nx11257, B1=>nx16519);
   modgen_ram_ix74_ix3927 : dff port map ( Q=>OPEN, QB=>nx11254, D=>nx1189, 
      CLK=>nx15483);
   modgen_ram_ix74_ix3963 : dff port map ( Q=>OPEN, QB=>nx11257, D=>nx1199, 
      CLK=>nx15483);
   ix1667 : oai22 port map ( Y=>nx1666, A0=>nx11261, A1=>nx16527, B0=>
      nx11264, B1=>nx16543);
   modgen_ram_ix74_ix3859 : dff port map ( Q=>OPEN, QB=>nx11261, D=>nx1179, 
      CLK=>nx15485);
   modgen_ram_ix74_ix3795 : dff port map ( Q=>OPEN, QB=>nx11264, D=>nx1169, 
      CLK=>nx15485);
   ix1649 : nand03 port map ( Y=>nx1648, A0=>nx11268, A1=>nx11278, A2=>
      nx11284);
   ix11269 : nor02_2x port map ( Y=>nx11268, A0=>nx1644, A1=>nx1636);
   ix1645 : nor04 port map ( Y=>nx1644, A0=>nx11271, A1=>address(4), A2=>
      address(5), A3=>nx15895);
   modgen_ram_ix74_ix3919 : dff port map ( Q=>OPEN, QB=>nx11271, D=>nx1159, 
      CLK=>nx15485);
   ix1637 : nor03_2x port map ( Y=>nx1636, A0=>nx11275, A1=>nx15819, A2=>
      nx15895);
   modgen_ram_ix74_ix3855 : dff port map ( Q=>OPEN, QB=>nx11275, D=>nx1149, 
      CLK=>nx15485);
   ix11279 : nand03 port map ( Y=>nx11278, A0=>modgen_ram_ix74_a_12_dup_1142, 
      A1=>nx16229, A2=>nx16567);
   modgen_ram_ix74_ix3915 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_1142, 
      QB=>nx11282, D=>nx1139, CLK=>nx15485);
   ix11285 : nand03 port map ( Y=>nx11284, A0=>modgen_ram_ix74_a_28_dup_1126, 
      A1=>nx16195, A2=>nx16567);
   modgen_ram_ix74_ix3851 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_1126, 
      QB=>nx11288, D=>nx1129, CLK=>nx15485);
   modgen_ram_ix74_ix3723 : dff port map ( Q=>OPEN, QB=>nx11293, D=>nx1119, 
      CLK=>nx15485);
   modgen_ram_ix74_ix3799 : dff port map ( Q=>OPEN, QB=>nx11297, D=>nx1109, 
      CLK=>nx15487);
   modgen_ram_ix74_ix3791 : dff port map ( Q=>OPEN, QB=>nx11301, D=>nx1099, 
      CLK=>nx15487);
   modgen_ram_ix74_ix3787 : dff port map ( Q=>OPEN, QB=>nx11304, D=>nx1089, 
      CLK=>nx15487);
   ix11308 : nor03_2x port map ( Y=>nx11307, A0=>nx1566, A1=>nx1558, A2=>
      nx1550);
   ix1567 : nor03_2x port map ( Y=>nx1566, A0=>nx11310, A1=>nx15851, A2=>
      nx15911);
   modgen_ram_ix74_ix3911 : dff port map ( Q=>OPEN, QB=>nx11310, D=>nx1079, 
      CLK=>nx15487);
   ix1559 : nor03_2x port map ( Y=>nx1558, A0=>nx11314, A1=>nx15419, A2=>
      nx15895);
   modgen_ram_ix74_ix3727 : dff port map ( Q=>OPEN, QB=>nx11314, D=>nx1069, 
      CLK=>nx15487);
   ix1551 : oai22 port map ( Y=>nx1550, A0=>nx11318, A1=>nx16643, B0=>
      nx11321, B1=>nx16659);
   modgen_ram_ix74_ix3735 : dff port map ( Q=>OPEN, QB=>nx11318, D=>nx1059, 
      CLK=>nx15487);
   modgen_ram_ix74_ix3731 : dff port map ( Q=>OPEN, QB=>nx11321, D=>nx1049, 
      CLK=>nx15487);
   ix1527 : oai22 port map ( Y=>nx1526, A0=>nx11328, A1=>nx16675, B0=>
      nx11331, B1=>nx16691);
   modgen_ram_ix74_ix3879 : dff port map ( Q=>OPEN, QB=>nx11328, D=>nx1029, 
      CLK=>nx15489);
   modgen_ram_ix74_ix3923 : dff port map ( Q=>OPEN, QB=>nx11331, D=>nx1039, 
      CLK=>nx15489);
   ix1509 : oai22 port map ( Y=>nx1508, A0=>nx11335, A1=>nx16707, B0=>
      nx11338, B1=>nx16723);
   modgen_ram_ix74_ix3939 : dff port map ( Q=>OPEN, QB=>nx11335, D=>nx1019, 
      CLK=>nx15489);
   modgen_ram_ix74_ix3875 : dff port map ( Q=>OPEN, QB=>nx11338, D=>nx1009, 
      CLK=>nx15489);
   ix11342 : nor03_2x port map ( Y=>nx11341, A0=>nx1486, A1=>nx1478, A2=>
      nx1470);
   ix1487 : nor03_2x port map ( Y=>nx1486, A0=>nx11344, A1=>nx15419, A2=>
      nx15753);
   modgen_ram_ix74_ix3747 : dff port map ( Q=>OPEN, QB=>nx11344, D=>nx999, 
      CLK=>nx15489);
   ix1479 : nor03_2x port map ( Y=>nx1478, A0=>nx11348, A1=>nx15851, A2=>
      nx15797);
   modgen_ram_ix74_ix3935 : dff port map ( Q=>OPEN, QB=>nx11348, D=>nx989, 
      CLK=>nx15489);
   ix1471 : oai22 port map ( Y=>nx1470, A0=>nx11352, A1=>nx16747, B0=>
      nx11355, B1=>nx16755);
   modgen_ram_ix74_ix3743 : dff port map ( Q=>OPEN, QB=>nx11352, D=>nx979, 
      CLK=>nx15489);
   modgen_ram_ix74_ix3931 : dff port map ( Q=>OPEN, QB=>nx11355, D=>nx969, 
      CLK=>nx15491);
   ix11359 : nor03_2x port map ( Y=>nx11358, A0=>nx1446, A1=>nx1438, A2=>
      nx1430);
   ix1447 : nor03_2x port map ( Y=>nx1446, A0=>nx11361, A1=>nx15761, A2=>
      nx15813);
   modgen_ram_ix74_ix3803 : dff port map ( Q=>OPEN, QB=>nx11361, D=>nx959, 
      CLK=>nx15491);
   ix1439 : nor03_2x port map ( Y=>nx1438, A0=>nx11365, A1=>nx15819, A2=>
      nx15797);
   modgen_ram_ix74_ix3871 : dff port map ( Q=>OPEN, QB=>nx11365, D=>nx949, 
      CLK=>nx15491);
   ix1431 : oai22 port map ( Y=>nx1430, A0=>nx11369, A1=>nx16771, B0=>
      nx11372, B1=>nx16787);
   modgen_ram_ix74_ix3867 : dff port map ( Q=>OPEN, QB=>nx11369, D=>nx939, 
      CLK=>nx15491);
   modgen_ram_ix74_ix3739 : dff port map ( Q=>OPEN, QB=>nx11372, D=>nx929, 
      CLK=>nx15491);
   ix11376 : nor03_2x port map ( Y=>nx11375, A0=>nx1408, A1=>nx1400, A2=>
      nx1392);
   ix1409 : nor03_2x port map ( Y=>nx1408, A0=>nx11378, A1=>nx15761, A2=>
      nx15799);
   modgen_ram_ix74_ix3807 : dff port map ( Q=>OPEN, QB=>nx11378, D=>nx919, 
      CLK=>nx15491);
   ix1401 : nor03_2x port map ( Y=>nx1400, A0=>nx11382, A1=>nx15763, A2=>
      nx15403);
   modgen_ram_ix74_ix3815 : dff port map ( Q=>OPEN, QB=>nx11382, D=>nx909, 
      CLK=>nx15491);
   ix1393 : oai22 port map ( Y=>nx1392, A0=>nx11386, A1=>nx16819, B0=>
      nx11389, B1=>nx16835);
   modgen_ram_ix74_ix3751 : dff port map ( Q=>OPEN, QB=>nx11386, D=>nx889, 
      CLK=>nx15493);
   modgen_ram_ix74_ix3811 : dff port map ( Q=>OPEN, QB=>nx11389, D=>nx899, 
      CLK=>nx15493);
   tri_data_out_2 : tri01 port map ( Y=>data_out(2), A=>nx11393, E=>
      write_out);
   ix2641 : oai22 port map ( Y=>nx2640, A0=>nx11399, A1=>nx16157, B0=>
      nx11404, B1=>nx16183);
   modgen_ram_ix74_ix3498 : dff port map ( Q=>OPEN, QB=>nx11399, D=>nx2159, 
      CLK=>nx15493);
   modgen_ram_ix74_ix3606 : dff port map ( Q=>OPEN, QB=>nx11404, D=>nx2149, 
      CLK=>nx15493);
   modgen_ram_ix74_ix3582 : dff port map ( Q=>OPEN, QB=>nx11408, D=>nx2129, 
      CLK=>nx15493);
   modgen_ram_ix74_ix3590 : dff port map ( Q=>OPEN, QB=>nx11411, D=>nx2139, 
      CLK=>nx15493);
   ix11415 : nor02_2x port map ( Y=>nx11414, A0=>nx2602, A1=>nx2584);
   ix2603 : oai33 port map ( Y=>nx2602, A0=>nx11417, A1=>nx15851, A2=>
      nx16093, B0=>nx11420, B1=>nx15419, B2=>nx16021);
   modgen_ram_ix74_ix3690 : dff port map ( Q=>OPEN, QB=>nx11417, D=>nx2109, 
      CLK=>nx15493);
   modgen_ram_ix74_ix3502 : dff port map ( Q=>OPEN, QB=>nx11420, D=>nx2119, 
      CLK=>nx15495);
   ix2585 : oai22 port map ( Y=>nx2584, A0=>nx11424, A1=>nx16259, B0=>
      nx11427, B1=>nx16275);
   modgen_ram_ix74_ix3626 : dff port map ( Q=>OPEN, QB=>nx11424, D=>nx2099, 
      CLK=>nx15495);
   modgen_ram_ix74_ix3562 : dff port map ( Q=>OPEN, QB=>nx11427, D=>nx2089, 
      CLK=>nx15495);
   ix11431 : nor03_2x port map ( Y=>nx11430, A0=>nx2560, A1=>nx2552, A2=>
      nx2544);
   ix2561 : nor03_2x port map ( Y=>nx2560, A0=>nx11433, A1=>nx15763, A2=>
      nx16061);
   modgen_ram_ix74_ix3518 : dff port map ( Q=>OPEN, QB=>nx11433, D=>nx2079, 
      CLK=>nx15495);
   ix2553 : nor03_2x port map ( Y=>nx2552, A0=>nx11437, A1=>nx15851, A2=>
      nx15403);
   modgen_ram_ix74_ix3686 : dff port map ( Q=>OPEN, QB=>nx11437, D=>nx2069, 
      CLK=>nx15495);
   ix2545 : oai33 port map ( Y=>nx2544, A0=>nx11441, A1=>nx15763, A2=>
      nx15911, B0=>nx11444, B1=>nx15419, B2=>nx16063);
   modgen_ram_ix74_ix3526 : dff port map ( Q=>OPEN, QB=>nx11441, D=>nx2049, 
      CLK=>nx15495);
   modgen_ram_ix74_ix3454 : dff port map ( Q=>OPEN, QB=>nx11444, D=>nx2059, 
      CLK=>nx15495);
   ix11448 : nor03_2x port map ( Y=>nx11447, A0=>nx2522, A1=>nx2514, A2=>
      nx2506);
   ix2523 : nor03_2x port map ( Y=>nx2522, A0=>nx11450, A1=>nx15763, A2=>
      nx16041);
   modgen_ram_ix74_ix3522 : dff port map ( Q=>OPEN, QB=>nx11450, D=>nx2039, 
      CLK=>nx15497);
   ix2515 : nor04 port map ( Y=>nx2514, A0=>nx11454, A1=>address(4), A2=>
      address(5), A3=>nx16063);
   modgen_ram_ix74_ix3646 : dff port map ( Q=>OPEN, QB=>nx11454, D=>nx2029, 
      CLK=>nx15497);
   ix2507 : oai22 port map ( Y=>nx2506, A0=>nx11458, A1=>nx16327, B0=>
      nx11461, B1=>nx16343);
   modgen_ram_ix74_ix3462 : dff port map ( Q=>OPEN, QB=>nx11458, D=>nx2009, 
      CLK=>nx15497);
   modgen_ram_ix74_ix3458 : dff port map ( Q=>OPEN, QB=>nx11461, D=>nx2019, 
      CLK=>nx15497);
   modgen_ram_ix74_ix3586 : dff port map ( Q=>OPEN, QB=>nx11468, D=>nx1999, 
      CLK=>nx15497);
   modgen_ram_ix74_ix3650 : dff port map ( Q=>OPEN, QB=>nx11472, D=>nx1989, 
      CLK=>nx15497);
   ix2465 : oai22 port map ( Y=>nx2464, A0=>nx11476, A1=>nx16359, B0=>
      nx11479, B1=>nx16375);
   modgen_ram_ix74_ix3630 : dff port map ( Q=>OPEN, QB=>nx11476, D=>nx1969, 
      CLK=>nx15497);
   modgen_ram_ix74_ix3566 : dff port map ( Q=>OPEN, QB=>nx11479, D=>nx1979, 
      CLK=>nx15499);
   modgen_ram_ix74_ix3694 : dff port map ( Q=>OPEN, QB=>nx11485, D=>nx1959, 
      CLK=>nx15499);
   modgen_ram_ix74_ix3506 : dff port map ( Q=>OPEN, QB=>nx11489, D=>nx1949, 
      CLK=>nx15499);
   ix2427 : oai22 port map ( Y=>nx2426, A0=>nx11493, A1=>nx16399, B0=>
      nx11496, B1=>nx16415);
   modgen_ram_ix74_ix3634 : dff port map ( Q=>OPEN, QB=>nx11493, D=>nx1929, 
      CLK=>nx15499);
   modgen_ram_ix74_ix3570 : dff port map ( Q=>OPEN, QB=>nx11496, D=>nx1939, 
      CLK=>nx15499);
   modgen_ram_ix74_ix3698 : dff port map ( Q=>OPEN, QB=>nx11502, D=>nx1919, 
      CLK=>nx15499);
   modgen_ram_ix74_ix3510 : dff port map ( Q=>OPEN, QB=>nx11506, D=>nx1909, 
      CLK=>nx15499);
   modgen_ram_ix74_ix3638 : dff port map ( Q=>OPEN, QB=>nx11510, D=>nx1889, 
      CLK=>nx15501);
   modgen_ram_ix74_ix3574 : dff port map ( Q=>OPEN, QB=>nx11513, D=>nx1899, 
      CLK=>nx15501);
   modgen_ram_ix74_ix3702 : dff port map ( Q=>OPEN, QB=>nx11519, D=>nx1879, 
      CLK=>nx15501);
   ix2357 : nor03_2x port map ( Y=>nx2356, A0=>nx11523, A1=>nx15421, A2=>
      nx15959);
   modgen_ram_ix74_ix3514 : dff port map ( Q=>OPEN, QB=>nx11523, D=>nx1869, 
      CLK=>nx15501);
   modgen_ram_ix74_ix3642 : dff port map ( Q=>OPEN, QB=>nx11527, D=>nx1849, 
      CLK=>nx15501);
   modgen_ram_ix74_ix3578 : dff port map ( Q=>OPEN, QB=>nx11530, D=>nx1859, 
      CLK=>nx15501);
   ix2323 : oai22 port map ( Y=>nx2322, A0=>nx11540, A1=>nx16511, B0=>
      nx11543, B1=>nx16519);
   modgen_ram_ix74_ix3670 : dff port map ( Q=>OPEN, QB=>nx11540, D=>nx1829, 
      CLK=>nx15501);
   modgen_ram_ix74_ix3706 : dff port map ( Q=>OPEN, QB=>nx11543, D=>nx1839, 
      CLK=>nx15503);
   ix2305 : oai22 port map ( Y=>nx2304, A0=>nx11547, A1=>nx16527, B0=>
      nx11550, B1=>nx16543);
   modgen_ram_ix74_ix3602 : dff port map ( Q=>OPEN, QB=>nx11547, D=>nx1819, 
      CLK=>nx15503);
   modgen_ram_ix74_ix3538 : dff port map ( Q=>OPEN, QB=>nx11550, D=>nx1809, 
      CLK=>nx15503);
   ix2287 : nand03 port map ( Y=>nx2286, A0=>nx11554, A1=>nx11564, A2=>
      nx11570);
   ix11555 : nor02_2x port map ( Y=>nx11554, A0=>nx2282, A1=>nx2274);
   ix2283 : nor04 port map ( Y=>nx2282, A0=>nx11557, A1=>address(4), A2=>
      address(5), A3=>nx15897);
   modgen_ram_ix74_ix3662 : dff port map ( Q=>OPEN, QB=>nx11557, D=>nx1799, 
      CLK=>nx15503);
   ix2275 : nor03_2x port map ( Y=>nx2274, A0=>nx11561, A1=>nx15821, A2=>
      nx15897);
   modgen_ram_ix74_ix3598 : dff port map ( Q=>OPEN, QB=>nx11561, D=>nx1789, 
      CLK=>nx15503);
   ix11565 : nand03 port map ( Y=>nx11564, A0=>modgen_ram_ix74_a_12_dup_1076, 
      A1=>nx16229, A2=>nx16569);
   modgen_ram_ix74_ix3658 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_1076, 
      QB=>nx11568, D=>nx1779, CLK=>nx15503);
   ix11571 : nand03 port map ( Y=>nx11570, A0=>modgen_ram_ix74_a_28_dup_1060, 
      A1=>nx16195, A2=>nx16569);
   modgen_ram_ix74_ix3594 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_1060, 
      QB=>nx11574, D=>nx1769, CLK=>nx15503);
   modgen_ram_ix74_ix3466 : dff port map ( Q=>OPEN, QB=>nx11579, D=>nx1759, 
      CLK=>nx15505);
   modgen_ram_ix74_ix3542 : dff port map ( Q=>OPEN, QB=>nx11583, D=>nx1749, 
      CLK=>nx15505);
   modgen_ram_ix74_ix3534 : dff port map ( Q=>OPEN, QB=>nx11587, D=>nx1739, 
      CLK=>nx15505);
   modgen_ram_ix74_ix3530 : dff port map ( Q=>OPEN, QB=>nx11590, D=>nx1729, 
      CLK=>nx15505);
   ix11594 : nor03_2x port map ( Y=>nx11593, A0=>nx2204, A1=>nx2196, A2=>
      nx2188);
   ix2205 : nor03_2x port map ( Y=>nx2204, A0=>nx11596, A1=>nx15851, A2=>
      nx15913);
   modgen_ram_ix74_ix3654 : dff port map ( Q=>OPEN, QB=>nx11596, D=>nx1719, 
      CLK=>nx15505);
   ix2197 : nor03_2x port map ( Y=>nx2196, A0=>nx11600, A1=>nx15421, A2=>
      nx15897);
   modgen_ram_ix74_ix3470 : dff port map ( Q=>OPEN, QB=>nx11600, D=>nx1709, 
      CLK=>nx15505);
   ix2189 : oai22 port map ( Y=>nx2188, A0=>nx11604, A1=>nx16643, B0=>
      nx11607, B1=>nx16659);
   modgen_ram_ix74_ix3478 : dff port map ( Q=>OPEN, QB=>nx11604, D=>nx1699, 
      CLK=>nx15505);
   modgen_ram_ix74_ix3474 : dff port map ( Q=>OPEN, QB=>nx11607, D=>nx1689, 
      CLK=>nx15507);
   ix2165 : oai22 port map ( Y=>nx2164, A0=>nx11614, A1=>nx16675, B0=>
      nx11617, B1=>nx16691);
   modgen_ram_ix74_ix3622 : dff port map ( Q=>OPEN, QB=>nx11614, D=>nx1669, 
      CLK=>nx15507);
   modgen_ram_ix74_ix3666 : dff port map ( Q=>OPEN, QB=>nx11617, D=>nx1679, 
      CLK=>nx15507);
   ix2147 : oai22 port map ( Y=>nx2146, A0=>nx11621, A1=>nx16707, B0=>
      nx11624, B1=>nx16723);
   modgen_ram_ix74_ix3682 : dff port map ( Q=>OPEN, QB=>nx11621, D=>nx1659, 
      CLK=>nx15507);
   modgen_ram_ix74_ix3618 : dff port map ( Q=>OPEN, QB=>nx11624, D=>nx1649, 
      CLK=>nx15507);
   ix11628 : nor03_2x port map ( Y=>nx11627, A0=>nx2124, A1=>nx2116, A2=>
      nx2108);
   ix2125 : nor03_2x port map ( Y=>nx2124, A0=>nx11630, A1=>nx15421, A2=>
      nx15753);
   modgen_ram_ix74_ix3490 : dff port map ( Q=>OPEN, QB=>nx11630, D=>nx1639, 
      CLK=>nx15507);
   ix2117 : nor03_2x port map ( Y=>nx2116, A0=>nx11634, A1=>nx15853, A2=>
      nx15799);
   modgen_ram_ix74_ix3678 : dff port map ( Q=>OPEN, QB=>nx11634, D=>nx1629, 
      CLK=>nx15507);
   ix2109 : oai22 port map ( Y=>nx2108, A0=>nx11638, A1=>nx16747, B0=>
      nx11641, B1=>nx16755);
   modgen_ram_ix74_ix3486 : dff port map ( Q=>OPEN, QB=>nx11638, D=>nx1619, 
      CLK=>nx15509);
   modgen_ram_ix74_ix3674 : dff port map ( Q=>OPEN, QB=>nx11641, D=>nx1609, 
      CLK=>nx15509);
   ix11645 : nor03_2x port map ( Y=>nx11644, A0=>nx2084, A1=>nx2076, A2=>
      nx2068);
   ix2085 : nor03_2x port map ( Y=>nx2084, A0=>nx11647, A1=>nx15763, A2=>
      nx15813);
   modgen_ram_ix74_ix3546 : dff port map ( Q=>OPEN, QB=>nx11647, D=>nx1599, 
      CLK=>nx15509);
   ix2077 : nor03_2x port map ( Y=>nx2076, A0=>nx11651, A1=>nx15821, A2=>
      nx15799);
   modgen_ram_ix74_ix3614 : dff port map ( Q=>OPEN, QB=>nx11651, D=>nx1589, 
      CLK=>nx15509);
   ix2069 : oai22 port map ( Y=>nx2068, A0=>nx11655, A1=>nx16771, B0=>
      nx11658, B1=>nx16787);
   modgen_ram_ix74_ix3610 : dff port map ( Q=>OPEN, QB=>nx11655, D=>nx1579, 
      CLK=>nx15509);
   modgen_ram_ix74_ix3482 : dff port map ( Q=>OPEN, QB=>nx11658, D=>nx1569, 
      CLK=>nx15509);
   ix11662 : nor03_2x port map ( Y=>nx11661, A0=>nx2046, A1=>nx2038, A2=>
      nx2030);
   ix2047 : nor03_2x port map ( Y=>nx2046, A0=>nx11664, A1=>nx15763, A2=>
      nx15799);
   modgen_ram_ix74_ix3550 : dff port map ( Q=>OPEN, QB=>nx11664, D=>nx1559, 
      CLK=>nx15509);
   ix2039 : nor03_2x port map ( Y=>nx2038, A0=>nx11668, A1=>nx15765, A2=>
      nx15403);
   modgen_ram_ix74_ix3558 : dff port map ( Q=>OPEN, QB=>nx11668, D=>nx1549, 
      CLK=>nx15511);
   ix2031 : oai22 port map ( Y=>nx2030, A0=>nx11672, A1=>nx16819, B0=>
      nx11675, B1=>nx16835);
   modgen_ram_ix74_ix3494 : dff port map ( Q=>OPEN, QB=>nx11672, D=>nx1529, 
      CLK=>nx15511);
   modgen_ram_ix74_ix3554 : dff port map ( Q=>OPEN, QB=>nx11675, D=>nx1539, 
      CLK=>nx15511);
   tri_data_out_3 : tri01 port map ( Y=>data_out(3), A=>nx11679, E=>
      write_out);
   ix3279 : oai22 port map ( Y=>nx3278, A0=>nx11685, A1=>nx16157, B0=>
      nx11690, B1=>nx16183);
   modgen_ram_ix74_ix3241 : dff port map ( Q=>OPEN, QB=>nx11685, D=>nx2799, 
      CLK=>nx15511);
   modgen_ram_ix74_ix3349 : dff port map ( Q=>OPEN, QB=>nx11690, D=>nx2789, 
      CLK=>nx15511);
   ix3261 : oai22 port map ( Y=>nx3260, A0=>nx11694, A1=>nx16201, B0=>
      nx11697, B1=>nx18957);
   modgen_ram_ix74_ix3325 : dff port map ( Q=>OPEN, QB=>nx11694, D=>nx2769, 
      CLK=>nx15511);
   modgen_ram_ix74_ix3333 : dff port map ( Q=>OPEN, QB=>nx11697, D=>nx2779, 
      CLK=>nx15511);
   ix11701 : nor02_2x port map ( Y=>nx11700, A0=>nx3240, A1=>nx3222);
   ix3241 : oai33 port map ( Y=>nx3240, A0=>nx11703, A1=>nx15853, A2=>
      nx16093, B0=>nx11706, B1=>nx15421, B2=>nx16023);
   modgen_ram_ix74_ix3433 : dff port map ( Q=>OPEN, QB=>nx11703, D=>nx2749, 
      CLK=>nx15513);
   modgen_ram_ix74_ix3245 : dff port map ( Q=>OPEN, QB=>nx11706, D=>nx2759, 
      CLK=>nx15513);
   ix3223 : oai22 port map ( Y=>nx3222, A0=>nx11710, A1=>nx16259, B0=>
      nx11713, B1=>nx16275);
   modgen_ram_ix74_ix3369 : dff port map ( Q=>OPEN, QB=>nx11710, D=>nx2739, 
      CLK=>nx15513);
   modgen_ram_ix74_ix3305 : dff port map ( Q=>OPEN, QB=>nx11713, D=>nx2729, 
      CLK=>nx15513);
   ix11717 : nor03_2x port map ( Y=>nx11716, A0=>nx3198, A1=>nx3190, A2=>
      nx3182);
   ix3199 : nor03_2x port map ( Y=>nx3198, A0=>nx11719, A1=>nx15765, A2=>
      nx16063);
   modgen_ram_ix74_ix3261 : dff port map ( Q=>OPEN, QB=>nx11719, D=>nx2719, 
      CLK=>nx15513);
   ix3191 : nor03_2x port map ( Y=>nx3190, A0=>nx11723, A1=>nx15853, A2=>
      nx15405);
   modgen_ram_ix74_ix3429 : dff port map ( Q=>OPEN, QB=>nx11723, D=>nx2709, 
      CLK=>nx15513);
   ix3183 : oai33 port map ( Y=>nx3182, A0=>nx11727, A1=>nx15765, A2=>
      nx15913, B0=>nx11730, B1=>nx15421, B2=>nx16063);
   modgen_ram_ix74_ix3269 : dff port map ( Q=>OPEN, QB=>nx11727, D=>nx2689, 
      CLK=>nx15513);
   modgen_ram_ix74_ix3197 : dff port map ( Q=>OPEN, QB=>nx11730, D=>nx2699, 
      CLK=>nx15515);
   ix11734 : nor03_2x port map ( Y=>nx11733, A0=>nx3160, A1=>nx3152, A2=>
      nx3144);
   ix3161 : nor03_2x port map ( Y=>nx3160, A0=>nx11736, A1=>nx15765, A2=>
      nx16041);
   modgen_ram_ix74_ix3265 : dff port map ( Q=>OPEN, QB=>nx11736, D=>nx2679, 
      CLK=>nx15515);
   ix3153 : nor04 port map ( Y=>nx3152, A0=>nx11740, A1=>address(4), A2=>
      address(5), A3=>nx16063);
   modgen_ram_ix74_ix3389 : dff port map ( Q=>OPEN, QB=>nx11740, D=>nx2669, 
      CLK=>nx15515);
   ix3145 : oai22 port map ( Y=>nx3144, A0=>nx11744, A1=>nx16327, B0=>
      nx11747, B1=>nx16343);
   modgen_ram_ix74_ix3205 : dff port map ( Q=>OPEN, QB=>nx11744, D=>nx2649, 
      CLK=>nx15515);
   modgen_ram_ix74_ix3201 : dff port map ( Q=>OPEN, QB=>nx11747, D=>nx2659, 
      CLK=>nx15515);
   modgen_ram_ix74_ix3329 : dff port map ( Q=>OPEN, QB=>nx11754, D=>nx2639, 
      CLK=>nx15515);
   modgen_ram_ix74_ix3393 : dff port map ( Q=>OPEN, QB=>nx11758, D=>nx2629, 
      CLK=>nx15515);
   ix3103 : oai22 port map ( Y=>nx3102, A0=>nx11762, A1=>nx16359, B0=>
      nx11765, B1=>nx16375);
   modgen_ram_ix74_ix3373 : dff port map ( Q=>OPEN, QB=>nx11762, D=>nx2609, 
      CLK=>nx15517);
   modgen_ram_ix74_ix3309 : dff port map ( Q=>OPEN, QB=>nx11765, D=>nx2619, 
      CLK=>nx15517);
   modgen_ram_ix74_ix3437 : dff port map ( Q=>OPEN, QB=>nx11771, D=>nx2599, 
      CLK=>nx15517);
   modgen_ram_ix74_ix3249 : dff port map ( Q=>OPEN, QB=>nx11775, D=>nx2589, 
      CLK=>nx15517);
   ix3065 : oai22 port map ( Y=>nx3064, A0=>nx11779, A1=>nx16399, B0=>
      nx11782, B1=>nx16415);
   modgen_ram_ix74_ix3377 : dff port map ( Q=>OPEN, QB=>nx11779, D=>nx2569, 
      CLK=>nx15517);
   modgen_ram_ix74_ix3313 : dff port map ( Q=>OPEN, QB=>nx11782, D=>nx2579, 
      CLK=>nx15517);
   modgen_ram_ix74_ix3441 : dff port map ( Q=>OPEN, QB=>nx11788, D=>nx2559, 
      CLK=>nx15517);
   modgen_ram_ix74_ix3253 : dff port map ( Q=>OPEN, QB=>nx11792, D=>nx2549, 
      CLK=>nx15519);
   ix3025 : oai22 port map ( Y=>nx3024, A0=>nx11796, A1=>nx16439, B0=>
      nx11799, B1=>nx16455);
   modgen_ram_ix74_ix3381 : dff port map ( Q=>OPEN, QB=>nx11796, D=>nx2529, 
      CLK=>nx15519);
   modgen_ram_ix74_ix3317 : dff port map ( Q=>OPEN, QB=>nx11799, D=>nx2539, 
      CLK=>nx15519);
   modgen_ram_ix74_ix3445 : dff port map ( Q=>OPEN, QB=>nx11805, D=>nx2519, 
      CLK=>nx15519);
   ix2995 : nor03_2x port map ( Y=>nx2994, A0=>nx11809, A1=>nx15423, A2=>
      nx15959);
   modgen_ram_ix74_ix3257 : dff port map ( Q=>OPEN, QB=>nx11809, D=>nx2509, 
      CLK=>nx15519);
   ix2987 : oai22 port map ( Y=>nx2986, A0=>nx11813, A1=>nx16479, B0=>
      nx11816, B1=>nx16495);
   modgen_ram_ix74_ix3385 : dff port map ( Q=>OPEN, QB=>nx11813, D=>nx2489, 
      CLK=>nx15519);
   modgen_ram_ix74_ix3321 : dff port map ( Q=>OPEN, QB=>nx11816, D=>nx2499, 
      CLK=>nx15519);
   ix2961 : oai22 port map ( Y=>nx2960, A0=>nx11826, A1=>nx16511, B0=>
      nx11829, B1=>nx16519);
   modgen_ram_ix74_ix3413 : dff port map ( Q=>OPEN, QB=>nx11826, D=>nx2469, 
      CLK=>nx15521);
   modgen_ram_ix74_ix3449 : dff port map ( Q=>OPEN, QB=>nx11829, D=>nx2479, 
      CLK=>nx15521);
   ix2943 : oai22 port map ( Y=>nx2942, A0=>nx11833, A1=>nx16527, B0=>
      nx11836, B1=>nx16543);
   modgen_ram_ix74_ix3345 : dff port map ( Q=>OPEN, QB=>nx11833, D=>nx2459, 
      CLK=>nx15521);
   modgen_ram_ix74_ix3281 : dff port map ( Q=>OPEN, QB=>nx11836, D=>nx2449, 
      CLK=>nx15521);
   ix2925 : nand03 port map ( Y=>nx2924, A0=>nx11840, A1=>nx11850, A2=>
      nx11856);
   ix11841 : nor02_2x port map ( Y=>nx11840, A0=>nx2920, A1=>nx2912);
   ix2921 : nor04 port map ( Y=>nx2920, A0=>nx11843, A1=>address(4), A2=>
      address(5), A3=>nx15897);
   modgen_ram_ix74_ix3405 : dff port map ( Q=>OPEN, QB=>nx11843, D=>nx2439, 
      CLK=>nx15521);
   ix2913 : nor03_2x port map ( Y=>nx2912, A0=>nx11847, A1=>nx15821, A2=>
      nx15897);
   modgen_ram_ix74_ix3341 : dff port map ( Q=>OPEN, QB=>nx11847, D=>nx2429, 
      CLK=>nx15521);
   ix11851 : nand03 port map ( Y=>nx11850, A0=>modgen_ram_ix74_a_12_dup_1011, 
      A1=>nx16229, A2=>nx16569);
   modgen_ram_ix74_ix3401 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_1011, 
      QB=>nx11854, D=>nx2419, CLK=>nx15521);
   ix11857 : nand03 port map ( Y=>nx11856, A0=>modgen_ram_ix74_a_28_dup_995, 
      A1=>nx16195, A2=>nx16569);
   modgen_ram_ix74_ix3337 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_995, 
      QB=>nx11860, D=>nx2409, CLK=>nx15523);
   ix11863 : nor03_2x port map ( Y=>nx11862, A0=>nx2880, A1=>nx2872, A2=>
      nx2864);
   ix2881 : nor03_2x port map ( Y=>nx2880, A0=>nx11865, A1=>nx15423, A2=>
      nx15929);
   modgen_ram_ix74_ix3209 : dff port map ( Q=>OPEN, QB=>nx11865, D=>nx2399, 
      CLK=>nx15523);
   ix2873 : nor03_2x port map ( Y=>nx2872, A0=>nx11869, A1=>nx15765, A2=>
      nx15889);
   modgen_ram_ix74_ix3285 : dff port map ( Q=>OPEN, QB=>nx11869, D=>nx2389, 
      CLK=>nx15523);
   ix2865 : oai22 port map ( Y=>nx2864, A0=>nx11873, A1=>nx16603, B0=>
      nx11876, B1=>nx16619);
   modgen_ram_ix74_ix3277 : dff port map ( Q=>OPEN, QB=>nx11873, D=>nx2379, 
      CLK=>nx15523);
   modgen_ram_ix74_ix3273 : dff port map ( Q=>OPEN, QB=>nx11876, D=>nx2369, 
      CLK=>nx15523);
   ix11880 : nor03_2x port map ( Y=>nx11879, A0=>nx2842, A1=>nx2834, A2=>
      nx2826);
   ix2843 : nor03_2x port map ( Y=>nx2842, A0=>nx11882, A1=>nx15853, A2=>
      nx15913);
   modgen_ram_ix74_ix3397 : dff port map ( Q=>OPEN, QB=>nx11882, D=>nx2359, 
      CLK=>nx15523);
   ix2835 : nor03_2x port map ( Y=>nx2834, A0=>nx11886, A1=>nx15423, A2=>
      nx15897);
   modgen_ram_ix74_ix3213 : dff port map ( Q=>OPEN, QB=>nx11886, D=>nx2349, 
      CLK=>nx15523);
   ix2827 : oai22 port map ( Y=>nx2826, A0=>nx11890, A1=>nx16643, B0=>
      nx11893, B1=>nx16659);
   modgen_ram_ix74_ix3221 : dff port map ( Q=>OPEN, QB=>nx11890, D=>nx2339, 
      CLK=>nx15525);
   modgen_ram_ix74_ix3217 : dff port map ( Q=>OPEN, QB=>nx11893, D=>nx2329, 
      CLK=>nx15525);
   ix2803 : oai22 port map ( Y=>nx2802, A0=>nx11900, A1=>nx16675, B0=>
      nx11903, B1=>nx16691);
   modgen_ram_ix74_ix3365 : dff port map ( Q=>OPEN, QB=>nx11900, D=>nx2309, 
      CLK=>nx15525);
   modgen_ram_ix74_ix3409 : dff port map ( Q=>OPEN, QB=>nx11903, D=>nx2319, 
      CLK=>nx15525);
   ix2785 : oai22 port map ( Y=>nx2784, A0=>nx11907, A1=>nx16707, B0=>
      nx11910, B1=>nx16723);
   modgen_ram_ix74_ix3425 : dff port map ( Q=>OPEN, QB=>nx11907, D=>nx2299, 
      CLK=>nx15525);
   modgen_ram_ix74_ix3361 : dff port map ( Q=>OPEN, QB=>nx11910, D=>nx2289, 
      CLK=>nx15525);
   ix11914 : nor03_2x port map ( Y=>nx11913, A0=>nx2762, A1=>nx2754, A2=>
      nx2746);
   ix2763 : nor03_2x port map ( Y=>nx2762, A0=>nx11916, A1=>nx15423, A2=>
      nx15753);
   modgen_ram_ix74_ix3233 : dff port map ( Q=>OPEN, QB=>nx11916, D=>nx2279, 
      CLK=>nx15525);
   ix2755 : nor03_2x port map ( Y=>nx2754, A0=>nx11920, A1=>nx15853, A2=>
      nx15799);
   modgen_ram_ix74_ix3421 : dff port map ( Q=>OPEN, QB=>nx11920, D=>nx2269, 
      CLK=>nx15527);
   ix2747 : oai22 port map ( Y=>nx2746, A0=>nx11924, A1=>nx16747, B0=>
      nx11927, B1=>nx16755);
   modgen_ram_ix74_ix3229 : dff port map ( Q=>OPEN, QB=>nx11924, D=>nx2259, 
      CLK=>nx15527);
   modgen_ram_ix74_ix3417 : dff port map ( Q=>OPEN, QB=>nx11927, D=>nx2249, 
      CLK=>nx15527);
   ix11931 : nor03_2x port map ( Y=>nx11930, A0=>nx2722, A1=>nx2714, A2=>
      nx2706);
   ix2723 : nor03_2x port map ( Y=>nx2722, A0=>nx11933, A1=>nx15765, A2=>
      nx15813);
   modgen_ram_ix74_ix3289 : dff port map ( Q=>OPEN, QB=>nx11933, D=>nx2239, 
      CLK=>nx15527);
   ix2715 : nor03_2x port map ( Y=>nx2714, A0=>nx11937, A1=>nx15821, A2=>
      nx15799);
   modgen_ram_ix74_ix3357 : dff port map ( Q=>OPEN, QB=>nx11937, D=>nx2229, 
      CLK=>nx15527);
   ix2707 : oai22 port map ( Y=>nx2706, A0=>nx11941, A1=>nx16771, B0=>
      nx11944, B1=>nx16787);
   modgen_ram_ix74_ix3353 : dff port map ( Q=>OPEN, QB=>nx11941, D=>nx2219, 
      CLK=>nx15527);
   modgen_ram_ix74_ix3225 : dff port map ( Q=>OPEN, QB=>nx11944, D=>nx2209, 
      CLK=>nx15527);
   ix11948 : nor03_2x port map ( Y=>nx11947, A0=>nx2684, A1=>nx2676, A2=>
      nx2668);
   ix2685 : nor03_2x port map ( Y=>nx2684, A0=>nx11950, A1=>nx15765, A2=>
      nx15799);
   modgen_ram_ix74_ix3293 : dff port map ( Q=>OPEN, QB=>nx11950, D=>nx2199, 
      CLK=>nx15529);
   ix2677 : nor03_2x port map ( Y=>nx2676, A0=>nx11954, A1=>nx15767, A2=>
      nx15405);
   modgen_ram_ix74_ix3301 : dff port map ( Q=>OPEN, QB=>nx11954, D=>nx2189, 
      CLK=>nx15529);
   ix2669 : oai22 port map ( Y=>nx2668, A0=>nx11958, A1=>nx16819, B0=>
      nx11961, B1=>nx16835);
   modgen_ram_ix74_ix3237 : dff port map ( Q=>OPEN, QB=>nx11958, D=>nx2169, 
      CLK=>nx15529);
   modgen_ram_ix74_ix3297 : dff port map ( Q=>OPEN, QB=>nx11961, D=>nx2179, 
      CLK=>nx15529);
   tri_data_out_4 : tri01 port map ( Y=>data_out(4), A=>nx11965, E=>
      write_out);
   ix3917 : oai22 port map ( Y=>nx3916, A0=>nx11971, A1=>nx16157, B0=>
      nx11976, B1=>nx16183);
   modgen_ram_ix74_ix2984 : dff port map ( Q=>OPEN, QB=>nx11971, D=>nx3439, 
      CLK=>nx15529);
   modgen_ram_ix74_ix3092 : dff port map ( Q=>OPEN, QB=>nx11976, D=>nx3429, 
      CLK=>nx15529);
   ix3899 : oai22 port map ( Y=>nx3898, A0=>nx11980, A1=>nx16201, B0=>
      nx11983, B1=>nx18957);
   modgen_ram_ix74_ix3068 : dff port map ( Q=>OPEN, QB=>nx11980, D=>nx3409, 
      CLK=>nx15529);
   modgen_ram_ix74_ix3076 : dff port map ( Q=>OPEN, QB=>nx11983, D=>nx3419, 
      CLK=>nx15531);
   ix11987 : nor02_2x port map ( Y=>nx11986, A0=>nx3878, A1=>nx3860);
   ix3879 : oai33 port map ( Y=>nx3878, A0=>nx11989, A1=>nx15853, A2=>
      nx16093, B0=>nx11992, B1=>nx15423, B2=>nx16023);
   modgen_ram_ix74_ix3176 : dff port map ( Q=>OPEN, QB=>nx11989, D=>nx3389, 
      CLK=>nx15531);
   modgen_ram_ix74_ix2988 : dff port map ( Q=>OPEN, QB=>nx11992, D=>nx3399, 
      CLK=>nx15531);
   ix3861 : oai22 port map ( Y=>nx3860, A0=>nx11996, A1=>nx16259, B0=>
      nx11999, B1=>nx16275);
   modgen_ram_ix74_ix3112 : dff port map ( Q=>OPEN, QB=>nx11996, D=>nx3379, 
      CLK=>nx15531);
   modgen_ram_ix74_ix3048 : dff port map ( Q=>OPEN, QB=>nx11999, D=>nx3369, 
      CLK=>nx15531);
   ix12003 : nor03_2x port map ( Y=>nx12002, A0=>nx3836, A1=>nx3828, A2=>
      nx3820);
   ix3837 : nor03_2x port map ( Y=>nx3836, A0=>nx12005, A1=>nx15767, A2=>
      nx16063);
   modgen_ram_ix74_ix3004 : dff port map ( Q=>OPEN, QB=>nx12005, D=>nx3359, 
      CLK=>nx15531);
   ix3829 : nor03_2x port map ( Y=>nx3828, A0=>nx12009, A1=>nx15855, A2=>
      nx15405);
   modgen_ram_ix74_ix3172 : dff port map ( Q=>OPEN, QB=>nx12009, D=>nx3349, 
      CLK=>nx15531);
   ix3821 : oai33 port map ( Y=>nx3820, A0=>nx12013, A1=>nx15767, A2=>
      nx15913, B0=>nx12016, B1=>nx15423, B2=>nx16063);
   modgen_ram_ix74_ix3012 : dff port map ( Q=>OPEN, QB=>nx12013, D=>nx3329, 
      CLK=>nx15533);
   modgen_ram_ix74_ix2940 : dff port map ( Q=>OPEN, QB=>nx12016, D=>nx3339, 
      CLK=>nx15533);
   ix12020 : nor03_2x port map ( Y=>nx12019, A0=>nx3798, A1=>nx3790, A2=>
      nx3782);
   ix3799 : nor03_2x port map ( Y=>nx3798, A0=>nx12022, A1=>nx15767, A2=>
      nx16041);
   modgen_ram_ix74_ix3008 : dff port map ( Q=>OPEN, QB=>nx12022, D=>nx3319, 
      CLK=>nx15533);
   ix3791 : nor04 port map ( Y=>nx3790, A0=>nx12026, A1=>address(4), A2=>
      address(5), A3=>nx16065);
   modgen_ram_ix74_ix3132 : dff port map ( Q=>OPEN, QB=>nx12026, D=>nx3309, 
      CLK=>nx15533);
   ix3783 : oai22 port map ( Y=>nx3782, A0=>nx12030, A1=>nx16327, B0=>
      nx12033, B1=>nx16343);
   modgen_ram_ix74_ix2948 : dff port map ( Q=>OPEN, QB=>nx12030, D=>nx3289, 
      CLK=>nx15533);
   modgen_ram_ix74_ix2944 : dff port map ( Q=>OPEN, QB=>nx12033, D=>nx3299, 
      CLK=>nx15533);
   modgen_ram_ix74_ix3072 : dff port map ( Q=>OPEN, QB=>nx12040, D=>nx3279, 
      CLK=>nx15533);
   modgen_ram_ix74_ix3136 : dff port map ( Q=>OPEN, QB=>nx12044, D=>nx3269, 
      CLK=>nx15535);
   ix3741 : oai22 port map ( Y=>nx3740, A0=>nx12048, A1=>nx16359, B0=>
      nx12051, B1=>nx16375);
   modgen_ram_ix74_ix3116 : dff port map ( Q=>OPEN, QB=>nx12048, D=>nx3249, 
      CLK=>nx15535);
   modgen_ram_ix74_ix3052 : dff port map ( Q=>OPEN, QB=>nx12051, D=>nx3259, 
      CLK=>nx15535);
   modgen_ram_ix74_ix3180 : dff port map ( Q=>OPEN, QB=>nx12057, D=>nx3239, 
      CLK=>nx15535);
   modgen_ram_ix74_ix2992 : dff port map ( Q=>OPEN, QB=>nx12061, D=>nx3229, 
      CLK=>nx15535);
   ix3703 : oai22 port map ( Y=>nx3702, A0=>nx12065, A1=>nx16399, B0=>
      nx12068, B1=>nx16415);
   modgen_ram_ix74_ix3120 : dff port map ( Q=>OPEN, QB=>nx12065, D=>nx3209, 
      CLK=>nx15535);
   modgen_ram_ix74_ix3056 : dff port map ( Q=>OPEN, QB=>nx12068, D=>nx3219, 
      CLK=>nx15535);
   modgen_ram_ix74_ix3184 : dff port map ( Q=>OPEN, QB=>nx12074, D=>nx3199, 
      CLK=>nx15537);
   modgen_ram_ix74_ix2996 : dff port map ( Q=>OPEN, QB=>nx12078, D=>nx3189, 
      CLK=>nx15537);
   ix3663 : oai22 port map ( Y=>nx3662, A0=>nx12082, A1=>nx16439, B0=>
      nx12085, B1=>nx16455);
   modgen_ram_ix74_ix3124 : dff port map ( Q=>OPEN, QB=>nx12082, D=>nx3169, 
      CLK=>nx15537);
   modgen_ram_ix74_ix3060 : dff port map ( Q=>OPEN, QB=>nx12085, D=>nx3179, 
      CLK=>nx15537);
   modgen_ram_ix74_ix3188 : dff port map ( Q=>OPEN, QB=>nx12091, D=>nx3159, 
      CLK=>nx15537);
   ix3633 : nor03_2x port map ( Y=>nx3632, A0=>nx12095, A1=>nx15425, A2=>
      nx15959);
   modgen_ram_ix74_ix3000 : dff port map ( Q=>OPEN, QB=>nx12095, D=>nx3149, 
      CLK=>nx15537);
   ix3625 : oai22 port map ( Y=>nx3624, A0=>nx12099, A1=>nx16479, B0=>
      nx12102, B1=>nx16495);
   modgen_ram_ix74_ix3128 : dff port map ( Q=>OPEN, QB=>nx12099, D=>nx3129, 
      CLK=>nx15537);
   modgen_ram_ix74_ix3064 : dff port map ( Q=>OPEN, QB=>nx12102, D=>nx3139, 
      CLK=>nx15539);
   ix3599 : oai22 port map ( Y=>nx3598, A0=>nx12112, A1=>nx16511, B0=>
      nx12115, B1=>nx16519);
   modgen_ram_ix74_ix3156 : dff port map ( Q=>OPEN, QB=>nx12112, D=>nx3109, 
      CLK=>nx15539);
   modgen_ram_ix74_ix3192 : dff port map ( Q=>OPEN, QB=>nx12115, D=>nx3119, 
      CLK=>nx15539);
   ix3581 : oai22 port map ( Y=>nx3580, A0=>nx12119, A1=>nx16527, B0=>
      nx12122, B1=>nx16543);
   modgen_ram_ix74_ix3088 : dff port map ( Q=>OPEN, QB=>nx12119, D=>nx3099, 
      CLK=>nx15539);
   modgen_ram_ix74_ix3024 : dff port map ( Q=>OPEN, QB=>nx12122, D=>nx3089, 
      CLK=>nx15539);
   ix3563 : nand03 port map ( Y=>nx3562, A0=>nx12126, A1=>nx12136, A2=>
      nx12142);
   ix12127 : nor02_2x port map ( Y=>nx12126, A0=>nx3558, A1=>nx3550);
   ix3559 : nor04 port map ( Y=>nx3558, A0=>nx12129, A1=>address(4), A2=>
      address(5), A3=>nx15897);
   modgen_ram_ix74_ix3148 : dff port map ( Q=>OPEN, QB=>nx12129, D=>nx3079, 
      CLK=>nx15539);
   ix3551 : nor03_2x port map ( Y=>nx3550, A0=>nx12133, A1=>nx15821, A2=>
      nx15899);
   modgen_ram_ix74_ix3084 : dff port map ( Q=>OPEN, QB=>nx12133, D=>nx3069, 
      CLK=>nx15539);
   ix12137 : nand03 port map ( Y=>nx12136, A0=>modgen_ram_ix74_a_12_dup_946, 
      A1=>nx16231, A2=>nx16569);
   modgen_ram_ix74_ix3144 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_946, 
      QB=>nx12140, D=>nx3059, CLK=>nx15541);
   ix12143 : nand03 port map ( Y=>nx12142, A0=>modgen_ram_ix74_a_28_dup_930, 
      A1=>nx16195, A2=>nx16569);
   modgen_ram_ix74_ix3080 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_930, 
      QB=>nx12146, D=>nx3049, CLK=>nx15541);
   ix12149 : nor03_2x port map ( Y=>nx12148, A0=>nx3518, A1=>nx3510, A2=>
      nx3502);
   ix3519 : nor03_2x port map ( Y=>nx3518, A0=>nx12151, A1=>nx15425, A2=>
      nx15929);
   modgen_ram_ix74_ix2952 : dff port map ( Q=>OPEN, QB=>nx12151, D=>nx3039, 
      CLK=>nx15541);
   ix3511 : nor03_2x port map ( Y=>nx3510, A0=>nx12155, A1=>nx15767, A2=>
      nx15889);
   modgen_ram_ix74_ix3028 : dff port map ( Q=>OPEN, QB=>nx12155, D=>nx3029, 
      CLK=>nx15541);
   ix3503 : oai22 port map ( Y=>nx3502, A0=>nx12159, A1=>nx16603, B0=>
      nx12162, B1=>nx16619);
   modgen_ram_ix74_ix3020 : dff port map ( Q=>OPEN, QB=>nx12159, D=>nx3019, 
      CLK=>nx15541);
   modgen_ram_ix74_ix3016 : dff port map ( Q=>OPEN, QB=>nx12162, D=>nx3009, 
      CLK=>nx15541);
   ix12166 : nor03_2x port map ( Y=>nx12165, A0=>nx3480, A1=>nx3472, A2=>
      nx3464);
   ix3481 : nor03_2x port map ( Y=>nx3480, A0=>nx12168, A1=>nx15855, A2=>
      nx15913);
   modgen_ram_ix74_ix3140 : dff port map ( Q=>OPEN, QB=>nx12168, D=>nx2999, 
      CLK=>nx15541);
   ix3473 : nor03_2x port map ( Y=>nx3472, A0=>nx12172, A1=>nx15425, A2=>
      nx15899);
   modgen_ram_ix74_ix2956 : dff port map ( Q=>OPEN, QB=>nx12172, D=>nx2989, 
      CLK=>nx15543);
   ix3465 : oai22 port map ( Y=>nx3464, A0=>nx12176, A1=>nx16643, B0=>
      nx12179, B1=>nx16659);
   modgen_ram_ix74_ix2964 : dff port map ( Q=>OPEN, QB=>nx12176, D=>nx2979, 
      CLK=>nx15543);
   modgen_ram_ix74_ix2960 : dff port map ( Q=>OPEN, QB=>nx12179, D=>nx2969, 
      CLK=>nx15543);
   ix3441 : oai22 port map ( Y=>nx3440, A0=>nx12186, A1=>nx16675, B0=>
      nx12189, B1=>nx16691);
   modgen_ram_ix74_ix3108 : dff port map ( Q=>OPEN, QB=>nx12186, D=>nx2949, 
      CLK=>nx15543);
   modgen_ram_ix74_ix3152 : dff port map ( Q=>OPEN, QB=>nx12189, D=>nx2959, 
      CLK=>nx15543);
   ix3423 : oai22 port map ( Y=>nx3422, A0=>nx12193, A1=>nx16707, B0=>
      nx12196, B1=>nx16723);
   modgen_ram_ix74_ix3168 : dff port map ( Q=>OPEN, QB=>nx12193, D=>nx2939, 
      CLK=>nx15543);
   modgen_ram_ix74_ix3104 : dff port map ( Q=>OPEN, QB=>nx12196, D=>nx2929, 
      CLK=>nx15543);
   ix12200 : nor03_2x port map ( Y=>nx12199, A0=>nx3400, A1=>nx3392, A2=>
      nx3384);
   ix3401 : nor03_2x port map ( Y=>nx3400, A0=>nx12202, A1=>nx15425, A2=>
      nx15753);
   modgen_ram_ix74_ix2976 : dff port map ( Q=>OPEN, QB=>nx12202, D=>nx2919, 
      CLK=>nx15545);
   ix3393 : nor03_2x port map ( Y=>nx3392, A0=>nx12206, A1=>nx15855, A2=>
      nx15801);
   modgen_ram_ix74_ix3164 : dff port map ( Q=>OPEN, QB=>nx12206, D=>nx2909, 
      CLK=>nx15545);
   ix3385 : oai22 port map ( Y=>nx3384, A0=>nx12210, A1=>nx16747, B0=>
      nx12213, B1=>nx16755);
   modgen_ram_ix74_ix2972 : dff port map ( Q=>OPEN, QB=>nx12210, D=>nx2899, 
      CLK=>nx15545);
   modgen_ram_ix74_ix3160 : dff port map ( Q=>OPEN, QB=>nx12213, D=>nx2889, 
      CLK=>nx15545);
   ix12217 : nor03_2x port map ( Y=>nx12216, A0=>nx3360, A1=>nx3352, A2=>
      nx3344);
   ix3361 : nor03_2x port map ( Y=>nx3360, A0=>nx12219, A1=>nx15767, A2=>
      nx15813);
   modgen_ram_ix74_ix3032 : dff port map ( Q=>OPEN, QB=>nx12219, D=>nx2879, 
      CLK=>nx15545);
   ix3353 : nor03_2x port map ( Y=>nx3352, A0=>nx12223, A1=>nx15823, A2=>
      nx15801);
   modgen_ram_ix74_ix3100 : dff port map ( Q=>OPEN, QB=>nx12223, D=>nx2869, 
      CLK=>nx15545);
   ix3345 : oai22 port map ( Y=>nx3344, A0=>nx12227, A1=>nx16771, B0=>
      nx12230, B1=>nx16787);
   modgen_ram_ix74_ix3096 : dff port map ( Q=>OPEN, QB=>nx12227, D=>nx2859, 
      CLK=>nx15545);
   modgen_ram_ix74_ix2968 : dff port map ( Q=>OPEN, QB=>nx12230, D=>nx2849, 
      CLK=>nx15547);
   ix12234 : nor03_2x port map ( Y=>nx12233, A0=>nx3322, A1=>nx3314, A2=>
      nx3306);
   ix3323 : nor03_2x port map ( Y=>nx3322, A0=>nx12236, A1=>nx15767, A2=>
      nx15801);
   modgen_ram_ix74_ix3036 : dff port map ( Q=>OPEN, QB=>nx12236, D=>nx2839, 
      CLK=>nx15547);
   ix3315 : nor03_2x port map ( Y=>nx3314, A0=>nx12240, A1=>nx15769, A2=>
      nx15405);
   modgen_ram_ix74_ix3044 : dff port map ( Q=>OPEN, QB=>nx12240, D=>nx2829, 
      CLK=>nx15547);
   ix3307 : oai22 port map ( Y=>nx3306, A0=>nx12244, A1=>nx16819, B0=>
      nx12247, B1=>nx16835);
   modgen_ram_ix74_ix2980 : dff port map ( Q=>OPEN, QB=>nx12244, D=>nx2809, 
      CLK=>nx15547);
   modgen_ram_ix74_ix3040 : dff port map ( Q=>OPEN, QB=>nx12247, D=>nx2819, 
      CLK=>nx15547);
   tri_data_out_5 : tri01 port map ( Y=>data_out(5), A=>nx12251, E=>
      write_out);
   ix4555 : oai22 port map ( Y=>nx4554, A0=>nx12257, A1=>nx16157, B0=>
      nx12262, B1=>nx16183);
   modgen_ram_ix74_ix2727 : dff port map ( Q=>OPEN, QB=>nx12257, D=>nx4079, 
      CLK=>nx15547);
   modgen_ram_ix74_ix2835 : dff port map ( Q=>OPEN, QB=>nx12262, D=>nx4069, 
      CLK=>nx15547);
   ix4537 : oai22 port map ( Y=>nx4536, A0=>nx12266, A1=>nx16201, B0=>
      nx12269, B1=>nx18957);
   modgen_ram_ix74_ix2811 : dff port map ( Q=>OPEN, QB=>nx12266, D=>nx4049, 
      CLK=>nx15549);
   modgen_ram_ix74_ix2819 : dff port map ( Q=>OPEN, QB=>nx12269, D=>nx4059, 
      CLK=>nx15549);
   ix12273 : nor02_2x port map ( Y=>nx12272, A0=>nx4516, A1=>nx4498);
   ix4517 : oai33 port map ( Y=>nx4516, A0=>nx12275, A1=>nx15855, A2=>
      nx16093, B0=>nx12278, B1=>nx15425, B2=>nx16023);
   modgen_ram_ix74_ix2919 : dff port map ( Q=>OPEN, QB=>nx12275, D=>nx4029, 
      CLK=>nx15549);
   modgen_ram_ix74_ix2731 : dff port map ( Q=>OPEN, QB=>nx12278, D=>nx4039, 
      CLK=>nx15549);
   ix4499 : oai22 port map ( Y=>nx4498, A0=>nx12282, A1=>nx16259, B0=>
      nx12285, B1=>nx16275);
   modgen_ram_ix74_ix2855 : dff port map ( Q=>OPEN, QB=>nx12282, D=>nx4019, 
      CLK=>nx15549);
   modgen_ram_ix74_ix2791 : dff port map ( Q=>OPEN, QB=>nx12285, D=>nx4009, 
      CLK=>nx15549);
   ix12289 : nor03_2x port map ( Y=>nx12288, A0=>nx4474, A1=>nx4466, A2=>
      nx4458);
   ix4475 : nor03_2x port map ( Y=>nx4474, A0=>nx12291, A1=>nx15769, A2=>
      nx16065);
   modgen_ram_ix74_ix2747 : dff port map ( Q=>OPEN, QB=>nx12291, D=>nx3999, 
      CLK=>nx15549);
   ix4467 : nor03_2x port map ( Y=>nx4466, A0=>nx12295, A1=>nx15855, A2=>
      nx15405);
   modgen_ram_ix74_ix2915 : dff port map ( Q=>OPEN, QB=>nx12295, D=>nx3989, 
      CLK=>nx15551);
   ix4459 : oai33 port map ( Y=>nx4458, A0=>nx12299, A1=>nx15769, A2=>
      nx15913, B0=>nx12302, B1=>nx15427, B2=>nx16065);
   modgen_ram_ix74_ix2755 : dff port map ( Q=>OPEN, QB=>nx12299, D=>nx3969, 
      CLK=>nx15551);
   modgen_ram_ix74_ix2683 : dff port map ( Q=>OPEN, QB=>nx12302, D=>nx3979, 
      CLK=>nx15551);
   ix12306 : nor03_2x port map ( Y=>nx12305, A0=>nx4436, A1=>nx4428, A2=>
      nx4420);
   ix4437 : nor03_2x port map ( Y=>nx4436, A0=>nx12308, A1=>nx15769, A2=>
      nx16043);
   modgen_ram_ix74_ix2751 : dff port map ( Q=>OPEN, QB=>nx12308, D=>nx3959, 
      CLK=>nx15551);
   ix4429 : nor04 port map ( Y=>nx4428, A0=>nx12312, A1=>address(4), A2=>
      address(5), A3=>nx16065);
   modgen_ram_ix74_ix2875 : dff port map ( Q=>OPEN, QB=>nx12312, D=>nx3949, 
      CLK=>nx15551);
   ix4421 : oai22 port map ( Y=>nx4420, A0=>nx12316, A1=>nx16327, B0=>
      nx12319, B1=>nx16343);
   modgen_ram_ix74_ix2691 : dff port map ( Q=>OPEN, QB=>nx12316, D=>nx3929, 
      CLK=>nx15551);
   modgen_ram_ix74_ix2687 : dff port map ( Q=>OPEN, QB=>nx12319, D=>nx3939, 
      CLK=>nx15551);
   modgen_ram_ix74_ix2815 : dff port map ( Q=>OPEN, QB=>nx12326, D=>nx3919, 
      CLK=>nx15553);
   modgen_ram_ix74_ix2879 : dff port map ( Q=>OPEN, QB=>nx12330, D=>nx3909, 
      CLK=>nx15553);
   ix4379 : oai22 port map ( Y=>nx4378, A0=>nx12334, A1=>nx16359, B0=>
      nx12337, B1=>nx16375);
   modgen_ram_ix74_ix2859 : dff port map ( Q=>OPEN, QB=>nx12334, D=>nx3889, 
      CLK=>nx15553);
   modgen_ram_ix74_ix2795 : dff port map ( Q=>OPEN, QB=>nx12337, D=>nx3899, 
      CLK=>nx15553);
   modgen_ram_ix74_ix2923 : dff port map ( Q=>OPEN, QB=>nx12343, D=>nx3879, 
      CLK=>nx15553);
   modgen_ram_ix74_ix2735 : dff port map ( Q=>OPEN, QB=>nx12347, D=>nx3869, 
      CLK=>nx15553);
   ix4341 : oai22 port map ( Y=>nx4340, A0=>nx12351, A1=>nx16399, B0=>
      nx12354, B1=>nx16415);
   modgen_ram_ix74_ix2863 : dff port map ( Q=>OPEN, QB=>nx12351, D=>nx3849, 
      CLK=>nx15553);
   modgen_ram_ix74_ix2799 : dff port map ( Q=>OPEN, QB=>nx12354, D=>nx3859, 
      CLK=>nx15555);
   modgen_ram_ix74_ix2927 : dff port map ( Q=>OPEN, QB=>nx12360, D=>nx3839, 
      CLK=>nx15555);
   modgen_ram_ix74_ix2739 : dff port map ( Q=>OPEN, QB=>nx12364, D=>nx3829, 
      CLK=>nx15555);
   ix4301 : oai22 port map ( Y=>nx4300, A0=>nx12368, A1=>nx16439, B0=>
      nx12371, B1=>nx16455);
   modgen_ram_ix74_ix2867 : dff port map ( Q=>OPEN, QB=>nx12368, D=>nx3809, 
      CLK=>nx15555);
   modgen_ram_ix74_ix2803 : dff port map ( Q=>OPEN, QB=>nx12371, D=>nx3819, 
      CLK=>nx15555);
   modgen_ram_ix74_ix2931 : dff port map ( Q=>OPEN, QB=>nx12377, D=>nx3799, 
      CLK=>nx15555);
   ix4271 : nor03_2x port map ( Y=>nx4270, A0=>nx12381, A1=>nx15427, A2=>
      nx15961);
   modgen_ram_ix74_ix2743 : dff port map ( Q=>OPEN, QB=>nx12381, D=>nx3789, 
      CLK=>nx15555);
   ix4263 : oai22 port map ( Y=>nx4262, A0=>nx12385, A1=>nx16479, B0=>
      nx12388, B1=>nx16495);
   modgen_ram_ix74_ix2871 : dff port map ( Q=>OPEN, QB=>nx12385, D=>nx3769, 
      CLK=>nx15557);
   modgen_ram_ix74_ix2807 : dff port map ( Q=>OPEN, QB=>nx12388, D=>nx3779, 
      CLK=>nx15557);
   ix4237 : oai22 port map ( Y=>nx4236, A0=>nx12398, A1=>nx16511, B0=>
      nx12401, B1=>nx16519);
   modgen_ram_ix74_ix2899 : dff port map ( Q=>OPEN, QB=>nx12398, D=>nx3749, 
      CLK=>nx15557);
   modgen_ram_ix74_ix2935 : dff port map ( Q=>OPEN, QB=>nx12401, D=>nx3759, 
      CLK=>nx15557);
   ix4219 : oai22 port map ( Y=>nx4218, A0=>nx12405, A1=>nx16527, B0=>
      nx12408, B1=>nx16543);
   modgen_ram_ix74_ix2831 : dff port map ( Q=>OPEN, QB=>nx12405, D=>nx3739, 
      CLK=>nx15557);
   modgen_ram_ix74_ix2767 : dff port map ( Q=>OPEN, QB=>nx12408, D=>nx3729, 
      CLK=>nx15557);
   ix4201 : nand03 port map ( Y=>nx4200, A0=>nx12412, A1=>nx12422, A2=>
      nx12428);
   ix12413 : nor02_2x port map ( Y=>nx12412, A0=>nx4196, A1=>nx4188);
   ix4197 : nor04 port map ( Y=>nx4196, A0=>nx12415, A1=>address(4), A2=>
      address(5), A3=>nx15899);
   modgen_ram_ix74_ix2891 : dff port map ( Q=>OPEN, QB=>nx12415, D=>nx3719, 
      CLK=>nx15557);
   ix4189 : nor03_2x port map ( Y=>nx4188, A0=>nx12419, A1=>nx15823, A2=>
      nx15899);
   modgen_ram_ix74_ix2827 : dff port map ( Q=>OPEN, QB=>nx12419, D=>nx3709, 
      CLK=>nx15559);
   ix12423 : nand03 port map ( Y=>nx12422, A0=>modgen_ram_ix74_a_12_dup_881, 
      A1=>nx16231, A2=>nx16569);
   modgen_ram_ix74_ix2887 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_881, 
      QB=>nx12426, D=>nx3699, CLK=>nx15559);
   ix12429 : nand03 port map ( Y=>nx12428, A0=>modgen_ram_ix74_a_28_dup_865, 
      A1=>nx16195, A2=>nx16571);
   modgen_ram_ix74_ix2823 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_865, 
      QB=>nx12432, D=>nx3689, CLK=>nx15559);
   ix12435 : nor03_2x port map ( Y=>nx12434, A0=>nx4156, A1=>nx4148, A2=>
      nx4140);
   ix4157 : nor03_2x port map ( Y=>nx4156, A0=>nx12437, A1=>nx15427, A2=>
      nx15929);
   modgen_ram_ix74_ix2695 : dff port map ( Q=>OPEN, QB=>nx12437, D=>nx3679, 
      CLK=>nx15559);
   ix4149 : nor03_2x port map ( Y=>nx4148, A0=>nx12441, A1=>nx15769, A2=>
      nx15889);
   modgen_ram_ix74_ix2771 : dff port map ( Q=>OPEN, QB=>nx12441, D=>nx3669, 
      CLK=>nx15559);
   ix4141 : oai22 port map ( Y=>nx4140, A0=>nx12445, A1=>nx16603, B0=>
      nx12448, B1=>nx16619);
   modgen_ram_ix74_ix2763 : dff port map ( Q=>OPEN, QB=>nx12445, D=>nx3659, 
      CLK=>nx15559);
   modgen_ram_ix74_ix2759 : dff port map ( Q=>OPEN, QB=>nx12448, D=>nx3649, 
      CLK=>nx15559);
   ix12452 : nor03_2x port map ( Y=>nx12451, A0=>nx4118, A1=>nx4110, A2=>
      nx4102);
   ix4119 : nor03_2x port map ( Y=>nx4118, A0=>nx12454, A1=>nx15857, A2=>
      nx15913);
   modgen_ram_ix74_ix2883 : dff port map ( Q=>OPEN, QB=>nx12454, D=>nx3639, 
      CLK=>nx15561);
   ix4111 : nor03_2x port map ( Y=>nx4110, A0=>nx12458, A1=>nx15427, A2=>
      nx15899);
   modgen_ram_ix74_ix2699 : dff port map ( Q=>OPEN, QB=>nx12458, D=>nx3629, 
      CLK=>nx15561);
   ix4103 : oai22 port map ( Y=>nx4102, A0=>nx12462, A1=>nx16643, B0=>
      nx12465, B1=>nx16659);
   modgen_ram_ix74_ix2707 : dff port map ( Q=>OPEN, QB=>nx12462, D=>nx3619, 
      CLK=>nx15561);
   modgen_ram_ix74_ix2703 : dff port map ( Q=>OPEN, QB=>nx12465, D=>nx3609, 
      CLK=>nx15561);
   ix4079 : oai22 port map ( Y=>nx4078, A0=>nx12472, A1=>nx16675, B0=>
      nx12475, B1=>nx16691);
   modgen_ram_ix74_ix2851 : dff port map ( Q=>OPEN, QB=>nx12472, D=>nx3589, 
      CLK=>nx15561);
   modgen_ram_ix74_ix2895 : dff port map ( Q=>OPEN, QB=>nx12475, D=>nx3599, 
      CLK=>nx15561);
   ix4061 : oai22 port map ( Y=>nx4060, A0=>nx12479, A1=>nx16707, B0=>
      nx12482, B1=>nx16723);
   modgen_ram_ix74_ix2911 : dff port map ( Q=>OPEN, QB=>nx12479, D=>nx3579, 
      CLK=>nx15561);
   modgen_ram_ix74_ix2847 : dff port map ( Q=>OPEN, QB=>nx12482, D=>nx3569, 
      CLK=>nx15563);
   ix12486 : nor03_2x port map ( Y=>nx12485, A0=>nx4038, A1=>nx4030, A2=>
      nx4022);
   ix4039 : nor03_2x port map ( Y=>nx4038, A0=>nx12488, A1=>nx15427, A2=>
      nx15753);
   modgen_ram_ix74_ix2719 : dff port map ( Q=>OPEN, QB=>nx12488, D=>nx3559, 
      CLK=>nx15563);
   ix4031 : nor03_2x port map ( Y=>nx4030, A0=>nx12492, A1=>nx15857, A2=>
      nx15801);
   modgen_ram_ix74_ix2907 : dff port map ( Q=>OPEN, QB=>nx12492, D=>nx3549, 
      CLK=>nx15563);
   ix4023 : oai22 port map ( Y=>nx4022, A0=>nx12496, A1=>nx16747, B0=>
      nx12499, B1=>nx16755);
   modgen_ram_ix74_ix2715 : dff port map ( Q=>OPEN, QB=>nx12496, D=>nx3539, 
      CLK=>nx15563);
   modgen_ram_ix74_ix2903 : dff port map ( Q=>OPEN, QB=>nx12499, D=>nx3529, 
      CLK=>nx15563);
   ix12503 : nor03_2x port map ( Y=>nx12502, A0=>nx3998, A1=>nx3990, A2=>
      nx3982);
   ix3999 : nor03_2x port map ( Y=>nx3998, A0=>nx12505, A1=>nx15769, A2=>
      nx15815);
   modgen_ram_ix74_ix2775 : dff port map ( Q=>OPEN, QB=>nx12505, D=>nx3519, 
      CLK=>nx15563);
   ix3991 : nor03_2x port map ( Y=>nx3990, A0=>nx12509, A1=>nx15823, A2=>
      nx15801);
   modgen_ram_ix74_ix2843 : dff port map ( Q=>OPEN, QB=>nx12509, D=>nx3509, 
      CLK=>nx15563);
   ix3983 : oai22 port map ( Y=>nx3982, A0=>nx12513, A1=>nx16771, B0=>
      nx12516, B1=>nx16787);
   modgen_ram_ix74_ix2839 : dff port map ( Q=>OPEN, QB=>nx12513, D=>nx3499, 
      CLK=>nx15565);
   modgen_ram_ix74_ix2711 : dff port map ( Q=>OPEN, QB=>nx12516, D=>nx3489, 
      CLK=>nx15565);
   ix12520 : nor03_2x port map ( Y=>nx12519, A0=>nx3960, A1=>nx3952, A2=>
      nx3944);
   ix3961 : nor03_2x port map ( Y=>nx3960, A0=>nx12522, A1=>nx15769, A2=>
      nx15801);
   modgen_ram_ix74_ix2779 : dff port map ( Q=>OPEN, QB=>nx12522, D=>nx3479, 
      CLK=>nx15565);
   ix3953 : nor03_2x port map ( Y=>nx3952, A0=>nx12526, A1=>nx15771, A2=>
      nx15405);
   modgen_ram_ix74_ix2787 : dff port map ( Q=>OPEN, QB=>nx12526, D=>nx3469, 
      CLK=>nx15565);
   ix3945 : oai22 port map ( Y=>nx3944, A0=>nx12530, A1=>nx16819, B0=>
      nx12533, B1=>nx16835);
   modgen_ram_ix74_ix2723 : dff port map ( Q=>OPEN, QB=>nx12530, D=>nx3449, 
      CLK=>nx15565);
   modgen_ram_ix74_ix2783 : dff port map ( Q=>OPEN, QB=>nx12533, D=>nx3459, 
      CLK=>nx15565);
   tri_data_out_6 : tri01 port map ( Y=>data_out(6), A=>nx12537, E=>
      write_out);
   ix5193 : oai22 port map ( Y=>nx5192, A0=>nx12543, A1=>nx16157, B0=>
      nx12548, B1=>nx16183);
   modgen_ram_ix74_ix2470 : dff port map ( Q=>OPEN, QB=>nx12543, D=>nx4719, 
      CLK=>nx15565);
   modgen_ram_ix74_ix2578 : dff port map ( Q=>OPEN, QB=>nx12548, D=>nx4709, 
      CLK=>nx15567);
   ix5175 : oai22 port map ( Y=>nx5174, A0=>nx12552, A1=>nx16201, B0=>
      nx12555, B1=>nx18957);
   modgen_ram_ix74_ix2554 : dff port map ( Q=>OPEN, QB=>nx12552, D=>nx4689, 
      CLK=>nx15567);
   modgen_ram_ix74_ix2562 : dff port map ( Q=>OPEN, QB=>nx12555, D=>nx4699, 
      CLK=>nx15567);
   ix12559 : nor02_2x port map ( Y=>nx12558, A0=>nx5154, A1=>nx5136);
   ix5155 : oai33 port map ( Y=>nx5154, A0=>nx12561, A1=>nx15857, A2=>
      nx16093, B0=>nx12564, B1=>nx15429, B2=>nx16023);
   modgen_ram_ix74_ix2662 : dff port map ( Q=>OPEN, QB=>nx12561, D=>nx4669, 
      CLK=>nx15567);
   modgen_ram_ix74_ix2474 : dff port map ( Q=>OPEN, QB=>nx12564, D=>nx4679, 
      CLK=>nx15567);
   ix5137 : oai22 port map ( Y=>nx5136, A0=>nx12568, A1=>nx16259, B0=>
      nx12571, B1=>nx16275);
   modgen_ram_ix74_ix2598 : dff port map ( Q=>OPEN, QB=>nx12568, D=>nx4659, 
      CLK=>nx15567);
   modgen_ram_ix74_ix2534 : dff port map ( Q=>OPEN, QB=>nx12571, D=>nx4649, 
      CLK=>nx15567);
   ix12575 : nor03_2x port map ( Y=>nx12574, A0=>nx5112, A1=>nx5104, A2=>
      nx5096);
   ix5113 : nor03_2x port map ( Y=>nx5112, A0=>nx12577, A1=>nx15771, A2=>
      nx16065);
   modgen_ram_ix74_ix2490 : dff port map ( Q=>OPEN, QB=>nx12577, D=>nx4639, 
      CLK=>nx15569);
   ix5105 : nor03_2x port map ( Y=>nx5104, A0=>nx12581, A1=>nx15857, A2=>
      nx15407);
   modgen_ram_ix74_ix2658 : dff port map ( Q=>OPEN, QB=>nx12581, D=>nx4629, 
      CLK=>nx15569);
   ix5097 : oai33 port map ( Y=>nx5096, A0=>nx12585, A1=>nx15771, A2=>
      nx15915, B0=>nx12588, B1=>nx15429, B2=>nx16065);
   modgen_ram_ix74_ix2498 : dff port map ( Q=>OPEN, QB=>nx12585, D=>nx4609, 
      CLK=>nx15569);
   modgen_ram_ix74_ix2426 : dff port map ( Q=>OPEN, QB=>nx12588, D=>nx4619, 
      CLK=>nx15569);
   ix12592 : nor03_2x port map ( Y=>nx12591, A0=>nx5074, A1=>nx5066, A2=>
      nx5058);
   ix5075 : nor03_2x port map ( Y=>nx5074, A0=>nx12594, A1=>nx15771, A2=>
      nx16043);
   modgen_ram_ix74_ix2494 : dff port map ( Q=>OPEN, QB=>nx12594, D=>nx4599, 
      CLK=>nx15569);
   ix5067 : nor04 port map ( Y=>nx5066, A0=>nx12598, A1=>address(4), A2=>
      address(5), A3=>nx16065);
   modgen_ram_ix74_ix2618 : dff port map ( Q=>OPEN, QB=>nx12598, D=>nx4589, 
      CLK=>nx15569);
   ix5059 : oai22 port map ( Y=>nx5058, A0=>nx12602, A1=>nx16327, B0=>
      nx12605, B1=>nx16343);
   modgen_ram_ix74_ix2434 : dff port map ( Q=>OPEN, QB=>nx12602, D=>nx4569, 
      CLK=>nx15569);
   modgen_ram_ix74_ix2430 : dff port map ( Q=>OPEN, QB=>nx12605, D=>nx4579, 
      CLK=>nx15571);
   modgen_ram_ix74_ix2558 : dff port map ( Q=>OPEN, QB=>nx12612, D=>nx4559, 
      CLK=>nx15571);
   modgen_ram_ix74_ix2622 : dff port map ( Q=>OPEN, QB=>nx12616, D=>nx4549, 
      CLK=>nx15571);
   ix5017 : oai22 port map ( Y=>nx5016, A0=>nx12620, A1=>nx16359, B0=>
      nx12623, B1=>nx16375);
   modgen_ram_ix74_ix2602 : dff port map ( Q=>OPEN, QB=>nx12620, D=>nx4529, 
      CLK=>nx15571);
   modgen_ram_ix74_ix2538 : dff port map ( Q=>OPEN, QB=>nx12623, D=>nx4539, 
      CLK=>nx15571);
   modgen_ram_ix74_ix2666 : dff port map ( Q=>OPEN, QB=>nx12629, D=>nx4519, 
      CLK=>nx15571);
   modgen_ram_ix74_ix2478 : dff port map ( Q=>OPEN, QB=>nx12633, D=>nx4509, 
      CLK=>nx15571);
   ix4979 : oai22 port map ( Y=>nx4978, A0=>nx12637, A1=>nx16399, B0=>
      nx12640, B1=>nx16415);
   modgen_ram_ix74_ix2606 : dff port map ( Q=>OPEN, QB=>nx12637, D=>nx4489, 
      CLK=>nx15573);
   modgen_ram_ix74_ix2542 : dff port map ( Q=>OPEN, QB=>nx12640, D=>nx4499, 
      CLK=>nx15573);
   modgen_ram_ix74_ix2670 : dff port map ( Q=>OPEN, QB=>nx12646, D=>nx4479, 
      CLK=>nx15573);
   modgen_ram_ix74_ix2482 : dff port map ( Q=>OPEN, QB=>nx12650, D=>nx4469, 
      CLK=>nx15573);
   ix4939 : oai22 port map ( Y=>nx4938, A0=>nx12654, A1=>nx16439, B0=>
      nx12657, B1=>nx16455);
   modgen_ram_ix74_ix2610 : dff port map ( Q=>OPEN, QB=>nx12654, D=>nx4449, 
      CLK=>nx15573);
   modgen_ram_ix74_ix2546 : dff port map ( Q=>OPEN, QB=>nx12657, D=>nx4459, 
      CLK=>nx15573);
   modgen_ram_ix74_ix2674 : dff port map ( Q=>OPEN, QB=>nx12663, D=>nx4439, 
      CLK=>nx15573);
   ix4909 : nor03_2x port map ( Y=>nx4908, A0=>nx12667, A1=>nx15429, A2=>
      nx15961);
   modgen_ram_ix74_ix2486 : dff port map ( Q=>OPEN, QB=>nx12667, D=>nx4429, 
      CLK=>nx15575);
   ix4901 : oai22 port map ( Y=>nx4900, A0=>nx12671, A1=>nx16479, B0=>
      nx12674, B1=>nx16495);
   modgen_ram_ix74_ix2614 : dff port map ( Q=>OPEN, QB=>nx12671, D=>nx4409, 
      CLK=>nx15575);
   modgen_ram_ix74_ix2550 : dff port map ( Q=>OPEN, QB=>nx12674, D=>nx4419, 
      CLK=>nx15575);
   ix4875 : oai22 port map ( Y=>nx4874, A0=>nx12684, A1=>nx16511, B0=>
      nx12687, B1=>nx16519);
   modgen_ram_ix74_ix2642 : dff port map ( Q=>OPEN, QB=>nx12684, D=>nx4389, 
      CLK=>nx15575);
   modgen_ram_ix74_ix2678 : dff port map ( Q=>OPEN, QB=>nx12687, D=>nx4399, 
      CLK=>nx15575);
   ix4857 : oai22 port map ( Y=>nx4856, A0=>nx12691, A1=>nx16527, B0=>
      nx12694, B1=>nx16543);
   modgen_ram_ix74_ix2574 : dff port map ( Q=>OPEN, QB=>nx12691, D=>nx4379, 
      CLK=>nx15575);
   modgen_ram_ix74_ix2510 : dff port map ( Q=>OPEN, QB=>nx12694, D=>nx4369, 
      CLK=>nx15575);
   ix4839 : nand03 port map ( Y=>nx4838, A0=>nx12698, A1=>nx12708, A2=>
      nx12714);
   ix12699 : nor02_2x port map ( Y=>nx12698, A0=>nx4834, A1=>nx4826);
   ix4835 : nor04 port map ( Y=>nx4834, A0=>nx12701, A1=>address(4), A2=>
      address(5), A3=>nx15899);
   modgen_ram_ix74_ix2634 : dff port map ( Q=>OPEN, QB=>nx12701, D=>nx4359, 
      CLK=>nx15577);
   ix4827 : nor03_2x port map ( Y=>nx4826, A0=>nx12705, A1=>nx15823, A2=>
      nx15899);
   modgen_ram_ix74_ix2570 : dff port map ( Q=>OPEN, QB=>nx12705, D=>nx4349, 
      CLK=>nx15577);
   ix12709 : nand03 port map ( Y=>nx12708, A0=>modgen_ram_ix74_a_12_dup_815, 
      A1=>nx16231, A2=>nx16571);
   modgen_ram_ix74_ix2630 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_815, 
      QB=>nx12712, D=>nx4339, CLK=>nx15577);
   ix12715 : nand03 port map ( Y=>nx12714, A0=>modgen_ram_ix74_a_28_dup_799, 
      A1=>nx16197, A2=>nx16571);
   modgen_ram_ix74_ix2566 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_799, 
      QB=>nx12718, D=>nx4329, CLK=>nx15577);
   ix12721 : nor03_2x port map ( Y=>nx12720, A0=>nx4794, A1=>nx4786, A2=>
      nx4778);
   ix4795 : nor03_2x port map ( Y=>nx4794, A0=>nx12723, A1=>nx15429, A2=>
      nx15931);
   modgen_ram_ix74_ix2438 : dff port map ( Q=>OPEN, QB=>nx12723, D=>nx4319, 
      CLK=>nx15577);
   ix4787 : nor03_2x port map ( Y=>nx4786, A0=>nx12727, A1=>nx15771, A2=>
      nx15891);
   modgen_ram_ix74_ix2514 : dff port map ( Q=>OPEN, QB=>nx12727, D=>nx4309, 
      CLK=>nx15577);
   ix4779 : oai22 port map ( Y=>nx4778, A0=>nx12731, A1=>nx16603, B0=>
      nx12734, B1=>nx16619);
   modgen_ram_ix74_ix2506 : dff port map ( Q=>OPEN, QB=>nx12731, D=>nx4299, 
      CLK=>nx15577);
   modgen_ram_ix74_ix2502 : dff port map ( Q=>OPEN, QB=>nx12734, D=>nx4289, 
      CLK=>nx15579);
   ix4757 : nor03_2x port map ( Y=>nx4756, A0=>nx12740, A1=>nx15857, A2=>
      nx15915);
   modgen_ram_ix74_ix2626 : dff port map ( Q=>OPEN, QB=>nx12740, D=>nx4279, 
      CLK=>nx15579);
   ix4749 : nor03_2x port map ( Y=>nx4748, A0=>nx12744, A1=>nx15429, A2=>
      nx15901);
   modgen_ram_ix74_ix2442 : dff port map ( Q=>OPEN, QB=>nx12744, D=>nx4269, 
      CLK=>nx15579);
   modgen_ram_ix74_ix2450 : dff port map ( Q=>OPEN, QB=>nx12748, D=>nx4259, 
      CLK=>nx15579);
   modgen_ram_ix74_ix2446 : dff port map ( Q=>OPEN, QB=>nx12751, D=>nx4249, 
      CLK=>nx15579);
   ix4717 : oai22 port map ( Y=>nx4716, A0=>nx12758, A1=>nx16675, B0=>
      nx12761, B1=>nx16691);
   modgen_ram_ix74_ix2594 : dff port map ( Q=>OPEN, QB=>nx12758, D=>nx4229, 
      CLK=>nx15579);
   modgen_ram_ix74_ix2638 : dff port map ( Q=>OPEN, QB=>nx12761, D=>nx4239, 
      CLK=>nx15579);
   ix4699 : oai22 port map ( Y=>nx4698, A0=>nx12765, A1=>nx16707, B0=>
      nx12768, B1=>nx16723);
   modgen_ram_ix74_ix2654 : dff port map ( Q=>OPEN, QB=>nx12765, D=>nx4219, 
      CLK=>nx15581);
   modgen_ram_ix74_ix2590 : dff port map ( Q=>OPEN, QB=>nx12768, D=>nx4209, 
      CLK=>nx15581);
   ix12772 : nor03_2x port map ( Y=>nx12771, A0=>nx4676, A1=>nx4668, A2=>
      nx4660);
   ix4677 : nor03_2x port map ( Y=>nx4676, A0=>nx12774, A1=>nx15431, A2=>
      nx15755);
   modgen_ram_ix74_ix2462 : dff port map ( Q=>OPEN, QB=>nx12774, D=>nx4199, 
      CLK=>nx15581);
   ix4669 : nor03_2x port map ( Y=>nx4668, A0=>nx12778, A1=>nx15857, A2=>
      nx15801);
   modgen_ram_ix74_ix2650 : dff port map ( Q=>OPEN, QB=>nx12778, D=>nx4189, 
      CLK=>nx15581);
   ix4661 : oai22 port map ( Y=>nx4660, A0=>nx12782, A1=>nx16747, B0=>
      nx12785, B1=>nx16755);
   modgen_ram_ix74_ix2458 : dff port map ( Q=>OPEN, QB=>nx12782, D=>nx4179, 
      CLK=>nx15581);
   modgen_ram_ix74_ix2646 : dff port map ( Q=>OPEN, QB=>nx12785, D=>nx4169, 
      CLK=>nx15581);
   ix12789 : nor03_2x port map ( Y=>nx12788, A0=>nx4636, A1=>nx4628, A2=>
      nx4620);
   ix4637 : nor03_2x port map ( Y=>nx4636, A0=>nx12791, A1=>nx15771, A2=>
      nx15815);
   modgen_ram_ix74_ix2518 : dff port map ( Q=>OPEN, QB=>nx12791, D=>nx4159, 
      CLK=>nx15581);
   ix4629 : nor03_2x port map ( Y=>nx4628, A0=>nx12795, A1=>nx15823, A2=>
      nx15803);
   modgen_ram_ix74_ix2586 : dff port map ( Q=>OPEN, QB=>nx12795, D=>nx4149, 
      CLK=>nx15583);
   ix4621 : oai22 port map ( Y=>nx4620, A0=>nx12799, A1=>nx16771, B0=>
      nx12802, B1=>nx16787);
   modgen_ram_ix74_ix2582 : dff port map ( Q=>OPEN, QB=>nx12799, D=>nx4139, 
      CLK=>nx15583);
   modgen_ram_ix74_ix2454 : dff port map ( Q=>OPEN, QB=>nx12802, D=>nx4129, 
      CLK=>nx15583);
   ix12806 : nor03_2x port map ( Y=>nx12805, A0=>nx4598, A1=>nx4590, A2=>
      nx4582);
   ix4599 : nor03_2x port map ( Y=>nx4598, A0=>nx12808, A1=>nx15771, A2=>
      nx15803);
   modgen_ram_ix74_ix2522 : dff port map ( Q=>OPEN, QB=>nx12808, D=>nx4119, 
      CLK=>nx15583);
   ix4591 : nor03_2x port map ( Y=>nx4590, A0=>nx12812, A1=>nx15773, A2=>
      nx15407);
   modgen_ram_ix74_ix2530 : dff port map ( Q=>OPEN, QB=>nx12812, D=>nx4109, 
      CLK=>nx15583);
   ix4583 : oai22 port map ( Y=>nx4582, A0=>nx12816, A1=>nx16819, B0=>
      nx12819, B1=>nx16835);
   modgen_ram_ix74_ix2466 : dff port map ( Q=>OPEN, QB=>nx12816, D=>nx4089, 
      CLK=>nx15583);
   modgen_ram_ix74_ix2526 : dff port map ( Q=>OPEN, QB=>nx12819, D=>nx4099, 
      CLK=>nx15583);
   tri_data_out_7 : tri01 port map ( Y=>data_out(7), A=>nx12823, E=>
      write_out);
   ix5831 : oai22 port map ( Y=>nx5830, A0=>nx12829, A1=>nx16159, B0=>
      nx12834, B1=>nx16185);
   modgen_ram_ix74_ix2213 : dff port map ( Q=>OPEN, QB=>nx12829, D=>nx5359, 
      CLK=>nx15585);
   modgen_ram_ix74_ix2321 : dff port map ( Q=>OPEN, QB=>nx12834, D=>nx5349, 
      CLK=>nx15585);
   ix5813 : oai22 port map ( Y=>nx5812, A0=>nx12838, A1=>nx16203, B0=>
      nx12841, B1=>nx18957);
   modgen_ram_ix74_ix2297 : dff port map ( Q=>OPEN, QB=>nx12838, D=>nx5329, 
      CLK=>nx15585);
   modgen_ram_ix74_ix2305 : dff port map ( Q=>OPEN, QB=>nx12841, D=>nx5339, 
      CLK=>nx15585);
   ix12845 : nor02_2x port map ( Y=>nx12844, A0=>nx5792, A1=>nx5774);
   ix5793 : oai33 port map ( Y=>nx5792, A0=>nx12847, A1=>nx15859, A2=>
      nx16095, B0=>nx12850, B1=>nx15431, B2=>nx16025);
   modgen_ram_ix74_ix2405 : dff port map ( Q=>OPEN, QB=>nx12847, D=>nx5309, 
      CLK=>nx15585);
   modgen_ram_ix74_ix2217 : dff port map ( Q=>OPEN, QB=>nx12850, D=>nx5319, 
      CLK=>nx15585);
   ix5775 : oai22 port map ( Y=>nx5774, A0=>nx12854, A1=>nx16261, B0=>
      nx12857, B1=>nx16277);
   modgen_ram_ix74_ix2341 : dff port map ( Q=>OPEN, QB=>nx12854, D=>nx5299, 
      CLK=>nx15585);
   modgen_ram_ix74_ix2277 : dff port map ( Q=>OPEN, QB=>nx12857, D=>nx5289, 
      CLK=>nx15587);
   ix12861 : nor03_2x port map ( Y=>nx12860, A0=>nx5750, A1=>nx5742, A2=>
      nx5734);
   ix5751 : nor03_2x port map ( Y=>nx5750, A0=>nx12863, A1=>nx15773, A2=>
      nx16067);
   modgen_ram_ix74_ix2233 : dff port map ( Q=>OPEN, QB=>nx12863, D=>nx5279, 
      CLK=>nx15587);
   ix5743 : nor03_2x port map ( Y=>nx5742, A0=>nx12867, A1=>nx15859, A2=>
      nx15407);
   modgen_ram_ix74_ix2401 : dff port map ( Q=>OPEN, QB=>nx12867, D=>nx5269, 
      CLK=>nx15587);
   ix5735 : oai33 port map ( Y=>nx5734, A0=>nx12871, A1=>nx15773, A2=>
      nx15915, B0=>nx12874, B1=>nx15431, B2=>nx16067);
   modgen_ram_ix74_ix2241 : dff port map ( Q=>OPEN, QB=>nx12871, D=>nx5249, 
      CLK=>nx15587);
   modgen_ram_ix74_ix2169 : dff port map ( Q=>OPEN, QB=>nx12874, D=>nx5259, 
      CLK=>nx15587);
   ix12878 : nor03_2x port map ( Y=>nx12877, A0=>nx5712, A1=>nx5704, A2=>
      nx5696);
   ix5713 : nor03_2x port map ( Y=>nx5712, A0=>nx12880, A1=>nx15773, A2=>
      nx16045);
   modgen_ram_ix74_ix2237 : dff port map ( Q=>OPEN, QB=>nx12880, D=>nx5239, 
      CLK=>nx15587);
   ix5705 : nor04 port map ( Y=>nx5704, A0=>nx12884, A1=>address(4), A2=>
      address(5), A3=>nx16067);
   modgen_ram_ix74_ix2361 : dff port map ( Q=>OPEN, QB=>nx12884, D=>nx5229, 
      CLK=>nx15587);
   ix5697 : oai22 port map ( Y=>nx5696, A0=>nx12888, A1=>nx16329, B0=>
      nx12891, B1=>nx16345);
   modgen_ram_ix74_ix2177 : dff port map ( Q=>OPEN, QB=>nx12888, D=>nx5209, 
      CLK=>nx15589);
   modgen_ram_ix74_ix2173 : dff port map ( Q=>OPEN, QB=>nx12891, D=>nx5219, 
      CLK=>nx15589);
   modgen_ram_ix74_ix2301 : dff port map ( Q=>OPEN, QB=>nx12898, D=>nx5199, 
      CLK=>nx15589);
   modgen_ram_ix74_ix2365 : dff port map ( Q=>OPEN, QB=>nx12902, D=>nx5189, 
      CLK=>nx15589);
   ix5655 : oai22 port map ( Y=>nx5654, A0=>nx12906, A1=>nx16361, B0=>
      nx12909, B1=>nx16377);
   modgen_ram_ix74_ix2345 : dff port map ( Q=>OPEN, QB=>nx12906, D=>nx5169, 
      CLK=>nx15589);
   modgen_ram_ix74_ix2281 : dff port map ( Q=>OPEN, QB=>nx12909, D=>nx5179, 
      CLK=>nx15589);
   modgen_ram_ix74_ix2409 : dff port map ( Q=>OPEN, QB=>nx12915, D=>nx5159, 
      CLK=>nx15589);
   modgen_ram_ix74_ix2221 : dff port map ( Q=>OPEN, QB=>nx12919, D=>nx5149, 
      CLK=>nx15591);
   ix5617 : oai22 port map ( Y=>nx5616, A0=>nx12923, A1=>nx16401, B0=>
      nx12926, B1=>nx16417);
   modgen_ram_ix74_ix2349 : dff port map ( Q=>OPEN, QB=>nx12923, D=>nx5129, 
      CLK=>nx15591);
   modgen_ram_ix74_ix2285 : dff port map ( Q=>OPEN, QB=>nx12926, D=>nx5139, 
      CLK=>nx15591);
   modgen_ram_ix74_ix2413 : dff port map ( Q=>OPEN, QB=>nx12932, D=>nx5119, 
      CLK=>nx15591);
   modgen_ram_ix74_ix2225 : dff port map ( Q=>OPEN, QB=>nx12936, D=>nx5109, 
      CLK=>nx15591);
   ix5577 : oai22 port map ( Y=>nx5576, A0=>nx12940, A1=>nx16441, B0=>
      nx12943, B1=>nx16457);
   modgen_ram_ix74_ix2353 : dff port map ( Q=>OPEN, QB=>nx12940, D=>nx5089, 
      CLK=>nx15591);
   modgen_ram_ix74_ix2289 : dff port map ( Q=>OPEN, QB=>nx12943, D=>nx5099, 
      CLK=>nx15591);
   modgen_ram_ix74_ix2417 : dff port map ( Q=>OPEN, QB=>nx12949, D=>nx5079, 
      CLK=>nx15593);
   ix5547 : nor03_2x port map ( Y=>nx5546, A0=>nx12953, A1=>nx15431, A2=>
      nx15961);
   modgen_ram_ix74_ix2229 : dff port map ( Q=>OPEN, QB=>nx12953, D=>nx5069, 
      CLK=>nx15593);
   ix5539 : oai22 port map ( Y=>nx5538, A0=>nx12957, A1=>nx16481, B0=>
      nx12960, B1=>nx16497);
   modgen_ram_ix74_ix2357 : dff port map ( Q=>OPEN, QB=>nx12957, D=>nx5049, 
      CLK=>nx15593);
   modgen_ram_ix74_ix2293 : dff port map ( Q=>OPEN, QB=>nx12960, D=>nx5059, 
      CLK=>nx15593);
   ix5513 : oai22 port map ( Y=>nx5512, A0=>nx12970, A1=>nx16513, B0=>
      nx12973, B1=>nx16521);
   modgen_ram_ix74_ix2385 : dff port map ( Q=>OPEN, QB=>nx12970, D=>nx5029, 
      CLK=>nx15593);
   modgen_ram_ix74_ix2421 : dff port map ( Q=>OPEN, QB=>nx12973, D=>nx5039, 
      CLK=>nx15593);
   ix5495 : oai22 port map ( Y=>nx5494, A0=>nx12977, A1=>nx16529, B0=>
      nx12980, B1=>nx16545);
   modgen_ram_ix74_ix2317 : dff port map ( Q=>OPEN, QB=>nx12977, D=>nx5019, 
      CLK=>nx15593);
   modgen_ram_ix74_ix2253 : dff port map ( Q=>OPEN, QB=>nx12980, D=>nx5009, 
      CLK=>nx15595);
   ix5477 : nand03 port map ( Y=>nx5476, A0=>nx12984, A1=>nx12994, A2=>
      nx13000);
   ix12985 : nor02_2x port map ( Y=>nx12984, A0=>nx5472, A1=>nx5464);
   ix5473 : nor04 port map ( Y=>nx5472, A0=>nx12987, A1=>address(4), A2=>
      address(5), A3=>nx15901);
   modgen_ram_ix74_ix2377 : dff port map ( Q=>OPEN, QB=>nx12987, D=>nx4999, 
      CLK=>nx15595);
   ix5465 : nor03_2x port map ( Y=>nx5464, A0=>nx12991, A1=>nx15825, A2=>
      nx15901);
   modgen_ram_ix74_ix2313 : dff port map ( Q=>OPEN, QB=>nx12991, D=>nx4989, 
      CLK=>nx15595);
   ix12995 : nand03 port map ( Y=>nx12994, A0=>modgen_ram_ix74_a_12_dup_750, 
      A1=>nx16231, A2=>nx16571);
   modgen_ram_ix74_ix2373 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_750, 
      QB=>nx12998, D=>nx4979, CLK=>nx15595);
   ix13001 : nand03 port map ( Y=>nx13000, A0=>modgen_ram_ix74_a_28_dup_734, 
      A1=>nx16197, A2=>nx16571);
   modgen_ram_ix74_ix2309 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_734, 
      QB=>nx13004, D=>nx4969, CLK=>nx15595);
   ix13007 : nor03_2x port map ( Y=>nx13006, A0=>nx5432, A1=>nx5424, A2=>
      nx5416);
   ix5433 : nor03_2x port map ( Y=>nx5432, A0=>nx13009, A1=>nx15431, A2=>
      nx15931);
   modgen_ram_ix74_ix2181 : dff port map ( Q=>OPEN, QB=>nx13009, D=>nx4959, 
      CLK=>nx15595);
   ix5425 : nor03_2x port map ( Y=>nx5424, A0=>nx13013, A1=>nx15773, A2=>
      nx15891);
   modgen_ram_ix74_ix2257 : dff port map ( Q=>OPEN, QB=>nx13013, D=>nx4949, 
      CLK=>nx15595);
   ix5417 : oai22 port map ( Y=>nx5416, A0=>nx13017, A1=>nx16605, B0=>
      nx13020, B1=>nx16621);
   modgen_ram_ix74_ix2249 : dff port map ( Q=>OPEN, QB=>nx13017, D=>nx4939, 
      CLK=>nx15597);
   modgen_ram_ix74_ix2245 : dff port map ( Q=>OPEN, QB=>nx13020, D=>nx4929, 
      CLK=>nx15597);
   ix13024 : nor03_2x port map ( Y=>nx13023, A0=>nx5394, A1=>nx5386, A2=>
      nx5378);
   ix5395 : nor03_2x port map ( Y=>nx5394, A0=>nx13026, A1=>nx15859, A2=>
      nx15915);
   modgen_ram_ix74_ix2369 : dff port map ( Q=>OPEN, QB=>nx13026, D=>nx4919, 
      CLK=>nx15597);
   ix5387 : nor03_2x port map ( Y=>nx5386, A0=>nx13030, A1=>nx15433, A2=>
      nx15901);
   modgen_ram_ix74_ix2185 : dff port map ( Q=>OPEN, QB=>nx13030, D=>nx4909, 
      CLK=>nx15597);
   ix5379 : oai22 port map ( Y=>nx5378, A0=>nx13034, A1=>nx16645, B0=>
      nx13037, B1=>nx16661);
   modgen_ram_ix74_ix2193 : dff port map ( Q=>OPEN, QB=>nx13034, D=>nx4899, 
      CLK=>nx15597);
   modgen_ram_ix74_ix2189 : dff port map ( Q=>OPEN, QB=>nx13037, D=>nx4889, 
      CLK=>nx15597);
   ix5355 : oai22 port map ( Y=>nx5354, A0=>nx13044, A1=>nx16677, B0=>
      nx13047, B1=>nx16693);
   modgen_ram_ix74_ix2337 : dff port map ( Q=>OPEN, QB=>nx13044, D=>nx4869, 
      CLK=>nx15597);
   modgen_ram_ix74_ix2381 : dff port map ( Q=>OPEN, QB=>nx13047, D=>nx4879, 
      CLK=>nx15599);
   ix5337 : oai22 port map ( Y=>nx5336, A0=>nx13051, A1=>nx16709, B0=>
      nx13054, B1=>nx16725);
   modgen_ram_ix74_ix2397 : dff port map ( Q=>OPEN, QB=>nx13051, D=>nx4859, 
      CLK=>nx15599);
   modgen_ram_ix74_ix2333 : dff port map ( Q=>OPEN, QB=>nx13054, D=>nx4849, 
      CLK=>nx15599);
   ix13058 : nor03_2x port map ( Y=>nx13057, A0=>nx5314, A1=>nx5306, A2=>
      nx5298);
   ix5315 : nor03_2x port map ( Y=>nx5314, A0=>nx13060, A1=>nx15433, A2=>
      nx15755);
   modgen_ram_ix74_ix2205 : dff port map ( Q=>OPEN, QB=>nx13060, D=>nx4839, 
      CLK=>nx15599);
   ix5307 : nor03_2x port map ( Y=>nx5306, A0=>nx13064, A1=>nx15859, A2=>
      nx15803);
   modgen_ram_ix74_ix2393 : dff port map ( Q=>OPEN, QB=>nx13064, D=>nx4829, 
      CLK=>nx15599);
   ix5299 : oai22 port map ( Y=>nx5298, A0=>nx13068, A1=>nx16749, B0=>
      nx13071, B1=>nx16757);
   modgen_ram_ix74_ix2201 : dff port map ( Q=>OPEN, QB=>nx13068, D=>nx4819, 
      CLK=>nx15599);
   modgen_ram_ix74_ix2389 : dff port map ( Q=>OPEN, QB=>nx13071, D=>nx4809, 
      CLK=>nx15599);
   ix13075 : nor03_2x port map ( Y=>nx13074, A0=>nx5274, A1=>nx5266, A2=>
      nx5258);
   ix5275 : nor03_2x port map ( Y=>nx5274, A0=>nx13077, A1=>nx15773, A2=>
      nx15815);
   modgen_ram_ix74_ix2261 : dff port map ( Q=>OPEN, QB=>nx13077, D=>nx4799, 
      CLK=>nx15601);
   ix5267 : nor03_2x port map ( Y=>nx5266, A0=>nx13081, A1=>nx15825, A2=>
      nx15803);
   modgen_ram_ix74_ix2329 : dff port map ( Q=>OPEN, QB=>nx13081, D=>nx4789, 
      CLK=>nx15601);
   ix5259 : oai22 port map ( Y=>nx5258, A0=>nx13085, A1=>nx16773, B0=>
      nx13088, B1=>nx16789);
   modgen_ram_ix74_ix2325 : dff port map ( Q=>OPEN, QB=>nx13085, D=>nx4779, 
      CLK=>nx15601);
   modgen_ram_ix74_ix2197 : dff port map ( Q=>OPEN, QB=>nx13088, D=>nx4769, 
      CLK=>nx15601);
   ix13092 : nor03_2x port map ( Y=>nx13091, A0=>nx5236, A1=>nx5228, A2=>
      nx5220);
   ix5237 : nor03_2x port map ( Y=>nx5236, A0=>nx13094, A1=>nx15773, A2=>
      nx15803);
   modgen_ram_ix74_ix2265 : dff port map ( Q=>OPEN, QB=>nx13094, D=>nx4759, 
      CLK=>nx15601);
   ix5229 : nor03_2x port map ( Y=>nx5228, A0=>nx13098, A1=>nx15775, A2=>
      nx15407);
   modgen_ram_ix74_ix2273 : dff port map ( Q=>OPEN, QB=>nx13098, D=>nx4749, 
      CLK=>nx15601);
   ix5221 : oai22 port map ( Y=>nx5220, A0=>nx13102, A1=>nx16821, B0=>
      nx13105, B1=>nx16837);
   modgen_ram_ix74_ix2209 : dff port map ( Q=>OPEN, QB=>nx13102, D=>nx4729, 
      CLK=>nx15601);
   modgen_ram_ix74_ix2269 : dff port map ( Q=>OPEN, QB=>nx13105, D=>nx4739, 
      CLK=>nx15603);
   tri_data_out_8 : tri01 port map ( Y=>data_out(8), A=>nx13109, E=>
      write_out);
   ix6469 : oai22 port map ( Y=>nx6468, A0=>nx13115, A1=>nx16159, B0=>
      nx13120, B1=>nx16185);
   modgen_ram_ix74_ix1956 : dff port map ( Q=>OPEN, QB=>nx13115, D=>nx5999, 
      CLK=>nx15603);
   modgen_ram_ix74_ix2064 : dff port map ( Q=>OPEN, QB=>nx13120, D=>nx5989, 
      CLK=>nx15603);
   ix6451 : oai22 port map ( Y=>nx6450, A0=>nx13124, A1=>nx16203, B0=>
      nx13127, B1=>nx18957);
   modgen_ram_ix74_ix2040 : dff port map ( Q=>OPEN, QB=>nx13124, D=>nx5969, 
      CLK=>nx15603);
   modgen_ram_ix74_ix2048 : dff port map ( Q=>OPEN, QB=>nx13127, D=>nx5979, 
      CLK=>nx15603);
   ix13131 : nor02_2x port map ( Y=>nx13130, A0=>nx6430, A1=>nx6412);
   ix6431 : oai33 port map ( Y=>nx6430, A0=>nx13133, A1=>nx15859, A2=>
      nx16095, B0=>nx13136, B1=>nx15433, B2=>nx16025);
   modgen_ram_ix74_ix2148 : dff port map ( Q=>OPEN, QB=>nx13133, D=>nx5949, 
      CLK=>nx15603);
   modgen_ram_ix74_ix1960 : dff port map ( Q=>OPEN, QB=>nx13136, D=>nx5959, 
      CLK=>nx15603);
   ix6413 : oai22 port map ( Y=>nx6412, A0=>nx13140, A1=>nx16261, B0=>
      nx13143, B1=>nx16277);
   modgen_ram_ix74_ix2084 : dff port map ( Q=>OPEN, QB=>nx13140, D=>nx5939, 
      CLK=>nx15605);
   modgen_ram_ix74_ix2020 : dff port map ( Q=>OPEN, QB=>nx13143, D=>nx5929, 
      CLK=>nx15605);
   ix13147 : nor03_2x port map ( Y=>nx13146, A0=>nx6388, A1=>nx6380, A2=>
      nx6372);
   ix6389 : nor03_2x port map ( Y=>nx6388, A0=>nx13149, A1=>nx15775, A2=>
      nx16067);
   modgen_ram_ix74_ix1976 : dff port map ( Q=>OPEN, QB=>nx13149, D=>nx5919, 
      CLK=>nx15605);
   ix6381 : nor03_2x port map ( Y=>nx6380, A0=>nx13153, A1=>nx15859, A2=>
      nx15407);
   modgen_ram_ix74_ix2144 : dff port map ( Q=>OPEN, QB=>nx13153, D=>nx5909, 
      CLK=>nx15605);
   ix6373 : oai33 port map ( Y=>nx6372, A0=>nx13157, A1=>nx15775, A2=>
      nx15915, B0=>nx13160, B1=>nx15433, B2=>nx16067);
   modgen_ram_ix74_ix1984 : dff port map ( Q=>OPEN, QB=>nx13157, D=>nx5889, 
      CLK=>nx15605);
   modgen_ram_ix74_ix1912 : dff port map ( Q=>OPEN, QB=>nx13160, D=>nx5899, 
      CLK=>nx15605);
   ix13164 : nor03_2x port map ( Y=>nx13163, A0=>nx6350, A1=>nx6342, A2=>
      nx6334);
   ix6351 : nor03_2x port map ( Y=>nx6350, A0=>nx13166, A1=>nx15775, A2=>
      nx16045);
   modgen_ram_ix74_ix1980 : dff port map ( Q=>OPEN, QB=>nx13166, D=>nx5879, 
      CLK=>nx15605);
   ix6343 : nor04 port map ( Y=>nx6342, A0=>nx13170, A1=>address(4), A2=>
      address(5), A3=>nx16067);
   modgen_ram_ix74_ix2104 : dff port map ( Q=>OPEN, QB=>nx13170, D=>nx5869, 
      CLK=>nx15607);
   ix6335 : oai22 port map ( Y=>nx6334, A0=>nx13174, A1=>nx16329, B0=>
      nx13177, B1=>nx16345);
   modgen_ram_ix74_ix1920 : dff port map ( Q=>OPEN, QB=>nx13174, D=>nx5849, 
      CLK=>nx15607);
   modgen_ram_ix74_ix1916 : dff port map ( Q=>OPEN, QB=>nx13177, D=>nx5859, 
      CLK=>nx15607);
   modgen_ram_ix74_ix2044 : dff port map ( Q=>OPEN, QB=>nx13184, D=>nx5839, 
      CLK=>nx15607);
   modgen_ram_ix74_ix2108 : dff port map ( Q=>OPEN, QB=>nx13188, D=>nx5829, 
      CLK=>nx15607);
   ix6293 : oai22 port map ( Y=>nx6292, A0=>nx13192, A1=>nx16361, B0=>
      nx13195, B1=>nx16377);
   modgen_ram_ix74_ix2088 : dff port map ( Q=>OPEN, QB=>nx13192, D=>nx5809, 
      CLK=>nx15607);
   modgen_ram_ix74_ix2024 : dff port map ( Q=>OPEN, QB=>nx13195, D=>nx5819, 
      CLK=>nx15607);
   modgen_ram_ix74_ix2152 : dff port map ( Q=>OPEN, QB=>nx13201, D=>nx5799, 
      CLK=>nx15609);
   modgen_ram_ix74_ix1964 : dff port map ( Q=>OPEN, QB=>nx13205, D=>nx5789, 
      CLK=>nx15609);
   ix6255 : oai22 port map ( Y=>nx6254, A0=>nx13209, A1=>nx16401, B0=>
      nx13212, B1=>nx16417);
   modgen_ram_ix74_ix2092 : dff port map ( Q=>OPEN, QB=>nx13209, D=>nx5769, 
      CLK=>nx15609);
   modgen_ram_ix74_ix2028 : dff port map ( Q=>OPEN, QB=>nx13212, D=>nx5779, 
      CLK=>nx15609);
   modgen_ram_ix74_ix2156 : dff port map ( Q=>OPEN, QB=>nx13218, D=>nx5759, 
      CLK=>nx15609);
   modgen_ram_ix74_ix1968 : dff port map ( Q=>OPEN, QB=>nx13222, D=>nx5749, 
      CLK=>nx15609);
   ix6215 : oai22 port map ( Y=>nx6214, A0=>nx13226, A1=>nx16441, B0=>
      nx13229, B1=>nx16457);
   modgen_ram_ix74_ix2096 : dff port map ( Q=>OPEN, QB=>nx13226, D=>nx5729, 
      CLK=>nx15609);
   modgen_ram_ix74_ix2032 : dff port map ( Q=>OPEN, QB=>nx13229, D=>nx5739, 
      CLK=>nx15611);
   modgen_ram_ix74_ix2160 : dff port map ( Q=>OPEN, QB=>nx13235, D=>nx5719, 
      CLK=>nx15611);
   ix6185 : nor03_2x port map ( Y=>nx6184, A0=>nx13239, A1=>nx15433, A2=>
      nx15961);
   modgen_ram_ix74_ix1972 : dff port map ( Q=>OPEN, QB=>nx13239, D=>nx5709, 
      CLK=>nx15611);
   ix6177 : oai22 port map ( Y=>nx6176, A0=>nx13243, A1=>nx16481, B0=>
      nx13246, B1=>nx16497);
   modgen_ram_ix74_ix2100 : dff port map ( Q=>OPEN, QB=>nx13243, D=>nx5689, 
      CLK=>nx15611);
   modgen_ram_ix74_ix2036 : dff port map ( Q=>OPEN, QB=>nx13246, D=>nx5699, 
      CLK=>nx15611);
   ix6151 : oai22 port map ( Y=>nx6150, A0=>nx13256, A1=>nx16513, B0=>
      nx13259, B1=>nx16521);
   modgen_ram_ix74_ix2128 : dff port map ( Q=>OPEN, QB=>nx13256, D=>nx5669, 
      CLK=>nx15611);
   modgen_ram_ix74_ix2164 : dff port map ( Q=>OPEN, QB=>nx13259, D=>nx5679, 
      CLK=>nx15611);
   ix6133 : oai22 port map ( Y=>nx6132, A0=>nx13263, A1=>nx16529, B0=>
      nx13266, B1=>nx16545);
   modgen_ram_ix74_ix2060 : dff port map ( Q=>OPEN, QB=>nx13263, D=>nx5659, 
      CLK=>nx15613);
   modgen_ram_ix74_ix1996 : dff port map ( Q=>OPEN, QB=>nx13266, D=>nx5649, 
      CLK=>nx15613);
   ix6115 : nand03 port map ( Y=>nx6114, A0=>nx13270, A1=>nx13280, A2=>
      nx13286);
   ix13271 : nor02_2x port map ( Y=>nx13270, A0=>nx6110, A1=>nx6102);
   ix6111 : nor04 port map ( Y=>nx6110, A0=>nx13273, A1=>address(4), A2=>
      address(5), A3=>nx15901);
   modgen_ram_ix74_ix2120 : dff port map ( Q=>OPEN, QB=>nx13273, D=>nx5639, 
      CLK=>nx15613);
   ix6103 : nor03_2x port map ( Y=>nx6102, A0=>nx13277, A1=>nx15825, A2=>
      nx15901);
   modgen_ram_ix74_ix2056 : dff port map ( Q=>OPEN, QB=>nx13277, D=>nx5629, 
      CLK=>nx15613);
   ix13281 : nand03 port map ( Y=>nx13280, A0=>modgen_ram_ix74_a_12_dup_685, 
      A1=>nx16231, A2=>nx16571);
   modgen_ram_ix74_ix2116 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_685, 
      QB=>nx13284, D=>nx5619, CLK=>nx15613);
   ix13287 : nand03 port map ( Y=>nx13286, A0=>modgen_ram_ix74_a_28_dup_669, 
      A1=>nx16197, A2=>nx16571);
   modgen_ram_ix74_ix2052 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_669, 
      QB=>nx13290, D=>nx5609, CLK=>nx15613);
   ix13293 : nor03_2x port map ( Y=>nx13292, A0=>nx6070, A1=>nx6062, A2=>
      nx6054);
   ix6071 : nor03_2x port map ( Y=>nx6070, A0=>nx13295, A1=>nx15435, A2=>
      nx15931);
   modgen_ram_ix74_ix1924 : dff port map ( Q=>OPEN, QB=>nx13295, D=>nx5599, 
      CLK=>nx15613);
   ix6063 : nor03_2x port map ( Y=>nx6062, A0=>nx13299, A1=>nx15775, A2=>
      nx15891);
   modgen_ram_ix74_ix2000 : dff port map ( Q=>OPEN, QB=>nx13299, D=>nx5589, 
      CLK=>nx15615);
   ix6055 : oai22 port map ( Y=>nx6054, A0=>nx13303, A1=>nx16605, B0=>
      nx13306, B1=>nx16621);
   modgen_ram_ix74_ix1992 : dff port map ( Q=>OPEN, QB=>nx13303, D=>nx5579, 
      CLK=>nx15615);
   modgen_ram_ix74_ix1988 : dff port map ( Q=>OPEN, QB=>nx13306, D=>nx5569, 
      CLK=>nx15615);
   ix13310 : nor03_2x port map ( Y=>nx13309, A0=>nx6032, A1=>nx6024, A2=>
      nx6016);
   ix6033 : nor03_2x port map ( Y=>nx6032, A0=>nx13312, A1=>nx15861, A2=>
      nx15915);
   modgen_ram_ix74_ix2112 : dff port map ( Q=>OPEN, QB=>nx13312, D=>nx5559, 
      CLK=>nx15615);
   ix6025 : nor03_2x port map ( Y=>nx6024, A0=>nx13316, A1=>nx15435, A2=>
      nx15901);
   modgen_ram_ix74_ix1928 : dff port map ( Q=>OPEN, QB=>nx13316, D=>nx5549, 
      CLK=>nx15615);
   ix6017 : oai22 port map ( Y=>nx6016, A0=>nx13320, A1=>nx16645, B0=>
      nx13323, B1=>nx16661);
   modgen_ram_ix74_ix1936 : dff port map ( Q=>OPEN, QB=>nx13320, D=>nx5539, 
      CLK=>nx15615);
   modgen_ram_ix74_ix1932 : dff port map ( Q=>OPEN, QB=>nx13323, D=>nx5529, 
      CLK=>nx15615);
   ix5993 : oai22 port map ( Y=>nx5992, A0=>nx13330, A1=>nx16677, B0=>
      nx13333, B1=>nx16693);
   modgen_ram_ix74_ix2080 : dff port map ( Q=>OPEN, QB=>nx13330, D=>nx5509, 
      CLK=>nx15617);
   modgen_ram_ix74_ix2124 : dff port map ( Q=>OPEN, QB=>nx13333, D=>nx5519, 
      CLK=>nx15617);
   ix5975 : oai22 port map ( Y=>nx5974, A0=>nx13337, A1=>nx16709, B0=>
      nx13340, B1=>nx16725);
   modgen_ram_ix74_ix2140 : dff port map ( Q=>OPEN, QB=>nx13337, D=>nx5499, 
      CLK=>nx15617);
   modgen_ram_ix74_ix2076 : dff port map ( Q=>OPEN, QB=>nx13340, D=>nx5489, 
      CLK=>nx15617);
   ix13344 : nor03_2x port map ( Y=>nx13343, A0=>nx5952, A1=>nx5944, A2=>
      nx5936);
   ix5953 : nor03_2x port map ( Y=>nx5952, A0=>nx13346, A1=>nx15435, A2=>
      nx15755);
   modgen_ram_ix74_ix1948 : dff port map ( Q=>OPEN, QB=>nx13346, D=>nx5479, 
      CLK=>nx15617);
   ix5945 : nor03_2x port map ( Y=>nx5944, A0=>nx13350, A1=>nx15861, A2=>
      nx15803);
   modgen_ram_ix74_ix2136 : dff port map ( Q=>OPEN, QB=>nx13350, D=>nx5469, 
      CLK=>nx15617);
   ix5937 : oai22 port map ( Y=>nx5936, A0=>nx13354, A1=>nx16749, B0=>
      nx13357, B1=>nx16757);
   modgen_ram_ix74_ix1944 : dff port map ( Q=>OPEN, QB=>nx13354, D=>nx5459, 
      CLK=>nx15617);
   modgen_ram_ix74_ix2132 : dff port map ( Q=>OPEN, QB=>nx13357, D=>nx5449, 
      CLK=>nx15619);
   ix13361 : nor03_2x port map ( Y=>nx13360, A0=>nx5912, A1=>nx5904, A2=>
      nx5896);
   ix5913 : nor03_2x port map ( Y=>nx5912, A0=>nx13363, A1=>nx15775, A2=>
      nx15815);
   modgen_ram_ix74_ix2004 : dff port map ( Q=>OPEN, QB=>nx13363, D=>nx5439, 
      CLK=>nx15619);
   ix5905 : nor03_2x port map ( Y=>nx5904, A0=>nx13367, A1=>nx15825, A2=>
      nx15803);
   modgen_ram_ix74_ix2072 : dff port map ( Q=>OPEN, QB=>nx13367, D=>nx5429, 
      CLK=>nx15619);
   ix5897 : oai22 port map ( Y=>nx5896, A0=>nx13371, A1=>nx16773, B0=>
      nx13374, B1=>nx16789);
   modgen_ram_ix74_ix2068 : dff port map ( Q=>OPEN, QB=>nx13371, D=>nx5419, 
      CLK=>nx15619);
   modgen_ram_ix74_ix1940 : dff port map ( Q=>OPEN, QB=>nx13374, D=>nx5409, 
      CLK=>nx15619);
   ix13378 : nor03_2x port map ( Y=>nx13377, A0=>nx5874, A1=>nx5866, A2=>
      nx5858);
   ix5875 : nor03_2x port map ( Y=>nx5874, A0=>nx13380, A1=>nx15775, A2=>
      nx15805);
   modgen_ram_ix74_ix2008 : dff port map ( Q=>OPEN, QB=>nx13380, D=>nx5399, 
      CLK=>nx15619);
   ix5867 : nor03_2x port map ( Y=>nx5866, A0=>nx13384, A1=>nx15777, A2=>
      nx15407);
   modgen_ram_ix74_ix2016 : dff port map ( Q=>OPEN, QB=>nx13384, D=>nx5389, 
      CLK=>nx15619);
   ix5859 : oai22 port map ( Y=>nx5858, A0=>nx13388, A1=>nx16821, B0=>
      nx13391, B1=>nx16837);
   modgen_ram_ix74_ix1952 : dff port map ( Q=>OPEN, QB=>nx13388, D=>nx5369, 
      CLK=>nx15621);
   modgen_ram_ix74_ix2012 : dff port map ( Q=>OPEN, QB=>nx13391, D=>nx5379, 
      CLK=>nx15621);
   tri_data_out_9 : tri01 port map ( Y=>data_out(9), A=>nx13395, E=>
      write_out);
   ix7107 : oai22 port map ( Y=>nx7106, A0=>nx13401, A1=>nx16159, B0=>
      nx13406, B1=>nx16185);
   modgen_ram_ix74_ix1699 : dff port map ( Q=>OPEN, QB=>nx13401, D=>nx6639, 
      CLK=>nx15621);
   modgen_ram_ix74_ix1807 : dff port map ( Q=>OPEN, QB=>nx13406, D=>nx6629, 
      CLK=>nx15621);
   ix7089 : oai22 port map ( Y=>nx7088, A0=>nx13410, A1=>nx16203, B0=>
      nx13413, B1=>nx18957);
   modgen_ram_ix74_ix1783 : dff port map ( Q=>OPEN, QB=>nx13410, D=>nx6609, 
      CLK=>nx15621);
   modgen_ram_ix74_ix1791 : dff port map ( Q=>OPEN, QB=>nx13413, D=>nx6619, 
      CLK=>nx15621);
   ix13417 : nor02_2x port map ( Y=>nx13416, A0=>nx7068, A1=>nx7050);
   ix7069 : oai33 port map ( Y=>nx7068, A0=>nx13419, A1=>nx15861, A2=>
      nx16095, B0=>nx13422, B1=>nx15435, B2=>nx16025);
   modgen_ram_ix74_ix1891 : dff port map ( Q=>OPEN, QB=>nx13419, D=>nx6589, 
      CLK=>nx15621);
   modgen_ram_ix74_ix1703 : dff port map ( Q=>OPEN, QB=>nx13422, D=>nx6599, 
      CLK=>nx15623);
   ix7051 : oai22 port map ( Y=>nx7050, A0=>nx13426, A1=>nx16261, B0=>
      nx13429, B1=>nx16277);
   modgen_ram_ix74_ix1827 : dff port map ( Q=>OPEN, QB=>nx13426, D=>nx6579, 
      CLK=>nx15623);
   modgen_ram_ix74_ix1763 : dff port map ( Q=>OPEN, QB=>nx13429, D=>nx6569, 
      CLK=>nx15623);
   ix13433 : nor03_2x port map ( Y=>nx13432, A0=>nx7026, A1=>nx7018, A2=>
      nx7010);
   ix7027 : nor03_2x port map ( Y=>nx7026, A0=>nx13435, A1=>nx15777, A2=>
      nx16067);
   modgen_ram_ix74_ix1719 : dff port map ( Q=>OPEN, QB=>nx13435, D=>nx6559, 
      CLK=>nx15623);
   ix7019 : nor03_2x port map ( Y=>nx7018, A0=>nx13439, A1=>nx15861, A2=>
      nx15409);
   modgen_ram_ix74_ix1887 : dff port map ( Q=>OPEN, QB=>nx13439, D=>nx6549, 
      CLK=>nx15623);
   ix7011 : oai33 port map ( Y=>nx7010, A0=>nx13443, A1=>nx15777, A2=>
      nx15915, B0=>nx13446, B1=>nx15435, B2=>nx16069);
   modgen_ram_ix74_ix1727 : dff port map ( Q=>OPEN, QB=>nx13443, D=>nx6529, 
      CLK=>nx15623);
   modgen_ram_ix74_ix1655 : dff port map ( Q=>OPEN, QB=>nx13446, D=>nx6539, 
      CLK=>nx15623);
   ix13450 : nor03_2x port map ( Y=>nx13449, A0=>nx6988, A1=>nx6980, A2=>
      nx6972);
   ix6989 : nor03_2x port map ( Y=>nx6988, A0=>nx13452, A1=>nx15777, A2=>
      nx16047);
   modgen_ram_ix74_ix1723 : dff port map ( Q=>OPEN, QB=>nx13452, D=>nx6519, 
      CLK=>nx15625);
   ix6981 : nor04 port map ( Y=>nx6980, A0=>nx13456, A1=>address(4), A2=>
      address(5), A3=>nx16069);
   modgen_ram_ix74_ix1847 : dff port map ( Q=>OPEN, QB=>nx13456, D=>nx6509, 
      CLK=>nx15625);
   ix6973 : oai22 port map ( Y=>nx6972, A0=>nx13460, A1=>nx16329, B0=>
      nx13463, B1=>nx16345);
   modgen_ram_ix74_ix1663 : dff port map ( Q=>OPEN, QB=>nx13460, D=>nx6489, 
      CLK=>nx15625);
   modgen_ram_ix74_ix1659 : dff port map ( Q=>OPEN, QB=>nx13463, D=>nx6499, 
      CLK=>nx15625);
   modgen_ram_ix74_ix1787 : dff port map ( Q=>OPEN, QB=>nx13470, D=>nx6479, 
      CLK=>nx15625);
   modgen_ram_ix74_ix1851 : dff port map ( Q=>OPEN, QB=>nx13474, D=>nx6469, 
      CLK=>nx15625);
   ix6931 : oai22 port map ( Y=>nx6930, A0=>nx13478, A1=>nx16361, B0=>
      nx13481, B1=>nx16377);
   modgen_ram_ix74_ix1831 : dff port map ( Q=>OPEN, QB=>nx13478, D=>nx6449, 
      CLK=>nx15625);
   modgen_ram_ix74_ix1767 : dff port map ( Q=>OPEN, QB=>nx13481, D=>nx6459, 
      CLK=>nx15627);
   modgen_ram_ix74_ix1895 : dff port map ( Q=>OPEN, QB=>nx13487, D=>nx6439, 
      CLK=>nx15627);
   modgen_ram_ix74_ix1707 : dff port map ( Q=>OPEN, QB=>nx13491, D=>nx6429, 
      CLK=>nx15627);
   ix6893 : oai22 port map ( Y=>nx6892, A0=>nx13495, A1=>nx16401, B0=>
      nx13498, B1=>nx16417);
   modgen_ram_ix74_ix1835 : dff port map ( Q=>OPEN, QB=>nx13495, D=>nx6409, 
      CLK=>nx15627);
   modgen_ram_ix74_ix1771 : dff port map ( Q=>OPEN, QB=>nx13498, D=>nx6419, 
      CLK=>nx15627);
   modgen_ram_ix74_ix1899 : dff port map ( Q=>OPEN, QB=>nx13504, D=>nx6399, 
      CLK=>nx15627);
   modgen_ram_ix74_ix1711 : dff port map ( Q=>OPEN, QB=>nx13508, D=>nx6389, 
      CLK=>nx15627);
   ix6853 : oai22 port map ( Y=>nx6852, A0=>nx13512, A1=>nx16441, B0=>
      nx13515, B1=>nx16457);
   modgen_ram_ix74_ix1839 : dff port map ( Q=>OPEN, QB=>nx13512, D=>nx6369, 
      CLK=>nx15629);
   modgen_ram_ix74_ix1775 : dff port map ( Q=>OPEN, QB=>nx13515, D=>nx6379, 
      CLK=>nx15629);
   modgen_ram_ix74_ix1903 : dff port map ( Q=>OPEN, QB=>nx13521, D=>nx6359, 
      CLK=>nx15629);
   ix6823 : nor03_2x port map ( Y=>nx6822, A0=>nx13525, A1=>nx15437, A2=>
      nx15961);
   modgen_ram_ix74_ix1715 : dff port map ( Q=>OPEN, QB=>nx13525, D=>nx6349, 
      CLK=>nx15629);
   ix6815 : oai22 port map ( Y=>nx6814, A0=>nx13529, A1=>nx16481, B0=>
      nx13532, B1=>nx16497);
   modgen_ram_ix74_ix1843 : dff port map ( Q=>OPEN, QB=>nx13529, D=>nx6329, 
      CLK=>nx15629);
   modgen_ram_ix74_ix1779 : dff port map ( Q=>OPEN, QB=>nx13532, D=>nx6339, 
      CLK=>nx15629);
   ix6789 : oai22 port map ( Y=>nx6788, A0=>nx13542, A1=>nx16513, B0=>
      nx13545, B1=>nx16521);
   modgen_ram_ix74_ix1871 : dff port map ( Q=>OPEN, QB=>nx13542, D=>nx6309, 
      CLK=>nx15629);
   modgen_ram_ix74_ix1907 : dff port map ( Q=>OPEN, QB=>nx13545, D=>nx6319, 
      CLK=>nx15631);
   ix6771 : oai22 port map ( Y=>nx6770, A0=>nx13549, A1=>nx16529, B0=>
      nx13552, B1=>nx16545);
   modgen_ram_ix74_ix1803 : dff port map ( Q=>OPEN, QB=>nx13549, D=>nx6299, 
      CLK=>nx15631);
   modgen_ram_ix74_ix1739 : dff port map ( Q=>OPEN, QB=>nx13552, D=>nx6289, 
      CLK=>nx15631);
   ix6753 : nand03 port map ( Y=>nx6752, A0=>nx13556, A1=>nx13566, A2=>
      nx13572);
   ix13557 : nor02_2x port map ( Y=>nx13556, A0=>nx6748, A1=>nx6740);
   ix6749 : nor04 port map ( Y=>nx6748, A0=>nx13559, A1=>address(4), A2=>
      address(5), A3=>nx15903);
   modgen_ram_ix74_ix1863 : dff port map ( Q=>OPEN, QB=>nx13559, D=>nx6279, 
      CLK=>nx15631);
   ix6741 : nor03_2x port map ( Y=>nx6740, A0=>nx13563, A1=>nx15827, A2=>
      nx15903);
   modgen_ram_ix74_ix1799 : dff port map ( Q=>OPEN, QB=>nx13563, D=>nx6269, 
      CLK=>nx15631);
   ix13567 : nand03 port map ( Y=>nx13566, A0=>modgen_ram_ix74_a_12_dup_620, 
      A1=>nx16231, A2=>nx16573);
   modgen_ram_ix74_ix1859 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_620, 
      QB=>nx13570, D=>nx6259, CLK=>nx15631);
   ix13573 : nand03 port map ( Y=>nx13572, A0=>modgen_ram_ix74_a_28_dup_604, 
      A1=>nx16197, A2=>nx16573);
   modgen_ram_ix74_ix1795 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_604, 
      QB=>nx13576, D=>nx6249, CLK=>nx15631);
   ix13579 : nor03_2x port map ( Y=>nx13578, A0=>nx6708, A1=>nx6700, A2=>
      nx6692);
   ix6709 : nor03_2x port map ( Y=>nx6708, A0=>nx13581, A1=>nx15437, A2=>
      nx15931);
   modgen_ram_ix74_ix1667 : dff port map ( Q=>OPEN, QB=>nx13581, D=>nx6239, 
      CLK=>nx15633);
   ix6701 : nor03_2x port map ( Y=>nx6700, A0=>nx13585, A1=>nx15777, A2=>
      nx15891);
   modgen_ram_ix74_ix1743 : dff port map ( Q=>OPEN, QB=>nx13585, D=>nx6229, 
      CLK=>nx15633);
   ix6693 : oai22 port map ( Y=>nx6692, A0=>nx13589, A1=>nx16605, B0=>
      nx13592, B1=>nx16621);
   modgen_ram_ix74_ix1735 : dff port map ( Q=>OPEN, QB=>nx13589, D=>nx6219, 
      CLK=>nx15633);
   modgen_ram_ix74_ix1731 : dff port map ( Q=>OPEN, QB=>nx13592, D=>nx6209, 
      CLK=>nx15633);
   ix13596 : nor03_2x port map ( Y=>nx13595, A0=>nx6670, A1=>nx6662, A2=>
      nx6654);
   ix6671 : nor03_2x port map ( Y=>nx6670, A0=>nx13598, A1=>nx15861, A2=>
      nx15917);
   modgen_ram_ix74_ix1855 : dff port map ( Q=>OPEN, QB=>nx13598, D=>nx6199, 
      CLK=>nx15633);
   ix6663 : nor03_2x port map ( Y=>nx6662, A0=>nx13602, A1=>nx15437, A2=>
      nx15903);
   modgen_ram_ix74_ix1671 : dff port map ( Q=>OPEN, QB=>nx13602, D=>nx6189, 
      CLK=>nx15633);
   ix6655 : oai22 port map ( Y=>nx6654, A0=>nx13606, A1=>nx16645, B0=>
      nx13609, B1=>nx16661);
   modgen_ram_ix74_ix1679 : dff port map ( Q=>OPEN, QB=>nx13606, D=>nx6179, 
      CLK=>nx15633);
   modgen_ram_ix74_ix1675 : dff port map ( Q=>OPEN, QB=>nx13609, D=>nx6169, 
      CLK=>nx15635);
   ix6631 : oai22 port map ( Y=>nx6630, A0=>nx13616, A1=>nx16677, B0=>
      nx13619, B1=>nx16693);
   modgen_ram_ix74_ix1823 : dff port map ( Q=>OPEN, QB=>nx13616, D=>nx6149, 
      CLK=>nx15635);
   modgen_ram_ix74_ix1867 : dff port map ( Q=>OPEN, QB=>nx13619, D=>nx6159, 
      CLK=>nx15635);
   ix6613 : oai22 port map ( Y=>nx6612, A0=>nx13623, A1=>nx16709, B0=>
      nx13626, B1=>nx16725);
   modgen_ram_ix74_ix1883 : dff port map ( Q=>OPEN, QB=>nx13623, D=>nx6139, 
      CLK=>nx15635);
   modgen_ram_ix74_ix1819 : dff port map ( Q=>OPEN, QB=>nx13626, D=>nx6129, 
      CLK=>nx15635);
   ix13630 : nor03_2x port map ( Y=>nx13629, A0=>nx6590, A1=>nx6582, A2=>
      nx6574);
   ix6591 : nor03_2x port map ( Y=>nx6590, A0=>nx13632, A1=>nx15437, A2=>
      nx15755);
   modgen_ram_ix74_ix1691 : dff port map ( Q=>OPEN, QB=>nx13632, D=>nx6119, 
      CLK=>nx15635);
   ix6583 : nor03_2x port map ( Y=>nx6582, A0=>nx13636, A1=>nx15863, A2=>
      nx15805);
   modgen_ram_ix74_ix1879 : dff port map ( Q=>OPEN, QB=>nx13636, D=>nx6109, 
      CLK=>nx15635);
   ix6575 : oai22 port map ( Y=>nx6574, A0=>nx13640, A1=>nx16749, B0=>
      nx13643, B1=>nx16757);
   modgen_ram_ix74_ix1687 : dff port map ( Q=>OPEN, QB=>nx13640, D=>nx6099, 
      CLK=>nx15637);
   modgen_ram_ix74_ix1875 : dff port map ( Q=>OPEN, QB=>nx13643, D=>nx6089, 
      CLK=>nx15637);
   ix13647 : nor03_2x port map ( Y=>nx13646, A0=>nx6550, A1=>nx6542, A2=>
      nx6534);
   ix6551 : nor03_2x port map ( Y=>nx6550, A0=>nx13649, A1=>nx15777, A2=>
      nx15815);
   modgen_ram_ix74_ix1747 : dff port map ( Q=>OPEN, QB=>nx13649, D=>nx6079, 
      CLK=>nx15637);
   ix6543 : nor03_2x port map ( Y=>nx6542, A0=>nx13653, A1=>nx15827, A2=>
      nx15805);
   modgen_ram_ix74_ix1815 : dff port map ( Q=>OPEN, QB=>nx13653, D=>nx6069, 
      CLK=>nx15637);
   ix6535 : oai22 port map ( Y=>nx6534, A0=>nx13657, A1=>nx16773, B0=>
      nx13660, B1=>nx16789);
   modgen_ram_ix74_ix1811 : dff port map ( Q=>OPEN, QB=>nx13657, D=>nx6059, 
      CLK=>nx15637);
   modgen_ram_ix74_ix1683 : dff port map ( Q=>OPEN, QB=>nx13660, D=>nx6049, 
      CLK=>nx15637);
   ix13664 : nor03_2x port map ( Y=>nx13663, A0=>nx6512, A1=>nx6504, A2=>
      nx6496);
   ix6513 : nor03_2x port map ( Y=>nx6512, A0=>nx13666, A1=>nx15777, A2=>
      nx15805);
   modgen_ram_ix74_ix1751 : dff port map ( Q=>OPEN, QB=>nx13666, D=>nx6039, 
      CLK=>nx15637);
   ix6505 : nor03_2x port map ( Y=>nx6504, A0=>nx13670, A1=>nx15779, A2=>
      nx15409);
   modgen_ram_ix74_ix1759 : dff port map ( Q=>OPEN, QB=>nx13670, D=>nx6029, 
      CLK=>nx15639);
   ix6497 : oai22 port map ( Y=>nx6496, A0=>nx13674, A1=>nx16821, B0=>
      nx13677, B1=>nx16837);
   modgen_ram_ix74_ix1695 : dff port map ( Q=>OPEN, QB=>nx13674, D=>nx6009, 
      CLK=>nx15639);
   modgen_ram_ix74_ix1755 : dff port map ( Q=>OPEN, QB=>nx13677, D=>nx6019, 
      CLK=>nx15639);
   tri_data_out_10 : tri01 port map ( Y=>data_out(10), A=>nx13681, E=>
      write_out);
   ix7745 : oai22 port map ( Y=>nx7744, A0=>nx13687, A1=>nx16159, B0=>
      nx13692, B1=>nx16185);
   modgen_ram_ix74_ix1442 : dff port map ( Q=>OPEN, QB=>nx13687, D=>nx7279, 
      CLK=>nx15639);
   modgen_ram_ix74_ix1550 : dff port map ( Q=>OPEN, QB=>nx13692, D=>nx7269, 
      CLK=>nx15639);
   ix7727 : oai22 port map ( Y=>nx7726, A0=>nx13696, A1=>nx16203, B0=>
      nx13699, B1=>nx18958);
   modgen_ram_ix74_ix1526 : dff port map ( Q=>OPEN, QB=>nx13696, D=>nx7249, 
      CLK=>nx15639);
   modgen_ram_ix74_ix1534 : dff port map ( Q=>OPEN, QB=>nx13699, D=>nx7259, 
      CLK=>nx15639);
   ix13703 : nor02_2x port map ( Y=>nx13702, A0=>nx7706, A1=>nx7688);
   ix7707 : oai33 port map ( Y=>nx7706, A0=>nx13705, A1=>nx15863, A2=>
      nx16095, B0=>nx13708, B1=>nx15437, B2=>nx16027);
   modgen_ram_ix74_ix1634 : dff port map ( Q=>OPEN, QB=>nx13705, D=>nx7229, 
      CLK=>nx15641);
   modgen_ram_ix74_ix1446 : dff port map ( Q=>OPEN, QB=>nx13708, D=>nx7239, 
      CLK=>nx15641);
   ix7689 : oai22 port map ( Y=>nx7688, A0=>nx13712, A1=>nx16261, B0=>
      nx13715, B1=>nx16277);
   modgen_ram_ix74_ix1570 : dff port map ( Q=>OPEN, QB=>nx13712, D=>nx7219, 
      CLK=>nx15641);
   modgen_ram_ix74_ix1506 : dff port map ( Q=>OPEN, QB=>nx13715, D=>nx7209, 
      CLK=>nx15641);
   ix13719 : nor03_2x port map ( Y=>nx13718, A0=>nx7664, A1=>nx7656, A2=>
      nx7648);
   ix7665 : nor03_2x port map ( Y=>nx7664, A0=>nx13721, A1=>nx15779, A2=>
      nx16069);
   modgen_ram_ix74_ix1462 : dff port map ( Q=>OPEN, QB=>nx13721, D=>nx7199, 
      CLK=>nx15641);
   ix7657 : nor03_2x port map ( Y=>nx7656, A0=>nx13725, A1=>nx15863, A2=>
      nx15409);
   modgen_ram_ix74_ix1630 : dff port map ( Q=>OPEN, QB=>nx13725, D=>nx7189, 
      CLK=>nx15641);
   ix7649 : oai33 port map ( Y=>nx7648, A0=>nx13729, A1=>nx15779, A2=>
      nx15917, B0=>nx13732, B1=>nx15437, B2=>nx16069);
   modgen_ram_ix74_ix1470 : dff port map ( Q=>OPEN, QB=>nx13729, D=>nx7169, 
      CLK=>nx15641);
   modgen_ram_ix74_ix1398 : dff port map ( Q=>OPEN, QB=>nx13732, D=>nx7179, 
      CLK=>nx15643);
   ix13736 : nor03_2x port map ( Y=>nx13735, A0=>nx7626, A1=>nx7618, A2=>
      nx7610);
   ix7627 : nor03_2x port map ( Y=>nx7626, A0=>nx13738, A1=>nx15779, A2=>
      nx16047);
   modgen_ram_ix74_ix1466 : dff port map ( Q=>OPEN, QB=>nx13738, D=>nx7159, 
      CLK=>nx15643);
   ix7619 : nor04 port map ( Y=>nx7618, A0=>nx13742, A1=>address(4), A2=>
      address(5), A3=>nx16069);
   modgen_ram_ix74_ix1590 : dff port map ( Q=>OPEN, QB=>nx13742, D=>nx7149, 
      CLK=>nx15643);
   ix7611 : oai22 port map ( Y=>nx7610, A0=>nx13746, A1=>nx16329, B0=>
      nx13749, B1=>nx16345);
   modgen_ram_ix74_ix1406 : dff port map ( Q=>OPEN, QB=>nx13746, D=>nx7129, 
      CLK=>nx15643);
   modgen_ram_ix74_ix1402 : dff port map ( Q=>OPEN, QB=>nx13749, D=>nx7139, 
      CLK=>nx15643);
   modgen_ram_ix74_ix1530 : dff port map ( Q=>OPEN, QB=>nx13756, D=>nx7119, 
      CLK=>nx15643);
   modgen_ram_ix74_ix1594 : dff port map ( Q=>OPEN, QB=>nx13760, D=>nx7109, 
      CLK=>nx15643);
   ix7569 : oai22 port map ( Y=>nx7568, A0=>nx13764, A1=>nx16361, B0=>
      nx13767, B1=>nx16377);
   modgen_ram_ix74_ix1574 : dff port map ( Q=>OPEN, QB=>nx13764, D=>nx7089, 
      CLK=>nx15645);
   modgen_ram_ix74_ix1510 : dff port map ( Q=>OPEN, QB=>nx13767, D=>nx7099, 
      CLK=>nx15645);
   modgen_ram_ix74_ix1638 : dff port map ( Q=>OPEN, QB=>nx13773, D=>nx7079, 
      CLK=>nx15645);
   modgen_ram_ix74_ix1450 : dff port map ( Q=>OPEN, QB=>nx13777, D=>nx7069, 
      CLK=>nx15645);
   ix7531 : oai22 port map ( Y=>nx7530, A0=>nx13781, A1=>nx16401, B0=>
      nx13784, B1=>nx16417);
   modgen_ram_ix74_ix1578 : dff port map ( Q=>OPEN, QB=>nx13781, D=>nx7049, 
      CLK=>nx15645);
   modgen_ram_ix74_ix1514 : dff port map ( Q=>OPEN, QB=>nx13784, D=>nx7059, 
      CLK=>nx15645);
   modgen_ram_ix74_ix1642 : dff port map ( Q=>OPEN, QB=>nx13790, D=>nx7039, 
      CLK=>nx15645);
   modgen_ram_ix74_ix1454 : dff port map ( Q=>OPEN, QB=>nx13794, D=>nx7029, 
      CLK=>nx15647);
   ix7491 : oai22 port map ( Y=>nx7490, A0=>nx13798, A1=>nx16441, B0=>
      nx13801, B1=>nx16457);
   modgen_ram_ix74_ix1582 : dff port map ( Q=>OPEN, QB=>nx13798, D=>nx7009, 
      CLK=>nx15647);
   modgen_ram_ix74_ix1518 : dff port map ( Q=>OPEN, QB=>nx13801, D=>nx7019, 
      CLK=>nx15647);
   modgen_ram_ix74_ix1646 : dff port map ( Q=>OPEN, QB=>nx13807, D=>nx6999, 
      CLK=>nx15647);
   ix7461 : nor03_2x port map ( Y=>nx7460, A0=>nx13811, A1=>nx15439, A2=>
      nx15961);
   modgen_ram_ix74_ix1458 : dff port map ( Q=>OPEN, QB=>nx13811, D=>nx6989, 
      CLK=>nx15647);
   ix7453 : oai22 port map ( Y=>nx7452, A0=>nx13815, A1=>nx16481, B0=>
      nx13818, B1=>nx16497);
   modgen_ram_ix74_ix1586 : dff port map ( Q=>OPEN, QB=>nx13815, D=>nx6969, 
      CLK=>nx15647);
   modgen_ram_ix74_ix1522 : dff port map ( Q=>OPEN, QB=>nx13818, D=>nx6979, 
      CLK=>nx15647);
   ix7427 : oai22 port map ( Y=>nx7426, A0=>nx13828, A1=>nx16513, B0=>
      nx13831, B1=>nx16521);
   modgen_ram_ix74_ix1614 : dff port map ( Q=>OPEN, QB=>nx13828, D=>nx6949, 
      CLK=>nx15649);
   modgen_ram_ix74_ix1650 : dff port map ( Q=>OPEN, QB=>nx13831, D=>nx6959, 
      CLK=>nx15649);
   ix7409 : oai22 port map ( Y=>nx7408, A0=>nx13835, A1=>nx16529, B0=>
      nx13838, B1=>nx16545);
   modgen_ram_ix74_ix1546 : dff port map ( Q=>OPEN, QB=>nx13835, D=>nx6939, 
      CLK=>nx15649);
   modgen_ram_ix74_ix1482 : dff port map ( Q=>OPEN, QB=>nx13838, D=>nx6929, 
      CLK=>nx15649);
   ix7391 : nand03 port map ( Y=>nx7390, A0=>nx13842, A1=>nx13852, A2=>
      nx13858);
   ix13843 : nor02_2x port map ( Y=>nx13842, A0=>nx7386, A1=>nx7378);
   ix7387 : nor04 port map ( Y=>nx7386, A0=>nx13845, A1=>address(4), A2=>
      address(5), A3=>nx15903);
   modgen_ram_ix74_ix1606 : dff port map ( Q=>OPEN, QB=>nx13845, D=>nx6919, 
      CLK=>nx15649);
   ix7379 : nor03_2x port map ( Y=>nx7378, A0=>nx13849, A1=>nx15827, A2=>
      nx15903);
   modgen_ram_ix74_ix1542 : dff port map ( Q=>OPEN, QB=>nx13849, D=>nx6909, 
      CLK=>nx15649);
   ix13853 : nand03 port map ( Y=>nx13852, A0=>modgen_ram_ix74_a_12_dup_554, 
      A1=>nx16231, A2=>nx16573);
   modgen_ram_ix74_ix1602 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_554, 
      QB=>nx13856, D=>nx6899, CLK=>nx15649);
   ix13859 : nand03 port map ( Y=>nx13858, A0=>modgen_ram_ix74_a_28_dup_538, 
      A1=>nx16197, A2=>nx16573);
   modgen_ram_ix74_ix1538 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_538, 
      QB=>nx13862, D=>nx6889, CLK=>nx15651);
   ix13865 : nor03_2x port map ( Y=>nx13864, A0=>nx7346, A1=>nx7338, A2=>
      nx7330);
   ix7347 : nor03_2x port map ( Y=>nx7346, A0=>nx13867, A1=>nx15439, A2=>
      nx15931);
   modgen_ram_ix74_ix1410 : dff port map ( Q=>OPEN, QB=>nx13867, D=>nx6879, 
      CLK=>nx15651);
   ix7339 : nor03_2x port map ( Y=>nx7338, A0=>nx13871, A1=>nx15779, A2=>
      nx15891);
   modgen_ram_ix74_ix1486 : dff port map ( Q=>OPEN, QB=>nx13871, D=>nx6869, 
      CLK=>nx15651);
   ix7331 : oai22 port map ( Y=>nx7330, A0=>nx13875, A1=>nx16605, B0=>
      nx13878, B1=>nx16621);
   modgen_ram_ix74_ix1478 : dff port map ( Q=>OPEN, QB=>nx13875, D=>nx6859, 
      CLK=>nx15651);
   modgen_ram_ix74_ix1474 : dff port map ( Q=>OPEN, QB=>nx13878, D=>nx6849, 
      CLK=>nx15651);
   ix13882 : nor03_2x port map ( Y=>nx13881, A0=>nx7308, A1=>nx7300, A2=>
      nx7292);
   ix7309 : nor03_2x port map ( Y=>nx7308, A0=>nx13884, A1=>nx15863, A2=>
      nx15917);
   modgen_ram_ix74_ix1598 : dff port map ( Q=>OPEN, QB=>nx13884, D=>nx6839, 
      CLK=>nx15651);
   ix7301 : nor03_2x port map ( Y=>nx7300, A0=>nx13888, A1=>nx15439, A2=>
      nx15903);
   modgen_ram_ix74_ix1414 : dff port map ( Q=>OPEN, QB=>nx13888, D=>nx6829, 
      CLK=>nx15651);
   ix7293 : oai22 port map ( Y=>nx7292, A0=>nx13892, A1=>nx16645, B0=>
      nx13895, B1=>nx16661);
   modgen_ram_ix74_ix1422 : dff port map ( Q=>OPEN, QB=>nx13892, D=>nx6819, 
      CLK=>nx15653);
   modgen_ram_ix74_ix1418 : dff port map ( Q=>OPEN, QB=>nx13895, D=>nx6809, 
      CLK=>nx15653);
   ix7269 : oai22 port map ( Y=>nx7268, A0=>nx13902, A1=>nx16677, B0=>
      nx13905, B1=>nx16693);
   modgen_ram_ix74_ix1566 : dff port map ( Q=>OPEN, QB=>nx13902, D=>nx6789, 
      CLK=>nx15653);
   modgen_ram_ix74_ix1610 : dff port map ( Q=>OPEN, QB=>nx13905, D=>nx6799, 
      CLK=>nx15653);
   ix7251 : oai22 port map ( Y=>nx7250, A0=>nx13909, A1=>nx16709, B0=>
      nx13912, B1=>nx16725);
   modgen_ram_ix74_ix1626 : dff port map ( Q=>OPEN, QB=>nx13909, D=>nx6779, 
      CLK=>nx15653);
   modgen_ram_ix74_ix1562 : dff port map ( Q=>OPEN, QB=>nx13912, D=>nx6769, 
      CLK=>nx15653);
   ix13916 : nor03_2x port map ( Y=>nx13915, A0=>nx7228, A1=>nx7220, A2=>
      nx7212);
   ix7229 : nor03_2x port map ( Y=>nx7228, A0=>nx13918, A1=>nx15439, A2=>
      nx15755);
   modgen_ram_ix74_ix1434 : dff port map ( Q=>OPEN, QB=>nx13918, D=>nx6759, 
      CLK=>nx15653);
   ix7221 : nor03_2x port map ( Y=>nx7220, A0=>nx13922, A1=>nx15863, A2=>
      nx15805);
   modgen_ram_ix74_ix1622 : dff port map ( Q=>OPEN, QB=>nx13922, D=>nx6749, 
      CLK=>nx15655);
   ix7213 : oai22 port map ( Y=>nx7212, A0=>nx13926, A1=>nx16749, B0=>
      nx13929, B1=>nx16757);
   modgen_ram_ix74_ix1430 : dff port map ( Q=>OPEN, QB=>nx13926, D=>nx6739, 
      CLK=>nx15655);
   modgen_ram_ix74_ix1618 : dff port map ( Q=>OPEN, QB=>nx13929, D=>nx6729, 
      CLK=>nx15655);
   ix13933 : nor03_2x port map ( Y=>nx13932, A0=>nx7188, A1=>nx7180, A2=>
      nx7172);
   ix7189 : nor03_2x port map ( Y=>nx7188, A0=>nx13935, A1=>nx15779, A2=>
      nx15815);
   modgen_ram_ix74_ix1490 : dff port map ( Q=>OPEN, QB=>nx13935, D=>nx6719, 
      CLK=>nx15655);
   ix7181 : nor03_2x port map ( Y=>nx7180, A0=>nx13939, A1=>nx15827, A2=>
      nx15805);
   modgen_ram_ix74_ix1558 : dff port map ( Q=>OPEN, QB=>nx13939, D=>nx6709, 
      CLK=>nx15655);
   ix7173 : oai22 port map ( Y=>nx7172, A0=>nx13943, A1=>nx16773, B0=>
      nx13946, B1=>nx16789);
   modgen_ram_ix74_ix1554 : dff port map ( Q=>OPEN, QB=>nx13943, D=>nx6699, 
      CLK=>nx15655);
   modgen_ram_ix74_ix1426 : dff port map ( Q=>OPEN, QB=>nx13946, D=>nx6689, 
      CLK=>nx15655);
   ix13950 : nor03_2x port map ( Y=>nx13949, A0=>nx7150, A1=>nx7142, A2=>
      nx7134);
   ix7151 : nor03_2x port map ( Y=>nx7150, A0=>nx13952, A1=>nx15779, A2=>
      nx15805);
   modgen_ram_ix74_ix1494 : dff port map ( Q=>OPEN, QB=>nx13952, D=>nx6679, 
      CLK=>nx15657);
   ix7143 : nor03_2x port map ( Y=>nx7142, A0=>nx13956, A1=>nx15781, A2=>
      nx15409);
   modgen_ram_ix74_ix1502 : dff port map ( Q=>OPEN, QB=>nx13956, D=>nx6669, 
      CLK=>nx15657);
   ix7135 : oai22 port map ( Y=>nx7134, A0=>nx13960, A1=>nx16821, B0=>
      nx13963, B1=>nx16837);
   modgen_ram_ix74_ix1438 : dff port map ( Q=>OPEN, QB=>nx13960, D=>nx6649, 
      CLK=>nx15657);
   modgen_ram_ix74_ix1498 : dff port map ( Q=>OPEN, QB=>nx13963, D=>nx6659, 
      CLK=>nx15657);
   tri_data_out_11 : tri01 port map ( Y=>data_out(11), A=>nx13967, E=>
      write_out);
   ix8383 : oai22 port map ( Y=>nx8382, A0=>nx13973, A1=>nx16159, B0=>
      nx13978, B1=>nx16185);
   modgen_ram_ix74_ix1185 : dff port map ( Q=>OPEN, QB=>nx13973, D=>nx7919, 
      CLK=>nx15657);
   modgen_ram_ix74_ix1293 : dff port map ( Q=>OPEN, QB=>nx13978, D=>nx7909, 
      CLK=>nx15657);
   ix8365 : oai22 port map ( Y=>nx8364, A0=>nx13982, A1=>nx16203, B0=>
      nx13985, B1=>nx18958);
   modgen_ram_ix74_ix1269 : dff port map ( Q=>OPEN, QB=>nx13982, D=>nx7889, 
      CLK=>nx15657);
   modgen_ram_ix74_ix1277 : dff port map ( Q=>OPEN, QB=>nx13985, D=>nx7899, 
      CLK=>nx15659);
   ix13989 : nor02_2x port map ( Y=>nx13988, A0=>nx8344, A1=>nx8326);
   ix8345 : oai33 port map ( Y=>nx8344, A0=>nx13991, A1=>nx15863, A2=>
      nx16095, B0=>nx13994, B1=>nx15439, B2=>nx16027);
   modgen_ram_ix74_ix1377 : dff port map ( Q=>OPEN, QB=>nx13991, D=>nx7869, 
      CLK=>nx15659);
   modgen_ram_ix74_ix1189 : dff port map ( Q=>OPEN, QB=>nx13994, D=>nx7879, 
      CLK=>nx15659);
   ix8327 : oai22 port map ( Y=>nx8326, A0=>nx13998, A1=>nx16261, B0=>
      nx14001, B1=>nx16277);
   modgen_ram_ix74_ix1313 : dff port map ( Q=>OPEN, QB=>nx13998, D=>nx7859, 
      CLK=>nx15659);
   modgen_ram_ix74_ix1249 : dff port map ( Q=>OPEN, QB=>nx14001, D=>nx7849, 
      CLK=>nx15659);
   ix14005 : nor03_2x port map ( Y=>nx14004, A0=>nx8302, A1=>nx8294, A2=>
      nx8286);
   ix8303 : nor03_2x port map ( Y=>nx8302, A0=>nx14007, A1=>nx15781, A2=>
      nx16069);
   modgen_ram_ix74_ix1205 : dff port map ( Q=>OPEN, QB=>nx14007, D=>nx7839, 
      CLK=>nx15659);
   ix8295 : nor03_2x port map ( Y=>nx8294, A0=>nx14011, A1=>nx15865, A2=>
      nx15409);
   modgen_ram_ix74_ix1373 : dff port map ( Q=>OPEN, QB=>nx14011, D=>nx7829, 
      CLK=>nx15659);
   ix8287 : oai33 port map ( Y=>nx8286, A0=>nx14015, A1=>nx15781, A2=>
      nx15917, B0=>nx14018, B1=>nx15439, B2=>nx16069);
   modgen_ram_ix74_ix1213 : dff port map ( Q=>OPEN, QB=>nx14015, D=>nx7809, 
      CLK=>nx15661);
   modgen_ram_ix74_ix1141 : dff port map ( Q=>OPEN, QB=>nx14018, D=>nx7819, 
      CLK=>nx15661);
   ix14022 : nor03_2x port map ( Y=>nx14021, A0=>nx8264, A1=>nx8256, A2=>
      nx8248);
   ix8265 : nor03_2x port map ( Y=>nx8264, A0=>nx14024, A1=>nx15781, A2=>
      nx16047);
   modgen_ram_ix74_ix1209 : dff port map ( Q=>OPEN, QB=>nx14024, D=>nx7799, 
      CLK=>nx15661);
   ix8257 : nor04 port map ( Y=>nx8256, A0=>nx14028, A1=>address(4), A2=>
      address(5), A3=>nx16071);
   modgen_ram_ix74_ix1333 : dff port map ( Q=>OPEN, QB=>nx14028, D=>nx7789, 
      CLK=>nx15661);
   ix8249 : oai22 port map ( Y=>nx8248, A0=>nx14032, A1=>nx16329, B0=>
      nx14035, B1=>nx16345);
   modgen_ram_ix74_ix1149 : dff port map ( Q=>OPEN, QB=>nx14032, D=>nx7769, 
      CLK=>nx15661);
   modgen_ram_ix74_ix1145 : dff port map ( Q=>OPEN, QB=>nx14035, D=>nx7779, 
      CLK=>nx15661);
   modgen_ram_ix74_ix1273 : dff port map ( Q=>OPEN, QB=>nx14042, D=>nx7759, 
      CLK=>nx15661);
   modgen_ram_ix74_ix1337 : dff port map ( Q=>OPEN, QB=>nx14046, D=>nx7749, 
      CLK=>nx15663);
   ix8207 : oai22 port map ( Y=>nx8206, A0=>nx14050, A1=>nx16361, B0=>
      nx14053, B1=>nx16377);
   modgen_ram_ix74_ix1317 : dff port map ( Q=>OPEN, QB=>nx14050, D=>nx7729, 
      CLK=>nx15663);
   modgen_ram_ix74_ix1253 : dff port map ( Q=>OPEN, QB=>nx14053, D=>nx7739, 
      CLK=>nx15663);
   modgen_ram_ix74_ix1381 : dff port map ( Q=>OPEN, QB=>nx14059, D=>nx7719, 
      CLK=>nx15663);
   modgen_ram_ix74_ix1193 : dff port map ( Q=>OPEN, QB=>nx14063, D=>nx7709, 
      CLK=>nx15663);
   ix8169 : oai22 port map ( Y=>nx8168, A0=>nx14067, A1=>nx16401, B0=>
      nx14070, B1=>nx16417);
   modgen_ram_ix74_ix1321 : dff port map ( Q=>OPEN, QB=>nx14067, D=>nx7689, 
      CLK=>nx15663);
   modgen_ram_ix74_ix1257 : dff port map ( Q=>OPEN, QB=>nx14070, D=>nx7699, 
      CLK=>nx15663);
   modgen_ram_ix74_ix1385 : dff port map ( Q=>OPEN, QB=>nx14076, D=>nx7679, 
      CLK=>nx15665);
   modgen_ram_ix74_ix1197 : dff port map ( Q=>OPEN, QB=>nx14080, D=>nx7669, 
      CLK=>nx15665);
   ix8129 : oai22 port map ( Y=>nx8128, A0=>nx14084, A1=>nx16441, B0=>
      nx14087, B1=>nx16457);
   modgen_ram_ix74_ix1325 : dff port map ( Q=>OPEN, QB=>nx14084, D=>nx7649, 
      CLK=>nx15665);
   modgen_ram_ix74_ix1261 : dff port map ( Q=>OPEN, QB=>nx14087, D=>nx7659, 
      CLK=>nx15665);
   modgen_ram_ix74_ix1389 : dff port map ( Q=>OPEN, QB=>nx14093, D=>nx7639, 
      CLK=>nx15665);
   ix8099 : nor03_2x port map ( Y=>nx8098, A0=>nx14097, A1=>nx15441, A2=>
      nx15961);
   modgen_ram_ix74_ix1201 : dff port map ( Q=>OPEN, QB=>nx14097, D=>nx7629, 
      CLK=>nx15665);
   ix8091 : oai22 port map ( Y=>nx8090, A0=>nx14101, A1=>nx16481, B0=>
      nx14104, B1=>nx16497);
   modgen_ram_ix74_ix1329 : dff port map ( Q=>OPEN, QB=>nx14101, D=>nx7609, 
      CLK=>nx15665);
   modgen_ram_ix74_ix1265 : dff port map ( Q=>OPEN, QB=>nx14104, D=>nx7619, 
      CLK=>nx15667);
   ix8065 : oai22 port map ( Y=>nx8064, A0=>nx14114, A1=>nx16513, B0=>
      nx14117, B1=>nx16521);
   modgen_ram_ix74_ix1357 : dff port map ( Q=>OPEN, QB=>nx14114, D=>nx7589, 
      CLK=>nx15667);
   modgen_ram_ix74_ix1393 : dff port map ( Q=>OPEN, QB=>nx14117, D=>nx7599, 
      CLK=>nx15667);
   ix8047 : oai22 port map ( Y=>nx8046, A0=>nx14121, A1=>nx16529, B0=>
      nx14124, B1=>nx16545);
   modgen_ram_ix74_ix1289 : dff port map ( Q=>OPEN, QB=>nx14121, D=>nx7579, 
      CLK=>nx15667);
   modgen_ram_ix74_ix1225 : dff port map ( Q=>OPEN, QB=>nx14124, D=>nx7569, 
      CLK=>nx15667);
   ix8029 : nand03 port map ( Y=>nx8028, A0=>nx14128, A1=>nx14138, A2=>
      nx14144);
   ix14129 : nor02_2x port map ( Y=>nx14128, A0=>nx8024, A1=>nx8016);
   ix8025 : nor04 port map ( Y=>nx8024, A0=>nx14131, A1=>address(4), A2=>
      address(5), A3=>nx15903);
   modgen_ram_ix74_ix1349 : dff port map ( Q=>OPEN, QB=>nx14131, D=>nx7559, 
      CLK=>nx15667);
   ix8017 : nor03_2x port map ( Y=>nx8016, A0=>nx14135, A1=>nx15827, A2=>
      nx15905);
   modgen_ram_ix74_ix1285 : dff port map ( Q=>OPEN, QB=>nx14135, D=>nx7549, 
      CLK=>nx15667);
   ix14139 : nand03 port map ( Y=>nx14138, A0=>modgen_ram_ix74_a_12_dup_489, 
      A1=>nx16233, A2=>nx16573);
   modgen_ram_ix74_ix1345 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_489, 
      QB=>nx14142, D=>nx7539, CLK=>nx15669);
   ix14145 : nand03 port map ( Y=>nx14144, A0=>modgen_ram_ix74_a_28_dup_473, 
      A1=>nx16197, A2=>nx16573);
   modgen_ram_ix74_ix1281 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_473, 
      QB=>nx14148, D=>nx7529, CLK=>nx15669);
   ix14151 : nor03_2x port map ( Y=>nx14150, A0=>nx7984, A1=>nx7976, A2=>
      nx7968);
   ix7985 : nor03_2x port map ( Y=>nx7984, A0=>nx14153, A1=>nx15441, A2=>
      nx15931);
   modgen_ram_ix74_ix1153 : dff port map ( Q=>OPEN, QB=>nx14153, D=>nx7519, 
      CLK=>nx15669);
   ix7977 : nor03_2x port map ( Y=>nx7976, A0=>nx14157, A1=>nx15781, A2=>
      nx15891);
   modgen_ram_ix74_ix1229 : dff port map ( Q=>OPEN, QB=>nx14157, D=>nx7509, 
      CLK=>nx15669);
   ix7969 : oai22 port map ( Y=>nx7968, A0=>nx14161, A1=>nx16605, B0=>
      nx14164, B1=>nx16621);
   modgen_ram_ix74_ix1221 : dff port map ( Q=>OPEN, QB=>nx14161, D=>nx7499, 
      CLK=>nx15669);
   modgen_ram_ix74_ix1217 : dff port map ( Q=>OPEN, QB=>nx14164, D=>nx7489, 
      CLK=>nx15669);
   ix14168 : nor03_2x port map ( Y=>nx14167, A0=>nx7946, A1=>nx7938, A2=>
      nx7930);
   ix7947 : nor03_2x port map ( Y=>nx7946, A0=>nx14170, A1=>nx15865, A2=>
      nx15917);
   modgen_ram_ix74_ix1341 : dff port map ( Q=>OPEN, QB=>nx14170, D=>nx7479, 
      CLK=>nx15669);
   ix7939 : nor03_2x port map ( Y=>nx7938, A0=>nx14174, A1=>nx15441, A2=>
      nx15905);
   modgen_ram_ix74_ix1157 : dff port map ( Q=>OPEN, QB=>nx14174, D=>nx7469, 
      CLK=>nx15671);
   ix7931 : oai22 port map ( Y=>nx7930, A0=>nx14178, A1=>nx16645, B0=>
      nx14181, B1=>nx16661);
   modgen_ram_ix74_ix1165 : dff port map ( Q=>OPEN, QB=>nx14178, D=>nx7459, 
      CLK=>nx15671);
   modgen_ram_ix74_ix1161 : dff port map ( Q=>OPEN, QB=>nx14181, D=>nx7449, 
      CLK=>nx15671);
   ix7907 : oai22 port map ( Y=>nx7906, A0=>nx14188, A1=>nx16677, B0=>
      nx14191, B1=>nx16693);
   modgen_ram_ix74_ix1309 : dff port map ( Q=>OPEN, QB=>nx14188, D=>nx7429, 
      CLK=>nx15671);
   modgen_ram_ix74_ix1353 : dff port map ( Q=>OPEN, QB=>nx14191, D=>nx7439, 
      CLK=>nx15671);
   ix7889 : oai22 port map ( Y=>nx7888, A0=>nx14195, A1=>nx16709, B0=>
      nx14198, B1=>nx16725);
   modgen_ram_ix74_ix1369 : dff port map ( Q=>OPEN, QB=>nx14195, D=>nx7419, 
      CLK=>nx15671);
   modgen_ram_ix74_ix1305 : dff port map ( Q=>OPEN, QB=>nx14198, D=>nx7409, 
      CLK=>nx15671);
   ix14202 : nor03_2x port map ( Y=>nx14201, A0=>nx7866, A1=>nx7858, A2=>
      nx7850);
   ix7867 : nor03_2x port map ( Y=>nx7866, A0=>nx14204, A1=>nx15441, A2=>
      nx15755);
   modgen_ram_ix74_ix1177 : dff port map ( Q=>OPEN, QB=>nx14204, D=>nx7399, 
      CLK=>nx15673);
   ix7859 : nor03_2x port map ( Y=>nx7858, A0=>nx14208, A1=>nx15865, A2=>
      nx15807);
   modgen_ram_ix74_ix1365 : dff port map ( Q=>OPEN, QB=>nx14208, D=>nx7389, 
      CLK=>nx15673);
   ix7851 : oai22 port map ( Y=>nx7850, A0=>nx14212, A1=>nx16749, B0=>
      nx14215, B1=>nx16757);
   modgen_ram_ix74_ix1173 : dff port map ( Q=>OPEN, QB=>nx14212, D=>nx7379, 
      CLK=>nx15673);
   modgen_ram_ix74_ix1361 : dff port map ( Q=>OPEN, QB=>nx14215, D=>nx7369, 
      CLK=>nx15673);
   ix14219 : nor03_2x port map ( Y=>nx14218, A0=>nx7826, A1=>nx7818, A2=>
      nx7810);
   ix7827 : nor03_2x port map ( Y=>nx7826, A0=>nx14221, A1=>nx15781, A2=>
      nx15815);
   modgen_ram_ix74_ix1233 : dff port map ( Q=>OPEN, QB=>nx14221, D=>nx7359, 
      CLK=>nx15673);
   ix7819 : nor03_2x port map ( Y=>nx7818, A0=>nx14225, A1=>nx15829, A2=>
      nx15807);
   modgen_ram_ix74_ix1301 : dff port map ( Q=>OPEN, QB=>nx14225, D=>nx7349, 
      CLK=>nx15673);
   ix7811 : oai22 port map ( Y=>nx7810, A0=>nx14229, A1=>nx16773, B0=>
      nx14232, B1=>nx16789);
   modgen_ram_ix74_ix1297 : dff port map ( Q=>OPEN, QB=>nx14229, D=>nx7339, 
      CLK=>nx15673);
   modgen_ram_ix74_ix1169 : dff port map ( Q=>OPEN, QB=>nx14232, D=>nx7329, 
      CLK=>nx15675);
   ix14236 : nor03_2x port map ( Y=>nx14235, A0=>nx7788, A1=>nx7780, A2=>
      nx7772);
   ix7789 : nor03_2x port map ( Y=>nx7788, A0=>nx14238, A1=>nx15781, A2=>
      nx15807);
   modgen_ram_ix74_ix1237 : dff port map ( Q=>OPEN, QB=>nx14238, D=>nx7319, 
      CLK=>nx15675);
   ix7781 : nor03_2x port map ( Y=>nx7780, A0=>nx14242, A1=>nx15783, A2=>
      nx15409);
   modgen_ram_ix74_ix1245 : dff port map ( Q=>OPEN, QB=>nx14242, D=>nx7309, 
      CLK=>nx15675);
   ix7773 : oai22 port map ( Y=>nx7772, A0=>nx14246, A1=>nx16821, B0=>
      nx14249, B1=>nx16837);
   modgen_ram_ix74_ix1181 : dff port map ( Q=>OPEN, QB=>nx14246, D=>nx7289, 
      CLK=>nx15675);
   modgen_ram_ix74_ix1241 : dff port map ( Q=>OPEN, QB=>nx14249, D=>nx7299, 
      CLK=>nx15675);
   tri_data_out_12 : tri01 port map ( Y=>data_out(12), A=>nx14253, E=>
      write_out);
   ix9021 : oai22 port map ( Y=>nx9020, A0=>nx14259, A1=>nx16159, B0=>
      nx14264, B1=>nx16185);
   modgen_ram_ix74_ix928 : dff port map ( Q=>OPEN, QB=>nx14259, D=>nx8559, 
      CLK=>nx15675);
   modgen_ram_ix74_ix1036 : dff port map ( Q=>OPEN, QB=>nx14264, D=>nx8549, 
      CLK=>nx15675);
   ix9003 : oai22 port map ( Y=>nx9002, A0=>nx14268, A1=>nx16203, B0=>
      nx14271, B1=>nx18958);
   modgen_ram_ix74_ix1012 : dff port map ( Q=>OPEN, QB=>nx14268, D=>nx8529, 
      CLK=>nx15677);
   modgen_ram_ix74_ix1020 : dff port map ( Q=>OPEN, QB=>nx14271, D=>nx8539, 
      CLK=>nx15677);
   ix14275 : nor02_2x port map ( Y=>nx14274, A0=>nx8982, A1=>nx8964);
   ix8983 : oai33 port map ( Y=>nx8982, A0=>nx14277, A1=>nx15865, A2=>
      nx16095, B0=>nx14280, B1=>nx15441, B2=>nx16027);
   modgen_ram_ix74_ix1120 : dff port map ( Q=>OPEN, QB=>nx14277, D=>nx8509, 
      CLK=>nx15677);
   modgen_ram_ix74_ix932 : dff port map ( Q=>OPEN, QB=>nx14280, D=>nx8519, 
      CLK=>nx15677);
   ix8965 : oai22 port map ( Y=>nx8964, A0=>nx14284, A1=>nx16261, B0=>
      nx14287, B1=>nx16277);
   modgen_ram_ix74_ix1056 : dff port map ( Q=>OPEN, QB=>nx14284, D=>nx8499, 
      CLK=>nx15677);
   modgen_ram_ix74_ix992 : dff port map ( Q=>OPEN, QB=>nx14287, D=>nx8489, 
      CLK=>nx15677);
   ix14291 : nor03_2x port map ( Y=>nx14290, A0=>nx8940, A1=>nx8932, A2=>
      nx8924);
   ix8941 : nor03_2x port map ( Y=>nx8940, A0=>nx14293, A1=>nx15783, A2=>
      nx16071);
   modgen_ram_ix74_ix948 : dff port map ( Q=>OPEN, QB=>nx14293, D=>nx8479, 
      CLK=>nx15677);
   ix8933 : nor03_2x port map ( Y=>nx8932, A0=>nx14297, A1=>nx15865, A2=>
      nx15411);
   modgen_ram_ix74_ix1116 : dff port map ( Q=>OPEN, QB=>nx14297, D=>nx8469, 
      CLK=>nx15679);
   ix8925 : oai33 port map ( Y=>nx8924, A0=>nx14301, A1=>nx15783, A2=>
      nx15917, B0=>nx14304, B1=>nx15443, B2=>nx16071);
   modgen_ram_ix74_ix956 : dff port map ( Q=>OPEN, QB=>nx14301, D=>nx8449, 
      CLK=>nx15679);
   modgen_ram_ix74_ix884 : dff port map ( Q=>OPEN, QB=>nx14304, D=>nx8459, 
      CLK=>nx15679);
   ix14308 : nor03_2x port map ( Y=>nx14307, A0=>nx8902, A1=>nx8894, A2=>
      nx8886);
   ix8903 : nor03_2x port map ( Y=>nx8902, A0=>nx14310, A1=>nx15783, A2=>
      nx16049);
   modgen_ram_ix74_ix952 : dff port map ( Q=>OPEN, QB=>nx14310, D=>nx8439, 
      CLK=>nx15679);
   ix8895 : nor04 port map ( Y=>nx8894, A0=>nx14314, A1=>address(4), A2=>
      address(5), A3=>nx16071);
   modgen_ram_ix74_ix1076 : dff port map ( Q=>OPEN, QB=>nx14314, D=>nx8429, 
      CLK=>nx15679);
   ix8887 : oai22 port map ( Y=>nx8886, A0=>nx14318, A1=>nx16329, B0=>
      nx14321, B1=>nx16345);
   modgen_ram_ix74_ix892 : dff port map ( Q=>OPEN, QB=>nx14318, D=>nx8409, 
      CLK=>nx15679);
   modgen_ram_ix74_ix888 : dff port map ( Q=>OPEN, QB=>nx14321, D=>nx8419, 
      CLK=>nx15679);
   modgen_ram_ix74_ix1016 : dff port map ( Q=>OPEN, QB=>nx14328, D=>nx8399, 
      CLK=>nx15681);
   modgen_ram_ix74_ix1080 : dff port map ( Q=>OPEN, QB=>nx14332, D=>nx8389, 
      CLK=>nx15681);
   ix8845 : oai22 port map ( Y=>nx8844, A0=>nx14336, A1=>nx16361, B0=>
      nx14339, B1=>nx16377);
   modgen_ram_ix74_ix1060 : dff port map ( Q=>OPEN, QB=>nx14336, D=>nx8369, 
      CLK=>nx15681);
   modgen_ram_ix74_ix996 : dff port map ( Q=>OPEN, QB=>nx14339, D=>nx8379, 
      CLK=>nx15681);
   modgen_ram_ix74_ix1124 : dff port map ( Q=>OPEN, QB=>nx14345, D=>nx8359, 
      CLK=>nx15681);
   modgen_ram_ix74_ix936 : dff port map ( Q=>OPEN, QB=>nx14349, D=>nx8349, 
      CLK=>nx15681);
   ix8807 : oai22 port map ( Y=>nx8806, A0=>nx14353, A1=>nx16401, B0=>
      nx14356, B1=>nx16417);
   modgen_ram_ix74_ix1064 : dff port map ( Q=>OPEN, QB=>nx14353, D=>nx8329, 
      CLK=>nx15681);
   modgen_ram_ix74_ix1000 : dff port map ( Q=>OPEN, QB=>nx14356, D=>nx8339, 
      CLK=>nx15683);
   modgen_ram_ix74_ix1128 : dff port map ( Q=>OPEN, QB=>nx14362, D=>nx8319, 
      CLK=>nx15683);
   modgen_ram_ix74_ix940 : dff port map ( Q=>OPEN, QB=>nx14366, D=>nx8309, 
      CLK=>nx15683);
   ix8767 : oai22 port map ( Y=>nx8766, A0=>nx14370, A1=>nx16441, B0=>
      nx14373, B1=>nx16457);
   modgen_ram_ix74_ix1068 : dff port map ( Q=>OPEN, QB=>nx14370, D=>nx8289, 
      CLK=>nx15683);
   modgen_ram_ix74_ix1004 : dff port map ( Q=>OPEN, QB=>nx14373, D=>nx8299, 
      CLK=>nx15683);
   modgen_ram_ix74_ix1132 : dff port map ( Q=>OPEN, QB=>nx14379, D=>nx8279, 
      CLK=>nx15683);
   ix8737 : nor03_2x port map ( Y=>nx8736, A0=>nx14383, A1=>nx15443, A2=>
      nx15963);
   modgen_ram_ix74_ix944 : dff port map ( Q=>OPEN, QB=>nx14383, D=>nx8269, 
      CLK=>nx15683);
   ix8729 : oai22 port map ( Y=>nx8728, A0=>nx14387, A1=>nx16481, B0=>
      nx14390, B1=>nx16497);
   modgen_ram_ix74_ix1072 : dff port map ( Q=>OPEN, QB=>nx14387, D=>nx8249, 
      CLK=>nx15685);
   modgen_ram_ix74_ix1008 : dff port map ( Q=>OPEN, QB=>nx14390, D=>nx8259, 
      CLK=>nx15685);
   ix8703 : oai22 port map ( Y=>nx8702, A0=>nx14400, A1=>nx16513, B0=>
      nx14403, B1=>nx16521);
   modgen_ram_ix74_ix1100 : dff port map ( Q=>OPEN, QB=>nx14400, D=>nx8229, 
      CLK=>nx15685);
   modgen_ram_ix74_ix1136 : dff port map ( Q=>OPEN, QB=>nx14403, D=>nx8239, 
      CLK=>nx15685);
   ix8685 : oai22 port map ( Y=>nx8684, A0=>nx14407, A1=>nx16529, B0=>
      nx14410, B1=>nx16545);
   modgen_ram_ix74_ix1032 : dff port map ( Q=>OPEN, QB=>nx14407, D=>nx8219, 
      CLK=>nx15685);
   modgen_ram_ix74_ix968 : dff port map ( Q=>OPEN, QB=>nx14410, D=>nx8209, 
      CLK=>nx15685);
   ix8667 : nand03 port map ( Y=>nx8666, A0=>nx14414, A1=>nx14424, A2=>
      nx14430);
   ix14415 : nor02_2x port map ( Y=>nx14414, A0=>nx8662, A1=>nx8654);
   ix8663 : nor04 port map ( Y=>nx8662, A0=>nx14417, A1=>address(4), A2=>
      address(5), A3=>nx15905);
   modgen_ram_ix74_ix1092 : dff port map ( Q=>OPEN, QB=>nx14417, D=>nx8199, 
      CLK=>nx15685);
   ix8655 : nor03_2x port map ( Y=>nx8654, A0=>nx14421, A1=>nx15829, A2=>
      nx15905);
   modgen_ram_ix74_ix1028 : dff port map ( Q=>OPEN, QB=>nx14421, D=>nx8189, 
      CLK=>nx15687);
   ix14425 : nand03 port map ( Y=>nx14424, A0=>modgen_ram_ix74_a_12_dup_424, 
      A1=>nx16233, A2=>nx16573);
   modgen_ram_ix74_ix1088 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_424, 
      QB=>nx14428, D=>nx8179, CLK=>nx15687);
   ix14431 : nand03 port map ( Y=>nx14430, A0=>modgen_ram_ix74_a_28_dup_408, 
      A1=>nx16197, A2=>nx16575);
   modgen_ram_ix74_ix1024 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_408, 
      QB=>nx14434, D=>nx8169, CLK=>nx15687);
   ix14437 : nor03_2x port map ( Y=>nx14436, A0=>nx8622, A1=>nx8614, A2=>
      nx8606);
   ix8623 : nor03_2x port map ( Y=>nx8622, A0=>nx14439, A1=>nx15443, A2=>
      nx15931);
   modgen_ram_ix74_ix896 : dff port map ( Q=>OPEN, QB=>nx14439, D=>nx8159, 
      CLK=>nx15687);
   ix8615 : nor03_2x port map ( Y=>nx8614, A0=>nx14443, A1=>nx15783, A2=>
      nx15891);
   modgen_ram_ix74_ix972 : dff port map ( Q=>OPEN, QB=>nx14443, D=>nx8149, 
      CLK=>nx15687);
   ix8607 : oai22 port map ( Y=>nx8606, A0=>nx14447, A1=>nx16605, B0=>
      nx14450, B1=>nx16621);
   modgen_ram_ix74_ix964 : dff port map ( Q=>OPEN, QB=>nx14447, D=>nx8139, 
      CLK=>nx15687);
   modgen_ram_ix74_ix960 : dff port map ( Q=>OPEN, QB=>nx14450, D=>nx8129, 
      CLK=>nx15687);
   ix14454 : nor03_2x port map ( Y=>nx14453, A0=>nx8584, A1=>nx8576, A2=>
      nx8568);
   ix8585 : nor03_2x port map ( Y=>nx8584, A0=>nx14456, A1=>nx15867, A2=>
      nx15917);
   modgen_ram_ix74_ix1084 : dff port map ( Q=>OPEN, QB=>nx14456, D=>nx8119, 
      CLK=>nx15689);
   ix8577 : nor03_2x port map ( Y=>nx8576, A0=>nx14460, A1=>nx15443, A2=>
      nx15905);
   modgen_ram_ix74_ix900 : dff port map ( Q=>OPEN, QB=>nx14460, D=>nx8109, 
      CLK=>nx15689);
   ix8569 : oai22 port map ( Y=>nx8568, A0=>nx14464, A1=>nx16645, B0=>
      nx14467, B1=>nx16661);
   modgen_ram_ix74_ix908 : dff port map ( Q=>OPEN, QB=>nx14464, D=>nx8099, 
      CLK=>nx15689);
   modgen_ram_ix74_ix904 : dff port map ( Q=>OPEN, QB=>nx14467, D=>nx8089, 
      CLK=>nx15689);
   ix8545 : oai22 port map ( Y=>nx8544, A0=>nx14474, A1=>nx16677, B0=>
      nx14477, B1=>nx16693);
   modgen_ram_ix74_ix1052 : dff port map ( Q=>OPEN, QB=>nx14474, D=>nx8069, 
      CLK=>nx15689);
   modgen_ram_ix74_ix1096 : dff port map ( Q=>OPEN, QB=>nx14477, D=>nx8079, 
      CLK=>nx15689);
   ix8527 : oai22 port map ( Y=>nx8526, A0=>nx14481, A1=>nx16709, B0=>
      nx14484, B1=>nx16725);
   modgen_ram_ix74_ix1112 : dff port map ( Q=>OPEN, QB=>nx14481, D=>nx8059, 
      CLK=>nx15689);
   modgen_ram_ix74_ix1048 : dff port map ( Q=>OPEN, QB=>nx14484, D=>nx8049, 
      CLK=>nx15691);
   ix14488 : nor03_2x port map ( Y=>nx14487, A0=>nx8504, A1=>nx8496, A2=>
      nx8488);
   ix8505 : nor03_2x port map ( Y=>nx8504, A0=>nx14490, A1=>nx15443, A2=>
      nx15757);
   modgen_ram_ix74_ix920 : dff port map ( Q=>OPEN, QB=>nx14490, D=>nx8039, 
      CLK=>nx15691);
   ix8497 : nor03_2x port map ( Y=>nx8496, A0=>nx14494, A1=>nx15867, A2=>
      nx15807);
   modgen_ram_ix74_ix1108 : dff port map ( Q=>OPEN, QB=>nx14494, D=>nx8029, 
      CLK=>nx15691);
   ix8489 : oai22 port map ( Y=>nx8488, A0=>nx14498, A1=>nx16749, B0=>
      nx14501, B1=>nx16757);
   modgen_ram_ix74_ix916 : dff port map ( Q=>OPEN, QB=>nx14498, D=>nx8019, 
      CLK=>nx15691);
   modgen_ram_ix74_ix1104 : dff port map ( Q=>OPEN, QB=>nx14501, D=>nx8009, 
      CLK=>nx15691);
   ix14505 : nor03_2x port map ( Y=>nx14504, A0=>nx8464, A1=>nx8456, A2=>
      nx8448);
   ix8465 : nor03_2x port map ( Y=>nx8464, A0=>nx14507, A1=>nx15783, A2=>
      nx15817);
   modgen_ram_ix74_ix976 : dff port map ( Q=>OPEN, QB=>nx14507, D=>nx7999, 
      CLK=>nx15691);
   ix8457 : nor03_2x port map ( Y=>nx8456, A0=>nx14511, A1=>nx15829, A2=>
      nx15807);
   modgen_ram_ix74_ix1044 : dff port map ( Q=>OPEN, QB=>nx14511, D=>nx7989, 
      CLK=>nx15691);
   ix8449 : oai22 port map ( Y=>nx8448, A0=>nx14515, A1=>nx16773, B0=>
      nx14518, B1=>nx16789);
   modgen_ram_ix74_ix1040 : dff port map ( Q=>OPEN, QB=>nx14515, D=>nx7979, 
      CLK=>nx15693);
   modgen_ram_ix74_ix912 : dff port map ( Q=>OPEN, QB=>nx14518, D=>nx7969, 
      CLK=>nx15693);
   ix14522 : nor03_2x port map ( Y=>nx14521, A0=>nx8426, A1=>nx8418, A2=>
      nx8410);
   ix8427 : nor03_2x port map ( Y=>nx8426, A0=>nx14524, A1=>nx15783, A2=>
      nx15807);
   modgen_ram_ix74_ix980 : dff port map ( Q=>OPEN, QB=>nx14524, D=>nx7959, 
      CLK=>nx15693);
   ix8419 : nor03_2x port map ( Y=>nx8418, A0=>nx14528, A1=>nx15785, A2=>
      nx15411);
   modgen_ram_ix74_ix988 : dff port map ( Q=>OPEN, QB=>nx14528, D=>nx7949, 
      CLK=>nx15693);
   ix8411 : oai22 port map ( Y=>nx8410, A0=>nx14532, A1=>nx16821, B0=>
      nx14535, B1=>nx16837);
   modgen_ram_ix74_ix924 : dff port map ( Q=>OPEN, QB=>nx14532, D=>nx7929, 
      CLK=>nx15693);
   modgen_ram_ix74_ix984 : dff port map ( Q=>OPEN, QB=>nx14535, D=>nx7939, 
      CLK=>nx15693);
   tri_data_out_13 : tri01 port map ( Y=>data_out(13), A=>nx14539, E=>
      write_out);
   ix9659 : oai22 port map ( Y=>nx9658, A0=>nx14545, A1=>nx16159, B0=>
      nx14550, B1=>nx16185);
   modgen_ram_ix74_ix671 : dff port map ( Q=>OPEN, QB=>nx14545, D=>nx9199, 
      CLK=>nx15693);
   modgen_ram_ix74_ix779 : dff port map ( Q=>OPEN, QB=>nx14550, D=>nx9189, 
      CLK=>nx15695);
   modgen_ram_ix74_ix755 : dff port map ( Q=>OPEN, QB=>nx14554, D=>nx9169, 
      CLK=>nx15695);
   modgen_ram_ix74_ix763 : dff port map ( Q=>OPEN, QB=>nx14557, D=>nx9179, 
      CLK=>nx15695);
   ix14561 : nor02_2x port map ( Y=>nx14560, A0=>nx9620, A1=>nx9602);
   ix9621 : oai33 port map ( Y=>nx9620, A0=>nx14563, A1=>nx15867, A2=>
      nx16095, B0=>nx14566, B1=>nx15445, B2=>nx16027);
   modgen_ram_ix74_ix863 : dff port map ( Q=>OPEN, QB=>nx14563, D=>nx9149, 
      CLK=>nx15695);
   modgen_ram_ix74_ix675 : dff port map ( Q=>OPEN, QB=>nx14566, D=>nx9159, 
      CLK=>nx15695);
   ix9603 : oai22 port map ( Y=>nx9602, A0=>nx14570, A1=>nx16261, B0=>
      nx14573, B1=>nx16277);
   modgen_ram_ix74_ix799 : dff port map ( Q=>OPEN, QB=>nx14570, D=>nx9139, 
      CLK=>nx15695);
   modgen_ram_ix74_ix735 : dff port map ( Q=>OPEN, QB=>nx14573, D=>nx9129, 
      CLK=>nx15695);
   ix14577 : nor03_2x port map ( Y=>nx14576, A0=>nx9578, A1=>nx9570, A2=>
      nx9562);
   ix9579 : nor03_2x port map ( Y=>nx9578, A0=>nx14579, A1=>nx15785, A2=>
      nx16071);
   modgen_ram_ix74_ix691 : dff port map ( Q=>OPEN, QB=>nx14579, D=>nx9119, 
      CLK=>nx15697);
   ix9571 : nor03_2x port map ( Y=>nx9570, A0=>nx14583, A1=>nx15867, A2=>
      nx15411);
   modgen_ram_ix74_ix859 : dff port map ( Q=>OPEN, QB=>nx14583, D=>nx9109, 
      CLK=>nx15697);
   ix9563 : oai33 port map ( Y=>nx9562, A0=>nx14587, A1=>nx15785, A2=>
      nx15919, B0=>nx14590, B1=>nx15445, B2=>nx16071);
   modgen_ram_ix74_ix699 : dff port map ( Q=>OPEN, QB=>nx14587, D=>nx9089, 
      CLK=>nx15697);
   modgen_ram_ix74_ix627 : dff port map ( Q=>OPEN, QB=>nx14590, D=>nx9099, 
      CLK=>nx15697);
   ix14594 : nor03_2x port map ( Y=>nx14593, A0=>nx9540, A1=>nx9532, A2=>
      nx9524);
   ix9541 : nor03_2x port map ( Y=>nx9540, A0=>nx14596, A1=>nx15785, A2=>
      nx16049);
   modgen_ram_ix74_ix695 : dff port map ( Q=>OPEN, QB=>nx14596, D=>nx9079, 
      CLK=>nx15697);
   ix9533 : nor04 port map ( Y=>nx9532, A0=>nx14600, A1=>address(4), A2=>
      address(5), A3=>nx16071);
   modgen_ram_ix74_ix819 : dff port map ( Q=>OPEN, QB=>nx14600, D=>nx9069, 
      CLK=>nx15697);
   ix9525 : oai22 port map ( Y=>nx9524, A0=>nx14604, A1=>nx16329, B0=>
      nx14607, B1=>nx16345);
   modgen_ram_ix74_ix635 : dff port map ( Q=>OPEN, QB=>nx14604, D=>nx9049, 
      CLK=>nx15697);
   modgen_ram_ix74_ix631 : dff port map ( Q=>OPEN, QB=>nx14607, D=>nx9059, 
      CLK=>nx15699);
   modgen_ram_ix74_ix759 : dff port map ( Q=>OPEN, QB=>nx14614, D=>nx9039, 
      CLK=>nx15699);
   modgen_ram_ix74_ix823 : dff port map ( Q=>OPEN, QB=>nx14618, D=>nx9029, 
      CLK=>nx15699);
   ix9483 : oai22 port map ( Y=>nx9482, A0=>nx14622, A1=>nx16361, B0=>
      nx14625, B1=>nx16377);
   modgen_ram_ix74_ix803 : dff port map ( Q=>OPEN, QB=>nx14622, D=>nx9009, 
      CLK=>nx15699);
   modgen_ram_ix74_ix739 : dff port map ( Q=>OPEN, QB=>nx14625, D=>nx9019, 
      CLK=>nx15699);
   modgen_ram_ix74_ix867 : dff port map ( Q=>OPEN, QB=>nx14631, D=>nx8999, 
      CLK=>nx15699);
   modgen_ram_ix74_ix679 : dff port map ( Q=>OPEN, QB=>nx14635, D=>nx8989, 
      CLK=>nx15699);
   ix9445 : oai22 port map ( Y=>nx9444, A0=>nx14639, A1=>nx16401, B0=>
      nx14642, B1=>nx16417);
   modgen_ram_ix74_ix807 : dff port map ( Q=>OPEN, QB=>nx14639, D=>nx8969, 
      CLK=>nx15701);
   modgen_ram_ix74_ix743 : dff port map ( Q=>OPEN, QB=>nx14642, D=>nx8979, 
      CLK=>nx15701);
   modgen_ram_ix74_ix871 : dff port map ( Q=>OPEN, QB=>nx14648, D=>nx8959, 
      CLK=>nx15701);
   modgen_ram_ix74_ix683 : dff port map ( Q=>OPEN, QB=>nx14652, D=>nx8949, 
      CLK=>nx15701);
   modgen_ram_ix74_ix811 : dff port map ( Q=>OPEN, QB=>nx14656, D=>nx8929, 
      CLK=>nx15701);
   modgen_ram_ix74_ix747 : dff port map ( Q=>OPEN, QB=>nx14659, D=>nx8939, 
      CLK=>nx15701);
   modgen_ram_ix74_ix875 : dff port map ( Q=>OPEN, QB=>nx14665, D=>nx8919, 
      CLK=>nx15701);
   ix9375 : nor03_2x port map ( Y=>nx9374, A0=>nx14669, A1=>nx15445, A2=>
      nx15963);
   modgen_ram_ix74_ix687 : dff port map ( Q=>OPEN, QB=>nx14669, D=>nx8909, 
      CLK=>nx15703);
   modgen_ram_ix74_ix815 : dff port map ( Q=>OPEN, QB=>nx14673, D=>nx8889, 
      CLK=>nx15703);
   modgen_ram_ix74_ix751 : dff port map ( Q=>OPEN, QB=>nx14676, D=>nx8899, 
      CLK=>nx15703);
   ix9341 : oai22 port map ( Y=>nx9340, A0=>nx14686, A1=>nx16513, B0=>
      nx14689, B1=>nx16521);
   modgen_ram_ix74_ix843 : dff port map ( Q=>OPEN, QB=>nx14686, D=>nx8869, 
      CLK=>nx15703);
   modgen_ram_ix74_ix879 : dff port map ( Q=>OPEN, QB=>nx14689, D=>nx8879, 
      CLK=>nx15703);
   ix9323 : oai22 port map ( Y=>nx9322, A0=>nx14693, A1=>nx16529, B0=>
      nx14696, B1=>nx16545);
   modgen_ram_ix74_ix775 : dff port map ( Q=>OPEN, QB=>nx14693, D=>nx8859, 
      CLK=>nx15703);
   modgen_ram_ix74_ix711 : dff port map ( Q=>OPEN, QB=>nx14696, D=>nx8849, 
      CLK=>nx15703);
   ix9305 : nand03 port map ( Y=>nx9304, A0=>nx14700, A1=>nx14710, A2=>
      nx14716);
   ix14701 : nor02_2x port map ( Y=>nx14700, A0=>nx9300, A1=>nx9292);
   ix9301 : nor04 port map ( Y=>nx9300, A0=>nx14703, A1=>address(4), A2=>
      address(5), A3=>nx15905);
   modgen_ram_ix74_ix835 : dff port map ( Q=>OPEN, QB=>nx14703, D=>nx8839, 
      CLK=>nx15705);
   ix9293 : nor03_2x port map ( Y=>nx9292, A0=>nx14707, A1=>nx15829, A2=>
      nx15905);
   modgen_ram_ix74_ix771 : dff port map ( Q=>OPEN, QB=>nx14707, D=>nx8829, 
      CLK=>nx15705);
   ix14711 : nand03 port map ( Y=>nx14710, A0=>modgen_ram_ix74_a_12_dup_358, 
      A1=>nx16233, A2=>nx16575);
   modgen_ram_ix74_ix831 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_358, 
      QB=>nx14714, D=>nx8819, CLK=>nx15705);
   ix14717 : nand03 port map ( Y=>nx14716, A0=>modgen_ram_ix74_a_28_dup_342, 
      A1=>nx16199, A2=>nx16575);
   modgen_ram_ix74_ix767 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_342, 
      QB=>nx14720, D=>nx8809, CLK=>nx15705);
   modgen_ram_ix74_ix639 : dff port map ( Q=>OPEN, QB=>nx14725, D=>nx8799, 
      CLK=>nx15705);
   modgen_ram_ix74_ix715 : dff port map ( Q=>OPEN, QB=>nx14729, D=>nx8789, 
      CLK=>nx15705);
   modgen_ram_ix74_ix707 : dff port map ( Q=>OPEN, QB=>nx14733, D=>nx8779, 
      CLK=>nx15705);
   modgen_ram_ix74_ix703 : dff port map ( Q=>OPEN, QB=>nx14736, D=>nx8769, 
      CLK=>nx15707);
   ix14740 : nor03_2x port map ( Y=>nx14739, A0=>nx9222, A1=>nx9214, A2=>
      nx9206);
   ix9223 : nor03_2x port map ( Y=>nx9222, A0=>nx14742, A1=>nx15867, A2=>
      nx15919);
   modgen_ram_ix74_ix827 : dff port map ( Q=>OPEN, QB=>nx14742, D=>nx8759, 
      CLK=>nx15707);
   ix9215 : nor03_2x port map ( Y=>nx9214, A0=>nx14746, A1=>nx15445, A2=>
      nx15907);
   modgen_ram_ix74_ix643 : dff port map ( Q=>OPEN, QB=>nx14746, D=>nx8749, 
      CLK=>nx15707);
   ix9207 : oai22 port map ( Y=>nx9206, A0=>nx14750, A1=>nx16645, B0=>
      nx14753, B1=>nx16661);
   modgen_ram_ix74_ix651 : dff port map ( Q=>OPEN, QB=>nx14750, D=>nx8739, 
      CLK=>nx15707);
   modgen_ram_ix74_ix647 : dff port map ( Q=>OPEN, QB=>nx14753, D=>nx8729, 
      CLK=>nx15707);
   ix9183 : oai22 port map ( Y=>nx9182, A0=>nx14760, A1=>nx16677, B0=>
      nx14763, B1=>nx16693);
   modgen_ram_ix74_ix795 : dff port map ( Q=>OPEN, QB=>nx14760, D=>nx8709, 
      CLK=>nx15707);
   modgen_ram_ix74_ix839 : dff port map ( Q=>OPEN, QB=>nx14763, D=>nx8719, 
      CLK=>nx15707);
   ix9165 : oai22 port map ( Y=>nx9164, A0=>nx14767, A1=>nx16709, B0=>
      nx14770, B1=>nx16725);
   modgen_ram_ix74_ix855 : dff port map ( Q=>OPEN, QB=>nx14767, D=>nx8699, 
      CLK=>nx15709);
   modgen_ram_ix74_ix791 : dff port map ( Q=>OPEN, QB=>nx14770, D=>nx8689, 
      CLK=>nx15709);
   ix14774 : nor03_2x port map ( Y=>nx14773, A0=>nx9142, A1=>nx9134, A2=>
      nx9126);
   ix9143 : nor03_2x port map ( Y=>nx9142, A0=>nx14776, A1=>nx15447, A2=>
      nx15757);
   modgen_ram_ix74_ix663 : dff port map ( Q=>OPEN, QB=>nx14776, D=>nx8679, 
      CLK=>nx15709);
   ix9135 : nor03_2x port map ( Y=>nx9134, A0=>nx14780, A1=>nx15867, A2=>
      nx15807);
   modgen_ram_ix74_ix851 : dff port map ( Q=>OPEN, QB=>nx14780, D=>nx8669, 
      CLK=>nx15709);
   ix9127 : oai22 port map ( Y=>nx9126, A0=>nx14784, A1=>nx16749, B0=>
      nx14787, B1=>nx16757);
   modgen_ram_ix74_ix659 : dff port map ( Q=>OPEN, QB=>nx14784, D=>nx8659, 
      CLK=>nx15709);
   modgen_ram_ix74_ix847 : dff port map ( Q=>OPEN, QB=>nx14787, D=>nx8649, 
      CLK=>nx15709);
   ix14791 : nor03_2x port map ( Y=>nx14790, A0=>nx9102, A1=>nx9094, A2=>
      nx9086);
   ix9103 : nor03_2x port map ( Y=>nx9102, A0=>nx14793, A1=>nx15785, A2=>
      nx15817);
   modgen_ram_ix74_ix719 : dff port map ( Q=>OPEN, QB=>nx14793, D=>nx8639, 
      CLK=>nx15709);
   ix9095 : nor03_2x port map ( Y=>nx9094, A0=>nx14797, A1=>nx15829, A2=>
      nx15809);
   modgen_ram_ix74_ix787 : dff port map ( Q=>OPEN, QB=>nx14797, D=>nx8629, 
      CLK=>nx15711);
   ix9087 : oai22 port map ( Y=>nx9086, A0=>nx14801, A1=>nx16773, B0=>
      nx14804, B1=>nx16789);
   modgen_ram_ix74_ix783 : dff port map ( Q=>OPEN, QB=>nx14801, D=>nx8619, 
      CLK=>nx15711);
   modgen_ram_ix74_ix655 : dff port map ( Q=>OPEN, QB=>nx14804, D=>nx8609, 
      CLK=>nx15711);
   ix14808 : nor03_2x port map ( Y=>nx14807, A0=>nx9064, A1=>nx9056, A2=>
      nx9048);
   ix9065 : nor03_2x port map ( Y=>nx9064, A0=>nx14810, A1=>nx15785, A2=>
      nx15809);
   modgen_ram_ix74_ix723 : dff port map ( Q=>OPEN, QB=>nx14810, D=>nx8599, 
      CLK=>nx15711);
   ix9057 : nor03_2x port map ( Y=>nx9056, A0=>nx14814, A1=>nx15787, A2=>
      nx15411);
   modgen_ram_ix74_ix731 : dff port map ( Q=>OPEN, QB=>nx14814, D=>nx8589, 
      CLK=>nx15711);
   ix9049 : oai22 port map ( Y=>nx9048, A0=>nx14818, A1=>nx16821, B0=>
      nx14821, B1=>nx16837);
   modgen_ram_ix74_ix667 : dff port map ( Q=>OPEN, QB=>nx14818, D=>nx8569, 
      CLK=>nx15711);
   modgen_ram_ix74_ix727 : dff port map ( Q=>OPEN, QB=>nx14821, D=>nx8579, 
      CLK=>nx15711);
   tri_data_out_14 : tri01 port map ( Y=>data_out(14), A=>nx14825, E=>
      write_out);
   ix10297 : oai22 port map ( Y=>nx10296, A0=>nx14831, A1=>nx16161, B0=>
      nx14836, B1=>nx16187);
   modgen_ram_ix74_ix414 : dff port map ( Q=>OPEN, QB=>nx14831, D=>nx9839, 
      CLK=>nx15713);
   modgen_ram_ix74_ix522 : dff port map ( Q=>OPEN, QB=>nx14836, D=>nx9829, 
      CLK=>nx15713);
   ix10279 : oai22 port map ( Y=>nx10278, A0=>nx14840, A1=>nx10555, B0=>
      nx14843, B1=>nx18958);
   modgen_ram_ix74_ix498 : dff port map ( Q=>OPEN, QB=>nx14840, D=>nx9809, 
      CLK=>nx15713);
   modgen_ram_ix74_ix506 : dff port map ( Q=>OPEN, QB=>nx14843, D=>nx9819, 
      CLK=>nx15713);
   ix14847 : nor02_2x port map ( Y=>nx14846, A0=>nx10258, A1=>nx10240);
   ix10259 : oai33 port map ( Y=>nx10258, A0=>nx14849, A1=>nx15869, A2=>
      nx16097, B0=>nx14852, B1=>nx15447, B2=>nx16029);
   modgen_ram_ix74_ix606 : dff port map ( Q=>OPEN, QB=>nx14849, D=>nx9789, 
      CLK=>nx15713);
   modgen_ram_ix74_ix418 : dff port map ( Q=>OPEN, QB=>nx14852, D=>nx9799, 
      CLK=>nx15713);
   ix10241 : oai22 port map ( Y=>nx10240, A0=>nx14856, A1=>nx16263, B0=>
      nx14859, B1=>nx16279);
   modgen_ram_ix74_ix542 : dff port map ( Q=>OPEN, QB=>nx14856, D=>nx9779, 
      CLK=>nx15713);
   modgen_ram_ix74_ix478 : dff port map ( Q=>OPEN, QB=>nx14859, D=>nx9769, 
      CLK=>nx15715);
   ix14863 : nor03_2x port map ( Y=>nx14862, A0=>nx10216, A1=>nx10208, A2=>
      nx10200);
   ix10217 : nor03_2x port map ( Y=>nx10216, A0=>nx14865, A1=>nx15787, A2=>
      nx16073);
   modgen_ram_ix74_ix434 : dff port map ( Q=>OPEN, QB=>nx14865, D=>nx9759, 
      CLK=>nx15715);
   ix10209 : nor03_2x port map ( Y=>nx10208, A0=>nx14869, A1=>nx15869, A2=>
      nx15411);
   modgen_ram_ix74_ix602 : dff port map ( Q=>OPEN, QB=>nx14869, D=>nx9749, 
      CLK=>nx15715);
   ix10201 : oai33 port map ( Y=>nx10200, A0=>nx14873, A1=>nx15787, A2=>
      nx15919, B0=>nx14876, B1=>nx15447, B2=>nx16073);
   modgen_ram_ix74_ix442 : dff port map ( Q=>OPEN, QB=>nx14873, D=>nx9729, 
      CLK=>nx15715);
   modgen_ram_ix74_ix370 : dff port map ( Q=>OPEN, QB=>nx14876, D=>nx9739, 
      CLK=>nx15715);
   ix14880 : nor03_2x port map ( Y=>nx14879, A0=>nx10178, A1=>nx10170, A2=>
      nx10162);
   ix10179 : nor03_2x port map ( Y=>nx10178, A0=>nx14882, A1=>nx15787, A2=>
      nx16051);
   modgen_ram_ix74_ix438 : dff port map ( Q=>OPEN, QB=>nx14882, D=>nx9719, 
      CLK=>nx15715);
   ix10171 : nor04 port map ( Y=>nx10170, A0=>nx14886, A1=>address(4), A2=>
      address(5), A3=>nx16073);
   modgen_ram_ix74_ix562 : dff port map ( Q=>OPEN, QB=>nx14886, D=>nx9709, 
      CLK=>nx15715);
   ix10163 : oai22 port map ( Y=>nx10162, A0=>nx14890, A1=>nx16331, B0=>
      nx14893, B1=>nx16347);
   modgen_ram_ix74_ix378 : dff port map ( Q=>OPEN, QB=>nx14890, D=>nx9689, 
      CLK=>nx15717);
   modgen_ram_ix74_ix374 : dff port map ( Q=>OPEN, QB=>nx14893, D=>nx9699, 
      CLK=>nx15717);
   modgen_ram_ix74_ix502 : dff port map ( Q=>OPEN, QB=>nx14900, D=>nx9679, 
      CLK=>nx15717);
   modgen_ram_ix74_ix566 : dff port map ( Q=>OPEN, QB=>nx14904, D=>nx9669, 
      CLK=>nx15717);
   ix10121 : oai22 port map ( Y=>nx10120, A0=>nx14908, A1=>nx16363, B0=>
      nx14911, B1=>nx16379);
   modgen_ram_ix74_ix546 : dff port map ( Q=>OPEN, QB=>nx14908, D=>nx9649, 
      CLK=>nx15717);
   modgen_ram_ix74_ix482 : dff port map ( Q=>OPEN, QB=>nx14911, D=>nx9659, 
      CLK=>nx15717);
   modgen_ram_ix74_ix610 : dff port map ( Q=>OPEN, QB=>nx14917, D=>nx9639, 
      CLK=>nx15717);
   modgen_ram_ix74_ix422 : dff port map ( Q=>OPEN, QB=>nx14921, D=>nx9629, 
      CLK=>nx15719);
   ix10083 : oai22 port map ( Y=>nx10082, A0=>nx14925, A1=>nx16403, B0=>
      nx14928, B1=>nx16419);
   modgen_ram_ix74_ix550 : dff port map ( Q=>OPEN, QB=>nx14925, D=>nx9609, 
      CLK=>nx15719);
   modgen_ram_ix74_ix486 : dff port map ( Q=>OPEN, QB=>nx14928, D=>nx9619, 
      CLK=>nx15719);
   modgen_ram_ix74_ix614 : dff port map ( Q=>OPEN, QB=>nx14934, D=>nx9599, 
      CLK=>nx15719);
   modgen_ram_ix74_ix426 : dff port map ( Q=>OPEN, QB=>nx14938, D=>nx9589, 
      CLK=>nx15719);
   ix10043 : oai22 port map ( Y=>nx10042, A0=>nx14942, A1=>nx16443, B0=>
      nx14945, B1=>nx16459);
   modgen_ram_ix74_ix554 : dff port map ( Q=>OPEN, QB=>nx14942, D=>nx9569, 
      CLK=>nx15719);
   modgen_ram_ix74_ix490 : dff port map ( Q=>OPEN, QB=>nx14945, D=>nx9579, 
      CLK=>nx15719);
   modgen_ram_ix74_ix618 : dff port map ( Q=>OPEN, QB=>nx14951, D=>nx9559, 
      CLK=>nx15721);
   ix10013 : nor03_2x port map ( Y=>nx10012, A0=>nx14955, A1=>nx15447, A2=>
      nx15963);
   modgen_ram_ix74_ix430 : dff port map ( Q=>OPEN, QB=>nx14955, D=>nx9549, 
      CLK=>nx15721);
   ix10005 : oai22 port map ( Y=>nx10004, A0=>nx14959, A1=>nx16483, B0=>
      nx14962, B1=>nx16499);
   modgen_ram_ix74_ix558 : dff port map ( Q=>OPEN, QB=>nx14959, D=>nx9529, 
      CLK=>nx15721);
   modgen_ram_ix74_ix494 : dff port map ( Q=>OPEN, QB=>nx14962, D=>nx9539, 
      CLK=>nx15721);
   ix9979 : oai22 port map ( Y=>nx9978, A0=>nx14972, A1=>nx16515, B0=>
      nx14975, B1=>nx16523);
   modgen_ram_ix74_ix586 : dff port map ( Q=>OPEN, QB=>nx14972, D=>nx9509, 
      CLK=>nx15721);
   modgen_ram_ix74_ix622 : dff port map ( Q=>OPEN, QB=>nx14975, D=>nx9519, 
      CLK=>nx15721);
   ix9961 : oai22 port map ( Y=>nx9960, A0=>nx14979, A1=>nx16531, B0=>
      nx14982, B1=>nx16547);
   modgen_ram_ix74_ix518 : dff port map ( Q=>OPEN, QB=>nx14979, D=>nx9499, 
      CLK=>nx15721);
   modgen_ram_ix74_ix454 : dff port map ( Q=>OPEN, QB=>nx14982, D=>nx9489, 
      CLK=>nx15723);
   ix9943 : nand03 port map ( Y=>nx9942, A0=>nx14986, A1=>nx14996, A2=>
      nx15002);
   ix14987 : nor02_2x port map ( Y=>nx14986, A0=>nx9938, A1=>nx9930);
   ix9939 : nor04 port map ( Y=>nx9938, A0=>nx14989, A1=>address(4), A2=>
      address(5), A3=>nx15907);
   modgen_ram_ix74_ix578 : dff port map ( Q=>OPEN, QB=>nx14989, D=>nx9479, 
      CLK=>nx15723);
   ix9931 : nor03_2x port map ( Y=>nx9930, A0=>nx14993, A1=>nx15831, A2=>
      nx15907);
   modgen_ram_ix74_ix514 : dff port map ( Q=>OPEN, QB=>nx14993, D=>nx9469, 
      CLK=>nx15723);
   ix14997 : nand03 port map ( Y=>nx14996, A0=>modgen_ram_ix74_a_12_dup_293, 
      A1=>nx16233, A2=>nx16575);
   modgen_ram_ix74_ix574 : dff port map ( Q=>modgen_ram_ix74_a_12_dup_293, 
      QB=>nx15000, D=>nx9459, CLK=>nx15723);
   ix15003 : nand03 port map ( Y=>nx15002, A0=>modgen_ram_ix74_a_28_dup_277, 
      A1=>nx16199, A2=>nx16575);
   modgen_ram_ix74_ix510 : dff port map ( Q=>modgen_ram_ix74_a_28_dup_277, 
      QB=>nx15006, D=>nx9449, CLK=>nx15723);
   ix15009 : nor03_2x port map ( Y=>nx15008, A0=>nx9898, A1=>nx9890, A2=>
      nx9882);
   ix9899 : nor03_2x port map ( Y=>nx9898, A0=>nx15011, A1=>nx15447, A2=>
      nx15933);
   modgen_ram_ix74_ix382 : dff port map ( Q=>OPEN, QB=>nx15011, D=>nx9439, 
      CLK=>nx15723);
   ix9891 : nor03_2x port map ( Y=>nx9890, A0=>nx15015, A1=>nx15787, A2=>
      nx15893);
   modgen_ram_ix74_ix458 : dff port map ( Q=>OPEN, QB=>nx15015, D=>nx9429, 
      CLK=>nx15723);
   ix9883 : oai22 port map ( Y=>nx9882, A0=>nx15019, A1=>nx16607, B0=>
      nx15022, B1=>nx16623);
   modgen_ram_ix74_ix450 : dff port map ( Q=>OPEN, QB=>nx15019, D=>nx9419, 
      CLK=>nx15725);
   modgen_ram_ix74_ix446 : dff port map ( Q=>OPEN, QB=>nx15022, D=>nx9409, 
      CLK=>nx15725);
   ix15026 : nor03_2x port map ( Y=>nx15025, A0=>nx9860, A1=>nx9852, A2=>
      nx9844);
   ix9861 : nor03_2x port map ( Y=>nx9860, A0=>nx15028, A1=>nx15869, A2=>
      nx15919);
   modgen_ram_ix74_ix570 : dff port map ( Q=>OPEN, QB=>nx15028, D=>nx9399, 
      CLK=>nx15725);
   ix9853 : nor03_2x port map ( Y=>nx9852, A0=>nx15032, A1=>nx15449, A2=>
      nx15907);
   modgen_ram_ix74_ix386 : dff port map ( Q=>OPEN, QB=>nx15032, D=>nx9389, 
      CLK=>nx15725);
   ix9845 : oai22 port map ( Y=>nx9844, A0=>nx15036, A1=>nx16647, B0=>
      nx15039, B1=>nx16663);
   modgen_ram_ix74_ix394 : dff port map ( Q=>OPEN, QB=>nx15036, D=>nx9379, 
      CLK=>nx15725);
   modgen_ram_ix74_ix390 : dff port map ( Q=>OPEN, QB=>nx15039, D=>nx9369, 
      CLK=>nx15725);
   ix9821 : oai22 port map ( Y=>nx9820, A0=>nx15046, A1=>nx16679, B0=>
      nx15049, B1=>nx16695);
   modgen_ram_ix74_ix538 : dff port map ( Q=>OPEN, QB=>nx15046, D=>nx9349, 
      CLK=>nx15725);
   modgen_ram_ix74_ix582 : dff port map ( Q=>OPEN, QB=>nx15049, D=>nx9359, 
      CLK=>nx15727);
   ix9803 : oai22 port map ( Y=>nx9802, A0=>nx15053, A1=>nx16711, B0=>
      nx15056, B1=>nx16727);
   modgen_ram_ix74_ix598 : dff port map ( Q=>OPEN, QB=>nx15053, D=>nx9339, 
      CLK=>nx15727);
   modgen_ram_ix74_ix534 : dff port map ( Q=>OPEN, QB=>nx15056, D=>nx9329, 
      CLK=>nx15727);
   ix15060 : nor03_2x port map ( Y=>nx15059, A0=>nx9780, A1=>nx9772, A2=>
      nx9764);
   ix9781 : nor03_2x port map ( Y=>nx9780, A0=>nx15062, A1=>nx15449, A2=>
      nx15757);
   modgen_ram_ix74_ix406 : dff port map ( Q=>OPEN, QB=>nx15062, D=>nx9319, 
      CLK=>nx15727);
   ix9773 : nor03_2x port map ( Y=>nx9772, A0=>nx15066, A1=>nx15869, A2=>
      nx15809);
   modgen_ram_ix74_ix594 : dff port map ( Q=>OPEN, QB=>nx15066, D=>nx9309, 
      CLK=>nx15727);
   ix9765 : oai22 port map ( Y=>nx9764, A0=>nx15070, A1=>nx16751, B0=>
      nx15073, B1=>nx16759);
   modgen_ram_ix74_ix402 : dff port map ( Q=>OPEN, QB=>nx15070, D=>nx9299, 
      CLK=>nx15727);
   modgen_ram_ix74_ix590 : dff port map ( Q=>OPEN, QB=>nx15073, D=>nx9289, 
      CLK=>nx15727);
   ix15077 : nor03_2x port map ( Y=>nx15076, A0=>nx9740, A1=>nx9732, A2=>
      nx9724);
   ix9741 : nor03_2x port map ( Y=>nx9740, A0=>nx15079, A1=>nx15787, A2=>
      nx15817);
   modgen_ram_ix74_ix462 : dff port map ( Q=>OPEN, QB=>nx15079, D=>nx9279, 
      CLK=>nx15729);
   ix9733 : nor03_2x port map ( Y=>nx9732, A0=>nx15083, A1=>nx15831, A2=>
      nx15809);
   modgen_ram_ix74_ix530 : dff port map ( Q=>OPEN, QB=>nx15083, D=>nx9269, 
      CLK=>nx15729);
   ix9725 : oai22 port map ( Y=>nx9724, A0=>nx15087, A1=>nx16775, B0=>
      nx15090, B1=>nx16791);
   modgen_ram_ix74_ix526 : dff port map ( Q=>OPEN, QB=>nx15087, D=>nx9259, 
      CLK=>nx15729);
   modgen_ram_ix74_ix398 : dff port map ( Q=>OPEN, QB=>nx15090, D=>nx9249, 
      CLK=>nx15729);
   ix15094 : nor03_2x port map ( Y=>nx15093, A0=>nx9702, A1=>nx9694, A2=>
      nx9686);
   ix9703 : nor03_2x port map ( Y=>nx9702, A0=>nx15096, A1=>nx15787, A2=>
      nx15809);
   modgen_ram_ix74_ix466 : dff port map ( Q=>OPEN, QB=>nx15096, D=>nx9239, 
      CLK=>nx15729);
   ix9695 : nor03_2x port map ( Y=>nx9694, A0=>nx15100, A1=>nx15789, A2=>
      nx15411);
   modgen_ram_ix74_ix474 : dff port map ( Q=>OPEN, QB=>nx15100, D=>nx9229, 
      CLK=>nx15729);
   ix9687 : oai22 port map ( Y=>nx9686, A0=>nx15104, A1=>nx16823, B0=>
      nx15107, B1=>nx16839);
   modgen_ram_ix74_ix410 : dff port map ( Q=>OPEN, QB=>nx15104, D=>nx9209, 
      CLK=>nx15729);
   modgen_ram_ix74_ix470 : dff port map ( Q=>OPEN, QB=>nx15107, D=>nx9219, 
      CLK=>nx15731);
   tri_data_out_15 : tri01 port map ( Y=>data_out(15), A=>nx15111, E=>
      write_out);
   ix10935 : oai22 port map ( Y=>nx10934, A0=>nx15117, A1=>nx16161, B0=>
      nx15122, B1=>nx16187);
   modgen_ram_ix74_ix155 : dff port map ( Q=>OPEN, QB=>nx15117, D=>nx10479, 
      CLK=>nx15731);
   modgen_ram_ix74_ix263 : dff port map ( Q=>OPEN, QB=>nx15122, D=>nx10469, 
      CLK=>nx15731);
   ix10917 : oai22 port map ( Y=>nx10916, A0=>nx15126, A1=>nx10555, B0=>
      nx15129, B1=>nx18958);
   modgen_ram_ix74_ix239 : dff port map ( Q=>OPEN, QB=>nx15126, D=>nx10449, 
      CLK=>nx15731);
   modgen_ram_ix74_ix247 : dff port map ( Q=>OPEN, QB=>nx15129, D=>nx10459, 
      CLK=>nx15731);
   ix15133 : nor02_2x port map ( Y=>nx15132, A0=>nx10896, A1=>nx10878);
   ix10897 : oai33 port map ( Y=>nx10896, A0=>nx15135, A1=>nx15869, A2=>
      nx16097, B0=>nx15138, B1=>nx15449, B2=>nx16029);
   modgen_ram_ix74_ix347 : dff port map ( Q=>OPEN, QB=>nx15135, D=>nx10429, 
      CLK=>nx15731);
   modgen_ram_ix74_ix159 : dff port map ( Q=>OPEN, QB=>nx15138, D=>nx10439, 
      CLK=>nx15731);
   ix10879 : oai22 port map ( Y=>nx10878, A0=>nx15142, A1=>nx16263, B0=>
      nx15145, B1=>nx16279);
   modgen_ram_ix74_ix283 : dff port map ( Q=>OPEN, QB=>nx15142, D=>nx10419, 
      CLK=>nx15733);
   modgen_ram_ix74_ix219 : dff port map ( Q=>OPEN, QB=>nx15145, D=>nx10409, 
      CLK=>nx15733);
   ix15149 : nor03_2x port map ( Y=>nx15148, A0=>nx10854, A1=>nx10846, A2=>
      nx10838);
   ix10855 : nor03_2x port map ( Y=>nx10854, A0=>nx15151, A1=>nx15789, A2=>
      nx16073);
   modgen_ram_ix74_ix175 : dff port map ( Q=>OPEN, QB=>nx15151, D=>nx10399, 
      CLK=>nx15733);
   ix10847 : nor03_2x port map ( Y=>nx10846, A0=>nx15155, A1=>nx15869, A2=>
      nx15413);
   modgen_ram_ix74_ix343 : dff port map ( Q=>OPEN, QB=>nx15155, D=>nx10389, 
      CLK=>nx15733);
   ix10839 : oai33 port map ( Y=>nx10838, A0=>nx15159, A1=>nx15789, A2=>
      nx15919, B0=>nx15162, B1=>nx15449, B2=>nx16073);
   modgen_ram_ix74_ix183 : dff port map ( Q=>OPEN, QB=>nx15159, D=>nx10369, 
      CLK=>nx15733);
   modgen_ram_ix74_ix111 : dff port map ( Q=>OPEN, QB=>nx15162, D=>nx10379, 
      CLK=>nx15733);
   ix15166 : nor03_2x port map ( Y=>nx15165, A0=>nx10816, A1=>nx10808, A2=>
      nx10800);
   ix10817 : nor03_2x port map ( Y=>nx10816, A0=>nx15168, A1=>nx15789, A2=>
      nx16051);
   modgen_ram_ix74_ix179 : dff port map ( Q=>OPEN, QB=>nx15168, D=>nx10359, 
      CLK=>nx15733);
   ix10809 : nor04 port map ( Y=>nx10808, A0=>nx15172, A1=>address(4), A2=>
      address(5), A3=>nx16073);
   modgen_ram_ix74_ix303 : dff port map ( Q=>OPEN, QB=>nx15172, D=>nx10349, 
      CLK=>nx15735);
   ix10801 : oai22 port map ( Y=>nx10800, A0=>nx15176, A1=>nx16331, B0=>
      nx15179, B1=>nx16347);
   modgen_ram_ix74_ix119 : dff port map ( Q=>OPEN, QB=>nx15176, D=>nx10329, 
      CLK=>nx15735);
   modgen_ram_ix74_ix115 : dff port map ( Q=>OPEN, QB=>nx15179, D=>nx10339, 
      CLK=>nx15735);
   modgen_ram_ix74_ix243 : dff port map ( Q=>OPEN, QB=>nx15186, D=>nx10319, 
      CLK=>nx15735);
   modgen_ram_ix74_ix307 : dff port map ( Q=>OPEN, QB=>nx15190, D=>nx10309, 
      CLK=>nx15735);
   ix10759 : oai22 port map ( Y=>nx10758, A0=>nx15194, A1=>nx16363, B0=>
      nx15197, B1=>nx16379);
   modgen_ram_ix74_ix287 : dff port map ( Q=>OPEN, QB=>nx15194, D=>nx10289, 
      CLK=>nx15735);
   modgen_ram_ix74_ix223 : dff port map ( Q=>OPEN, QB=>nx15197, D=>nx10299, 
      CLK=>nx15735);
   modgen_ram_ix74_ix351 : dff port map ( Q=>OPEN, QB=>nx15203, D=>nx10279, 
      CLK=>nx15737);
   modgen_ram_ix74_ix163 : dff port map ( Q=>OPEN, QB=>nx15207, D=>nx10269, 
      CLK=>nx15737);
   ix10721 : oai22 port map ( Y=>nx10720, A0=>nx15211, A1=>nx16403, B0=>
      nx15214, B1=>nx16419);
   modgen_ram_ix74_ix291 : dff port map ( Q=>OPEN, QB=>nx15211, D=>nx10249, 
      CLK=>nx15737);
   modgen_ram_ix74_ix227 : dff port map ( Q=>OPEN, QB=>nx15214, D=>nx10259, 
      CLK=>nx15737);
   modgen_ram_ix74_ix355 : dff port map ( Q=>OPEN, QB=>nx15220, D=>nx10239, 
      CLK=>nx15737);
   modgen_ram_ix74_ix167 : dff port map ( Q=>OPEN, QB=>nx15224, D=>nx10229, 
      CLK=>nx15737);
   ix10681 : oai22 port map ( Y=>nx10680, A0=>nx15228, A1=>nx16443, B0=>
      nx15231, B1=>nx16459);
   modgen_ram_ix74_ix295 : dff port map ( Q=>OPEN, QB=>nx15228, D=>nx10209, 
      CLK=>nx15737);
   modgen_ram_ix74_ix231 : dff port map ( Q=>OPEN, QB=>nx15231, D=>nx10219, 
      CLK=>nx15739);
   modgen_ram_ix74_ix359 : dff port map ( Q=>OPEN, QB=>nx15237, D=>nx10199, 
      CLK=>nx15739);
   ix10651 : nor03_2x port map ( Y=>nx10650, A0=>nx15241, A1=>nx15449, A2=>
      nx15963);
   modgen_ram_ix74_ix171 : dff port map ( Q=>OPEN, QB=>nx15241, D=>nx10189, 
      CLK=>nx15739);
   ix10643 : oai22 port map ( Y=>nx10642, A0=>nx15245, A1=>nx16483, B0=>
      nx15248, B1=>nx16499);
   modgen_ram_ix74_ix299 : dff port map ( Q=>OPEN, QB=>nx15245, D=>nx10169, 
      CLK=>nx15739);
   modgen_ram_ix74_ix235 : dff port map ( Q=>OPEN, QB=>nx15248, D=>nx10179, 
      CLK=>nx15739);
   ix10617 : oai22 port map ( Y=>nx10616, A0=>nx15258, A1=>nx16515, B0=>
      nx15261, B1=>nx16523);
   modgen_ram_ix74_ix327 : dff port map ( Q=>OPEN, QB=>nx15258, D=>nx10149, 
      CLK=>nx15739);
   modgen_ram_ix74_ix363 : dff port map ( Q=>OPEN, QB=>nx15261, D=>nx10159, 
      CLK=>nx15739);
   ix10599 : oai22 port map ( Y=>nx10598, A0=>nx15265, A1=>nx16531, B0=>
      nx15268, B1=>nx16547);
   modgen_ram_ix74_ix259 : dff port map ( Q=>OPEN, QB=>nx15265, D=>nx10139, 
      CLK=>nx15741);
   modgen_ram_ix74_ix195 : dff port map ( Q=>OPEN, QB=>nx15268, D=>nx10129, 
      CLK=>nx15741);
   ix10581 : nand03 port map ( Y=>nx10580, A0=>nx15272, A1=>nx15282, A2=>
      nx15288);
   ix15273 : nor02_2x port map ( Y=>nx15272, A0=>nx10576, A1=>nx10568);
   ix10577 : nor04 port map ( Y=>nx10576, A0=>nx15275, A1=>address(4), A2=>
      address(5), A3=>nx15907);
   modgen_ram_ix74_ix319 : dff port map ( Q=>OPEN, QB=>nx15275, D=>nx10119, 
      CLK=>nx15741);
   ix10569 : nor03_2x port map ( Y=>nx10568, A0=>nx15279, A1=>nx15831, A2=>
      nx15907);
   modgen_ram_ix74_ix255 : dff port map ( Q=>OPEN, QB=>nx15279, D=>nx10109, 
      CLK=>nx15741);
   ix15283 : nand03 port map ( Y=>nx15282, A0=>modgen_ram_ix74_a_12, A1=>
      nx16233, A2=>nx16575);
   modgen_ram_ix74_ix315 : dff port map ( Q=>modgen_ram_ix74_a_12, QB=>
      nx15286, D=>nx10099, CLK=>nx15741);
   ix15289 : nand03 port map ( Y=>nx15288, A0=>modgen_ram_ix74_a_28, A1=>
      nx16199, A2=>nx16575);
   modgen_ram_ix74_ix251 : dff port map ( Q=>modgen_ram_ix74_a_28, QB=>
      nx15292, D=>nx10089, CLK=>nx15741);
   ix15295 : nor03_2x port map ( Y=>nx15294, A0=>nx10536, A1=>nx10528, A2=>
      nx10520);
   ix10537 : nor03_2x port map ( Y=>nx10536, A0=>nx15297, A1=>nx15451, A2=>
      nx15933);
   modgen_ram_ix74_ix123 : dff port map ( Q=>OPEN, QB=>nx15297, D=>nx10079, 
      CLK=>nx15741);
   ix10529 : nor03_2x port map ( Y=>nx10528, A0=>nx15301, A1=>nx15789, A2=>
      nx15893);
   modgen_ram_ix74_ix199 : dff port map ( Q=>OPEN, QB=>nx15301, D=>nx10069, 
      CLK=>nx15743);
   ix10521 : oai22 port map ( Y=>nx10520, A0=>nx15305, A1=>nx16607, B0=>
      nx15308, B1=>nx16623);
   modgen_ram_ix74_ix191 : dff port map ( Q=>OPEN, QB=>nx15305, D=>nx10059, 
      CLK=>nx15743);
   modgen_ram_ix74_ix187 : dff port map ( Q=>OPEN, QB=>nx15308, D=>nx10049, 
      CLK=>nx15743);
   ix15312 : nor03_2x port map ( Y=>nx15311, A0=>nx10498, A1=>nx10490, A2=>
      nx10482);
   ix10499 : nor03_2x port map ( Y=>nx10498, A0=>nx15314, A1=>nx15871, A2=>
      nx15919);
   modgen_ram_ix74_ix311 : dff port map ( Q=>OPEN, QB=>nx15314, D=>nx10039, 
      CLK=>nx15743);
   ix10491 : nor03_2x port map ( Y=>nx10490, A0=>nx15318, A1=>nx15451, A2=>
      nx15907);
   modgen_ram_ix74_ix127 : dff port map ( Q=>OPEN, QB=>nx15318, D=>nx10029, 
      CLK=>nx15743);
   ix10483 : oai22 port map ( Y=>nx10482, A0=>nx15322, A1=>nx16647, B0=>
      nx15325, B1=>nx16663);
   modgen_ram_ix74_ix135 : dff port map ( Q=>OPEN, QB=>nx15322, D=>nx10019, 
      CLK=>nx15743);
   modgen_ram_ix74_ix131 : dff port map ( Q=>OPEN, QB=>nx15325, D=>nx10009, 
      CLK=>nx15743);
   ix10459 : oai22 port map ( Y=>nx10458, A0=>nx15332, A1=>nx16679, B0=>
      nx15335, B1=>nx16695);
   modgen_ram_ix74_ix279 : dff port map ( Q=>OPEN, QB=>nx15332, D=>nx9989, 
      CLK=>nx15745);
   modgen_ram_ix74_ix323 : dff port map ( Q=>OPEN, QB=>nx15335, D=>nx9999, 
      CLK=>nx15745);
   ix10441 : oai22 port map ( Y=>nx10440, A0=>nx15339, A1=>nx16711, B0=>
      nx15342, B1=>nx16727);
   modgen_ram_ix74_ix339 : dff port map ( Q=>OPEN, QB=>nx15339, D=>nx9979, 
      CLK=>nx15745);
   modgen_ram_ix74_ix275 : dff port map ( Q=>OPEN, QB=>nx15342, D=>nx9969, 
      CLK=>nx15745);
   ix15346 : nor03_2x port map ( Y=>nx15345, A0=>nx10418, A1=>nx10410, A2=>
      nx10402);
   ix10419 : nor03_2x port map ( Y=>nx10418, A0=>nx15348, A1=>nx15451, A2=>
      nx15757);
   modgen_ram_ix74_ix147 : dff port map ( Q=>OPEN, QB=>nx15348, D=>nx9959, 
      CLK=>nx15745);
   ix10411 : nor03_2x port map ( Y=>nx10410, A0=>nx15352, A1=>nx15871, A2=>
      nx15809);
   modgen_ram_ix74_ix335 : dff port map ( Q=>OPEN, QB=>nx15352, D=>nx9949, 
      CLK=>nx15745);
   ix10403 : oai22 port map ( Y=>nx10402, A0=>nx15356, A1=>nx16751, B0=>
      nx15359, B1=>nx16759);
   modgen_ram_ix74_ix143 : dff port map ( Q=>OPEN, QB=>nx15356, D=>nx9939, 
      CLK=>nx15745);
   modgen_ram_ix74_ix331 : dff port map ( Q=>OPEN, QB=>nx15359, D=>nx9929, 
      CLK=>nx15747);
   ix15363 : nor03_2x port map ( Y=>nx15362, A0=>nx10378, A1=>nx10370, A2=>
      nx10362);
   ix10379 : nor03_2x port map ( Y=>nx10378, A0=>nx15365, A1=>nx15789, A2=>
      nx15817);
   modgen_ram_ix74_ix203 : dff port map ( Q=>OPEN, QB=>nx15365, D=>nx9919, 
      CLK=>nx15747);
   ix10371 : nor03_2x port map ( Y=>nx10370, A0=>nx15369, A1=>nx15831, A2=>
      nx15809);
   modgen_ram_ix74_ix271 : dff port map ( Q=>OPEN, QB=>nx15369, D=>nx9909, 
      CLK=>nx15747);
   ix10363 : oai22 port map ( Y=>nx10362, A0=>nx15373, A1=>nx16775, B0=>
      nx15376, B1=>nx16791);
   modgen_ram_ix74_ix267 : dff port map ( Q=>OPEN, QB=>nx15373, D=>nx9899, 
      CLK=>nx15747);
   modgen_ram_ix74_ix139 : dff port map ( Q=>OPEN, QB=>nx15376, D=>nx9889, 
      CLK=>nx15747);
   ix15380 : nor03_2x port map ( Y=>nx15379, A0=>nx10340, A1=>nx10332, A2=>
      nx10324);
   ix10341 : nor03_2x port map ( Y=>nx10340, A0=>nx15382, A1=>nx15789, A2=>
      nx98);
   modgen_ram_ix74_ix207 : dff port map ( Q=>OPEN, QB=>nx15382, D=>nx9879, 
      CLK=>nx15747);
   ix10333 : nor03_2x port map ( Y=>nx10332, A0=>nx15386, A1=>nx15791, A2=>
      nx15413);
   modgen_ram_ix74_ix215 : dff port map ( Q=>OPEN, QB=>nx15386, D=>nx9869, 
      CLK=>nx15747);
   ix10325 : oai22 port map ( Y=>nx10324, A0=>nx15390, A1=>nx16823, B0=>
      nx15393, B1=>nx16839);
   modgen_ram_ix74_ix151 : dff port map ( Q=>OPEN, QB=>nx15390, D=>nx9849, 
      CLK=>nx15749);
   modgen_ram_ix74_ix211 : dff port map ( Q=>OPEN, QB=>nx15393, D=>nx9859, 
      CLK=>nx15749);
   ix15400 : inv01 port map ( Y=>nx15401, A=>nx8);
   ix15402 : inv02 port map ( Y=>nx15403, A=>nx15401);
   ix15404 : inv02 port map ( Y=>nx15405, A=>nx15401);
   ix15406 : inv02 port map ( Y=>nx15407, A=>nx15401);
   ix15408 : inv02 port map ( Y=>nx15409, A=>nx15401);
   ix15410 : inv02 port map ( Y=>nx15411, A=>nx15401);
   ix15412 : inv02 port map ( Y=>nx15413, A=>nx15401);
   ix15414 : buf02 port map ( Y=>nx15415, A=>nx17153);
   ix15416 : buf02 port map ( Y=>nx15417, A=>nx17153);
   ix15418 : buf02 port map ( Y=>nx15419, A=>nx17153);
   ix15420 : buf02 port map ( Y=>nx15421, A=>nx17153);
   ix15422 : buf02 port map ( Y=>nx15423, A=>nx17153);
   ix15424 : buf02 port map ( Y=>nx15425, A=>nx17153);
   ix15426 : buf02 port map ( Y=>nx15427, A=>nx17153);
   ix15428 : buf02 port map ( Y=>nx15429, A=>nx17155);
   ix15430 : buf02 port map ( Y=>nx15431, A=>nx17155);
   ix15432 : buf02 port map ( Y=>nx15433, A=>nx17155);
   ix15434 : buf02 port map ( Y=>nx15435, A=>nx17155);
   ix15436 : buf02 port map ( Y=>nx15437, A=>nx17155);
   ix15438 : buf02 port map ( Y=>nx15439, A=>nx17155);
   ix15440 : buf02 port map ( Y=>nx15441, A=>nx17155);
   ix15442 : buf02 port map ( Y=>nx15443, A=>nx14);
   ix15444 : buf02 port map ( Y=>nx15445, A=>nx14);
   ix15446 : buf02 port map ( Y=>nx15447, A=>nx14);
   ix15448 : buf02 port map ( Y=>nx15449, A=>nx14);
   ix15450 : buf02 port map ( Y=>nx15451, A=>nx14);
   ix15452 : nor02_2x port map ( Y=>nx15453, A0=>nx10514, A1=>nx15415);
   ix15454 : nor02_2x port map ( Y=>nx15455, A0=>nx10514, A1=>nx15415);
   ix15456 : inv02 port map ( Y=>nx15457, A=>clk);
   ix15458 : inv02 port map ( Y=>nx15459, A=>clk);
   ix15460 : inv02 port map ( Y=>nx15461, A=>clk);
   ix15462 : inv02 port map ( Y=>nx15463, A=>clk);
   ix15464 : inv02 port map ( Y=>nx15465, A=>clk);
   ix15466 : inv02 port map ( Y=>nx15467, A=>clk);
   ix15468 : inv02 port map ( Y=>nx15469, A=>clk);
   ix15470 : inv02 port map ( Y=>nx15471, A=>clk);
   ix15472 : inv02 port map ( Y=>nx15473, A=>clk);
   ix15474 : inv02 port map ( Y=>nx15475, A=>clk);
   ix15476 : inv02 port map ( Y=>nx15477, A=>clk);
   ix15478 : inv02 port map ( Y=>nx15479, A=>clk);
   ix15480 : inv02 port map ( Y=>nx15481, A=>clk);
   ix15482 : inv02 port map ( Y=>nx15483, A=>clk);
   ix15484 : inv02 port map ( Y=>nx15485, A=>clk);
   ix15486 : inv02 port map ( Y=>nx15487, A=>clk);
   ix15488 : inv02 port map ( Y=>nx15489, A=>clk);
   ix15490 : inv02 port map ( Y=>nx15491, A=>clk);
   ix15492 : inv02 port map ( Y=>nx15493, A=>clk);
   ix15494 : inv02 port map ( Y=>nx15495, A=>clk);
   ix15496 : inv02 port map ( Y=>nx15497, A=>clk);
   ix15498 : inv02 port map ( Y=>nx15499, A=>clk);
   ix15500 : inv02 port map ( Y=>nx15501, A=>clk);
   ix15502 : inv02 port map ( Y=>nx15503, A=>clk);
   ix15504 : inv02 port map ( Y=>nx15505, A=>clk);
   ix15506 : inv02 port map ( Y=>nx15507, A=>clk);
   ix15508 : inv02 port map ( Y=>nx15509, A=>clk);
   ix15510 : inv02 port map ( Y=>nx15511, A=>clk);
   ix15512 : inv02 port map ( Y=>nx15513, A=>clk);
   ix15514 : inv02 port map ( Y=>nx15515, A=>clk);
   ix15516 : inv02 port map ( Y=>nx15517, A=>clk);
   ix15518 : inv02 port map ( Y=>nx15519, A=>clk);
   ix15520 : inv02 port map ( Y=>nx15521, A=>clk);
   ix15522 : inv02 port map ( Y=>nx15523, A=>clk);
   ix15524 : inv02 port map ( Y=>nx15525, A=>clk);
   ix15526 : inv02 port map ( Y=>nx15527, A=>clk);
   ix15528 : inv02 port map ( Y=>nx15529, A=>clk);
   ix15530 : inv02 port map ( Y=>nx15531, A=>clk);
   ix15532 : inv02 port map ( Y=>nx15533, A=>clk);
   ix15534 : inv02 port map ( Y=>nx15535, A=>clk);
   ix15536 : inv02 port map ( Y=>nx15537, A=>clk);
   ix15538 : inv02 port map ( Y=>nx15539, A=>clk);
   ix15540 : inv02 port map ( Y=>nx15541, A=>clk);
   ix15542 : inv02 port map ( Y=>nx15543, A=>clk);
   ix15544 : inv02 port map ( Y=>nx15545, A=>clk);
   ix15546 : inv02 port map ( Y=>nx15547, A=>clk);
   ix15548 : inv02 port map ( Y=>nx15549, A=>clk);
   ix15550 : inv02 port map ( Y=>nx15551, A=>clk);
   ix15552 : inv02 port map ( Y=>nx15553, A=>clk);
   ix15554 : inv02 port map ( Y=>nx15555, A=>clk);
   ix15556 : inv02 port map ( Y=>nx15557, A=>clk);
   ix15558 : inv02 port map ( Y=>nx15559, A=>clk);
   ix15560 : inv02 port map ( Y=>nx15561, A=>clk);
   ix15562 : inv02 port map ( Y=>nx15563, A=>clk);
   ix15564 : inv02 port map ( Y=>nx15565, A=>clk);
   ix15566 : inv02 port map ( Y=>nx15567, A=>clk);
   ix15568 : inv02 port map ( Y=>nx15569, A=>clk);
   ix15570 : inv02 port map ( Y=>nx15571, A=>clk);
   ix15572 : inv02 port map ( Y=>nx15573, A=>clk);
   ix15574 : inv02 port map ( Y=>nx15575, A=>clk);
   ix15576 : inv02 port map ( Y=>nx15577, A=>clk);
   ix15578 : inv02 port map ( Y=>nx15579, A=>clk);
   ix15580 : inv02 port map ( Y=>nx15581, A=>clk);
   ix15582 : inv02 port map ( Y=>nx15583, A=>clk);
   ix15584 : inv02 port map ( Y=>nx15585, A=>clk);
   ix15586 : inv02 port map ( Y=>nx15587, A=>clk);
   ix15588 : inv02 port map ( Y=>nx15589, A=>clk);
   ix15590 : inv02 port map ( Y=>nx15591, A=>clk);
   ix15592 : inv02 port map ( Y=>nx15593, A=>clk);
   ix15594 : inv02 port map ( Y=>nx15595, A=>clk);
   ix15596 : inv02 port map ( Y=>nx15597, A=>clk);
   ix15598 : inv02 port map ( Y=>nx15599, A=>clk);
   ix15600 : inv02 port map ( Y=>nx15601, A=>clk);
   ix15602 : inv02 port map ( Y=>nx15603, A=>clk);
   ix15604 : inv02 port map ( Y=>nx15605, A=>clk);
   ix15606 : inv02 port map ( Y=>nx15607, A=>clk);
   ix15608 : inv02 port map ( Y=>nx15609, A=>clk);
   ix15610 : inv02 port map ( Y=>nx15611, A=>clk);
   ix15612 : inv02 port map ( Y=>nx15613, A=>clk);
   ix15614 : inv02 port map ( Y=>nx15615, A=>clk);
   ix15616 : inv02 port map ( Y=>nx15617, A=>clk);
   ix15618 : inv02 port map ( Y=>nx15619, A=>clk);
   ix15620 : inv02 port map ( Y=>nx15621, A=>clk);
   ix15622 : inv02 port map ( Y=>nx15623, A=>clk);
   ix15624 : inv02 port map ( Y=>nx15625, A=>clk);
   ix15626 : inv02 port map ( Y=>nx15627, A=>clk);
   ix15628 : inv02 port map ( Y=>nx15629, A=>clk);
   ix15630 : inv02 port map ( Y=>nx15631, A=>clk);
   ix15632 : inv02 port map ( Y=>nx15633, A=>clk);
   ix15634 : inv02 port map ( Y=>nx15635, A=>clk);
   ix15636 : inv02 port map ( Y=>nx15637, A=>clk);
   ix15638 : inv02 port map ( Y=>nx15639, A=>clk);
   ix15640 : inv02 port map ( Y=>nx15641, A=>clk);
   ix15642 : inv02 port map ( Y=>nx15643, A=>clk);
   ix15644 : inv02 port map ( Y=>nx15645, A=>clk);
   ix15646 : inv02 port map ( Y=>nx15647, A=>clk);
   ix15648 : inv02 port map ( Y=>nx15649, A=>clk);
   ix15650 : inv02 port map ( Y=>nx15651, A=>clk);
   ix15652 : inv02 port map ( Y=>nx15653, A=>clk);
   ix15654 : inv02 port map ( Y=>nx15655, A=>clk);
   ix15656 : inv02 port map ( Y=>nx15657, A=>clk);
   ix15658 : inv02 port map ( Y=>nx15659, A=>clk);
   ix15660 : inv02 port map ( Y=>nx15661, A=>clk);
   ix15662 : inv02 port map ( Y=>nx15663, A=>clk);
   ix15664 : inv02 port map ( Y=>nx15665, A=>clk);
   ix15666 : inv02 port map ( Y=>nx15667, A=>clk);
   ix15668 : inv02 port map ( Y=>nx15669, A=>clk);
   ix15670 : inv02 port map ( Y=>nx15671, A=>clk);
   ix15672 : inv02 port map ( Y=>nx15673, A=>clk);
   ix15674 : inv02 port map ( Y=>nx15675, A=>clk);
   ix15676 : inv02 port map ( Y=>nx15677, A=>clk);
   ix15678 : inv02 port map ( Y=>nx15679, A=>clk);
   ix15680 : inv02 port map ( Y=>nx15681, A=>clk);
   ix15682 : inv02 port map ( Y=>nx15683, A=>clk);
   ix15684 : inv02 port map ( Y=>nx15685, A=>clk);
   ix15686 : inv02 port map ( Y=>nx15687, A=>clk);
   ix15688 : inv02 port map ( Y=>nx15689, A=>clk);
   ix15690 : inv02 port map ( Y=>nx15691, A=>clk);
   ix15692 : inv02 port map ( Y=>nx15693, A=>clk);
   ix15694 : inv02 port map ( Y=>nx15695, A=>clk);
   ix15696 : inv02 port map ( Y=>nx15697, A=>clk);
   ix15698 : inv02 port map ( Y=>nx15699, A=>clk);
   ix15700 : inv02 port map ( Y=>nx15701, A=>clk);
   ix15702 : inv02 port map ( Y=>nx15703, A=>clk);
   ix15704 : inv02 port map ( Y=>nx15705, A=>clk);
   ix15706 : inv02 port map ( Y=>nx15707, A=>clk);
   ix15708 : inv02 port map ( Y=>nx15709, A=>clk);
   ix15710 : inv02 port map ( Y=>nx15711, A=>clk);
   ix15712 : inv02 port map ( Y=>nx15713, A=>clk);
   ix15714 : inv02 port map ( Y=>nx15715, A=>clk);
   ix15716 : inv02 port map ( Y=>nx15717, A=>clk);
   ix15718 : inv02 port map ( Y=>nx15719, A=>clk);
   ix15720 : inv02 port map ( Y=>nx15721, A=>clk);
   ix15722 : inv02 port map ( Y=>nx15723, A=>clk);
   ix15724 : inv02 port map ( Y=>nx15725, A=>clk);
   ix15726 : inv02 port map ( Y=>nx15727, A=>clk);
   ix15728 : inv02 port map ( Y=>nx15729, A=>clk);
   ix15730 : inv02 port map ( Y=>nx15731, A=>clk);
   ix15732 : inv02 port map ( Y=>nx15733, A=>clk);
   ix15734 : inv02 port map ( Y=>nx15735, A=>clk);
   ix15736 : inv02 port map ( Y=>nx15737, A=>clk);
   ix15738 : inv02 port map ( Y=>nx15739, A=>clk);
   ix15740 : inv02 port map ( Y=>nx15741, A=>clk);
   ix15742 : inv02 port map ( Y=>nx15743, A=>clk);
   ix15744 : inv02 port map ( Y=>nx15745, A=>clk);
   ix15746 : inv02 port map ( Y=>nx15747, A=>clk);
   ix15748 : inv02 port map ( Y=>nx15749, A=>clk);
   ix15750 : inv01 port map ( Y=>nx15751, A=>nx44);
   ix15752 : inv02 port map ( Y=>nx15753, A=>nx15751);
   ix15754 : inv02 port map ( Y=>nx15755, A=>nx15751);
   ix15756 : inv02 port map ( Y=>nx15757, A=>nx15751);
   ix15758 : buf02 port map ( Y=>nx15759, A=>nx17157);
   ix15760 : buf02 port map ( Y=>nx15761, A=>nx17157);
   ix15762 : buf02 port map ( Y=>nx15763, A=>nx17157);
   ix15764 : buf02 port map ( Y=>nx15765, A=>nx17157);
   ix15766 : buf02 port map ( Y=>nx15767, A=>nx17157);
   ix15768 : buf02 port map ( Y=>nx15769, A=>nx17157);
   ix15770 : buf02 port map ( Y=>nx15771, A=>nx17157);
   ix15772 : buf02 port map ( Y=>nx15773, A=>nx17159);
   ix15774 : buf02 port map ( Y=>nx15775, A=>nx17159);
   ix15776 : buf02 port map ( Y=>nx15777, A=>nx17159);
   ix15778 : buf02 port map ( Y=>nx15779, A=>nx17159);
   ix15780 : buf02 port map ( Y=>nx15781, A=>nx17159);
   ix15782 : buf02 port map ( Y=>nx15783, A=>nx17159);
   ix15784 : buf02 port map ( Y=>nx15785, A=>nx17159);
   ix15786 : buf02 port map ( Y=>nx15787, A=>nx48);
   ix15788 : buf02 port map ( Y=>nx15789, A=>nx48);
   ix15790 : buf02 port map ( Y=>nx15791, A=>nx48);
   ix15792 : nor02_2x port map ( Y=>nx15793, A0=>nx10514, A1=>nx15759);
   ix15796 : inv04 port map ( Y=>nx15797, A=>nx17143);
   ix15798 : inv04 port map ( Y=>nx15799, A=>nx17143);
   ix15800 : inv04 port map ( Y=>nx15801, A=>nx17143);
   ix15802 : inv04 port map ( Y=>nx15803, A=>nx17143);
   ix15804 : inv04 port map ( Y=>nx15805, A=>nx17143);
   ix15806 : inv04 port map ( Y=>nx15807, A=>nx17143);
   ix15808 : inv04 port map ( Y=>nx15809, A=>nx17143);
   ix15812 : buf04 port map ( Y=>nx15813, A=>nx128);
   ix15814 : buf04 port map ( Y=>nx15815, A=>nx128);
   ix15816 : buf04 port map ( Y=>nx15817, A=>nx128);
   ix15818 : buf02 port map ( Y=>nx15819, A=>nx150);
   ix15820 : buf02 port map ( Y=>nx15821, A=>nx150);
   ix15822 : buf02 port map ( Y=>nx15823, A=>nx150);
   ix15824 : buf02 port map ( Y=>nx15825, A=>nx150);
   ix15826 : buf02 port map ( Y=>nx15827, A=>nx150);
   ix15828 : buf02 port map ( Y=>nx15829, A=>nx150);
   ix15830 : buf02 port map ( Y=>nx15831, A=>nx150);
   ix15848 : inv04 port map ( Y=>nx15849, A=>nx16233);
   ix15850 : inv04 port map ( Y=>nx15851, A=>nx16233);
   ix15852 : inv04 port map ( Y=>nx15853, A=>nx16235);
   ix15854 : inv04 port map ( Y=>nx15855, A=>nx16235);
   ix15856 : inv04 port map ( Y=>nx15857, A=>nx16235);
   ix15858 : inv04 port map ( Y=>nx15859, A=>nx16235);
   ix15860 : inv04 port map ( Y=>nx15861, A=>nx16235);
   ix15862 : inv04 port map ( Y=>nx15863, A=>nx16235);
   ix15864 : inv04 port map ( Y=>nx15865, A=>nx16235);
   ix15866 : inv04 port map ( Y=>nx15867, A=>nx16237);
   ix15868 : inv04 port map ( Y=>nx15869, A=>nx16237);
   ix15870 : inv04 port map ( Y=>nx15871, A=>nx16237);
   ix15888 : buf04 port map ( Y=>nx15889, A=>nx404);
   ix15890 : buf04 port map ( Y=>nx15891, A=>nx404);
   ix15892 : buf04 port map ( Y=>nx15893, A=>nx404);
   ix15894 : buf02 port map ( Y=>nx15895, A=>nx426);
   ix15896 : buf02 port map ( Y=>nx15897, A=>nx426);
   ix15898 : buf02 port map ( Y=>nx15899, A=>nx426);
   ix15900 : buf02 port map ( Y=>nx15901, A=>nx426);
   ix15902 : buf02 port map ( Y=>nx15903, A=>nx426);
   ix15904 : buf02 port map ( Y=>nx15905, A=>nx426);
   ix15906 : buf02 port map ( Y=>nx15907, A=>nx426);
   ix15908 : inv01 port map ( Y=>nx15909, A=>nx452);
   ix15910 : inv02 port map ( Y=>nx15911, A=>nx15909);
   ix15912 : inv02 port map ( Y=>nx15913, A=>nx15909);
   ix15914 : inv02 port map ( Y=>nx15915, A=>nx15909);
   ix15916 : inv02 port map ( Y=>nx15917, A=>nx15909);
   ix15918 : inv02 port map ( Y=>nx15919, A=>nx15909);
   ix15928 : buf04 port map ( Y=>nx15929, A=>nx476);
   ix15930 : buf04 port map ( Y=>nx15931, A=>nx476);
   ix15932 : buf04 port map ( Y=>nx15933, A=>nx476);
   ix15958 : buf04 port map ( Y=>nx15959, A=>nx694);
   ix15960 : buf04 port map ( Y=>nx15961, A=>nx694);
   ix15962 : buf04 port map ( Y=>nx15963, A=>nx694);
   ix15980 : inv02 port map ( Y=>nx15981, A=>nx780);
   ix15982 : inv04 port map ( Y=>nx15983, A=>nx15981);
   ix15984 : inv04 port map ( Y=>nx15985, A=>nx15981);
   ix15986 : inv04 port map ( Y=>nx15987, A=>nx15981);
   ix15988 : inv04 port map ( Y=>nx15989, A=>nx15981);
   ix15990 : inv04 port map ( Y=>nx15991, A=>nx15981);
   ix16000 : buf02 port map ( Y=>nx16001, A=>nx860);
   ix16002 : buf02 port map ( Y=>nx16003, A=>nx860);
   ix16004 : buf02 port map ( Y=>nx16005, A=>nx860);
   ix16006 : buf02 port map ( Y=>nx16007, A=>nx860);
   ix16008 : buf02 port map ( Y=>nx16009, A=>nx860);
   ix16018 : inv01 port map ( Y=>nx16019, A=>nx942);
   ix16020 : inv02 port map ( Y=>nx16021, A=>nx16019);
   ix16022 : inv02 port map ( Y=>nx16023, A=>nx16019);
   ix16024 : inv02 port map ( Y=>nx16025, A=>nx16019);
   ix16026 : inv02 port map ( Y=>nx16027, A=>nx16019);
   ix16028 : inv02 port map ( Y=>nx16029, A=>nx16019);
   ix16038 : buf02 port map ( Y=>nx16039, A=>nx1004);
   ix16040 : buf02 port map ( Y=>nx16041, A=>nx1004);
   ix16042 : buf02 port map ( Y=>nx16043, A=>nx1004);
   ix16044 : buf02 port map ( Y=>nx16045, A=>nx1004);
   ix16046 : buf02 port map ( Y=>nx16047, A=>nx1004);
   ix16048 : buf02 port map ( Y=>nx16049, A=>nx1004);
   ix16050 : buf02 port map ( Y=>nx16051, A=>nx1004);
   ix16060 : buf02 port map ( Y=>nx16061, A=>nx1088);
   ix16062 : buf02 port map ( Y=>nx16063, A=>nx1088);
   ix16064 : buf02 port map ( Y=>nx16065, A=>nx1088);
   ix16066 : buf02 port map ( Y=>nx16067, A=>nx1088);
   ix16068 : buf02 port map ( Y=>nx16069, A=>nx1088);
   ix16070 : buf02 port map ( Y=>nx16071, A=>nx1088);
   ix16072 : buf02 port map ( Y=>nx16073, A=>nx1088);
   ix16092 : inv02 port map ( Y=>nx16093, A=>nx16091);
   ix16094 : inv02 port map ( Y=>nx16095, A=>nx16091);
   ix16096 : inv02 port map ( Y=>nx16097, A=>nx16091);
   ix16122 : inv02 port map ( Y=>nx16123, A=>data_in(0));
   ix16124 : inv02 port map ( Y=>nx16125, A=>data_in(0));
   ix16126 : inv02 port map ( Y=>nx16127, A=>data_in(0));
   ix16128 : inv02 port map ( Y=>nx16129, A=>data_in(0));
   ix16130 : inv02 port map ( Y=>nx16131, A=>data_in(0));
   ix16132 : inv02 port map ( Y=>nx16133, A=>data_in(0));
   ix16134 : inv02 port map ( Y=>nx16135, A=>data_in(0));
   ix16136 : inv02 port map ( Y=>nx16137, A=>data_in(0));
   ix16138 : inv02 port map ( Y=>nx16139, A=>data_in(0));
   ix16140 : inv02 port map ( Y=>nx16141, A=>data_in(0));
   ix16154 : inv01 port map ( Y=>nx16155, A=>nx10519);
   ix16156 : inv02 port map ( Y=>nx16157, A=>nx16155);
   ix16158 : inv02 port map ( Y=>nx16159, A=>nx16155);
   ix16160 : inv02 port map ( Y=>nx16161, A=>nx16155);
   ix16162 : nor02_2x port map ( Y=>nx16163, A0=>nx10507, A1=>address(3));
   ix16164 : nor02_2x port map ( Y=>nx16165, A0=>nx10507, A1=>address(3));
   ix16166 : nor02_2x port map ( Y=>nx16167, A0=>address(2), A1=>nx10537);
   ix16168 : nor02_2x port map ( Y=>nx16169, A0=>address(2), A1=>nx10537);
   ix16170 : inv02 port map ( Y=>nx16171, A=>address(1));
   ix16172 : inv02 port map ( Y=>nx16173, A=>address(1));
   ix16174 : inv02 port map ( Y=>nx16175, A=>address(1));
   ix16176 : buf02 port map ( Y=>nx16177, A=>nx10541);
   ix16178 : buf02 port map ( Y=>nx16179, A=>nx10541);
   ix16180 : inv01 port map ( Y=>nx16181, A=>nx10543);
   ix16182 : inv02 port map ( Y=>nx16183, A=>nx16181);
   ix16184 : inv02 port map ( Y=>nx16185, A=>nx16181);
   ix16186 : inv02 port map ( Y=>nx16187, A=>nx16181);
   ix16190 : inv02 port map ( Y=>nx16191, A=>nx17301);
   ix16194 : inv02 port map ( Y=>nx16195, A=>nx17301);
   ix16196 : inv02 port map ( Y=>nx16197, A=>nx17301);
   ix16198 : inv02 port map ( Y=>nx16199, A=>nx17301);
   ix16212 : inv02 port map ( Y=>nx16213, A=>address(0));
   ix16214 : inv02 port map ( Y=>nx16215, A=>address(0));
   ix16224 : inv04 port map ( Y=>nx16225, A=>nx17179);
   ix16226 : inv04 port map ( Y=>nx16227, A=>nx17179);
   ix16228 : inv04 port map ( Y=>nx16229, A=>nx17179);
   ix16230 : inv04 port map ( Y=>nx16231, A=>nx17179);
   ix16232 : inv04 port map ( Y=>nx16233, A=>nx17179);
   ix16234 : inv04 port map ( Y=>nx16235, A=>nx17179);
   ix16236 : inv04 port map ( Y=>nx16237, A=>nx17179);
   ix16246 : nor02_2x port map ( Y=>nx16247, A0=>address(2), A1=>address(3)
   );
   ix16258 : inv02 port map ( Y=>nx16259, A=>nx16257);
   ix16260 : inv02 port map ( Y=>nx16261, A=>nx16257);
   ix16262 : inv02 port map ( Y=>nx16263, A=>nx16257);
   ix16272 : inv01 port map ( Y=>nx16273, A=>nx10611);
   ix16274 : inv02 port map ( Y=>nx16275, A=>nx16273);
   ix16276 : inv02 port map ( Y=>nx16277, A=>nx16273);
   ix16278 : inv02 port map ( Y=>nx16279, A=>nx16273);
   ix16280 : nor02_2x port map ( Y=>nx16281, A0=>address(4), A1=>nx10525);
   ix16324 : inv01 port map ( Y=>nx16325, A=>nx10679);
   ix16326 : inv02 port map ( Y=>nx16327, A=>nx16325);
   ix16328 : inv02 port map ( Y=>nx16329, A=>nx16325);
   ix16330 : inv02 port map ( Y=>nx16331, A=>nx16325);
   ix16340 : inv01 port map ( Y=>nx16341, A=>nx10686);
   ix16342 : inv02 port map ( Y=>nx16343, A=>nx16341);
   ix16344 : inv02 port map ( Y=>nx16345, A=>nx16341);
   ix16346 : inv02 port map ( Y=>nx16347, A=>nx16341);
   ix16356 : inv01 port map ( Y=>nx16357, A=>nx10711);
   ix16358 : inv02 port map ( Y=>nx16359, A=>nx16357);
   ix16360 : inv02 port map ( Y=>nx16361, A=>nx16357);
   ix16362 : inv02 port map ( Y=>nx16363, A=>nx16357);
   ix16372 : inv01 port map ( Y=>nx16373, A=>nx10719);
   ix16374 : inv02 port map ( Y=>nx16375, A=>nx16373);
   ix16376 : inv02 port map ( Y=>nx16377, A=>nx16373);
   ix16378 : inv02 port map ( Y=>nx16379, A=>nx16373);
   ix16396 : inv01 port map ( Y=>nx16397, A=>nx10749);
   ix16398 : inv02 port map ( Y=>nx16399, A=>nx16397);
   ix16400 : inv02 port map ( Y=>nx16401, A=>nx16397);
   ix16402 : inv02 port map ( Y=>nx16403, A=>nx16397);
   ix16412 : inv01 port map ( Y=>nx16413, A=>nx10757);
   ix16414 : inv02 port map ( Y=>nx16415, A=>nx16413);
   ix16416 : inv02 port map ( Y=>nx16417, A=>nx16413);
   ix16418 : inv02 port map ( Y=>nx16419, A=>nx16413);
   ix16436 : inv01 port map ( Y=>nx16437, A=>nx10787);
   ix16442 : inv02 port map ( Y=>nx16443, A=>nx16437);
   ix16452 : inv01 port map ( Y=>nx16453, A=>nx10795);
   ix16458 : inv02 port map ( Y=>nx16459, A=>nx16453);
   ix16476 : inv01 port map ( Y=>nx16477, A=>nx10823);
   ix16482 : inv02 port map ( Y=>nx16483, A=>nx16477);
   ix16492 : inv01 port map ( Y=>nx16493, A=>nx10831);
   ix16498 : inv02 port map ( Y=>nx16499, A=>nx16493);
   ix16508 : inv01 port map ( Y=>nx16509, A=>nx10850);
   ix16510 : inv02 port map ( Y=>nx16511, A=>nx16509);
   ix16512 : inv02 port map ( Y=>nx16513, A=>nx16509);
   ix16514 : inv02 port map ( Y=>nx16515, A=>nx16509);
   ix16516 : inv01 port map ( Y=>nx16517, A=>nx10857);
   ix16518 : inv02 port map ( Y=>nx16519, A=>nx16517);
   ix16520 : inv02 port map ( Y=>nx16521, A=>nx16517);
   ix16522 : inv02 port map ( Y=>nx16523, A=>nx16517);
   ix16524 : inv01 port map ( Y=>nx16525, A=>nx10866);
   ix16526 : inv02 port map ( Y=>nx16527, A=>nx16525);
   ix16528 : inv02 port map ( Y=>nx16529, A=>nx16525);
   ix16530 : inv02 port map ( Y=>nx16531, A=>nx16525);
   ix16540 : inv01 port map ( Y=>nx16541, A=>nx10877);
   ix16542 : inv02 port map ( Y=>nx16543, A=>nx16541);
   ix16544 : inv02 port map ( Y=>nx16545, A=>nx16541);
   ix16546 : inv02 port map ( Y=>nx16547, A=>nx16541);
   ix16566 : inv02 port map ( Y=>nx16567, A=>nx17457);
   ix16568 : inv02 port map ( Y=>nx16569, A=>nx17457);
   ix16570 : inv02 port map ( Y=>nx16571, A=>nx17457);
   ix16572 : inv02 port map ( Y=>nx16573, A=>nx17457);
   ix16574 : inv02 port map ( Y=>nx16575, A=>nx17457);
   ix16600 : inv01 port map ( Y=>nx16601, A=>nx10941);
   ix16606 : inv02 port map ( Y=>nx16607, A=>nx16601);
   ix16616 : inv01 port map ( Y=>nx16617, A=>nx10949);
   ix16618 : inv02 port map ( Y=>nx16619, A=>nx16617);
   ix16620 : inv02 port map ( Y=>nx16621, A=>nx16617);
   ix16622 : inv02 port map ( Y=>nx16623, A=>nx16617);
   ix16640 : inv01 port map ( Y=>nx16641, A=>nx10970);
   ix16642 : inv02 port map ( Y=>nx16643, A=>nx16641);
   ix16644 : inv02 port map ( Y=>nx16645, A=>nx16641);
   ix16646 : inv02 port map ( Y=>nx16647, A=>nx16641);
   ix16656 : inv01 port map ( Y=>nx16657, A=>nx10977);
   ix16658 : inv02 port map ( Y=>nx16659, A=>nx16657);
   ix16660 : inv02 port map ( Y=>nx16661, A=>nx16657);
   ix16662 : inv02 port map ( Y=>nx16663, A=>nx16657);
   ix16672 : inv01 port map ( Y=>nx16673, A=>nx10990);
   ix16674 : inv02 port map ( Y=>nx16675, A=>nx16673);
   ix16676 : inv02 port map ( Y=>nx16677, A=>nx16673);
   ix16678 : inv02 port map ( Y=>nx16679, A=>nx16673);
   ix16688 : inv01 port map ( Y=>nx16689, A=>nx10997);
   ix16690 : inv02 port map ( Y=>nx16691, A=>nx16689);
   ix16692 : inv02 port map ( Y=>nx16693, A=>nx16689);
   ix16694 : inv02 port map ( Y=>nx16695, A=>nx16689);
   ix16706 : inv02 port map ( Y=>nx16707, A=>nx16705);
   ix16708 : inv02 port map ( Y=>nx16709, A=>nx16705);
   ix16710 : inv02 port map ( Y=>nx16711, A=>nx16705);
   ix16722 : inv02 port map ( Y=>nx16723, A=>nx16721);
   ix16724 : inv02 port map ( Y=>nx16725, A=>nx16721);
   ix16726 : inv02 port map ( Y=>nx16727, A=>nx16721);
   ix16744 : inv01 port map ( Y=>nx16745, A=>nx11039);
   ix16746 : inv02 port map ( Y=>nx16747, A=>nx16745);
   ix16748 : inv02 port map ( Y=>nx16749, A=>nx16745);
   ix16750 : inv02 port map ( Y=>nx16751, A=>nx16745);
   ix16754 : inv02 port map ( Y=>nx16755, A=>nx16753);
   ix16756 : inv02 port map ( Y=>nx16757, A=>nx16753);
   ix16758 : inv02 port map ( Y=>nx16759, A=>nx16753);
   ix16770 : inv02 port map ( Y=>nx16771, A=>nx16769);
   ix16772 : inv02 port map ( Y=>nx16773, A=>nx16769);
   ix16774 : inv02 port map ( Y=>nx16775, A=>nx16769);
   ix16784 : inv01 port map ( Y=>nx16785, A=>nx11075);
   ix16786 : inv02 port map ( Y=>nx16787, A=>nx16785);
   ix16788 : inv02 port map ( Y=>nx16789, A=>nx16785);
   ix16790 : inv02 port map ( Y=>nx16791, A=>nx16785);
   ix16816 : inv01 port map ( Y=>nx16817, A=>nx11097);
   ix16818 : inv02 port map ( Y=>nx16819, A=>nx16817);
   ix16820 : inv02 port map ( Y=>nx16821, A=>nx16817);
   ix16822 : inv02 port map ( Y=>nx16823, A=>nx16817);
   ix16832 : inv01 port map ( Y=>nx16833, A=>nx11104);
   ix16834 : inv02 port map ( Y=>nx16835, A=>nx16833);
   ix16836 : inv02 port map ( Y=>nx16837, A=>nx16833);
   ix16838 : inv02 port map ( Y=>nx16839, A=>nx16833);
   ix16840 : inv02 port map ( Y=>nx16841, A=>data_in(1));
   ix16842 : inv02 port map ( Y=>nx16843, A=>data_in(1));
   ix16844 : inv02 port map ( Y=>nx16845, A=>data_in(1));
   ix16846 : inv02 port map ( Y=>nx16847, A=>data_in(1));
   ix16848 : inv02 port map ( Y=>nx16849, A=>data_in(1));
   ix16850 : inv02 port map ( Y=>nx16851, A=>data_in(1));
   ix16852 : inv02 port map ( Y=>nx16853, A=>data_in(1));
   ix16854 : inv02 port map ( Y=>nx16855, A=>data_in(1));
   ix16856 : inv02 port map ( Y=>nx16857, A=>data_in(1));
   ix16858 : inv02 port map ( Y=>nx16859, A=>data_in(1));
   ix16860 : inv02 port map ( Y=>nx16861, A=>data_in(2));
   ix16862 : inv02 port map ( Y=>nx16863, A=>data_in(2));
   ix16864 : inv02 port map ( Y=>nx16865, A=>data_in(2));
   ix16866 : inv02 port map ( Y=>nx16867, A=>data_in(2));
   ix16868 : inv02 port map ( Y=>nx16869, A=>data_in(2));
   ix16870 : inv02 port map ( Y=>nx16871, A=>data_in(2));
   ix16872 : inv02 port map ( Y=>nx16873, A=>data_in(2));
   ix16874 : inv02 port map ( Y=>nx16875, A=>data_in(2));
   ix16876 : inv02 port map ( Y=>nx16877, A=>data_in(2));
   ix16878 : inv02 port map ( Y=>nx16879, A=>data_in(2));
   ix16880 : inv02 port map ( Y=>nx16881, A=>data_in(3));
   ix16882 : inv02 port map ( Y=>nx16883, A=>data_in(3));
   ix16884 : inv02 port map ( Y=>nx16885, A=>data_in(3));
   ix16886 : inv02 port map ( Y=>nx16887, A=>data_in(3));
   ix16888 : inv02 port map ( Y=>nx16889, A=>data_in(3));
   ix16890 : inv02 port map ( Y=>nx16891, A=>data_in(3));
   ix16892 : inv02 port map ( Y=>nx16893, A=>data_in(3));
   ix16894 : inv02 port map ( Y=>nx16895, A=>data_in(3));
   ix16896 : inv02 port map ( Y=>nx16897, A=>data_in(3));
   ix16898 : inv02 port map ( Y=>nx16899, A=>data_in(3));
   ix16900 : inv02 port map ( Y=>nx16901, A=>data_in(4));
   ix16902 : inv02 port map ( Y=>nx16903, A=>data_in(4));
   ix16904 : inv02 port map ( Y=>nx16905, A=>data_in(4));
   ix16906 : inv02 port map ( Y=>nx16907, A=>data_in(4));
   ix16908 : inv02 port map ( Y=>nx16909, A=>data_in(4));
   ix16910 : inv02 port map ( Y=>nx16911, A=>data_in(4));
   ix16912 : inv02 port map ( Y=>nx16913, A=>data_in(4));
   ix16914 : inv02 port map ( Y=>nx16915, A=>data_in(4));
   ix16916 : inv02 port map ( Y=>nx16917, A=>data_in(4));
   ix16918 : inv02 port map ( Y=>nx16919, A=>data_in(4));
   ix16920 : inv02 port map ( Y=>nx16921, A=>data_in(5));
   ix16922 : inv02 port map ( Y=>nx16923, A=>data_in(5));
   ix16924 : inv02 port map ( Y=>nx16925, A=>data_in(5));
   ix16926 : inv02 port map ( Y=>nx16927, A=>data_in(5));
   ix16928 : inv02 port map ( Y=>nx16929, A=>data_in(5));
   ix16930 : inv02 port map ( Y=>nx16931, A=>data_in(5));
   ix16932 : inv02 port map ( Y=>nx16933, A=>data_in(5));
   ix16934 : inv02 port map ( Y=>nx16935, A=>data_in(5));
   ix16936 : inv02 port map ( Y=>nx16937, A=>data_in(5));
   ix16938 : inv02 port map ( Y=>nx16939, A=>data_in(5));
   ix16940 : inv02 port map ( Y=>nx16941, A=>data_in(6));
   ix16942 : inv02 port map ( Y=>nx16943, A=>data_in(6));
   ix16944 : inv02 port map ( Y=>nx16945, A=>data_in(6));
   ix16946 : inv02 port map ( Y=>nx16947, A=>data_in(6));
   ix16948 : inv02 port map ( Y=>nx16949, A=>data_in(6));
   ix16950 : inv02 port map ( Y=>nx16951, A=>data_in(6));
   ix16952 : inv02 port map ( Y=>nx16953, A=>data_in(6));
   ix16954 : inv02 port map ( Y=>nx16955, A=>data_in(6));
   ix16956 : inv02 port map ( Y=>nx16957, A=>data_in(6));
   ix16958 : inv02 port map ( Y=>nx16959, A=>data_in(6));
   ix16960 : inv02 port map ( Y=>nx16961, A=>data_in(7));
   ix16962 : inv02 port map ( Y=>nx16963, A=>data_in(7));
   ix16964 : inv02 port map ( Y=>nx16965, A=>data_in(7));
   ix16966 : inv02 port map ( Y=>nx16967, A=>data_in(7));
   ix16968 : inv02 port map ( Y=>nx16969, A=>data_in(7));
   ix16970 : inv02 port map ( Y=>nx16971, A=>data_in(7));
   ix16972 : inv02 port map ( Y=>nx16973, A=>data_in(7));
   ix16974 : inv02 port map ( Y=>nx16975, A=>data_in(7));
   ix16976 : inv02 port map ( Y=>nx16977, A=>data_in(7));
   ix16978 : inv02 port map ( Y=>nx16979, A=>data_in(7));
   ix16980 : inv02 port map ( Y=>nx16981, A=>data_in(8));
   ix16982 : inv02 port map ( Y=>nx16983, A=>data_in(8));
   ix16984 : inv02 port map ( Y=>nx16985, A=>data_in(8));
   ix16986 : inv02 port map ( Y=>nx16987, A=>data_in(8));
   ix16988 : inv02 port map ( Y=>nx16989, A=>data_in(8));
   ix16990 : inv02 port map ( Y=>nx16991, A=>data_in(8));
   ix16992 : inv02 port map ( Y=>nx16993, A=>data_in(8));
   ix16994 : inv02 port map ( Y=>nx16995, A=>data_in(8));
   ix16996 : inv02 port map ( Y=>nx16997, A=>data_in(8));
   ix16998 : inv02 port map ( Y=>nx16999, A=>data_in(8));
   ix17000 : inv02 port map ( Y=>nx17001, A=>data_in(9));
   ix17002 : inv02 port map ( Y=>nx17003, A=>data_in(9));
   ix17004 : inv02 port map ( Y=>nx17005, A=>data_in(9));
   ix17006 : inv02 port map ( Y=>nx17007, A=>data_in(9));
   ix17008 : inv02 port map ( Y=>nx17009, A=>data_in(9));
   ix17010 : inv02 port map ( Y=>nx17011, A=>data_in(9));
   ix17012 : inv02 port map ( Y=>nx17013, A=>data_in(9));
   ix17014 : inv02 port map ( Y=>nx17015, A=>data_in(9));
   ix17016 : inv02 port map ( Y=>nx17017, A=>data_in(9));
   ix17018 : inv02 port map ( Y=>nx17019, A=>data_in(9));
   ix17020 : inv02 port map ( Y=>nx17021, A=>data_in(10));
   ix17022 : inv02 port map ( Y=>nx17023, A=>data_in(10));
   ix17024 : inv02 port map ( Y=>nx17025, A=>data_in(10));
   ix17026 : inv02 port map ( Y=>nx17027, A=>data_in(10));
   ix17028 : inv02 port map ( Y=>nx17029, A=>data_in(10));
   ix17030 : inv02 port map ( Y=>nx17031, A=>data_in(10));
   ix17032 : inv02 port map ( Y=>nx17033, A=>data_in(10));
   ix17034 : inv02 port map ( Y=>nx17035, A=>data_in(10));
   ix17036 : inv02 port map ( Y=>nx17037, A=>data_in(10));
   ix17038 : inv02 port map ( Y=>nx17039, A=>data_in(10));
   ix17040 : inv02 port map ( Y=>nx17041, A=>data_in(11));
   ix17042 : inv02 port map ( Y=>nx17043, A=>data_in(11));
   ix17044 : inv02 port map ( Y=>nx17045, A=>data_in(11));
   ix17046 : inv02 port map ( Y=>nx17047, A=>data_in(11));
   ix17048 : inv02 port map ( Y=>nx17049, A=>data_in(11));
   ix17050 : inv02 port map ( Y=>nx17051, A=>data_in(11));
   ix17052 : inv02 port map ( Y=>nx17053, A=>data_in(11));
   ix17054 : inv02 port map ( Y=>nx17055, A=>data_in(11));
   ix17056 : inv02 port map ( Y=>nx17057, A=>data_in(11));
   ix17058 : inv02 port map ( Y=>nx17059, A=>data_in(11));
   ix17060 : inv02 port map ( Y=>nx17061, A=>data_in(12));
   ix17062 : inv02 port map ( Y=>nx17063, A=>data_in(12));
   ix17064 : inv02 port map ( Y=>nx17065, A=>data_in(12));
   ix17066 : inv02 port map ( Y=>nx17067, A=>data_in(12));
   ix17068 : inv02 port map ( Y=>nx17069, A=>data_in(12));
   ix17070 : inv02 port map ( Y=>nx17071, A=>data_in(12));
   ix17072 : inv02 port map ( Y=>nx17073, A=>data_in(12));
   ix17074 : inv02 port map ( Y=>nx17075, A=>data_in(12));
   ix17076 : inv02 port map ( Y=>nx17077, A=>data_in(12));
   ix17078 : inv02 port map ( Y=>nx17079, A=>data_in(12));
   ix17080 : inv02 port map ( Y=>nx17081, A=>data_in(13));
   ix17082 : inv02 port map ( Y=>nx17083, A=>data_in(13));
   ix17084 : inv02 port map ( Y=>nx17085, A=>data_in(13));
   ix17086 : inv02 port map ( Y=>nx17087, A=>data_in(13));
   ix17088 : inv02 port map ( Y=>nx17089, A=>data_in(13));
   ix17090 : inv02 port map ( Y=>nx17091, A=>data_in(13));
   ix17092 : inv02 port map ( Y=>nx17093, A=>data_in(13));
   ix17094 : inv02 port map ( Y=>nx17095, A=>data_in(13));
   ix17096 : inv02 port map ( Y=>nx17097, A=>data_in(13));
   ix17098 : inv02 port map ( Y=>nx17099, A=>data_in(13));
   ix17100 : inv02 port map ( Y=>nx17101, A=>data_in(14));
   ix17102 : inv02 port map ( Y=>nx17103, A=>data_in(14));
   ix17104 : inv02 port map ( Y=>nx17105, A=>data_in(14));
   ix17106 : inv02 port map ( Y=>nx17107, A=>data_in(14));
   ix17108 : inv02 port map ( Y=>nx17109, A=>data_in(14));
   ix17110 : inv02 port map ( Y=>nx17111, A=>data_in(14));
   ix17112 : inv02 port map ( Y=>nx17113, A=>data_in(14));
   ix17114 : inv02 port map ( Y=>nx17115, A=>data_in(14));
   ix17116 : inv02 port map ( Y=>nx17117, A=>data_in(14));
   ix17118 : inv02 port map ( Y=>nx17119, A=>data_in(14));
   ix17120 : inv02 port map ( Y=>nx17121, A=>data_in(15));
   ix17122 : inv02 port map ( Y=>nx17123, A=>data_in(15));
   ix17124 : inv02 port map ( Y=>nx17125, A=>data_in(15));
   ix17126 : inv02 port map ( Y=>nx17127, A=>data_in(15));
   ix17128 : inv02 port map ( Y=>nx17129, A=>data_in(15));
   ix17130 : inv02 port map ( Y=>nx17131, A=>data_in(15));
   ix17132 : inv02 port map ( Y=>nx17133, A=>data_in(15));
   ix17134 : inv02 port map ( Y=>nx17135, A=>data_in(15));
   ix17136 : inv02 port map ( Y=>nx17137, A=>data_in(15));
   ix17138 : inv02 port map ( Y=>nx17139, A=>data_in(15));
   ix17140 : buf02 port map ( Y=>nx17141, A=>nx14);
   ix17142 : inv04 port map ( Y=>nx17143, A=>nx98);
   ix17146 : inv02 port map ( Y=>nx17147, A=>nx17301);
   ix17152 : nand02 port map ( Y=>nx17153, A0=>address(4), A1=>address(5));
   ix17154 : nand02 port map ( Y=>nx17155, A0=>address(4), A1=>address(5));
   ix17156 : nand02 port map ( Y=>nx17157, A0=>nx10523, A1=>address(5));
   ix17158 : nand02 port map ( Y=>nx17159, A0=>nx10523, A1=>address(5));
   ix880 : mux21 port map ( Y=>nx879, A0=>nx10497, A1=>nx16123, S0=>nx17295
   );
   ix870 : mux21 port map ( Y=>nx869, A0=>nx16123, A1=>nx10529, S0=>nx17289
   );
   ix850 : mux21 port map ( Y=>nx849, A0=>nx16123, A1=>nx10548, S0=>nx17277
   );
   ix860 : mux21 port map ( Y=>nx859, A0=>nx16123, A1=>nx10559, S0=>nx17283
   );
   ix830 : mux21 port map ( Y=>nx829, A0=>nx10574, A1=>nx16123, S0=>nx17305
   );
   ix1211 : nor02_2x port map ( Y=>nx16091, A0=>nx17165, A1=>nx18926);
   ix17164 : inv01 port map ( Y=>nx17165, A=>nx16163);
   ix840 : mux21 port map ( Y=>nx839, A0=>nx10584, A1=>nx16123, S0=>nx17311
   );
   ix820 : mux21 port map ( Y=>nx819, A0=>nx10595, A1=>nx16123, S0=>nx17317
   );
   ix10602 : nor03_2x port map ( Y=>nx16257, A0=>nx17301, A1=>nx17165, A2=>
      nx18927);
   ix810 : mux21 port map ( Y=>nx809, A0=>nx10603, A1=>nx16125, S0=>nx17323
   );
   ix800 : mux21 port map ( Y=>nx799, A0=>nx16125, A1=>nx10619, S0=>nx17271
   );
   ix790 : mux21 port map ( Y=>nx789, A0=>nx10629, A1=>nx16125, S0=>nx17329
   );
   ix770 : mux21 port map ( Y=>nx769, A0=>nx10637, A1=>nx16125, S0=>nx17335
   );
   ix780 : mux21 port map ( Y=>nx779, A0=>nx10645, A1=>nx16125, S0=>nx17341
   );
   ix760 : mux21 port map ( Y=>nx759, A0=>nx10654, A1=>nx16125, S0=>nx17347
   );
   ix750 : mux21 port map ( Y=>nx749, A0=>nx16125, A1=>nx10666, S0=>nx17265
   );
   ix730 : mux21 port map ( Y=>nx729, A0=>nx10674, A1=>nx16127, S0=>nx17353
   );
   ix740 : mux21 port map ( Y=>nx739, A0=>nx10681, A1=>nx16127, S0=>nx17359
   );
   ix720 : mux21 port map ( Y=>nx719, A0=>nx16127, A1=>nx10692, S0=>nx17259
   );
   ix710 : mux21 port map ( Y=>nx709, A0=>nx10699, A1=>nx16127, S0=>nx17365
   );
   ix690 : mux21 port map ( Y=>nx689, A0=>nx16127, A1=>nx10706, S0=>nx17253
   );
   ix700 : mux21 port map ( Y=>nx699, A0=>nx10713, A1=>nx16127, S0=>nx17371
   );
   ix680 : mux21 port map ( Y=>nx679, A0=>nx10724, A1=>nx16127, S0=>nx17377
   );
   ix670 : mux21 port map ( Y=>nx669, A0=>nx10731, A1=>nx16129, S0=>nx17383
   );
   ix650 : mux21 port map ( Y=>nx649, A0=>nx16129, A1=>nx10744, S0=>nx17247
   );
   ix660 : mux21 port map ( Y=>nx659, A0=>nx10751, A1=>nx16129, S0=>nx17389
   );
   ix640 : mux21 port map ( Y=>nx639, A0=>nx10762, A1=>nx16129, S0=>nx17395
   );
   ix630 : mux21 port map ( Y=>nx629, A0=>nx10769, A1=>nx16129, S0=>nx17401
   );
   ix610 : mux21 port map ( Y=>nx609, A0=>nx16129, A1=>nx10783, S0=>nx17241
   );
   ix620 : mux21 port map ( Y=>nx619, A0=>nx10789, A1=>nx16129, S0=>nx17407
   );
   ix600 : mux21 port map ( Y=>nx599, A0=>nx10801, A1=>nx16131, S0=>nx17413
   );
   ix590 : mux21 port map ( Y=>nx589, A0=>nx10807, A1=>nx16131, S0=>nx17419
   );
   ix570 : mux21 port map ( Y=>nx569, A0=>nx16131, A1=>nx10817, S0=>nx17235
   );
   ix580 : mux21 port map ( Y=>nx579, A0=>nx10825, A1=>nx16131, S0=>nx17425
   );
   ix550 : mux21 port map ( Y=>nx549, A0=>nx10841, A1=>nx16131, S0=>nx17431
   );
   ix560 : mux21 port map ( Y=>nx559, A0=>nx16131, A1=>nx10852, S0=>nx17229
   );
   ix540 : mux21 port map ( Y=>nx539, A0=>nx16131, A1=>nx10861, S0=>nx17223
   );
   ix530 : mux21 port map ( Y=>nx529, A0=>nx10869, A1=>nx16133, S0=>nx17437
   );
   ix520 : mux21 port map ( Y=>nx519, A0=>nx10884, A1=>nx16133, S0=>nx17443
   );
   ix510 : mux21 port map ( Y=>nx509, A0=>nx16133, A1=>nx10893, S0=>nx17217
   );
   ix500 : mux21 port map ( Y=>nx499, A0=>nx10903, A1=>nx16133, S0=>nx17451
   );
   ix10906 : nor03_2x port map ( Y=>nx16557, A0=>nx17457, A1=>nx10514, A2=>
      nx218);
   ix490 : mux21 port map ( Y=>nx489, A0=>nx16133, A1=>nx10913, S0=>nx17211
   );
   ix480 : mux21 port map ( Y=>nx479, A0=>nx10922, A1=>nx16133, S0=>nx17463
   );
   ix10926 : nor02_2x port map ( Y=>nx16577, A0=>nx17457, A1=>nx17167);
   ix17166 : inv01 port map ( Y=>nx17167, A=>nx15455);
   ix470 : mux21 port map ( Y=>nx469, A0=>nx10928, A1=>nx16133, S0=>nx17469
   );
   ix460 : mux21 port map ( Y=>nx459, A0=>nx10935, A1=>nx16135, S0=>nx17475
   );
   ix450 : mux21 port map ( Y=>nx449, A0=>nx10943, A1=>nx16135, S0=>nx17483
   );
   ix10948 : nor03_2x port map ( Y=>nx16609, A0=>nx17459, A1=>nx10514, A2=>
      nx17169);
   ix17168 : inv01 port map ( Y=>nx17169, A=>nx16283);
   ix440 : mux21 port map ( Y=>nx439, A0=>nx16135, A1=>nx10954, S0=>nx17205
   );
   ix430 : mux21 port map ( Y=>nx429, A0=>nx10959, A1=>nx16135, S0=>nx17489
   );
   ix420 : mux21 port map ( Y=>nx419, A0=>nx10965, A1=>nx16135, S0=>nx17495
   );
   ix410 : mux21 port map ( Y=>nx409, A0=>nx10972, A1=>nx16135, S0=>nx17501
   );
   ix390 : mux21 port map ( Y=>nx389, A0=>nx10983, A1=>nx16135, S0=>nx17507
   );
   ix400 : mux21 port map ( Y=>nx399, A0=>nx10992, A1=>nx16137, S0=>nx17513
   );
   ix380 : mux21 port map ( Y=>nx379, A0=>nx11000, A1=>nx16137, S0=>nx17519
   );
   ix11006 : nor03_2x port map ( Y=>nx16705, A0=>nx218, A1=>nx17171, A2=>
      nx17173);
   ix17170 : inv01 port map ( Y=>nx17171, A=>nx16165);
   ix17172 : inv01 port map ( Y=>nx17173, A=>nx10663);
   ix370 : mux21 port map ( Y=>nx369, A0=>nx11007, A1=>nx16137, S0=>nx17525
   );
   ix11015 : nor03_2x port map ( Y=>nx16721, A0=>nx17303, A1=>nx17171, A2=>
      nx17173);
   ix360 : mux21 port map ( Y=>nx359, A0=>nx11019, A1=>nx16137, S0=>nx17531
   );
   ix350 : mux21 port map ( Y=>nx349, A0=>nx16137, A1=>nx11026, S0=>nx17199
   );
   ix340 : mux21 port map ( Y=>nx339, A0=>nx11032, A1=>nx16137, S0=>nx17537
   );
   ix330 : mux21 port map ( Y=>nx329, A0=>nx16137, A1=>nx11041, S0=>nx17193
   );
   ix11047 : nor03_2x port map ( Y=>nx16753, A0=>nx218, A1=>nx17175, A2=>
      nx122);
   ix17174 : inv01 port map ( Y=>nx17175, A=>nx16169);
   ix320 : mux21 port map ( Y=>nx319, A0=>nx11051, A1=>nx16139, S0=>nx17543
   );
   ix310 : mux21 port map ( Y=>nx309, A0=>nx16139, A1=>nx11059, S0=>nx17187
   );
   ix300 : mux21 port map ( Y=>nx299, A0=>nx16139, A1=>nx11064, S0=>nx17181
   );
   ix11069 : nor03_2x port map ( Y=>nx16769, A0=>nx17303, A1=>nx17175, A2=>
      nx122);
   ix290 : mux21 port map ( Y=>nx289, A0=>nx11070, A1=>nx16139, S0=>nx17549
   );
   ix280 : mux21 port map ( Y=>nx279, A0=>nx11080, A1=>nx16139, S0=>nx17555
   );
   ix270 : mux21 port map ( Y=>nx269, A0=>nx11086, A1=>nx16139, S0=>nx17561
   );
   ix250 : mux21 port map ( Y=>nx249, A0=>nx11092, A1=>nx16139, S0=>nx17567
   );
   ix260 : mux21 port map ( Y=>nx259, A0=>nx11099, A1=>nx16141, S0=>nx17573
   );
   ix1520 : mux21 port map ( Y=>nx1519, A0=>nx11113, A1=>nx16841, S0=>
      nx17295);
   ix1510 : mux21 port map ( Y=>nx1509, A0=>nx16841, A1=>nx11118, S0=>
      nx17289);
   ix1490 : mux21 port map ( Y=>nx1489, A0=>nx16841, A1=>nx11122, S0=>
      nx17277);
   ix1500 : mux21 port map ( Y=>nx1499, A0=>nx16841, A1=>nx11125, S0=>
      nx17283);
   ix1470 : mux21 port map ( Y=>nx1469, A0=>nx11131, A1=>nx16841, S0=>
      nx17305);
   ix1480 : mux21 port map ( Y=>nx1479, A0=>nx11134, A1=>nx16841, S0=>
      nx17311);
   ix1460 : mux21 port map ( Y=>nx1459, A0=>nx11138, A1=>nx16841, S0=>
      nx17317);
   ix1450 : mux21 port map ( Y=>nx1449, A0=>nx11141, A1=>nx16843, S0=>
      nx17323);
   ix1440 : mux21 port map ( Y=>nx1439, A0=>nx16843, A1=>nx11147, S0=>
      nx17271);
   ix1430 : mux21 port map ( Y=>nx1429, A0=>nx11151, A1=>nx16843, S0=>
      nx17329);
   ix1410 : mux21 port map ( Y=>nx1409, A0=>nx11155, A1=>nx16843, S0=>
      nx17335);
   ix1420 : mux21 port map ( Y=>nx1419, A0=>nx11158, A1=>nx16843, S0=>
      nx17341);
   ix1400 : mux21 port map ( Y=>nx1399, A0=>nx11164, A1=>nx16843, S0=>
      nx17347);
   ix1390 : mux21 port map ( Y=>nx1389, A0=>nx16843, A1=>nx11168, S0=>
      nx17265);
   ix1370 : mux21 port map ( Y=>nx1369, A0=>nx11172, A1=>nx16845, S0=>
      nx17353);
   ix1380 : mux21 port map ( Y=>nx1379, A0=>nx11175, A1=>nx16845, S0=>
      nx17359);
   ix1360 : mux21 port map ( Y=>nx1359, A0=>nx16845, A1=>nx11182, S0=>
      nx17259);
   ix1350 : mux21 port map ( Y=>nx1349, A0=>nx11186, A1=>nx16845, S0=>
      nx17365);
   ix1330 : mux21 port map ( Y=>nx1329, A0=>nx16845, A1=>nx11190, S0=>
      nx17253);
   ix1340 : mux21 port map ( Y=>nx1339, A0=>nx11193, A1=>nx16845, S0=>
      nx17371);
   ix1320 : mux21 port map ( Y=>nx1319, A0=>nx11199, A1=>nx16845, S0=>
      nx17377);
   ix1310 : mux21 port map ( Y=>nx1309, A0=>nx11203, A1=>nx16847, S0=>
      nx17383);
   ix1290 : mux21 port map ( Y=>nx1289, A0=>nx16847, A1=>nx11207, S0=>
      nx17247);
   ix1300 : mux21 port map ( Y=>nx1299, A0=>nx11210, A1=>nx16847, S0=>
      nx17389);
   ix1280 : mux21 port map ( Y=>nx1279, A0=>nx11216, A1=>nx16847, S0=>
      nx17395);
   ix1270 : mux21 port map ( Y=>nx1269, A0=>nx11220, A1=>nx16847, S0=>
      nx17401);
   ix1250 : mux21 port map ( Y=>nx1249, A0=>nx16847, A1=>nx11224, S0=>
      nx17241);
   ix1260 : mux21 port map ( Y=>nx1259, A0=>nx11227, A1=>nx16847, S0=>
      nx17407);
   ix1240 : mux21 port map ( Y=>nx1239, A0=>nx11233, A1=>nx16849, S0=>
      nx17413);
   ix1230 : mux21 port map ( Y=>nx1229, A0=>nx11237, A1=>nx16849, S0=>
      nx17419);
   ix1210 : mux21 port map ( Y=>nx1209, A0=>nx16849, A1=>nx11241, S0=>
      nx17235);
   ix1220 : mux21 port map ( Y=>nx1219, A0=>nx11244, A1=>nx16849, S0=>
      nx17425);
   ix1190 : mux21 port map ( Y=>nx1189, A0=>nx11254, A1=>nx16849, S0=>
      nx17431);
   ix1200 : mux21 port map ( Y=>nx1199, A0=>nx16849, A1=>nx11257, S0=>
      nx17229);
   ix1180 : mux21 port map ( Y=>nx1179, A0=>nx16849, A1=>nx11261, S0=>
      nx17223);
   ix1170 : mux21 port map ( Y=>nx1169, A0=>nx11264, A1=>nx16851, S0=>
      nx17437);
   ix1160 : mux21 port map ( Y=>nx1159, A0=>nx11271, A1=>nx16851, S0=>
      nx17443);
   ix1150 : mux21 port map ( Y=>nx1149, A0=>nx16851, A1=>nx11275, S0=>
      nx17217);
   ix1140 : mux21 port map ( Y=>nx1139, A0=>nx11282, A1=>nx16851, S0=>
      nx17451);
   ix1130 : mux21 port map ( Y=>nx1129, A0=>nx16851, A1=>nx11288, S0=>
      nx17211);
   ix1120 : mux21 port map ( Y=>nx1119, A0=>nx11293, A1=>nx16851, S0=>
      nx17463);
   ix1110 : mux21 port map ( Y=>nx1109, A0=>nx11297, A1=>nx16851, S0=>
      nx17469);
   ix1100 : mux21 port map ( Y=>nx1099, A0=>nx11301, A1=>nx16853, S0=>
      nx17475);
   ix1090 : mux21 port map ( Y=>nx1089, A0=>nx11304, A1=>nx16853, S0=>
      nx17483);
   ix1080 : mux21 port map ( Y=>nx1079, A0=>nx16853, A1=>nx11310, S0=>
      nx17205);
   ix1070 : mux21 port map ( Y=>nx1069, A0=>nx11314, A1=>nx16853, S0=>
      nx17489);
   ix1060 : mux21 port map ( Y=>nx1059, A0=>nx11318, A1=>nx16853, S0=>
      nx17495);
   ix1050 : mux21 port map ( Y=>nx1049, A0=>nx11321, A1=>nx16853, S0=>
      nx17501);
   ix1030 : mux21 port map ( Y=>nx1029, A0=>nx11328, A1=>nx16853, S0=>
      nx17507);
   ix1040 : mux21 port map ( Y=>nx1039, A0=>nx11331, A1=>nx16855, S0=>
      nx17513);
   ix1020 : mux21 port map ( Y=>nx1019, A0=>nx11335, A1=>nx16855, S0=>
      nx17519);
   ix1010 : mux21 port map ( Y=>nx1009, A0=>nx11338, A1=>nx16855, S0=>
      nx17525);
   ix1000 : mux21 port map ( Y=>nx999, A0=>nx11344, A1=>nx16855, S0=>nx17531
   );
   ix990 : mux21 port map ( Y=>nx989, A0=>nx16855, A1=>nx11348, S0=>nx17199
   );
   ix980 : mux21 port map ( Y=>nx979, A0=>nx11352, A1=>nx16855, S0=>nx17537
   );
   ix970 : mux21 port map ( Y=>nx969, A0=>nx16855, A1=>nx11355, S0=>nx17193
   );
   ix960 : mux21 port map ( Y=>nx959, A0=>nx11361, A1=>nx16857, S0=>nx17543
   );
   ix950 : mux21 port map ( Y=>nx949, A0=>nx16857, A1=>nx11365, S0=>nx17187
   );
   ix940 : mux21 port map ( Y=>nx939, A0=>nx16857, A1=>nx11369, S0=>nx17181
   );
   ix930 : mux21 port map ( Y=>nx929, A0=>nx11372, A1=>nx16857, S0=>nx17549
   );
   ix920 : mux21 port map ( Y=>nx919, A0=>nx11378, A1=>nx16857, S0=>nx17555
   );
   ix910 : mux21 port map ( Y=>nx909, A0=>nx11382, A1=>nx16857, S0=>nx17561
   );
   ix890 : mux21 port map ( Y=>nx889, A0=>nx11386, A1=>nx16857, S0=>nx17567
   );
   ix900 : mux21 port map ( Y=>nx899, A0=>nx11389, A1=>nx16859, S0=>nx17573
   );
   ix2160 : mux21 port map ( Y=>nx2159, A0=>nx11399, A1=>nx16861, S0=>
      nx17295);
   ix2150 : mux21 port map ( Y=>nx2149, A0=>nx16861, A1=>nx11404, S0=>
      nx17289);
   ix2130 : mux21 port map ( Y=>nx2129, A0=>nx16861, A1=>nx11408, S0=>
      nx17277);
   ix2140 : mux21 port map ( Y=>nx2139, A0=>nx16861, A1=>nx11411, S0=>
      nx17283);
   ix2110 : mux21 port map ( Y=>nx2109, A0=>nx11417, A1=>nx16861, S0=>
      nx17305);
   ix2120 : mux21 port map ( Y=>nx2119, A0=>nx11420, A1=>nx16861, S0=>
      nx17311);
   ix2100 : mux21 port map ( Y=>nx2099, A0=>nx11424, A1=>nx16861, S0=>
      nx17317);
   ix2090 : mux21 port map ( Y=>nx2089, A0=>nx11427, A1=>nx16863, S0=>
      nx17323);
   ix2080 : mux21 port map ( Y=>nx2079, A0=>nx16863, A1=>nx11433, S0=>
      nx17271);
   ix2070 : mux21 port map ( Y=>nx2069, A0=>nx11437, A1=>nx16863, S0=>
      nx17329);
   ix2050 : mux21 port map ( Y=>nx2049, A0=>nx11441, A1=>nx16863, S0=>
      nx17335);
   ix2060 : mux21 port map ( Y=>nx2059, A0=>nx11444, A1=>nx16863, S0=>
      nx17341);
   ix2040 : mux21 port map ( Y=>nx2039, A0=>nx11450, A1=>nx16863, S0=>
      nx17347);
   ix2030 : mux21 port map ( Y=>nx2029, A0=>nx16863, A1=>nx11454, S0=>
      nx17265);
   ix2010 : mux21 port map ( Y=>nx2009, A0=>nx11458, A1=>nx16865, S0=>
      nx17353);
   ix2020 : mux21 port map ( Y=>nx2019, A0=>nx11461, A1=>nx16865, S0=>
      nx17359);
   ix2000 : mux21 port map ( Y=>nx1999, A0=>nx16865, A1=>nx11468, S0=>
      nx17259);
   ix1990 : mux21 port map ( Y=>nx1989, A0=>nx11472, A1=>nx16865, S0=>
      nx17365);
   ix1970 : mux21 port map ( Y=>nx1969, A0=>nx16865, A1=>nx11476, S0=>
      nx17253);
   ix1980 : mux21 port map ( Y=>nx1979, A0=>nx11479, A1=>nx16865, S0=>
      nx17371);
   ix1960 : mux21 port map ( Y=>nx1959, A0=>nx11485, A1=>nx16865, S0=>
      nx17377);
   ix1950 : mux21 port map ( Y=>nx1949, A0=>nx11489, A1=>nx16867, S0=>
      nx17383);
   ix1930 : mux21 port map ( Y=>nx1929, A0=>nx16867, A1=>nx11493, S0=>
      nx17247);
   ix1940 : mux21 port map ( Y=>nx1939, A0=>nx11496, A1=>nx16867, S0=>
      nx17389);
   ix1920 : mux21 port map ( Y=>nx1919, A0=>nx11502, A1=>nx16867, S0=>
      nx17395);
   ix1910 : mux21 port map ( Y=>nx1909, A0=>nx11506, A1=>nx16867, S0=>
      nx17401);
   ix1890 : mux21 port map ( Y=>nx1889, A0=>nx16867, A1=>nx11510, S0=>
      nx17241);
   ix1900 : mux21 port map ( Y=>nx1899, A0=>nx11513, A1=>nx16867, S0=>
      nx17407);
   ix1880 : mux21 port map ( Y=>nx1879, A0=>nx11519, A1=>nx16869, S0=>
      nx17413);
   ix1870 : mux21 port map ( Y=>nx1869, A0=>nx11523, A1=>nx16869, S0=>
      nx17419);
   ix1850 : mux21 port map ( Y=>nx1849, A0=>nx16869, A1=>nx11527, S0=>
      nx17235);
   ix1860 : mux21 port map ( Y=>nx1859, A0=>nx11530, A1=>nx16869, S0=>
      nx17425);
   ix1830 : mux21 port map ( Y=>nx1829, A0=>nx11540, A1=>nx16869, S0=>
      nx17431);
   ix1840 : mux21 port map ( Y=>nx1839, A0=>nx16869, A1=>nx11543, S0=>
      nx17229);
   ix1820 : mux21 port map ( Y=>nx1819, A0=>nx16869, A1=>nx11547, S0=>
      nx17223);
   ix1810 : mux21 port map ( Y=>nx1809, A0=>nx11550, A1=>nx16871, S0=>
      nx17437);
   ix1800 : mux21 port map ( Y=>nx1799, A0=>nx11557, A1=>nx16871, S0=>
      nx17443);
   ix1790 : mux21 port map ( Y=>nx1789, A0=>nx16871, A1=>nx11561, S0=>
      nx17217);
   ix1780 : mux21 port map ( Y=>nx1779, A0=>nx11568, A1=>nx16871, S0=>
      nx17451);
   ix1770 : mux21 port map ( Y=>nx1769, A0=>nx16871, A1=>nx11574, S0=>
      nx17211);
   ix1760 : mux21 port map ( Y=>nx1759, A0=>nx11579, A1=>nx16871, S0=>
      nx17463);
   ix1750 : mux21 port map ( Y=>nx1749, A0=>nx11583, A1=>nx16871, S0=>
      nx17469);
   ix1740 : mux21 port map ( Y=>nx1739, A0=>nx11587, A1=>nx16873, S0=>
      nx17475);
   ix1730 : mux21 port map ( Y=>nx1729, A0=>nx11590, A1=>nx16873, S0=>
      nx17483);
   ix1720 : mux21 port map ( Y=>nx1719, A0=>nx16873, A1=>nx11596, S0=>
      nx17205);
   ix1710 : mux21 port map ( Y=>nx1709, A0=>nx11600, A1=>nx16873, S0=>
      nx17489);
   ix1700 : mux21 port map ( Y=>nx1699, A0=>nx11604, A1=>nx16873, S0=>
      nx17495);
   ix1690 : mux21 port map ( Y=>nx1689, A0=>nx11607, A1=>nx16873, S0=>
      nx17501);
   ix1670 : mux21 port map ( Y=>nx1669, A0=>nx11614, A1=>nx16873, S0=>
      nx17507);
   ix1680 : mux21 port map ( Y=>nx1679, A0=>nx11617, A1=>nx16875, S0=>
      nx17513);
   ix1660 : mux21 port map ( Y=>nx1659, A0=>nx11621, A1=>nx16875, S0=>
      nx17519);
   ix1650 : mux21 port map ( Y=>nx1649, A0=>nx11624, A1=>nx16875, S0=>
      nx17525);
   ix1640 : mux21 port map ( Y=>nx1639, A0=>nx11630, A1=>nx16875, S0=>
      nx17531);
   ix1630 : mux21 port map ( Y=>nx1629, A0=>nx16875, A1=>nx11634, S0=>
      nx17199);
   ix1620 : mux21 port map ( Y=>nx1619, A0=>nx11638, A1=>nx16875, S0=>
      nx17537);
   ix1610 : mux21 port map ( Y=>nx1609, A0=>nx16875, A1=>nx11641, S0=>
      nx17193);
   ix1600 : mux21 port map ( Y=>nx1599, A0=>nx11647, A1=>nx16877, S0=>
      nx17543);
   ix1590 : mux21 port map ( Y=>nx1589, A0=>nx16877, A1=>nx11651, S0=>
      nx17187);
   ix1580 : mux21 port map ( Y=>nx1579, A0=>nx16877, A1=>nx11655, S0=>
      nx17181);
   ix1570 : mux21 port map ( Y=>nx1569, A0=>nx11658, A1=>nx16877, S0=>
      nx17549);
   ix1560 : mux21 port map ( Y=>nx1559, A0=>nx11664, A1=>nx16877, S0=>
      nx17555);
   ix1550 : mux21 port map ( Y=>nx1549, A0=>nx11668, A1=>nx16877, S0=>
      nx17561);
   ix1530 : mux21 port map ( Y=>nx1529, A0=>nx11672, A1=>nx16877, S0=>
      nx17567);
   ix1540 : mux21 port map ( Y=>nx1539, A0=>nx11675, A1=>nx16879, S0=>
      nx17573);
   ix2800 : mux21 port map ( Y=>nx2799, A0=>nx11685, A1=>nx16881, S0=>
      nx17295);
   ix2790 : mux21 port map ( Y=>nx2789, A0=>nx16881, A1=>nx11690, S0=>
      nx17289);
   ix2770 : mux21 port map ( Y=>nx2769, A0=>nx16881, A1=>nx11694, S0=>
      nx17277);
   ix2780 : mux21 port map ( Y=>nx2779, A0=>nx16881, A1=>nx11697, S0=>
      nx17283);
   ix2750 : mux21 port map ( Y=>nx2749, A0=>nx11703, A1=>nx16881, S0=>
      nx17305);
   ix2760 : mux21 port map ( Y=>nx2759, A0=>nx11706, A1=>nx16881, S0=>
      nx17311);
   ix2740 : mux21 port map ( Y=>nx2739, A0=>nx11710, A1=>nx16881, S0=>
      nx17317);
   ix2730 : mux21 port map ( Y=>nx2729, A0=>nx11713, A1=>nx16883, S0=>
      nx17323);
   ix2720 : mux21 port map ( Y=>nx2719, A0=>nx16883, A1=>nx11719, S0=>
      nx17271);
   ix2710 : mux21 port map ( Y=>nx2709, A0=>nx11723, A1=>nx16883, S0=>
      nx17329);
   ix2690 : mux21 port map ( Y=>nx2689, A0=>nx11727, A1=>nx16883, S0=>
      nx17335);
   ix2700 : mux21 port map ( Y=>nx2699, A0=>nx11730, A1=>nx16883, S0=>
      nx17341);
   ix2680 : mux21 port map ( Y=>nx2679, A0=>nx11736, A1=>nx16883, S0=>
      nx17347);
   ix2670 : mux21 port map ( Y=>nx2669, A0=>nx16883, A1=>nx11740, S0=>
      nx17265);
   ix2650 : mux21 port map ( Y=>nx2649, A0=>nx11744, A1=>nx16885, S0=>
      nx17353);
   ix2660 : mux21 port map ( Y=>nx2659, A0=>nx11747, A1=>nx16885, S0=>
      nx17359);
   ix2640 : mux21 port map ( Y=>nx2639, A0=>nx16885, A1=>nx11754, S0=>
      nx17259);
   ix2630 : mux21 port map ( Y=>nx2629, A0=>nx11758, A1=>nx16885, S0=>
      nx17365);
   ix2610 : mux21 port map ( Y=>nx2609, A0=>nx16885, A1=>nx11762, S0=>
      nx17253);
   ix2620 : mux21 port map ( Y=>nx2619, A0=>nx11765, A1=>nx16885, S0=>
      nx17371);
   ix2600 : mux21 port map ( Y=>nx2599, A0=>nx11771, A1=>nx16885, S0=>
      nx17377);
   ix2590 : mux21 port map ( Y=>nx2589, A0=>nx11775, A1=>nx16887, S0=>
      nx17383);
   ix2570 : mux21 port map ( Y=>nx2569, A0=>nx16887, A1=>nx11779, S0=>
      nx17247);
   ix2580 : mux21 port map ( Y=>nx2579, A0=>nx11782, A1=>nx16887, S0=>
      nx17389);
   ix2560 : mux21 port map ( Y=>nx2559, A0=>nx11788, A1=>nx16887, S0=>
      nx17395);
   ix2550 : mux21 port map ( Y=>nx2549, A0=>nx11792, A1=>nx16887, S0=>
      nx17401);
   ix2530 : mux21 port map ( Y=>nx2529, A0=>nx16887, A1=>nx11796, S0=>
      nx17241);
   ix2540 : mux21 port map ( Y=>nx2539, A0=>nx11799, A1=>nx16887, S0=>
      nx17407);
   ix2520 : mux21 port map ( Y=>nx2519, A0=>nx11805, A1=>nx16889, S0=>
      nx17413);
   ix2510 : mux21 port map ( Y=>nx2509, A0=>nx11809, A1=>nx16889, S0=>
      nx17419);
   ix2490 : mux21 port map ( Y=>nx2489, A0=>nx16889, A1=>nx11813, S0=>
      nx17235);
   ix2500 : mux21 port map ( Y=>nx2499, A0=>nx11816, A1=>nx16889, S0=>
      nx17425);
   ix2470 : mux21 port map ( Y=>nx2469, A0=>nx11826, A1=>nx16889, S0=>
      nx17431);
   ix2480 : mux21 port map ( Y=>nx2479, A0=>nx16889, A1=>nx11829, S0=>
      nx17229);
   ix2460 : mux21 port map ( Y=>nx2459, A0=>nx16889, A1=>nx11833, S0=>
      nx17223);
   ix2450 : mux21 port map ( Y=>nx2449, A0=>nx11836, A1=>nx16891, S0=>
      nx17437);
   ix2440 : mux21 port map ( Y=>nx2439, A0=>nx11843, A1=>nx16891, S0=>
      nx17443);
   ix2430 : mux21 port map ( Y=>nx2429, A0=>nx16891, A1=>nx11847, S0=>
      nx17217);
   ix2420 : mux21 port map ( Y=>nx2419, A0=>nx11854, A1=>nx16891, S0=>
      nx17451);
   ix2410 : mux21 port map ( Y=>nx2409, A0=>nx16891, A1=>nx11860, S0=>
      nx17211);
   ix2400 : mux21 port map ( Y=>nx2399, A0=>nx11865, A1=>nx16891, S0=>
      nx17463);
   ix2390 : mux21 port map ( Y=>nx2389, A0=>nx11869, A1=>nx16891, S0=>
      nx17469);
   ix2380 : mux21 port map ( Y=>nx2379, A0=>nx11873, A1=>nx16893, S0=>
      nx17475);
   ix2370 : mux21 port map ( Y=>nx2369, A0=>nx11876, A1=>nx16893, S0=>
      nx17483);
   ix2360 : mux21 port map ( Y=>nx2359, A0=>nx16893, A1=>nx11882, S0=>
      nx17205);
   ix2350 : mux21 port map ( Y=>nx2349, A0=>nx11886, A1=>nx16893, S0=>
      nx17489);
   ix2340 : mux21 port map ( Y=>nx2339, A0=>nx11890, A1=>nx16893, S0=>
      nx17495);
   ix2330 : mux21 port map ( Y=>nx2329, A0=>nx11893, A1=>nx16893, S0=>
      nx17501);
   ix2310 : mux21 port map ( Y=>nx2309, A0=>nx11900, A1=>nx16893, S0=>
      nx17507);
   ix2320 : mux21 port map ( Y=>nx2319, A0=>nx11903, A1=>nx16895, S0=>
      nx17513);
   ix2300 : mux21 port map ( Y=>nx2299, A0=>nx11907, A1=>nx16895, S0=>
      nx17519);
   ix2290 : mux21 port map ( Y=>nx2289, A0=>nx11910, A1=>nx16895, S0=>
      nx17525);
   ix2280 : mux21 port map ( Y=>nx2279, A0=>nx11916, A1=>nx16895, S0=>
      nx17531);
   ix2270 : mux21 port map ( Y=>nx2269, A0=>nx16895, A1=>nx11920, S0=>
      nx17199);
   ix2260 : mux21 port map ( Y=>nx2259, A0=>nx11924, A1=>nx16895, S0=>
      nx17537);
   ix2250 : mux21 port map ( Y=>nx2249, A0=>nx16895, A1=>nx11927, S0=>
      nx17193);
   ix2240 : mux21 port map ( Y=>nx2239, A0=>nx11933, A1=>nx16897, S0=>
      nx17543);
   ix2230 : mux21 port map ( Y=>nx2229, A0=>nx16897, A1=>nx11937, S0=>
      nx17187);
   ix2220 : mux21 port map ( Y=>nx2219, A0=>nx16897, A1=>nx11941, S0=>
      nx17181);
   ix2210 : mux21 port map ( Y=>nx2209, A0=>nx11944, A1=>nx16897, S0=>
      nx17549);
   ix2200 : mux21 port map ( Y=>nx2199, A0=>nx11950, A1=>nx16897, S0=>
      nx17555);
   ix2190 : mux21 port map ( Y=>nx2189, A0=>nx11954, A1=>nx16897, S0=>
      nx17561);
   ix2170 : mux21 port map ( Y=>nx2169, A0=>nx11958, A1=>nx16897, S0=>
      nx17567);
   ix2180 : mux21 port map ( Y=>nx2179, A0=>nx11961, A1=>nx16899, S0=>
      nx17573);
   ix3440 : mux21 port map ( Y=>nx3439, A0=>nx11971, A1=>nx16901, S0=>
      nx17295);
   ix3430 : mux21 port map ( Y=>nx3429, A0=>nx16901, A1=>nx11976, S0=>
      nx17289);
   ix3410 : mux21 port map ( Y=>nx3409, A0=>nx16901, A1=>nx11980, S0=>
      nx17277);
   ix3420 : mux21 port map ( Y=>nx3419, A0=>nx16901, A1=>nx11983, S0=>
      nx17283);
   ix3390 : mux21 port map ( Y=>nx3389, A0=>nx11989, A1=>nx16901, S0=>
      nx17305);
   ix3400 : mux21 port map ( Y=>nx3399, A0=>nx11992, A1=>nx16901, S0=>
      nx17311);
   ix3380 : mux21 port map ( Y=>nx3379, A0=>nx11996, A1=>nx16901, S0=>
      nx17317);
   ix3370 : mux21 port map ( Y=>nx3369, A0=>nx11999, A1=>nx16903, S0=>
      nx17323);
   ix3360 : mux21 port map ( Y=>nx3359, A0=>nx16903, A1=>nx12005, S0=>
      nx17271);
   ix3350 : mux21 port map ( Y=>nx3349, A0=>nx12009, A1=>nx16903, S0=>
      nx17329);
   ix3330 : mux21 port map ( Y=>nx3329, A0=>nx12013, A1=>nx16903, S0=>
      nx17335);
   ix3340 : mux21 port map ( Y=>nx3339, A0=>nx12016, A1=>nx16903, S0=>
      nx17341);
   ix3320 : mux21 port map ( Y=>nx3319, A0=>nx12022, A1=>nx16903, S0=>
      nx17347);
   ix3310 : mux21 port map ( Y=>nx3309, A0=>nx16903, A1=>nx12026, S0=>
      nx17265);
   ix3290 : mux21 port map ( Y=>nx3289, A0=>nx12030, A1=>nx16905, S0=>
      nx17353);
   ix3300 : mux21 port map ( Y=>nx3299, A0=>nx12033, A1=>nx16905, S0=>
      nx17359);
   ix3280 : mux21 port map ( Y=>nx3279, A0=>nx16905, A1=>nx12040, S0=>
      nx17259);
   ix3270 : mux21 port map ( Y=>nx3269, A0=>nx12044, A1=>nx16905, S0=>
      nx17365);
   ix3250 : mux21 port map ( Y=>nx3249, A0=>nx16905, A1=>nx12048, S0=>
      nx17253);
   ix3260 : mux21 port map ( Y=>nx3259, A0=>nx12051, A1=>nx16905, S0=>
      nx17371);
   ix3240 : mux21 port map ( Y=>nx3239, A0=>nx12057, A1=>nx16905, S0=>
      nx17377);
   ix3230 : mux21 port map ( Y=>nx3229, A0=>nx12061, A1=>nx16907, S0=>
      nx17383);
   ix3210 : mux21 port map ( Y=>nx3209, A0=>nx16907, A1=>nx12065, S0=>
      nx17247);
   ix3220 : mux21 port map ( Y=>nx3219, A0=>nx12068, A1=>nx16907, S0=>
      nx17389);
   ix3200 : mux21 port map ( Y=>nx3199, A0=>nx12074, A1=>nx16907, S0=>
      nx17395);
   ix3190 : mux21 port map ( Y=>nx3189, A0=>nx12078, A1=>nx16907, S0=>
      nx17401);
   ix3170 : mux21 port map ( Y=>nx3169, A0=>nx16907, A1=>nx12082, S0=>
      nx17241);
   ix3180 : mux21 port map ( Y=>nx3179, A0=>nx12085, A1=>nx16907, S0=>
      nx17407);
   ix3160 : mux21 port map ( Y=>nx3159, A0=>nx12091, A1=>nx16909, S0=>
      nx17413);
   ix3150 : mux21 port map ( Y=>nx3149, A0=>nx12095, A1=>nx16909, S0=>
      nx17419);
   ix3130 : mux21 port map ( Y=>nx3129, A0=>nx16909, A1=>nx12099, S0=>
      nx17235);
   ix3140 : mux21 port map ( Y=>nx3139, A0=>nx12102, A1=>nx16909, S0=>
      nx17425);
   ix3110 : mux21 port map ( Y=>nx3109, A0=>nx12112, A1=>nx16909, S0=>
      nx17431);
   ix3120 : mux21 port map ( Y=>nx3119, A0=>nx16909, A1=>nx12115, S0=>
      nx17229);
   ix3100 : mux21 port map ( Y=>nx3099, A0=>nx16909, A1=>nx12119, S0=>
      nx17223);
   ix3090 : mux21 port map ( Y=>nx3089, A0=>nx12122, A1=>nx16911, S0=>
      nx17437);
   ix3080 : mux21 port map ( Y=>nx3079, A0=>nx12129, A1=>nx16911, S0=>
      nx17443);
   ix3070 : mux21 port map ( Y=>nx3069, A0=>nx16911, A1=>nx12133, S0=>
      nx17217);
   ix3060 : mux21 port map ( Y=>nx3059, A0=>nx12140, A1=>nx16911, S0=>
      nx17451);
   ix3050 : mux21 port map ( Y=>nx3049, A0=>nx16911, A1=>nx12146, S0=>
      nx17211);
   ix3040 : mux21 port map ( Y=>nx3039, A0=>nx12151, A1=>nx16911, S0=>
      nx17463);
   ix3030 : mux21 port map ( Y=>nx3029, A0=>nx12155, A1=>nx16911, S0=>
      nx17469);
   ix3020 : mux21 port map ( Y=>nx3019, A0=>nx12159, A1=>nx16913, S0=>
      nx17475);
   ix3010 : mux21 port map ( Y=>nx3009, A0=>nx12162, A1=>nx16913, S0=>
      nx17483);
   ix3000 : mux21 port map ( Y=>nx2999, A0=>nx16913, A1=>nx12168, S0=>
      nx17205);
   ix2990 : mux21 port map ( Y=>nx2989, A0=>nx12172, A1=>nx16913, S0=>
      nx17489);
   ix2980 : mux21 port map ( Y=>nx2979, A0=>nx12176, A1=>nx16913, S0=>
      nx17495);
   ix2970 : mux21 port map ( Y=>nx2969, A0=>nx12179, A1=>nx16913, S0=>
      nx17501);
   ix2950 : mux21 port map ( Y=>nx2949, A0=>nx12186, A1=>nx16913, S0=>
      nx17507);
   ix2960 : mux21 port map ( Y=>nx2959, A0=>nx12189, A1=>nx16915, S0=>
      nx17513);
   ix2940 : mux21 port map ( Y=>nx2939, A0=>nx12193, A1=>nx16915, S0=>
      nx17519);
   ix2930 : mux21 port map ( Y=>nx2929, A0=>nx12196, A1=>nx16915, S0=>
      nx17525);
   ix2920 : mux21 port map ( Y=>nx2919, A0=>nx12202, A1=>nx16915, S0=>
      nx17531);
   ix2910 : mux21 port map ( Y=>nx2909, A0=>nx16915, A1=>nx12206, S0=>
      nx17199);
   ix2900 : mux21 port map ( Y=>nx2899, A0=>nx12210, A1=>nx16915, S0=>
      nx17537);
   ix2890 : mux21 port map ( Y=>nx2889, A0=>nx16915, A1=>nx12213, S0=>
      nx17193);
   ix2880 : mux21 port map ( Y=>nx2879, A0=>nx12219, A1=>nx16917, S0=>
      nx17543);
   ix2870 : mux21 port map ( Y=>nx2869, A0=>nx16917, A1=>nx12223, S0=>
      nx17187);
   ix2860 : mux21 port map ( Y=>nx2859, A0=>nx16917, A1=>nx12227, S0=>
      nx17181);
   ix2850 : mux21 port map ( Y=>nx2849, A0=>nx12230, A1=>nx16917, S0=>
      nx17549);
   ix2840 : mux21 port map ( Y=>nx2839, A0=>nx12236, A1=>nx16917, S0=>
      nx17555);
   ix2830 : mux21 port map ( Y=>nx2829, A0=>nx12240, A1=>nx16917, S0=>
      nx17561);
   ix2810 : mux21 port map ( Y=>nx2809, A0=>nx12244, A1=>nx16917, S0=>
      nx17567);
   ix2820 : mux21 port map ( Y=>nx2819, A0=>nx12247, A1=>nx16919, S0=>
      nx17573);
   ix4080 : mux21 port map ( Y=>nx4079, A0=>nx12257, A1=>nx16921, S0=>
      nx17295);
   ix4070 : mux21 port map ( Y=>nx4069, A0=>nx16921, A1=>nx12262, S0=>
      nx17289);
   ix4050 : mux21 port map ( Y=>nx4049, A0=>nx16921, A1=>nx12266, S0=>
      nx17277);
   ix4060 : mux21 port map ( Y=>nx4059, A0=>nx16921, A1=>nx12269, S0=>
      nx17283);
   ix4030 : mux21 port map ( Y=>nx4029, A0=>nx12275, A1=>nx16921, S0=>
      nx17305);
   ix4040 : mux21 port map ( Y=>nx4039, A0=>nx12278, A1=>nx16921, S0=>
      nx17311);
   ix4020 : mux21 port map ( Y=>nx4019, A0=>nx12282, A1=>nx16921, S0=>
      nx17317);
   ix4010 : mux21 port map ( Y=>nx4009, A0=>nx12285, A1=>nx16923, S0=>
      nx17323);
   ix4000 : mux21 port map ( Y=>nx3999, A0=>nx16923, A1=>nx12291, S0=>
      nx17271);
   ix3990 : mux21 port map ( Y=>nx3989, A0=>nx12295, A1=>nx16923, S0=>
      nx17329);
   ix3970 : mux21 port map ( Y=>nx3969, A0=>nx12299, A1=>nx16923, S0=>
      nx17335);
   ix3980 : mux21 port map ( Y=>nx3979, A0=>nx12302, A1=>nx16923, S0=>
      nx17341);
   ix3960 : mux21 port map ( Y=>nx3959, A0=>nx12308, A1=>nx16923, S0=>
      nx17347);
   ix3950 : mux21 port map ( Y=>nx3949, A0=>nx16923, A1=>nx12312, S0=>
      nx17265);
   ix3930 : mux21 port map ( Y=>nx3929, A0=>nx12316, A1=>nx16925, S0=>
      nx17353);
   ix3940 : mux21 port map ( Y=>nx3939, A0=>nx12319, A1=>nx16925, S0=>
      nx17359);
   ix3920 : mux21 port map ( Y=>nx3919, A0=>nx16925, A1=>nx12326, S0=>
      nx17259);
   ix3910 : mux21 port map ( Y=>nx3909, A0=>nx12330, A1=>nx16925, S0=>
      nx17365);
   ix3890 : mux21 port map ( Y=>nx3889, A0=>nx16925, A1=>nx12334, S0=>
      nx17253);
   ix3900 : mux21 port map ( Y=>nx3899, A0=>nx12337, A1=>nx16925, S0=>
      nx17371);
   ix3880 : mux21 port map ( Y=>nx3879, A0=>nx12343, A1=>nx16925, S0=>
      nx17377);
   ix3870 : mux21 port map ( Y=>nx3869, A0=>nx12347, A1=>nx16927, S0=>
      nx17383);
   ix3850 : mux21 port map ( Y=>nx3849, A0=>nx16927, A1=>nx12351, S0=>
      nx17247);
   ix3860 : mux21 port map ( Y=>nx3859, A0=>nx12354, A1=>nx16927, S0=>
      nx17389);
   ix3840 : mux21 port map ( Y=>nx3839, A0=>nx12360, A1=>nx16927, S0=>
      nx17395);
   ix3830 : mux21 port map ( Y=>nx3829, A0=>nx12364, A1=>nx16927, S0=>
      nx17401);
   ix3810 : mux21 port map ( Y=>nx3809, A0=>nx16927, A1=>nx12368, S0=>
      nx17241);
   ix3820 : mux21 port map ( Y=>nx3819, A0=>nx12371, A1=>nx16927, S0=>
      nx17407);
   ix3800 : mux21 port map ( Y=>nx3799, A0=>nx12377, A1=>nx16929, S0=>
      nx17413);
   ix3790 : mux21 port map ( Y=>nx3789, A0=>nx12381, A1=>nx16929, S0=>
      nx17419);
   ix3770 : mux21 port map ( Y=>nx3769, A0=>nx16929, A1=>nx12385, S0=>
      nx17235);
   ix3780 : mux21 port map ( Y=>nx3779, A0=>nx12388, A1=>nx16929, S0=>
      nx17425);
   ix3750 : mux21 port map ( Y=>nx3749, A0=>nx12398, A1=>nx16929, S0=>
      nx17431);
   ix3760 : mux21 port map ( Y=>nx3759, A0=>nx16929, A1=>nx12401, S0=>
      nx17229);
   ix3740 : mux21 port map ( Y=>nx3739, A0=>nx16929, A1=>nx12405, S0=>
      nx17223);
   ix3730 : mux21 port map ( Y=>nx3729, A0=>nx12408, A1=>nx16931, S0=>
      nx17437);
   ix3720 : mux21 port map ( Y=>nx3719, A0=>nx12415, A1=>nx16931, S0=>
      nx17443);
   ix3710 : mux21 port map ( Y=>nx3709, A0=>nx16931, A1=>nx12419, S0=>
      nx17217);
   ix3700 : mux21 port map ( Y=>nx3699, A0=>nx12426, A1=>nx16931, S0=>
      nx17451);
   ix3690 : mux21 port map ( Y=>nx3689, A0=>nx16931, A1=>nx12432, S0=>
      nx17211);
   ix3680 : mux21 port map ( Y=>nx3679, A0=>nx12437, A1=>nx16931, S0=>
      nx17463);
   ix3670 : mux21 port map ( Y=>nx3669, A0=>nx12441, A1=>nx16931, S0=>
      nx17469);
   ix3660 : mux21 port map ( Y=>nx3659, A0=>nx12445, A1=>nx16933, S0=>
      nx17475);
   ix3650 : mux21 port map ( Y=>nx3649, A0=>nx12448, A1=>nx16933, S0=>
      nx17483);
   ix3640 : mux21 port map ( Y=>nx3639, A0=>nx16933, A1=>nx12454, S0=>
      nx17205);
   ix3630 : mux21 port map ( Y=>nx3629, A0=>nx12458, A1=>nx16933, S0=>
      nx17489);
   ix3620 : mux21 port map ( Y=>nx3619, A0=>nx12462, A1=>nx16933, S0=>
      nx17495);
   ix3610 : mux21 port map ( Y=>nx3609, A0=>nx12465, A1=>nx16933, S0=>
      nx17501);
   ix3590 : mux21 port map ( Y=>nx3589, A0=>nx12472, A1=>nx16933, S0=>
      nx17507);
   ix3600 : mux21 port map ( Y=>nx3599, A0=>nx12475, A1=>nx16935, S0=>
      nx17513);
   ix3580 : mux21 port map ( Y=>nx3579, A0=>nx12479, A1=>nx16935, S0=>
      nx17519);
   ix3570 : mux21 port map ( Y=>nx3569, A0=>nx12482, A1=>nx16935, S0=>
      nx17525);
   ix3560 : mux21 port map ( Y=>nx3559, A0=>nx12488, A1=>nx16935, S0=>
      nx17531);
   ix3550 : mux21 port map ( Y=>nx3549, A0=>nx16935, A1=>nx12492, S0=>
      nx17199);
   ix3540 : mux21 port map ( Y=>nx3539, A0=>nx12496, A1=>nx16935, S0=>
      nx17537);
   ix3530 : mux21 port map ( Y=>nx3529, A0=>nx16935, A1=>nx12499, S0=>
      nx17193);
   ix3520 : mux21 port map ( Y=>nx3519, A0=>nx12505, A1=>nx16937, S0=>
      nx17543);
   ix3510 : mux21 port map ( Y=>nx3509, A0=>nx16937, A1=>nx12509, S0=>
      nx17187);
   ix3500 : mux21 port map ( Y=>nx3499, A0=>nx16937, A1=>nx12513, S0=>
      nx17181);
   ix3490 : mux21 port map ( Y=>nx3489, A0=>nx12516, A1=>nx16937, S0=>
      nx17549);
   ix3480 : mux21 port map ( Y=>nx3479, A0=>nx12522, A1=>nx16937, S0=>
      nx17555);
   ix3470 : mux21 port map ( Y=>nx3469, A0=>nx12526, A1=>nx16937, S0=>
      nx17561);
   ix3450 : mux21 port map ( Y=>nx3449, A0=>nx12530, A1=>nx16937, S0=>
      nx17567);
   ix3460 : mux21 port map ( Y=>nx3459, A0=>nx12533, A1=>nx16939, S0=>
      nx17573);
   ix4720 : mux21 port map ( Y=>nx4719, A0=>nx12543, A1=>nx16941, S0=>
      nx17295);
   ix4710 : mux21 port map ( Y=>nx4709, A0=>nx16941, A1=>nx12548, S0=>
      nx17289);
   ix4690 : mux21 port map ( Y=>nx4689, A0=>nx16941, A1=>nx12552, S0=>
      nx17277);
   ix4700 : mux21 port map ( Y=>nx4699, A0=>nx16941, A1=>nx12555, S0=>
      nx17283);
   ix4670 : mux21 port map ( Y=>nx4669, A0=>nx12561, A1=>nx16941, S0=>
      nx17305);
   ix4680 : mux21 port map ( Y=>nx4679, A0=>nx12564, A1=>nx16941, S0=>
      nx17311);
   ix4660 : mux21 port map ( Y=>nx4659, A0=>nx12568, A1=>nx16941, S0=>
      nx17317);
   ix4650 : mux21 port map ( Y=>nx4649, A0=>nx12571, A1=>nx16943, S0=>
      nx17323);
   ix4640 : mux21 port map ( Y=>nx4639, A0=>nx16943, A1=>nx12577, S0=>
      nx17271);
   ix4630 : mux21 port map ( Y=>nx4629, A0=>nx12581, A1=>nx16943, S0=>
      nx17329);
   ix4610 : mux21 port map ( Y=>nx4609, A0=>nx12585, A1=>nx16943, S0=>
      nx17335);
   ix4620 : mux21 port map ( Y=>nx4619, A0=>nx12588, A1=>nx16943, S0=>
      nx17341);
   ix4600 : mux21 port map ( Y=>nx4599, A0=>nx12594, A1=>nx16943, S0=>
      nx17347);
   ix4590 : mux21 port map ( Y=>nx4589, A0=>nx16943, A1=>nx12598, S0=>
      nx17265);
   ix4570 : mux21 port map ( Y=>nx4569, A0=>nx12602, A1=>nx16945, S0=>
      nx17353);
   ix4580 : mux21 port map ( Y=>nx4579, A0=>nx12605, A1=>nx16945, S0=>
      nx17359);
   ix4560 : mux21 port map ( Y=>nx4559, A0=>nx16945, A1=>nx12612, S0=>
      nx17259);
   ix4550 : mux21 port map ( Y=>nx4549, A0=>nx12616, A1=>nx16945, S0=>
      nx17365);
   ix4530 : mux21 port map ( Y=>nx4529, A0=>nx16945, A1=>nx12620, S0=>
      nx17253);
   ix4540 : mux21 port map ( Y=>nx4539, A0=>nx12623, A1=>nx16945, S0=>
      nx17371);
   ix4520 : mux21 port map ( Y=>nx4519, A0=>nx12629, A1=>nx16945, S0=>
      nx17377);
   ix4510 : mux21 port map ( Y=>nx4509, A0=>nx12633, A1=>nx16947, S0=>
      nx17383);
   ix4490 : mux21 port map ( Y=>nx4489, A0=>nx16947, A1=>nx12637, S0=>
      nx17247);
   ix4500 : mux21 port map ( Y=>nx4499, A0=>nx12640, A1=>nx16947, S0=>
      nx17389);
   ix4480 : mux21 port map ( Y=>nx4479, A0=>nx12646, A1=>nx16947, S0=>
      nx17395);
   ix4470 : mux21 port map ( Y=>nx4469, A0=>nx12650, A1=>nx16947, S0=>
      nx17401);
   ix4450 : mux21 port map ( Y=>nx4449, A0=>nx16947, A1=>nx12654, S0=>
      nx17241);
   ix4460 : mux21 port map ( Y=>nx4459, A0=>nx12657, A1=>nx16947, S0=>
      nx17407);
   ix4440 : mux21 port map ( Y=>nx4439, A0=>nx12663, A1=>nx16949, S0=>
      nx17413);
   ix4430 : mux21 port map ( Y=>nx4429, A0=>nx12667, A1=>nx16949, S0=>
      nx17419);
   ix4410 : mux21 port map ( Y=>nx4409, A0=>nx16949, A1=>nx12671, S0=>
      nx17235);
   ix4420 : mux21 port map ( Y=>nx4419, A0=>nx12674, A1=>nx16949, S0=>
      nx17425);
   ix4390 : mux21 port map ( Y=>nx4389, A0=>nx12684, A1=>nx16949, S0=>
      nx17431);
   ix4400 : mux21 port map ( Y=>nx4399, A0=>nx16949, A1=>nx12687, S0=>
      nx17229);
   ix4380 : mux21 port map ( Y=>nx4379, A0=>nx16949, A1=>nx12691, S0=>
      nx17223);
   ix4370 : mux21 port map ( Y=>nx4369, A0=>nx12694, A1=>nx16951, S0=>
      nx17437);
   ix4360 : mux21 port map ( Y=>nx4359, A0=>nx12701, A1=>nx16951, S0=>
      nx17443);
   ix4350 : mux21 port map ( Y=>nx4349, A0=>nx16951, A1=>nx12705, S0=>
      nx17217);
   ix4340 : mux21 port map ( Y=>nx4339, A0=>nx12712, A1=>nx16951, S0=>
      nx17451);
   ix4330 : mux21 port map ( Y=>nx4329, A0=>nx16951, A1=>nx12718, S0=>
      nx17211);
   ix4320 : mux21 port map ( Y=>nx4319, A0=>nx12723, A1=>nx16951, S0=>
      nx17463);
   ix4310 : mux21 port map ( Y=>nx4309, A0=>nx12727, A1=>nx16951, S0=>
      nx17469);
   ix4300 : mux21 port map ( Y=>nx4299, A0=>nx12731, A1=>nx16953, S0=>
      nx17475);
   ix4290 : mux21 port map ( Y=>nx4289, A0=>nx12734, A1=>nx16953, S0=>
      nx17483);
   ix4280 : mux21 port map ( Y=>nx4279, A0=>nx16953, A1=>nx12740, S0=>
      nx17205);
   ix4270 : mux21 port map ( Y=>nx4269, A0=>nx12744, A1=>nx16953, S0=>
      nx17489);
   ix4260 : mux21 port map ( Y=>nx4259, A0=>nx12748, A1=>nx16953, S0=>
      nx17495);
   ix4250 : mux21 port map ( Y=>nx4249, A0=>nx12751, A1=>nx16953, S0=>
      nx17501);
   ix4230 : mux21 port map ( Y=>nx4229, A0=>nx12758, A1=>nx16953, S0=>
      nx17507);
   ix4240 : mux21 port map ( Y=>nx4239, A0=>nx12761, A1=>nx16955, S0=>
      nx17513);
   ix4220 : mux21 port map ( Y=>nx4219, A0=>nx12765, A1=>nx16955, S0=>
      nx17519);
   ix4210 : mux21 port map ( Y=>nx4209, A0=>nx12768, A1=>nx16955, S0=>
      nx17525);
   ix4200 : mux21 port map ( Y=>nx4199, A0=>nx12774, A1=>nx16955, S0=>
      nx17531);
   ix4190 : mux21 port map ( Y=>nx4189, A0=>nx16955, A1=>nx12778, S0=>
      nx17199);
   ix4180 : mux21 port map ( Y=>nx4179, A0=>nx12782, A1=>nx16955, S0=>
      nx17537);
   ix4170 : mux21 port map ( Y=>nx4169, A0=>nx16955, A1=>nx12785, S0=>
      nx17193);
   ix4160 : mux21 port map ( Y=>nx4159, A0=>nx12791, A1=>nx16957, S0=>
      nx17543);
   ix4150 : mux21 port map ( Y=>nx4149, A0=>nx16957, A1=>nx12795, S0=>
      nx17187);
   ix4140 : mux21 port map ( Y=>nx4139, A0=>nx16957, A1=>nx12799, S0=>
      nx17181);
   ix4130 : mux21 port map ( Y=>nx4129, A0=>nx12802, A1=>nx16957, S0=>
      nx17549);
   ix4120 : mux21 port map ( Y=>nx4119, A0=>nx12808, A1=>nx16957, S0=>
      nx17555);
   ix4110 : mux21 port map ( Y=>nx4109, A0=>nx12812, A1=>nx16957, S0=>
      nx17561);
   ix4090 : mux21 port map ( Y=>nx4089, A0=>nx12816, A1=>nx16957, S0=>
      nx17567);
   ix4100 : mux21 port map ( Y=>nx4099, A0=>nx12819, A1=>nx16959, S0=>
      nx17573);
   ix5360 : mux21 port map ( Y=>nx5359, A0=>nx12829, A1=>nx16961, S0=>
      nx17297);
   ix5350 : mux21 port map ( Y=>nx5349, A0=>nx16961, A1=>nx12834, S0=>
      nx17291);
   ix5330 : mux21 port map ( Y=>nx5329, A0=>nx16961, A1=>nx12838, S0=>
      nx17279);
   ix5340 : mux21 port map ( Y=>nx5339, A0=>nx16961, A1=>nx12841, S0=>
      nx17285);
   ix5310 : mux21 port map ( Y=>nx5309, A0=>nx12847, A1=>nx16961, S0=>
      nx17307);
   ix5320 : mux21 port map ( Y=>nx5319, A0=>nx12850, A1=>nx16961, S0=>
      nx17313);
   ix5300 : mux21 port map ( Y=>nx5299, A0=>nx12854, A1=>nx16961, S0=>
      nx17319);
   ix5290 : mux21 port map ( Y=>nx5289, A0=>nx12857, A1=>nx16963, S0=>
      nx17325);
   ix5280 : mux21 port map ( Y=>nx5279, A0=>nx16963, A1=>nx12863, S0=>
      nx17273);
   ix5270 : mux21 port map ( Y=>nx5269, A0=>nx12867, A1=>nx16963, S0=>
      nx17331);
   ix5250 : mux21 port map ( Y=>nx5249, A0=>nx12871, A1=>nx16963, S0=>
      nx17337);
   ix5260 : mux21 port map ( Y=>nx5259, A0=>nx12874, A1=>nx16963, S0=>
      nx17343);
   ix5240 : mux21 port map ( Y=>nx5239, A0=>nx12880, A1=>nx16963, S0=>
      nx17349);
   ix5230 : mux21 port map ( Y=>nx5229, A0=>nx16963, A1=>nx12884, S0=>
      nx17267);
   ix5210 : mux21 port map ( Y=>nx5209, A0=>nx12888, A1=>nx16965, S0=>
      nx17355);
   ix5220 : mux21 port map ( Y=>nx5219, A0=>nx12891, A1=>nx16965, S0=>
      nx17361);
   ix5200 : mux21 port map ( Y=>nx5199, A0=>nx16965, A1=>nx12898, S0=>
      nx17261);
   ix5190 : mux21 port map ( Y=>nx5189, A0=>nx12902, A1=>nx16965, S0=>
      nx17367);
   ix5170 : mux21 port map ( Y=>nx5169, A0=>nx16965, A1=>nx12906, S0=>
      nx17255);
   ix5180 : mux21 port map ( Y=>nx5179, A0=>nx12909, A1=>nx16965, S0=>
      nx17373);
   ix5160 : mux21 port map ( Y=>nx5159, A0=>nx12915, A1=>nx16965, S0=>
      nx17379);
   ix5150 : mux21 port map ( Y=>nx5149, A0=>nx12919, A1=>nx16967, S0=>
      nx17385);
   ix5130 : mux21 port map ( Y=>nx5129, A0=>nx16967, A1=>nx12923, S0=>
      nx17249);
   ix5140 : mux21 port map ( Y=>nx5139, A0=>nx12926, A1=>nx16967, S0=>
      nx17391);
   ix5120 : mux21 port map ( Y=>nx5119, A0=>nx12932, A1=>nx16967, S0=>
      nx17397);
   ix5110 : mux21 port map ( Y=>nx5109, A0=>nx12936, A1=>nx16967, S0=>
      nx17403);
   ix5090 : mux21 port map ( Y=>nx5089, A0=>nx16967, A1=>nx12940, S0=>
      nx17243);
   ix5100 : mux21 port map ( Y=>nx5099, A0=>nx12943, A1=>nx16967, S0=>
      nx17409);
   ix5080 : mux21 port map ( Y=>nx5079, A0=>nx12949, A1=>nx16969, S0=>
      nx17415);
   ix5070 : mux21 port map ( Y=>nx5069, A0=>nx12953, A1=>nx16969, S0=>
      nx17421);
   ix5050 : mux21 port map ( Y=>nx5049, A0=>nx16969, A1=>nx12957, S0=>
      nx17237);
   ix5060 : mux21 port map ( Y=>nx5059, A0=>nx12960, A1=>nx16969, S0=>
      nx17427);
   ix5030 : mux21 port map ( Y=>nx5029, A0=>nx12970, A1=>nx16969, S0=>
      nx17433);
   ix5040 : mux21 port map ( Y=>nx5039, A0=>nx16969, A1=>nx12973, S0=>
      nx17231);
   ix5020 : mux21 port map ( Y=>nx5019, A0=>nx16969, A1=>nx12977, S0=>
      nx17225);
   ix5010 : mux21 port map ( Y=>nx5009, A0=>nx12980, A1=>nx16971, S0=>
      nx17439);
   ix5000 : mux21 port map ( Y=>nx4999, A0=>nx12987, A1=>nx16971, S0=>
      nx17445);
   ix4990 : mux21 port map ( Y=>nx4989, A0=>nx16971, A1=>nx12991, S0=>
      nx17219);
   ix4980 : mux21 port map ( Y=>nx4979, A0=>nx12998, A1=>nx16971, S0=>
      nx17453);
   ix4970 : mux21 port map ( Y=>nx4969, A0=>nx16971, A1=>nx13004, S0=>
      nx17213);
   ix4960 : mux21 port map ( Y=>nx4959, A0=>nx13009, A1=>nx16971, S0=>
      nx17465);
   ix4950 : mux21 port map ( Y=>nx4949, A0=>nx13013, A1=>nx16971, S0=>
      nx17471);
   ix4940 : mux21 port map ( Y=>nx4939, A0=>nx13017, A1=>nx16973, S0=>
      nx17477);
   ix4930 : mux21 port map ( Y=>nx4929, A0=>nx13020, A1=>nx16973, S0=>
      nx17485);
   ix4920 : mux21 port map ( Y=>nx4919, A0=>nx16973, A1=>nx13026, S0=>
      nx17207);
   ix4910 : mux21 port map ( Y=>nx4909, A0=>nx13030, A1=>nx16973, S0=>
      nx17491);
   ix4900 : mux21 port map ( Y=>nx4899, A0=>nx13034, A1=>nx16973, S0=>
      nx17497);
   ix4890 : mux21 port map ( Y=>nx4889, A0=>nx13037, A1=>nx16973, S0=>
      nx17503);
   ix4870 : mux21 port map ( Y=>nx4869, A0=>nx13044, A1=>nx16973, S0=>
      nx17509);
   ix4880 : mux21 port map ( Y=>nx4879, A0=>nx13047, A1=>nx16975, S0=>
      nx17515);
   ix4860 : mux21 port map ( Y=>nx4859, A0=>nx13051, A1=>nx16975, S0=>
      nx17521);
   ix4850 : mux21 port map ( Y=>nx4849, A0=>nx13054, A1=>nx16975, S0=>
      nx17527);
   ix4840 : mux21 port map ( Y=>nx4839, A0=>nx13060, A1=>nx16975, S0=>
      nx17533);
   ix4830 : mux21 port map ( Y=>nx4829, A0=>nx16975, A1=>nx13064, S0=>
      nx17201);
   ix4820 : mux21 port map ( Y=>nx4819, A0=>nx13068, A1=>nx16975, S0=>
      nx17539);
   ix4810 : mux21 port map ( Y=>nx4809, A0=>nx16975, A1=>nx13071, S0=>
      nx17195);
   ix4800 : mux21 port map ( Y=>nx4799, A0=>nx13077, A1=>nx16977, S0=>
      nx17545);
   ix4790 : mux21 port map ( Y=>nx4789, A0=>nx16977, A1=>nx13081, S0=>
      nx17189);
   ix4780 : mux21 port map ( Y=>nx4779, A0=>nx16977, A1=>nx13085, S0=>
      nx17183);
   ix4770 : mux21 port map ( Y=>nx4769, A0=>nx13088, A1=>nx16977, S0=>
      nx17551);
   ix4760 : mux21 port map ( Y=>nx4759, A0=>nx13094, A1=>nx16977, S0=>
      nx17557);
   ix4750 : mux21 port map ( Y=>nx4749, A0=>nx13098, A1=>nx16977, S0=>
      nx17563);
   ix4730 : mux21 port map ( Y=>nx4729, A0=>nx13102, A1=>nx16977, S0=>
      nx17569);
   ix4740 : mux21 port map ( Y=>nx4739, A0=>nx13105, A1=>nx16979, S0=>
      nx17575);
   ix6000 : mux21 port map ( Y=>nx5999, A0=>nx13115, A1=>nx16981, S0=>
      nx17297);
   ix5990 : mux21 port map ( Y=>nx5989, A0=>nx16981, A1=>nx13120, S0=>
      nx17291);
   ix5970 : mux21 port map ( Y=>nx5969, A0=>nx16981, A1=>nx13124, S0=>
      nx17279);
   ix5980 : mux21 port map ( Y=>nx5979, A0=>nx16981, A1=>nx13127, S0=>
      nx17285);
   ix5950 : mux21 port map ( Y=>nx5949, A0=>nx13133, A1=>nx16981, S0=>
      nx17307);
   ix5960 : mux21 port map ( Y=>nx5959, A0=>nx13136, A1=>nx16981, S0=>
      nx17313);
   ix5940 : mux21 port map ( Y=>nx5939, A0=>nx13140, A1=>nx16981, S0=>
      nx17319);
   ix5930 : mux21 port map ( Y=>nx5929, A0=>nx13143, A1=>nx16983, S0=>
      nx17325);
   ix5920 : mux21 port map ( Y=>nx5919, A0=>nx16983, A1=>nx13149, S0=>
      nx17273);
   ix5910 : mux21 port map ( Y=>nx5909, A0=>nx13153, A1=>nx16983, S0=>
      nx17331);
   ix5890 : mux21 port map ( Y=>nx5889, A0=>nx13157, A1=>nx16983, S0=>
      nx17337);
   ix5900 : mux21 port map ( Y=>nx5899, A0=>nx13160, A1=>nx16983, S0=>
      nx17343);
   ix5880 : mux21 port map ( Y=>nx5879, A0=>nx13166, A1=>nx16983, S0=>
      nx17349);
   ix5870 : mux21 port map ( Y=>nx5869, A0=>nx16983, A1=>nx13170, S0=>
      nx17267);
   ix5850 : mux21 port map ( Y=>nx5849, A0=>nx13174, A1=>nx16985, S0=>
      nx17355);
   ix5860 : mux21 port map ( Y=>nx5859, A0=>nx13177, A1=>nx16985, S0=>
      nx17361);
   ix5840 : mux21 port map ( Y=>nx5839, A0=>nx16985, A1=>nx13184, S0=>
      nx17261);
   ix5830 : mux21 port map ( Y=>nx5829, A0=>nx13188, A1=>nx16985, S0=>
      nx17367);
   ix5810 : mux21 port map ( Y=>nx5809, A0=>nx16985, A1=>nx13192, S0=>
      nx17255);
   ix5820 : mux21 port map ( Y=>nx5819, A0=>nx13195, A1=>nx16985, S0=>
      nx17373);
   ix5800 : mux21 port map ( Y=>nx5799, A0=>nx13201, A1=>nx16985, S0=>
      nx17379);
   ix5790 : mux21 port map ( Y=>nx5789, A0=>nx13205, A1=>nx16987, S0=>
      nx17385);
   ix5770 : mux21 port map ( Y=>nx5769, A0=>nx16987, A1=>nx13209, S0=>
      nx17249);
   ix5780 : mux21 port map ( Y=>nx5779, A0=>nx13212, A1=>nx16987, S0=>
      nx17391);
   ix5760 : mux21 port map ( Y=>nx5759, A0=>nx13218, A1=>nx16987, S0=>
      nx17397);
   ix5750 : mux21 port map ( Y=>nx5749, A0=>nx13222, A1=>nx16987, S0=>
      nx17403);
   ix5730 : mux21 port map ( Y=>nx5729, A0=>nx16987, A1=>nx13226, S0=>
      nx17243);
   ix5740 : mux21 port map ( Y=>nx5739, A0=>nx13229, A1=>nx16987, S0=>
      nx17409);
   ix5720 : mux21 port map ( Y=>nx5719, A0=>nx13235, A1=>nx16989, S0=>
      nx17415);
   ix5710 : mux21 port map ( Y=>nx5709, A0=>nx13239, A1=>nx16989, S0=>
      nx17421);
   ix5690 : mux21 port map ( Y=>nx5689, A0=>nx16989, A1=>nx13243, S0=>
      nx17237);
   ix5700 : mux21 port map ( Y=>nx5699, A0=>nx13246, A1=>nx16989, S0=>
      nx17427);
   ix5670 : mux21 port map ( Y=>nx5669, A0=>nx13256, A1=>nx16989, S0=>
      nx17433);
   ix5680 : mux21 port map ( Y=>nx5679, A0=>nx16989, A1=>nx13259, S0=>
      nx17231);
   ix5660 : mux21 port map ( Y=>nx5659, A0=>nx16989, A1=>nx13263, S0=>
      nx17225);
   ix5650 : mux21 port map ( Y=>nx5649, A0=>nx13266, A1=>nx16991, S0=>
      nx17439);
   ix5640 : mux21 port map ( Y=>nx5639, A0=>nx13273, A1=>nx16991, S0=>
      nx17445);
   ix5630 : mux21 port map ( Y=>nx5629, A0=>nx16991, A1=>nx13277, S0=>
      nx17219);
   ix5620 : mux21 port map ( Y=>nx5619, A0=>nx13284, A1=>nx16991, S0=>
      nx17453);
   ix5610 : mux21 port map ( Y=>nx5609, A0=>nx16991, A1=>nx13290, S0=>
      nx17213);
   ix5600 : mux21 port map ( Y=>nx5599, A0=>nx13295, A1=>nx16991, S0=>
      nx17465);
   ix5590 : mux21 port map ( Y=>nx5589, A0=>nx13299, A1=>nx16991, S0=>
      nx17471);
   ix5580 : mux21 port map ( Y=>nx5579, A0=>nx13303, A1=>nx16993, S0=>
      nx17477);
   ix5570 : mux21 port map ( Y=>nx5569, A0=>nx13306, A1=>nx16993, S0=>
      nx17485);
   ix5560 : mux21 port map ( Y=>nx5559, A0=>nx16993, A1=>nx13312, S0=>
      nx17207);
   ix5550 : mux21 port map ( Y=>nx5549, A0=>nx13316, A1=>nx16993, S0=>
      nx17491);
   ix5540 : mux21 port map ( Y=>nx5539, A0=>nx13320, A1=>nx16993, S0=>
      nx17497);
   ix5530 : mux21 port map ( Y=>nx5529, A0=>nx13323, A1=>nx16993, S0=>
      nx17503);
   ix5510 : mux21 port map ( Y=>nx5509, A0=>nx13330, A1=>nx16993, S0=>
      nx17509);
   ix5520 : mux21 port map ( Y=>nx5519, A0=>nx13333, A1=>nx16995, S0=>
      nx17515);
   ix5500 : mux21 port map ( Y=>nx5499, A0=>nx13337, A1=>nx16995, S0=>
      nx17521);
   ix5490 : mux21 port map ( Y=>nx5489, A0=>nx13340, A1=>nx16995, S0=>
      nx17527);
   ix5480 : mux21 port map ( Y=>nx5479, A0=>nx13346, A1=>nx16995, S0=>
      nx17533);
   ix5470 : mux21 port map ( Y=>nx5469, A0=>nx16995, A1=>nx13350, S0=>
      nx17201);
   ix5460 : mux21 port map ( Y=>nx5459, A0=>nx13354, A1=>nx16995, S0=>
      nx17539);
   ix5450 : mux21 port map ( Y=>nx5449, A0=>nx16995, A1=>nx13357, S0=>
      nx17195);
   ix5440 : mux21 port map ( Y=>nx5439, A0=>nx13363, A1=>nx16997, S0=>
      nx17545);
   ix5430 : mux21 port map ( Y=>nx5429, A0=>nx16997, A1=>nx13367, S0=>
      nx17189);
   ix5420 : mux21 port map ( Y=>nx5419, A0=>nx16997, A1=>nx13371, S0=>
      nx17183);
   ix5410 : mux21 port map ( Y=>nx5409, A0=>nx13374, A1=>nx16997, S0=>
      nx17551);
   ix5400 : mux21 port map ( Y=>nx5399, A0=>nx13380, A1=>nx16997, S0=>
      nx17557);
   ix5390 : mux21 port map ( Y=>nx5389, A0=>nx13384, A1=>nx16997, S0=>
      nx17563);
   ix5370 : mux21 port map ( Y=>nx5369, A0=>nx13388, A1=>nx16997, S0=>
      nx17569);
   ix5380 : mux21 port map ( Y=>nx5379, A0=>nx13391, A1=>nx16999, S0=>
      nx17575);
   ix6640 : mux21 port map ( Y=>nx6639, A0=>nx13401, A1=>nx17001, S0=>
      nx17297);
   ix6630 : mux21 port map ( Y=>nx6629, A0=>nx17001, A1=>nx13406, S0=>
      nx17291);
   ix6610 : mux21 port map ( Y=>nx6609, A0=>nx17001, A1=>nx13410, S0=>
      nx17279);
   ix6620 : mux21 port map ( Y=>nx6619, A0=>nx17001, A1=>nx13413, S0=>
      nx17285);
   ix6590 : mux21 port map ( Y=>nx6589, A0=>nx13419, A1=>nx17001, S0=>
      nx17307);
   ix6600 : mux21 port map ( Y=>nx6599, A0=>nx13422, A1=>nx17001, S0=>
      nx17313);
   ix6580 : mux21 port map ( Y=>nx6579, A0=>nx13426, A1=>nx17001, S0=>
      nx17319);
   ix6570 : mux21 port map ( Y=>nx6569, A0=>nx13429, A1=>nx17003, S0=>
      nx17325);
   ix6560 : mux21 port map ( Y=>nx6559, A0=>nx17003, A1=>nx13435, S0=>
      nx17273);
   ix6550 : mux21 port map ( Y=>nx6549, A0=>nx13439, A1=>nx17003, S0=>
      nx17331);
   ix6530 : mux21 port map ( Y=>nx6529, A0=>nx13443, A1=>nx17003, S0=>
      nx17337);
   ix6540 : mux21 port map ( Y=>nx6539, A0=>nx13446, A1=>nx17003, S0=>
      nx17343);
   ix6520 : mux21 port map ( Y=>nx6519, A0=>nx13452, A1=>nx17003, S0=>
      nx17349);
   ix6510 : mux21 port map ( Y=>nx6509, A0=>nx17003, A1=>nx13456, S0=>
      nx17267);
   ix6490 : mux21 port map ( Y=>nx6489, A0=>nx13460, A1=>nx17005, S0=>
      nx17355);
   ix6500 : mux21 port map ( Y=>nx6499, A0=>nx13463, A1=>nx17005, S0=>
      nx17361);
   ix6480 : mux21 port map ( Y=>nx6479, A0=>nx17005, A1=>nx13470, S0=>
      nx17261);
   ix6470 : mux21 port map ( Y=>nx6469, A0=>nx13474, A1=>nx17005, S0=>
      nx17367);
   ix6450 : mux21 port map ( Y=>nx6449, A0=>nx17005, A1=>nx13478, S0=>
      nx17255);
   ix6460 : mux21 port map ( Y=>nx6459, A0=>nx13481, A1=>nx17005, S0=>
      nx17373);
   ix6440 : mux21 port map ( Y=>nx6439, A0=>nx13487, A1=>nx17005, S0=>
      nx17379);
   ix6430 : mux21 port map ( Y=>nx6429, A0=>nx13491, A1=>nx17007, S0=>
      nx17385);
   ix6410 : mux21 port map ( Y=>nx6409, A0=>nx17007, A1=>nx13495, S0=>
      nx17249);
   ix6420 : mux21 port map ( Y=>nx6419, A0=>nx13498, A1=>nx17007, S0=>
      nx17391);
   ix6400 : mux21 port map ( Y=>nx6399, A0=>nx13504, A1=>nx17007, S0=>
      nx17397);
   ix6390 : mux21 port map ( Y=>nx6389, A0=>nx13508, A1=>nx17007, S0=>
      nx17403);
   ix6370 : mux21 port map ( Y=>nx6369, A0=>nx17007, A1=>nx13512, S0=>
      nx17243);
   ix6380 : mux21 port map ( Y=>nx6379, A0=>nx13515, A1=>nx17007, S0=>
      nx17409);
   ix6360 : mux21 port map ( Y=>nx6359, A0=>nx13521, A1=>nx17009, S0=>
      nx17415);
   ix6350 : mux21 port map ( Y=>nx6349, A0=>nx13525, A1=>nx17009, S0=>
      nx17421);
   ix6330 : mux21 port map ( Y=>nx6329, A0=>nx17009, A1=>nx13529, S0=>
      nx17237);
   ix6340 : mux21 port map ( Y=>nx6339, A0=>nx13532, A1=>nx17009, S0=>
      nx17427);
   ix6310 : mux21 port map ( Y=>nx6309, A0=>nx13542, A1=>nx17009, S0=>
      nx17433);
   ix6320 : mux21 port map ( Y=>nx6319, A0=>nx17009, A1=>nx13545, S0=>
      nx17231);
   ix6300 : mux21 port map ( Y=>nx6299, A0=>nx17009, A1=>nx13549, S0=>
      nx17225);
   ix6290 : mux21 port map ( Y=>nx6289, A0=>nx13552, A1=>nx17011, S0=>
      nx17439);
   ix6280 : mux21 port map ( Y=>nx6279, A0=>nx13559, A1=>nx17011, S0=>
      nx17445);
   ix6270 : mux21 port map ( Y=>nx6269, A0=>nx17011, A1=>nx13563, S0=>
      nx17219);
   ix6260 : mux21 port map ( Y=>nx6259, A0=>nx13570, A1=>nx17011, S0=>
      nx17453);
   ix6250 : mux21 port map ( Y=>nx6249, A0=>nx17011, A1=>nx13576, S0=>
      nx17213);
   ix6240 : mux21 port map ( Y=>nx6239, A0=>nx13581, A1=>nx17011, S0=>
      nx17465);
   ix6230 : mux21 port map ( Y=>nx6229, A0=>nx13585, A1=>nx17011, S0=>
      nx17471);
   ix6220 : mux21 port map ( Y=>nx6219, A0=>nx13589, A1=>nx17013, S0=>
      nx17477);
   ix6210 : mux21 port map ( Y=>nx6209, A0=>nx13592, A1=>nx17013, S0=>
      nx17485);
   ix6200 : mux21 port map ( Y=>nx6199, A0=>nx17013, A1=>nx13598, S0=>
      nx17207);
   ix6190 : mux21 port map ( Y=>nx6189, A0=>nx13602, A1=>nx17013, S0=>
      nx17491);
   ix6180 : mux21 port map ( Y=>nx6179, A0=>nx13606, A1=>nx17013, S0=>
      nx17497);
   ix6170 : mux21 port map ( Y=>nx6169, A0=>nx13609, A1=>nx17013, S0=>
      nx17503);
   ix6150 : mux21 port map ( Y=>nx6149, A0=>nx13616, A1=>nx17013, S0=>
      nx17509);
   ix6160 : mux21 port map ( Y=>nx6159, A0=>nx13619, A1=>nx17015, S0=>
      nx17515);
   ix6140 : mux21 port map ( Y=>nx6139, A0=>nx13623, A1=>nx17015, S0=>
      nx17521);
   ix6130 : mux21 port map ( Y=>nx6129, A0=>nx13626, A1=>nx17015, S0=>
      nx17527);
   ix6120 : mux21 port map ( Y=>nx6119, A0=>nx13632, A1=>nx17015, S0=>
      nx17533);
   ix6110 : mux21 port map ( Y=>nx6109, A0=>nx17015, A1=>nx13636, S0=>
      nx17201);
   ix6100 : mux21 port map ( Y=>nx6099, A0=>nx13640, A1=>nx17015, S0=>
      nx17539);
   ix6090 : mux21 port map ( Y=>nx6089, A0=>nx17015, A1=>nx13643, S0=>
      nx17195);
   ix6080 : mux21 port map ( Y=>nx6079, A0=>nx13649, A1=>nx17017, S0=>
      nx17545);
   ix6070 : mux21 port map ( Y=>nx6069, A0=>nx17017, A1=>nx13653, S0=>
      nx17189);
   ix6060 : mux21 port map ( Y=>nx6059, A0=>nx17017, A1=>nx13657, S0=>
      nx17183);
   ix6050 : mux21 port map ( Y=>nx6049, A0=>nx13660, A1=>nx17017, S0=>
      nx17551);
   ix6040 : mux21 port map ( Y=>nx6039, A0=>nx13666, A1=>nx17017, S0=>
      nx17557);
   ix6030 : mux21 port map ( Y=>nx6029, A0=>nx13670, A1=>nx17017, S0=>
      nx17563);
   ix6010 : mux21 port map ( Y=>nx6009, A0=>nx13674, A1=>nx17017, S0=>
      nx17569);
   ix6020 : mux21 port map ( Y=>nx6019, A0=>nx13677, A1=>nx17019, S0=>
      nx17575);
   ix7280 : mux21 port map ( Y=>nx7279, A0=>nx13687, A1=>nx17021, S0=>
      nx17297);
   ix7270 : mux21 port map ( Y=>nx7269, A0=>nx17021, A1=>nx13692, S0=>
      nx17291);
   ix7250 : mux21 port map ( Y=>nx7249, A0=>nx17021, A1=>nx13696, S0=>
      nx17279);
   ix7260 : mux21 port map ( Y=>nx7259, A0=>nx17021, A1=>nx13699, S0=>
      nx17285);
   ix7230 : mux21 port map ( Y=>nx7229, A0=>nx13705, A1=>nx17021, S0=>
      nx17307);
   ix7240 : mux21 port map ( Y=>nx7239, A0=>nx13708, A1=>nx17021, S0=>
      nx17313);
   ix7220 : mux21 port map ( Y=>nx7219, A0=>nx13712, A1=>nx17021, S0=>
      nx17319);
   ix7210 : mux21 port map ( Y=>nx7209, A0=>nx13715, A1=>nx17023, S0=>
      nx17325);
   ix7200 : mux21 port map ( Y=>nx7199, A0=>nx17023, A1=>nx13721, S0=>
      nx17273);
   ix7190 : mux21 port map ( Y=>nx7189, A0=>nx13725, A1=>nx17023, S0=>
      nx17331);
   ix7170 : mux21 port map ( Y=>nx7169, A0=>nx13729, A1=>nx17023, S0=>
      nx17337);
   ix7180 : mux21 port map ( Y=>nx7179, A0=>nx13732, A1=>nx17023, S0=>
      nx17343);
   ix7160 : mux21 port map ( Y=>nx7159, A0=>nx13738, A1=>nx17023, S0=>
      nx17349);
   ix7150 : mux21 port map ( Y=>nx7149, A0=>nx17023, A1=>nx13742, S0=>
      nx17267);
   ix7130 : mux21 port map ( Y=>nx7129, A0=>nx13746, A1=>nx17025, S0=>
      nx17355);
   ix7140 : mux21 port map ( Y=>nx7139, A0=>nx13749, A1=>nx17025, S0=>
      nx17361);
   ix7120 : mux21 port map ( Y=>nx7119, A0=>nx17025, A1=>nx13756, S0=>
      nx17261);
   ix7110 : mux21 port map ( Y=>nx7109, A0=>nx13760, A1=>nx17025, S0=>
      nx17367);
   ix7090 : mux21 port map ( Y=>nx7089, A0=>nx17025, A1=>nx13764, S0=>
      nx17255);
   ix7100 : mux21 port map ( Y=>nx7099, A0=>nx13767, A1=>nx17025, S0=>
      nx17373);
   ix7080 : mux21 port map ( Y=>nx7079, A0=>nx13773, A1=>nx17025, S0=>
      nx17379);
   ix7070 : mux21 port map ( Y=>nx7069, A0=>nx13777, A1=>nx17027, S0=>
      nx17385);
   ix7050 : mux21 port map ( Y=>nx7049, A0=>nx17027, A1=>nx13781, S0=>
      nx17249);
   ix7060 : mux21 port map ( Y=>nx7059, A0=>nx13784, A1=>nx17027, S0=>
      nx17391);
   ix7040 : mux21 port map ( Y=>nx7039, A0=>nx13790, A1=>nx17027, S0=>
      nx17397);
   ix7030 : mux21 port map ( Y=>nx7029, A0=>nx13794, A1=>nx17027, S0=>
      nx17403);
   ix7010 : mux21 port map ( Y=>nx7009, A0=>nx17027, A1=>nx13798, S0=>
      nx17243);
   ix7020 : mux21 port map ( Y=>nx7019, A0=>nx13801, A1=>nx17027, S0=>
      nx17409);
   ix7000 : mux21 port map ( Y=>nx6999, A0=>nx13807, A1=>nx17029, S0=>
      nx17415);
   ix6990 : mux21 port map ( Y=>nx6989, A0=>nx13811, A1=>nx17029, S0=>
      nx17421);
   ix6970 : mux21 port map ( Y=>nx6969, A0=>nx17029, A1=>nx13815, S0=>
      nx17237);
   ix6980 : mux21 port map ( Y=>nx6979, A0=>nx13818, A1=>nx17029, S0=>
      nx17427);
   ix6950 : mux21 port map ( Y=>nx6949, A0=>nx13828, A1=>nx17029, S0=>
      nx17433);
   ix6960 : mux21 port map ( Y=>nx6959, A0=>nx17029, A1=>nx13831, S0=>
      nx17231);
   ix6940 : mux21 port map ( Y=>nx6939, A0=>nx17029, A1=>nx13835, S0=>
      nx17225);
   ix6930 : mux21 port map ( Y=>nx6929, A0=>nx13838, A1=>nx17031, S0=>
      nx17439);
   ix6920 : mux21 port map ( Y=>nx6919, A0=>nx13845, A1=>nx17031, S0=>
      nx17445);
   ix6910 : mux21 port map ( Y=>nx6909, A0=>nx17031, A1=>nx13849, S0=>
      nx17219);
   ix6900 : mux21 port map ( Y=>nx6899, A0=>nx13856, A1=>nx17031, S0=>
      nx17453);
   ix6890 : mux21 port map ( Y=>nx6889, A0=>nx17031, A1=>nx13862, S0=>
      nx17213);
   ix6880 : mux21 port map ( Y=>nx6879, A0=>nx13867, A1=>nx17031, S0=>
      nx17465);
   ix6870 : mux21 port map ( Y=>nx6869, A0=>nx13871, A1=>nx17031, S0=>
      nx17471);
   ix6860 : mux21 port map ( Y=>nx6859, A0=>nx13875, A1=>nx17033, S0=>
      nx17477);
   ix6850 : mux21 port map ( Y=>nx6849, A0=>nx13878, A1=>nx17033, S0=>
      nx17485);
   ix6840 : mux21 port map ( Y=>nx6839, A0=>nx17033, A1=>nx13884, S0=>
      nx17207);
   ix6830 : mux21 port map ( Y=>nx6829, A0=>nx13888, A1=>nx17033, S0=>
      nx17491);
   ix6820 : mux21 port map ( Y=>nx6819, A0=>nx13892, A1=>nx17033, S0=>
      nx17497);
   ix6810 : mux21 port map ( Y=>nx6809, A0=>nx13895, A1=>nx17033, S0=>
      nx17503);
   ix6790 : mux21 port map ( Y=>nx6789, A0=>nx13902, A1=>nx17033, S0=>
      nx17509);
   ix6800 : mux21 port map ( Y=>nx6799, A0=>nx13905, A1=>nx17035, S0=>
      nx17515);
   ix6780 : mux21 port map ( Y=>nx6779, A0=>nx13909, A1=>nx17035, S0=>
      nx17521);
   ix6770 : mux21 port map ( Y=>nx6769, A0=>nx13912, A1=>nx17035, S0=>
      nx17527);
   ix6760 : mux21 port map ( Y=>nx6759, A0=>nx13918, A1=>nx17035, S0=>
      nx17533);
   ix6750 : mux21 port map ( Y=>nx6749, A0=>nx17035, A1=>nx13922, S0=>
      nx17201);
   ix6740 : mux21 port map ( Y=>nx6739, A0=>nx13926, A1=>nx17035, S0=>
      nx17539);
   ix6730 : mux21 port map ( Y=>nx6729, A0=>nx17035, A1=>nx13929, S0=>
      nx17195);
   ix6720 : mux21 port map ( Y=>nx6719, A0=>nx13935, A1=>nx17037, S0=>
      nx17545);
   ix6710 : mux21 port map ( Y=>nx6709, A0=>nx17037, A1=>nx13939, S0=>
      nx17189);
   ix6700 : mux21 port map ( Y=>nx6699, A0=>nx17037, A1=>nx13943, S0=>
      nx17183);
   ix6690 : mux21 port map ( Y=>nx6689, A0=>nx13946, A1=>nx17037, S0=>
      nx17551);
   ix6680 : mux21 port map ( Y=>nx6679, A0=>nx13952, A1=>nx17037, S0=>
      nx17557);
   ix6670 : mux21 port map ( Y=>nx6669, A0=>nx13956, A1=>nx17037, S0=>
      nx17563);
   ix6650 : mux21 port map ( Y=>nx6649, A0=>nx13960, A1=>nx17037, S0=>
      nx17569);
   ix6660 : mux21 port map ( Y=>nx6659, A0=>nx13963, A1=>nx17039, S0=>
      nx17575);
   ix7920 : mux21 port map ( Y=>nx7919, A0=>nx13973, A1=>nx17041, S0=>
      nx17297);
   ix7910 : mux21 port map ( Y=>nx7909, A0=>nx17041, A1=>nx13978, S0=>
      nx17291);
   ix7890 : mux21 port map ( Y=>nx7889, A0=>nx17041, A1=>nx13982, S0=>
      nx17279);
   ix7900 : mux21 port map ( Y=>nx7899, A0=>nx17041, A1=>nx13985, S0=>
      nx17285);
   ix7870 : mux21 port map ( Y=>nx7869, A0=>nx13991, A1=>nx17041, S0=>
      nx17307);
   ix7880 : mux21 port map ( Y=>nx7879, A0=>nx13994, A1=>nx17041, S0=>
      nx17313);
   ix7860 : mux21 port map ( Y=>nx7859, A0=>nx13998, A1=>nx17041, S0=>
      nx17319);
   ix7850 : mux21 port map ( Y=>nx7849, A0=>nx14001, A1=>nx17043, S0=>
      nx17325);
   ix7840 : mux21 port map ( Y=>nx7839, A0=>nx17043, A1=>nx14007, S0=>
      nx17273);
   ix7830 : mux21 port map ( Y=>nx7829, A0=>nx14011, A1=>nx17043, S0=>
      nx17331);
   ix7810 : mux21 port map ( Y=>nx7809, A0=>nx14015, A1=>nx17043, S0=>
      nx17337);
   ix7820 : mux21 port map ( Y=>nx7819, A0=>nx14018, A1=>nx17043, S0=>
      nx17343);
   ix7800 : mux21 port map ( Y=>nx7799, A0=>nx14024, A1=>nx17043, S0=>
      nx17349);
   ix7790 : mux21 port map ( Y=>nx7789, A0=>nx17043, A1=>nx14028, S0=>
      nx17267);
   ix7770 : mux21 port map ( Y=>nx7769, A0=>nx14032, A1=>nx17045, S0=>
      nx17355);
   ix7780 : mux21 port map ( Y=>nx7779, A0=>nx14035, A1=>nx17045, S0=>
      nx17361);
   ix7760 : mux21 port map ( Y=>nx7759, A0=>nx17045, A1=>nx14042, S0=>
      nx17261);
   ix7750 : mux21 port map ( Y=>nx7749, A0=>nx14046, A1=>nx17045, S0=>
      nx17367);
   ix7730 : mux21 port map ( Y=>nx7729, A0=>nx17045, A1=>nx14050, S0=>
      nx17255);
   ix7740 : mux21 port map ( Y=>nx7739, A0=>nx14053, A1=>nx17045, S0=>
      nx17373);
   ix7720 : mux21 port map ( Y=>nx7719, A0=>nx14059, A1=>nx17045, S0=>
      nx17379);
   ix7710 : mux21 port map ( Y=>nx7709, A0=>nx14063, A1=>nx17047, S0=>
      nx17385);
   ix7690 : mux21 port map ( Y=>nx7689, A0=>nx17047, A1=>nx14067, S0=>
      nx17249);
   ix7700 : mux21 port map ( Y=>nx7699, A0=>nx14070, A1=>nx17047, S0=>
      nx17391);
   ix7680 : mux21 port map ( Y=>nx7679, A0=>nx14076, A1=>nx17047, S0=>
      nx17397);
   ix7670 : mux21 port map ( Y=>nx7669, A0=>nx14080, A1=>nx17047, S0=>
      nx17403);
   ix7650 : mux21 port map ( Y=>nx7649, A0=>nx17047, A1=>nx14084, S0=>
      nx17243);
   ix7660 : mux21 port map ( Y=>nx7659, A0=>nx14087, A1=>nx17047, S0=>
      nx17409);
   ix7640 : mux21 port map ( Y=>nx7639, A0=>nx14093, A1=>nx17049, S0=>
      nx17415);
   ix7630 : mux21 port map ( Y=>nx7629, A0=>nx14097, A1=>nx17049, S0=>
      nx17421);
   ix7610 : mux21 port map ( Y=>nx7609, A0=>nx17049, A1=>nx14101, S0=>
      nx17237);
   ix7620 : mux21 port map ( Y=>nx7619, A0=>nx14104, A1=>nx17049, S0=>
      nx17427);
   ix7590 : mux21 port map ( Y=>nx7589, A0=>nx14114, A1=>nx17049, S0=>
      nx17433);
   ix7600 : mux21 port map ( Y=>nx7599, A0=>nx17049, A1=>nx14117, S0=>
      nx17231);
   ix7580 : mux21 port map ( Y=>nx7579, A0=>nx17049, A1=>nx14121, S0=>
      nx17225);
   ix7570 : mux21 port map ( Y=>nx7569, A0=>nx14124, A1=>nx17051, S0=>
      nx17439);
   ix7560 : mux21 port map ( Y=>nx7559, A0=>nx14131, A1=>nx17051, S0=>
      nx17445);
   ix7550 : mux21 port map ( Y=>nx7549, A0=>nx17051, A1=>nx14135, S0=>
      nx17219);
   ix7540 : mux21 port map ( Y=>nx7539, A0=>nx14142, A1=>nx17051, S0=>
      nx17453);
   ix7530 : mux21 port map ( Y=>nx7529, A0=>nx17051, A1=>nx14148, S0=>
      nx17213);
   ix7520 : mux21 port map ( Y=>nx7519, A0=>nx14153, A1=>nx17051, S0=>
      nx17465);
   ix7510 : mux21 port map ( Y=>nx7509, A0=>nx14157, A1=>nx17051, S0=>
      nx17471);
   ix7500 : mux21 port map ( Y=>nx7499, A0=>nx14161, A1=>nx17053, S0=>
      nx17477);
   ix7490 : mux21 port map ( Y=>nx7489, A0=>nx14164, A1=>nx17053, S0=>
      nx17485);
   ix7480 : mux21 port map ( Y=>nx7479, A0=>nx17053, A1=>nx14170, S0=>
      nx17207);
   ix7470 : mux21 port map ( Y=>nx7469, A0=>nx14174, A1=>nx17053, S0=>
      nx17491);
   ix7460 : mux21 port map ( Y=>nx7459, A0=>nx14178, A1=>nx17053, S0=>
      nx17497);
   ix7450 : mux21 port map ( Y=>nx7449, A0=>nx14181, A1=>nx17053, S0=>
      nx17503);
   ix7430 : mux21 port map ( Y=>nx7429, A0=>nx14188, A1=>nx17053, S0=>
      nx17509);
   ix7440 : mux21 port map ( Y=>nx7439, A0=>nx14191, A1=>nx17055, S0=>
      nx17515);
   ix7420 : mux21 port map ( Y=>nx7419, A0=>nx14195, A1=>nx17055, S0=>
      nx17521);
   ix7410 : mux21 port map ( Y=>nx7409, A0=>nx14198, A1=>nx17055, S0=>
      nx17527);
   ix7400 : mux21 port map ( Y=>nx7399, A0=>nx14204, A1=>nx17055, S0=>
      nx17533);
   ix7390 : mux21 port map ( Y=>nx7389, A0=>nx17055, A1=>nx14208, S0=>
      nx17201);
   ix7380 : mux21 port map ( Y=>nx7379, A0=>nx14212, A1=>nx17055, S0=>
      nx17539);
   ix7370 : mux21 port map ( Y=>nx7369, A0=>nx17055, A1=>nx14215, S0=>
      nx17195);
   ix7360 : mux21 port map ( Y=>nx7359, A0=>nx14221, A1=>nx17057, S0=>
      nx17545);
   ix7350 : mux21 port map ( Y=>nx7349, A0=>nx17057, A1=>nx14225, S0=>
      nx17189);
   ix7340 : mux21 port map ( Y=>nx7339, A0=>nx17057, A1=>nx14229, S0=>
      nx17183);
   ix7330 : mux21 port map ( Y=>nx7329, A0=>nx14232, A1=>nx17057, S0=>
      nx17551);
   ix7320 : mux21 port map ( Y=>nx7319, A0=>nx14238, A1=>nx17057, S0=>
      nx17557);
   ix7310 : mux21 port map ( Y=>nx7309, A0=>nx14242, A1=>nx17057, S0=>
      nx17563);
   ix7290 : mux21 port map ( Y=>nx7289, A0=>nx14246, A1=>nx17057, S0=>
      nx17569);
   ix7300 : mux21 port map ( Y=>nx7299, A0=>nx14249, A1=>nx17059, S0=>
      nx17575);
   ix8560 : mux21 port map ( Y=>nx8559, A0=>nx14259, A1=>nx17061, S0=>
      nx17297);
   ix8550 : mux21 port map ( Y=>nx8549, A0=>nx17061, A1=>nx14264, S0=>
      nx17291);
   ix8530 : mux21 port map ( Y=>nx8529, A0=>nx17061, A1=>nx14268, S0=>
      nx17279);
   ix8540 : mux21 port map ( Y=>nx8539, A0=>nx17061, A1=>nx14271, S0=>
      nx17285);
   ix8510 : mux21 port map ( Y=>nx8509, A0=>nx14277, A1=>nx17061, S0=>
      nx17307);
   ix8520 : mux21 port map ( Y=>nx8519, A0=>nx14280, A1=>nx17061, S0=>
      nx17313);
   ix8500 : mux21 port map ( Y=>nx8499, A0=>nx14284, A1=>nx17061, S0=>
      nx17319);
   ix8490 : mux21 port map ( Y=>nx8489, A0=>nx14287, A1=>nx17063, S0=>
      nx17325);
   ix8480 : mux21 port map ( Y=>nx8479, A0=>nx17063, A1=>nx14293, S0=>
      nx17273);
   ix8470 : mux21 port map ( Y=>nx8469, A0=>nx14297, A1=>nx17063, S0=>
      nx17331);
   ix8450 : mux21 port map ( Y=>nx8449, A0=>nx14301, A1=>nx17063, S0=>
      nx17337);
   ix8460 : mux21 port map ( Y=>nx8459, A0=>nx14304, A1=>nx17063, S0=>
      nx17343);
   ix8440 : mux21 port map ( Y=>nx8439, A0=>nx14310, A1=>nx17063, S0=>
      nx17349);
   ix8430 : mux21 port map ( Y=>nx8429, A0=>nx17063, A1=>nx14314, S0=>
      nx17267);
   ix8410 : mux21 port map ( Y=>nx8409, A0=>nx14318, A1=>nx17065, S0=>
      nx17355);
   ix8420 : mux21 port map ( Y=>nx8419, A0=>nx14321, A1=>nx17065, S0=>
      nx17361);
   ix8400 : mux21 port map ( Y=>nx8399, A0=>nx17065, A1=>nx14328, S0=>
      nx17261);
   ix8390 : mux21 port map ( Y=>nx8389, A0=>nx14332, A1=>nx17065, S0=>
      nx17367);
   ix8370 : mux21 port map ( Y=>nx8369, A0=>nx17065, A1=>nx14336, S0=>
      nx17255);
   ix8380 : mux21 port map ( Y=>nx8379, A0=>nx14339, A1=>nx17065, S0=>
      nx17373);
   ix8360 : mux21 port map ( Y=>nx8359, A0=>nx14345, A1=>nx17065, S0=>
      nx17379);
   ix8350 : mux21 port map ( Y=>nx8349, A0=>nx14349, A1=>nx17067, S0=>
      nx17385);
   ix8330 : mux21 port map ( Y=>nx8329, A0=>nx17067, A1=>nx14353, S0=>
      nx17249);
   ix8340 : mux21 port map ( Y=>nx8339, A0=>nx14356, A1=>nx17067, S0=>
      nx17391);
   ix8320 : mux21 port map ( Y=>nx8319, A0=>nx14362, A1=>nx17067, S0=>
      nx17397);
   ix8310 : mux21 port map ( Y=>nx8309, A0=>nx14366, A1=>nx17067, S0=>
      nx17403);
   ix8290 : mux21 port map ( Y=>nx8289, A0=>nx17067, A1=>nx14370, S0=>
      nx17243);
   ix8300 : mux21 port map ( Y=>nx8299, A0=>nx14373, A1=>nx17067, S0=>
      nx17409);
   ix8280 : mux21 port map ( Y=>nx8279, A0=>nx14379, A1=>nx17069, S0=>
      nx17415);
   ix8270 : mux21 port map ( Y=>nx8269, A0=>nx14383, A1=>nx17069, S0=>
      nx17421);
   ix8250 : mux21 port map ( Y=>nx8249, A0=>nx17069, A1=>nx14387, S0=>
      nx17237);
   ix8260 : mux21 port map ( Y=>nx8259, A0=>nx14390, A1=>nx17069, S0=>
      nx17427);
   ix8230 : mux21 port map ( Y=>nx8229, A0=>nx14400, A1=>nx17069, S0=>
      nx17433);
   ix8240 : mux21 port map ( Y=>nx8239, A0=>nx17069, A1=>nx14403, S0=>
      nx17231);
   ix8220 : mux21 port map ( Y=>nx8219, A0=>nx17069, A1=>nx14407, S0=>
      nx17225);
   ix8210 : mux21 port map ( Y=>nx8209, A0=>nx14410, A1=>nx17071, S0=>
      nx17439);
   ix8200 : mux21 port map ( Y=>nx8199, A0=>nx14417, A1=>nx17071, S0=>
      nx17445);
   ix8190 : mux21 port map ( Y=>nx8189, A0=>nx17071, A1=>nx14421, S0=>
      nx17219);
   ix8180 : mux21 port map ( Y=>nx8179, A0=>nx14428, A1=>nx17071, S0=>
      nx17453);
   ix8170 : mux21 port map ( Y=>nx8169, A0=>nx17071, A1=>nx14434, S0=>
      nx17213);
   ix8160 : mux21 port map ( Y=>nx8159, A0=>nx14439, A1=>nx17071, S0=>
      nx17465);
   ix8150 : mux21 port map ( Y=>nx8149, A0=>nx14443, A1=>nx17071, S0=>
      nx17471);
   ix8140 : mux21 port map ( Y=>nx8139, A0=>nx14447, A1=>nx17073, S0=>
      nx17477);
   ix8130 : mux21 port map ( Y=>nx8129, A0=>nx14450, A1=>nx17073, S0=>
      nx17485);
   ix8120 : mux21 port map ( Y=>nx8119, A0=>nx17073, A1=>nx14456, S0=>
      nx17207);
   ix8110 : mux21 port map ( Y=>nx8109, A0=>nx14460, A1=>nx17073, S0=>
      nx17491);
   ix8100 : mux21 port map ( Y=>nx8099, A0=>nx14464, A1=>nx17073, S0=>
      nx17497);
   ix8090 : mux21 port map ( Y=>nx8089, A0=>nx14467, A1=>nx17073, S0=>
      nx17503);
   ix8070 : mux21 port map ( Y=>nx8069, A0=>nx14474, A1=>nx17073, S0=>
      nx17509);
   ix8080 : mux21 port map ( Y=>nx8079, A0=>nx14477, A1=>nx17075, S0=>
      nx17515);
   ix8060 : mux21 port map ( Y=>nx8059, A0=>nx14481, A1=>nx17075, S0=>
      nx17521);
   ix8050 : mux21 port map ( Y=>nx8049, A0=>nx14484, A1=>nx17075, S0=>
      nx17527);
   ix8040 : mux21 port map ( Y=>nx8039, A0=>nx14490, A1=>nx17075, S0=>
      nx17533);
   ix8030 : mux21 port map ( Y=>nx8029, A0=>nx17075, A1=>nx14494, S0=>
      nx17201);
   ix8020 : mux21 port map ( Y=>nx8019, A0=>nx14498, A1=>nx17075, S0=>
      nx17539);
   ix8010 : mux21 port map ( Y=>nx8009, A0=>nx17075, A1=>nx14501, S0=>
      nx17195);
   ix8000 : mux21 port map ( Y=>nx7999, A0=>nx14507, A1=>nx17077, S0=>
      nx17545);
   ix7990 : mux21 port map ( Y=>nx7989, A0=>nx17077, A1=>nx14511, S0=>
      nx17189);
   ix7980 : mux21 port map ( Y=>nx7979, A0=>nx17077, A1=>nx14515, S0=>
      nx17183);
   ix7970 : mux21 port map ( Y=>nx7969, A0=>nx14518, A1=>nx17077, S0=>
      nx17551);
   ix7960 : mux21 port map ( Y=>nx7959, A0=>nx14524, A1=>nx17077, S0=>
      nx17557);
   ix7950 : mux21 port map ( Y=>nx7949, A0=>nx14528, A1=>nx17077, S0=>
      nx17563);
   ix7930 : mux21 port map ( Y=>nx7929, A0=>nx14532, A1=>nx17077, S0=>
      nx17569);
   ix7940 : mux21 port map ( Y=>nx7939, A0=>nx14535, A1=>nx17079, S0=>
      nx17575);
   ix9200 : mux21 port map ( Y=>nx9199, A0=>nx14545, A1=>nx17081, S0=>
      nx17297);
   ix9190 : mux21 port map ( Y=>nx9189, A0=>nx17081, A1=>nx14550, S0=>
      nx17291);
   ix9170 : mux21 port map ( Y=>nx9169, A0=>nx17081, A1=>nx14554, S0=>
      nx17279);
   ix9180 : mux21 port map ( Y=>nx9179, A0=>nx17081, A1=>nx14557, S0=>
      nx17285);
   ix9150 : mux21 port map ( Y=>nx9149, A0=>nx14563, A1=>nx17081, S0=>
      nx17307);
   ix9160 : mux21 port map ( Y=>nx9159, A0=>nx14566, A1=>nx17081, S0=>
      nx17313);
   ix9140 : mux21 port map ( Y=>nx9139, A0=>nx14570, A1=>nx17081, S0=>
      nx17319);
   ix9130 : mux21 port map ( Y=>nx9129, A0=>nx14573, A1=>nx17083, S0=>
      nx17325);
   ix9120 : mux21 port map ( Y=>nx9119, A0=>nx17083, A1=>nx14579, S0=>
      nx17273);
   ix9110 : mux21 port map ( Y=>nx9109, A0=>nx14583, A1=>nx17083, S0=>
      nx17331);
   ix9090 : mux21 port map ( Y=>nx9089, A0=>nx14587, A1=>nx17083, S0=>
      nx17337);
   ix9100 : mux21 port map ( Y=>nx9099, A0=>nx14590, A1=>nx17083, S0=>
      nx17343);
   ix9080 : mux21 port map ( Y=>nx9079, A0=>nx14596, A1=>nx17083, S0=>
      nx17349);
   ix9070 : mux21 port map ( Y=>nx9069, A0=>nx17083, A1=>nx14600, S0=>
      nx17267);
   ix9050 : mux21 port map ( Y=>nx9049, A0=>nx14604, A1=>nx17085, S0=>
      nx17355);
   ix9060 : mux21 port map ( Y=>nx9059, A0=>nx14607, A1=>nx17085, S0=>
      nx17361);
   ix9040 : mux21 port map ( Y=>nx9039, A0=>nx17085, A1=>nx14614, S0=>
      nx17261);
   ix9030 : mux21 port map ( Y=>nx9029, A0=>nx14618, A1=>nx17085, S0=>
      nx17367);
   ix9010 : mux21 port map ( Y=>nx9009, A0=>nx17085, A1=>nx14622, S0=>
      nx17255);
   ix9020 : mux21 port map ( Y=>nx9019, A0=>nx14625, A1=>nx17085, S0=>
      nx17373);
   ix9000 : mux21 port map ( Y=>nx8999, A0=>nx14631, A1=>nx17085, S0=>
      nx17379);
   ix8990 : mux21 port map ( Y=>nx8989, A0=>nx14635, A1=>nx17087, S0=>
      nx17385);
   ix8970 : mux21 port map ( Y=>nx8969, A0=>nx17087, A1=>nx14639, S0=>
      nx17249);
   ix8980 : mux21 port map ( Y=>nx8979, A0=>nx14642, A1=>nx17087, S0=>
      nx17391);
   ix8960 : mux21 port map ( Y=>nx8959, A0=>nx14648, A1=>nx17087, S0=>
      nx17397);
   ix8950 : mux21 port map ( Y=>nx8949, A0=>nx14652, A1=>nx17087, S0=>
      nx17403);
   ix8930 : mux21 port map ( Y=>nx8929, A0=>nx17087, A1=>nx14656, S0=>
      nx17243);
   ix8940 : mux21 port map ( Y=>nx8939, A0=>nx14659, A1=>nx17087, S0=>
      nx17409);
   ix8920 : mux21 port map ( Y=>nx8919, A0=>nx14665, A1=>nx17089, S0=>
      nx17415);
   ix8910 : mux21 port map ( Y=>nx8909, A0=>nx14669, A1=>nx17089, S0=>
      nx17421);
   ix8890 : mux21 port map ( Y=>nx8889, A0=>nx17089, A1=>nx14673, S0=>
      nx17237);
   ix8900 : mux21 port map ( Y=>nx8899, A0=>nx14676, A1=>nx17089, S0=>
      nx17427);
   ix8870 : mux21 port map ( Y=>nx8869, A0=>nx14686, A1=>nx17089, S0=>
      nx17433);
   ix8880 : mux21 port map ( Y=>nx8879, A0=>nx17089, A1=>nx14689, S0=>
      nx17231);
   ix8860 : mux21 port map ( Y=>nx8859, A0=>nx17089, A1=>nx14693, S0=>
      nx17225);
   ix8850 : mux21 port map ( Y=>nx8849, A0=>nx14696, A1=>nx17091, S0=>
      nx17439);
   ix8840 : mux21 port map ( Y=>nx8839, A0=>nx14703, A1=>nx17091, S0=>
      nx17445);
   ix8830 : mux21 port map ( Y=>nx8829, A0=>nx17091, A1=>nx14707, S0=>
      nx17219);
   ix8820 : mux21 port map ( Y=>nx8819, A0=>nx14714, A1=>nx17091, S0=>
      nx17453);
   ix8810 : mux21 port map ( Y=>nx8809, A0=>nx17091, A1=>nx14720, S0=>
      nx17213);
   ix8800 : mux21 port map ( Y=>nx8799, A0=>nx14725, A1=>nx17091, S0=>
      nx17465);
   ix8790 : mux21 port map ( Y=>nx8789, A0=>nx14729, A1=>nx17091, S0=>
      nx17471);
   ix8780 : mux21 port map ( Y=>nx8779, A0=>nx14733, A1=>nx17093, S0=>
      nx17477);
   ix8770 : mux21 port map ( Y=>nx8769, A0=>nx14736, A1=>nx17093, S0=>
      nx17485);
   ix8760 : mux21 port map ( Y=>nx8759, A0=>nx17093, A1=>nx14742, S0=>
      nx17207);
   ix8750 : mux21 port map ( Y=>nx8749, A0=>nx14746, A1=>nx17093, S0=>
      nx17491);
   ix8740 : mux21 port map ( Y=>nx8739, A0=>nx14750, A1=>nx17093, S0=>
      nx17497);
   ix8730 : mux21 port map ( Y=>nx8729, A0=>nx14753, A1=>nx17093, S0=>
      nx17503);
   ix8710 : mux21 port map ( Y=>nx8709, A0=>nx14760, A1=>nx17093, S0=>
      nx17509);
   ix8720 : mux21 port map ( Y=>nx8719, A0=>nx14763, A1=>nx17095, S0=>
      nx17515);
   ix8700 : mux21 port map ( Y=>nx8699, A0=>nx14767, A1=>nx17095, S0=>
      nx17521);
   ix8690 : mux21 port map ( Y=>nx8689, A0=>nx14770, A1=>nx17095, S0=>
      nx17527);
   ix8680 : mux21 port map ( Y=>nx8679, A0=>nx14776, A1=>nx17095, S0=>
      nx17533);
   ix8670 : mux21 port map ( Y=>nx8669, A0=>nx17095, A1=>nx14780, S0=>
      nx17201);
   ix8660 : mux21 port map ( Y=>nx8659, A0=>nx14784, A1=>nx17095, S0=>
      nx17539);
   ix8650 : mux21 port map ( Y=>nx8649, A0=>nx17095, A1=>nx14787, S0=>
      nx17195);
   ix8640 : mux21 port map ( Y=>nx8639, A0=>nx14793, A1=>nx17097, S0=>
      nx17545);
   ix8630 : mux21 port map ( Y=>nx8629, A0=>nx17097, A1=>nx14797, S0=>
      nx17189);
   ix8620 : mux21 port map ( Y=>nx8619, A0=>nx17097, A1=>nx14801, S0=>
      nx17183);
   ix8610 : mux21 port map ( Y=>nx8609, A0=>nx14804, A1=>nx17097, S0=>
      nx17551);
   ix8600 : mux21 port map ( Y=>nx8599, A0=>nx14810, A1=>nx17097, S0=>
      nx17557);
   ix8590 : mux21 port map ( Y=>nx8589, A0=>nx14814, A1=>nx17097, S0=>
      nx17563);
   ix8570 : mux21 port map ( Y=>nx8569, A0=>nx14818, A1=>nx17097, S0=>
      nx17569);
   ix8580 : mux21 port map ( Y=>nx8579, A0=>nx14821, A1=>nx17099, S0=>
      nx17575);
   ix9840 : mux21 port map ( Y=>nx9839, A0=>nx14831, A1=>nx17101, S0=>
      nx17299);
   ix9830 : mux21 port map ( Y=>nx9829, A0=>nx17101, A1=>nx14836, S0=>
      nx17293);
   ix9810 : mux21 port map ( Y=>nx9809, A0=>nx17101, A1=>nx14840, S0=>
      nx17281);
   ix9820 : mux21 port map ( Y=>nx9819, A0=>nx17101, A1=>nx14843, S0=>
      nx17287);
   ix9790 : mux21 port map ( Y=>nx9789, A0=>nx14849, A1=>nx17101, S0=>
      nx17309);
   ix9800 : mux21 port map ( Y=>nx9799, A0=>nx14852, A1=>nx17101, S0=>
      nx17315);
   ix9780 : mux21 port map ( Y=>nx9779, A0=>nx14856, A1=>nx17101, S0=>
      nx17321);
   ix9770 : mux21 port map ( Y=>nx9769, A0=>nx14859, A1=>nx17103, S0=>
      nx17327);
   ix9760 : mux21 port map ( Y=>nx9759, A0=>nx17103, A1=>nx14865, S0=>
      nx17275);
   ix9750 : mux21 port map ( Y=>nx9749, A0=>nx14869, A1=>nx17103, S0=>
      nx17333);
   ix9730 : mux21 port map ( Y=>nx9729, A0=>nx14873, A1=>nx17103, S0=>
      nx17339);
   ix9740 : mux21 port map ( Y=>nx9739, A0=>nx14876, A1=>nx17103, S0=>
      nx17345);
   ix9720 : mux21 port map ( Y=>nx9719, A0=>nx14882, A1=>nx17103, S0=>
      nx17351);
   ix9710 : mux21 port map ( Y=>nx9709, A0=>nx17103, A1=>nx14886, S0=>
      nx17269);
   ix9690 : mux21 port map ( Y=>nx9689, A0=>nx14890, A1=>nx17105, S0=>
      nx17357);
   ix9700 : mux21 port map ( Y=>nx9699, A0=>nx14893, A1=>nx17105, S0=>
      nx17363);
   ix9680 : mux21 port map ( Y=>nx9679, A0=>nx17105, A1=>nx14900, S0=>
      nx17263);
   ix9670 : mux21 port map ( Y=>nx9669, A0=>nx14904, A1=>nx17105, S0=>
      nx17369);
   ix9650 : mux21 port map ( Y=>nx9649, A0=>nx17105, A1=>nx14908, S0=>
      nx17257);
   ix9660 : mux21 port map ( Y=>nx9659, A0=>nx14911, A1=>nx17105, S0=>
      nx17375);
   ix9640 : mux21 port map ( Y=>nx9639, A0=>nx14917, A1=>nx17105, S0=>
      nx17381);
   ix9630 : mux21 port map ( Y=>nx9629, A0=>nx14921, A1=>nx17107, S0=>
      nx17387);
   ix9610 : mux21 port map ( Y=>nx9609, A0=>nx17107, A1=>nx14925, S0=>
      nx17251);
   ix9620 : mux21 port map ( Y=>nx9619, A0=>nx14928, A1=>nx17107, S0=>
      nx17393);
   ix9600 : mux21 port map ( Y=>nx9599, A0=>nx14934, A1=>nx17107, S0=>
      nx17399);
   ix9590 : mux21 port map ( Y=>nx9589, A0=>nx14938, A1=>nx17107, S0=>
      nx17405);
   ix9570 : mux21 port map ( Y=>nx9569, A0=>nx17107, A1=>nx14942, S0=>
      nx17245);
   ix9580 : mux21 port map ( Y=>nx9579, A0=>nx14945, A1=>nx17107, S0=>
      nx17411);
   ix9560 : mux21 port map ( Y=>nx9559, A0=>nx14951, A1=>nx17109, S0=>
      nx17417);
   ix9550 : mux21 port map ( Y=>nx9549, A0=>nx14955, A1=>nx17109, S0=>
      nx17423);
   ix9530 : mux21 port map ( Y=>nx9529, A0=>nx17109, A1=>nx14959, S0=>
      nx17239);
   ix9540 : mux21 port map ( Y=>nx9539, A0=>nx14962, A1=>nx17109, S0=>
      nx17429);
   ix9510 : mux21 port map ( Y=>nx9509, A0=>nx14972, A1=>nx17109, S0=>
      nx17435);
   ix9520 : mux21 port map ( Y=>nx9519, A0=>nx17109, A1=>nx14975, S0=>
      nx17233);
   ix9500 : mux21 port map ( Y=>nx9499, A0=>nx17109, A1=>nx14979, S0=>
      nx17227);
   ix9490 : mux21 port map ( Y=>nx9489, A0=>nx14982, A1=>nx17111, S0=>
      nx17441);
   ix9480 : mux21 port map ( Y=>nx9479, A0=>nx14989, A1=>nx17111, S0=>
      nx17447);
   ix9470 : mux21 port map ( Y=>nx9469, A0=>nx17111, A1=>nx14993, S0=>
      nx17221);
   ix9460 : mux21 port map ( Y=>nx9459, A0=>nx15000, A1=>nx17111, S0=>
      nx17455);
   ix9450 : mux21 port map ( Y=>nx9449, A0=>nx17111, A1=>nx15006, S0=>
      nx17215);
   ix9440 : mux21 port map ( Y=>nx9439, A0=>nx15011, A1=>nx17111, S0=>
      nx17467);
   ix9430 : mux21 port map ( Y=>nx9429, A0=>nx15015, A1=>nx17111, S0=>
      nx17473);
   ix9420 : mux21 port map ( Y=>nx9419, A0=>nx15019, A1=>nx17113, S0=>
      nx17479);
   ix9410 : mux21 port map ( Y=>nx9409, A0=>nx15022, A1=>nx17113, S0=>
      nx17487);
   ix9400 : mux21 port map ( Y=>nx9399, A0=>nx17113, A1=>nx15028, S0=>
      nx17209);
   ix9390 : mux21 port map ( Y=>nx9389, A0=>nx15032, A1=>nx17113, S0=>
      nx17493);
   ix9380 : mux21 port map ( Y=>nx9379, A0=>nx15036, A1=>nx17113, S0=>
      nx17499);
   ix9370 : mux21 port map ( Y=>nx9369, A0=>nx15039, A1=>nx17113, S0=>
      nx17505);
   ix9350 : mux21 port map ( Y=>nx9349, A0=>nx15046, A1=>nx17113, S0=>
      nx17511);
   ix9360 : mux21 port map ( Y=>nx9359, A0=>nx15049, A1=>nx17115, S0=>
      nx17517);
   ix9340 : mux21 port map ( Y=>nx9339, A0=>nx15053, A1=>nx17115, S0=>
      nx17523);
   ix9330 : mux21 port map ( Y=>nx9329, A0=>nx15056, A1=>nx17115, S0=>
      nx17529);
   ix9320 : mux21 port map ( Y=>nx9319, A0=>nx15062, A1=>nx17115, S0=>
      nx17535);
   ix9310 : mux21 port map ( Y=>nx9309, A0=>nx17115, A1=>nx15066, S0=>
      nx17203);
   ix9300 : mux21 port map ( Y=>nx9299, A0=>nx15070, A1=>nx17115, S0=>
      nx17541);
   ix9290 : mux21 port map ( Y=>nx9289, A0=>nx17115, A1=>nx15073, S0=>
      nx17197);
   ix9280 : mux21 port map ( Y=>nx9279, A0=>nx15079, A1=>nx17117, S0=>
      nx17547);
   ix9270 : mux21 port map ( Y=>nx9269, A0=>nx17117, A1=>nx15083, S0=>
      nx17191);
   ix9260 : mux21 port map ( Y=>nx9259, A0=>nx17117, A1=>nx15087, S0=>
      nx17185);
   ix9250 : mux21 port map ( Y=>nx9249, A0=>nx15090, A1=>nx17117, S0=>
      nx17553);
   ix9240 : mux21 port map ( Y=>nx9239, A0=>nx15096, A1=>nx17117, S0=>
      nx17559);
   ix9230 : mux21 port map ( Y=>nx9229, A0=>nx15100, A1=>nx17117, S0=>
      nx17565);
   ix9210 : mux21 port map ( Y=>nx9209, A0=>nx15104, A1=>nx17117, S0=>
      nx17571);
   ix9220 : mux21 port map ( Y=>nx9219, A0=>nx15107, A1=>nx17119, S0=>
      nx17577);
   ix10480 : mux21 port map ( Y=>nx10479, A0=>nx15117, A1=>nx17121, S0=>
      nx17299);
   ix10470 : mux21 port map ( Y=>nx10469, A0=>nx17121, A1=>nx15122, S0=>
      nx17293);
   ix10450 : mux21 port map ( Y=>nx10449, A0=>nx17121, A1=>nx15126, S0=>
      nx17281);
   ix10460 : mux21 port map ( Y=>nx10459, A0=>nx17121, A1=>nx15129, S0=>
      nx17287);
   ix10430 : mux21 port map ( Y=>nx10429, A0=>nx15135, A1=>nx17121, S0=>
      nx17309);
   ix10440 : mux21 port map ( Y=>nx10439, A0=>nx15138, A1=>nx17121, S0=>
      nx17315);
   ix10420 : mux21 port map ( Y=>nx10419, A0=>nx15142, A1=>nx17121, S0=>
      nx17321);
   ix10410 : mux21 port map ( Y=>nx10409, A0=>nx15145, A1=>nx17123, S0=>
      nx17327);
   ix10400 : mux21 port map ( Y=>nx10399, A0=>nx17123, A1=>nx15151, S0=>
      nx17275);
   ix10390 : mux21 port map ( Y=>nx10389, A0=>nx15155, A1=>nx17123, S0=>
      nx17333);
   ix10370 : mux21 port map ( Y=>nx10369, A0=>nx15159, A1=>nx17123, S0=>
      nx17339);
   ix10380 : mux21 port map ( Y=>nx10379, A0=>nx15162, A1=>nx17123, S0=>
      nx17345);
   ix10360 : mux21 port map ( Y=>nx10359, A0=>nx15168, A1=>nx17123, S0=>
      nx17351);
   ix10350 : mux21 port map ( Y=>nx10349, A0=>nx17123, A1=>nx15172, S0=>
      nx17269);
   ix10330 : mux21 port map ( Y=>nx10329, A0=>nx15176, A1=>nx17125, S0=>
      nx17357);
   ix10340 : mux21 port map ( Y=>nx10339, A0=>nx15179, A1=>nx17125, S0=>
      nx17363);
   ix10320 : mux21 port map ( Y=>nx10319, A0=>nx17125, A1=>nx15186, S0=>
      nx17263);
   ix10310 : mux21 port map ( Y=>nx10309, A0=>nx15190, A1=>nx17125, S0=>
      nx17369);
   ix10290 : mux21 port map ( Y=>nx10289, A0=>nx17125, A1=>nx15194, S0=>
      nx17257);
   ix10300 : mux21 port map ( Y=>nx10299, A0=>nx15197, A1=>nx17125, S0=>
      nx17375);
   ix10280 : mux21 port map ( Y=>nx10279, A0=>nx15203, A1=>nx17125, S0=>
      nx17381);
   ix10270 : mux21 port map ( Y=>nx10269, A0=>nx15207, A1=>nx17127, S0=>
      nx17387);
   ix10250 : mux21 port map ( Y=>nx10249, A0=>nx17127, A1=>nx15211, S0=>
      nx17251);
   ix10260 : mux21 port map ( Y=>nx10259, A0=>nx15214, A1=>nx17127, S0=>
      nx17393);
   ix10240 : mux21 port map ( Y=>nx10239, A0=>nx15220, A1=>nx17127, S0=>
      nx17399);
   ix10230 : mux21 port map ( Y=>nx10229, A0=>nx15224, A1=>nx17127, S0=>
      nx17405);
   ix10210 : mux21 port map ( Y=>nx10209, A0=>nx17127, A1=>nx15228, S0=>
      nx17245);
   ix10220 : mux21 port map ( Y=>nx10219, A0=>nx15231, A1=>nx17127, S0=>
      nx17411);
   ix10200 : mux21 port map ( Y=>nx10199, A0=>nx15237, A1=>nx17129, S0=>
      nx17417);
   ix10190 : mux21 port map ( Y=>nx10189, A0=>nx15241, A1=>nx17129, S0=>
      nx17423);
   ix10170 : mux21 port map ( Y=>nx10169, A0=>nx17129, A1=>nx15245, S0=>
      nx17239);
   ix10180 : mux21 port map ( Y=>nx10179, A0=>nx15248, A1=>nx17129, S0=>
      nx17429);
   ix10150 : mux21 port map ( Y=>nx10149, A0=>nx15258, A1=>nx17129, S0=>
      nx17435);
   ix10160 : mux21 port map ( Y=>nx10159, A0=>nx17129, A1=>nx15261, S0=>
      nx17233);
   ix10140 : mux21 port map ( Y=>nx10139, A0=>nx17129, A1=>nx15265, S0=>
      nx17227);
   ix10130 : mux21 port map ( Y=>nx10129, A0=>nx15268, A1=>nx17131, S0=>
      nx17441);
   ix10120 : mux21 port map ( Y=>nx10119, A0=>nx15275, A1=>nx17131, S0=>
      nx17447);
   ix10110 : mux21 port map ( Y=>nx10109, A0=>nx17131, A1=>nx15279, S0=>
      nx17221);
   ix10100 : mux21 port map ( Y=>nx10099, A0=>nx15286, A1=>nx17131, S0=>
      nx17455);
   ix10090 : mux21 port map ( Y=>nx10089, A0=>nx17131, A1=>nx15292, S0=>
      nx17215);
   ix10080 : mux21 port map ( Y=>nx10079, A0=>nx15297, A1=>nx17131, S0=>
      nx17467);
   ix10070 : mux21 port map ( Y=>nx10069, A0=>nx15301, A1=>nx17131, S0=>
      nx17473);
   ix10060 : mux21 port map ( Y=>nx10059, A0=>nx15305, A1=>nx17133, S0=>
      nx17479);
   ix10050 : mux21 port map ( Y=>nx10049, A0=>nx15308, A1=>nx17133, S0=>
      nx17487);
   ix10040 : mux21 port map ( Y=>nx10039, A0=>nx17133, A1=>nx15314, S0=>
      nx17209);
   ix10030 : mux21 port map ( Y=>nx10029, A0=>nx15318, A1=>nx17133, S0=>
      nx17493);
   ix10020 : mux21 port map ( Y=>nx10019, A0=>nx15322, A1=>nx17133, S0=>
      nx17499);
   ix10010 : mux21 port map ( Y=>nx10009, A0=>nx15325, A1=>nx17133, S0=>
      nx17505);
   ix9990 : mux21 port map ( Y=>nx9989, A0=>nx15332, A1=>nx17133, S0=>
      nx17511);
   ix10000 : mux21 port map ( Y=>nx9999, A0=>nx15335, A1=>nx17135, S0=>
      nx17517);
   ix9980 : mux21 port map ( Y=>nx9979, A0=>nx15339, A1=>nx17135, S0=>
      nx17523);
   ix9970 : mux21 port map ( Y=>nx9969, A0=>nx15342, A1=>nx17135, S0=>
      nx17529);
   ix9960 : mux21 port map ( Y=>nx9959, A0=>nx15348, A1=>nx17135, S0=>
      nx17535);
   ix9950 : mux21 port map ( Y=>nx9949, A0=>nx17135, A1=>nx15352, S0=>
      nx17203);
   ix9940 : mux21 port map ( Y=>nx9939, A0=>nx15356, A1=>nx17135, S0=>
      nx17541);
   ix9930 : mux21 port map ( Y=>nx9929, A0=>nx17135, A1=>nx15359, S0=>
      nx17197);
   ix9920 : mux21 port map ( Y=>nx9919, A0=>nx15365, A1=>nx17137, S0=>
      nx17547);
   ix9910 : mux21 port map ( Y=>nx9909, A0=>nx17137, A1=>nx15369, S0=>
      nx17191);
   ix9900 : mux21 port map ( Y=>nx9899, A0=>nx17137, A1=>nx15373, S0=>
      nx17185);
   ix9890 : mux21 port map ( Y=>nx9889, A0=>nx15376, A1=>nx17137, S0=>
      nx17553);
   ix9880 : mux21 port map ( Y=>nx9879, A0=>nx15382, A1=>nx17137, S0=>
      nx17559);
   ix9870 : mux21 port map ( Y=>nx9869, A0=>nx15386, A1=>nx17137, S0=>
      nx17565);
   ix9850 : mux21 port map ( Y=>nx9849, A0=>nx15390, A1=>nx17137, S0=>
      nx17571);
   ix9860 : mux21 port map ( Y=>nx9859, A0=>nx15393, A1=>nx17139, S0=>
      nx17577);
   ix17178 : inv04 port map ( Y=>nx17179, A=>nx10579);
   ix17180 : inv02 port map ( Y=>nx17181, A=>nx158);
   ix17182 : inv02 port map ( Y=>nx17183, A=>nx158);
   ix17184 : inv02 port map ( Y=>nx17185, A=>nx158);
   ix17186 : inv02 port map ( Y=>nx17187, A=>nx178);
   ix17188 : inv02 port map ( Y=>nx17189, A=>nx178);
   ix17190 : inv02 port map ( Y=>nx17191, A=>nx178);
   ix17192 : inv02 port map ( Y=>nx17193, A=>nx226);
   ix17194 : inv02 port map ( Y=>nx17195, A=>nx226);
   ix17196 : inv02 port map ( Y=>nx17197, A=>nx226);
   ix17198 : inv02 port map ( Y=>nx17199, A=>nx264);
   ix17200 : inv02 port map ( Y=>nx17201, A=>nx264);
   ix17202 : inv02 port map ( Y=>nx17203, A=>nx264);
   ix17204 : inv02 port map ( Y=>nx17205, A=>nx456);
   ix17206 : inv02 port map ( Y=>nx17207, A=>nx456);
   ix17208 : inv02 port map ( Y=>nx17209, A=>nx456);
   ix17210 : inv02 port map ( Y=>nx17211, A=>nx560);
   ix17212 : inv02 port map ( Y=>nx17213, A=>nx560);
   ix17214 : inv02 port map ( Y=>nx17215, A=>nx560);
   ix17216 : inv02 port map ( Y=>nx17217, A=>nx598);
   ix17218 : inv02 port map ( Y=>nx17219, A=>nx598);
   ix17220 : inv02 port map ( Y=>nx17221, A=>nx598);
   ix17222 : inv02 port map ( Y=>nx17223, A=>nx656);
   ix17224 : inv02 port map ( Y=>nx17225, A=>nx656);
   ix17226 : inv02 port map ( Y=>nx17227, A=>nx656);
   ix17228 : inv02 port map ( Y=>nx17229, A=>nx698);
   ix17230 : inv02 port map ( Y=>nx17231, A=>nx698);
   ix17232 : inv02 port map ( Y=>nx17233, A=>nx698);
   ix17234 : inv02 port map ( Y=>nx17235, A=>nx726);
   ix17236 : inv02 port map ( Y=>nx17237, A=>nx726);
   ix17238 : inv02 port map ( Y=>nx17239, A=>nx726);
   ix17240 : inv02 port map ( Y=>nx17241, A=>nx806);
   ix17242 : inv02 port map ( Y=>nx17243, A=>nx806);
   ix17244 : inv02 port map ( Y=>nx17245, A=>nx806);
   ix17246 : inv02 port map ( Y=>nx17247, A=>nx888);
   ix17248 : inv02 port map ( Y=>nx17249, A=>nx888);
   ix17250 : inv02 port map ( Y=>nx17251, A=>nx888);
   ix17252 : inv02 port map ( Y=>nx17253, A=>nx968);
   ix17254 : inv02 port map ( Y=>nx17255, A=>nx968);
   ix17256 : inv02 port map ( Y=>nx17257, A=>nx968);
   ix17258 : inv02 port map ( Y=>nx17259, A=>nx1026);
   ix17260 : inv02 port map ( Y=>nx17261, A=>nx1026);
   ix17262 : inv02 port map ( Y=>nx17263, A=>nx1026);
   ix17264 : inv02 port map ( Y=>nx17265, A=>nx1092);
   ix17266 : inv02 port map ( Y=>nx17267, A=>nx1092);
   ix17268 : inv02 port map ( Y=>nx17269, A=>nx1092);
   ix17270 : inv02 port map ( Y=>nx17271, A=>nx1188);
   ix17272 : inv02 port map ( Y=>nx17273, A=>nx1188);
   ix17274 : inv02 port map ( Y=>nx17275, A=>nx1188);
   ix17276 : inv02 port map ( Y=>nx17277, A=>nx1292);
   ix17278 : inv02 port map ( Y=>nx17279, A=>nx1292);
   ix17280 : inv02 port map ( Y=>nx17281, A=>nx1292);
   ix17282 : inv02 port map ( Y=>nx17283, A=>nx1310);
   ix17284 : inv02 port map ( Y=>nx17285, A=>nx1310);
   ix17286 : inv02 port map ( Y=>nx17287, A=>nx1310);
   ix17288 : inv02 port map ( Y=>nx17289, A=>nx1330);
   ix17290 : inv02 port map ( Y=>nx17291, A=>nx1330);
   ix17292 : inv02 port map ( Y=>nx17293, A=>nx1330);
   ix17294 : inv02 port map ( Y=>nx17295, A=>nx10503);
   ix17296 : inv02 port map ( Y=>nx17297, A=>nx10503);
   ix17298 : inv02 port map ( Y=>nx17299, A=>nx10503);
   ix17302 : inv02 port map ( Y=>nx17303, A=>nx10545);
   ix17304 : inv02 port map ( Y=>nx17305, A=>nx10577);
   ix17306 : inv02 port map ( Y=>nx17307, A=>nx10577);
   ix17308 : inv02 port map ( Y=>nx17309, A=>nx10577);
   ix17310 : inv02 port map ( Y=>nx17311, A=>nx10587);
   ix17312 : inv02 port map ( Y=>nx17313, A=>nx10587);
   ix17314 : inv02 port map ( Y=>nx17315, A=>nx10587);
   ix17316 : inv02 port map ( Y=>nx17317, A=>nx10599);
   ix17318 : inv02 port map ( Y=>nx17319, A=>nx10599);
   ix17320 : inv02 port map ( Y=>nx17321, A=>nx10599);
   ix17322 : inv02 port map ( Y=>nx17323, A=>nx10607);
   ix17324 : inv02 port map ( Y=>nx17325, A=>nx10607);
   ix17326 : inv02 port map ( Y=>nx17327, A=>nx10607);
   ix17328 : inv02 port map ( Y=>nx17329, A=>nx10633);
   ix17330 : inv02 port map ( Y=>nx17331, A=>nx10633);
   ix17332 : inv02 port map ( Y=>nx17333, A=>nx10633);
   ix17334 : inv02 port map ( Y=>nx17335, A=>nx10641);
   ix17336 : inv02 port map ( Y=>nx17337, A=>nx10641);
   ix17338 : inv02 port map ( Y=>nx17339, A=>nx10641);
   ix17340 : inv02 port map ( Y=>nx17341, A=>nx10648);
   ix17342 : inv02 port map ( Y=>nx17343, A=>nx10648);
   ix17344 : inv02 port map ( Y=>nx17345, A=>nx10648);
   ix17346 : inv02 port map ( Y=>nx17347, A=>nx10657);
   ix17348 : inv02 port map ( Y=>nx17349, A=>nx10657);
   ix17350 : inv02 port map ( Y=>nx17351, A=>nx10657);
   ix17352 : inv02 port map ( Y=>nx17353, A=>nx10677);
   ix17354 : inv02 port map ( Y=>nx17355, A=>nx10677);
   ix17356 : inv02 port map ( Y=>nx17357, A=>nx10677);
   ix17358 : inv02 port map ( Y=>nx17359, A=>nx10684);
   ix17360 : inv02 port map ( Y=>nx17361, A=>nx10684);
   ix17362 : inv02 port map ( Y=>nx17363, A=>nx10684);
   ix17364 : inv02 port map ( Y=>nx17365, A=>nx10703);
   ix17366 : inv02 port map ( Y=>nx17367, A=>nx10703);
   ix17368 : inv02 port map ( Y=>nx17369, A=>nx10703);
   ix17370 : inv02 port map ( Y=>nx17371, A=>nx10716);
   ix17372 : inv02 port map ( Y=>nx17373, A=>nx10716);
   ix17374 : inv02 port map ( Y=>nx17375, A=>nx10716);
   ix17376 : inv02 port map ( Y=>nx17377, A=>nx10727);
   ix17378 : inv02 port map ( Y=>nx17379, A=>nx10727);
   ix17380 : inv02 port map ( Y=>nx17381, A=>nx10727);
   ix17382 : inv02 port map ( Y=>nx17383, A=>nx10734);
   ix17384 : inv02 port map ( Y=>nx17385, A=>nx10734);
   ix17386 : inv02 port map ( Y=>nx17387, A=>nx10734);
   ix17388 : inv02 port map ( Y=>nx17389, A=>nx10754);
   ix17390 : inv02 port map ( Y=>nx17391, A=>nx10754);
   ix17392 : inv02 port map ( Y=>nx17393, A=>nx10754);
   ix17394 : inv02 port map ( Y=>nx17395, A=>nx10765);
   ix17396 : inv02 port map ( Y=>nx17397, A=>nx10765);
   ix17398 : inv02 port map ( Y=>nx17399, A=>nx10765);
   ix17400 : inv02 port map ( Y=>nx17401, A=>nx10772);
   ix17402 : inv02 port map ( Y=>nx17403, A=>nx10772);
   ix17404 : inv02 port map ( Y=>nx17405, A=>nx10772);
   ix17406 : inv02 port map ( Y=>nx17407, A=>nx10793);
   ix17408 : inv02 port map ( Y=>nx17409, A=>nx10793);
   ix17410 : inv02 port map ( Y=>nx17411, A=>nx10793);
   ix17412 : inv02 port map ( Y=>nx17413, A=>nx10804);
   ix17414 : inv02 port map ( Y=>nx17415, A=>nx10804);
   ix17416 : inv02 port map ( Y=>nx17417, A=>nx10804);
   ix17418 : inv02 port map ( Y=>nx17419, A=>nx10811);
   ix17420 : inv02 port map ( Y=>nx17421, A=>nx10811);
   ix17422 : inv02 port map ( Y=>nx17423, A=>nx10811);
   ix17424 : inv02 port map ( Y=>nx17425, A=>nx10829);
   ix17426 : inv02 port map ( Y=>nx17427, A=>nx10829);
   ix17428 : inv02 port map ( Y=>nx17429, A=>nx10829);
   ix17430 : inv02 port map ( Y=>nx17431, A=>nx10844);
   ix17432 : inv02 port map ( Y=>nx17433, A=>nx10844);
   ix17434 : inv02 port map ( Y=>nx17435, A=>nx10844);
   ix17436 : inv02 port map ( Y=>nx17437, A=>nx10872);
   ix17438 : inv02 port map ( Y=>nx17439, A=>nx10872);
   ix17440 : inv02 port map ( Y=>nx17441, A=>nx10872);
   ix17442 : inv02 port map ( Y=>nx17443, A=>nx10887);
   ix17444 : inv02 port map ( Y=>nx17445, A=>nx10887);
   ix17446 : inv02 port map ( Y=>nx17447, A=>nx10887);
   ix17448 : inv01 port map ( Y=>nx17449, A=>nx16557);
   ix17450 : inv02 port map ( Y=>nx17451, A=>nx17449);
   ix17452 : inv02 port map ( Y=>nx17453, A=>nx17449);
   ix17454 : inv02 port map ( Y=>nx17455, A=>nx17449);
   ix17456 : inv02 port map ( Y=>nx17457, A=>nx10907);
   ix17458 : inv02 port map ( Y=>nx17459, A=>nx10907);
   ix17460 : inv01 port map ( Y=>nx17461, A=>nx16577);
   ix17462 : inv02 port map ( Y=>nx17463, A=>nx17461);
   ix17464 : inv02 port map ( Y=>nx17465, A=>nx17461);
   ix17466 : inv02 port map ( Y=>nx17467, A=>nx17461);
   ix17468 : inv02 port map ( Y=>nx17469, A=>nx10931);
   ix17470 : inv02 port map ( Y=>nx17471, A=>nx10931);
   ix17472 : inv02 port map ( Y=>nx17473, A=>nx10931);
   ix17474 : inv02 port map ( Y=>nx17475, A=>nx10939);
   ix17476 : inv02 port map ( Y=>nx17477, A=>nx10939);
   ix17478 : inv02 port map ( Y=>nx17479, A=>nx10939);
   ix17480 : inv01 port map ( Y=>nx17481, A=>nx16609);
   ix17482 : inv02 port map ( Y=>nx17483, A=>nx17481);
   ix17484 : inv02 port map ( Y=>nx17485, A=>nx17481);
   ix17486 : inv02 port map ( Y=>nx17487, A=>nx17481);
   ix17488 : inv02 port map ( Y=>nx17489, A=>nx10962);
   ix17490 : inv02 port map ( Y=>nx17491, A=>nx10962);
   ix17492 : inv02 port map ( Y=>nx17493, A=>nx10962);
   ix17494 : inv02 port map ( Y=>nx17495, A=>nx10968);
   ix17496 : inv02 port map ( Y=>nx17497, A=>nx10968);
   ix17498 : inv02 port map ( Y=>nx17499, A=>nx10968);
   ix17500 : inv02 port map ( Y=>nx17501, A=>nx10975);
   ix17502 : inv02 port map ( Y=>nx17503, A=>nx10975);
   ix17504 : inv02 port map ( Y=>nx17505, A=>nx10975);
   ix17506 : inv02 port map ( Y=>nx17507, A=>nx10986);
   ix17508 : inv02 port map ( Y=>nx17509, A=>nx10986);
   ix17510 : inv02 port map ( Y=>nx17511, A=>nx10986);
   ix17512 : inv02 port map ( Y=>nx17513, A=>nx10995);
   ix17514 : inv02 port map ( Y=>nx17515, A=>nx10995);
   ix17516 : inv02 port map ( Y=>nx17517, A=>nx10995);
   ix17518 : inv02 port map ( Y=>nx17519, A=>nx11003);
   ix17520 : inv02 port map ( Y=>nx17521, A=>nx11003);
   ix17522 : inv02 port map ( Y=>nx17523, A=>nx11003);
   ix17524 : inv02 port map ( Y=>nx17525, A=>nx11010);
   ix17526 : inv02 port map ( Y=>nx17527, A=>nx11010);
   ix17528 : inv02 port map ( Y=>nx17529, A=>nx11010);
   ix17530 : inv02 port map ( Y=>nx17531, A=>nx11022);
   ix17532 : inv02 port map ( Y=>nx17533, A=>nx11022);
   ix17534 : inv02 port map ( Y=>nx17535, A=>nx11022);
   ix17536 : inv02 port map ( Y=>nx17537, A=>nx11035);
   ix17538 : inv02 port map ( Y=>nx17539, A=>nx11035);
   ix17540 : inv02 port map ( Y=>nx17541, A=>nx11035);
   ix17542 : inv02 port map ( Y=>nx17543, A=>nx11054);
   ix17544 : inv02 port map ( Y=>nx17545, A=>nx11054);
   ix17546 : inv02 port map ( Y=>nx17547, A=>nx11054);
   ix17548 : inv02 port map ( Y=>nx17549, A=>nx11073);
   ix17550 : inv02 port map ( Y=>nx17551, A=>nx11073);
   ix17552 : inv02 port map ( Y=>nx17553, A=>nx11073);
   ix17554 : inv02 port map ( Y=>nx17555, A=>nx11083);
   ix17556 : inv02 port map ( Y=>nx17557, A=>nx11083);
   ix17558 : inv02 port map ( Y=>nx17559, A=>nx11083);
   ix17560 : inv02 port map ( Y=>nx17561, A=>nx11089);
   ix17562 : inv02 port map ( Y=>nx17563, A=>nx11089);
   ix17564 : inv02 port map ( Y=>nx17565, A=>nx11089);
   ix17566 : inv02 port map ( Y=>nx17567, A=>nx11095);
   ix17568 : inv02 port map ( Y=>nx17569, A=>nx11095);
   ix17570 : inv02 port map ( Y=>nx17571, A=>nx11095);
   ix17572 : inv02 port map ( Y=>nx17573, A=>nx11102);
   ix17574 : inv02 port map ( Y=>nx17575, A=>nx11102);
   ix17576 : inv02 port map ( Y=>nx17577, A=>nx11102);
   ix18959 : nor02ii port map ( Y=>nx18578, A0=>nx7268, A1=>nx13915);
   ix18960 : inv01 port map ( Y=>nx18579, A=>nx7250);
   reg_nx7274 : nand04_2x port map ( Y=>nx7274, A0=>nx18578, A1=>nx13949, A2
      =>nx13932, A3=>nx18579);
   ix18961 : inv02 port map ( Y=>nx18580, A=>address(4));
   ix18962 : inv02 port map ( Y=>nx18581, A=>address(5));
   ix18963 : inv01 port map ( Y=>nx18582, A=>nx16007);
   ix18964 : inv01 port map ( Y=>nx18583, A=>nx13790);
   ix18965 : inv01 port map ( Y=>nx18584, A=>nx15989);
   ix18966 : inv01 port map ( Y=>nx18585, A=>nx13794);
   ix18967 : inv01 port map ( Y=>nx18586, A=>nx15439);
   ix18968 : aoi43 port map ( Y=>nx18587, A0=>nx18580, A1=>nx18581, A2=>
      nx18582, A3=>nx18583, B0=>nx18584, B1=>nx18585, B2=>nx18586);
   reg_NOT_nx7538 : or03 port map ( Y=>NOT_nx7538, A0=>nx16007, A1=>nx13777, 
      A2=>nx15437);
   ix18969 : inv01 port map ( Y=>nx18588, A=>nx7744);
   ix18970 : nand04_2x port map ( Y=>nx18589, A0=>nx18587, A1=>NOT_nx7538, 
      A2=>nx13718, A3=>nx18588);
   ix18971 : oai43 port map ( Y=>nx18590, A0=>address(4), A1=>address(5), A2
      =>nx13773, A3=>nx16027, B0=>nx15989, B1=>nx13807, B2=>nx15863);
   ix18972 : inv01 port map ( Y=>nx18591, A=>nx18590);
   reg_NOT_nx7576 : or04 port map ( Y=>NOT_nx7576, A0=>address(4), A1=>
      address(5), A2=>nx16047, A3=>nx13760);
   ix18973 : nor02ii port map ( Y=>nx18592, A0=>nx7490, A1=>nx13864);
   ix18974 : nor02_2x port map ( Y=>nx18593, A0=>nx7726, A1=>nx7452);
   ix18975 : nand04_2x port map ( Y=>nx18594, A0=>nx18591, A1=>NOT_nx7576, 
      A2=>nx18592, A3=>nx18593);
   ix18976 : nor03_2x port map ( Y=>nx18595, A0=>nx7408, A1=>nx7426, A2=>
      nx7390);
   ix18977 : or03 port map ( Y=>nx18596, A0=>nx16047, A1=>nx13756, A2=>
      nx15827);
   ix18978 : inv01 port map ( Y=>nx18597, A=>nx7460);
   ix18979 : and03 port map ( Y=>nx18598, A0=>nx18596, A1=>nx13735, A2=>
      nx18597);
   ix18980 : nor02ii port map ( Y=>nx18599, A0=>nx7568, A1=>nx13881);
   ix18981 : nor02ii port map ( Y=>nx18600, A0=>nx7530, A1=>nx13702);
   ix18982 : nand04_2x port map ( Y=>nx18601, A0=>nx18595, A1=>nx18598, A2=>
      nx18599, A3=>nx18600);
   reg_nx13681 : nor04_2x port map ( Y=>nx13681, A0=>nx7274, A1=>nx18589, A2
      =>nx18594, A3=>nx18601);
   ix18983 : nor02ii port map ( Y=>nx18602, A0=>nx3440, A1=>nx12199);
   ix18984 : inv01 port map ( Y=>nx18603, A=>nx3422);
   reg_nx3446 : nand04_2x port map ( Y=>nx3446, A0=>nx18602, A1=>nx12233, A2
      =>nx12216, A3=>nx18603);
   ix18985 : inv02 port map ( Y=>nx18604, A=>address(4));
   ix18986 : inv02 port map ( Y=>nx18605, A=>address(5));
   ix18987 : inv01 port map ( Y=>nx18606, A=>nx16003);
   ix18988 : inv01 port map ( Y=>nx18607, A=>nx12074);
   ix18989 : inv01 port map ( Y=>nx18608, A=>nx15985);
   ix18990 : inv01 port map ( Y=>nx18609, A=>nx15425);
   ix18991 : inv01 port map ( Y=>nx18610, A=>nx12078);
   ix18992 : aoi43 port map ( Y=>nx18611, A0=>nx18604, A1=>nx18605, A2=>
      nx18606, A3=>nx18607, B0=>nx18608, B1=>nx18609, B2=>nx18610);
   reg_NOT_nx3710 : or03 port map ( Y=>NOT_nx3710, A0=>nx16003, A1=>nx15425, 
      A2=>nx12061);
   ix18993 : inv01 port map ( Y=>nx18612, A=>nx3916);
   ix18994 : nand04_2x port map ( Y=>nx18613, A0=>nx18611, A1=>NOT_nx3710, 
      A2=>nx12002, A3=>nx18612);
   ix18995 : oai43 port map ( Y=>nx18614, A0=>address(4), A1=>address(5), A2
      =>nx12057, A3=>nx16023, B0=>nx15985, B1=>nx12091, B2=>nx15855);
   ix18996 : inv01 port map ( Y=>nx18615, A=>nx18614);
   reg_NOT_nx3748 : or04 port map ( Y=>NOT_nx3748, A0=>address(4), A1=>
      address(5), A2=>nx16043, A3=>nx12044);
   ix18997 : nor02ii port map ( Y=>nx18616, A0=>nx3662, A1=>nx12148);
   ix18998 : nor02_2x port map ( Y=>nx18617, A0=>nx3898, A1=>nx3624);
   ix18999 : nand04_2x port map ( Y=>nx18618, A0=>nx18615, A1=>NOT_nx3748, 
      A2=>nx18616, A3=>nx18617);
   ix19000 : nor03_2x port map ( Y=>nx18619, A0=>nx3580, A1=>nx3598, A2=>
      nx3562);
   ix19001 : or03 port map ( Y=>nx18620, A0=>nx16043, A1=>nx12040, A2=>
      nx15821);
   ix19002 : inv01 port map ( Y=>nx18621, A=>nx3632);
   ix19003 : and03 port map ( Y=>nx18622, A0=>nx18620, A1=>nx12165, A2=>
      nx18621);
   ix19004 : nor02ii port map ( Y=>nx18623, A0=>nx3740, A1=>nx12019);
   ix19005 : nor02ii port map ( Y=>nx18624, A0=>nx3702, A1=>nx11986);
   ix19006 : nand04_2x port map ( Y=>nx18625, A0=>nx18619, A1=>nx18622, A2=>
      nx18623, A3=>nx18624);
   reg_nx11965 : nor04_2x port map ( Y=>nx11965, A0=>nx3446, A1=>nx18613, A2
      =>nx18618, A3=>nx18625);
   ix19007 : nor02ii port map ( Y=>nx18626, A0=>nx8544, A1=>nx14487);
   ix19008 : inv01 port map ( Y=>nx18627, A=>nx8526);
   reg_nx8550 : nand04_2x port map ( Y=>nx8550, A0=>nx18626, A1=>nx14521, A2
      =>nx14504, A3=>nx18627);
   ix19009 : inv02 port map ( Y=>nx18628, A=>address(4));
   ix19010 : inv02 port map ( Y=>nx18629, A=>address(5));
   ix19011 : inv01 port map ( Y=>nx18630, A=>nx16007);
   ix19012 : inv01 port map ( Y=>nx18631, A=>nx14362);
   ix19013 : inv01 port map ( Y=>nx18632, A=>nx15989);
   ix19014 : inv01 port map ( Y=>nx18633, A=>nx15443);
   ix19015 : inv01 port map ( Y=>nx18634, A=>nx14366);
   ix19016 : aoi43 port map ( Y=>nx18635, A0=>nx18628, A1=>nx18629, A2=>
      nx18630, A3=>nx18631, B0=>nx18632, B1=>nx18633, B2=>nx18634);
   reg_NOT_nx8814 : or03 port map ( Y=>NOT_nx8814, A0=>nx16007, A1=>nx15443, 
      A2=>nx14349);
   ix19017 : inv01 port map ( Y=>nx18636, A=>nx9020);
   ix19018 : nand04_2x port map ( Y=>nx18637, A0=>nx18635, A1=>NOT_nx8814, 
      A2=>nx14290, A3=>nx18636);
   ix19019 : oai43 port map ( Y=>nx18638, A0=>address(4), A1=>address(5), A2
      =>nx14345, A3=>nx16027, B0=>nx15989, B1=>nx14379, B2=>nx15865);
   ix19020 : inv01 port map ( Y=>nx18639, A=>nx18638);
   reg_NOT_nx8852 : or04 port map ( Y=>NOT_nx8852, A0=>address(4), A1=>
      address(5), A2=>nx16049, A3=>nx14332);
   ix19021 : nor02ii port map ( Y=>nx18640, A0=>nx8766, A1=>nx14436);
   ix19022 : nor02_2x port map ( Y=>nx18641, A0=>nx9002, A1=>nx8728);
   ix19023 : nand04_2x port map ( Y=>nx18642, A0=>nx18639, A1=>NOT_nx8852, 
      A2=>nx18640, A3=>nx18641);
   ix19024 : nor03_2x port map ( Y=>nx18643, A0=>nx8684, A1=>nx8702, A2=>
      nx8666);
   ix19025 : or03 port map ( Y=>nx18644, A0=>nx16049, A1=>nx14328, A2=>
      nx15829);
   ix19026 : inv01 port map ( Y=>nx18645, A=>nx8736);
   ix19027 : and03 port map ( Y=>nx18646, A0=>nx18644, A1=>nx14453, A2=>
      nx18645);
   ix19028 : nor02ii port map ( Y=>nx18647, A0=>nx8844, A1=>nx14307);
   ix19029 : nor02ii port map ( Y=>nx18648, A0=>nx8806, A1=>nx14274);
   ix19030 : nand04_2x port map ( Y=>nx18649, A0=>nx18643, A1=>nx18646, A2=>
      nx18647, A3=>nx18648);
   reg_nx14253 : nor04_2x port map ( Y=>nx14253, A0=>nx8550, A1=>nx18637, A2
      =>nx18642, A3=>nx18649);
   ix19031 : nor02ii port map ( Y=>nx18650, A0=>nx2802, A1=>nx11913);
   ix19032 : inv01 port map ( Y=>nx18651, A=>nx2784);
   reg_nx2808 : nand04_2x port map ( Y=>nx2808, A0=>nx18650, A1=>nx11947, A2
      =>nx11930, A3=>nx18651);
   ix19033 : inv02 port map ( Y=>nx18652, A=>address(4));
   ix19034 : inv02 port map ( Y=>nx18653, A=>address(5));
   ix19035 : inv01 port map ( Y=>nx18654, A=>nx16003);
   ix19036 : inv01 port map ( Y=>nx18655, A=>nx11788);
   ix19037 : inv01 port map ( Y=>nx18656, A=>nx15985);
   ix19038 : inv01 port map ( Y=>nx18657, A=>nx11792);
   ix19039 : inv01 port map ( Y=>nx18658, A=>nx15423);
   ix19040 : aoi43 port map ( Y=>nx18659, A0=>nx18652, A1=>nx18653, A2=>
      nx18654, A3=>nx18655, B0=>nx18656, B1=>nx18657, B2=>nx18658);
   reg_NOT_nx3072 : or03 port map ( Y=>NOT_nx3072, A0=>nx16003, A1=>nx11775, 
      A2=>nx15421);
   ix19041 : inv01 port map ( Y=>nx18660, A=>nx3278);
   ix19042 : nand04_2x port map ( Y=>nx18661, A0=>nx18659, A1=>NOT_nx3072, 
      A2=>nx11716, A3=>nx18660);
   ix19043 : oai43 port map ( Y=>nx18662, A0=>address(4), A1=>address(5), A2
      =>nx11771, A3=>nx16023, B0=>nx15985, B1=>nx11805, B2=>nx15853);
   ix19044 : inv01 port map ( Y=>nx18663, A=>nx18662);
   reg_NOT_nx3110 : or04 port map ( Y=>NOT_nx3110, A0=>address(4), A1=>
      address(5), A2=>nx16041, A3=>nx11758);
   ix19045 : nor02ii port map ( Y=>nx18664, A0=>nx3024, A1=>nx11862);
   ix19046 : nor02_2x port map ( Y=>nx18665, A0=>nx3260, A1=>nx2986);
   ix19047 : nand04_2x port map ( Y=>nx18666, A0=>nx18663, A1=>NOT_nx3110, 
      A2=>nx18664, A3=>nx18665);
   ix19048 : nor03_2x port map ( Y=>nx18667, A0=>nx2942, A1=>nx2960, A2=>
      nx2924);
   ix19049 : or03 port map ( Y=>nx18668, A0=>nx16041, A1=>nx11754, A2=>
      nx15821);
   ix19050 : inv01 port map ( Y=>nx18669, A=>nx2994);
   ix19051 : and03 port map ( Y=>nx18670, A0=>nx18668, A1=>nx11733, A2=>
      nx18669);
   ix19052 : nor02ii port map ( Y=>nx18671, A0=>nx3102, A1=>nx11879);
   ix19053 : nor02ii port map ( Y=>nx18672, A0=>nx3064, A1=>nx11700);
   ix19054 : nand04_2x port map ( Y=>nx18673, A0=>nx18667, A1=>nx18670, A2=>
      nx18671, A3=>nx18672);
   reg_nx11679 : nor04_2x port map ( Y=>nx11679, A0=>nx2808, A1=>nx18661, A2
      =>nx18666, A3=>nx18673);
   ix19055 : nor02ii port map ( Y=>nx18674, A0=>nx6630, A1=>nx13629);
   ix19056 : inv01 port map ( Y=>nx18675, A=>nx6612);
   reg_nx6636 : nand04_2x port map ( Y=>nx6636, A0=>nx18674, A1=>nx13663, A2
      =>nx13646, A3=>nx18675);
   ix19057 : inv02 port map ( Y=>nx18676, A=>address(4));
   ix19058 : inv02 port map ( Y=>nx18677, A=>address(5));
   ix19059 : inv01 port map ( Y=>nx18678, A=>nx16005);
   ix19060 : inv01 port map ( Y=>nx18679, A=>nx13504);
   ix19061 : inv01 port map ( Y=>nx18680, A=>nx15987);
   ix19062 : inv01 port map ( Y=>nx18681, A=>nx15435);
   ix19063 : inv01 port map ( Y=>nx18682, A=>nx13508);
   ix19064 : aoi43 port map ( Y=>nx18683, A0=>nx18676, A1=>nx18677, A2=>
      nx18678, A3=>nx18679, B0=>nx18680, B1=>nx18681, B2=>nx18682);
   reg_NOT_nx6900 : or03 port map ( Y=>NOT_nx6900, A0=>nx16005, A1=>nx15435, 
      A2=>nx13491);
   ix19065 : inv01 port map ( Y=>nx18684, A=>nx7106);
   ix19066 : nand04_2x port map ( Y=>nx18685, A0=>nx18683, A1=>NOT_nx6900, 
      A2=>nx13432, A3=>nx18684);
   ix19067 : oai43 port map ( Y=>nx18686, A0=>address(4), A1=>address(5), A2
      =>nx13487, A3=>nx16025, B0=>nx15987, B1=>nx13521, B2=>nx15861);
   ix19068 : inv01 port map ( Y=>nx18687, A=>nx18686);
   reg_NOT_nx6938 : or04 port map ( Y=>NOT_nx6938, A0=>address(4), A1=>
      address(5), A2=>nx16047, A3=>nx13474);
   ix19069 : nor02ii port map ( Y=>nx18688, A0=>nx6852, A1=>nx13578);
   ix19070 : nor02_2x port map ( Y=>nx18689, A0=>nx7088, A1=>nx6814);
   ix19071 : nand04_2x port map ( Y=>nx18690, A0=>nx18687, A1=>NOT_nx6938, 
      A2=>nx18688, A3=>nx18689);
   ix19072 : nor03_2x port map ( Y=>nx18691, A0=>nx6770, A1=>nx6788, A2=>
      nx6752);
   ix19073 : or03 port map ( Y=>nx18692, A0=>nx16047, A1=>nx13470, A2=>
      nx15825);
   ix19074 : inv01 port map ( Y=>nx18693, A=>nx6822);
   ix19075 : and03 port map ( Y=>nx18694, A0=>nx18692, A1=>nx13449, A2=>
      nx18693);
   ix19076 : nor02ii port map ( Y=>nx18695, A0=>nx6930, A1=>nx13595);
   ix19077 : nor02ii port map ( Y=>nx18696, A0=>nx6892, A1=>nx13416);
   ix19078 : nand04_2x port map ( Y=>nx18697, A0=>nx18691, A1=>nx18694, A2=>
      nx18695, A3=>nx18696);
   reg_nx13395 : nor04_2x port map ( Y=>nx13395, A0=>nx6636, A1=>nx18685, A2
      =>nx18690, A3=>nx18697);
   ix19079 : nor02ii port map ( Y=>nx18698, A0=>nx7906, A1=>nx14201);
   ix19080 : inv01 port map ( Y=>nx18699, A=>nx7888);
   reg_nx7912 : nand04_2x port map ( Y=>nx7912, A0=>nx18698, A1=>nx14235, A2
      =>nx14218, A3=>nx18699);
   ix19081 : inv02 port map ( Y=>nx18700, A=>address(4));
   ix19082 : inv02 port map ( Y=>nx18701, A=>address(5));
   ix19083 : inv01 port map ( Y=>nx18702, A=>nx16007);
   ix19084 : inv01 port map ( Y=>nx18703, A=>nx14076);
   ix19085 : inv01 port map ( Y=>nx18704, A=>nx15989);
   ix19086 : inv01 port map ( Y=>nx18705, A=>nx15441);
   ix19087 : inv01 port map ( Y=>nx18706, A=>nx14080);
   ix19088 : aoi43 port map ( Y=>nx18707, A0=>nx18700, A1=>nx18701, A2=>
      nx18702, A3=>nx18703, B0=>nx18704, B1=>nx18705, B2=>nx18706);
   reg_NOT_nx8176 : or03 port map ( Y=>NOT_nx8176, A0=>nx16007, A1=>nx15441, 
      A2=>nx14063);
   ix19089 : inv01 port map ( Y=>nx18708, A=>nx8382);
   ix19090 : nand04_2x port map ( Y=>nx18709, A0=>nx18707, A1=>NOT_nx8176, 
      A2=>nx14004, A3=>nx18708);
   ix19091 : oai43 port map ( Y=>nx18710, A0=>address(4), A1=>address(5), A2
      =>nx14059, A3=>nx16027, B0=>nx15989, B1=>nx14093, B2=>nx15865);
   ix19092 : inv01 port map ( Y=>nx18711, A=>nx18710);
   reg_NOT_nx8214 : or04 port map ( Y=>NOT_nx8214, A0=>address(4), A1=>
      address(5), A2=>nx16049, A3=>nx14046);
   ix19093 : nor02ii port map ( Y=>nx18712, A0=>nx8128, A1=>nx14150);
   ix19094 : nor02_2x port map ( Y=>nx18713, A0=>nx8364, A1=>nx8090);
   ix19095 : nand04_2x port map ( Y=>nx18714, A0=>nx18711, A1=>NOT_nx8214, 
      A2=>nx18712, A3=>nx18713);
   ix19096 : nor03_2x port map ( Y=>nx18715, A0=>nx8046, A1=>nx8064, A2=>
      nx8028);
   ix19097 : or03 port map ( Y=>nx18716, A0=>nx16049, A1=>nx14042, A2=>
      nx15827);
   ix19098 : inv01 port map ( Y=>nx18717, A=>nx8098);
   ix19099 : and03 port map ( Y=>nx18718, A0=>nx18716, A1=>nx14167, A2=>
      nx18717);
   ix19100 : nor02ii port map ( Y=>nx18719, A0=>nx8206, A1=>nx14021);
   ix19101 : nor02ii port map ( Y=>nx18720, A0=>nx8168, A1=>nx13988);
   ix19102 : nand04_2x port map ( Y=>nx18721, A0=>nx18715, A1=>nx18718, A2=>
      nx18719, A3=>nx18720);
   reg_nx13967 : nor04_2x port map ( Y=>nx13967, A0=>nx7912, A1=>nx18709, A2
      =>nx18714, A3=>nx18721);
   ix19103 : nor02ii port map ( Y=>nx18722, A0=>nx4078, A1=>nx12485);
   ix19104 : inv01 port map ( Y=>nx18723, A=>nx4060);
   reg_nx4084 : nand04_2x port map ( Y=>nx4084, A0=>nx18722, A1=>nx12519, A2
      =>nx12502, A3=>nx18723);
   ix19105 : inv02 port map ( Y=>nx18724, A=>address(4));
   ix19106 : inv02 port map ( Y=>nx18725, A=>address(5));
   ix19107 : inv01 port map ( Y=>nx18726, A=>nx16003);
   ix19108 : inv01 port map ( Y=>nx18727, A=>nx12360);
   ix19109 : inv01 port map ( Y=>nx18728, A=>nx15985);
   ix19110 : inv01 port map ( Y=>nx18729, A=>nx15427);
   ix19111 : inv01 port map ( Y=>nx18730, A=>nx12364);
   ix19112 : aoi43 port map ( Y=>nx18731, A0=>nx18724, A1=>nx18725, A2=>
      nx18726, A3=>nx18727, B0=>nx18728, B1=>nx18729, B2=>nx18730);
   reg_NOT_nx4348 : or03 port map ( Y=>NOT_nx4348, A0=>nx16003, A1=>nx15427, 
      A2=>nx12347);
   ix19113 : inv01 port map ( Y=>nx18732, A=>nx4554);
   ix19114 : nand04_2x port map ( Y=>nx18733, A0=>nx18731, A1=>NOT_nx4348, 
      A2=>nx12288, A3=>nx18732);
   ix19115 : oai43 port map ( Y=>nx18734, A0=>address(4), A1=>address(5), A2
      =>nx12343, A3=>nx16023, B0=>nx15985, B1=>nx12377, B2=>nx15855);
   ix19116 : inv01 port map ( Y=>nx18735, A=>nx18734);
   reg_NOT_nx4386 : or04 port map ( Y=>NOT_nx4386, A0=>address(4), A1=>
      address(5), A2=>nx16043, A3=>nx12330);
   ix19117 : nor02ii port map ( Y=>nx18736, A0=>nx4300, A1=>nx12434);
   ix19118 : nor02_2x port map ( Y=>nx18737, A0=>nx4536, A1=>nx4262);
   ix19119 : nand04_2x port map ( Y=>nx18738, A0=>nx18735, A1=>NOT_nx4386, 
      A2=>nx18736, A3=>nx18737);
   ix19120 : nor03_2x port map ( Y=>nx18739, A0=>nx4218, A1=>nx4236, A2=>
      nx4200);
   ix19121 : or03 port map ( Y=>nx18740, A0=>nx16043, A1=>nx12326, A2=>
      nx15823);
   ix19122 : inv01 port map ( Y=>nx18741, A=>nx4270);
   ix19123 : and03 port map ( Y=>nx18742, A0=>nx18740, A1=>nx12451, A2=>
      nx18741);
   ix19124 : nor02ii port map ( Y=>nx18743, A0=>nx4378, A1=>nx12305);
   ix19125 : nor02ii port map ( Y=>nx18744, A0=>nx4340, A1=>nx12272);
   ix19126 : nand04_2x port map ( Y=>nx18745, A0=>nx18739, A1=>nx18742, A2=>
      nx18743, A3=>nx18744);
   reg_nx12251 : nor04_2x port map ( Y=>nx12251, A0=>nx4084, A1=>nx18733, A2
      =>nx18738, A3=>nx18745);
   ix19127 : nor02ii port map ( Y=>nx18746, A0=>nx2164, A1=>nx11627);
   ix19128 : inv01 port map ( Y=>nx18747, A=>nx2146);
   reg_nx2170 : nand04_2x port map ( Y=>nx2170, A0=>nx18746, A1=>nx11661, A2
      =>nx11644, A3=>nx18747);
   ix19129 : inv02 port map ( Y=>nx18748, A=>address(4));
   ix19130 : inv02 port map ( Y=>nx18749, A=>address(5));
   ix19131 : inv01 port map ( Y=>nx18750, A=>nx16001);
   ix19132 : inv01 port map ( Y=>nx18751, A=>nx11502);
   ix19133 : inv01 port map ( Y=>nx18752, A=>nx15983);
   ix19134 : inv01 port map ( Y=>nx18753, A=>nx15419);
   ix19135 : inv01 port map ( Y=>nx18754, A=>nx11506);
   ix19136 : aoi43 port map ( Y=>nx18755, A0=>nx18748, A1=>nx18749, A2=>
      nx18750, A3=>nx18751, B0=>nx18752, B1=>nx18753, B2=>nx18754);
   reg_NOT_nx2434 : or03 port map ( Y=>NOT_nx2434, A0=>nx16001, A1=>nx15419, 
      A2=>nx11489);
   ix19137 : inv01 port map ( Y=>nx18756, A=>nx2640);
   ix19138 : nand04_2x port map ( Y=>nx18757, A0=>nx18755, A1=>NOT_nx2434, 
      A2=>nx11430, A3=>nx18756);
   ix19139 : nor03_2x port map ( Y=>nx18758, A0=>nx2304, A1=>nx2322, A2=>
      nx2286);
   reg_NOT_nx2364 : or03 port map ( Y=>NOT_nx2364, A0=>nx15983, A1=>nx11519, 
      A2=>nx15851);
   ix19140 : or03 port map ( Y=>nx18759, A0=>nx16041, A1=>nx11468, A2=>
      nx15819);
   ix19141 : nor02ii port map ( Y=>nx18760, A0=>nx2356, A1=>nx11447);
   ix19142 : nand04_2x port map ( Y=>nx18761, A0=>nx18758, A1=>NOT_nx2364, 
      A2=>nx18759, A3=>nx18760);
   reg_NOT_nx2472 : or04 port map ( Y=>NOT_nx2472, A0=>address(4), A1=>
      address(5), A2=>nx16041, A3=>nx11472);
   reg_NOT_nx2442 : or04 port map ( Y=>NOT_nx2442, A0=>address(4), A1=>
      address(5), A2=>nx11485, A3=>nx16021);
   ix19143 : inv01 port map ( Y=>nx18762, A=>nx11593);
   ix19144 : inv01 port map ( Y=>nx18763, A=>nx11414);
   ix19145 : nor04_2x port map ( Y=>nx18764, A0=>nx18762, A1=>nx2464, A2=>
      nx18763, A3=>nx2426);
   ix19146 : nand04_2x port map ( Y=>nx18765, A0=>NOT_nx2472, A1=>nx18932, 
      A2=>NOT_nx2442, A3=>nx18764);
   reg_nx11393 : nor04_2x port map ( Y=>nx11393, A0=>nx2170, A1=>nx18757, A2
      =>nx18761, A3=>nx18765);
   ix19147 : nor02ii port map ( Y=>nx18766, A0=>nx5354, A1=>nx13057);
   ix19148 : inv01 port map ( Y=>nx18767, A=>nx5336);
   reg_nx5360 : nand04_2x port map ( Y=>nx5360, A0=>nx18766, A1=>nx13091, A2
      =>nx13074, A3=>nx18767);
   ix19149 : inv02 port map ( Y=>nx18768, A=>address(4));
   ix19150 : inv02 port map ( Y=>nx18769, A=>address(5));
   ix19151 : inv01 port map ( Y=>nx18770, A=>nx16005);
   ix19152 : inv01 port map ( Y=>nx18771, A=>nx12932);
   ix19153 : inv01 port map ( Y=>nx18772, A=>nx15987);
   ix19154 : inv01 port map ( Y=>nx18773, A=>nx15431);
   ix19155 : inv01 port map ( Y=>nx18774, A=>nx12936);
   ix19156 : aoi43 port map ( Y=>nx18775, A0=>nx18768, A1=>nx18769, A2=>
      nx18770, A3=>nx18771, B0=>nx18772, B1=>nx18773, B2=>nx18774);
   reg_NOT_nx5624 : or03 port map ( Y=>NOT_nx5624, A0=>nx16005, A1=>nx15431, 
      A2=>nx12919);
   ix19157 : inv01 port map ( Y=>nx18776, A=>nx5830);
   ix19158 : nand04_2x port map ( Y=>nx18777, A0=>nx18775, A1=>NOT_nx5624, 
      A2=>nx12860, A3=>nx18776);
   ix19159 : oai43 port map ( Y=>nx18778, A0=>address(4), A1=>address(5), A2
      =>nx12915, A3=>nx16025, B0=>nx15987, B1=>nx12949, B2=>nx15859);
   ix19160 : inv01 port map ( Y=>nx18779, A=>nx18778);
   reg_NOT_nx5662 : or04 port map ( Y=>NOT_nx5662, A0=>address(4), A1=>
      address(5), A2=>nx16045, A3=>nx12902);
   ix19161 : nor02ii port map ( Y=>nx18780, A0=>nx5576, A1=>nx13006);
   ix19162 : nor02_2x port map ( Y=>nx18781, A0=>nx5812, A1=>nx5538);
   ix19163 : nand04_2x port map ( Y=>nx18782, A0=>nx18779, A1=>NOT_nx5662, 
      A2=>nx18780, A3=>nx18781);
   ix19164 : nor03_2x port map ( Y=>nx18783, A0=>nx5494, A1=>nx5512, A2=>
      nx5476);
   ix19165 : or03 port map ( Y=>nx18784, A0=>nx16045, A1=>nx12898, A2=>
      nx15825);
   ix19166 : inv01 port map ( Y=>nx18785, A=>nx5546);
   ix19167 : and03 port map ( Y=>nx18786, A0=>nx18784, A1=>nx13023, A2=>
      nx18785);
   ix19168 : nor02ii port map ( Y=>nx18787, A0=>nx5654, A1=>nx12877);
   ix19169 : nor02ii port map ( Y=>nx18788, A0=>nx5616, A1=>nx12844);
   ix19170 : nand04_2x port map ( Y=>nx18789, A0=>nx18783, A1=>nx18786, A2=>
      nx18787, A3=>nx18788);
   reg_nx12823 : nor04_2x port map ( Y=>nx12823, A0=>nx5360, A1=>nx18777, A2
      =>nx18782, A3=>nx18789);
   ix19171 : nor02ii port map ( Y=>nx18790, A0=>nx5992, A1=>nx13343);
   ix19172 : inv01 port map ( Y=>nx18791, A=>nx5974);
   reg_nx5998 : nand04_2x port map ( Y=>nx5998, A0=>nx18790, A1=>nx13377, A2
      =>nx13360, A3=>nx18791);
   ix19173 : inv02 port map ( Y=>nx18792, A=>address(4));
   ix19174 : inv02 port map ( Y=>nx18793, A=>address(5));
   ix19175 : inv01 port map ( Y=>nx18794, A=>nx16005);
   ix19176 : inv01 port map ( Y=>nx18795, A=>nx13218);
   ix19177 : inv01 port map ( Y=>nx18796, A=>nx15987);
   ix19178 : inv01 port map ( Y=>nx18797, A=>nx15433);
   ix19179 : inv01 port map ( Y=>nx18798, A=>nx13222);
   ix19180 : aoi43 port map ( Y=>nx18799, A0=>nx18792, A1=>nx18793, A2=>
      nx18794, A3=>nx18795, B0=>nx18796, B1=>nx18797, B2=>nx18798);
   reg_NOT_nx6262 : or03 port map ( Y=>NOT_nx6262, A0=>nx16005, A1=>nx15433, 
      A2=>nx13205);
   ix19181 : inv01 port map ( Y=>nx18800, A=>nx6468);
   ix19182 : nand04_2x port map ( Y=>nx18801, A0=>nx18799, A1=>NOT_nx6262, 
      A2=>nx13146, A3=>nx18800);
   ix19183 : oai43 port map ( Y=>nx18802, A0=>address(4), A1=>address(5), A2
      =>nx13201, A3=>nx16025, B0=>nx15987, B1=>nx13235, B2=>nx15861);
   ix19184 : inv01 port map ( Y=>nx18803, A=>nx18802);
   reg_NOT_nx6300 : or04 port map ( Y=>NOT_nx6300, A0=>address(4), A1=>
      address(5), A2=>nx16045, A3=>nx13188);
   ix19185 : nor02ii port map ( Y=>nx18804, A0=>nx6214, A1=>nx13292);
   ix19186 : nor02_2x port map ( Y=>nx18805, A0=>nx6450, A1=>nx6176);
   ix19187 : nand04_2x port map ( Y=>nx18806, A0=>nx18803, A1=>NOT_nx6300, 
      A2=>nx18804, A3=>nx18805);
   ix19188 : nor03_2x port map ( Y=>nx18807, A0=>nx6132, A1=>nx6150, A2=>
      nx6114);
   ix19189 : or03 port map ( Y=>nx18808, A0=>nx16045, A1=>nx13184, A2=>
      nx15825);
   ix19190 : inv01 port map ( Y=>nx18809, A=>nx6184);
   ix19191 : and03 port map ( Y=>nx18810, A0=>nx18808, A1=>nx13309, A2=>
      nx18809);
   ix19192 : nor02ii port map ( Y=>nx18811, A0=>nx6292, A1=>nx13163);
   ix19193 : nor02ii port map ( Y=>nx18812, A0=>nx6254, A1=>nx13130);
   ix19194 : nand04_2x port map ( Y=>nx18813, A0=>nx18807, A1=>nx18810, A2=>
      nx18811, A3=>nx18812);
   reg_nx13109 : nor04_2x port map ( Y=>nx13109, A0=>nx5998, A1=>nx18801, A2
      =>nx18806, A3=>nx18813);
   ix19195 : nor02ii port map ( Y=>nx18814, A0=>nx4716, A1=>nx12771);
   ix19196 : inv01 port map ( Y=>nx18815, A=>nx4698);
   reg_nx4722 : nand04_2x port map ( Y=>nx4722, A0=>nx18814, A1=>nx12805, A2
      =>nx12788, A3=>nx18815);
   ix19197 : nor03_2x port map ( Y=>nx18816, A0=>nx15985, A1=>nx15429, A2=>
      nx12650);
   ix19198 : nor03_2x port map ( Y=>nx18817, A0=>nx16043, A1=>nx12612, A2=>
      nx15823);
   ix19199 : inv01 port map ( Y=>nx18818, A=>nx12737);
   ix19200 : nor04_2x port map ( Y=>nx18819, A0=>nx18816, A1=>nx18817, A2=>
      nx18818, A3=>nx4908);
   reg_NOT_nx4986 : or03 port map ( Y=>NOT_nx4986, A0=>nx16003, A1=>nx15429, 
      A2=>nx12633);
   ix19201 : inv01 port map ( Y=>nx18820, A=>nx5192);
   ix19202 : nand04_2x port map ( Y=>nx18821, A0=>nx18819, A1=>NOT_nx4986, 
      A2=>nx12574, A3=>nx18820);
   ix19203 : oai43 port map ( Y=>nx18822, A0=>nx12629, A1=>nx16025, A2=>
      address(4), A3=>address(5), B0=>nx15987, B1=>nx12663, B2=>nx15857);
   ix19204 : inv01 port map ( Y=>nx18823, A=>nx18822);
   reg_NOT_nx5024 : or04 port map ( Y=>NOT_nx5024, A0=>address(4), A1=>
      address(5), A2=>nx12616, A3=>nx16045);
   ix19205 : nor02ii port map ( Y=>nx18824, A0=>nx4938, A1=>nx12720);
   ix19206 : nor02_2x port map ( Y=>nx18825, A0=>nx5174, A1=>nx4900);
   ix19207 : nand04_2x port map ( Y=>nx18826, A0=>nx18823, A1=>NOT_nx5024, 
      A2=>nx18824, A3=>nx18825);
   ix19208 : nor03_2x port map ( Y=>nx18827, A0=>nx4856, A1=>nx4874, A2=>
      nx4838);
   reg_NOT_nx4954 : or04 port map ( Y=>NOT_nx4954, A0=>address(4), A1=>
      address(5), A2=>nx12646, A3=>nx16005);
   ix19209 : nor02ii port map ( Y=>nx18828, A0=>nx5016, A1=>nx12591);
   ix19210 : nor02ii port map ( Y=>nx18829, A0=>nx4978, A1=>nx12558);
   ix19211 : nand04_2x port map ( Y=>nx18830, A0=>nx18827, A1=>NOT_nx4954, 
      A2=>nx18828, A3=>nx18829);
   reg_nx12537 : nor04_2x port map ( Y=>nx12537, A0=>nx4722, A1=>nx18821, A2
      =>nx18826, A3=>nx18830);
   ix19212 : nor02ii port map ( Y=>nx18831, A0=>nx378, A1=>nx11016);
   ix19213 : inv01 port map ( Y=>nx18832, A=>nx338);
   reg_nx384 : nand04_2x port map ( Y=>nx384, A0=>nx18831, A1=>nx11077, A2=>
      nx11048, A3=>nx18832);
   ix19214 : inv02 port map ( Y=>nx18833, A=>address(4));
   ix19215 : inv02 port map ( Y=>nx18834, A=>address(5));
   ix19216 : inv01 port map ( Y=>nx18835, A=>nx16001);
   ix19217 : inv01 port map ( Y=>nx18836, A=>nx10762);
   ix19218 : inv01 port map ( Y=>nx18837, A=>nx15983);
   ix19219 : inv01 port map ( Y=>nx18838, A=>nx17141);
   ix19220 : inv01 port map ( Y=>nx18839, A=>nx10769);
   ix19221 : aoi43 port map ( Y=>nx18840, A0=>nx18833, A1=>nx18834, A2=>
      nx18835, A3=>nx18836, B0=>nx18837, B1=>nx18838, B2=>nx18839);
   reg_NOT_nx940 : or03 port map ( Y=>NOT_nx940, A0=>nx16001, A1=>nx17141, 
      A2=>nx10731);
   ix19222 : inv01 port map ( Y=>nx18841, A=>nx1364);
   ix19223 : nand04_2x port map ( Y=>nx18842, A0=>nx18840, A1=>NOT_nx940, A2
      =>nx10615, A3=>nx18841);
   ix19224 : nor03_2x port map ( Y=>nx18843, A0=>nx672, A1=>nx714, A2=>nx634
   );
   reg_NOT_nx798 : or03 port map ( Y=>NOT_nx798, A0=>nx15983, A1=>nx10801, 
      A2=>nx15849);
   ix19225 : or03 port map ( Y=>nx18844, A0=>nx16039, A1=>nx10692, A2=>
      nx15819);
   ix19226 : nor02ii port map ( Y=>nx18845, A0=>nx778, A1=>nx10651);
   ix19227 : nand04_2x port map ( Y=>nx18846, A0=>nx18843, A1=>NOT_nx798, A2
      =>nx18844, A3=>nx18845);
   reg_NOT_nx1022 : or04 port map ( Y=>NOT_nx1022, A0=>address(4), A1=>
      address(5), A2=>nx16039, A3=>nx10699);
   reg_NOT_nx960 : or04 port map ( Y=>NOT_nx960, A0=>address(4), A1=>
      address(5), A2=>nx10724, A3=>nx16021);
   ix19228 : inv01 port map ( Y=>nx18847, A=>nx10951);
   ix19229 : inv01 port map ( Y=>nx18848, A=>nx10571);
   ix19230 : nor04_2x port map ( Y=>nx18849, A0=>nx18847, A1=>nx1002, A2=>
      nx18848, A3=>nx922);
   ix19231 : nand04_2x port map ( Y=>nx18850, A0=>NOT_nx1022, A1=>nx18948, 
      A2=>NOT_nx960, A3=>nx18849);
   reg_nx10491 : nor04_2x port map ( Y=>nx10491, A0=>nx384, A1=>nx18842, A2
      =>nx18846, A3=>nx18850);
   ix19232 : nor02ii port map ( Y=>nx18851, A0=>nx1526, A1=>nx11341);
   ix19233 : inv01 port map ( Y=>nx18852, A=>nx1508);
   reg_nx1532 : nand04_2x port map ( Y=>nx1532, A0=>nx18851, A1=>nx11375, A2
      =>nx11358, A3=>nx18852);
   ix19234 : inv02 port map ( Y=>nx18853, A=>address(4));
   ix19235 : inv02 port map ( Y=>nx18854, A=>address(5));
   ix19236 : inv01 port map ( Y=>nx18855, A=>nx16001);
   ix19237 : inv01 port map ( Y=>nx18856, A=>nx11216);
   ix19238 : inv01 port map ( Y=>nx18857, A=>nx15983);
   ix19239 : inv01 port map ( Y=>nx18858, A=>nx15417);
   ix19240 : inv01 port map ( Y=>nx18859, A=>nx11220);
   ix19241 : aoi43 port map ( Y=>nx18860, A0=>nx18853, A1=>nx18854, A2=>
      nx18855, A3=>nx18856, B0=>nx18857, B1=>nx18858, B2=>nx18859);
   reg_NOT_nx1796 : or03 port map ( Y=>NOT_nx1796, A0=>nx16001, A1=>nx15417, 
      A2=>nx11203);
   ix19242 : inv01 port map ( Y=>nx18861, A=>nx2002);
   ix19243 : nand04_2x port map ( Y=>nx18862, A0=>nx18860, A1=>NOT_nx1796, 
      A2=>nx11144, A3=>nx18861);
   ix19244 : nor03_2x port map ( Y=>nx18863, A0=>nx1666, A1=>nx1684, A2=>
      nx1648);
   reg_NOT_nx1726 : or03 port map ( Y=>NOT_nx1726, A0=>nx15983, A1=>nx11233, 
      A2=>nx15851);
   ix19245 : or03 port map ( Y=>nx18864, A0=>nx16039, A1=>nx11182, A2=>
      nx15819);
   ix19246 : nor02ii port map ( Y=>nx18865, A0=>nx1718, A1=>nx11161);
   ix19247 : nand04_2x port map ( Y=>nx18866, A0=>nx18863, A1=>NOT_nx1726, 
      A2=>nx18864, A3=>nx18865);
   reg_NOT_nx1834 : or04 port map ( Y=>NOT_nx1834, A0=>address(4), A1=>
      address(5), A2=>nx16039, A3=>nx11186);
   reg_NOT_nx1804 : or04 port map ( Y=>NOT_nx1804, A0=>address(4), A1=>
      address(5), A2=>nx11199, A3=>nx16021);
   ix19248 : inv01 port map ( Y=>nx18867, A=>nx11307);
   ix19249 : inv01 port map ( Y=>nx18868, A=>nx11128);
   ix19250 : nor04_2x port map ( Y=>nx18869, A0=>nx18867, A1=>nx1826, A2=>
      nx18868, A3=>nx1788);
   ix19251 : nand04_2x port map ( Y=>nx18870, A0=>NOT_nx1834, A1=>nx18940, 
      A2=>NOT_nx1804, A3=>nx18869);
   reg_nx11107 : nor04_2x port map ( Y=>nx11107, A0=>nx1532, A1=>nx18862, A2
      =>nx18866, A3=>nx18870);
   ix19252 : nor02ii port map ( Y=>nx18871, A0=>nx9182, A1=>nx14773);
   ix19253 : inv01 port map ( Y=>nx18872, A=>nx9164);
   reg_nx9188 : nand04_2x port map ( Y=>nx9188, A0=>nx18871, A1=>nx14807, A2
      =>nx14790, A3=>nx18872);
   ix19254 : oai33 port map ( Y=>nx18873, A0=>nx15991, A1=>nx14665, A2=>
      nx15867, B0=>nx15989, B1=>nx15445, B2=>nx14652);
   ix19255 : inv01 port map ( Y=>nx18874, A=>nx18873);
   reg_NOT_nx9452 : or03 port map ( Y=>NOT_nx9452, A0=>nx16007, A1=>nx15445, 
      A2=>nx14635);
   ix19256 : inv01 port map ( Y=>nx18875, A=>nx9658);
   ix19257 : nand04_2x port map ( Y=>nx18876, A0=>nx18874, A1=>NOT_nx9452, 
      A2=>nx14576, A3=>nx18875);
   ix19258 : nor03_2x port map ( Y=>nx18877, A0=>nx9322, A1=>nx9340, A2=>
      nx9304);
   reg_NOT_nx9420 : or04 port map ( Y=>NOT_nx9420, A0=>address(4), A1=>
      address(5), A2=>nx14648, A3=>nx16009);
   ix19259 : or03 port map ( Y=>nx18878, A0=>nx16049, A1=>nx14614, A2=>
      nx15829);
   ix19260 : nor02ii port map ( Y=>nx18879, A0=>nx9374, A1=>nx14739);
   ix19261 : nand04_2x port map ( Y=>nx18880, A0=>nx18877, A1=>NOT_nx9420, 
      A2=>nx18878, A3=>nx18879);
   ix19262 : nor04_2x port map ( Y=>nx18881, A0=>address(4), A1=>address(5), 
      A2=>nx14618, A3=>nx16051);
   ix19263 : nor04_2x port map ( Y=>nx18882, A0=>address(4), A1=>address(5), 
      A2=>nx14631, A3=>nx16029);
   ix19264 : nor02_2x port map ( Y=>nx18883, A0=>nx18881, A1=>nx18882);
   ix19265 : nor02ii port map ( Y=>nx18884, A0=>nx9482, A1=>nx14593);
   ix19266 : nor02ii port map ( Y=>nx18885, A0=>nx9444, A1=>nx14560);
   ix19267 : nand04_2x port map ( Y=>nx18886, A0=>nx18883, A1=>nx18953, A2=>
      nx18884, A3=>nx18885);
   reg_nx14539 : nor04_2x port map ( Y=>nx14539, A0=>nx9188, A1=>nx18876, A2
      =>nx18880, A3=>nx18886);
   ix19268 : inv01 port map ( Y=>nx18887, A=>nx15362);
   ix19269 : nor03_2x port map ( Y=>nx18888, A0=>nx10458, A1=>nx18887, A2=>
      nx10440);
   reg_nx10464 : nand03_2x port map ( Y=>nx10464, A0=>nx18888, A1=>nx15345, 
      A2=>nx15379);
   ix19270 : nor03_2x port map ( Y=>nx18889, A0=>nx16009, A1=>nx15207, A2=>
      nx15449);
   ix19271 : inv01 port map ( Y=>nx18890, A=>nx15311);
   ix19272 : nor03_2x port map ( Y=>nx18891, A0=>nx18889, A1=>nx18890, A2=>
      nx10934);
   reg_NOT_nx10688 : or03 port map ( Y=>NOT_nx10688, A0=>nx15991, A1=>
      nx15449, A2=>nx15224);
   ix19273 : or03 port map ( Y=>nx18892, A0=>nx16051, A1=>nx15186, A2=>
      nx15831);
   ix19274 : nor02ii port map ( Y=>nx18893, A0=>nx10650, A1=>nx15165);
   ix19275 : nand04_2x port map ( Y=>nx18894, A0=>nx18891, A1=>NOT_nx10688, 
      A2=>nx18892, A3=>nx18893);
   ix19276 : nor02_2x port map ( Y=>nx18895, A0=>address(4), A1=>address(5)
   );
   ix19277 : nor02_2x port map ( Y=>nx18896, A0=>nx15203, A1=>nx16029);
   ix19278 : nor02_2x port map ( Y=>nx18897, A0=>nx16051, A1=>nx15190);
   ix19279 : oai43 port map ( Y=>nx18898, A0=>address(4), A1=>address(5), A2
      =>nx16009, A3=>nx15220, B0=>nx15991, B1=>nx15237, B2=>nx15871);
   ix19280 : ao221 port map ( Y=>nx18899, A0=>nx18895, A1=>nx18896, B0=>
      nx18895, B1=>nx18897, C0=>nx18898);
   ix19281 : nor03_2x port map ( Y=>nx18900, A0=>nx10580, A1=>nx10616, A2=>
      nx10598);
   ix19282 : nor04_2x port map ( Y=>nx18901, A0=>nx10680, A1=>nx10642, A2=>
      nx10916, A3=>nx10720);
   ix19283 : and02 port map ( Y=>nx18902, A0=>nx15148, A1=>nx15294);
   ix19284 : nor02ii port map ( Y=>nx18903, A0=>nx10758, A1=>nx15132);
   ix19285 : nand04_2x port map ( Y=>nx18904, A0=>nx18900, A1=>nx18901, A2=>
      nx18902, A3=>nx18903);
   reg_nx15111 : nor04_2x port map ( Y=>nx15111, A0=>nx10464, A1=>nx18894, 
      A2=>nx18899, A3=>nx18904);
   ix19286 : nor02ii port map ( Y=>nx18905, A0=>nx9820, A1=>nx15059);
   ix19287 : inv01 port map ( Y=>nx18906, A=>nx9802);
   reg_nx9826 : nand04_2x port map ( Y=>nx9826, A0=>nx18905, A1=>nx15093, A2
      =>nx15076, A3=>nx18906);
   ix19288 : nor03_2x port map ( Y=>nx18907, A0=>nx15991, A1=>nx15447, A2=>
      nx14938);
   ix19289 : nor03_2x port map ( Y=>nx18908, A0=>nx16051, A1=>nx14900, A2=>
      nx15831);
   ix19290 : inv01 port map ( Y=>nx18909, A=>nx14879);
   ix19291 : nor04_2x port map ( Y=>nx18910, A0=>nx18907, A1=>nx18908, A2=>
      nx18909, A3=>nx10012);
   reg_NOT_nx10090 : or03 port map ( Y=>NOT_nx10090, A0=>nx16009, A1=>
      nx15447, A2=>nx14921);
   ix19292 : inv01 port map ( Y=>nx18911, A=>nx10296);
   ix19293 : nand04_2x port map ( Y=>nx18912, A0=>nx18910, A1=>NOT_nx10090, 
      A2=>nx14862, A3=>nx18911);
   ix19294 : nor02_2x port map ( Y=>nx18913, A0=>address(4), A1=>address(5)
   );
   ix19295 : nor02_2x port map ( Y=>nx18914, A0=>nx14917, A1=>nx16029);
   ix19296 : nor02_2x port map ( Y=>nx18915, A0=>nx16051, A1=>nx14904);
   ix19297 : oai43 port map ( Y=>nx18916, A0=>address(4), A1=>address(5), A2
      =>nx16009, A3=>nx14934, B0=>nx15991, B1=>nx14951, B2=>nx15869);
   ix19298 : ao221 port map ( Y=>nx18917, A0=>nx18913, A1=>nx18914, B0=>
      nx18913, B1=>nx18915, C0=>nx18916);
   ix19299 : nor03_2x port map ( Y=>nx18918, A0=>nx9942, A1=>nx9978, A2=>
      nx9960);
   ix19300 : inv01 port map ( Y=>nx18919, A=>nx15025);
   ix19301 : nor04_2x port map ( Y=>nx18920, A0=>nx18919, A1=>nx10004, A2=>
      nx10278, A3=>nx10042);
   ix19302 : nor02_2x port map ( Y=>nx18921, A0=>nx10120, A1=>nx10082);
   ix19303 : and03 port map ( Y=>nx18922, A0=>nx18921, A1=>nx14846, A2=>
      nx15008);
   ix19304 : nand03_2x port map ( Y=>nx18923, A0=>nx18918, A1=>nx18920, A2=>
      nx18922);
   reg_nx14825 : nor04_2x port map ( Y=>nx14825, A0=>nx9826, A1=>nx18912, A2
      =>nx18917, A3=>nx18923);
   reg_nx10545 : nor02ii port map ( Y=>nx10545, A0=>address(5), A1=>
      address(4));
   ix19305 : inv01 port map ( Y=>nx18924, A=>address(5));
   reg_nx17301 : nand02_2x port map ( Y=>nx17301, A0=>address(4), A1=>
      nx18924);
   reg_nx10523 : inv01 port map ( Y=>nx10523, A=>address(4));
   reg_nx10511 : nor02_2x port map ( Y=>nx10511, A0=>address(0), A1=>
      address(1));
   reg_nx16283 : nor02ii port map ( Y=>nx16283, A0=>address(4), A1=>
      address(5));
   reg_nx10949 : nand04_2x port map ( Y=>nx10949, A0=>nx18956, A1=>nx19343, 
      A2=>address(2), A3=>address(3));
   reg_nx10525 : inv01 port map ( Y=>nx10525, A=>address(5));
   reg_nx17177 : inv01 port map ( Y=>nx17177, A=>nx18956);
   reg_nx16151 : inv01 port map ( Y=>nx16151, A=>nx18956);
   ix19306 : inv01 port map ( Y=>nx18925, A=>nx18956);
   ix19307 : inv01 port map ( Y=>nx18926, A=>nx18956);
   ix19308 : inv01 port map ( Y=>nx18927, A=>nx18956);
   ix19309 : inv01 port map ( Y=>nx18928, A=>nx10557);
   ix19310 : inv01 port map ( Y=>nx18929, A=>nx16191);
   reg_nx2622 : oai32 port map ( Y=>nx2622, A0=>nx18928, A1=>nx18929, A2=>
      nx11408, B0=>nx18958, B1=>nx11411);
   ix19311 : oai322 port map ( Y=>nx18930, A0=>nx15889, A1=>nx11583, A2=>
      nx15763, B0=>nx16495, B1=>nx11530, C0=>nx16479, C1=>nx11527);
   reg_nx2226 : oai22 port map ( Y=>nx2226, A0=>nx16603, A1=>nx11587, B0=>
      nx11590, B1=>nx16619);
   ix19312 : oai322 port map ( Y=>nx18931, A0=>nx15929, A1=>nx11579, A2=>
      nx15421, B0=>nx16455, B1=>nx11513, C0=>nx16439, C1=>nx11510);
   ix19313 : nor04_2x port map ( Y=>nx18932, A0=>nx2622, A1=>nx18930, A2=>
      nx2226, A3=>nx18931);
   ix19314 : nand02_2x port map ( Y=>nx18933, A0=>nx17147, A1=>nx10567);
   ix19315 : inv01 port map ( Y=>nx18934, A=>address(2));
   ix19316 : inv02 port map ( Y=>nx18935, A=>address(3));
   ix19317 : inv01 port map ( Y=>nx18936, A=>nx10557);
   ix19318 : inv01 port map ( Y=>nx18937, A=>nx16191);
   reg_nx1984 : oai43 port map ( Y=>nx1984, A0=>nx18933, A1=>nx11125, A2=>
      nx18934, A3=>nx18935, B0=>nx18936, B1=>nx18937, B2=>nx11122);
   ix19319 : oai322 port map ( Y=>nx18938, A0=>nx15889, A1=>nx11297, A2=>
      nx15761, B0=>nx16495, B1=>nx11244, C0=>nx16479, C1=>nx11241);
   reg_nx1588 : oai22 port map ( Y=>nx1588, A0=>nx16603, A1=>nx11301, B0=>
      nx11304, B1=>nx16619);
   ix19320 : oai322 port map ( Y=>nx18939, A0=>nx15929, A1=>nx11293, A2=>
      nx15419, B0=>nx16455, B1=>nx11227, C0=>nx16439, C1=>nx11224);
   ix19321 : nor04_2x port map ( Y=>nx18940, A0=>nx1984, A1=>nx18938, A2=>
      nx1588, A3=>nx18939);
   ix19322 : nand02_2x port map ( Y=>nx18941, A0=>nx17147, A1=>nx10567);
   ix19323 : inv01 port map ( Y=>nx18942, A=>address(2));
   ix19324 : inv02 port map ( Y=>nx18943, A=>address(3));
   ix19325 : inv01 port map ( Y=>nx18944, A=>nx10557);
   ix19326 : inv01 port map ( Y=>nx18945, A=>nx16191);
   reg_nx1326 : oai43 port map ( Y=>nx1326, A0=>nx18941, A1=>nx10559, A2=>
      nx18942, A3=>nx18943, B0=>nx18944, B1=>nx18945, B2=>nx10548);
   reg_nx16495 : inv02 port map ( Y=>nx16495, A=>nx16493);
   reg_nx16479 : inv02 port map ( Y=>nx16479, A=>nx16477);
   ix19327 : oai322 port map ( Y=>nx18946, A0=>nx15889, A1=>nx10928, A2=>
      nx15759, B0=>nx16495, B1=>nx10825, C0=>nx16479, C1=>nx10817);
   reg_nx16603 : inv02 port map ( Y=>nx16603, A=>nx16601);
   reg_nx514 : oai22 port map ( Y=>nx514, A0=>nx16603, A1=>nx10935, B0=>
      nx10943, B1=>nx16619);
   reg_nx16455 : inv02 port map ( Y=>nx16455, A=>nx16453);
   reg_nx16439 : inv02 port map ( Y=>nx16439, A=>nx16437);
   ix19328 : oai322 port map ( Y=>nx18947, A0=>nx15929, A1=>nx10922, A2=>
      nx17141, B0=>nx16455, B1=>nx10789, C0=>nx16439, C1=>nx10783);
   ix19329 : nor04_2x port map ( Y=>nx18948, A0=>nx1326, A1=>nx18946, A2=>
      nx514, A3=>nx18947);
   reg_nx16201 : nand02_2x port map ( Y=>nx16201, A0=>nx16191, A1=>nx10557);
   reg_nx10565 : nand04_2x port map ( Y=>nx10565, A0=>address(2), A1=>
      address(3), A2=>nx17147, A3=>nx10567);
   ix19330 : inv01 port map ( Y=>nx18949, A=>nx10557);
   ix19331 : inv01 port map ( Y=>nx18950, A=>nx16191);
   reg_nx9640 : oai32 port map ( Y=>nx9640, A0=>nx18949, A1=>nx18950, A2=>
      nx14554, B0=>nx18958, B1=>nx14557);
   reg_nx16497 : inv02 port map ( Y=>nx16497, A=>nx16493);
   reg_nx16481 : inv02 port map ( Y=>nx16481, A=>nx16477);
   ix19332 : oai322 port map ( Y=>nx18951, A0=>nx15893, A1=>nx14729, A2=>
      nx15785, B0=>nx16497, B1=>nx14676, C0=>nx16481, C1=>nx14673);
   reg_nx16605 : inv02 port map ( Y=>nx16605, A=>nx16601);
   reg_nx9244 : oai22 port map ( Y=>nx9244, A0=>nx16605, A1=>nx14733, B0=>
      nx14736, B1=>nx16621);
   reg_nx16457 : inv02 port map ( Y=>nx16457, A=>nx16453);
   reg_nx16441 : inv02 port map ( Y=>nx16441, A=>nx16437);
   ix19333 : oai322 port map ( Y=>nx18952, A0=>nx15933, A1=>nx14725, A2=>
      nx15445, B0=>nx16457, B1=>nx14659, C0=>nx16441, C1=>nx14656);
   ix19334 : nor04_2x port map ( Y=>nx18953, A0=>nx9640, A1=>nx18951, A2=>
      nx9244, A3=>nx18952);
   reg_nx16203 : nand02_2x port map ( Y=>nx16203, A0=>nx16191, A1=>nx10557);
   ix19335 : oai22 port map ( Y=>nx18954, A0=>nx12748, A1=>nx16643, B0=>
      nx12751, B1=>nx16659);
   reg_nx12737 : nor03_2x port map ( Y=>nx12737, A0=>nx18954, A1=>nx4756, A2
      =>nx4748);
   ix19336 : buf16 port map ( Y=>nx18955, A=>nx10511);
   ix19337 : buf16 port map ( Y=>nx18956, A=>nx10511);
   ix19338 : buf16 port map ( Y=>nx18957, A=>nx10565);
   ix19339 : buf16 port map ( Y=>nx18958, A=>nx10565);
   ix19340 : inv02 port map ( Y=>nx19341, A=>nx17303);
   ix19342 : inv02 port map ( Y=>nx19343, A=>nx17169);
end Behavioral ;

