
-- 
-- Definition of  DCNNChip
-- 
--      Sun May 12 02:11:27 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Queue_5 is
   port (
      d : IN std_logic_vector (15 DOWNTO 0) ;
      q_0_15 : OUT std_logic ;
      q_0_14 : OUT std_logic ;
      q_0_13 : OUT std_logic ;
      q_0_12 : OUT std_logic ;
      q_0_11 : OUT std_logic ;
      q_0_10 : OUT std_logic ;
      q_0_9 : OUT std_logic ;
      q_0_8 : OUT std_logic ;
      q_0_7 : OUT std_logic ;
      q_0_6 : OUT std_logic ;
      q_0_5 : OUT std_logic ;
      q_0_4 : OUT std_logic ;
      q_0_3 : OUT std_logic ;
      q_0_2 : OUT std_logic ;
      q_0_1 : OUT std_logic ;
      q_0_0 : OUT std_logic ;
      q_1_15 : OUT std_logic ;
      q_1_14 : OUT std_logic ;
      q_1_13 : OUT std_logic ;
      q_1_12 : OUT std_logic ;
      q_1_11 : OUT std_logic ;
      q_1_10 : OUT std_logic ;
      q_1_9 : OUT std_logic ;
      q_1_8 : OUT std_logic ;
      q_1_7 : OUT std_logic ;
      q_1_6 : OUT std_logic ;
      q_1_5 : OUT std_logic ;
      q_1_4 : OUT std_logic ;
      q_1_3 : OUT std_logic ;
      q_1_2 : OUT std_logic ;
      q_1_1 : OUT std_logic ;
      q_1_0 : OUT std_logic ;
      q_2_15 : OUT std_logic ;
      q_2_14 : OUT std_logic ;
      q_2_13 : OUT std_logic ;
      q_2_12 : OUT std_logic ;
      q_2_11 : OUT std_logic ;
      q_2_10 : OUT std_logic ;
      q_2_9 : OUT std_logic ;
      q_2_8 : OUT std_logic ;
      q_2_7 : OUT std_logic ;
      q_2_6 : OUT std_logic ;
      q_2_5 : OUT std_logic ;
      q_2_4 : OUT std_logic ;
      q_2_3 : OUT std_logic ;
      q_2_2 : OUT std_logic ;
      q_2_1 : OUT std_logic ;
      q_2_0 : OUT std_logic ;
      q_3_15 : OUT std_logic ;
      q_3_14 : OUT std_logic ;
      q_3_13 : OUT std_logic ;
      q_3_12 : OUT std_logic ;
      q_3_11 : OUT std_logic ;
      q_3_10 : OUT std_logic ;
      q_3_9 : OUT std_logic ;
      q_3_8 : OUT std_logic ;
      q_3_7 : OUT std_logic ;
      q_3_6 : OUT std_logic ;
      q_3_5 : OUT std_logic ;
      q_3_4 : OUT std_logic ;
      q_3_3 : OUT std_logic ;
      q_3_2 : OUT std_logic ;
      q_3_1 : OUT std_logic ;
      q_3_0 : OUT std_logic ;
      q_4_15 : OUT std_logic ;
      q_4_14 : OUT std_logic ;
      q_4_13 : OUT std_logic ;
      q_4_12 : OUT std_logic ;
      q_4_11 : OUT std_logic ;
      q_4_10 : OUT std_logic ;
      q_4_9 : OUT std_logic ;
      q_4_8 : OUT std_logic ;
      q_4_7 : OUT std_logic ;
      q_4_6 : OUT std_logic ;
      q_4_5 : OUT std_logic ;
      q_4_4 : OUT std_logic ;
      q_4_3 : OUT std_logic ;
      q_4_2 : OUT std_logic ;
      q_4_1 : OUT std_logic ;
      q_4_0 : OUT std_logic ;
      clk : IN std_logic ;
      load : IN std_logic ;
      reset : IN std_logic) ;
end Queue_5 ;

architecture Dataflow of Queue_5 is
   signal q_0_15_EXMPLR, q_0_14_EXMPLR, q_0_13_EXMPLR, q_0_12_EXMPLR, 
      q_0_11_EXMPLR, q_0_10_EXMPLR, q_0_9_EXMPLR, q_0_8_EXMPLR, q_0_7_EXMPLR, 
      q_0_6_EXMPLR, q_0_5_EXMPLR, q_0_4_EXMPLR, q_0_3_EXMPLR, q_0_2_EXMPLR, 
      q_0_1_EXMPLR, q_0_0_EXMPLR, q_1_15_EXMPLR, q_1_14_EXMPLR, 
      q_1_13_EXMPLR, q_1_12_EXMPLR, q_1_11_EXMPLR, q_1_10_EXMPLR, 
      q_1_9_EXMPLR, q_1_8_EXMPLR, q_1_7_EXMPLR, q_1_6_EXMPLR, q_1_5_EXMPLR, 
      q_1_4_EXMPLR, q_1_3_EXMPLR, q_1_2_EXMPLR, q_1_1_EXMPLR, q_1_0_EXMPLR, 
      q_2_15_EXMPLR, q_2_14_EXMPLR, q_2_13_EXMPLR, q_2_12_EXMPLR, 
      q_2_11_EXMPLR, q_2_10_EXMPLR, q_2_9_EXMPLR, q_2_8_EXMPLR, q_2_7_EXMPLR, 
      q_2_6_EXMPLR, q_2_5_EXMPLR, q_2_4_EXMPLR, q_2_3_EXMPLR, q_2_2_EXMPLR, 
      q_2_1_EXMPLR, q_2_0_EXMPLR, q_3_15_EXMPLR, q_3_14_EXMPLR, 
      q_3_13_EXMPLR, q_3_12_EXMPLR, q_3_11_EXMPLR, q_3_10_EXMPLR, 
      q_3_9_EXMPLR, q_3_8_EXMPLR, q_3_7_EXMPLR, q_3_6_EXMPLR, q_3_5_EXMPLR, 
      q_3_4_EXMPLR, q_3_3_EXMPLR, q_3_2_EXMPLR, q_3_1_EXMPLR, q_3_0_EXMPLR, 
      q_4_15_EXMPLR, q_4_14_EXMPLR, q_4_13_EXMPLR, q_4_12_EXMPLR, 
      q_4_11_EXMPLR, q_4_10_EXMPLR, q_4_9_EXMPLR, q_4_8_EXMPLR, q_4_7_EXMPLR, 
      q_4_6_EXMPLR, q_4_5_EXMPLR, q_4_4_EXMPLR, q_4_3_EXMPLR, q_4_2_EXMPLR, 
      q_4_1_EXMPLR, q_4_0_EXMPLR, nx393, nx403, nx413, nx423, nx433, nx443, 
      nx453, nx463, nx473, nx483, nx493, nx503, nx513, nx523, nx533, nx543, 
      nx553, nx563, nx573, nx583, nx593, nx603, nx613, nx623, nx633, nx643, 
      nx653, nx663, nx673, nx683, nx693, nx703, nx713, nx723, nx733, nx743, 
      nx753, nx763, nx773, nx783, nx793, nx803, nx813, nx823, nx833, nx843, 
      nx853, nx863, nx873, nx883, nx893, nx903, nx913, nx923, nx933, nx943, 
      nx953, nx963, nx973, nx983, nx993, nx1003, nx1013, nx1023, nx1033, 
      nx1043, nx1053, nx1063, nx1073, nx1083, nx1093, nx1103, nx1113, nx1123, 
      nx1133, nx1143, nx1153, nx1163, nx1173, nx1183, nx1440, nx1442, nx1444, 
      nx1446, nx1448, nx1450, nx1452, nx1454, nx1456, nx1458, nx1460, nx1462, 
      nx1466, nx1468, nx1470, nx1472, nx1474, nx1476, nx1478, nx1480, nx1482, 
      nx1484, nx1486, nx1488, nx1492, nx1494, nx1496, nx1498, nx1500, nx1502, 
      nx1504, nx1506, nx1508, nx1510, nx1512, nx1514, nx1516, nx1518, nx1520, 
      nx1522, nx1524, nx1526: std_logic ;

begin
   q_0_15 <= q_0_15_EXMPLR ;
   q_0_14 <= q_0_14_EXMPLR ;
   q_0_13 <= q_0_13_EXMPLR ;
   q_0_12 <= q_0_12_EXMPLR ;
   q_0_11 <= q_0_11_EXMPLR ;
   q_0_10 <= q_0_10_EXMPLR ;
   q_0_9 <= q_0_9_EXMPLR ;
   q_0_8 <= q_0_8_EXMPLR ;
   q_0_7 <= q_0_7_EXMPLR ;
   q_0_6 <= q_0_6_EXMPLR ;
   q_0_5 <= q_0_5_EXMPLR ;
   q_0_4 <= q_0_4_EXMPLR ;
   q_0_3 <= q_0_3_EXMPLR ;
   q_0_2 <= q_0_2_EXMPLR ;
   q_0_1 <= q_0_1_EXMPLR ;
   q_0_0 <= q_0_0_EXMPLR ;
   q_1_15 <= q_1_15_EXMPLR ;
   q_1_14 <= q_1_14_EXMPLR ;
   q_1_13 <= q_1_13_EXMPLR ;
   q_1_12 <= q_1_12_EXMPLR ;
   q_1_11 <= q_1_11_EXMPLR ;
   q_1_10 <= q_1_10_EXMPLR ;
   q_1_9 <= q_1_9_EXMPLR ;
   q_1_8 <= q_1_8_EXMPLR ;
   q_1_7 <= q_1_7_EXMPLR ;
   q_1_6 <= q_1_6_EXMPLR ;
   q_1_5 <= q_1_5_EXMPLR ;
   q_1_4 <= q_1_4_EXMPLR ;
   q_1_3 <= q_1_3_EXMPLR ;
   q_1_2 <= q_1_2_EXMPLR ;
   q_1_1 <= q_1_1_EXMPLR ;
   q_1_0 <= q_1_0_EXMPLR ;
   q_2_15 <= q_2_15_EXMPLR ;
   q_2_14 <= q_2_14_EXMPLR ;
   q_2_13 <= q_2_13_EXMPLR ;
   q_2_12 <= q_2_12_EXMPLR ;
   q_2_11 <= q_2_11_EXMPLR ;
   q_2_10 <= q_2_10_EXMPLR ;
   q_2_9 <= q_2_9_EXMPLR ;
   q_2_8 <= q_2_8_EXMPLR ;
   q_2_7 <= q_2_7_EXMPLR ;
   q_2_6 <= q_2_6_EXMPLR ;
   q_2_5 <= q_2_5_EXMPLR ;
   q_2_4 <= q_2_4_EXMPLR ;
   q_2_3 <= q_2_3_EXMPLR ;
   q_2_2 <= q_2_2_EXMPLR ;
   q_2_1 <= q_2_1_EXMPLR ;
   q_2_0 <= q_2_0_EXMPLR ;
   q_3_15 <= q_3_15_EXMPLR ;
   q_3_14 <= q_3_14_EXMPLR ;
   q_3_13 <= q_3_13_EXMPLR ;
   q_3_12 <= q_3_12_EXMPLR ;
   q_3_11 <= q_3_11_EXMPLR ;
   q_3_10 <= q_3_10_EXMPLR ;
   q_3_9 <= q_3_9_EXMPLR ;
   q_3_8 <= q_3_8_EXMPLR ;
   q_3_7 <= q_3_7_EXMPLR ;
   q_3_6 <= q_3_6_EXMPLR ;
   q_3_5 <= q_3_5_EXMPLR ;
   q_3_4 <= q_3_4_EXMPLR ;
   q_3_3 <= q_3_3_EXMPLR ;
   q_3_2 <= q_3_2_EXMPLR ;
   q_3_1 <= q_3_1_EXMPLR ;
   q_3_0 <= q_3_0_EXMPLR ;
   q_4_15 <= q_4_15_EXMPLR ;
   q_4_14 <= q_4_14_EXMPLR ;
   q_4_13 <= q_4_13_EXMPLR ;
   q_4_12 <= q_4_12_EXMPLR ;
   q_4_11 <= q_4_11_EXMPLR ;
   q_4_10 <= q_4_10_EXMPLR ;
   q_4_9 <= q_4_9_EXMPLR ;
   q_4_8 <= q_4_8_EXMPLR ;
   q_4_7 <= q_4_7_EXMPLR ;
   q_4_6 <= q_4_6_EXMPLR ;
   q_4_5 <= q_4_5_EXMPLR ;
   q_4_4 <= q_4_4_EXMPLR ;
   q_4_3 <= q_4_3_EXMPLR ;
   q_4_2 <= q_4_2_EXMPLR ;
   q_4_1 <= q_4_1_EXMPLR ;
   q_4_0 <= q_4_0_EXMPLR ;
   gen_regs_4_regi_reg_q_0 : dffr port map ( Q=>q_4_0_EXMPLR, QB=>OPEN, D=>
      nx433, CLK=>nx1492, R=>nx1466);
   ix434 : mux21_ni port map ( Y=>nx433, A0=>q_4_0_EXMPLR, A1=>q_3_0_EXMPLR, 
      S0=>nx1440);
   gen_regs_3_regi_reg_q_0 : dffr port map ( Q=>q_3_0_EXMPLR, QB=>OPEN, D=>
      nx423, CLK=>nx1492, R=>nx1466);
   ix424 : mux21_ni port map ( Y=>nx423, A0=>q_3_0_EXMPLR, A1=>q_2_0_EXMPLR, 
      S0=>nx1440);
   gen_regs_2_regi_reg_q_0 : dffr port map ( Q=>q_2_0_EXMPLR, QB=>OPEN, D=>
      nx413, CLK=>nx1492, R=>nx1466);
   ix414 : mux21_ni port map ( Y=>nx413, A0=>q_2_0_EXMPLR, A1=>q_1_0_EXMPLR, 
      S0=>nx1440);
   gen_regs_1_regi_reg_q_0 : dffr port map ( Q=>q_1_0_EXMPLR, QB=>OPEN, D=>
      nx403, CLK=>nx1492, R=>nx1466);
   ix404 : mux21_ni port map ( Y=>nx403, A0=>q_1_0_EXMPLR, A1=>q_0_0_EXMPLR, 
      S0=>nx1440);
   reg0_reg_q_0 : dffr port map ( Q=>q_0_0_EXMPLR, QB=>OPEN, D=>nx393, CLK=>
      nx1492, R=>nx1466);
   ix394 : mux21_ni port map ( Y=>nx393, A0=>q_0_0_EXMPLR, A1=>d(0), S0=>
      nx1440);
   gen_regs_4_regi_reg_q_1 : dffr port map ( Q=>q_4_1_EXMPLR, QB=>OPEN, D=>
      nx483, CLK=>nx1494, R=>nx1468);
   ix484 : mux21_ni port map ( Y=>nx483, A0=>q_4_1_EXMPLR, A1=>q_3_1_EXMPLR, 
      S0=>nx1442);
   gen_regs_3_regi_reg_q_1 : dffr port map ( Q=>q_3_1_EXMPLR, QB=>OPEN, D=>
      nx473, CLK=>nx1494, R=>nx1468);
   ix474 : mux21_ni port map ( Y=>nx473, A0=>q_3_1_EXMPLR, A1=>q_2_1_EXMPLR, 
      S0=>nx1442);
   gen_regs_2_regi_reg_q_1 : dffr port map ( Q=>q_2_1_EXMPLR, QB=>OPEN, D=>
      nx463, CLK=>nx1494, R=>nx1468);
   ix464 : mux21_ni port map ( Y=>nx463, A0=>q_2_1_EXMPLR, A1=>q_1_1_EXMPLR, 
      S0=>nx1442);
   gen_regs_1_regi_reg_q_1 : dffr port map ( Q=>q_1_1_EXMPLR, QB=>OPEN, D=>
      nx453, CLK=>nx1492, R=>nx1466);
   ix454 : mux21_ni port map ( Y=>nx453, A0=>q_1_1_EXMPLR, A1=>q_0_1_EXMPLR, 
      S0=>nx1440);
   reg0_reg_q_1 : dffr port map ( Q=>q_0_1_EXMPLR, QB=>OPEN, D=>nx443, CLK=>
      nx1492, R=>nx1466);
   ix444 : mux21_ni port map ( Y=>nx443, A0=>q_0_1_EXMPLR, A1=>d(1), S0=>
      nx1440);
   gen_regs_4_regi_reg_q_2 : dffr port map ( Q=>q_4_2_EXMPLR, QB=>OPEN, D=>
      nx533, CLK=>nx1496, R=>nx1470);
   ix534 : mux21_ni port map ( Y=>nx533, A0=>q_4_2_EXMPLR, A1=>q_3_2_EXMPLR, 
      S0=>nx1444);
   gen_regs_3_regi_reg_q_2 : dffr port map ( Q=>q_3_2_EXMPLR, QB=>OPEN, D=>
      nx523, CLK=>nx1494, R=>nx1468);
   ix524 : mux21_ni port map ( Y=>nx523, A0=>q_3_2_EXMPLR, A1=>q_2_2_EXMPLR, 
      S0=>nx1442);
   gen_regs_2_regi_reg_q_2 : dffr port map ( Q=>q_2_2_EXMPLR, QB=>OPEN, D=>
      nx513, CLK=>nx1494, R=>nx1468);
   ix514 : mux21_ni port map ( Y=>nx513, A0=>q_2_2_EXMPLR, A1=>q_1_2_EXMPLR, 
      S0=>nx1442);
   gen_regs_1_regi_reg_q_2 : dffr port map ( Q=>q_1_2_EXMPLR, QB=>OPEN, D=>
      nx503, CLK=>nx1494, R=>nx1468);
   ix504 : mux21_ni port map ( Y=>nx503, A0=>q_1_2_EXMPLR, A1=>q_0_2_EXMPLR, 
      S0=>nx1442);
   reg0_reg_q_2 : dffr port map ( Q=>q_0_2_EXMPLR, QB=>OPEN, D=>nx493, CLK=>
      nx1494, R=>nx1468);
   ix494 : mux21_ni port map ( Y=>nx493, A0=>q_0_2_EXMPLR, A1=>d(2), S0=>
      nx1442);
   gen_regs_4_regi_reg_q_3 : dffr port map ( Q=>q_4_3_EXMPLR, QB=>OPEN, D=>
      nx583, CLK=>nx1496, R=>nx1470);
   ix584 : mux21_ni port map ( Y=>nx583, A0=>q_4_3_EXMPLR, A1=>q_3_3_EXMPLR, 
      S0=>nx1444);
   gen_regs_3_regi_reg_q_3 : dffr port map ( Q=>q_3_3_EXMPLR, QB=>OPEN, D=>
      nx573, CLK=>nx1496, R=>nx1470);
   ix574 : mux21_ni port map ( Y=>nx573, A0=>q_3_3_EXMPLR, A1=>q_2_3_EXMPLR, 
      S0=>nx1444);
   gen_regs_2_regi_reg_q_3 : dffr port map ( Q=>q_2_3_EXMPLR, QB=>OPEN, D=>
      nx563, CLK=>nx1496, R=>nx1470);
   ix564 : mux21_ni port map ( Y=>nx563, A0=>q_2_3_EXMPLR, A1=>q_1_3_EXMPLR, 
      S0=>nx1444);
   gen_regs_1_regi_reg_q_3 : dffr port map ( Q=>q_1_3_EXMPLR, QB=>OPEN, D=>
      nx553, CLK=>nx1496, R=>nx1470);
   ix554 : mux21_ni port map ( Y=>nx553, A0=>q_1_3_EXMPLR, A1=>q_0_3_EXMPLR, 
      S0=>nx1444);
   reg0_reg_q_3 : dffr port map ( Q=>q_0_3_EXMPLR, QB=>OPEN, D=>nx543, CLK=>
      nx1496, R=>nx1470);
   ix544 : mux21_ni port map ( Y=>nx543, A0=>q_0_3_EXMPLR, A1=>d(3), S0=>
      nx1444);
   gen_regs_4_regi_reg_q_4 : dffr port map ( Q=>q_4_4_EXMPLR, QB=>OPEN, D=>
      nx633, CLK=>nx1498, R=>nx1472);
   ix634 : mux21_ni port map ( Y=>nx633, A0=>q_4_4_EXMPLR, A1=>q_3_4_EXMPLR, 
      S0=>nx1446);
   gen_regs_3_regi_reg_q_4 : dffr port map ( Q=>q_3_4_EXMPLR, QB=>OPEN, D=>
      nx623, CLK=>nx1498, R=>nx1472);
   ix624 : mux21_ni port map ( Y=>nx623, A0=>q_3_4_EXMPLR, A1=>q_2_4_EXMPLR, 
      S0=>nx1446);
   gen_regs_2_regi_reg_q_4 : dffr port map ( Q=>q_2_4_EXMPLR, QB=>OPEN, D=>
      nx613, CLK=>nx1498, R=>nx1472);
   ix614 : mux21_ni port map ( Y=>nx613, A0=>q_2_4_EXMPLR, A1=>q_1_4_EXMPLR, 
      S0=>nx1446);
   gen_regs_1_regi_reg_q_4 : dffr port map ( Q=>q_1_4_EXMPLR, QB=>OPEN, D=>
      nx603, CLK=>nx1498, R=>nx1472);
   ix604 : mux21_ni port map ( Y=>nx603, A0=>q_1_4_EXMPLR, A1=>q_0_4_EXMPLR, 
      S0=>nx1446);
   reg0_reg_q_4 : dffr port map ( Q=>q_0_4_EXMPLR, QB=>OPEN, D=>nx593, CLK=>
      nx1496, R=>nx1470);
   ix594 : mux21_ni port map ( Y=>nx593, A0=>q_0_4_EXMPLR, A1=>d(4), S0=>
      nx1444);
   gen_regs_4_regi_reg_q_5 : dffr port map ( Q=>q_4_5_EXMPLR, QB=>OPEN, D=>
      nx683, CLK=>nx1500, R=>nx1474);
   ix684 : mux21_ni port map ( Y=>nx683, A0=>q_4_5_EXMPLR, A1=>q_3_5_EXMPLR, 
      S0=>nx1448);
   gen_regs_3_regi_reg_q_5 : dffr port map ( Q=>q_3_5_EXMPLR, QB=>OPEN, D=>
      nx673, CLK=>nx1500, R=>nx1474);
   ix674 : mux21_ni port map ( Y=>nx673, A0=>q_3_5_EXMPLR, A1=>q_2_5_EXMPLR, 
      S0=>nx1448);
   gen_regs_2_regi_reg_q_5 : dffr port map ( Q=>q_2_5_EXMPLR, QB=>OPEN, D=>
      nx663, CLK=>nx1498, R=>nx1472);
   ix664 : mux21_ni port map ( Y=>nx663, A0=>q_2_5_EXMPLR, A1=>q_1_5_EXMPLR, 
      S0=>nx1446);
   gen_regs_1_regi_reg_q_5 : dffr port map ( Q=>q_1_5_EXMPLR, QB=>OPEN, D=>
      nx653, CLK=>nx1498, R=>nx1472);
   ix654 : mux21_ni port map ( Y=>nx653, A0=>q_1_5_EXMPLR, A1=>q_0_5_EXMPLR, 
      S0=>nx1446);
   reg0_reg_q_5 : dffr port map ( Q=>q_0_5_EXMPLR, QB=>OPEN, D=>nx643, CLK=>
      nx1498, R=>nx1472);
   ix644 : mux21_ni port map ( Y=>nx643, A0=>q_0_5_EXMPLR, A1=>d(5), S0=>
      nx1446);
   gen_regs_4_regi_reg_q_6 : dffr port map ( Q=>q_4_6_EXMPLR, QB=>OPEN, D=>
      nx733, CLK=>nx1500, R=>nx1474);
   ix734 : mux21_ni port map ( Y=>nx733, A0=>q_4_6_EXMPLR, A1=>q_3_6_EXMPLR, 
      S0=>nx1448);
   gen_regs_3_regi_reg_q_6 : dffr port map ( Q=>q_3_6_EXMPLR, QB=>OPEN, D=>
      nx723, CLK=>nx1500, R=>nx1474);
   ix724 : mux21_ni port map ( Y=>nx723, A0=>q_3_6_EXMPLR, A1=>q_2_6_EXMPLR, 
      S0=>nx1448);
   gen_regs_2_regi_reg_q_6 : dffr port map ( Q=>q_2_6_EXMPLR, QB=>OPEN, D=>
      nx713, CLK=>nx1500, R=>nx1474);
   ix714 : mux21_ni port map ( Y=>nx713, A0=>q_2_6_EXMPLR, A1=>q_1_6_EXMPLR, 
      S0=>nx1448);
   gen_regs_1_regi_reg_q_6 : dffr port map ( Q=>q_1_6_EXMPLR, QB=>OPEN, D=>
      nx703, CLK=>nx1500, R=>nx1474);
   ix704 : mux21_ni port map ( Y=>nx703, A0=>q_1_6_EXMPLR, A1=>q_0_6_EXMPLR, 
      S0=>nx1448);
   reg0_reg_q_6 : dffr port map ( Q=>q_0_6_EXMPLR, QB=>OPEN, D=>nx693, CLK=>
      nx1500, R=>nx1474);
   ix694 : mux21_ni port map ( Y=>nx693, A0=>q_0_6_EXMPLR, A1=>d(6), S0=>
      nx1448);
   gen_regs_4_regi_reg_q_7 : dffr port map ( Q=>q_4_7_EXMPLR, QB=>OPEN, D=>
      nx783, CLK=>nx1502, R=>nx1476);
   ix784 : mux21_ni port map ( Y=>nx783, A0=>q_4_7_EXMPLR, A1=>q_3_7_EXMPLR, 
      S0=>nx1450);
   gen_regs_3_regi_reg_q_7 : dffr port map ( Q=>q_3_7_EXMPLR, QB=>OPEN, D=>
      nx773, CLK=>nx1502, R=>nx1476);
   ix774 : mux21_ni port map ( Y=>nx773, A0=>q_3_7_EXMPLR, A1=>q_2_7_EXMPLR, 
      S0=>nx1450);
   gen_regs_2_regi_reg_q_7 : dffr port map ( Q=>q_2_7_EXMPLR, QB=>OPEN, D=>
      nx763, CLK=>nx1502, R=>nx1476);
   ix764 : mux21_ni port map ( Y=>nx763, A0=>q_2_7_EXMPLR, A1=>q_1_7_EXMPLR, 
      S0=>nx1450);
   gen_regs_1_regi_reg_q_7 : dffr port map ( Q=>q_1_7_EXMPLR, QB=>OPEN, D=>
      nx753, CLK=>nx1502, R=>nx1476);
   ix754 : mux21_ni port map ( Y=>nx753, A0=>q_1_7_EXMPLR, A1=>q_0_7_EXMPLR, 
      S0=>nx1450);
   reg0_reg_q_7 : dffr port map ( Q=>q_0_7_EXMPLR, QB=>OPEN, D=>nx743, CLK=>
      nx1502, R=>nx1476);
   ix744 : mux21_ni port map ( Y=>nx743, A0=>q_0_7_EXMPLR, A1=>d(7), S0=>
      nx1450);
   gen_regs_4_regi_reg_q_8 : dffr port map ( Q=>q_4_8_EXMPLR, QB=>OPEN, D=>
      nx833, CLK=>nx1504, R=>nx1478);
   ix834 : mux21_ni port map ( Y=>nx833, A0=>q_4_8_EXMPLR, A1=>q_3_8_EXMPLR, 
      S0=>nx1452);
   gen_regs_3_regi_reg_q_8 : dffr port map ( Q=>q_3_8_EXMPLR, QB=>OPEN, D=>
      nx823, CLK=>nx1504, R=>nx1478);
   ix824 : mux21_ni port map ( Y=>nx823, A0=>q_3_8_EXMPLR, A1=>q_2_8_EXMPLR, 
      S0=>nx1452);
   gen_regs_2_regi_reg_q_8 : dffr port map ( Q=>q_2_8_EXMPLR, QB=>OPEN, D=>
      nx813, CLK=>nx1504, R=>nx1478);
   ix814 : mux21_ni port map ( Y=>nx813, A0=>q_2_8_EXMPLR, A1=>q_1_8_EXMPLR, 
      S0=>nx1452);
   gen_regs_1_regi_reg_q_8 : dffr port map ( Q=>q_1_8_EXMPLR, QB=>OPEN, D=>
      nx803, CLK=>nx1502, R=>nx1476);
   ix804 : mux21_ni port map ( Y=>nx803, A0=>q_1_8_EXMPLR, A1=>q_0_8_EXMPLR, 
      S0=>nx1450);
   reg0_reg_q_8 : dffr port map ( Q=>q_0_8_EXMPLR, QB=>OPEN, D=>nx793, CLK=>
      nx1502, R=>nx1476);
   ix794 : mux21_ni port map ( Y=>nx793, A0=>q_0_8_EXMPLR, A1=>d(8), S0=>
      nx1450);
   gen_regs_4_regi_reg_q_9 : dffr port map ( Q=>q_4_9_EXMPLR, QB=>OPEN, D=>
      nx883, CLK=>nx1506, R=>nx1480);
   ix884 : mux21_ni port map ( Y=>nx883, A0=>q_4_9_EXMPLR, A1=>q_3_9_EXMPLR, 
      S0=>nx1454);
   gen_regs_3_regi_reg_q_9 : dffr port map ( Q=>q_3_9_EXMPLR, QB=>OPEN, D=>
      nx873, CLK=>nx1504, R=>nx1478);
   ix874 : mux21_ni port map ( Y=>nx873, A0=>q_3_9_EXMPLR, A1=>q_2_9_EXMPLR, 
      S0=>nx1452);
   gen_regs_2_regi_reg_q_9 : dffr port map ( Q=>q_2_9_EXMPLR, QB=>OPEN, D=>
      nx863, CLK=>nx1504, R=>nx1478);
   ix864 : mux21_ni port map ( Y=>nx863, A0=>q_2_9_EXMPLR, A1=>q_1_9_EXMPLR, 
      S0=>nx1452);
   gen_regs_1_regi_reg_q_9 : dffr port map ( Q=>q_1_9_EXMPLR, QB=>OPEN, D=>
      nx853, CLK=>nx1504, R=>nx1478);
   ix854 : mux21_ni port map ( Y=>nx853, A0=>q_1_9_EXMPLR, A1=>q_0_9_EXMPLR, 
      S0=>nx1452);
   reg0_reg_q_9 : dffr port map ( Q=>q_0_9_EXMPLR, QB=>OPEN, D=>nx843, CLK=>
      nx1504, R=>nx1478);
   ix844 : mux21_ni port map ( Y=>nx843, A0=>q_0_9_EXMPLR, A1=>d(9), S0=>
      nx1452);
   gen_regs_4_regi_reg_q_10 : dffr port map ( Q=>q_4_10_EXMPLR, QB=>OPEN, D
      =>nx933, CLK=>nx1506, R=>nx1480);
   ix934 : mux21_ni port map ( Y=>nx933, A0=>q_4_10_EXMPLR, A1=>
      q_3_10_EXMPLR, S0=>nx1454);
   gen_regs_3_regi_reg_q_10 : dffr port map ( Q=>q_3_10_EXMPLR, QB=>OPEN, D
      =>nx923, CLK=>nx1506, R=>nx1480);
   ix924 : mux21_ni port map ( Y=>nx923, A0=>q_3_10_EXMPLR, A1=>
      q_2_10_EXMPLR, S0=>nx1454);
   gen_regs_2_regi_reg_q_10 : dffr port map ( Q=>q_2_10_EXMPLR, QB=>OPEN, D
      =>nx913, CLK=>nx1506, R=>nx1480);
   ix914 : mux21_ni port map ( Y=>nx913, A0=>q_2_10_EXMPLR, A1=>
      q_1_10_EXMPLR, S0=>nx1454);
   gen_regs_1_regi_reg_q_10 : dffr port map ( Q=>q_1_10_EXMPLR, QB=>OPEN, D
      =>nx903, CLK=>nx1506, R=>nx1480);
   ix904 : mux21_ni port map ( Y=>nx903, A0=>q_1_10_EXMPLR, A1=>
      q_0_10_EXMPLR, S0=>nx1454);
   reg0_reg_q_10 : dffr port map ( Q=>q_0_10_EXMPLR, QB=>OPEN, D=>nx893, CLK
      =>nx1506, R=>nx1480);
   ix894 : mux21_ni port map ( Y=>nx893, A0=>q_0_10_EXMPLR, A1=>d(10), S0=>
      nx1454);
   gen_regs_4_regi_reg_q_11 : dffr port map ( Q=>q_4_11_EXMPLR, QB=>OPEN, D
      =>nx983, CLK=>nx1508, R=>nx1482);
   ix984 : mux21_ni port map ( Y=>nx983, A0=>q_4_11_EXMPLR, A1=>
      q_3_11_EXMPLR, S0=>nx1456);
   gen_regs_3_regi_reg_q_11 : dffr port map ( Q=>q_3_11_EXMPLR, QB=>OPEN, D
      =>nx973, CLK=>nx1508, R=>nx1482);
   ix974 : mux21_ni port map ( Y=>nx973, A0=>q_3_11_EXMPLR, A1=>
      q_2_11_EXMPLR, S0=>nx1456);
   gen_regs_2_regi_reg_q_11 : dffr port map ( Q=>q_2_11_EXMPLR, QB=>OPEN, D
      =>nx963, CLK=>nx1508, R=>nx1482);
   ix964 : mux21_ni port map ( Y=>nx963, A0=>q_2_11_EXMPLR, A1=>
      q_1_11_EXMPLR, S0=>nx1456);
   gen_regs_1_regi_reg_q_11 : dffr port map ( Q=>q_1_11_EXMPLR, QB=>OPEN, D
      =>nx953, CLK=>nx1508, R=>nx1482);
   ix954 : mux21_ni port map ( Y=>nx953, A0=>q_1_11_EXMPLR, A1=>
      q_0_11_EXMPLR, S0=>nx1456);
   reg0_reg_q_11 : dffr port map ( Q=>q_0_11_EXMPLR, QB=>OPEN, D=>nx943, CLK
      =>nx1506, R=>nx1480);
   ix944 : mux21_ni port map ( Y=>nx943, A0=>q_0_11_EXMPLR, A1=>d(11), S0=>
      nx1454);
   gen_regs_4_regi_reg_q_12 : dffr port map ( Q=>q_4_12_EXMPLR, QB=>OPEN, D
      =>nx1033, CLK=>nx1510, R=>nx1484);
   ix1034 : mux21_ni port map ( Y=>nx1033, A0=>q_4_12_EXMPLR, A1=>
      q_3_12_EXMPLR, S0=>nx1458);
   gen_regs_3_regi_reg_q_12 : dffr port map ( Q=>q_3_12_EXMPLR, QB=>OPEN, D
      =>nx1023, CLK=>nx1510, R=>nx1484);
   ix1024 : mux21_ni port map ( Y=>nx1023, A0=>q_3_12_EXMPLR, A1=>
      q_2_12_EXMPLR, S0=>nx1458);
   gen_regs_2_regi_reg_q_12 : dffr port map ( Q=>q_2_12_EXMPLR, QB=>OPEN, D
      =>nx1013, CLK=>nx1508, R=>nx1482);
   ix1014 : mux21_ni port map ( Y=>nx1013, A0=>q_2_12_EXMPLR, A1=>
      q_1_12_EXMPLR, S0=>nx1456);
   gen_regs_1_regi_reg_q_12 : dffr port map ( Q=>q_1_12_EXMPLR, QB=>OPEN, D
      =>nx1003, CLK=>nx1508, R=>nx1482);
   ix1004 : mux21_ni port map ( Y=>nx1003, A0=>q_1_12_EXMPLR, A1=>
      q_0_12_EXMPLR, S0=>nx1456);
   reg0_reg_q_12 : dffr port map ( Q=>q_0_12_EXMPLR, QB=>OPEN, D=>nx993, CLK
      =>nx1508, R=>nx1482);
   ix994 : mux21_ni port map ( Y=>nx993, A0=>q_0_12_EXMPLR, A1=>d(12), S0=>
      nx1456);
   gen_regs_4_regi_reg_q_13 : dffr port map ( Q=>q_4_13_EXMPLR, QB=>OPEN, D
      =>nx1083, CLK=>nx1510, R=>nx1484);
   ix1084 : mux21_ni port map ( Y=>nx1083, A0=>q_4_13_EXMPLR, A1=>
      q_3_13_EXMPLR, S0=>nx1458);
   gen_regs_3_regi_reg_q_13 : dffr port map ( Q=>q_3_13_EXMPLR, QB=>OPEN, D
      =>nx1073, CLK=>nx1510, R=>nx1484);
   ix1074 : mux21_ni port map ( Y=>nx1073, A0=>q_3_13_EXMPLR, A1=>
      q_2_13_EXMPLR, S0=>nx1458);
   gen_regs_2_regi_reg_q_13 : dffr port map ( Q=>q_2_13_EXMPLR, QB=>OPEN, D
      =>nx1063, CLK=>nx1510, R=>nx1484);
   ix1064 : mux21_ni port map ( Y=>nx1063, A0=>q_2_13_EXMPLR, A1=>
      q_1_13_EXMPLR, S0=>nx1458);
   gen_regs_1_regi_reg_q_13 : dffr port map ( Q=>q_1_13_EXMPLR, QB=>OPEN, D
      =>nx1053, CLK=>nx1510, R=>nx1484);
   ix1054 : mux21_ni port map ( Y=>nx1053, A0=>q_1_13_EXMPLR, A1=>
      q_0_13_EXMPLR, S0=>nx1458);
   reg0_reg_q_13 : dffr port map ( Q=>q_0_13_EXMPLR, QB=>OPEN, D=>nx1043, 
      CLK=>nx1510, R=>nx1484);
   ix1044 : mux21_ni port map ( Y=>nx1043, A0=>q_0_13_EXMPLR, A1=>d(13), S0
      =>nx1458);
   gen_regs_4_regi_reg_q_14 : dffr port map ( Q=>q_4_14_EXMPLR, QB=>OPEN, D
      =>nx1133, CLK=>nx1512, R=>nx1486);
   ix1134 : mux21_ni port map ( Y=>nx1133, A0=>q_4_14_EXMPLR, A1=>
      q_3_14_EXMPLR, S0=>nx1460);
   gen_regs_3_regi_reg_q_14 : dffr port map ( Q=>q_3_14_EXMPLR, QB=>OPEN, D
      =>nx1123, CLK=>nx1512, R=>nx1486);
   ix1124 : mux21_ni port map ( Y=>nx1123, A0=>q_3_14_EXMPLR, A1=>
      q_2_14_EXMPLR, S0=>nx1460);
   gen_regs_2_regi_reg_q_14 : dffr port map ( Q=>q_2_14_EXMPLR, QB=>OPEN, D
      =>nx1113, CLK=>nx1512, R=>nx1486);
   ix1114 : mux21_ni port map ( Y=>nx1113, A0=>q_2_14_EXMPLR, A1=>
      q_1_14_EXMPLR, S0=>nx1460);
   gen_regs_1_regi_reg_q_14 : dffr port map ( Q=>q_1_14_EXMPLR, QB=>OPEN, D
      =>nx1103, CLK=>nx1512, R=>nx1486);
   ix1104 : mux21_ni port map ( Y=>nx1103, A0=>q_1_14_EXMPLR, A1=>
      q_0_14_EXMPLR, S0=>nx1460);
   reg0_reg_q_14 : dffr port map ( Q=>q_0_14_EXMPLR, QB=>OPEN, D=>nx1093, 
      CLK=>nx1512, R=>nx1486);
   ix1094 : mux21_ni port map ( Y=>nx1093, A0=>q_0_14_EXMPLR, A1=>d(14), S0
      =>nx1460);
   gen_regs_4_regi_reg_q_15 : dffr port map ( Q=>q_4_15_EXMPLR, QB=>OPEN, D
      =>nx1183, CLK=>nx1514, R=>nx1488);
   ix1184 : mux21_ni port map ( Y=>nx1183, A0=>q_4_15_EXMPLR, A1=>
      q_3_15_EXMPLR, S0=>nx1462);
   gen_regs_3_regi_reg_q_15 : dffr port map ( Q=>q_3_15_EXMPLR, QB=>OPEN, D
      =>nx1173, CLK=>nx1514, R=>nx1488);
   ix1174 : mux21_ni port map ( Y=>nx1173, A0=>q_3_15_EXMPLR, A1=>
      q_2_15_EXMPLR, S0=>nx1462);
   gen_regs_2_regi_reg_q_15 : dffr port map ( Q=>q_2_15_EXMPLR, QB=>OPEN, D
      =>nx1163, CLK=>nx1514, R=>nx1488);
   ix1164 : mux21_ni port map ( Y=>nx1163, A0=>q_2_15_EXMPLR, A1=>
      q_1_15_EXMPLR, S0=>nx1462);
   gen_regs_1_regi_reg_q_15 : dffr port map ( Q=>q_1_15_EXMPLR, QB=>OPEN, D
      =>nx1153, CLK=>nx1512, R=>nx1486);
   ix1154 : mux21_ni port map ( Y=>nx1153, A0=>q_1_15_EXMPLR, A1=>
      q_0_15_EXMPLR, S0=>nx1460);
   reg0_reg_q_15 : dffr port map ( Q=>q_0_15_EXMPLR, QB=>OPEN, D=>nx1143, 
      CLK=>nx1512, R=>nx1486);
   ix1144 : mux21_ni port map ( Y=>nx1143, A0=>q_0_15_EXMPLR, A1=>d(15), S0
      =>nx1460);
   ix1439 : inv02 port map ( Y=>nx1440, A=>nx1516);
   ix1441 : inv02 port map ( Y=>nx1442, A=>nx1516);
   ix1443 : inv02 port map ( Y=>nx1444, A=>nx1516);
   ix1445 : inv02 port map ( Y=>nx1446, A=>nx1516);
   ix1447 : inv02 port map ( Y=>nx1448, A=>nx1516);
   ix1449 : inv02 port map ( Y=>nx1450, A=>nx1516);
   ix1451 : inv02 port map ( Y=>nx1452, A=>nx1516);
   ix1453 : inv02 port map ( Y=>nx1454, A=>nx1518);
   ix1455 : inv02 port map ( Y=>nx1456, A=>nx1518);
   ix1457 : inv02 port map ( Y=>nx1458, A=>nx1518);
   ix1459 : inv02 port map ( Y=>nx1460, A=>nx1518);
   ix1461 : inv02 port map ( Y=>nx1462, A=>nx1518);
   ix1465 : inv02 port map ( Y=>nx1466, A=>nx1520);
   ix1467 : inv02 port map ( Y=>nx1468, A=>nx1520);
   ix1469 : inv02 port map ( Y=>nx1470, A=>nx1520);
   ix1471 : inv02 port map ( Y=>nx1472, A=>nx1520);
   ix1473 : inv02 port map ( Y=>nx1474, A=>nx1520);
   ix1475 : inv02 port map ( Y=>nx1476, A=>nx1520);
   ix1477 : inv02 port map ( Y=>nx1478, A=>nx1520);
   ix1479 : inv02 port map ( Y=>nx1480, A=>nx1522);
   ix1481 : inv02 port map ( Y=>nx1482, A=>nx1522);
   ix1483 : inv02 port map ( Y=>nx1484, A=>nx1522);
   ix1485 : inv02 port map ( Y=>nx1486, A=>nx1522);
   ix1487 : inv02 port map ( Y=>nx1488, A=>nx1522);
   ix1491 : inv02 port map ( Y=>nx1492, A=>nx1524);
   ix1493 : inv02 port map ( Y=>nx1494, A=>nx1524);
   ix1495 : inv02 port map ( Y=>nx1496, A=>nx1524);
   ix1497 : inv02 port map ( Y=>nx1498, A=>nx1524);
   ix1499 : inv02 port map ( Y=>nx1500, A=>nx1524);
   ix1501 : inv02 port map ( Y=>nx1502, A=>nx1524);
   ix1503 : inv02 port map ( Y=>nx1504, A=>nx1524);
   ix1505 : inv02 port map ( Y=>nx1506, A=>nx1526);
   ix1507 : inv02 port map ( Y=>nx1508, A=>nx1526);
   ix1509 : inv02 port map ( Y=>nx1510, A=>nx1526);
   ix1511 : inv02 port map ( Y=>nx1512, A=>nx1526);
   ix1513 : inv02 port map ( Y=>nx1514, A=>nx1526);
   ix1515 : inv02 port map ( Y=>nx1516, A=>load);
   ix1517 : inv02 port map ( Y=>nx1518, A=>load);
   ix1519 : inv02 port map ( Y=>nx1520, A=>reset);
   ix1521 : inv02 port map ( Y=>nx1522, A=>reset);
   ix1523 : inv02 port map ( Y=>nx1524, A=>clk);
   ix1525 : inv02 port map ( Y=>nx1526, A=>clk);
end Dataflow ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Cache_5_16_28_5 is
   port (
      in_word : IN std_logic_vector (15 DOWNTO 0) ;
      cache_in_sel : IN std_logic_vector (4 DOWNTO 0) ;
      cache_out_sel : IN std_logic_vector (4 DOWNTO 0) ;
      decoder_enable : IN std_logic ;
      out_column_0_15 : OUT std_logic ;
      out_column_0_14 : OUT std_logic ;
      out_column_0_13 : OUT std_logic ;
      out_column_0_12 : OUT std_logic ;
      out_column_0_11 : OUT std_logic ;
      out_column_0_10 : OUT std_logic ;
      out_column_0_9 : OUT std_logic ;
      out_column_0_8 : OUT std_logic ;
      out_column_0_7 : OUT std_logic ;
      out_column_0_6 : OUT std_logic ;
      out_column_0_5 : OUT std_logic ;
      out_column_0_4 : OUT std_logic ;
      out_column_0_3 : OUT std_logic ;
      out_column_0_2 : OUT std_logic ;
      out_column_0_1 : OUT std_logic ;
      out_column_0_0 : OUT std_logic ;
      out_column_1_15 : OUT std_logic ;
      out_column_1_14 : OUT std_logic ;
      out_column_1_13 : OUT std_logic ;
      out_column_1_12 : OUT std_logic ;
      out_column_1_11 : OUT std_logic ;
      out_column_1_10 : OUT std_logic ;
      out_column_1_9 : OUT std_logic ;
      out_column_1_8 : OUT std_logic ;
      out_column_1_7 : OUT std_logic ;
      out_column_1_6 : OUT std_logic ;
      out_column_1_5 : OUT std_logic ;
      out_column_1_4 : OUT std_logic ;
      out_column_1_3 : OUT std_logic ;
      out_column_1_2 : OUT std_logic ;
      out_column_1_1 : OUT std_logic ;
      out_column_1_0 : OUT std_logic ;
      out_column_2_15 : OUT std_logic ;
      out_column_2_14 : OUT std_logic ;
      out_column_2_13 : OUT std_logic ;
      out_column_2_12 : OUT std_logic ;
      out_column_2_11 : OUT std_logic ;
      out_column_2_10 : OUT std_logic ;
      out_column_2_9 : OUT std_logic ;
      out_column_2_8 : OUT std_logic ;
      out_column_2_7 : OUT std_logic ;
      out_column_2_6 : OUT std_logic ;
      out_column_2_5 : OUT std_logic ;
      out_column_2_4 : OUT std_logic ;
      out_column_2_3 : OUT std_logic ;
      out_column_2_2 : OUT std_logic ;
      out_column_2_1 : OUT std_logic ;
      out_column_2_0 : OUT std_logic ;
      out_column_3_15 : OUT std_logic ;
      out_column_3_14 : OUT std_logic ;
      out_column_3_13 : OUT std_logic ;
      out_column_3_12 : OUT std_logic ;
      out_column_3_11 : OUT std_logic ;
      out_column_3_10 : OUT std_logic ;
      out_column_3_9 : OUT std_logic ;
      out_column_3_8 : OUT std_logic ;
      out_column_3_7 : OUT std_logic ;
      out_column_3_6 : OUT std_logic ;
      out_column_3_5 : OUT std_logic ;
      out_column_3_4 : OUT std_logic ;
      out_column_3_3 : OUT std_logic ;
      out_column_3_2 : OUT std_logic ;
      out_column_3_1 : OUT std_logic ;
      out_column_3_0 : OUT std_logic ;
      out_column_4_15 : OUT std_logic ;
      out_column_4_14 : OUT std_logic ;
      out_column_4_13 : OUT std_logic ;
      out_column_4_12 : OUT std_logic ;
      out_column_4_11 : OUT std_logic ;
      out_column_4_10 : OUT std_logic ;
      out_column_4_9 : OUT std_logic ;
      out_column_4_8 : OUT std_logic ;
      out_column_4_7 : OUT std_logic ;
      out_column_4_6 : OUT std_logic ;
      out_column_4_5 : OUT std_logic ;
      out_column_4_4 : OUT std_logic ;
      out_column_4_3 : OUT std_logic ;
      out_column_4_2 : OUT std_logic ;
      out_column_4_1 : OUT std_logic ;
      out_column_4_0 : OUT std_logic ;
      clk : IN std_logic ;
      reset : IN std_logic) ;
end Cache_5_16_28_5 ;

architecture Dataflow of Cache_5_16_28_5 is
   component Queue_5
      port (
         d : IN std_logic_vector (15 DOWNTO 0) ;
         q_0_15 : OUT std_logic ;
         q_0_14 : OUT std_logic ;
         q_0_13 : OUT std_logic ;
         q_0_12 : OUT std_logic ;
         q_0_11 : OUT std_logic ;
         q_0_10 : OUT std_logic ;
         q_0_9 : OUT std_logic ;
         q_0_8 : OUT std_logic ;
         q_0_7 : OUT std_logic ;
         q_0_6 : OUT std_logic ;
         q_0_5 : OUT std_logic ;
         q_0_4 : OUT std_logic ;
         q_0_3 : OUT std_logic ;
         q_0_2 : OUT std_logic ;
         q_0_1 : OUT std_logic ;
         q_0_0 : OUT std_logic ;
         q_1_15 : OUT std_logic ;
         q_1_14 : OUT std_logic ;
         q_1_13 : OUT std_logic ;
         q_1_12 : OUT std_logic ;
         q_1_11 : OUT std_logic ;
         q_1_10 : OUT std_logic ;
         q_1_9 : OUT std_logic ;
         q_1_8 : OUT std_logic ;
         q_1_7 : OUT std_logic ;
         q_1_6 : OUT std_logic ;
         q_1_5 : OUT std_logic ;
         q_1_4 : OUT std_logic ;
         q_1_3 : OUT std_logic ;
         q_1_2 : OUT std_logic ;
         q_1_1 : OUT std_logic ;
         q_1_0 : OUT std_logic ;
         q_2_15 : OUT std_logic ;
         q_2_14 : OUT std_logic ;
         q_2_13 : OUT std_logic ;
         q_2_12 : OUT std_logic ;
         q_2_11 : OUT std_logic ;
         q_2_10 : OUT std_logic ;
         q_2_9 : OUT std_logic ;
         q_2_8 : OUT std_logic ;
         q_2_7 : OUT std_logic ;
         q_2_6 : OUT std_logic ;
         q_2_5 : OUT std_logic ;
         q_2_4 : OUT std_logic ;
         q_2_3 : OUT std_logic ;
         q_2_2 : OUT std_logic ;
         q_2_1 : OUT std_logic ;
         q_2_0 : OUT std_logic ;
         q_3_15 : OUT std_logic ;
         q_3_14 : OUT std_logic ;
         q_3_13 : OUT std_logic ;
         q_3_12 : OUT std_logic ;
         q_3_11 : OUT std_logic ;
         q_3_10 : OUT std_logic ;
         q_3_9 : OUT std_logic ;
         q_3_8 : OUT std_logic ;
         q_3_7 : OUT std_logic ;
         q_3_6 : OUT std_logic ;
         q_3_5 : OUT std_logic ;
         q_3_4 : OUT std_logic ;
         q_3_3 : OUT std_logic ;
         q_3_2 : OUT std_logic ;
         q_3_1 : OUT std_logic ;
         q_3_0 : OUT std_logic ;
         q_4_15 : OUT std_logic ;
         q_4_14 : OUT std_logic ;
         q_4_13 : OUT std_logic ;
         q_4_12 : OUT std_logic ;
         q_4_11 : OUT std_logic ;
         q_4_10 : OUT std_logic ;
         q_4_9 : OUT std_logic ;
         q_4_8 : OUT std_logic ;
         q_4_7 : OUT std_logic ;
         q_4_6 : OUT std_logic ;
         q_4_5 : OUT std_logic ;
         q_4_4 : OUT std_logic ;
         q_4_3 : OUT std_logic ;
         q_4_2 : OUT std_logic ;
         q_4_1 : OUT std_logic ;
         q_4_0 : OUT std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         reset : IN std_logic) ;
   end component ;
   signal que_out_0_0_15, que_out_0_0_14, que_out_0_0_13, que_out_0_0_12, 
      que_out_0_0_11, que_out_0_0_10, que_out_0_0_9, que_out_0_0_8, 
      que_out_0_0_7, que_out_0_0_6, que_out_0_0_5, que_out_0_0_4, 
      que_out_0_0_3, que_out_0_0_2, que_out_0_0_1, que_out_0_0_0, 
      que_out_0_1_15, que_out_0_1_14, que_out_0_1_13, que_out_0_1_12, 
      que_out_0_1_11, que_out_0_1_10, que_out_0_1_9, que_out_0_1_8, 
      que_out_0_1_7, que_out_0_1_6, que_out_0_1_5, que_out_0_1_4, 
      que_out_0_1_3, que_out_0_1_2, que_out_0_1_1, que_out_0_1_0, 
      que_out_0_2_15, que_out_0_2_14, que_out_0_2_13, que_out_0_2_12, 
      que_out_0_2_11, que_out_0_2_10, que_out_0_2_9, que_out_0_2_8, 
      que_out_0_2_7, que_out_0_2_6, que_out_0_2_5, que_out_0_2_4, 
      que_out_0_2_3, que_out_0_2_2, que_out_0_2_1, que_out_0_2_0, 
      que_out_0_3_15, que_out_0_3_14, que_out_0_3_13, que_out_0_3_12, 
      que_out_0_3_11, que_out_0_3_10, que_out_0_3_9, que_out_0_3_8, 
      que_out_0_3_7, que_out_0_3_6, que_out_0_3_5, que_out_0_3_4, 
      que_out_0_3_3, que_out_0_3_2, que_out_0_3_1, que_out_0_3_0, 
      que_out_0_4_15, que_out_0_4_14, que_out_0_4_13, que_out_0_4_12, 
      que_out_0_4_11, que_out_0_4_10, que_out_0_4_9, que_out_0_4_8, 
      que_out_0_4_7, que_out_0_4_6, que_out_0_4_5, que_out_0_4_4, 
      que_out_0_4_3, que_out_0_4_2, que_out_0_4_1, que_out_0_4_0, 
      que_out_1_0_15, que_out_1_0_14, que_out_1_0_13, que_out_1_0_12, 
      que_out_1_0_11, que_out_1_0_10, que_out_1_0_9, que_out_1_0_8, 
      que_out_1_0_7, que_out_1_0_6, que_out_1_0_5, que_out_1_0_4, 
      que_out_1_0_3, que_out_1_0_2, que_out_1_0_1, que_out_1_0_0, 
      que_out_1_1_15, que_out_1_1_14, que_out_1_1_13, que_out_1_1_12, 
      que_out_1_1_11, que_out_1_1_10, que_out_1_1_9, que_out_1_1_8, 
      que_out_1_1_7, que_out_1_1_6, que_out_1_1_5, que_out_1_1_4, 
      que_out_1_1_3, que_out_1_1_2, que_out_1_1_1, que_out_1_1_0, 
      que_out_1_2_15, que_out_1_2_14, que_out_1_2_13, que_out_1_2_12, 
      que_out_1_2_11, que_out_1_2_10, que_out_1_2_9, que_out_1_2_8, 
      que_out_1_2_7, que_out_1_2_6, que_out_1_2_5, que_out_1_2_4, 
      que_out_1_2_3, que_out_1_2_2, que_out_1_2_1, que_out_1_2_0, 
      que_out_1_3_15, que_out_1_3_14, que_out_1_3_13, que_out_1_3_12, 
      que_out_1_3_11, que_out_1_3_10, que_out_1_3_9, que_out_1_3_8, 
      que_out_1_3_7, que_out_1_3_6, que_out_1_3_5, que_out_1_3_4, 
      que_out_1_3_3, que_out_1_3_2, que_out_1_3_1, que_out_1_3_0, 
      que_out_1_4_15, que_out_1_4_14, que_out_1_4_13, que_out_1_4_12, 
      que_out_1_4_11, que_out_1_4_10, que_out_1_4_9, que_out_1_4_8, 
      que_out_1_4_7, que_out_1_4_6, que_out_1_4_5, que_out_1_4_4, 
      que_out_1_4_3, que_out_1_4_2, que_out_1_4_1, que_out_1_4_0, 
      que_out_2_0_15, que_out_2_0_14, que_out_2_0_13, que_out_2_0_12, 
      que_out_2_0_11, que_out_2_0_10, que_out_2_0_9, que_out_2_0_8, 
      que_out_2_0_7, que_out_2_0_6, que_out_2_0_5, que_out_2_0_4, 
      que_out_2_0_3, que_out_2_0_2, que_out_2_0_1, que_out_2_0_0, 
      que_out_2_1_15, que_out_2_1_14, que_out_2_1_13, que_out_2_1_12, 
      que_out_2_1_11, que_out_2_1_10, que_out_2_1_9, que_out_2_1_8, 
      que_out_2_1_7, que_out_2_1_6, que_out_2_1_5, que_out_2_1_4, 
      que_out_2_1_3, que_out_2_1_2, que_out_2_1_1, que_out_2_1_0, 
      que_out_2_2_15, que_out_2_2_14, que_out_2_2_13, que_out_2_2_12, 
      que_out_2_2_11, que_out_2_2_10, que_out_2_2_9, que_out_2_2_8, 
      que_out_2_2_7, que_out_2_2_6, que_out_2_2_5, que_out_2_2_4, 
      que_out_2_2_3, que_out_2_2_2, que_out_2_2_1, que_out_2_2_0, 
      que_out_2_3_15, que_out_2_3_14, que_out_2_3_13, que_out_2_3_12, 
      que_out_2_3_11, que_out_2_3_10, que_out_2_3_9, que_out_2_3_8, 
      que_out_2_3_7, que_out_2_3_6, que_out_2_3_5, que_out_2_3_4, 
      que_out_2_3_3, que_out_2_3_2, que_out_2_3_1, que_out_2_3_0, 
      que_out_2_4_15, que_out_2_4_14, que_out_2_4_13, que_out_2_4_12, 
      que_out_2_4_11, que_out_2_4_10, que_out_2_4_9, que_out_2_4_8, 
      que_out_2_4_7, que_out_2_4_6, que_out_2_4_5, que_out_2_4_4, 
      que_out_2_4_3, que_out_2_4_2, que_out_2_4_1, que_out_2_4_0, 
      que_out_3_0_15, que_out_3_0_14, que_out_3_0_13, que_out_3_0_12, 
      que_out_3_0_11, que_out_3_0_10, que_out_3_0_9, que_out_3_0_8, 
      que_out_3_0_7, que_out_3_0_6, que_out_3_0_5, que_out_3_0_4, 
      que_out_3_0_3, que_out_3_0_2, que_out_3_0_1, que_out_3_0_0, 
      que_out_3_1_15, que_out_3_1_14, que_out_3_1_13, que_out_3_1_12, 
      que_out_3_1_11, que_out_3_1_10, que_out_3_1_9, que_out_3_1_8, 
      que_out_3_1_7, que_out_3_1_6, que_out_3_1_5, que_out_3_1_4, 
      que_out_3_1_3, que_out_3_1_2, que_out_3_1_1, que_out_3_1_0, 
      que_out_3_2_15, que_out_3_2_14, que_out_3_2_13, que_out_3_2_12, 
      que_out_3_2_11, que_out_3_2_10, que_out_3_2_9, que_out_3_2_8, 
      que_out_3_2_7, que_out_3_2_6, que_out_3_2_5, que_out_3_2_4, 
      que_out_3_2_3, que_out_3_2_2, que_out_3_2_1, que_out_3_2_0, 
      que_out_3_3_15, que_out_3_3_14, que_out_3_3_13, que_out_3_3_12, 
      que_out_3_3_11, que_out_3_3_10, que_out_3_3_9, que_out_3_3_8, 
      que_out_3_3_7, que_out_3_3_6, que_out_3_3_5, que_out_3_3_4, 
      que_out_3_3_3, que_out_3_3_2, que_out_3_3_1, que_out_3_3_0, 
      que_out_3_4_15, que_out_3_4_14, que_out_3_4_13, que_out_3_4_12, 
      que_out_3_4_11, que_out_3_4_10, que_out_3_4_9, que_out_3_4_8, 
      que_out_3_4_7, que_out_3_4_6, que_out_3_4_5, que_out_3_4_4, 
      que_out_3_4_3, que_out_3_4_2, que_out_3_4_1, que_out_3_4_0, 
      que_out_4_0_15, que_out_4_0_14, que_out_4_0_13, que_out_4_0_12, 
      que_out_4_0_11, que_out_4_0_10, que_out_4_0_9, que_out_4_0_8, 
      que_out_4_0_7, que_out_4_0_6, que_out_4_0_5, que_out_4_0_4, 
      que_out_4_0_3, que_out_4_0_2, que_out_4_0_1, que_out_4_0_0, 
      que_out_4_1_15, que_out_4_1_14, que_out_4_1_13, que_out_4_1_12, 
      que_out_4_1_11, que_out_4_1_10, que_out_4_1_9, que_out_4_1_8, 
      que_out_4_1_7, que_out_4_1_6, que_out_4_1_5, que_out_4_1_4, 
      que_out_4_1_3, que_out_4_1_2, que_out_4_1_1, que_out_4_1_0, 
      que_out_4_2_15, que_out_4_2_14, que_out_4_2_13, que_out_4_2_12, 
      que_out_4_2_11, que_out_4_2_10, que_out_4_2_9, que_out_4_2_8, 
      que_out_4_2_7, que_out_4_2_6, que_out_4_2_5, que_out_4_2_4, 
      que_out_4_2_3, que_out_4_2_2, que_out_4_2_1, que_out_4_2_0, 
      que_out_4_3_15, que_out_4_3_14, que_out_4_3_13, que_out_4_3_12, 
      que_out_4_3_11, que_out_4_3_10, que_out_4_3_9, que_out_4_3_8, 
      que_out_4_3_7, que_out_4_3_6, que_out_4_3_5, que_out_4_3_4, 
      que_out_4_3_3, que_out_4_3_2, que_out_4_3_1, que_out_4_3_0, 
      que_out_4_4_15, que_out_4_4_14, que_out_4_4_13, que_out_4_4_12, 
      que_out_4_4_11, que_out_4_4_10, que_out_4_4_9, que_out_4_4_8, 
      que_out_4_4_7, que_out_4_4_6, que_out_4_4_5, que_out_4_4_4, 
      que_out_4_4_3, que_out_4_4_2, que_out_4_4_1, que_out_4_4_0, 
      que_out_5_0_15, que_out_5_0_14, que_out_5_0_13, que_out_5_0_12, 
      que_out_5_0_11, que_out_5_0_10, que_out_5_0_9, que_out_5_0_8, 
      que_out_5_0_7, que_out_5_0_6, que_out_5_0_5, que_out_5_0_4, 
      que_out_5_0_3, que_out_5_0_2, que_out_5_0_1, que_out_5_0_0, 
      que_out_5_1_15, que_out_5_1_14, que_out_5_1_13, que_out_5_1_12, 
      que_out_5_1_11, que_out_5_1_10, que_out_5_1_9, que_out_5_1_8, 
      que_out_5_1_7, que_out_5_1_6, que_out_5_1_5, que_out_5_1_4, 
      que_out_5_1_3, que_out_5_1_2, que_out_5_1_1, que_out_5_1_0, 
      que_out_5_2_15, que_out_5_2_14, que_out_5_2_13, que_out_5_2_12, 
      que_out_5_2_11, que_out_5_2_10, que_out_5_2_9, que_out_5_2_8, 
      que_out_5_2_7, que_out_5_2_6, que_out_5_2_5, que_out_5_2_4, 
      que_out_5_2_3, que_out_5_2_2, que_out_5_2_1, que_out_5_2_0, 
      que_out_5_3_15, que_out_5_3_14, que_out_5_3_13, que_out_5_3_12, 
      que_out_5_3_11, que_out_5_3_10, que_out_5_3_9, que_out_5_3_8, 
      que_out_5_3_7, que_out_5_3_6, que_out_5_3_5, que_out_5_3_4, 
      que_out_5_3_3, que_out_5_3_2, que_out_5_3_1, que_out_5_3_0, 
      que_out_5_4_15, que_out_5_4_14, que_out_5_4_13, que_out_5_4_12, 
      que_out_5_4_11, que_out_5_4_10, que_out_5_4_9, que_out_5_4_8, 
      que_out_5_4_7, que_out_5_4_6, que_out_5_4_5, que_out_5_4_4, 
      que_out_5_4_3, que_out_5_4_2, que_out_5_4_1, que_out_5_4_0, 
      que_out_6_0_15, que_out_6_0_14, que_out_6_0_13, que_out_6_0_12, 
      que_out_6_0_11, que_out_6_0_10, que_out_6_0_9, que_out_6_0_8, 
      que_out_6_0_7, que_out_6_0_6, que_out_6_0_5, que_out_6_0_4, 
      que_out_6_0_3, que_out_6_0_2, que_out_6_0_1, que_out_6_0_0, 
      que_out_6_1_15, que_out_6_1_14, que_out_6_1_13, que_out_6_1_12, 
      que_out_6_1_11, que_out_6_1_10, que_out_6_1_9, que_out_6_1_8, 
      que_out_6_1_7, que_out_6_1_6, que_out_6_1_5, que_out_6_1_4, 
      que_out_6_1_3, que_out_6_1_2, que_out_6_1_1, que_out_6_1_0, 
      que_out_6_2_15, que_out_6_2_14, que_out_6_2_13, que_out_6_2_12, 
      que_out_6_2_11, que_out_6_2_10, que_out_6_2_9, que_out_6_2_8, 
      que_out_6_2_7, que_out_6_2_6, que_out_6_2_5, que_out_6_2_4, 
      que_out_6_2_3, que_out_6_2_2, que_out_6_2_1, que_out_6_2_0, 
      que_out_6_3_15, que_out_6_3_14, que_out_6_3_13, que_out_6_3_12, 
      que_out_6_3_11, que_out_6_3_10, que_out_6_3_9, que_out_6_3_8, 
      que_out_6_3_7, que_out_6_3_6, que_out_6_3_5, que_out_6_3_4, 
      que_out_6_3_3, que_out_6_3_2, que_out_6_3_1, que_out_6_3_0, 
      que_out_6_4_15, que_out_6_4_14, que_out_6_4_13, que_out_6_4_12, 
      que_out_6_4_11, que_out_6_4_10, que_out_6_4_9, que_out_6_4_8, 
      que_out_6_4_7, que_out_6_4_6, que_out_6_4_5, que_out_6_4_4, 
      que_out_6_4_3, que_out_6_4_2, que_out_6_4_1, que_out_6_4_0, 
      que_out_7_0_15, que_out_7_0_14, que_out_7_0_13, que_out_7_0_12, 
      que_out_7_0_11, que_out_7_0_10, que_out_7_0_9, que_out_7_0_8, 
      que_out_7_0_7, que_out_7_0_6, que_out_7_0_5, que_out_7_0_4, 
      que_out_7_0_3, que_out_7_0_2, que_out_7_0_1, que_out_7_0_0, 
      que_out_7_1_15, que_out_7_1_14, que_out_7_1_13, que_out_7_1_12, 
      que_out_7_1_11, que_out_7_1_10, que_out_7_1_9, que_out_7_1_8, 
      que_out_7_1_7, que_out_7_1_6, que_out_7_1_5, que_out_7_1_4, 
      que_out_7_1_3, que_out_7_1_2, que_out_7_1_1, que_out_7_1_0, 
      que_out_7_2_15, que_out_7_2_14, que_out_7_2_13, que_out_7_2_12, 
      que_out_7_2_11, que_out_7_2_10, que_out_7_2_9, que_out_7_2_8, 
      que_out_7_2_7, que_out_7_2_6, que_out_7_2_5, que_out_7_2_4, 
      que_out_7_2_3, que_out_7_2_2, que_out_7_2_1, que_out_7_2_0, 
      que_out_7_3_15, que_out_7_3_14, que_out_7_3_13, que_out_7_3_12, 
      que_out_7_3_11, que_out_7_3_10, que_out_7_3_9, que_out_7_3_8, 
      que_out_7_3_7, que_out_7_3_6, que_out_7_3_5, que_out_7_3_4, 
      que_out_7_3_3, que_out_7_3_2, que_out_7_3_1, que_out_7_3_0, 
      que_out_7_4_15, que_out_7_4_14, que_out_7_4_13, que_out_7_4_12, 
      que_out_7_4_11, que_out_7_4_10, que_out_7_4_9, que_out_7_4_8, 
      que_out_7_4_7, que_out_7_4_6, que_out_7_4_5, que_out_7_4_4, 
      que_out_7_4_3, que_out_7_4_2, que_out_7_4_1, que_out_7_4_0, 
      que_out_8_0_15, que_out_8_0_14, que_out_8_0_13, que_out_8_0_12, 
      que_out_8_0_11, que_out_8_0_10, que_out_8_0_9, que_out_8_0_8, 
      que_out_8_0_7, que_out_8_0_6, que_out_8_0_5, que_out_8_0_4, 
      que_out_8_0_3, que_out_8_0_2, que_out_8_0_1, que_out_8_0_0, 
      que_out_8_1_15, que_out_8_1_14, que_out_8_1_13, que_out_8_1_12, 
      que_out_8_1_11, que_out_8_1_10, que_out_8_1_9, que_out_8_1_8, 
      que_out_8_1_7, que_out_8_1_6, que_out_8_1_5, que_out_8_1_4, 
      que_out_8_1_3, que_out_8_1_2, que_out_8_1_1, que_out_8_1_0, 
      que_out_8_2_15, que_out_8_2_14, que_out_8_2_13, que_out_8_2_12, 
      que_out_8_2_11, que_out_8_2_10, que_out_8_2_9, que_out_8_2_8, 
      que_out_8_2_7, que_out_8_2_6, que_out_8_2_5, que_out_8_2_4, 
      que_out_8_2_3, que_out_8_2_2, que_out_8_2_1, que_out_8_2_0, 
      que_out_8_3_15, que_out_8_3_14, que_out_8_3_13, que_out_8_3_12, 
      que_out_8_3_11, que_out_8_3_10, que_out_8_3_9, que_out_8_3_8, 
      que_out_8_3_7, que_out_8_3_6, que_out_8_3_5, que_out_8_3_4, 
      que_out_8_3_3, que_out_8_3_2, que_out_8_3_1, que_out_8_3_0, 
      que_out_8_4_15, que_out_8_4_14, que_out_8_4_13, que_out_8_4_12, 
      que_out_8_4_11, que_out_8_4_10, que_out_8_4_9, que_out_8_4_8, 
      que_out_8_4_7, que_out_8_4_6, que_out_8_4_5, que_out_8_4_4, 
      que_out_8_4_3, que_out_8_4_2, que_out_8_4_1, que_out_8_4_0, 
      que_out_9_0_15, que_out_9_0_14, que_out_9_0_13, que_out_9_0_12, 
      que_out_9_0_11, que_out_9_0_10, que_out_9_0_9, que_out_9_0_8, 
      que_out_9_0_7, que_out_9_0_6, que_out_9_0_5, que_out_9_0_4, 
      que_out_9_0_3, que_out_9_0_2, que_out_9_0_1, que_out_9_0_0, 
      que_out_9_1_15, que_out_9_1_14, que_out_9_1_13, que_out_9_1_12, 
      que_out_9_1_11, que_out_9_1_10, que_out_9_1_9, que_out_9_1_8, 
      que_out_9_1_7, que_out_9_1_6, que_out_9_1_5, que_out_9_1_4, 
      que_out_9_1_3, que_out_9_1_2, que_out_9_1_1, que_out_9_1_0, 
      que_out_9_2_15, que_out_9_2_14, que_out_9_2_13, que_out_9_2_12, 
      que_out_9_2_11, que_out_9_2_10, que_out_9_2_9, que_out_9_2_8, 
      que_out_9_2_7, que_out_9_2_6, que_out_9_2_5, que_out_9_2_4, 
      que_out_9_2_3, que_out_9_2_2, que_out_9_2_1, que_out_9_2_0, 
      que_out_9_3_15, que_out_9_3_14, que_out_9_3_13, que_out_9_3_12, 
      que_out_9_3_11, que_out_9_3_10, que_out_9_3_9, que_out_9_3_8, 
      que_out_9_3_7, que_out_9_3_6, que_out_9_3_5, que_out_9_3_4, 
      que_out_9_3_3, que_out_9_3_2, que_out_9_3_1, que_out_9_3_0, 
      que_out_9_4_15, que_out_9_4_14, que_out_9_4_13, que_out_9_4_12, 
      que_out_9_4_11, que_out_9_4_10, que_out_9_4_9, que_out_9_4_8, 
      que_out_9_4_7, que_out_9_4_6, que_out_9_4_5, que_out_9_4_4, 
      que_out_9_4_3, que_out_9_4_2, que_out_9_4_1, que_out_9_4_0, 
      que_out_10_0_15, que_out_10_0_14, que_out_10_0_13, que_out_10_0_12, 
      que_out_10_0_11, que_out_10_0_10, que_out_10_0_9, que_out_10_0_8, 
      que_out_10_0_7, que_out_10_0_6, que_out_10_0_5, que_out_10_0_4, 
      que_out_10_0_3, que_out_10_0_2, que_out_10_0_1, que_out_10_0_0, 
      que_out_10_1_15, que_out_10_1_14, que_out_10_1_13, que_out_10_1_12, 
      que_out_10_1_11, que_out_10_1_10, que_out_10_1_9, que_out_10_1_8, 
      que_out_10_1_7, que_out_10_1_6, que_out_10_1_5, que_out_10_1_4, 
      que_out_10_1_3, que_out_10_1_2, que_out_10_1_1, que_out_10_1_0, 
      que_out_10_2_15, que_out_10_2_14, que_out_10_2_13, que_out_10_2_12, 
      que_out_10_2_11, que_out_10_2_10, que_out_10_2_9, que_out_10_2_8, 
      que_out_10_2_7, que_out_10_2_6, que_out_10_2_5, que_out_10_2_4, 
      que_out_10_2_3, que_out_10_2_2, que_out_10_2_1, que_out_10_2_0, 
      que_out_10_3_15, que_out_10_3_14, que_out_10_3_13, que_out_10_3_12, 
      que_out_10_3_11, que_out_10_3_10, que_out_10_3_9, que_out_10_3_8, 
      que_out_10_3_7, que_out_10_3_6, que_out_10_3_5, que_out_10_3_4, 
      que_out_10_3_3, que_out_10_3_2, que_out_10_3_1, que_out_10_3_0, 
      que_out_10_4_15, que_out_10_4_14, que_out_10_4_13, que_out_10_4_12, 
      que_out_10_4_11, que_out_10_4_10, que_out_10_4_9, que_out_10_4_8, 
      que_out_10_4_7, que_out_10_4_6, que_out_10_4_5, que_out_10_4_4, 
      que_out_10_4_3, que_out_10_4_2, que_out_10_4_1, que_out_10_4_0, 
      que_out_11_0_15, que_out_11_0_14, que_out_11_0_13, que_out_11_0_12, 
      que_out_11_0_11, que_out_11_0_10, que_out_11_0_9, que_out_11_0_8, 
      que_out_11_0_7, que_out_11_0_6, que_out_11_0_5, que_out_11_0_4, 
      que_out_11_0_3, que_out_11_0_2, que_out_11_0_1, que_out_11_0_0, 
      que_out_11_1_15, que_out_11_1_14, que_out_11_1_13, que_out_11_1_12, 
      que_out_11_1_11, que_out_11_1_10, que_out_11_1_9, que_out_11_1_8, 
      que_out_11_1_7, que_out_11_1_6, que_out_11_1_5, que_out_11_1_4, 
      que_out_11_1_3, que_out_11_1_2, que_out_11_1_1, que_out_11_1_0, 
      que_out_11_2_15, que_out_11_2_14, que_out_11_2_13, que_out_11_2_12, 
      que_out_11_2_11, que_out_11_2_10, que_out_11_2_9, que_out_11_2_8, 
      que_out_11_2_7, que_out_11_2_6, que_out_11_2_5, que_out_11_2_4, 
      que_out_11_2_3, que_out_11_2_2, que_out_11_2_1, que_out_11_2_0, 
      que_out_11_3_15, que_out_11_3_14, que_out_11_3_13, que_out_11_3_12, 
      que_out_11_3_11, que_out_11_3_10, que_out_11_3_9, que_out_11_3_8, 
      que_out_11_3_7, que_out_11_3_6, que_out_11_3_5, que_out_11_3_4, 
      que_out_11_3_3, que_out_11_3_2, que_out_11_3_1, que_out_11_3_0, 
      que_out_11_4_15, que_out_11_4_14, que_out_11_4_13, que_out_11_4_12, 
      que_out_11_4_11, que_out_11_4_10, que_out_11_4_9, que_out_11_4_8, 
      que_out_11_4_7, que_out_11_4_6, que_out_11_4_5, que_out_11_4_4, 
      que_out_11_4_3, que_out_11_4_2, que_out_11_4_1, que_out_11_4_0, 
      que_out_12_0_15, que_out_12_0_14, que_out_12_0_13, que_out_12_0_12, 
      que_out_12_0_11, que_out_12_0_10, que_out_12_0_9, que_out_12_0_8, 
      que_out_12_0_7, que_out_12_0_6, que_out_12_0_5, que_out_12_0_4, 
      que_out_12_0_3, que_out_12_0_2, que_out_12_0_1, que_out_12_0_0, 
      que_out_12_1_15, que_out_12_1_14, que_out_12_1_13, que_out_12_1_12, 
      que_out_12_1_11, que_out_12_1_10, que_out_12_1_9, que_out_12_1_8, 
      que_out_12_1_7, que_out_12_1_6, que_out_12_1_5, que_out_12_1_4, 
      que_out_12_1_3, que_out_12_1_2, que_out_12_1_1, que_out_12_1_0, 
      que_out_12_2_15, que_out_12_2_14, que_out_12_2_13, que_out_12_2_12, 
      que_out_12_2_11, que_out_12_2_10, que_out_12_2_9, que_out_12_2_8, 
      que_out_12_2_7, que_out_12_2_6, que_out_12_2_5, que_out_12_2_4, 
      que_out_12_2_3, que_out_12_2_2, que_out_12_2_1, que_out_12_2_0, 
      que_out_12_3_15, que_out_12_3_14, que_out_12_3_13, que_out_12_3_12, 
      que_out_12_3_11, que_out_12_3_10, que_out_12_3_9, que_out_12_3_8, 
      que_out_12_3_7, que_out_12_3_6, que_out_12_3_5, que_out_12_3_4, 
      que_out_12_3_3, que_out_12_3_2, que_out_12_3_1, que_out_12_3_0, 
      que_out_12_4_15, que_out_12_4_14, que_out_12_4_13, que_out_12_4_12, 
      que_out_12_4_11, que_out_12_4_10, que_out_12_4_9, que_out_12_4_8, 
      que_out_12_4_7, que_out_12_4_6, que_out_12_4_5, que_out_12_4_4, 
      que_out_12_4_3, que_out_12_4_2, que_out_12_4_1, que_out_12_4_0, 
      que_out_13_0_15, que_out_13_0_14, que_out_13_0_13, que_out_13_0_12, 
      que_out_13_0_11, que_out_13_0_10, que_out_13_0_9, que_out_13_0_8, 
      que_out_13_0_7, que_out_13_0_6, que_out_13_0_5, que_out_13_0_4, 
      que_out_13_0_3, que_out_13_0_2, que_out_13_0_1, que_out_13_0_0, 
      que_out_13_1_15, que_out_13_1_14, que_out_13_1_13, que_out_13_1_12, 
      que_out_13_1_11, que_out_13_1_10, que_out_13_1_9, que_out_13_1_8, 
      que_out_13_1_7, que_out_13_1_6, que_out_13_1_5, que_out_13_1_4, 
      que_out_13_1_3, que_out_13_1_2, que_out_13_1_1, que_out_13_1_0, 
      que_out_13_2_15, que_out_13_2_14, que_out_13_2_13, que_out_13_2_12, 
      que_out_13_2_11, que_out_13_2_10, que_out_13_2_9, que_out_13_2_8, 
      que_out_13_2_7, que_out_13_2_6, que_out_13_2_5, que_out_13_2_4, 
      que_out_13_2_3, que_out_13_2_2, que_out_13_2_1, que_out_13_2_0, 
      que_out_13_3_15, que_out_13_3_14, que_out_13_3_13, que_out_13_3_12, 
      que_out_13_3_11, que_out_13_3_10, que_out_13_3_9, que_out_13_3_8, 
      que_out_13_3_7, que_out_13_3_6, que_out_13_3_5, que_out_13_3_4, 
      que_out_13_3_3, que_out_13_3_2, que_out_13_3_1, que_out_13_3_0, 
      que_out_13_4_15, que_out_13_4_14, que_out_13_4_13, que_out_13_4_12, 
      que_out_13_4_11, que_out_13_4_10, que_out_13_4_9, que_out_13_4_8, 
      que_out_13_4_7, que_out_13_4_6, que_out_13_4_5, que_out_13_4_4, 
      que_out_13_4_3, que_out_13_4_2, que_out_13_4_1, que_out_13_4_0, 
      que_out_14_0_15, que_out_14_0_14, que_out_14_0_13, que_out_14_0_12, 
      que_out_14_0_11, que_out_14_0_10, que_out_14_0_9, que_out_14_0_8, 
      que_out_14_0_7, que_out_14_0_6, que_out_14_0_5, que_out_14_0_4, 
      que_out_14_0_3, que_out_14_0_2, que_out_14_0_1, que_out_14_0_0, 
      que_out_14_1_15, que_out_14_1_14, que_out_14_1_13, que_out_14_1_12, 
      que_out_14_1_11, que_out_14_1_10, que_out_14_1_9, que_out_14_1_8, 
      que_out_14_1_7, que_out_14_1_6, que_out_14_1_5, que_out_14_1_4, 
      que_out_14_1_3, que_out_14_1_2, que_out_14_1_1, que_out_14_1_0, 
      que_out_14_2_15, que_out_14_2_14, que_out_14_2_13, que_out_14_2_12, 
      que_out_14_2_11, que_out_14_2_10, que_out_14_2_9, que_out_14_2_8, 
      que_out_14_2_7, que_out_14_2_6, que_out_14_2_5, que_out_14_2_4, 
      que_out_14_2_3, que_out_14_2_2, que_out_14_2_1, que_out_14_2_0, 
      que_out_14_3_15, que_out_14_3_14, que_out_14_3_13, que_out_14_3_12, 
      que_out_14_3_11, que_out_14_3_10, que_out_14_3_9, que_out_14_3_8, 
      que_out_14_3_7, que_out_14_3_6, que_out_14_3_5, que_out_14_3_4, 
      que_out_14_3_3, que_out_14_3_2, que_out_14_3_1, que_out_14_3_0, 
      que_out_14_4_15, que_out_14_4_14, que_out_14_4_13, que_out_14_4_12, 
      que_out_14_4_11, que_out_14_4_10, que_out_14_4_9, que_out_14_4_8, 
      que_out_14_4_7, que_out_14_4_6, que_out_14_4_5, que_out_14_4_4, 
      que_out_14_4_3, que_out_14_4_2, que_out_14_4_1, que_out_14_4_0, 
      que_out_15_0_15, que_out_15_0_14, que_out_15_0_13, que_out_15_0_12, 
      que_out_15_0_11, que_out_15_0_10, que_out_15_0_9, que_out_15_0_8, 
      que_out_15_0_7, que_out_15_0_6, que_out_15_0_5, que_out_15_0_4, 
      que_out_15_0_3, que_out_15_0_2, que_out_15_0_1, que_out_15_0_0, 
      que_out_15_1_15, que_out_15_1_14, que_out_15_1_13, que_out_15_1_12, 
      que_out_15_1_11, que_out_15_1_10, que_out_15_1_9, que_out_15_1_8, 
      que_out_15_1_7, que_out_15_1_6, que_out_15_1_5, que_out_15_1_4, 
      que_out_15_1_3, que_out_15_1_2, que_out_15_1_1, que_out_15_1_0, 
      que_out_15_2_15, que_out_15_2_14, que_out_15_2_13, que_out_15_2_12, 
      que_out_15_2_11, que_out_15_2_10, que_out_15_2_9, que_out_15_2_8, 
      que_out_15_2_7, que_out_15_2_6, que_out_15_2_5, que_out_15_2_4, 
      que_out_15_2_3, que_out_15_2_2, que_out_15_2_1, que_out_15_2_0, 
      que_out_15_3_15, que_out_15_3_14, que_out_15_3_13, que_out_15_3_12, 
      que_out_15_3_11, que_out_15_3_10, que_out_15_3_9, que_out_15_3_8, 
      que_out_15_3_7, que_out_15_3_6, que_out_15_3_5, que_out_15_3_4, 
      que_out_15_3_3, que_out_15_3_2, que_out_15_3_1, que_out_15_3_0, 
      que_out_15_4_15, que_out_15_4_14, que_out_15_4_13, que_out_15_4_12, 
      que_out_15_4_11, que_out_15_4_10, que_out_15_4_9, que_out_15_4_8, 
      que_out_15_4_7, que_out_15_4_6, que_out_15_4_5, que_out_15_4_4, 
      que_out_15_4_3, que_out_15_4_2, que_out_15_4_1, que_out_15_4_0, 
      que_out_16_0_15, que_out_16_0_14, que_out_16_0_13, que_out_16_0_12, 
      que_out_16_0_11, que_out_16_0_10, que_out_16_0_9, que_out_16_0_8, 
      que_out_16_0_7, que_out_16_0_6, que_out_16_0_5, que_out_16_0_4, 
      que_out_16_0_3, que_out_16_0_2, que_out_16_0_1, que_out_16_0_0, 
      que_out_16_1_15, que_out_16_1_14, que_out_16_1_13, que_out_16_1_12, 
      que_out_16_1_11, que_out_16_1_10, que_out_16_1_9, que_out_16_1_8, 
      que_out_16_1_7, que_out_16_1_6, que_out_16_1_5, que_out_16_1_4, 
      que_out_16_1_3, que_out_16_1_2, que_out_16_1_1, que_out_16_1_0, 
      que_out_16_2_15, que_out_16_2_14, que_out_16_2_13, que_out_16_2_12, 
      que_out_16_2_11, que_out_16_2_10, que_out_16_2_9, que_out_16_2_8, 
      que_out_16_2_7, que_out_16_2_6, que_out_16_2_5, que_out_16_2_4, 
      que_out_16_2_3, que_out_16_2_2, que_out_16_2_1, que_out_16_2_0, 
      que_out_16_3_15, que_out_16_3_14, que_out_16_3_13, que_out_16_3_12, 
      que_out_16_3_11, que_out_16_3_10, que_out_16_3_9, que_out_16_3_8, 
      que_out_16_3_7, que_out_16_3_6, que_out_16_3_5, que_out_16_3_4, 
      que_out_16_3_3, que_out_16_3_2, que_out_16_3_1, que_out_16_3_0, 
      que_out_16_4_15, que_out_16_4_14, que_out_16_4_13, que_out_16_4_12, 
      que_out_16_4_11, que_out_16_4_10, que_out_16_4_9, que_out_16_4_8, 
      que_out_16_4_7, que_out_16_4_6, que_out_16_4_5, que_out_16_4_4, 
      que_out_16_4_3, que_out_16_4_2, que_out_16_4_1, que_out_16_4_0, 
      que_out_17_0_15, que_out_17_0_14, que_out_17_0_13, que_out_17_0_12, 
      que_out_17_0_11, que_out_17_0_10, que_out_17_0_9, que_out_17_0_8, 
      que_out_17_0_7, que_out_17_0_6, que_out_17_0_5, que_out_17_0_4, 
      que_out_17_0_3, que_out_17_0_2, que_out_17_0_1, que_out_17_0_0, 
      que_out_17_1_15, que_out_17_1_14, que_out_17_1_13, que_out_17_1_12, 
      que_out_17_1_11, que_out_17_1_10, que_out_17_1_9, que_out_17_1_8, 
      que_out_17_1_7, que_out_17_1_6, que_out_17_1_5, que_out_17_1_4, 
      que_out_17_1_3, que_out_17_1_2, que_out_17_1_1, que_out_17_1_0, 
      que_out_17_2_15, que_out_17_2_14, que_out_17_2_13, que_out_17_2_12, 
      que_out_17_2_11, que_out_17_2_10, que_out_17_2_9, que_out_17_2_8, 
      que_out_17_2_7, que_out_17_2_6, que_out_17_2_5, que_out_17_2_4, 
      que_out_17_2_3, que_out_17_2_2, que_out_17_2_1, que_out_17_2_0, 
      que_out_17_3_15, que_out_17_3_14, que_out_17_3_13, que_out_17_3_12, 
      que_out_17_3_11, que_out_17_3_10, que_out_17_3_9, que_out_17_3_8, 
      que_out_17_3_7, que_out_17_3_6, que_out_17_3_5, que_out_17_3_4, 
      que_out_17_3_3, que_out_17_3_2, que_out_17_3_1, que_out_17_3_0, 
      que_out_17_4_15, que_out_17_4_14, que_out_17_4_13, que_out_17_4_12, 
      que_out_17_4_11, que_out_17_4_10, que_out_17_4_9, que_out_17_4_8, 
      que_out_17_4_7, que_out_17_4_6, que_out_17_4_5, que_out_17_4_4, 
      que_out_17_4_3, que_out_17_4_2, que_out_17_4_1, que_out_17_4_0, 
      que_out_18_0_15, que_out_18_0_14, que_out_18_0_13, que_out_18_0_12, 
      que_out_18_0_11, que_out_18_0_10, que_out_18_0_9, que_out_18_0_8, 
      que_out_18_0_7, que_out_18_0_6, que_out_18_0_5, que_out_18_0_4, 
      que_out_18_0_3, que_out_18_0_2, que_out_18_0_1, que_out_18_0_0, 
      que_out_18_1_15, que_out_18_1_14, que_out_18_1_13, que_out_18_1_12, 
      que_out_18_1_11, que_out_18_1_10, que_out_18_1_9, que_out_18_1_8, 
      que_out_18_1_7, que_out_18_1_6, que_out_18_1_5, que_out_18_1_4, 
      que_out_18_1_3, que_out_18_1_2, que_out_18_1_1, que_out_18_1_0, 
      que_out_18_2_15, que_out_18_2_14, que_out_18_2_13, que_out_18_2_12, 
      que_out_18_2_11, que_out_18_2_10, que_out_18_2_9, que_out_18_2_8, 
      que_out_18_2_7, que_out_18_2_6, que_out_18_2_5, que_out_18_2_4, 
      que_out_18_2_3, que_out_18_2_2, que_out_18_2_1, que_out_18_2_0, 
      que_out_18_3_15, que_out_18_3_14, que_out_18_3_13, que_out_18_3_12, 
      que_out_18_3_11, que_out_18_3_10, que_out_18_3_9, que_out_18_3_8, 
      que_out_18_3_7, que_out_18_3_6, que_out_18_3_5, que_out_18_3_4, 
      que_out_18_3_3, que_out_18_3_2, que_out_18_3_1, que_out_18_3_0, 
      que_out_18_4_15, que_out_18_4_14, que_out_18_4_13, que_out_18_4_12, 
      que_out_18_4_11, que_out_18_4_10, que_out_18_4_9, que_out_18_4_8, 
      que_out_18_4_7, que_out_18_4_6, que_out_18_4_5, que_out_18_4_4, 
      que_out_18_4_3, que_out_18_4_2, que_out_18_4_1, que_out_18_4_0, 
      que_out_19_0_15, que_out_19_0_14, que_out_19_0_13, que_out_19_0_12, 
      que_out_19_0_11, que_out_19_0_10, que_out_19_0_9, que_out_19_0_8, 
      que_out_19_0_7, que_out_19_0_6, que_out_19_0_5, que_out_19_0_4, 
      que_out_19_0_3, que_out_19_0_2, que_out_19_0_1, que_out_19_0_0, 
      que_out_19_1_15, que_out_19_1_14, que_out_19_1_13, que_out_19_1_12, 
      que_out_19_1_11, que_out_19_1_10, que_out_19_1_9, que_out_19_1_8, 
      que_out_19_1_7, que_out_19_1_6, que_out_19_1_5, que_out_19_1_4, 
      que_out_19_1_3, que_out_19_1_2, que_out_19_1_1, que_out_19_1_0, 
      que_out_19_2_15, que_out_19_2_14, que_out_19_2_13, que_out_19_2_12, 
      que_out_19_2_11, que_out_19_2_10, que_out_19_2_9, que_out_19_2_8, 
      que_out_19_2_7, que_out_19_2_6, que_out_19_2_5, que_out_19_2_4, 
      que_out_19_2_3, que_out_19_2_2, que_out_19_2_1, que_out_19_2_0, 
      que_out_19_3_15, que_out_19_3_14, que_out_19_3_13, que_out_19_3_12, 
      que_out_19_3_11, que_out_19_3_10, que_out_19_3_9, que_out_19_3_8, 
      que_out_19_3_7, que_out_19_3_6, que_out_19_3_5, que_out_19_3_4, 
      que_out_19_3_3, que_out_19_3_2, que_out_19_3_1, que_out_19_3_0, 
      que_out_19_4_15, que_out_19_4_14, que_out_19_4_13, que_out_19_4_12, 
      que_out_19_4_11, que_out_19_4_10, que_out_19_4_9, que_out_19_4_8, 
      que_out_19_4_7, que_out_19_4_6, que_out_19_4_5, que_out_19_4_4, 
      que_out_19_4_3, que_out_19_4_2, que_out_19_4_1, que_out_19_4_0, 
      que_out_20_0_15, que_out_20_0_14, que_out_20_0_13, que_out_20_0_12, 
      que_out_20_0_11, que_out_20_0_10, que_out_20_0_9, que_out_20_0_8, 
      que_out_20_0_7, que_out_20_0_6, que_out_20_0_5, que_out_20_0_4, 
      que_out_20_0_3, que_out_20_0_2, que_out_20_0_1, que_out_20_0_0, 
      que_out_20_1_15, que_out_20_1_14, que_out_20_1_13, que_out_20_1_12, 
      que_out_20_1_11, que_out_20_1_10, que_out_20_1_9, que_out_20_1_8, 
      que_out_20_1_7, que_out_20_1_6, que_out_20_1_5, que_out_20_1_4, 
      que_out_20_1_3, que_out_20_1_2, que_out_20_1_1, que_out_20_1_0, 
      que_out_20_2_15, que_out_20_2_14, que_out_20_2_13, que_out_20_2_12, 
      que_out_20_2_11, que_out_20_2_10, que_out_20_2_9, que_out_20_2_8, 
      que_out_20_2_7, que_out_20_2_6, que_out_20_2_5, que_out_20_2_4, 
      que_out_20_2_3, que_out_20_2_2, que_out_20_2_1, que_out_20_2_0, 
      que_out_20_3_15, que_out_20_3_14, que_out_20_3_13, que_out_20_3_12, 
      que_out_20_3_11, que_out_20_3_10, que_out_20_3_9, que_out_20_3_8, 
      que_out_20_3_7, que_out_20_3_6, que_out_20_3_5, que_out_20_3_4, 
      que_out_20_3_3, que_out_20_3_2, que_out_20_3_1, que_out_20_3_0, 
      que_out_20_4_15, que_out_20_4_14, que_out_20_4_13, que_out_20_4_12, 
      que_out_20_4_11, que_out_20_4_10, que_out_20_4_9, que_out_20_4_8, 
      que_out_20_4_7, que_out_20_4_6, que_out_20_4_5, que_out_20_4_4, 
      que_out_20_4_3, que_out_20_4_2, que_out_20_4_1, que_out_20_4_0, 
      que_out_21_0_15, que_out_21_0_14, que_out_21_0_13, que_out_21_0_12, 
      que_out_21_0_11, que_out_21_0_10, que_out_21_0_9, que_out_21_0_8, 
      que_out_21_0_7, que_out_21_0_6, que_out_21_0_5, que_out_21_0_4, 
      que_out_21_0_3, que_out_21_0_2, que_out_21_0_1, que_out_21_0_0, 
      que_out_21_1_15, que_out_21_1_14, que_out_21_1_13, que_out_21_1_12, 
      que_out_21_1_11, que_out_21_1_10, que_out_21_1_9, que_out_21_1_8, 
      que_out_21_1_7, que_out_21_1_6, que_out_21_1_5, que_out_21_1_4, 
      que_out_21_1_3, que_out_21_1_2, que_out_21_1_1, que_out_21_1_0, 
      que_out_21_2_15, que_out_21_2_14, que_out_21_2_13, que_out_21_2_12, 
      que_out_21_2_11, que_out_21_2_10, que_out_21_2_9, que_out_21_2_8, 
      que_out_21_2_7, que_out_21_2_6, que_out_21_2_5, que_out_21_2_4, 
      que_out_21_2_3, que_out_21_2_2, que_out_21_2_1, que_out_21_2_0, 
      que_out_21_3_15, que_out_21_3_14, que_out_21_3_13, que_out_21_3_12, 
      que_out_21_3_11, que_out_21_3_10, que_out_21_3_9, que_out_21_3_8, 
      que_out_21_3_7, que_out_21_3_6, que_out_21_3_5, que_out_21_3_4, 
      que_out_21_3_3, que_out_21_3_2, que_out_21_3_1, que_out_21_3_0, 
      que_out_21_4_15, que_out_21_4_14, que_out_21_4_13, que_out_21_4_12, 
      que_out_21_4_11, que_out_21_4_10, que_out_21_4_9, que_out_21_4_8, 
      que_out_21_4_7, que_out_21_4_6, que_out_21_4_5, que_out_21_4_4, 
      que_out_21_4_3, que_out_21_4_2, que_out_21_4_1, que_out_21_4_0, 
      que_out_22_0_15, que_out_22_0_14, que_out_22_0_13, que_out_22_0_12, 
      que_out_22_0_11, que_out_22_0_10, que_out_22_0_9, que_out_22_0_8, 
      que_out_22_0_7, que_out_22_0_6, que_out_22_0_5, que_out_22_0_4, 
      que_out_22_0_3, que_out_22_0_2, que_out_22_0_1, que_out_22_0_0, 
      que_out_22_1_15, que_out_22_1_14, que_out_22_1_13, que_out_22_1_12, 
      que_out_22_1_11, que_out_22_1_10, que_out_22_1_9, que_out_22_1_8, 
      que_out_22_1_7, que_out_22_1_6, que_out_22_1_5, que_out_22_1_4, 
      que_out_22_1_3, que_out_22_1_2, que_out_22_1_1, que_out_22_1_0, 
      que_out_22_2_15, que_out_22_2_14, que_out_22_2_13, que_out_22_2_12, 
      que_out_22_2_11, que_out_22_2_10, que_out_22_2_9, que_out_22_2_8, 
      que_out_22_2_7, que_out_22_2_6, que_out_22_2_5, que_out_22_2_4, 
      que_out_22_2_3, que_out_22_2_2, que_out_22_2_1, que_out_22_2_0, 
      que_out_22_3_15, que_out_22_3_14, que_out_22_3_13, que_out_22_3_12, 
      que_out_22_3_11, que_out_22_3_10, que_out_22_3_9, que_out_22_3_8, 
      que_out_22_3_7, que_out_22_3_6, que_out_22_3_5, que_out_22_3_4, 
      que_out_22_3_3, que_out_22_3_2, que_out_22_3_1, que_out_22_3_0, 
      que_out_22_4_15, que_out_22_4_14, que_out_22_4_13, que_out_22_4_12, 
      que_out_22_4_11, que_out_22_4_10, que_out_22_4_9, que_out_22_4_8, 
      que_out_22_4_7, que_out_22_4_6, que_out_22_4_5, que_out_22_4_4, 
      que_out_22_4_3, que_out_22_4_2, que_out_22_4_1, que_out_22_4_0, 
      que_out_23_0_15, que_out_23_0_14, que_out_23_0_13, que_out_23_0_12, 
      que_out_23_0_11, que_out_23_0_10, que_out_23_0_9, que_out_23_0_8, 
      que_out_23_0_7, que_out_23_0_6, que_out_23_0_5, que_out_23_0_4, 
      que_out_23_0_3, que_out_23_0_2, que_out_23_0_1, que_out_23_0_0, 
      que_out_23_1_15, que_out_23_1_14, que_out_23_1_13, que_out_23_1_12, 
      que_out_23_1_11, que_out_23_1_10, que_out_23_1_9, que_out_23_1_8, 
      que_out_23_1_7, que_out_23_1_6, que_out_23_1_5, que_out_23_1_4, 
      que_out_23_1_3, que_out_23_1_2, que_out_23_1_1, que_out_23_1_0, 
      que_out_23_2_15, que_out_23_2_14, que_out_23_2_13, que_out_23_2_12, 
      que_out_23_2_11, que_out_23_2_10, que_out_23_2_9, que_out_23_2_8, 
      que_out_23_2_7, que_out_23_2_6, que_out_23_2_5, que_out_23_2_4, 
      que_out_23_2_3, que_out_23_2_2, que_out_23_2_1, que_out_23_2_0, 
      que_out_23_3_15, que_out_23_3_14, que_out_23_3_13, que_out_23_3_12, 
      que_out_23_3_11, que_out_23_3_10, que_out_23_3_9, que_out_23_3_8, 
      que_out_23_3_7, que_out_23_3_6, que_out_23_3_5, que_out_23_3_4, 
      que_out_23_3_3, que_out_23_3_2, que_out_23_3_1, que_out_23_3_0, 
      que_out_23_4_15, que_out_23_4_14, que_out_23_4_13, que_out_23_4_12, 
      que_out_23_4_11, que_out_23_4_10, que_out_23_4_9, que_out_23_4_8, 
      que_out_23_4_7, que_out_23_4_6, que_out_23_4_5, que_out_23_4_4, 
      que_out_23_4_3, que_out_23_4_2, que_out_23_4_1, que_out_23_4_0, 
      que_out_24_0_15, que_out_24_0_14, que_out_24_0_13, que_out_24_0_12, 
      que_out_24_0_11, que_out_24_0_10, que_out_24_0_9, que_out_24_0_8, 
      que_out_24_0_7, que_out_24_0_6, que_out_24_0_5, que_out_24_0_4, 
      que_out_24_0_3, que_out_24_0_2, que_out_24_0_1, que_out_24_0_0, 
      que_out_24_1_15, que_out_24_1_14, que_out_24_1_13, que_out_24_1_12, 
      que_out_24_1_11, que_out_24_1_10, que_out_24_1_9, que_out_24_1_8, 
      que_out_24_1_7, que_out_24_1_6, que_out_24_1_5, que_out_24_1_4, 
      que_out_24_1_3, que_out_24_1_2, que_out_24_1_1, que_out_24_1_0, 
      que_out_24_2_15, que_out_24_2_14, que_out_24_2_13, que_out_24_2_12, 
      que_out_24_2_11, que_out_24_2_10, que_out_24_2_9, que_out_24_2_8, 
      que_out_24_2_7, que_out_24_2_6, que_out_24_2_5, que_out_24_2_4, 
      que_out_24_2_3, que_out_24_2_2, que_out_24_2_1, que_out_24_2_0, 
      que_out_24_3_15, que_out_24_3_14, que_out_24_3_13, que_out_24_3_12, 
      que_out_24_3_11, que_out_24_3_10, que_out_24_3_9, que_out_24_3_8, 
      que_out_24_3_7, que_out_24_3_6, que_out_24_3_5, que_out_24_3_4, 
      que_out_24_3_3, que_out_24_3_2, que_out_24_3_1, que_out_24_3_0, 
      que_out_24_4_15, que_out_24_4_14, que_out_24_4_13, que_out_24_4_12, 
      que_out_24_4_11, que_out_24_4_10, que_out_24_4_9, que_out_24_4_8, 
      que_out_24_4_7, que_out_24_4_6, que_out_24_4_5, que_out_24_4_4, 
      que_out_24_4_3, que_out_24_4_2, que_out_24_4_1, que_out_24_4_0, 
      que_out_25_0_15, que_out_25_0_14, que_out_25_0_13, que_out_25_0_12, 
      que_out_25_0_11, que_out_25_0_10, que_out_25_0_9, que_out_25_0_8, 
      que_out_25_0_7, que_out_25_0_6, que_out_25_0_5, que_out_25_0_4, 
      que_out_25_0_3, que_out_25_0_2, que_out_25_0_1, que_out_25_0_0, 
      que_out_25_1_15, que_out_25_1_14, que_out_25_1_13, que_out_25_1_12, 
      que_out_25_1_11, que_out_25_1_10, que_out_25_1_9, que_out_25_1_8, 
      que_out_25_1_7, que_out_25_1_6, que_out_25_1_5, que_out_25_1_4, 
      que_out_25_1_3, que_out_25_1_2, que_out_25_1_1, que_out_25_1_0, 
      que_out_25_2_15, que_out_25_2_14, que_out_25_2_13, que_out_25_2_12, 
      que_out_25_2_11, que_out_25_2_10, que_out_25_2_9, que_out_25_2_8, 
      que_out_25_2_7, que_out_25_2_6, que_out_25_2_5, que_out_25_2_4, 
      que_out_25_2_3, que_out_25_2_2, que_out_25_2_1, que_out_25_2_0, 
      que_out_25_3_15, que_out_25_3_14, que_out_25_3_13, que_out_25_3_12, 
      que_out_25_3_11, que_out_25_3_10, que_out_25_3_9, que_out_25_3_8, 
      que_out_25_3_7, que_out_25_3_6, que_out_25_3_5, que_out_25_3_4, 
      que_out_25_3_3, que_out_25_3_2, que_out_25_3_1, que_out_25_3_0, 
      que_out_25_4_15, que_out_25_4_14, que_out_25_4_13, que_out_25_4_12, 
      que_out_25_4_11, que_out_25_4_10, que_out_25_4_9, que_out_25_4_8, 
      que_out_25_4_7, que_out_25_4_6, que_out_25_4_5, que_out_25_4_4, 
      que_out_25_4_3, que_out_25_4_2, que_out_25_4_1, que_out_25_4_0, 
      que_out_26_0_15, que_out_26_0_14, que_out_26_0_13, que_out_26_0_12, 
      que_out_26_0_11, que_out_26_0_10, que_out_26_0_9, que_out_26_0_8, 
      que_out_26_0_7, que_out_26_0_6, que_out_26_0_5, que_out_26_0_4, 
      que_out_26_0_3, que_out_26_0_2, que_out_26_0_1, que_out_26_0_0, 
      que_out_26_1_15, que_out_26_1_14, que_out_26_1_13, que_out_26_1_12, 
      que_out_26_1_11, que_out_26_1_10, que_out_26_1_9, que_out_26_1_8, 
      que_out_26_1_7, que_out_26_1_6, que_out_26_1_5, que_out_26_1_4, 
      que_out_26_1_3, que_out_26_1_2, que_out_26_1_1, que_out_26_1_0, 
      que_out_26_2_15, que_out_26_2_14, que_out_26_2_13, que_out_26_2_12, 
      que_out_26_2_11, que_out_26_2_10, que_out_26_2_9, que_out_26_2_8, 
      que_out_26_2_7, que_out_26_2_6, que_out_26_2_5, que_out_26_2_4, 
      que_out_26_2_3, que_out_26_2_2, que_out_26_2_1, que_out_26_2_0, 
      que_out_26_3_15, que_out_26_3_14, que_out_26_3_13, que_out_26_3_12, 
      que_out_26_3_11, que_out_26_3_10, que_out_26_3_9, que_out_26_3_8, 
      que_out_26_3_7, que_out_26_3_6, que_out_26_3_5, que_out_26_3_4, 
      que_out_26_3_3, que_out_26_3_2, que_out_26_3_1, que_out_26_3_0, 
      que_out_26_4_15, que_out_26_4_14, que_out_26_4_13, que_out_26_4_12, 
      que_out_26_4_11, que_out_26_4_10, que_out_26_4_9, que_out_26_4_8, 
      que_out_26_4_7, que_out_26_4_6, que_out_26_4_5, que_out_26_4_4, 
      que_out_26_4_3, que_out_26_4_2, que_out_26_4_1, que_out_26_4_0, 
      que_out_27_0_15, que_out_27_0_14, que_out_27_0_13, que_out_27_0_12, 
      que_out_27_0_11, que_out_27_0_10, que_out_27_0_9, que_out_27_0_8, 
      que_out_27_0_7, que_out_27_0_6, que_out_27_0_5, que_out_27_0_4, 
      que_out_27_0_3, que_out_27_0_2, que_out_27_0_1, que_out_27_0_0, 
      que_out_27_1_15, que_out_27_1_14, que_out_27_1_13, que_out_27_1_12, 
      que_out_27_1_11, que_out_27_1_10, que_out_27_1_9, que_out_27_1_8, 
      que_out_27_1_7, que_out_27_1_6, que_out_27_1_5, que_out_27_1_4, 
      que_out_27_1_3, que_out_27_1_2, que_out_27_1_1, que_out_27_1_0, 
      que_out_27_2_15, que_out_27_2_14, que_out_27_2_13, que_out_27_2_12, 
      que_out_27_2_11, que_out_27_2_10, que_out_27_2_9, que_out_27_2_8, 
      que_out_27_2_7, que_out_27_2_6, que_out_27_2_5, que_out_27_2_4, 
      que_out_27_2_3, que_out_27_2_2, que_out_27_2_1, que_out_27_2_0, 
      que_out_27_3_15, que_out_27_3_14, que_out_27_3_13, que_out_27_3_12, 
      que_out_27_3_11, que_out_27_3_10, que_out_27_3_9, que_out_27_3_8, 
      que_out_27_3_7, que_out_27_3_6, que_out_27_3_5, que_out_27_3_4, 
      que_out_27_3_3, que_out_27_3_2, que_out_27_3_1, que_out_27_3_0, 
      que_out_27_4_15, que_out_27_4_14, que_out_27_4_13, que_out_27_4_12, 
      que_out_27_4_11, que_out_27_4_10, que_out_27_4_9, que_out_27_4_8, 
      que_out_27_4_7, que_out_27_4_6, que_out_27_4_5, que_out_27_4_4, 
      que_out_27_4_3, que_out_27_4_2, que_out_27_4_1, que_out_27_4_0, 
      sel_que_27, sel_que_26, sel_que_25, sel_que_24, sel_que_23, sel_que_22, 
      sel_que_21, sel_que_20, sel_que_19, sel_que_18, sel_que_17, sel_que_16, 
      sel_que_15, sel_que_14, sel_que_13, sel_que_12, sel_que_11, sel_que_10, 
      sel_que_9, sel_que_8, sel_que_7, sel_que_6, sel_que_5, sel_que_4, 
      sel_que_3, sel_que_2, sel_que_1, sel_que_0, nx12, nx14, nx28, nx30, 
      nx42, nx48, nx62, nx64, nx68, nx74, nx82, nx88, nx90, nx94, nx100, 
      nx104, nx114, nx118, nx122, nx130, nx136, nx144, nx150, nx158, nx166, 
      nx172, nx180, nx188, nx192, nx200, nx206, nx214, nx222, nx226, nx230, 
      nx238, nx268, nx294, nx322, nx348, nx378, nx404, nx432, nx458, nx488, 
      nx514, nx542, nx568, nx598, nx624, nx652, nx678, nx708, nx734, nx762, 
      nx788, nx818, nx844, nx872, nx898, nx928, nx954, nx982, nx1008, nx1038, 
      nx1064, nx1092, nx1118, nx1148, nx1174, nx1202, nx1228, nx1258, nx1284, 
      nx1312, nx1338, nx1368, nx1394, nx1422, nx1448, nx1478, nx1504, nx1532, 
      nx1558, nx1588, nx1614, nx1642, nx1668, nx1698, nx1724, nx1752, nx1778, 
      nx1808, nx1834, nx1862, nx1888, nx1918, nx1944, nx1972, nx1998, nx2028, 
      nx2054, nx2082, nx2108, nx2138, nx2164, nx2192, nx2218, nx2248, nx2274, 
      nx2302, nx2328, nx2358, nx2384, nx2412, nx2438, nx2468, nx2494, nx2522, 
      nx2548, nx2578, nx2604, nx2632, nx2658, nx2688, nx2714, nx2742, nx2768, 
      nx2798, nx2824, nx2852, nx2878, nx2908, nx2934, nx2962, nx2988, nx3018, 
      nx3044, nx3072, nx3098, nx3128, nx3154, nx3182, nx3208, nx3238, nx3264, 
      nx3292, nx3318, nx3348, nx3374, nx3402, nx3428, nx3458, nx3484, nx3512, 
      nx3538, nx3568, nx3594, nx3622, nx3648, nx3678, nx3704, nx3732, nx3758, 
      nx3788, nx3814, nx3842, nx3868, nx3898, nx3924, nx3952, nx3978, nx4008, 
      nx4034, nx4062, nx4088, nx4118, nx4144, nx4172, nx4198, nx4228, nx4254, 
      nx4282, nx4308, nx4338, nx4364, nx4392, nx4418, nx4448, nx4474, nx4502, 
      nx4528, nx4558, nx4584, nx4612, nx4638, nx4668, nx4694, nx4722, nx4748, 
      nx4778, nx4804, nx4832, nx4858, nx4888, nx4914, nx4942, nx4968, nx4998, 
      nx5024, nx5052, nx5078, nx5108, nx5134, nx5162, nx5188, nx5218, nx5244, 
      nx5272, nx5298, nx5328, nx5354, nx5382, nx5408, nx5438, nx5464, nx5492, 
      nx5518, nx5548, nx5574, nx5602, nx5628, nx5658, nx5684, nx5712, nx5738, 
      nx5768, nx5794, nx5822, nx5848, nx5878, nx5904, nx5932, nx5958, nx5988, 
      nx6014, nx6042, nx6068, nx6098, nx6124, nx6152, nx6178, nx6208, nx6234, 
      nx6262, nx6288, nx6318, nx6344, nx6372, nx6398, nx6428, nx6454, nx6482, 
      nx6508, nx6538, nx6564, nx6592, nx6618, nx6648, nx6674, nx6702, nx6728, 
      nx6758, nx6784, nx6812, nx6838, nx6868, nx6894, nx6922, nx6948, nx6978, 
      nx7004, nx7032, nx7058, nx7088, nx7114, nx7142, nx7168, nx7198, nx7224, 
      nx7252, nx7278, nx7308, nx7334, nx7362, nx7388, nx7418, nx7444, nx7472, 
      nx7498, nx7528, nx7554, nx7582, nx7608, nx7638, nx7664, nx7692, nx7718, 
      nx7748, nx7774, nx7802, nx7828, nx7858, nx7884, nx7912, nx7938, nx7968, 
      nx7994, nx8022, nx8048, nx8078, nx8104, nx8132, nx8158, nx8188, nx8214, 
      nx8242, nx8268, nx8298, nx8324, nx8352, nx8378, nx8408, nx8434, nx8462, 
      nx8488, nx8518, nx8544, nx8572, nx8598, nx8628, nx8654, nx8682, nx8708, 
      nx8738, nx8764, nx8792, nx8818, nx8848, nx8874, nx8902, nx8928, nx8938, 
      nx9038, nx6829, nx6833, nx6835, nx6839, nx6843, nx6847, nx6875, nx6885, 
      nx6889, nx6893, nx6897, nx6901, nx6905, nx6915, nx6927, nx6931, nx6933, 
      nx6937, nx6939, nx6943, nx6945, nx6949, nx6951, nx6955, nx6957, nx6961, 
      nx6965, nx6967, nx6971, nx6977, nx6985, nx6991, nx6999, nx7007, nx7017, 
      nx7029, nx7037, nx7043, nx7053, nx7055, nx7057, nx7061, nx7063, nx7065, 
      nx7069, nx7071, nx7073, nx7077, nx7079, nx7081, nx7087, nx7089, nx7091, 
      nx7095, nx7097, nx7099, nx7103, nx7105, nx7107, nx7111, nx7113, nx7115, 
      nx7121, nx7123, nx7125, nx7129, nx7131, nx7133, nx7137, nx7139, nx7141, 
      nx7145, nx7147, nx7149, nx7155, nx7157, nx7159, nx7163, nx7165, nx7167, 
      nx7171, nx7173, nx7175, nx7179, nx7181, nx7183, nx7189, nx7191, nx7193, 
      nx7197, nx7199, nx7201, nx7205, nx7207, nx7209, nx7213, nx7215, nx7217, 
      nx7223, nx7225, nx7227, nx7231, nx7233, nx7235, nx7239, nx7241, nx7243, 
      nx7247, nx7249, nx7251, nx7257, nx7259, nx7261, nx7265, nx7267, nx7269, 
      nx7273, nx7275, nx7277, nx7281, nx7283, nx7285, nx7291, nx7293, nx7295, 
      nx7299, nx7301, nx7303, nx7307, nx7309, nx7311, nx7315, nx7317, nx7319, 
      nx7325, nx7327, nx7329, nx7333, nx7335, nx7337, nx7341, nx7343, nx7345, 
      nx7349, nx7351, nx7353, nx7359, nx7361, nx7363, nx7367, nx7369, nx7371, 
      nx7375, nx7377, nx7379, nx7383, nx7385, nx7387, nx7393, nx7395, nx7397, 
      nx7401, nx7403, nx7405, nx7409, nx7411, nx7413, nx7417, nx7419, nx7421, 
      nx7427, nx7429, nx7431, nx7435, nx7437, nx7439, nx7443, nx7445, nx7447, 
      nx7451, nx7453, nx7455, nx7461, nx7463, nx7465, nx7469, nx7471, nx7473, 
      nx7477, nx7479, nx7481, nx7485, nx7487, nx7489, nx7495, nx7497, nx7499, 
      nx7503, nx7505, nx7507, nx7511, nx7513, nx7515, nx7519, nx7521, nx7523, 
      nx7529, nx7531, nx7533, nx7537, nx7539, nx7541, nx7545, nx7547, nx7549, 
      nx7553, nx7555, nx7557, nx7563, nx7565, nx7567, nx7571, nx7573, nx7575, 
      nx7579, nx7581, nx7583, nx7587, nx7589, nx7591, nx7597, nx7599, nx7601, 
      nx7605, nx7607, nx7609, nx7613, nx7615, nx7617, nx7621, nx7623, nx7625, 
      nx7631, nx7633, nx7635, nx7639, nx7641, nx7643, nx7647, nx7649, nx7651, 
      nx7655, nx7657, nx7659, nx7665, nx7667, nx7669, nx7673, nx7675, nx7677, 
      nx7681, nx7683, nx7685, nx7689, nx7691, nx7693, nx7699, nx7701, nx7703, 
      nx7707, nx7709, nx7711, nx7715, nx7717, nx7719, nx7723, nx7725, nx7727, 
      nx7733, nx7735, nx7737, nx7741, nx7743, nx7745, nx7749, nx7751, nx7753, 
      nx7757, nx7759, nx7761, nx7767, nx7769, nx7771, nx7775, nx7777, nx7779, 
      nx7783, nx7785, nx7787, nx7791, nx7793, nx7795, nx7801, nx7803, nx7805, 
      nx7809, nx7811, nx7813, nx7817, nx7819, nx7821, nx7825, nx7827, nx7829, 
      nx7835, nx7837, nx7839, nx7843, nx7845, nx7847, nx7851, nx7853, nx7855, 
      nx7859, nx7861, nx7863, nx7869, nx7871, nx7873, nx7877, nx7879, nx7881, 
      nx7885, nx7887, nx7889, nx7893, nx7895, nx7897, nx7903, nx7905, nx7907, 
      nx7911, nx7913, nx7915, nx7919, nx7921, nx7923, nx7927, nx7929, nx7931, 
      nx7937, nx7939, nx7941, nx7945, nx7947, nx7949, nx7953, nx7955, nx7957, 
      nx7961, nx7963, nx7965, nx7971, nx7973, nx7975, nx7979, nx7981, nx7983, 
      nx7987, nx7989, nx7991, nx7995, nx7997, nx7999, nx8005, nx8007, nx8009, 
      nx8013, nx8015, nx8017, nx8021, nx8023, nx8025, nx8029, nx8031, nx8033, 
      nx8039, nx8041, nx8043, nx8047, nx8049, nx8051, nx8055, nx8057, nx8059, 
      nx8063, nx8065, nx8067, nx8073, nx8075, nx8077, nx8081, nx8083, nx8085, 
      nx8089, nx8091, nx8093, nx8097, nx8099, nx8101, nx8107, nx8109, nx8111, 
      nx8115, nx8117, nx8119, nx8123, nx8125, nx8127, nx8131, nx8133, nx8135, 
      nx8141, nx8143, nx8145, nx8149, nx8151, nx8153, nx8157, nx8159, nx8161, 
      nx8165, nx8167, nx8169, nx8175, nx8177, nx8179, nx8183, nx8185, nx8187, 
      nx8191, nx8193, nx8195, nx8199, nx8201, nx8203, nx8209, nx8211, nx8213, 
      nx8217, nx8219, nx8221, nx8225, nx8227, nx8229, nx8233, nx8235, nx8237, 
      nx8243, nx8245, nx8247, nx8251, nx8253, nx8255, nx8259, nx8261, nx8263, 
      nx8267, nx8269, nx8271, nx8277, nx8279, nx8281, nx8285, nx8287, nx8289, 
      nx8293, nx8295, nx8297, nx8301, nx8303, nx8305, nx8311, nx8313, nx8315, 
      nx8319, nx8321, nx8323, nx8327, nx8329, nx8331, nx8335, nx8337, nx8339, 
      nx8345, nx8347, nx8349, nx8353, nx8355, nx8357, nx8361, nx8363, nx8365, 
      nx8369, nx8371, nx8373, nx8379, nx8381, nx8383, nx8387, nx8389, nx8391, 
      nx8395, nx8397, nx8399, nx8403, nx8405, nx8407, nx8413, nx8415, nx8417, 
      nx8421, nx8423, nx8425, nx8429, nx8431, nx8433, nx8437, nx8439, nx8441, 
      nx8447, nx8449, nx8451, nx8455, nx8457, nx8459, nx8463, nx8465, nx8467, 
      nx8471, nx8473, nx8475, nx8481, nx8483, nx8485, nx8489, nx8491, nx8493, 
      nx8497, nx8499, nx8501, nx8505, nx8507, nx8509, nx8515, nx8517, nx8519, 
      nx8523, nx8525, nx8527, nx8531, nx8533, nx8535, nx8539, nx8541, nx8543, 
      nx8549, nx8551, nx8553, nx8557, nx8559, nx8561, nx8565, nx8567, nx8569, 
      nx8573, nx8575, nx8577, nx8583, nx8585, nx8587, nx8591, nx8593, nx8595, 
      nx8599, nx8601, nx8603, nx8607, nx8609, nx8611, nx8617, nx8619, nx8621, 
      nx8625, nx8627, nx8629, nx8633, nx8635, nx8637, nx8641, nx8643, nx8645, 
      nx8651, nx8653, nx8655, nx8659, nx8661, nx8663, nx8667, nx8669, nx8671, 
      nx8675, nx8677, nx8679, nx8685, nx8687, nx8689, nx8693, nx8695, nx8697, 
      nx8701, nx8703, nx8705, nx8709, nx8711, nx8713, nx8719, nx8721, nx8723, 
      nx8727, nx8729, nx8731, nx8735, nx8737, nx8739, nx8743, nx8745, nx8747, 
      nx8753, nx8755, nx8757, nx8761, nx8763, nx8765, nx8769, nx8771, nx8773, 
      nx8777, nx8779, nx8781, nx8787, nx8789, nx8791, nx8795, nx8797, nx8799, 
      nx8803, nx8805, nx8807, nx8811, nx8813, nx8815, nx8821, nx8823, nx8825, 
      nx8829, nx8831, nx8833, nx8837, nx8839, nx8841, nx8845, nx8847, nx8849, 
      nx8855, nx8857, nx8859, nx8863, nx8865, nx8867, nx8871, nx8873, nx8875, 
      nx8879, nx8881, nx8883, nx8889, nx8891, nx8893, nx8897, nx8899, nx8901, 
      nx8905, nx8907, nx8909, nx8913, nx8915, nx8917, nx8923, nx8925, nx8927, 
      nx8931, nx8933, nx8935, nx8939, nx8941, nx8943, nx8947, nx8949, nx8951, 
      nx8955, nx8957, nx8959, nx8963, nx8965, nx8967, nx8970, nx8973, nx8975, 
      nx8978, nx8981, nx8983, nx8989, nx8991, nx8993, nx8997, nx8999, nx9001, 
      nx9005, nx9007, nx9009, nx9013, nx9015, nx9017, nx9023, nx9025, nx9027, 
      nx9031, nx9033, nx9035, nx9039, nx9041, nx9043, nx9047, nx9049, nx9051, 
      nx9057, nx9059, nx9061, nx9065, nx9067, nx9069, nx9073, nx9075, nx9077, 
      nx9081, nx9083, nx9085, nx9090, nx9093, nx9095, nx9098, nx9101, nx9103, 
      nx9106, nx9108, nx9110, nx9113, nx9115, nx9117, nx9121, nx9123, nx9125, 
      nx9128, nx9130, nx9132, nx9135, nx9137, nx9139, nx9142, nx9144, nx9146, 
      nx9150, nx9152, nx9154, nx9157, nx9159, nx9161, nx9164, nx9166, nx9168, 
      nx9171, nx9173, nx9175, nx9179, nx9181, nx9183, nx9186, nx9188, nx9190, 
      nx9193, nx9195, nx9197, nx9200, nx9202, nx9204, nx9208, nx9210, nx9212, 
      nx9215, nx9217, nx9219, nx9222, nx9224, nx9226, nx9229, nx9231, nx9233, 
      nx9237, nx9239, nx9241, nx9244, nx9246, nx9248, nx9251, nx9253, nx9255, 
      nx9258, nx9260, nx9262, nx9266, nx9268, nx9270, nx9273, nx9275, nx9277, 
      nx9280, nx9282, nx9284, nx9287, nx9289, nx9291, nx9295, nx9297, nx9299, 
      nx9302, nx9304, nx9306, nx9309, nx9311, nx9313, nx9316, nx9318, nx9320, 
      nx9324, nx9326, nx9328, nx9331, nx9333, nx9335, nx9338, nx9340, nx9342, 
      nx9345, nx9347, nx9349, nx9353, nx9355, nx9357, nx9360, nx9362, nx9364, 
      nx9367, nx9369, nx9371, nx9374, nx9376, nx9378, nx9382, nx9384, nx9386, 
      nx9389, nx9391, nx9393, nx9396, nx9398, nx9400, nx9403, nx9405, nx9407, 
      nx9411, nx9413, nx9415, nx9418, nx9420, nx9422, nx9425, nx9427, nx9429, 
      nx9432, nx9434, nx9436, nx9440, nx9442, nx9444, nx9447, nx9449, nx9451, 
      nx9454, nx9456, nx9458, nx9461, nx9463, nx9465, nx9469, nx9471, nx9473, 
      nx9476, nx9478, nx9480, nx9483, nx9485, nx9487, nx9490, nx9492, nx9494, 
      nx9498, nx9500, nx9502, nx9505, nx9507, nx9509, nx9512, nx9514, nx9516, 
      nx9519, nx9521, nx9523, nx9527, nx9529, nx9531, nx9534, nx9536, nx9538, 
      nx9541, nx9543, nx9545, nx9548, nx9550, nx9552, nx9556, nx9558, nx9560, 
      nx9563, nx9565, nx9567, nx9570, nx9572, nx9574, nx9577, nx9579, nx9581, 
      nx9585, nx9587, nx9589, nx9592, nx9594, nx9596, nx9599, nx9601, nx9603, 
      nx9606, nx9608, nx9610, nx9614, nx9616, nx9618, nx9621, nx9623, nx9625, 
      nx9628, nx9630, nx9632, nx9635, nx9637, nx9639, nx9648, nx9650, nx9652, 
      nx9654, nx9656, nx9658, nx9660, nx9662, nx9664, nx9666, nx9668, nx9670, 
      nx9674, nx9676, nx9678, nx9680, nx9682, nx9684, nx9686, nx9688, nx9690, 
      nx9692, nx9694, nx9696, nx9700, nx9702, nx9704, nx9706, nx9708, nx9710, 
      nx9712, nx9714, nx9716, nx9718, nx9720, nx9722, nx9726, nx9728, nx9730, 
      nx9732, nx9734, nx9736, nx9738, nx9740, nx9742, nx9744, nx9746, nx9748, 
      nx9752, nx9754, nx9756, nx9758, nx9760, nx9762, nx9764, nx9766, nx9768, 
      nx9770, nx9772, nx9774, nx9778, nx9780, nx9782, nx9784, nx9786, nx9788, 
      nx9790, nx9792, nx9794, nx9796, nx9798, nx9800, nx9804, nx9806, nx9808, 
      nx9810, nx9812, nx9814, nx9816, nx9818, nx9820, nx9822, nx9824, nx9826, 
      nx9830, nx9832, nx9834, nx9836, nx9838, nx9840, nx9842, nx9844, nx9846, 
      nx9848, nx9850, nx9852, nx9856, nx9858, nx9860, nx9862, nx9864, nx9866, 
      nx9868, nx9870, nx9872, nx9874, nx9876, nx9878, nx9882, nx9884, nx9886, 
      nx9888, nx9890, nx9892, nx9894, nx9896, nx9898, nx9900, nx9902, nx9904, 
      nx9908, nx9910, nx9912, nx9914, nx9916, nx9918, nx9920, nx9922, nx9924, 
      nx9926, nx9928, nx9930, nx9934, nx9936, nx9938, nx9940, nx9942, nx9944, 
      nx9946, nx9948, nx9950, nx9952, nx9954, nx9956, nx9960, nx9962, nx9964, 
      nx9966, nx9968, nx9970, nx9972, nx9974, nx9976, nx9978, nx9980, nx9982, 
      nx9986, nx9988, nx9990, nx9992, nx9994, nx9996, nx9998, nx10000, 
      nx10002, nx10004, nx10006, nx10008, nx10012, nx10014, nx10016, nx10018, 
      nx10020, nx10022, nx10024, nx10026, nx10028, nx10030, nx10032, nx10034, 
      nx10038, nx10040, nx10042, nx10044, nx10046, nx10048, nx10050, nx10052, 
      nx10054, nx10056, nx10058, nx10060, nx10064, nx10066, nx10068, nx10070, 
      nx10072, nx10074, nx10076, nx10078, nx10080, nx10082, nx10084, nx10086, 
      nx10090, nx10092, nx10094, nx10096, nx10098, nx10100, nx10102, nx10104, 
      nx10106, nx10108, nx10110, nx10112, nx10116, nx10118, nx10120, nx10122, 
      nx10124, nx10126, nx10128, nx10130, nx10132, nx10134, nx10136, nx10138, 
      nx10142, nx10144, nx10146, nx10148, nx10150, nx10152, nx10154, nx10156, 
      nx10158, nx10160, nx10162, nx10164, nx10168, nx10170, nx10172, nx10174, 
      nx10176, nx10178, nx10180, nx10182, nx10184, nx10186, nx10188, nx10190, 
      nx10194, nx10196, nx10198, nx10200, nx10202, nx10204, nx10206, nx10208, 
      nx10210, nx10212, nx10214, nx10216, nx10220, nx10222, nx10224, nx10226, 
      nx10228, nx10230, nx10232, nx10234, nx10236, nx10238, nx10240, nx10242, 
      nx10246, nx10248, nx10250, nx10252, nx10254, nx10256, nx10258, nx10260, 
      nx10262, nx10264, nx10266, nx10268, nx10272, nx10274, nx10276, nx10278, 
      nx10280, nx10282, nx10284, nx10286, nx10288, nx10290, nx10292, nx10294, 
      nx10298, nx10300, nx10302, nx10304, nx10306, nx10308, nx10310, nx10312, 
      nx10314, nx10316, nx10318, nx10320, nx10324, nx10326, nx10328, nx10330, 
      nx10332, nx10334, nx10336, nx10338, nx10340, nx10342, nx10344, nx10346, 
      nx10350, nx10352, nx10354, nx10356, nx10358, nx10360, nx10362, nx10364, 
      nx10366, nx10368, nx10370, nx10372, nx10374, nx10376, nx10378, nx10380, 
      nx10382, nx10384, nx10386, nx10388, nx10390, nx10392, nx10394, nx10396, 
      nx10398, nx10400, nx10402, nx10404, nx10406, nx10408, nx10410, nx10412, 
      nx10414, nx10416, nx10418, nx10420, nx10422, nx10424, nx10426, nx10428, 
      nx10430, nx10432, nx10434, nx10436, nx10438, nx10440, nx10442, nx10444, 
      nx10446, nx10448, nx10450, nx10452, nx10454, nx10456, nx10458, nx10460, 
      nx10462, nx10464, nx10466, nx10468, nx10470, nx10472, nx10474, nx10476, 
      nx10478, nx10480, nx10482, nx10484, nx10486, nx10488, nx10494, nx10496, 
      nx10498, nx10500, nx10502, nx10504, nx10506, nx10508, nx10510, nx10512, 
      nx10514, nx10516, nx10518, nx10520, nx10522, nx10524, nx10526, nx10528, 
      nx10530, nx10532, nx10534, nx10536, nx10538, nx10540, nx10542, nx10544, 
      nx10546, nx10548, nx10550, nx10552, nx10554, nx10556, nx10558, nx10560, 
      nx10562, nx10564, nx10566, nx10568, nx10570, nx10572, nx10574, nx10576, 
      nx10578, nx10580, nx10582, nx10584, nx10586, nx10588, nx10590, nx10592, 
      nx10594, nx10596, nx10598, nx10600, nx10602, nx10604, nx10606, nx10608, 
      nx10610, nx10612, nx10614, nx10616, nx10618, nx10620, nx10622, nx10624, 
      nx10626, nx10628, nx10630, nx10632, nx10634, nx10636, nx10638, nx10640, 
      nx10642, nx10644, nx10646, nx10648, nx10650, nx10652, nx10654, nx10656, 
      nx10658, nx10660, nx10662, nx10664, nx10666, nx10668, nx10690, nx10692, 
      nx10694, nx10696, nx10698, nx10700, nx10702, nx10704, nx10706, nx10708, 
      nx10710, nx10712, nx10714, nx10716, nx10718, nx10720, nx10722, nx10724, 
      nx10726, nx10728, nx10730, nx10732, nx10734, nx10736, nx10742, nx10744, 
      nx10746, nx10748: std_logic ;

begin
   gen_queues_0_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_0_0_15, q_0_14=>que_out_0_0_14, q_0_13=>
      que_out_0_0_13, q_0_12=>que_out_0_0_12, q_0_11=>que_out_0_0_11, q_0_10
      =>que_out_0_0_10, q_0_9=>que_out_0_0_9, q_0_8=>que_out_0_0_8, q_0_7=>
      que_out_0_0_7, q_0_6=>que_out_0_0_6, q_0_5=>que_out_0_0_5, q_0_4=>
      que_out_0_0_4, q_0_3=>que_out_0_0_3, q_0_2=>que_out_0_0_2, q_0_1=>
      que_out_0_0_1, q_0_0=>que_out_0_0_0, q_1_15=>que_out_0_1_15, q_1_14=>
      que_out_0_1_14, q_1_13=>que_out_0_1_13, q_1_12=>que_out_0_1_12, q_1_11
      =>que_out_0_1_11, q_1_10=>que_out_0_1_10, q_1_9=>que_out_0_1_9, q_1_8
      =>que_out_0_1_8, q_1_7=>que_out_0_1_7, q_1_6=>que_out_0_1_6, q_1_5=>
      que_out_0_1_5, q_1_4=>que_out_0_1_4, q_1_3=>que_out_0_1_3, q_1_2=>
      que_out_0_1_2, q_1_1=>que_out_0_1_1, q_1_0=>que_out_0_1_0, q_2_15=>
      que_out_0_2_15, q_2_14=>que_out_0_2_14, q_2_13=>que_out_0_2_13, q_2_12
      =>que_out_0_2_12, q_2_11=>que_out_0_2_11, q_2_10=>que_out_0_2_10, 
      q_2_9=>que_out_0_2_9, q_2_8=>que_out_0_2_8, q_2_7=>que_out_0_2_7, 
      q_2_6=>que_out_0_2_6, q_2_5=>que_out_0_2_5, q_2_4=>que_out_0_2_4, 
      q_2_3=>que_out_0_2_3, q_2_2=>que_out_0_2_2, q_2_1=>que_out_0_2_1, 
      q_2_0=>que_out_0_2_0, q_3_15=>que_out_0_3_15, q_3_14=>que_out_0_3_14, 
      q_3_13=>que_out_0_3_13, q_3_12=>que_out_0_3_12, q_3_11=>que_out_0_3_11, 
      q_3_10=>que_out_0_3_10, q_3_9=>que_out_0_3_9, q_3_8=>que_out_0_3_8, 
      q_3_7=>que_out_0_3_7, q_3_6=>que_out_0_3_6, q_3_5=>que_out_0_3_5, 
      q_3_4=>que_out_0_3_4, q_3_3=>que_out_0_3_3, q_3_2=>que_out_0_3_2, 
      q_3_1=>que_out_0_3_1, q_3_0=>que_out_0_3_0, q_4_15=>que_out_0_4_15, 
      q_4_14=>que_out_0_4_14, q_4_13=>que_out_0_4_13, q_4_12=>que_out_0_4_12, 
      q_4_11=>que_out_0_4_11, q_4_10=>que_out_0_4_10, q_4_9=>que_out_0_4_9, 
      q_4_8=>que_out_0_4_8, q_4_7=>que_out_0_4_7, q_4_6=>que_out_0_4_6, 
      q_4_5=>que_out_0_4_5, q_4_4=>que_out_0_4_4, q_4_3=>que_out_0_4_3, 
      q_4_2=>que_out_0_4_2, q_4_1=>que_out_0_4_1, q_4_0=>que_out_0_4_0, clk
      =>nx10714, load=>sel_que_0, reset=>nx10690);
   gen_queues_1_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_1_0_15, q_0_14=>que_out_1_0_14, q_0_13=>
      que_out_1_0_13, q_0_12=>que_out_1_0_12, q_0_11=>que_out_1_0_11, q_0_10
      =>que_out_1_0_10, q_0_9=>que_out_1_0_9, q_0_8=>que_out_1_0_8, q_0_7=>
      que_out_1_0_7, q_0_6=>que_out_1_0_6, q_0_5=>que_out_1_0_5, q_0_4=>
      que_out_1_0_4, q_0_3=>que_out_1_0_3, q_0_2=>que_out_1_0_2, q_0_1=>
      que_out_1_0_1, q_0_0=>que_out_1_0_0, q_1_15=>que_out_1_1_15, q_1_14=>
      que_out_1_1_14, q_1_13=>que_out_1_1_13, q_1_12=>que_out_1_1_12, q_1_11
      =>que_out_1_1_11, q_1_10=>que_out_1_1_10, q_1_9=>que_out_1_1_9, q_1_8
      =>que_out_1_1_8, q_1_7=>que_out_1_1_7, q_1_6=>que_out_1_1_6, q_1_5=>
      que_out_1_1_5, q_1_4=>que_out_1_1_4, q_1_3=>que_out_1_1_3, q_1_2=>
      que_out_1_1_2, q_1_1=>que_out_1_1_1, q_1_0=>que_out_1_1_0, q_2_15=>
      que_out_1_2_15, q_2_14=>que_out_1_2_14, q_2_13=>que_out_1_2_13, q_2_12
      =>que_out_1_2_12, q_2_11=>que_out_1_2_11, q_2_10=>que_out_1_2_10, 
      q_2_9=>que_out_1_2_9, q_2_8=>que_out_1_2_8, q_2_7=>que_out_1_2_7, 
      q_2_6=>que_out_1_2_6, q_2_5=>que_out_1_2_5, q_2_4=>que_out_1_2_4, 
      q_2_3=>que_out_1_2_3, q_2_2=>que_out_1_2_2, q_2_1=>que_out_1_2_1, 
      q_2_0=>que_out_1_2_0, q_3_15=>que_out_1_3_15, q_3_14=>que_out_1_3_14, 
      q_3_13=>que_out_1_3_13, q_3_12=>que_out_1_3_12, q_3_11=>que_out_1_3_11, 
      q_3_10=>que_out_1_3_10, q_3_9=>que_out_1_3_9, q_3_8=>que_out_1_3_8, 
      q_3_7=>que_out_1_3_7, q_3_6=>que_out_1_3_6, q_3_5=>que_out_1_3_5, 
      q_3_4=>que_out_1_3_4, q_3_3=>que_out_1_3_3, q_3_2=>que_out_1_3_2, 
      q_3_1=>que_out_1_3_1, q_3_0=>que_out_1_3_0, q_4_15=>que_out_1_4_15, 
      q_4_14=>que_out_1_4_14, q_4_13=>que_out_1_4_13, q_4_12=>que_out_1_4_12, 
      q_4_11=>que_out_1_4_11, q_4_10=>que_out_1_4_10, q_4_9=>que_out_1_4_9, 
      q_4_8=>que_out_1_4_8, q_4_7=>que_out_1_4_7, q_4_6=>que_out_1_4_6, 
      q_4_5=>que_out_1_4_5, q_4_4=>que_out_1_4_4, q_4_3=>que_out_1_4_3, 
      q_4_2=>que_out_1_4_2, q_4_1=>que_out_1_4_1, q_4_0=>que_out_1_4_0, clk
      =>nx10714, load=>sel_que_1, reset=>nx10690);
   gen_queues_2_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_2_0_15, q_0_14=>que_out_2_0_14, q_0_13=>
      que_out_2_0_13, q_0_12=>que_out_2_0_12, q_0_11=>que_out_2_0_11, q_0_10
      =>que_out_2_0_10, q_0_9=>que_out_2_0_9, q_0_8=>que_out_2_0_8, q_0_7=>
      que_out_2_0_7, q_0_6=>que_out_2_0_6, q_0_5=>que_out_2_0_5, q_0_4=>
      que_out_2_0_4, q_0_3=>que_out_2_0_3, q_0_2=>que_out_2_0_2, q_0_1=>
      que_out_2_0_1, q_0_0=>que_out_2_0_0, q_1_15=>que_out_2_1_15, q_1_14=>
      que_out_2_1_14, q_1_13=>que_out_2_1_13, q_1_12=>que_out_2_1_12, q_1_11
      =>que_out_2_1_11, q_1_10=>que_out_2_1_10, q_1_9=>que_out_2_1_9, q_1_8
      =>que_out_2_1_8, q_1_7=>que_out_2_1_7, q_1_6=>que_out_2_1_6, q_1_5=>
      que_out_2_1_5, q_1_4=>que_out_2_1_4, q_1_3=>que_out_2_1_3, q_1_2=>
      que_out_2_1_2, q_1_1=>que_out_2_1_1, q_1_0=>que_out_2_1_0, q_2_15=>
      que_out_2_2_15, q_2_14=>que_out_2_2_14, q_2_13=>que_out_2_2_13, q_2_12
      =>que_out_2_2_12, q_2_11=>que_out_2_2_11, q_2_10=>que_out_2_2_10, 
      q_2_9=>que_out_2_2_9, q_2_8=>que_out_2_2_8, q_2_7=>que_out_2_2_7, 
      q_2_6=>que_out_2_2_6, q_2_5=>que_out_2_2_5, q_2_4=>que_out_2_2_4, 
      q_2_3=>que_out_2_2_3, q_2_2=>que_out_2_2_2, q_2_1=>que_out_2_2_1, 
      q_2_0=>que_out_2_2_0, q_3_15=>que_out_2_3_15, q_3_14=>que_out_2_3_14, 
      q_3_13=>que_out_2_3_13, q_3_12=>que_out_2_3_12, q_3_11=>que_out_2_3_11, 
      q_3_10=>que_out_2_3_10, q_3_9=>que_out_2_3_9, q_3_8=>que_out_2_3_8, 
      q_3_7=>que_out_2_3_7, q_3_6=>que_out_2_3_6, q_3_5=>que_out_2_3_5, 
      q_3_4=>que_out_2_3_4, q_3_3=>que_out_2_3_3, q_3_2=>que_out_2_3_2, 
      q_3_1=>que_out_2_3_1, q_3_0=>que_out_2_3_0, q_4_15=>que_out_2_4_15, 
      q_4_14=>que_out_2_4_14, q_4_13=>que_out_2_4_13, q_4_12=>que_out_2_4_12, 
      q_4_11=>que_out_2_4_11, q_4_10=>que_out_2_4_10, q_4_9=>que_out_2_4_9, 
      q_4_8=>que_out_2_4_8, q_4_7=>que_out_2_4_7, q_4_6=>que_out_2_4_6, 
      q_4_5=>que_out_2_4_5, q_4_4=>que_out_2_4_4, q_4_3=>que_out_2_4_3, 
      q_4_2=>que_out_2_4_2, q_4_1=>que_out_2_4_1, q_4_0=>que_out_2_4_0, clk
      =>nx10714, load=>sel_que_2, reset=>nx10690);
   gen_queues_3_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_3_0_15, q_0_14=>que_out_3_0_14, q_0_13=>
      que_out_3_0_13, q_0_12=>que_out_3_0_12, q_0_11=>que_out_3_0_11, q_0_10
      =>que_out_3_0_10, q_0_9=>que_out_3_0_9, q_0_8=>que_out_3_0_8, q_0_7=>
      que_out_3_0_7, q_0_6=>que_out_3_0_6, q_0_5=>que_out_3_0_5, q_0_4=>
      que_out_3_0_4, q_0_3=>que_out_3_0_3, q_0_2=>que_out_3_0_2, q_0_1=>
      que_out_3_0_1, q_0_0=>que_out_3_0_0, q_1_15=>que_out_3_1_15, q_1_14=>
      que_out_3_1_14, q_1_13=>que_out_3_1_13, q_1_12=>que_out_3_1_12, q_1_11
      =>que_out_3_1_11, q_1_10=>que_out_3_1_10, q_1_9=>que_out_3_1_9, q_1_8
      =>que_out_3_1_8, q_1_7=>que_out_3_1_7, q_1_6=>que_out_3_1_6, q_1_5=>
      que_out_3_1_5, q_1_4=>que_out_3_1_4, q_1_3=>que_out_3_1_3, q_1_2=>
      que_out_3_1_2, q_1_1=>que_out_3_1_1, q_1_0=>que_out_3_1_0, q_2_15=>
      que_out_3_2_15, q_2_14=>que_out_3_2_14, q_2_13=>que_out_3_2_13, q_2_12
      =>que_out_3_2_12, q_2_11=>que_out_3_2_11, q_2_10=>que_out_3_2_10, 
      q_2_9=>que_out_3_2_9, q_2_8=>que_out_3_2_8, q_2_7=>que_out_3_2_7, 
      q_2_6=>que_out_3_2_6, q_2_5=>que_out_3_2_5, q_2_4=>que_out_3_2_4, 
      q_2_3=>que_out_3_2_3, q_2_2=>que_out_3_2_2, q_2_1=>que_out_3_2_1, 
      q_2_0=>que_out_3_2_0, q_3_15=>que_out_3_3_15, q_3_14=>que_out_3_3_14, 
      q_3_13=>que_out_3_3_13, q_3_12=>que_out_3_3_12, q_3_11=>que_out_3_3_11, 
      q_3_10=>que_out_3_3_10, q_3_9=>que_out_3_3_9, q_3_8=>que_out_3_3_8, 
      q_3_7=>que_out_3_3_7, q_3_6=>que_out_3_3_6, q_3_5=>que_out_3_3_5, 
      q_3_4=>que_out_3_3_4, q_3_3=>que_out_3_3_3, q_3_2=>que_out_3_3_2, 
      q_3_1=>que_out_3_3_1, q_3_0=>que_out_3_3_0, q_4_15=>que_out_3_4_15, 
      q_4_14=>que_out_3_4_14, q_4_13=>que_out_3_4_13, q_4_12=>que_out_3_4_12, 
      q_4_11=>que_out_3_4_11, q_4_10=>que_out_3_4_10, q_4_9=>que_out_3_4_9, 
      q_4_8=>que_out_3_4_8, q_4_7=>que_out_3_4_7, q_4_6=>que_out_3_4_6, 
      q_4_5=>que_out_3_4_5, q_4_4=>que_out_3_4_4, q_4_3=>que_out_3_4_3, 
      q_4_2=>que_out_3_4_2, q_4_1=>que_out_3_4_1, q_4_0=>que_out_3_4_0, clk
      =>nx10716, load=>sel_que_3, reset=>nx10692);
   gen_queues_4_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_4_0_15, q_0_14=>que_out_4_0_14, q_0_13=>
      que_out_4_0_13, q_0_12=>que_out_4_0_12, q_0_11=>que_out_4_0_11, q_0_10
      =>que_out_4_0_10, q_0_9=>que_out_4_0_9, q_0_8=>que_out_4_0_8, q_0_7=>
      que_out_4_0_7, q_0_6=>que_out_4_0_6, q_0_5=>que_out_4_0_5, q_0_4=>
      que_out_4_0_4, q_0_3=>que_out_4_0_3, q_0_2=>que_out_4_0_2, q_0_1=>
      que_out_4_0_1, q_0_0=>que_out_4_0_0, q_1_15=>que_out_4_1_15, q_1_14=>
      que_out_4_1_14, q_1_13=>que_out_4_1_13, q_1_12=>que_out_4_1_12, q_1_11
      =>que_out_4_1_11, q_1_10=>que_out_4_1_10, q_1_9=>que_out_4_1_9, q_1_8
      =>que_out_4_1_8, q_1_7=>que_out_4_1_7, q_1_6=>que_out_4_1_6, q_1_5=>
      que_out_4_1_5, q_1_4=>que_out_4_1_4, q_1_3=>que_out_4_1_3, q_1_2=>
      que_out_4_1_2, q_1_1=>que_out_4_1_1, q_1_0=>que_out_4_1_0, q_2_15=>
      que_out_4_2_15, q_2_14=>que_out_4_2_14, q_2_13=>que_out_4_2_13, q_2_12
      =>que_out_4_2_12, q_2_11=>que_out_4_2_11, q_2_10=>que_out_4_2_10, 
      q_2_9=>que_out_4_2_9, q_2_8=>que_out_4_2_8, q_2_7=>que_out_4_2_7, 
      q_2_6=>que_out_4_2_6, q_2_5=>que_out_4_2_5, q_2_4=>que_out_4_2_4, 
      q_2_3=>que_out_4_2_3, q_2_2=>que_out_4_2_2, q_2_1=>que_out_4_2_1, 
      q_2_0=>que_out_4_2_0, q_3_15=>que_out_4_3_15, q_3_14=>que_out_4_3_14, 
      q_3_13=>que_out_4_3_13, q_3_12=>que_out_4_3_12, q_3_11=>que_out_4_3_11, 
      q_3_10=>que_out_4_3_10, q_3_9=>que_out_4_3_9, q_3_8=>que_out_4_3_8, 
      q_3_7=>que_out_4_3_7, q_3_6=>que_out_4_3_6, q_3_5=>que_out_4_3_5, 
      q_3_4=>que_out_4_3_4, q_3_3=>que_out_4_3_3, q_3_2=>que_out_4_3_2, 
      q_3_1=>que_out_4_3_1, q_3_0=>que_out_4_3_0, q_4_15=>que_out_4_4_15, 
      q_4_14=>que_out_4_4_14, q_4_13=>que_out_4_4_13, q_4_12=>que_out_4_4_12, 
      q_4_11=>que_out_4_4_11, q_4_10=>que_out_4_4_10, q_4_9=>que_out_4_4_9, 
      q_4_8=>que_out_4_4_8, q_4_7=>que_out_4_4_7, q_4_6=>que_out_4_4_6, 
      q_4_5=>que_out_4_4_5, q_4_4=>que_out_4_4_4, q_4_3=>que_out_4_4_3, 
      q_4_2=>que_out_4_4_2, q_4_1=>que_out_4_4_1, q_4_0=>que_out_4_4_0, clk
      =>nx10716, load=>sel_que_4, reset=>nx10692);
   gen_queues_5_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_5_0_15, q_0_14=>que_out_5_0_14, q_0_13=>
      que_out_5_0_13, q_0_12=>que_out_5_0_12, q_0_11=>que_out_5_0_11, q_0_10
      =>que_out_5_0_10, q_0_9=>que_out_5_0_9, q_0_8=>que_out_5_0_8, q_0_7=>
      que_out_5_0_7, q_0_6=>que_out_5_0_6, q_0_5=>que_out_5_0_5, q_0_4=>
      que_out_5_0_4, q_0_3=>que_out_5_0_3, q_0_2=>que_out_5_0_2, q_0_1=>
      que_out_5_0_1, q_0_0=>que_out_5_0_0, q_1_15=>que_out_5_1_15, q_1_14=>
      que_out_5_1_14, q_1_13=>que_out_5_1_13, q_1_12=>que_out_5_1_12, q_1_11
      =>que_out_5_1_11, q_1_10=>que_out_5_1_10, q_1_9=>que_out_5_1_9, q_1_8
      =>que_out_5_1_8, q_1_7=>que_out_5_1_7, q_1_6=>que_out_5_1_6, q_1_5=>
      que_out_5_1_5, q_1_4=>que_out_5_1_4, q_1_3=>que_out_5_1_3, q_1_2=>
      que_out_5_1_2, q_1_1=>que_out_5_1_1, q_1_0=>que_out_5_1_0, q_2_15=>
      que_out_5_2_15, q_2_14=>que_out_5_2_14, q_2_13=>que_out_5_2_13, q_2_12
      =>que_out_5_2_12, q_2_11=>que_out_5_2_11, q_2_10=>que_out_5_2_10, 
      q_2_9=>que_out_5_2_9, q_2_8=>que_out_5_2_8, q_2_7=>que_out_5_2_7, 
      q_2_6=>que_out_5_2_6, q_2_5=>que_out_5_2_5, q_2_4=>que_out_5_2_4, 
      q_2_3=>que_out_5_2_3, q_2_2=>que_out_5_2_2, q_2_1=>que_out_5_2_1, 
      q_2_0=>que_out_5_2_0, q_3_15=>que_out_5_3_15, q_3_14=>que_out_5_3_14, 
      q_3_13=>que_out_5_3_13, q_3_12=>que_out_5_3_12, q_3_11=>que_out_5_3_11, 
      q_3_10=>que_out_5_3_10, q_3_9=>que_out_5_3_9, q_3_8=>que_out_5_3_8, 
      q_3_7=>que_out_5_3_7, q_3_6=>que_out_5_3_6, q_3_5=>que_out_5_3_5, 
      q_3_4=>que_out_5_3_4, q_3_3=>que_out_5_3_3, q_3_2=>que_out_5_3_2, 
      q_3_1=>que_out_5_3_1, q_3_0=>que_out_5_3_0, q_4_15=>que_out_5_4_15, 
      q_4_14=>que_out_5_4_14, q_4_13=>que_out_5_4_13, q_4_12=>que_out_5_4_12, 
      q_4_11=>que_out_5_4_11, q_4_10=>que_out_5_4_10, q_4_9=>que_out_5_4_9, 
      q_4_8=>que_out_5_4_8, q_4_7=>que_out_5_4_7, q_4_6=>que_out_5_4_6, 
      q_4_5=>que_out_5_4_5, q_4_4=>que_out_5_4_4, q_4_3=>que_out_5_4_3, 
      q_4_2=>que_out_5_4_2, q_4_1=>que_out_5_4_1, q_4_0=>que_out_5_4_0, clk
      =>nx10716, load=>sel_que_5, reset=>nx10692);
   gen_queues_6_que : Queue_5 port map ( d(15)=>nx10512, d(14)=>nx10522, 
      d(13)=>nx10532, d(12)=>nx10542, d(11)=>nx10552, d(10)=>nx10562, d(9)=>
      nx10572, d(8)=>nx10582, d(7)=>nx10592, d(6)=>nx10602, d(5)=>nx10612, 
      d(4)=>nx10622, d(3)=>nx10632, d(2)=>nx10642, d(1)=>nx10652, d(0)=>
      nx10662, q_0_15=>que_out_6_0_15, q_0_14=>que_out_6_0_14, q_0_13=>
      que_out_6_0_13, q_0_12=>que_out_6_0_12, q_0_11=>que_out_6_0_11, q_0_10
      =>que_out_6_0_10, q_0_9=>que_out_6_0_9, q_0_8=>que_out_6_0_8, q_0_7=>
      que_out_6_0_7, q_0_6=>que_out_6_0_6, q_0_5=>que_out_6_0_5, q_0_4=>
      que_out_6_0_4, q_0_3=>que_out_6_0_3, q_0_2=>que_out_6_0_2, q_0_1=>
      que_out_6_0_1, q_0_0=>que_out_6_0_0, q_1_15=>que_out_6_1_15, q_1_14=>
      que_out_6_1_14, q_1_13=>que_out_6_1_13, q_1_12=>que_out_6_1_12, q_1_11
      =>que_out_6_1_11, q_1_10=>que_out_6_1_10, q_1_9=>que_out_6_1_9, q_1_8
      =>que_out_6_1_8, q_1_7=>que_out_6_1_7, q_1_6=>que_out_6_1_6, q_1_5=>
      que_out_6_1_5, q_1_4=>que_out_6_1_4, q_1_3=>que_out_6_1_3, q_1_2=>
      que_out_6_1_2, q_1_1=>que_out_6_1_1, q_1_0=>que_out_6_1_0, q_2_15=>
      que_out_6_2_15, q_2_14=>que_out_6_2_14, q_2_13=>que_out_6_2_13, q_2_12
      =>que_out_6_2_12, q_2_11=>que_out_6_2_11, q_2_10=>que_out_6_2_10, 
      q_2_9=>que_out_6_2_9, q_2_8=>que_out_6_2_8, q_2_7=>que_out_6_2_7, 
      q_2_6=>que_out_6_2_6, q_2_5=>que_out_6_2_5, q_2_4=>que_out_6_2_4, 
      q_2_3=>que_out_6_2_3, q_2_2=>que_out_6_2_2, q_2_1=>que_out_6_2_1, 
      q_2_0=>que_out_6_2_0, q_3_15=>que_out_6_3_15, q_3_14=>que_out_6_3_14, 
      q_3_13=>que_out_6_3_13, q_3_12=>que_out_6_3_12, q_3_11=>que_out_6_3_11, 
      q_3_10=>que_out_6_3_10, q_3_9=>que_out_6_3_9, q_3_8=>que_out_6_3_8, 
      q_3_7=>que_out_6_3_7, q_3_6=>que_out_6_3_6, q_3_5=>que_out_6_3_5, 
      q_3_4=>que_out_6_3_4, q_3_3=>que_out_6_3_3, q_3_2=>que_out_6_3_2, 
      q_3_1=>que_out_6_3_1, q_3_0=>que_out_6_3_0, q_4_15=>que_out_6_4_15, 
      q_4_14=>que_out_6_4_14, q_4_13=>que_out_6_4_13, q_4_12=>que_out_6_4_12, 
      q_4_11=>que_out_6_4_11, q_4_10=>que_out_6_4_10, q_4_9=>que_out_6_4_9, 
      q_4_8=>que_out_6_4_8, q_4_7=>que_out_6_4_7, q_4_6=>que_out_6_4_6, 
      q_4_5=>que_out_6_4_5, q_4_4=>que_out_6_4_4, q_4_3=>que_out_6_4_3, 
      q_4_2=>que_out_6_4_2, q_4_1=>que_out_6_4_1, q_4_0=>que_out_6_4_0, clk
      =>nx10718, load=>sel_que_6, reset=>nx10694);
   gen_queues_7_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_7_0_15, q_0_14=>que_out_7_0_14, q_0_13=>
      que_out_7_0_13, q_0_12=>que_out_7_0_12, q_0_11=>que_out_7_0_11, q_0_10
      =>que_out_7_0_10, q_0_9=>que_out_7_0_9, q_0_8=>que_out_7_0_8, q_0_7=>
      que_out_7_0_7, q_0_6=>que_out_7_0_6, q_0_5=>que_out_7_0_5, q_0_4=>
      que_out_7_0_4, q_0_3=>que_out_7_0_3, q_0_2=>que_out_7_0_2, q_0_1=>
      que_out_7_0_1, q_0_0=>que_out_7_0_0, q_1_15=>que_out_7_1_15, q_1_14=>
      que_out_7_1_14, q_1_13=>que_out_7_1_13, q_1_12=>que_out_7_1_12, q_1_11
      =>que_out_7_1_11, q_1_10=>que_out_7_1_10, q_1_9=>que_out_7_1_9, q_1_8
      =>que_out_7_1_8, q_1_7=>que_out_7_1_7, q_1_6=>que_out_7_1_6, q_1_5=>
      que_out_7_1_5, q_1_4=>que_out_7_1_4, q_1_3=>que_out_7_1_3, q_1_2=>
      que_out_7_1_2, q_1_1=>que_out_7_1_1, q_1_0=>que_out_7_1_0, q_2_15=>
      que_out_7_2_15, q_2_14=>que_out_7_2_14, q_2_13=>que_out_7_2_13, q_2_12
      =>que_out_7_2_12, q_2_11=>que_out_7_2_11, q_2_10=>que_out_7_2_10, 
      q_2_9=>que_out_7_2_9, q_2_8=>que_out_7_2_8, q_2_7=>que_out_7_2_7, 
      q_2_6=>que_out_7_2_6, q_2_5=>que_out_7_2_5, q_2_4=>que_out_7_2_4, 
      q_2_3=>que_out_7_2_3, q_2_2=>que_out_7_2_2, q_2_1=>que_out_7_2_1, 
      q_2_0=>que_out_7_2_0, q_3_15=>que_out_7_3_15, q_3_14=>que_out_7_3_14, 
      q_3_13=>que_out_7_3_13, q_3_12=>que_out_7_3_12, q_3_11=>que_out_7_3_11, 
      q_3_10=>que_out_7_3_10, q_3_9=>que_out_7_3_9, q_3_8=>que_out_7_3_8, 
      q_3_7=>que_out_7_3_7, q_3_6=>que_out_7_3_6, q_3_5=>que_out_7_3_5, 
      q_3_4=>que_out_7_3_4, q_3_3=>que_out_7_3_3, q_3_2=>que_out_7_3_2, 
      q_3_1=>que_out_7_3_1, q_3_0=>que_out_7_3_0, q_4_15=>que_out_7_4_15, 
      q_4_14=>que_out_7_4_14, q_4_13=>que_out_7_4_13, q_4_12=>que_out_7_4_12, 
      q_4_11=>que_out_7_4_11, q_4_10=>que_out_7_4_10, q_4_9=>que_out_7_4_9, 
      q_4_8=>que_out_7_4_8, q_4_7=>que_out_7_4_7, q_4_6=>que_out_7_4_6, 
      q_4_5=>que_out_7_4_5, q_4_4=>que_out_7_4_4, q_4_3=>que_out_7_4_3, 
      q_4_2=>que_out_7_4_2, q_4_1=>que_out_7_4_1, q_4_0=>que_out_7_4_0, clk
      =>nx10720, load=>sel_que_7, reset=>nx10696);
   gen_queues_8_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_8_0_15, q_0_14=>que_out_8_0_14, q_0_13=>
      que_out_8_0_13, q_0_12=>que_out_8_0_12, q_0_11=>que_out_8_0_11, q_0_10
      =>que_out_8_0_10, q_0_9=>que_out_8_0_9, q_0_8=>que_out_8_0_8, q_0_7=>
      que_out_8_0_7, q_0_6=>que_out_8_0_6, q_0_5=>que_out_8_0_5, q_0_4=>
      que_out_8_0_4, q_0_3=>que_out_8_0_3, q_0_2=>que_out_8_0_2, q_0_1=>
      que_out_8_0_1, q_0_0=>que_out_8_0_0, q_1_15=>que_out_8_1_15, q_1_14=>
      que_out_8_1_14, q_1_13=>que_out_8_1_13, q_1_12=>que_out_8_1_12, q_1_11
      =>que_out_8_1_11, q_1_10=>que_out_8_1_10, q_1_9=>que_out_8_1_9, q_1_8
      =>que_out_8_1_8, q_1_7=>que_out_8_1_7, q_1_6=>que_out_8_1_6, q_1_5=>
      que_out_8_1_5, q_1_4=>que_out_8_1_4, q_1_3=>que_out_8_1_3, q_1_2=>
      que_out_8_1_2, q_1_1=>que_out_8_1_1, q_1_0=>que_out_8_1_0, q_2_15=>
      que_out_8_2_15, q_2_14=>que_out_8_2_14, q_2_13=>que_out_8_2_13, q_2_12
      =>que_out_8_2_12, q_2_11=>que_out_8_2_11, q_2_10=>que_out_8_2_10, 
      q_2_9=>que_out_8_2_9, q_2_8=>que_out_8_2_8, q_2_7=>que_out_8_2_7, 
      q_2_6=>que_out_8_2_6, q_2_5=>que_out_8_2_5, q_2_4=>que_out_8_2_4, 
      q_2_3=>que_out_8_2_3, q_2_2=>que_out_8_2_2, q_2_1=>que_out_8_2_1, 
      q_2_0=>que_out_8_2_0, q_3_15=>que_out_8_3_15, q_3_14=>que_out_8_3_14, 
      q_3_13=>que_out_8_3_13, q_3_12=>que_out_8_3_12, q_3_11=>que_out_8_3_11, 
      q_3_10=>que_out_8_3_10, q_3_9=>que_out_8_3_9, q_3_8=>que_out_8_3_8, 
      q_3_7=>que_out_8_3_7, q_3_6=>que_out_8_3_6, q_3_5=>que_out_8_3_5, 
      q_3_4=>que_out_8_3_4, q_3_3=>que_out_8_3_3, q_3_2=>que_out_8_3_2, 
      q_3_1=>que_out_8_3_1, q_3_0=>que_out_8_3_0, q_4_15=>que_out_8_4_15, 
      q_4_14=>que_out_8_4_14, q_4_13=>que_out_8_4_13, q_4_12=>que_out_8_4_12, 
      q_4_11=>que_out_8_4_11, q_4_10=>que_out_8_4_10, q_4_9=>que_out_8_4_9, 
      q_4_8=>que_out_8_4_8, q_4_7=>que_out_8_4_7, q_4_6=>que_out_8_4_6, 
      q_4_5=>que_out_8_4_5, q_4_4=>que_out_8_4_4, q_4_3=>que_out_8_4_3, 
      q_4_2=>que_out_8_4_2, q_4_1=>que_out_8_4_1, q_4_0=>que_out_8_4_0, clk
      =>nx10720, load=>sel_que_8, reset=>nx10696);
   gen_queues_9_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_9_0_15, q_0_14=>que_out_9_0_14, q_0_13=>
      que_out_9_0_13, q_0_12=>que_out_9_0_12, q_0_11=>que_out_9_0_11, q_0_10
      =>que_out_9_0_10, q_0_9=>que_out_9_0_9, q_0_8=>que_out_9_0_8, q_0_7=>
      que_out_9_0_7, q_0_6=>que_out_9_0_6, q_0_5=>que_out_9_0_5, q_0_4=>
      que_out_9_0_4, q_0_3=>que_out_9_0_3, q_0_2=>que_out_9_0_2, q_0_1=>
      que_out_9_0_1, q_0_0=>que_out_9_0_0, q_1_15=>que_out_9_1_15, q_1_14=>
      que_out_9_1_14, q_1_13=>que_out_9_1_13, q_1_12=>que_out_9_1_12, q_1_11
      =>que_out_9_1_11, q_1_10=>que_out_9_1_10, q_1_9=>que_out_9_1_9, q_1_8
      =>que_out_9_1_8, q_1_7=>que_out_9_1_7, q_1_6=>que_out_9_1_6, q_1_5=>
      que_out_9_1_5, q_1_4=>que_out_9_1_4, q_1_3=>que_out_9_1_3, q_1_2=>
      que_out_9_1_2, q_1_1=>que_out_9_1_1, q_1_0=>que_out_9_1_0, q_2_15=>
      que_out_9_2_15, q_2_14=>que_out_9_2_14, q_2_13=>que_out_9_2_13, q_2_12
      =>que_out_9_2_12, q_2_11=>que_out_9_2_11, q_2_10=>que_out_9_2_10, 
      q_2_9=>que_out_9_2_9, q_2_8=>que_out_9_2_8, q_2_7=>que_out_9_2_7, 
      q_2_6=>que_out_9_2_6, q_2_5=>que_out_9_2_5, q_2_4=>que_out_9_2_4, 
      q_2_3=>que_out_9_2_3, q_2_2=>que_out_9_2_2, q_2_1=>que_out_9_2_1, 
      q_2_0=>que_out_9_2_0, q_3_15=>que_out_9_3_15, q_3_14=>que_out_9_3_14, 
      q_3_13=>que_out_9_3_13, q_3_12=>que_out_9_3_12, q_3_11=>que_out_9_3_11, 
      q_3_10=>que_out_9_3_10, q_3_9=>que_out_9_3_9, q_3_8=>que_out_9_3_8, 
      q_3_7=>que_out_9_3_7, q_3_6=>que_out_9_3_6, q_3_5=>que_out_9_3_5, 
      q_3_4=>que_out_9_3_4, q_3_3=>que_out_9_3_3, q_3_2=>que_out_9_3_2, 
      q_3_1=>que_out_9_3_1, q_3_0=>que_out_9_3_0, q_4_15=>que_out_9_4_15, 
      q_4_14=>que_out_9_4_14, q_4_13=>que_out_9_4_13, q_4_12=>que_out_9_4_12, 
      q_4_11=>que_out_9_4_11, q_4_10=>que_out_9_4_10, q_4_9=>que_out_9_4_9, 
      q_4_8=>que_out_9_4_8, q_4_7=>que_out_9_4_7, q_4_6=>que_out_9_4_6, 
      q_4_5=>que_out_9_4_5, q_4_4=>que_out_9_4_4, q_4_3=>que_out_9_4_3, 
      q_4_2=>que_out_9_4_2, q_4_1=>que_out_9_4_1, q_4_0=>que_out_9_4_0, clk
      =>nx10720, load=>sel_que_9, reset=>nx10696);
   gen_queues_10_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_10_0_15, q_0_14=>que_out_10_0_14, q_0_13=>
      que_out_10_0_13, q_0_12=>que_out_10_0_12, q_0_11=>que_out_10_0_11, 
      q_0_10=>que_out_10_0_10, q_0_9=>que_out_10_0_9, q_0_8=>que_out_10_0_8, 
      q_0_7=>que_out_10_0_7, q_0_6=>que_out_10_0_6, q_0_5=>que_out_10_0_5, 
      q_0_4=>que_out_10_0_4, q_0_3=>que_out_10_0_3, q_0_2=>que_out_10_0_2, 
      q_0_1=>que_out_10_0_1, q_0_0=>que_out_10_0_0, q_1_15=>que_out_10_1_15, 
      q_1_14=>que_out_10_1_14, q_1_13=>que_out_10_1_13, q_1_12=>
      que_out_10_1_12, q_1_11=>que_out_10_1_11, q_1_10=>que_out_10_1_10, 
      q_1_9=>que_out_10_1_9, q_1_8=>que_out_10_1_8, q_1_7=>que_out_10_1_7, 
      q_1_6=>que_out_10_1_6, q_1_5=>que_out_10_1_5, q_1_4=>que_out_10_1_4, 
      q_1_3=>que_out_10_1_3, q_1_2=>que_out_10_1_2, q_1_1=>que_out_10_1_1, 
      q_1_0=>que_out_10_1_0, q_2_15=>que_out_10_2_15, q_2_14=>
      que_out_10_2_14, q_2_13=>que_out_10_2_13, q_2_12=>que_out_10_2_12, 
      q_2_11=>que_out_10_2_11, q_2_10=>que_out_10_2_10, q_2_9=>
      que_out_10_2_9, q_2_8=>que_out_10_2_8, q_2_7=>que_out_10_2_7, q_2_6=>
      que_out_10_2_6, q_2_5=>que_out_10_2_5, q_2_4=>que_out_10_2_4, q_2_3=>
      que_out_10_2_3, q_2_2=>que_out_10_2_2, q_2_1=>que_out_10_2_1, q_2_0=>
      que_out_10_2_0, q_3_15=>que_out_10_3_15, q_3_14=>que_out_10_3_14, 
      q_3_13=>que_out_10_3_13, q_3_12=>que_out_10_3_12, q_3_11=>
      que_out_10_3_11, q_3_10=>que_out_10_3_10, q_3_9=>que_out_10_3_9, q_3_8
      =>que_out_10_3_8, q_3_7=>que_out_10_3_7, q_3_6=>que_out_10_3_6, q_3_5
      =>que_out_10_3_5, q_3_4=>que_out_10_3_4, q_3_3=>que_out_10_3_3, q_3_2
      =>que_out_10_3_2, q_3_1=>que_out_10_3_1, q_3_0=>que_out_10_3_0, q_4_15
      =>que_out_10_4_15, q_4_14=>que_out_10_4_14, q_4_13=>que_out_10_4_13, 
      q_4_12=>que_out_10_4_12, q_4_11=>que_out_10_4_11, q_4_10=>
      que_out_10_4_10, q_4_9=>que_out_10_4_9, q_4_8=>que_out_10_4_8, q_4_7=>
      que_out_10_4_7, q_4_6=>que_out_10_4_6, q_4_5=>que_out_10_4_5, q_4_4=>
      que_out_10_4_4, q_4_3=>que_out_10_4_3, q_4_2=>que_out_10_4_2, q_4_1=>
      que_out_10_4_1, q_4_0=>que_out_10_4_0, clk=>nx10722, load=>sel_que_10, 
      reset=>nx10698);
   gen_queues_11_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_11_0_15, q_0_14=>que_out_11_0_14, q_0_13=>
      que_out_11_0_13, q_0_12=>que_out_11_0_12, q_0_11=>que_out_11_0_11, 
      q_0_10=>que_out_11_0_10, q_0_9=>que_out_11_0_9, q_0_8=>que_out_11_0_8, 
      q_0_7=>que_out_11_0_7, q_0_6=>que_out_11_0_6, q_0_5=>que_out_11_0_5, 
      q_0_4=>que_out_11_0_4, q_0_3=>que_out_11_0_3, q_0_2=>que_out_11_0_2, 
      q_0_1=>que_out_11_0_1, q_0_0=>que_out_11_0_0, q_1_15=>que_out_11_1_15, 
      q_1_14=>que_out_11_1_14, q_1_13=>que_out_11_1_13, q_1_12=>
      que_out_11_1_12, q_1_11=>que_out_11_1_11, q_1_10=>que_out_11_1_10, 
      q_1_9=>que_out_11_1_9, q_1_8=>que_out_11_1_8, q_1_7=>que_out_11_1_7, 
      q_1_6=>que_out_11_1_6, q_1_5=>que_out_11_1_5, q_1_4=>que_out_11_1_4, 
      q_1_3=>que_out_11_1_3, q_1_2=>que_out_11_1_2, q_1_1=>que_out_11_1_1, 
      q_1_0=>que_out_11_1_0, q_2_15=>que_out_11_2_15, q_2_14=>
      que_out_11_2_14, q_2_13=>que_out_11_2_13, q_2_12=>que_out_11_2_12, 
      q_2_11=>que_out_11_2_11, q_2_10=>que_out_11_2_10, q_2_9=>
      que_out_11_2_9, q_2_8=>que_out_11_2_8, q_2_7=>que_out_11_2_7, q_2_6=>
      que_out_11_2_6, q_2_5=>que_out_11_2_5, q_2_4=>que_out_11_2_4, q_2_3=>
      que_out_11_2_3, q_2_2=>que_out_11_2_2, q_2_1=>que_out_11_2_1, q_2_0=>
      que_out_11_2_0, q_3_15=>que_out_11_3_15, q_3_14=>que_out_11_3_14, 
      q_3_13=>que_out_11_3_13, q_3_12=>que_out_11_3_12, q_3_11=>
      que_out_11_3_11, q_3_10=>que_out_11_3_10, q_3_9=>que_out_11_3_9, q_3_8
      =>que_out_11_3_8, q_3_7=>que_out_11_3_7, q_3_6=>que_out_11_3_6, q_3_5
      =>que_out_11_3_5, q_3_4=>que_out_11_3_4, q_3_3=>que_out_11_3_3, q_3_2
      =>que_out_11_3_2, q_3_1=>que_out_11_3_1, q_3_0=>que_out_11_3_0, q_4_15
      =>que_out_11_4_15, q_4_14=>que_out_11_4_14, q_4_13=>que_out_11_4_13, 
      q_4_12=>que_out_11_4_12, q_4_11=>que_out_11_4_11, q_4_10=>
      que_out_11_4_10, q_4_9=>que_out_11_4_9, q_4_8=>que_out_11_4_8, q_4_7=>
      que_out_11_4_7, q_4_6=>que_out_11_4_6, q_4_5=>que_out_11_4_5, q_4_4=>
      que_out_11_4_4, q_4_3=>que_out_11_4_3, q_4_2=>que_out_11_4_2, q_4_1=>
      que_out_11_4_1, q_4_0=>que_out_11_4_0, clk=>nx10722, load=>sel_que_11, 
      reset=>nx10698);
   gen_queues_12_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_12_0_15, q_0_14=>que_out_12_0_14, q_0_13=>
      que_out_12_0_13, q_0_12=>que_out_12_0_12, q_0_11=>que_out_12_0_11, 
      q_0_10=>que_out_12_0_10, q_0_9=>que_out_12_0_9, q_0_8=>que_out_12_0_8, 
      q_0_7=>que_out_12_0_7, q_0_6=>que_out_12_0_6, q_0_5=>que_out_12_0_5, 
      q_0_4=>que_out_12_0_4, q_0_3=>que_out_12_0_3, q_0_2=>que_out_12_0_2, 
      q_0_1=>que_out_12_0_1, q_0_0=>que_out_12_0_0, q_1_15=>que_out_12_1_15, 
      q_1_14=>que_out_12_1_14, q_1_13=>que_out_12_1_13, q_1_12=>
      que_out_12_1_12, q_1_11=>que_out_12_1_11, q_1_10=>que_out_12_1_10, 
      q_1_9=>que_out_12_1_9, q_1_8=>que_out_12_1_8, q_1_7=>que_out_12_1_7, 
      q_1_6=>que_out_12_1_6, q_1_5=>que_out_12_1_5, q_1_4=>que_out_12_1_4, 
      q_1_3=>que_out_12_1_3, q_1_2=>que_out_12_1_2, q_1_1=>que_out_12_1_1, 
      q_1_0=>que_out_12_1_0, q_2_15=>que_out_12_2_15, q_2_14=>
      que_out_12_2_14, q_2_13=>que_out_12_2_13, q_2_12=>que_out_12_2_12, 
      q_2_11=>que_out_12_2_11, q_2_10=>que_out_12_2_10, q_2_9=>
      que_out_12_2_9, q_2_8=>que_out_12_2_8, q_2_7=>que_out_12_2_7, q_2_6=>
      que_out_12_2_6, q_2_5=>que_out_12_2_5, q_2_4=>que_out_12_2_4, q_2_3=>
      que_out_12_2_3, q_2_2=>que_out_12_2_2, q_2_1=>que_out_12_2_1, q_2_0=>
      que_out_12_2_0, q_3_15=>que_out_12_3_15, q_3_14=>que_out_12_3_14, 
      q_3_13=>que_out_12_3_13, q_3_12=>que_out_12_3_12, q_3_11=>
      que_out_12_3_11, q_3_10=>que_out_12_3_10, q_3_9=>que_out_12_3_9, q_3_8
      =>que_out_12_3_8, q_3_7=>que_out_12_3_7, q_3_6=>que_out_12_3_6, q_3_5
      =>que_out_12_3_5, q_3_4=>que_out_12_3_4, q_3_3=>que_out_12_3_3, q_3_2
      =>que_out_12_3_2, q_3_1=>que_out_12_3_1, q_3_0=>que_out_12_3_0, q_4_15
      =>que_out_12_4_15, q_4_14=>que_out_12_4_14, q_4_13=>que_out_12_4_13, 
      q_4_12=>que_out_12_4_12, q_4_11=>que_out_12_4_11, q_4_10=>
      que_out_12_4_10, q_4_9=>que_out_12_4_9, q_4_8=>que_out_12_4_8, q_4_7=>
      que_out_12_4_7, q_4_6=>que_out_12_4_6, q_4_5=>que_out_12_4_5, q_4_4=>
      que_out_12_4_4, q_4_3=>que_out_12_4_3, q_4_2=>que_out_12_4_2, q_4_1=>
      que_out_12_4_1, q_4_0=>que_out_12_4_0, clk=>nx10722, load=>sel_que_12, 
      reset=>nx10698);
   gen_queues_13_que : Queue_5 port map ( d(15)=>nx10514, d(14)=>nx10524, 
      d(13)=>nx10534, d(12)=>nx10544, d(11)=>nx10554, d(10)=>nx10564, d(9)=>
      nx10574, d(8)=>nx10584, d(7)=>nx10594, d(6)=>nx10604, d(5)=>nx10614, 
      d(4)=>nx10624, d(3)=>nx10634, d(2)=>nx10644, d(1)=>nx10654, d(0)=>
      nx10664, q_0_15=>que_out_13_0_15, q_0_14=>que_out_13_0_14, q_0_13=>
      que_out_13_0_13, q_0_12=>que_out_13_0_12, q_0_11=>que_out_13_0_11, 
      q_0_10=>que_out_13_0_10, q_0_9=>que_out_13_0_9, q_0_8=>que_out_13_0_8, 
      q_0_7=>que_out_13_0_7, q_0_6=>que_out_13_0_6, q_0_5=>que_out_13_0_5, 
      q_0_4=>que_out_13_0_4, q_0_3=>que_out_13_0_3, q_0_2=>que_out_13_0_2, 
      q_0_1=>que_out_13_0_1, q_0_0=>que_out_13_0_0, q_1_15=>que_out_13_1_15, 
      q_1_14=>que_out_13_1_14, q_1_13=>que_out_13_1_13, q_1_12=>
      que_out_13_1_12, q_1_11=>que_out_13_1_11, q_1_10=>que_out_13_1_10, 
      q_1_9=>que_out_13_1_9, q_1_8=>que_out_13_1_8, q_1_7=>que_out_13_1_7, 
      q_1_6=>que_out_13_1_6, q_1_5=>que_out_13_1_5, q_1_4=>que_out_13_1_4, 
      q_1_3=>que_out_13_1_3, q_1_2=>que_out_13_1_2, q_1_1=>que_out_13_1_1, 
      q_1_0=>que_out_13_1_0, q_2_15=>que_out_13_2_15, q_2_14=>
      que_out_13_2_14, q_2_13=>que_out_13_2_13, q_2_12=>que_out_13_2_12, 
      q_2_11=>que_out_13_2_11, q_2_10=>que_out_13_2_10, q_2_9=>
      que_out_13_2_9, q_2_8=>que_out_13_2_8, q_2_7=>que_out_13_2_7, q_2_6=>
      que_out_13_2_6, q_2_5=>que_out_13_2_5, q_2_4=>que_out_13_2_4, q_2_3=>
      que_out_13_2_3, q_2_2=>que_out_13_2_2, q_2_1=>que_out_13_2_1, q_2_0=>
      que_out_13_2_0, q_3_15=>que_out_13_3_15, q_3_14=>que_out_13_3_14, 
      q_3_13=>que_out_13_3_13, q_3_12=>que_out_13_3_12, q_3_11=>
      que_out_13_3_11, q_3_10=>que_out_13_3_10, q_3_9=>que_out_13_3_9, q_3_8
      =>que_out_13_3_8, q_3_7=>que_out_13_3_7, q_3_6=>que_out_13_3_6, q_3_5
      =>que_out_13_3_5, q_3_4=>que_out_13_3_4, q_3_3=>que_out_13_3_3, q_3_2
      =>que_out_13_3_2, q_3_1=>que_out_13_3_1, q_3_0=>que_out_13_3_0, q_4_15
      =>que_out_13_4_15, q_4_14=>que_out_13_4_14, q_4_13=>que_out_13_4_13, 
      q_4_12=>que_out_13_4_12, q_4_11=>que_out_13_4_11, q_4_10=>
      que_out_13_4_10, q_4_9=>que_out_13_4_9, q_4_8=>que_out_13_4_8, q_4_7=>
      que_out_13_4_7, q_4_6=>que_out_13_4_6, q_4_5=>que_out_13_4_5, q_4_4=>
      que_out_13_4_4, q_4_3=>que_out_13_4_3, q_4_2=>que_out_13_4_2, q_4_1=>
      que_out_13_4_1, q_4_0=>que_out_13_4_0, clk=>nx10724, load=>sel_que_13, 
      reset=>nx10700);
   gen_queues_14_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_14_0_15, q_0_14=>que_out_14_0_14, q_0_13=>
      que_out_14_0_13, q_0_12=>que_out_14_0_12, q_0_11=>que_out_14_0_11, 
      q_0_10=>que_out_14_0_10, q_0_9=>que_out_14_0_9, q_0_8=>que_out_14_0_8, 
      q_0_7=>que_out_14_0_7, q_0_6=>que_out_14_0_6, q_0_5=>que_out_14_0_5, 
      q_0_4=>que_out_14_0_4, q_0_3=>que_out_14_0_3, q_0_2=>que_out_14_0_2, 
      q_0_1=>que_out_14_0_1, q_0_0=>que_out_14_0_0, q_1_15=>que_out_14_1_15, 
      q_1_14=>que_out_14_1_14, q_1_13=>que_out_14_1_13, q_1_12=>
      que_out_14_1_12, q_1_11=>que_out_14_1_11, q_1_10=>que_out_14_1_10, 
      q_1_9=>que_out_14_1_9, q_1_8=>que_out_14_1_8, q_1_7=>que_out_14_1_7, 
      q_1_6=>que_out_14_1_6, q_1_5=>que_out_14_1_5, q_1_4=>que_out_14_1_4, 
      q_1_3=>que_out_14_1_3, q_1_2=>que_out_14_1_2, q_1_1=>que_out_14_1_1, 
      q_1_0=>que_out_14_1_0, q_2_15=>que_out_14_2_15, q_2_14=>
      que_out_14_2_14, q_2_13=>que_out_14_2_13, q_2_12=>que_out_14_2_12, 
      q_2_11=>que_out_14_2_11, q_2_10=>que_out_14_2_10, q_2_9=>
      que_out_14_2_9, q_2_8=>que_out_14_2_8, q_2_7=>que_out_14_2_7, q_2_6=>
      que_out_14_2_6, q_2_5=>que_out_14_2_5, q_2_4=>que_out_14_2_4, q_2_3=>
      que_out_14_2_3, q_2_2=>que_out_14_2_2, q_2_1=>que_out_14_2_1, q_2_0=>
      que_out_14_2_0, q_3_15=>que_out_14_3_15, q_3_14=>que_out_14_3_14, 
      q_3_13=>que_out_14_3_13, q_3_12=>que_out_14_3_12, q_3_11=>
      que_out_14_3_11, q_3_10=>que_out_14_3_10, q_3_9=>que_out_14_3_9, q_3_8
      =>que_out_14_3_8, q_3_7=>que_out_14_3_7, q_3_6=>que_out_14_3_6, q_3_5
      =>que_out_14_3_5, q_3_4=>que_out_14_3_4, q_3_3=>que_out_14_3_3, q_3_2
      =>que_out_14_3_2, q_3_1=>que_out_14_3_1, q_3_0=>que_out_14_3_0, q_4_15
      =>que_out_14_4_15, q_4_14=>que_out_14_4_14, q_4_13=>que_out_14_4_13, 
      q_4_12=>que_out_14_4_12, q_4_11=>que_out_14_4_11, q_4_10=>
      que_out_14_4_10, q_4_9=>que_out_14_4_9, q_4_8=>que_out_14_4_8, q_4_7=>
      que_out_14_4_7, q_4_6=>que_out_14_4_6, q_4_5=>que_out_14_4_5, q_4_4=>
      que_out_14_4_4, q_4_3=>que_out_14_4_3, q_4_2=>que_out_14_4_2, q_4_1=>
      que_out_14_4_1, q_4_0=>que_out_14_4_0, clk=>nx10726, load=>sel_que_14, 
      reset=>nx10702);
   gen_queues_15_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_15_0_15, q_0_14=>que_out_15_0_14, q_0_13=>
      que_out_15_0_13, q_0_12=>que_out_15_0_12, q_0_11=>que_out_15_0_11, 
      q_0_10=>que_out_15_0_10, q_0_9=>que_out_15_0_9, q_0_8=>que_out_15_0_8, 
      q_0_7=>que_out_15_0_7, q_0_6=>que_out_15_0_6, q_0_5=>que_out_15_0_5, 
      q_0_4=>que_out_15_0_4, q_0_3=>que_out_15_0_3, q_0_2=>que_out_15_0_2, 
      q_0_1=>que_out_15_0_1, q_0_0=>que_out_15_0_0, q_1_15=>que_out_15_1_15, 
      q_1_14=>que_out_15_1_14, q_1_13=>que_out_15_1_13, q_1_12=>
      que_out_15_1_12, q_1_11=>que_out_15_1_11, q_1_10=>que_out_15_1_10, 
      q_1_9=>que_out_15_1_9, q_1_8=>que_out_15_1_8, q_1_7=>que_out_15_1_7, 
      q_1_6=>que_out_15_1_6, q_1_5=>que_out_15_1_5, q_1_4=>que_out_15_1_4, 
      q_1_3=>que_out_15_1_3, q_1_2=>que_out_15_1_2, q_1_1=>que_out_15_1_1, 
      q_1_0=>que_out_15_1_0, q_2_15=>que_out_15_2_15, q_2_14=>
      que_out_15_2_14, q_2_13=>que_out_15_2_13, q_2_12=>que_out_15_2_12, 
      q_2_11=>que_out_15_2_11, q_2_10=>que_out_15_2_10, q_2_9=>
      que_out_15_2_9, q_2_8=>que_out_15_2_8, q_2_7=>que_out_15_2_7, q_2_6=>
      que_out_15_2_6, q_2_5=>que_out_15_2_5, q_2_4=>que_out_15_2_4, q_2_3=>
      que_out_15_2_3, q_2_2=>que_out_15_2_2, q_2_1=>que_out_15_2_1, q_2_0=>
      que_out_15_2_0, q_3_15=>que_out_15_3_15, q_3_14=>que_out_15_3_14, 
      q_3_13=>que_out_15_3_13, q_3_12=>que_out_15_3_12, q_3_11=>
      que_out_15_3_11, q_3_10=>que_out_15_3_10, q_3_9=>que_out_15_3_9, q_3_8
      =>que_out_15_3_8, q_3_7=>que_out_15_3_7, q_3_6=>que_out_15_3_6, q_3_5
      =>que_out_15_3_5, q_3_4=>que_out_15_3_4, q_3_3=>que_out_15_3_3, q_3_2
      =>que_out_15_3_2, q_3_1=>que_out_15_3_1, q_3_0=>que_out_15_3_0, q_4_15
      =>que_out_15_4_15, q_4_14=>que_out_15_4_14, q_4_13=>que_out_15_4_13, 
      q_4_12=>que_out_15_4_12, q_4_11=>que_out_15_4_11, q_4_10=>
      que_out_15_4_10, q_4_9=>que_out_15_4_9, q_4_8=>que_out_15_4_8, q_4_7=>
      que_out_15_4_7, q_4_6=>que_out_15_4_6, q_4_5=>que_out_15_4_5, q_4_4=>
      que_out_15_4_4, q_4_3=>que_out_15_4_3, q_4_2=>que_out_15_4_2, q_4_1=>
      que_out_15_4_1, q_4_0=>que_out_15_4_0, clk=>nx10726, load=>sel_que_15, 
      reset=>nx10702);
   gen_queues_16_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_16_0_15, q_0_14=>que_out_16_0_14, q_0_13=>
      que_out_16_0_13, q_0_12=>que_out_16_0_12, q_0_11=>que_out_16_0_11, 
      q_0_10=>que_out_16_0_10, q_0_9=>que_out_16_0_9, q_0_8=>que_out_16_0_8, 
      q_0_7=>que_out_16_0_7, q_0_6=>que_out_16_0_6, q_0_5=>que_out_16_0_5, 
      q_0_4=>que_out_16_0_4, q_0_3=>que_out_16_0_3, q_0_2=>que_out_16_0_2, 
      q_0_1=>que_out_16_0_1, q_0_0=>que_out_16_0_0, q_1_15=>que_out_16_1_15, 
      q_1_14=>que_out_16_1_14, q_1_13=>que_out_16_1_13, q_1_12=>
      que_out_16_1_12, q_1_11=>que_out_16_1_11, q_1_10=>que_out_16_1_10, 
      q_1_9=>que_out_16_1_9, q_1_8=>que_out_16_1_8, q_1_7=>que_out_16_1_7, 
      q_1_6=>que_out_16_1_6, q_1_5=>que_out_16_1_5, q_1_4=>que_out_16_1_4, 
      q_1_3=>que_out_16_1_3, q_1_2=>que_out_16_1_2, q_1_1=>que_out_16_1_1, 
      q_1_0=>que_out_16_1_0, q_2_15=>que_out_16_2_15, q_2_14=>
      que_out_16_2_14, q_2_13=>que_out_16_2_13, q_2_12=>que_out_16_2_12, 
      q_2_11=>que_out_16_2_11, q_2_10=>que_out_16_2_10, q_2_9=>
      que_out_16_2_9, q_2_8=>que_out_16_2_8, q_2_7=>que_out_16_2_7, q_2_6=>
      que_out_16_2_6, q_2_5=>que_out_16_2_5, q_2_4=>que_out_16_2_4, q_2_3=>
      que_out_16_2_3, q_2_2=>que_out_16_2_2, q_2_1=>que_out_16_2_1, q_2_0=>
      que_out_16_2_0, q_3_15=>que_out_16_3_15, q_3_14=>que_out_16_3_14, 
      q_3_13=>que_out_16_3_13, q_3_12=>que_out_16_3_12, q_3_11=>
      que_out_16_3_11, q_3_10=>que_out_16_3_10, q_3_9=>que_out_16_3_9, q_3_8
      =>que_out_16_3_8, q_3_7=>que_out_16_3_7, q_3_6=>que_out_16_3_6, q_3_5
      =>que_out_16_3_5, q_3_4=>que_out_16_3_4, q_3_3=>que_out_16_3_3, q_3_2
      =>que_out_16_3_2, q_3_1=>que_out_16_3_1, q_3_0=>que_out_16_3_0, q_4_15
      =>que_out_16_4_15, q_4_14=>que_out_16_4_14, q_4_13=>que_out_16_4_13, 
      q_4_12=>que_out_16_4_12, q_4_11=>que_out_16_4_11, q_4_10=>
      que_out_16_4_10, q_4_9=>que_out_16_4_9, q_4_8=>que_out_16_4_8, q_4_7=>
      que_out_16_4_7, q_4_6=>que_out_16_4_6, q_4_5=>que_out_16_4_5, q_4_4=>
      que_out_16_4_4, q_4_3=>que_out_16_4_3, q_4_2=>que_out_16_4_2, q_4_1=>
      que_out_16_4_1, q_4_0=>que_out_16_4_0, clk=>nx10726, load=>sel_que_16, 
      reset=>nx10702);
   gen_queues_17_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_17_0_15, q_0_14=>que_out_17_0_14, q_0_13=>
      que_out_17_0_13, q_0_12=>que_out_17_0_12, q_0_11=>que_out_17_0_11, 
      q_0_10=>que_out_17_0_10, q_0_9=>que_out_17_0_9, q_0_8=>que_out_17_0_8, 
      q_0_7=>que_out_17_0_7, q_0_6=>que_out_17_0_6, q_0_5=>que_out_17_0_5, 
      q_0_4=>que_out_17_0_4, q_0_3=>que_out_17_0_3, q_0_2=>que_out_17_0_2, 
      q_0_1=>que_out_17_0_1, q_0_0=>que_out_17_0_0, q_1_15=>que_out_17_1_15, 
      q_1_14=>que_out_17_1_14, q_1_13=>que_out_17_1_13, q_1_12=>
      que_out_17_1_12, q_1_11=>que_out_17_1_11, q_1_10=>que_out_17_1_10, 
      q_1_9=>que_out_17_1_9, q_1_8=>que_out_17_1_8, q_1_7=>que_out_17_1_7, 
      q_1_6=>que_out_17_1_6, q_1_5=>que_out_17_1_5, q_1_4=>que_out_17_1_4, 
      q_1_3=>que_out_17_1_3, q_1_2=>que_out_17_1_2, q_1_1=>que_out_17_1_1, 
      q_1_0=>que_out_17_1_0, q_2_15=>que_out_17_2_15, q_2_14=>
      que_out_17_2_14, q_2_13=>que_out_17_2_13, q_2_12=>que_out_17_2_12, 
      q_2_11=>que_out_17_2_11, q_2_10=>que_out_17_2_10, q_2_9=>
      que_out_17_2_9, q_2_8=>que_out_17_2_8, q_2_7=>que_out_17_2_7, q_2_6=>
      que_out_17_2_6, q_2_5=>que_out_17_2_5, q_2_4=>que_out_17_2_4, q_2_3=>
      que_out_17_2_3, q_2_2=>que_out_17_2_2, q_2_1=>que_out_17_2_1, q_2_0=>
      que_out_17_2_0, q_3_15=>que_out_17_3_15, q_3_14=>que_out_17_3_14, 
      q_3_13=>que_out_17_3_13, q_3_12=>que_out_17_3_12, q_3_11=>
      que_out_17_3_11, q_3_10=>que_out_17_3_10, q_3_9=>que_out_17_3_9, q_3_8
      =>que_out_17_3_8, q_3_7=>que_out_17_3_7, q_3_6=>que_out_17_3_6, q_3_5
      =>que_out_17_3_5, q_3_4=>que_out_17_3_4, q_3_3=>que_out_17_3_3, q_3_2
      =>que_out_17_3_2, q_3_1=>que_out_17_3_1, q_3_0=>que_out_17_3_0, q_4_15
      =>que_out_17_4_15, q_4_14=>que_out_17_4_14, q_4_13=>que_out_17_4_13, 
      q_4_12=>que_out_17_4_12, q_4_11=>que_out_17_4_11, q_4_10=>
      que_out_17_4_10, q_4_9=>que_out_17_4_9, q_4_8=>que_out_17_4_8, q_4_7=>
      que_out_17_4_7, q_4_6=>que_out_17_4_6, q_4_5=>que_out_17_4_5, q_4_4=>
      que_out_17_4_4, q_4_3=>que_out_17_4_3, q_4_2=>que_out_17_4_2, q_4_1=>
      que_out_17_4_1, q_4_0=>que_out_17_4_0, clk=>nx10728, load=>sel_que_17, 
      reset=>nx10704);
   gen_queues_18_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_18_0_15, q_0_14=>que_out_18_0_14, q_0_13=>
      que_out_18_0_13, q_0_12=>que_out_18_0_12, q_0_11=>que_out_18_0_11, 
      q_0_10=>que_out_18_0_10, q_0_9=>que_out_18_0_9, q_0_8=>que_out_18_0_8, 
      q_0_7=>que_out_18_0_7, q_0_6=>que_out_18_0_6, q_0_5=>que_out_18_0_5, 
      q_0_4=>que_out_18_0_4, q_0_3=>que_out_18_0_3, q_0_2=>que_out_18_0_2, 
      q_0_1=>que_out_18_0_1, q_0_0=>que_out_18_0_0, q_1_15=>que_out_18_1_15, 
      q_1_14=>que_out_18_1_14, q_1_13=>que_out_18_1_13, q_1_12=>
      que_out_18_1_12, q_1_11=>que_out_18_1_11, q_1_10=>que_out_18_1_10, 
      q_1_9=>que_out_18_1_9, q_1_8=>que_out_18_1_8, q_1_7=>que_out_18_1_7, 
      q_1_6=>que_out_18_1_6, q_1_5=>que_out_18_1_5, q_1_4=>que_out_18_1_4, 
      q_1_3=>que_out_18_1_3, q_1_2=>que_out_18_1_2, q_1_1=>que_out_18_1_1, 
      q_1_0=>que_out_18_1_0, q_2_15=>que_out_18_2_15, q_2_14=>
      que_out_18_2_14, q_2_13=>que_out_18_2_13, q_2_12=>que_out_18_2_12, 
      q_2_11=>que_out_18_2_11, q_2_10=>que_out_18_2_10, q_2_9=>
      que_out_18_2_9, q_2_8=>que_out_18_2_8, q_2_7=>que_out_18_2_7, q_2_6=>
      que_out_18_2_6, q_2_5=>que_out_18_2_5, q_2_4=>que_out_18_2_4, q_2_3=>
      que_out_18_2_3, q_2_2=>que_out_18_2_2, q_2_1=>que_out_18_2_1, q_2_0=>
      que_out_18_2_0, q_3_15=>que_out_18_3_15, q_3_14=>que_out_18_3_14, 
      q_3_13=>que_out_18_3_13, q_3_12=>que_out_18_3_12, q_3_11=>
      que_out_18_3_11, q_3_10=>que_out_18_3_10, q_3_9=>que_out_18_3_9, q_3_8
      =>que_out_18_3_8, q_3_7=>que_out_18_3_7, q_3_6=>que_out_18_3_6, q_3_5
      =>que_out_18_3_5, q_3_4=>que_out_18_3_4, q_3_3=>que_out_18_3_3, q_3_2
      =>que_out_18_3_2, q_3_1=>que_out_18_3_1, q_3_0=>que_out_18_3_0, q_4_15
      =>que_out_18_4_15, q_4_14=>que_out_18_4_14, q_4_13=>que_out_18_4_13, 
      q_4_12=>que_out_18_4_12, q_4_11=>que_out_18_4_11, q_4_10=>
      que_out_18_4_10, q_4_9=>que_out_18_4_9, q_4_8=>que_out_18_4_8, q_4_7=>
      que_out_18_4_7, q_4_6=>que_out_18_4_6, q_4_5=>que_out_18_4_5, q_4_4=>
      que_out_18_4_4, q_4_3=>que_out_18_4_3, q_4_2=>que_out_18_4_2, q_4_1=>
      que_out_18_4_1, q_4_0=>que_out_18_4_0, clk=>nx10728, load=>sel_que_18, 
      reset=>nx10704);
   gen_queues_19_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_19_0_15, q_0_14=>que_out_19_0_14, q_0_13=>
      que_out_19_0_13, q_0_12=>que_out_19_0_12, q_0_11=>que_out_19_0_11, 
      q_0_10=>que_out_19_0_10, q_0_9=>que_out_19_0_9, q_0_8=>que_out_19_0_8, 
      q_0_7=>que_out_19_0_7, q_0_6=>que_out_19_0_6, q_0_5=>que_out_19_0_5, 
      q_0_4=>que_out_19_0_4, q_0_3=>que_out_19_0_3, q_0_2=>que_out_19_0_2, 
      q_0_1=>que_out_19_0_1, q_0_0=>que_out_19_0_0, q_1_15=>que_out_19_1_15, 
      q_1_14=>que_out_19_1_14, q_1_13=>que_out_19_1_13, q_1_12=>
      que_out_19_1_12, q_1_11=>que_out_19_1_11, q_1_10=>que_out_19_1_10, 
      q_1_9=>que_out_19_1_9, q_1_8=>que_out_19_1_8, q_1_7=>que_out_19_1_7, 
      q_1_6=>que_out_19_1_6, q_1_5=>que_out_19_1_5, q_1_4=>que_out_19_1_4, 
      q_1_3=>que_out_19_1_3, q_1_2=>que_out_19_1_2, q_1_1=>que_out_19_1_1, 
      q_1_0=>que_out_19_1_0, q_2_15=>que_out_19_2_15, q_2_14=>
      que_out_19_2_14, q_2_13=>que_out_19_2_13, q_2_12=>que_out_19_2_12, 
      q_2_11=>que_out_19_2_11, q_2_10=>que_out_19_2_10, q_2_9=>
      que_out_19_2_9, q_2_8=>que_out_19_2_8, q_2_7=>que_out_19_2_7, q_2_6=>
      que_out_19_2_6, q_2_5=>que_out_19_2_5, q_2_4=>que_out_19_2_4, q_2_3=>
      que_out_19_2_3, q_2_2=>que_out_19_2_2, q_2_1=>que_out_19_2_1, q_2_0=>
      que_out_19_2_0, q_3_15=>que_out_19_3_15, q_3_14=>que_out_19_3_14, 
      q_3_13=>que_out_19_3_13, q_3_12=>que_out_19_3_12, q_3_11=>
      que_out_19_3_11, q_3_10=>que_out_19_3_10, q_3_9=>que_out_19_3_9, q_3_8
      =>que_out_19_3_8, q_3_7=>que_out_19_3_7, q_3_6=>que_out_19_3_6, q_3_5
      =>que_out_19_3_5, q_3_4=>que_out_19_3_4, q_3_3=>que_out_19_3_3, q_3_2
      =>que_out_19_3_2, q_3_1=>que_out_19_3_1, q_3_0=>que_out_19_3_0, q_4_15
      =>que_out_19_4_15, q_4_14=>que_out_19_4_14, q_4_13=>que_out_19_4_13, 
      q_4_12=>que_out_19_4_12, q_4_11=>que_out_19_4_11, q_4_10=>
      que_out_19_4_10, q_4_9=>que_out_19_4_9, q_4_8=>que_out_19_4_8, q_4_7=>
      que_out_19_4_7, q_4_6=>que_out_19_4_6, q_4_5=>que_out_19_4_5, q_4_4=>
      que_out_19_4_4, q_4_3=>que_out_19_4_3, q_4_2=>que_out_19_4_2, q_4_1=>
      que_out_19_4_1, q_4_0=>que_out_19_4_0, clk=>nx10728, load=>sel_que_19, 
      reset=>nx10704);
   gen_queues_20_que : Queue_5 port map ( d(15)=>nx10516, d(14)=>nx10526, 
      d(13)=>nx10536, d(12)=>nx10546, d(11)=>nx10556, d(10)=>nx10566, d(9)=>
      nx10576, d(8)=>nx10586, d(7)=>nx10596, d(6)=>nx10606, d(5)=>nx10616, 
      d(4)=>nx10626, d(3)=>nx10636, d(2)=>nx10646, d(1)=>nx10656, d(0)=>
      nx10666, q_0_15=>que_out_20_0_15, q_0_14=>que_out_20_0_14, q_0_13=>
      que_out_20_0_13, q_0_12=>que_out_20_0_12, q_0_11=>que_out_20_0_11, 
      q_0_10=>que_out_20_0_10, q_0_9=>que_out_20_0_9, q_0_8=>que_out_20_0_8, 
      q_0_7=>que_out_20_0_7, q_0_6=>que_out_20_0_6, q_0_5=>que_out_20_0_5, 
      q_0_4=>que_out_20_0_4, q_0_3=>que_out_20_0_3, q_0_2=>que_out_20_0_2, 
      q_0_1=>que_out_20_0_1, q_0_0=>que_out_20_0_0, q_1_15=>que_out_20_1_15, 
      q_1_14=>que_out_20_1_14, q_1_13=>que_out_20_1_13, q_1_12=>
      que_out_20_1_12, q_1_11=>que_out_20_1_11, q_1_10=>que_out_20_1_10, 
      q_1_9=>que_out_20_1_9, q_1_8=>que_out_20_1_8, q_1_7=>que_out_20_1_7, 
      q_1_6=>que_out_20_1_6, q_1_5=>que_out_20_1_5, q_1_4=>que_out_20_1_4, 
      q_1_3=>que_out_20_1_3, q_1_2=>que_out_20_1_2, q_1_1=>que_out_20_1_1, 
      q_1_0=>que_out_20_1_0, q_2_15=>que_out_20_2_15, q_2_14=>
      que_out_20_2_14, q_2_13=>que_out_20_2_13, q_2_12=>que_out_20_2_12, 
      q_2_11=>que_out_20_2_11, q_2_10=>que_out_20_2_10, q_2_9=>
      que_out_20_2_9, q_2_8=>que_out_20_2_8, q_2_7=>que_out_20_2_7, q_2_6=>
      que_out_20_2_6, q_2_5=>que_out_20_2_5, q_2_4=>que_out_20_2_4, q_2_3=>
      que_out_20_2_3, q_2_2=>que_out_20_2_2, q_2_1=>que_out_20_2_1, q_2_0=>
      que_out_20_2_0, q_3_15=>que_out_20_3_15, q_3_14=>que_out_20_3_14, 
      q_3_13=>que_out_20_3_13, q_3_12=>que_out_20_3_12, q_3_11=>
      que_out_20_3_11, q_3_10=>que_out_20_3_10, q_3_9=>que_out_20_3_9, q_3_8
      =>que_out_20_3_8, q_3_7=>que_out_20_3_7, q_3_6=>que_out_20_3_6, q_3_5
      =>que_out_20_3_5, q_3_4=>que_out_20_3_4, q_3_3=>que_out_20_3_3, q_3_2
      =>que_out_20_3_2, q_3_1=>que_out_20_3_1, q_3_0=>que_out_20_3_0, q_4_15
      =>que_out_20_4_15, q_4_14=>que_out_20_4_14, q_4_13=>que_out_20_4_13, 
      q_4_12=>que_out_20_4_12, q_4_11=>que_out_20_4_11, q_4_10=>
      que_out_20_4_10, q_4_9=>que_out_20_4_9, q_4_8=>que_out_20_4_8, q_4_7=>
      que_out_20_4_7, q_4_6=>que_out_20_4_6, q_4_5=>que_out_20_4_5, q_4_4=>
      que_out_20_4_4, q_4_3=>que_out_20_4_3, q_4_2=>que_out_20_4_2, q_4_1=>
      que_out_20_4_1, q_4_0=>que_out_20_4_0, clk=>nx10730, load=>sel_que_20, 
      reset=>nx10706);
   gen_queues_21_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_21_0_15, q_0_14=>que_out_21_0_14, q_0_13=>
      que_out_21_0_13, q_0_12=>que_out_21_0_12, q_0_11=>que_out_21_0_11, 
      q_0_10=>que_out_21_0_10, q_0_9=>que_out_21_0_9, q_0_8=>que_out_21_0_8, 
      q_0_7=>que_out_21_0_7, q_0_6=>que_out_21_0_6, q_0_5=>que_out_21_0_5, 
      q_0_4=>que_out_21_0_4, q_0_3=>que_out_21_0_3, q_0_2=>que_out_21_0_2, 
      q_0_1=>que_out_21_0_1, q_0_0=>que_out_21_0_0, q_1_15=>que_out_21_1_15, 
      q_1_14=>que_out_21_1_14, q_1_13=>que_out_21_1_13, q_1_12=>
      que_out_21_1_12, q_1_11=>que_out_21_1_11, q_1_10=>que_out_21_1_10, 
      q_1_9=>que_out_21_1_9, q_1_8=>que_out_21_1_8, q_1_7=>que_out_21_1_7, 
      q_1_6=>que_out_21_1_6, q_1_5=>que_out_21_1_5, q_1_4=>que_out_21_1_4, 
      q_1_3=>que_out_21_1_3, q_1_2=>que_out_21_1_2, q_1_1=>que_out_21_1_1, 
      q_1_0=>que_out_21_1_0, q_2_15=>que_out_21_2_15, q_2_14=>
      que_out_21_2_14, q_2_13=>que_out_21_2_13, q_2_12=>que_out_21_2_12, 
      q_2_11=>que_out_21_2_11, q_2_10=>que_out_21_2_10, q_2_9=>
      que_out_21_2_9, q_2_8=>que_out_21_2_8, q_2_7=>que_out_21_2_7, q_2_6=>
      que_out_21_2_6, q_2_5=>que_out_21_2_5, q_2_4=>que_out_21_2_4, q_2_3=>
      que_out_21_2_3, q_2_2=>que_out_21_2_2, q_2_1=>que_out_21_2_1, q_2_0=>
      que_out_21_2_0, q_3_15=>que_out_21_3_15, q_3_14=>que_out_21_3_14, 
      q_3_13=>que_out_21_3_13, q_3_12=>que_out_21_3_12, q_3_11=>
      que_out_21_3_11, q_3_10=>que_out_21_3_10, q_3_9=>que_out_21_3_9, q_3_8
      =>que_out_21_3_8, q_3_7=>que_out_21_3_7, q_3_6=>que_out_21_3_6, q_3_5
      =>que_out_21_3_5, q_3_4=>que_out_21_3_4, q_3_3=>que_out_21_3_3, q_3_2
      =>que_out_21_3_2, q_3_1=>que_out_21_3_1, q_3_0=>que_out_21_3_0, q_4_15
      =>que_out_21_4_15, q_4_14=>que_out_21_4_14, q_4_13=>que_out_21_4_13, 
      q_4_12=>que_out_21_4_12, q_4_11=>que_out_21_4_11, q_4_10=>
      que_out_21_4_10, q_4_9=>que_out_21_4_9, q_4_8=>que_out_21_4_8, q_4_7=>
      que_out_21_4_7, q_4_6=>que_out_21_4_6, q_4_5=>que_out_21_4_5, q_4_4=>
      que_out_21_4_4, q_4_3=>que_out_21_4_3, q_4_2=>que_out_21_4_2, q_4_1=>
      que_out_21_4_1, q_4_0=>que_out_21_4_0, clk=>nx10732, load=>sel_que_21, 
      reset=>nx10708);
   gen_queues_22_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_22_0_15, q_0_14=>que_out_22_0_14, q_0_13=>
      que_out_22_0_13, q_0_12=>que_out_22_0_12, q_0_11=>que_out_22_0_11, 
      q_0_10=>que_out_22_0_10, q_0_9=>que_out_22_0_9, q_0_8=>que_out_22_0_8, 
      q_0_7=>que_out_22_0_7, q_0_6=>que_out_22_0_6, q_0_5=>que_out_22_0_5, 
      q_0_4=>que_out_22_0_4, q_0_3=>que_out_22_0_3, q_0_2=>que_out_22_0_2, 
      q_0_1=>que_out_22_0_1, q_0_0=>que_out_22_0_0, q_1_15=>que_out_22_1_15, 
      q_1_14=>que_out_22_1_14, q_1_13=>que_out_22_1_13, q_1_12=>
      que_out_22_1_12, q_1_11=>que_out_22_1_11, q_1_10=>que_out_22_1_10, 
      q_1_9=>que_out_22_1_9, q_1_8=>que_out_22_1_8, q_1_7=>que_out_22_1_7, 
      q_1_6=>que_out_22_1_6, q_1_5=>que_out_22_1_5, q_1_4=>que_out_22_1_4, 
      q_1_3=>que_out_22_1_3, q_1_2=>que_out_22_1_2, q_1_1=>que_out_22_1_1, 
      q_1_0=>que_out_22_1_0, q_2_15=>que_out_22_2_15, q_2_14=>
      que_out_22_2_14, q_2_13=>que_out_22_2_13, q_2_12=>que_out_22_2_12, 
      q_2_11=>que_out_22_2_11, q_2_10=>que_out_22_2_10, q_2_9=>
      que_out_22_2_9, q_2_8=>que_out_22_2_8, q_2_7=>que_out_22_2_7, q_2_6=>
      que_out_22_2_6, q_2_5=>que_out_22_2_5, q_2_4=>que_out_22_2_4, q_2_3=>
      que_out_22_2_3, q_2_2=>que_out_22_2_2, q_2_1=>que_out_22_2_1, q_2_0=>
      que_out_22_2_0, q_3_15=>que_out_22_3_15, q_3_14=>que_out_22_3_14, 
      q_3_13=>que_out_22_3_13, q_3_12=>que_out_22_3_12, q_3_11=>
      que_out_22_3_11, q_3_10=>que_out_22_3_10, q_3_9=>que_out_22_3_9, q_3_8
      =>que_out_22_3_8, q_3_7=>que_out_22_3_7, q_3_6=>que_out_22_3_6, q_3_5
      =>que_out_22_3_5, q_3_4=>que_out_22_3_4, q_3_3=>que_out_22_3_3, q_3_2
      =>que_out_22_3_2, q_3_1=>que_out_22_3_1, q_3_0=>que_out_22_3_0, q_4_15
      =>que_out_22_4_15, q_4_14=>que_out_22_4_14, q_4_13=>que_out_22_4_13, 
      q_4_12=>que_out_22_4_12, q_4_11=>que_out_22_4_11, q_4_10=>
      que_out_22_4_10, q_4_9=>que_out_22_4_9, q_4_8=>que_out_22_4_8, q_4_7=>
      que_out_22_4_7, q_4_6=>que_out_22_4_6, q_4_5=>que_out_22_4_5, q_4_4=>
      que_out_22_4_4, q_4_3=>que_out_22_4_3, q_4_2=>que_out_22_4_2, q_4_1=>
      que_out_22_4_1, q_4_0=>que_out_22_4_0, clk=>nx10732, load=>sel_que_22, 
      reset=>nx10708);
   gen_queues_23_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_23_0_15, q_0_14=>que_out_23_0_14, q_0_13=>
      que_out_23_0_13, q_0_12=>que_out_23_0_12, q_0_11=>que_out_23_0_11, 
      q_0_10=>que_out_23_0_10, q_0_9=>que_out_23_0_9, q_0_8=>que_out_23_0_8, 
      q_0_7=>que_out_23_0_7, q_0_6=>que_out_23_0_6, q_0_5=>que_out_23_0_5, 
      q_0_4=>que_out_23_0_4, q_0_3=>que_out_23_0_3, q_0_2=>que_out_23_0_2, 
      q_0_1=>que_out_23_0_1, q_0_0=>que_out_23_0_0, q_1_15=>que_out_23_1_15, 
      q_1_14=>que_out_23_1_14, q_1_13=>que_out_23_1_13, q_1_12=>
      que_out_23_1_12, q_1_11=>que_out_23_1_11, q_1_10=>que_out_23_1_10, 
      q_1_9=>que_out_23_1_9, q_1_8=>que_out_23_1_8, q_1_7=>que_out_23_1_7, 
      q_1_6=>que_out_23_1_6, q_1_5=>que_out_23_1_5, q_1_4=>que_out_23_1_4, 
      q_1_3=>que_out_23_1_3, q_1_2=>que_out_23_1_2, q_1_1=>que_out_23_1_1, 
      q_1_0=>que_out_23_1_0, q_2_15=>que_out_23_2_15, q_2_14=>
      que_out_23_2_14, q_2_13=>que_out_23_2_13, q_2_12=>que_out_23_2_12, 
      q_2_11=>que_out_23_2_11, q_2_10=>que_out_23_2_10, q_2_9=>
      que_out_23_2_9, q_2_8=>que_out_23_2_8, q_2_7=>que_out_23_2_7, q_2_6=>
      que_out_23_2_6, q_2_5=>que_out_23_2_5, q_2_4=>que_out_23_2_4, q_2_3=>
      que_out_23_2_3, q_2_2=>que_out_23_2_2, q_2_1=>que_out_23_2_1, q_2_0=>
      que_out_23_2_0, q_3_15=>que_out_23_3_15, q_3_14=>que_out_23_3_14, 
      q_3_13=>que_out_23_3_13, q_3_12=>que_out_23_3_12, q_3_11=>
      que_out_23_3_11, q_3_10=>que_out_23_3_10, q_3_9=>que_out_23_3_9, q_3_8
      =>que_out_23_3_8, q_3_7=>que_out_23_3_7, q_3_6=>que_out_23_3_6, q_3_5
      =>que_out_23_3_5, q_3_4=>que_out_23_3_4, q_3_3=>que_out_23_3_3, q_3_2
      =>que_out_23_3_2, q_3_1=>que_out_23_3_1, q_3_0=>que_out_23_3_0, q_4_15
      =>que_out_23_4_15, q_4_14=>que_out_23_4_14, q_4_13=>que_out_23_4_13, 
      q_4_12=>que_out_23_4_12, q_4_11=>que_out_23_4_11, q_4_10=>
      que_out_23_4_10, q_4_9=>que_out_23_4_9, q_4_8=>que_out_23_4_8, q_4_7=>
      que_out_23_4_7, q_4_6=>que_out_23_4_6, q_4_5=>que_out_23_4_5, q_4_4=>
      que_out_23_4_4, q_4_3=>que_out_23_4_3, q_4_2=>que_out_23_4_2, q_4_1=>
      que_out_23_4_1, q_4_0=>que_out_23_4_0, clk=>nx10732, load=>sel_que_23, 
      reset=>nx10708);
   gen_queues_24_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_24_0_15, q_0_14=>que_out_24_0_14, q_0_13=>
      que_out_24_0_13, q_0_12=>que_out_24_0_12, q_0_11=>que_out_24_0_11, 
      q_0_10=>que_out_24_0_10, q_0_9=>que_out_24_0_9, q_0_8=>que_out_24_0_8, 
      q_0_7=>que_out_24_0_7, q_0_6=>que_out_24_0_6, q_0_5=>que_out_24_0_5, 
      q_0_4=>que_out_24_0_4, q_0_3=>que_out_24_0_3, q_0_2=>que_out_24_0_2, 
      q_0_1=>que_out_24_0_1, q_0_0=>que_out_24_0_0, q_1_15=>que_out_24_1_15, 
      q_1_14=>que_out_24_1_14, q_1_13=>que_out_24_1_13, q_1_12=>
      que_out_24_1_12, q_1_11=>que_out_24_1_11, q_1_10=>que_out_24_1_10, 
      q_1_9=>que_out_24_1_9, q_1_8=>que_out_24_1_8, q_1_7=>que_out_24_1_7, 
      q_1_6=>que_out_24_1_6, q_1_5=>que_out_24_1_5, q_1_4=>que_out_24_1_4, 
      q_1_3=>que_out_24_1_3, q_1_2=>que_out_24_1_2, q_1_1=>que_out_24_1_1, 
      q_1_0=>que_out_24_1_0, q_2_15=>que_out_24_2_15, q_2_14=>
      que_out_24_2_14, q_2_13=>que_out_24_2_13, q_2_12=>que_out_24_2_12, 
      q_2_11=>que_out_24_2_11, q_2_10=>que_out_24_2_10, q_2_9=>
      que_out_24_2_9, q_2_8=>que_out_24_2_8, q_2_7=>que_out_24_2_7, q_2_6=>
      que_out_24_2_6, q_2_5=>que_out_24_2_5, q_2_4=>que_out_24_2_4, q_2_3=>
      que_out_24_2_3, q_2_2=>que_out_24_2_2, q_2_1=>que_out_24_2_1, q_2_0=>
      que_out_24_2_0, q_3_15=>que_out_24_3_15, q_3_14=>que_out_24_3_14, 
      q_3_13=>que_out_24_3_13, q_3_12=>que_out_24_3_12, q_3_11=>
      que_out_24_3_11, q_3_10=>que_out_24_3_10, q_3_9=>que_out_24_3_9, q_3_8
      =>que_out_24_3_8, q_3_7=>que_out_24_3_7, q_3_6=>que_out_24_3_6, q_3_5
      =>que_out_24_3_5, q_3_4=>que_out_24_3_4, q_3_3=>que_out_24_3_3, q_3_2
      =>que_out_24_3_2, q_3_1=>que_out_24_3_1, q_3_0=>que_out_24_3_0, q_4_15
      =>que_out_24_4_15, q_4_14=>que_out_24_4_14, q_4_13=>que_out_24_4_13, 
      q_4_12=>que_out_24_4_12, q_4_11=>que_out_24_4_11, q_4_10=>
      que_out_24_4_10, q_4_9=>que_out_24_4_9, q_4_8=>que_out_24_4_8, q_4_7=>
      que_out_24_4_7, q_4_6=>que_out_24_4_6, q_4_5=>que_out_24_4_5, q_4_4=>
      que_out_24_4_4, q_4_3=>que_out_24_4_3, q_4_2=>que_out_24_4_2, q_4_1=>
      que_out_24_4_1, q_4_0=>que_out_24_4_0, clk=>nx10734, load=>sel_que_24, 
      reset=>nx10710);
   gen_queues_25_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_25_0_15, q_0_14=>que_out_25_0_14, q_0_13=>
      que_out_25_0_13, q_0_12=>que_out_25_0_12, q_0_11=>que_out_25_0_11, 
      q_0_10=>que_out_25_0_10, q_0_9=>que_out_25_0_9, q_0_8=>que_out_25_0_8, 
      q_0_7=>que_out_25_0_7, q_0_6=>que_out_25_0_6, q_0_5=>que_out_25_0_5, 
      q_0_4=>que_out_25_0_4, q_0_3=>que_out_25_0_3, q_0_2=>que_out_25_0_2, 
      q_0_1=>que_out_25_0_1, q_0_0=>que_out_25_0_0, q_1_15=>que_out_25_1_15, 
      q_1_14=>que_out_25_1_14, q_1_13=>que_out_25_1_13, q_1_12=>
      que_out_25_1_12, q_1_11=>que_out_25_1_11, q_1_10=>que_out_25_1_10, 
      q_1_9=>que_out_25_1_9, q_1_8=>que_out_25_1_8, q_1_7=>que_out_25_1_7, 
      q_1_6=>que_out_25_1_6, q_1_5=>que_out_25_1_5, q_1_4=>que_out_25_1_4, 
      q_1_3=>que_out_25_1_3, q_1_2=>que_out_25_1_2, q_1_1=>que_out_25_1_1, 
      q_1_0=>que_out_25_1_0, q_2_15=>que_out_25_2_15, q_2_14=>
      que_out_25_2_14, q_2_13=>que_out_25_2_13, q_2_12=>que_out_25_2_12, 
      q_2_11=>que_out_25_2_11, q_2_10=>que_out_25_2_10, q_2_9=>
      que_out_25_2_9, q_2_8=>que_out_25_2_8, q_2_7=>que_out_25_2_7, q_2_6=>
      que_out_25_2_6, q_2_5=>que_out_25_2_5, q_2_4=>que_out_25_2_4, q_2_3=>
      que_out_25_2_3, q_2_2=>que_out_25_2_2, q_2_1=>que_out_25_2_1, q_2_0=>
      que_out_25_2_0, q_3_15=>que_out_25_3_15, q_3_14=>que_out_25_3_14, 
      q_3_13=>que_out_25_3_13, q_3_12=>que_out_25_3_12, q_3_11=>
      que_out_25_3_11, q_3_10=>que_out_25_3_10, q_3_9=>que_out_25_3_9, q_3_8
      =>que_out_25_3_8, q_3_7=>que_out_25_3_7, q_3_6=>que_out_25_3_6, q_3_5
      =>que_out_25_3_5, q_3_4=>que_out_25_3_4, q_3_3=>que_out_25_3_3, q_3_2
      =>que_out_25_3_2, q_3_1=>que_out_25_3_1, q_3_0=>que_out_25_3_0, q_4_15
      =>que_out_25_4_15, q_4_14=>que_out_25_4_14, q_4_13=>que_out_25_4_13, 
      q_4_12=>que_out_25_4_12, q_4_11=>que_out_25_4_11, q_4_10=>
      que_out_25_4_10, q_4_9=>que_out_25_4_9, q_4_8=>que_out_25_4_8, q_4_7=>
      que_out_25_4_7, q_4_6=>que_out_25_4_6, q_4_5=>que_out_25_4_5, q_4_4=>
      que_out_25_4_4, q_4_3=>que_out_25_4_3, q_4_2=>que_out_25_4_2, q_4_1=>
      que_out_25_4_1, q_4_0=>que_out_25_4_0, clk=>nx10734, load=>sel_que_25, 
      reset=>nx10710);
   gen_queues_26_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_26_0_15, q_0_14=>que_out_26_0_14, q_0_13=>
      que_out_26_0_13, q_0_12=>que_out_26_0_12, q_0_11=>que_out_26_0_11, 
      q_0_10=>que_out_26_0_10, q_0_9=>que_out_26_0_9, q_0_8=>que_out_26_0_8, 
      q_0_7=>que_out_26_0_7, q_0_6=>que_out_26_0_6, q_0_5=>que_out_26_0_5, 
      q_0_4=>que_out_26_0_4, q_0_3=>que_out_26_0_3, q_0_2=>que_out_26_0_2, 
      q_0_1=>que_out_26_0_1, q_0_0=>que_out_26_0_0, q_1_15=>que_out_26_1_15, 
      q_1_14=>que_out_26_1_14, q_1_13=>que_out_26_1_13, q_1_12=>
      que_out_26_1_12, q_1_11=>que_out_26_1_11, q_1_10=>que_out_26_1_10, 
      q_1_9=>que_out_26_1_9, q_1_8=>que_out_26_1_8, q_1_7=>que_out_26_1_7, 
      q_1_6=>que_out_26_1_6, q_1_5=>que_out_26_1_5, q_1_4=>que_out_26_1_4, 
      q_1_3=>que_out_26_1_3, q_1_2=>que_out_26_1_2, q_1_1=>que_out_26_1_1, 
      q_1_0=>que_out_26_1_0, q_2_15=>que_out_26_2_15, q_2_14=>
      que_out_26_2_14, q_2_13=>que_out_26_2_13, q_2_12=>que_out_26_2_12, 
      q_2_11=>que_out_26_2_11, q_2_10=>que_out_26_2_10, q_2_9=>
      que_out_26_2_9, q_2_8=>que_out_26_2_8, q_2_7=>que_out_26_2_7, q_2_6=>
      que_out_26_2_6, q_2_5=>que_out_26_2_5, q_2_4=>que_out_26_2_4, q_2_3=>
      que_out_26_2_3, q_2_2=>que_out_26_2_2, q_2_1=>que_out_26_2_1, q_2_0=>
      que_out_26_2_0, q_3_15=>que_out_26_3_15, q_3_14=>que_out_26_3_14, 
      q_3_13=>que_out_26_3_13, q_3_12=>que_out_26_3_12, q_3_11=>
      que_out_26_3_11, q_3_10=>que_out_26_3_10, q_3_9=>que_out_26_3_9, q_3_8
      =>que_out_26_3_8, q_3_7=>que_out_26_3_7, q_3_6=>que_out_26_3_6, q_3_5
      =>que_out_26_3_5, q_3_4=>que_out_26_3_4, q_3_3=>que_out_26_3_3, q_3_2
      =>que_out_26_3_2, q_3_1=>que_out_26_3_1, q_3_0=>que_out_26_3_0, q_4_15
      =>que_out_26_4_15, q_4_14=>que_out_26_4_14, q_4_13=>que_out_26_4_13, 
      q_4_12=>que_out_26_4_12, q_4_11=>que_out_26_4_11, q_4_10=>
      que_out_26_4_10, q_4_9=>que_out_26_4_9, q_4_8=>que_out_26_4_8, q_4_7=>
      que_out_26_4_7, q_4_6=>que_out_26_4_6, q_4_5=>que_out_26_4_5, q_4_4=>
      que_out_26_4_4, q_4_3=>que_out_26_4_3, q_4_2=>que_out_26_4_2, q_4_1=>
      que_out_26_4_1, q_4_0=>que_out_26_4_0, clk=>nx10734, load=>sel_que_26, 
      reset=>nx10710);
   gen_queues_27_que : Queue_5 port map ( d(15)=>nx10518, d(14)=>nx10528, 
      d(13)=>nx10538, d(12)=>nx10548, d(11)=>nx10558, d(10)=>nx10568, d(9)=>
      nx10578, d(8)=>nx10588, d(7)=>nx10598, d(6)=>nx10608, d(5)=>nx10618, 
      d(4)=>nx10628, d(3)=>nx10638, d(2)=>nx10648, d(1)=>nx10658, d(0)=>
      nx10668, q_0_15=>que_out_27_0_15, q_0_14=>que_out_27_0_14, q_0_13=>
      que_out_27_0_13, q_0_12=>que_out_27_0_12, q_0_11=>que_out_27_0_11, 
      q_0_10=>que_out_27_0_10, q_0_9=>que_out_27_0_9, q_0_8=>que_out_27_0_8, 
      q_0_7=>que_out_27_0_7, q_0_6=>que_out_27_0_6, q_0_5=>que_out_27_0_5, 
      q_0_4=>que_out_27_0_4, q_0_3=>que_out_27_0_3, q_0_2=>que_out_27_0_2, 
      q_0_1=>que_out_27_0_1, q_0_0=>que_out_27_0_0, q_1_15=>que_out_27_1_15, 
      q_1_14=>que_out_27_1_14, q_1_13=>que_out_27_1_13, q_1_12=>
      que_out_27_1_12, q_1_11=>que_out_27_1_11, q_1_10=>que_out_27_1_10, 
      q_1_9=>que_out_27_1_9, q_1_8=>que_out_27_1_8, q_1_7=>que_out_27_1_7, 
      q_1_6=>que_out_27_1_6, q_1_5=>que_out_27_1_5, q_1_4=>que_out_27_1_4, 
      q_1_3=>que_out_27_1_3, q_1_2=>que_out_27_1_2, q_1_1=>que_out_27_1_1, 
      q_1_0=>que_out_27_1_0, q_2_15=>que_out_27_2_15, q_2_14=>
      que_out_27_2_14, q_2_13=>que_out_27_2_13, q_2_12=>que_out_27_2_12, 
      q_2_11=>que_out_27_2_11, q_2_10=>que_out_27_2_10, q_2_9=>
      que_out_27_2_9, q_2_8=>que_out_27_2_8, q_2_7=>que_out_27_2_7, q_2_6=>
      que_out_27_2_6, q_2_5=>que_out_27_2_5, q_2_4=>que_out_27_2_4, q_2_3=>
      que_out_27_2_3, q_2_2=>que_out_27_2_2, q_2_1=>que_out_27_2_1, q_2_0=>
      que_out_27_2_0, q_3_15=>que_out_27_3_15, q_3_14=>que_out_27_3_14, 
      q_3_13=>que_out_27_3_13, q_3_12=>que_out_27_3_12, q_3_11=>
      que_out_27_3_11, q_3_10=>que_out_27_3_10, q_3_9=>que_out_27_3_9, q_3_8
      =>que_out_27_3_8, q_3_7=>que_out_27_3_7, q_3_6=>que_out_27_3_6, q_3_5
      =>que_out_27_3_5, q_3_4=>que_out_27_3_4, q_3_3=>que_out_27_3_3, q_3_2
      =>que_out_27_3_2, q_3_1=>que_out_27_3_1, q_3_0=>que_out_27_3_0, q_4_15
      =>que_out_27_4_15, q_4_14=>que_out_27_4_14, q_4_13=>que_out_27_4_13, 
      q_4_12=>que_out_27_4_12, q_4_11=>que_out_27_4_11, q_4_10=>
      que_out_27_4_10, q_4_9=>que_out_27_4_9, q_4_8=>que_out_27_4_8, q_4_7=>
      que_out_27_4_7, q_4_6=>que_out_27_4_6, q_4_5=>que_out_27_4_5, q_4_4=>
      que_out_27_4_4, q_4_3=>que_out_27_4_3, q_4_2=>que_out_27_4_2, q_4_1=>
      que_out_27_4_1, q_4_0=>que_out_27_4_0, clk=>nx10736, load=>sel_que_27, 
      reset=>nx10712);
   ix6830 : nand03 port map ( Y=>nx6829, A0=>nx8938, A1=>nx6833, A2=>nx6835
   );
   ix8939 : nor02ii port map ( Y=>nx8938, A0=>cache_in_sel(4), A1=>
      decoder_enable);
   ix6834 : inv01 port map ( Y=>nx6833, A=>cache_in_sel(1));
   ix6836 : inv01 port map ( Y=>nx6835, A=>cache_in_sel(0));
   ix6840 : nand03 port map ( Y=>nx6839, A0=>nx8938, A1=>nx6833, A2=>nx10508
   );
   ix6844 : nand03 port map ( Y=>nx6843, A0=>nx8938, A1=>nx10506, A2=>nx6835
   );
   ix6848 : nand03 port map ( Y=>nx6847, A0=>nx8938, A1=>nx10506, A2=>
      nx10508);
   ix9023 : nor02_2x port map ( Y=>sel_que_12, A0=>nx6875, A1=>nx6829);
   ix6876 : nand02 port map ( Y=>nx6875, A0=>cache_in_sel(3), A1=>
      cache_in_sel(2));
   ix9025 : nor02_2x port map ( Y=>sel_que_13, A0=>nx6875, A1=>nx6839);
   ix9027 : nor02_2x port map ( Y=>sel_que_14, A0=>nx6843, A1=>nx6875);
   ix9029 : nor02_2x port map ( Y=>sel_que_15, A0=>nx6875, A1=>nx6847);
   ix9043 : and02 port map ( Y=>sel_que_16, A0=>nx6885, A1=>nx9038);
   ix6886 : nor02_2x port map ( Y=>nx6885, A0=>cache_in_sel(2), A1=>
      cache_in_sel(3));
   ix9039 : nor03_2x port map ( Y=>nx9038, A0=>nx6889, A1=>nx10506, A2=>
      nx10508);
   ix6890 : nand02 port map ( Y=>nx6889, A0=>cache_in_sel(4), A1=>
      decoder_enable);
   ix6894 : nand04 port map ( Y=>nx6893, A0=>cache_in_sel(4), A1=>
      decoder_enable, A2=>nx6833, A3=>nx10508);
   ix6898 : nand04 port map ( Y=>nx6897, A0=>cache_in_sel(4), A1=>
      decoder_enable, A2=>nx10506, A3=>nx6835);
   ix6902 : nand04 port map ( Y=>nx6901, A0=>cache_in_sel(4), A1=>
      decoder_enable, A2=>nx10506, A3=>nx10508);
   ix9075 : and02 port map ( Y=>sel_que_20, A0=>nx6905, A1=>nx9038);
   ix9091 : and02 port map ( Y=>sel_que_24, A0=>nx6915, A1=>nx9038);
   ix243 : or04 port map ( Y=>out_column_4_0, A0=>nx238, A1=>nx188, A2=>
      nx130, A3=>nx82);
   ix239 : nand03 port map ( Y=>nx238, A0=>nx6927, A1=>nx6951, A2=>nx6967);
   ix6928 : aoi222 port map ( Y=>nx6927, A0=>que_out_10_4_0, A1=>nx10298, B0
      =>que_out_6_4_0, B1=>nx10350, C0=>que_out_9_4_0, C1=>nx10324);
   ix6932 : nand02_2x port map ( Y=>nx6931, A0=>cache_out_sel(3), A1=>nx6933
   );
   ix6934 : inv01 port map ( Y=>nx6933, A=>cache_out_sel(0));
   ix6938 : inv01 port map ( Y=>nx6937, A=>cache_out_sel(4));
   ix6940 : inv02 port map ( Y=>nx6939, A=>cache_out_sel(2));
   ix6946 : nand03 port map ( Y=>nx6945, A0=>nx10502, A1=>nx6937, A2=>
      nx10498);
   ix227 : nor04 port map ( Y=>nx226, A0=>nx6949, A1=>nx10502, A2=>nx10494, 
      A3=>nx10498);
   ix6950 : nand02_2x port map ( Y=>nx6949, A0=>cache_out_sel(3), A1=>
      cache_out_sel(0));
   ix6952 : aoi22 port map ( Y=>nx6951, A0=>que_out_5_4_0, A1=>nx10246, B0=>
      que_out_18_4_0, B1=>nx10272);
   ix6956 : nand02 port map ( Y=>nx6955, A0=>nx6957, A1=>cache_out_sel(0));
   ix6958 : inv01 port map ( Y=>nx6957, A=>cache_out_sel(3));
   ix6962 : inv01 port map ( Y=>nx6961, A=>cache_out_sel(1));
   ix215 : nor03_2x port map ( Y=>nx214, A0=>nx6965, A1=>nx10498, A2=>nx6943
   );
   ix6966 : nand02_2x port map ( Y=>nx6965, A0=>nx10494, A1=>nx10504);
   ix6968 : aoi22 port map ( Y=>nx6967, A0=>que_out_17_4_0, A1=>nx10220, B0
      =>que_out_20_4_0, B1=>nx10194);
   ix201 : nor03_2x port map ( Y=>nx200, A0=>nx6971, A1=>nx10498, A2=>
      nx10374);
   ix6972 : nand02_2x port map ( Y=>nx6971, A0=>nx10496, A1=>nx6961);
   ix193 : nor03_2x port map ( Y=>nx192, A0=>nx6971, A1=>nx6939, A2=>nx6943
   );
   ix189 : nand03 port map ( Y=>nx188, A0=>nx6977, A1=>nx6985, A2=>nx6991);
   ix6978 : aoi222 port map ( Y=>nx6977, A0=>que_out_19_4_0, A1=>nx10168, B0
      =>que_out_21_4_0, B1=>nx10142, C0=>que_out_8_4_0, C1=>nx10116);
   ix181 : nor03_2x port map ( Y=>nx180, A0=>nx6965, A1=>nx10498, A2=>
      nx10374);
   ix173 : nor03_2x port map ( Y=>nx172, A0=>nx6971, A1=>nx6939, A2=>nx10374
   );
   ix167 : nor04 port map ( Y=>nx166, A0=>nx6931, A1=>nx10502, A2=>nx10494, 
      A3=>nx10498);
   ix6986 : aoi22 port map ( Y=>nx6985, A0=>que_out_25_4_0, A1=>nx10064, B0
      =>que_out_16_4_0, B1=>nx10090);
   ix151 : nor02_2x port map ( Y=>nx150, A0=>nx6949, A1=>nx6971);
   ix159 : nor03_2x port map ( Y=>nx158, A0=>nx6971, A1=>nx10498, A2=>nx6943
   );
   ix6992 : aoi22 port map ( Y=>nx6991, A0=>que_out_24_4_0, A1=>nx10038, B0
      =>que_out_22_4_0, B1=>nx10012);
   ix145 : nor02_2x port map ( Y=>nx144, A0=>nx6971, A1=>nx6931);
   ix137 : nor03_2x port map ( Y=>nx136, A0=>nx6965, A1=>nx6939, A2=>nx6943
   );
   ix131 : nand03 port map ( Y=>nx130, A0=>nx6999, A1=>nx7007, A2=>nx7017);
   ix7000 : aoi222 port map ( Y=>nx6999, A0=>que_out_15_4_0, A1=>nx9960, B0
      =>que_out_3_4_0, B1=>nx9986, C0=>que_out_23_4_0, C1=>nx9934);
   ix119 : nor02_2x port map ( Y=>nx118, A0=>nx6949, A1=>nx6945);
   ix115 : nor03_2x port map ( Y=>nx114, A0=>nx6965, A1=>nx6939, A2=>nx10374
   );
   ix7008 : aoi22 port map ( Y=>nx7007, A0=>que_out_27_4_0, A1=>nx9908, B0=>
      que_out_4_4_0, B1=>nx9882);
   ix105 : nor02_2x port map ( Y=>nx104, A0=>nx6949, A1=>nx6965);
   ix101 : and02 port map ( Y=>nx100, A0=>nx88, A1=>nx28);
   ix89 : nor02_2x port map ( Y=>nx88, A0=>cache_out_sel(3), A1=>
      cache_out_sel(0));
   ix29 : nor03_2x port map ( Y=>nx28, A0=>nx10502, A1=>nx10494, A2=>nx6939
   );
   ix7018 : aoi22 port map ( Y=>nx7017, A0=>que_out_0_4_0, A1=>nx9830, B0=>
      que_out_2_4_0, B1=>nx9856);
   ix91 : and02 port map ( Y=>nx90, A0=>nx88, A1=>nx12);
   ix13 : nor03_2x port map ( Y=>nx12, A0=>nx10504, A1=>nx10494, A2=>nx10500
   );
   ix95 : and02 port map ( Y=>nx94, A0=>nx88, A1=>nx62);
   ix63 : nor03_2x port map ( Y=>nx62, A0=>nx6961, A1=>nx10494, A2=>nx10500
   );
   ix83 : nand03 port map ( Y=>nx82, A0=>nx7029, A1=>nx7037, A2=>nx7043);
   ix7030 : aoi222 port map ( Y=>nx7029, A0=>que_out_26_4_0, A1=>nx9804, B0
      =>que_out_14_4_0, B1=>nx9778, C0=>que_out_11_4_0, C1=>nx9752);
   ix75 : nor02_2x port map ( Y=>nx74, A0=>nx6965, A1=>nx6931);
   ix69 : nor02_2x port map ( Y=>nx68, A0=>nx6931, A1=>nx6945);
   ix7038 : aoi22 port map ( Y=>nx7037, A0=>que_out_13_4_0, A1=>nx9726, B0=>
      que_out_7_4_0, B1=>nx9700);
   ix43 : nor02_2x port map ( Y=>nx42, A0=>nx10374, A1=>nx6945);
   ix7044 : aoi22 port map ( Y=>nx7043, A0=>que_out_12_4_0, A1=>nx9674, B0=>
      que_out_1_4_0, B1=>nx9648);
   ix15 : nor04 port map ( Y=>nx14, A0=>nx10376, A1=>nx10504, A2=>nx10494, 
      A3=>nx10500);
   ix353 : or04 port map ( Y=>out_column_4_1, A0=>nx348, A1=>nx322, A2=>
      nx294, A3=>nx268);
   ix349 : nand03 port map ( Y=>nx348, A0=>nx7053, A1=>nx7055, A2=>nx7057);
   ix7054 : aoi222 port map ( Y=>nx7053, A0=>que_out_10_4_1, A1=>nx10298, B0
      =>que_out_6_4_1, B1=>nx10350, C0=>que_out_9_4_1, C1=>nx10324);
   ix7056 : aoi22 port map ( Y=>nx7055, A0=>que_out_5_4_1, A1=>nx10246, B0=>
      que_out_18_4_1, B1=>nx10272);
   ix7058 : aoi22 port map ( Y=>nx7057, A0=>que_out_17_4_1, A1=>nx10220, B0
      =>que_out_20_4_1, B1=>nx10194);
   ix323 : nand03 port map ( Y=>nx322, A0=>nx7061, A1=>nx7063, A2=>nx7065);
   ix7062 : aoi222 port map ( Y=>nx7061, A0=>que_out_19_4_1, A1=>nx10168, B0
      =>que_out_21_4_1, B1=>nx10142, C0=>que_out_8_4_1, C1=>nx10116);
   ix7064 : aoi22 port map ( Y=>nx7063, A0=>que_out_25_4_1, A1=>nx10064, B0
      =>que_out_16_4_1, B1=>nx10090);
   ix7066 : aoi22 port map ( Y=>nx7065, A0=>que_out_24_4_1, A1=>nx10038, B0
      =>que_out_22_4_1, B1=>nx10012);
   ix295 : nand03 port map ( Y=>nx294, A0=>nx7069, A1=>nx7071, A2=>nx7073);
   ix7070 : aoi222 port map ( Y=>nx7069, A0=>que_out_15_4_1, A1=>nx9960, B0
      =>que_out_3_4_1, B1=>nx9986, C0=>que_out_23_4_1, C1=>nx9934);
   ix7072 : aoi22 port map ( Y=>nx7071, A0=>que_out_27_4_1, A1=>nx9908, B0=>
      que_out_4_4_1, B1=>nx9882);
   ix7074 : aoi22 port map ( Y=>nx7073, A0=>que_out_0_4_1, A1=>nx9830, B0=>
      que_out_2_4_1, B1=>nx9856);
   ix269 : nand03 port map ( Y=>nx268, A0=>nx7077, A1=>nx7079, A2=>nx7081);
   ix7078 : aoi222 port map ( Y=>nx7077, A0=>que_out_26_4_1, A1=>nx9804, B0
      =>que_out_14_4_1, B1=>nx9778, C0=>que_out_11_4_1, C1=>nx9752);
   ix7080 : aoi22 port map ( Y=>nx7079, A0=>que_out_13_4_1, A1=>nx9726, B0=>
      que_out_7_4_1, B1=>nx9700);
   ix7082 : aoi22 port map ( Y=>nx7081, A0=>que_out_12_4_1, A1=>nx9674, B0=>
      que_out_1_4_1, B1=>nx9648);
   ix463 : or04 port map ( Y=>out_column_4_2, A0=>nx458, A1=>nx432, A2=>
      nx404, A3=>nx378);
   ix459 : nand03 port map ( Y=>nx458, A0=>nx7087, A1=>nx7089, A2=>nx7091);
   ix7088 : aoi222 port map ( Y=>nx7087, A0=>que_out_10_4_2, A1=>nx10298, B0
      =>que_out_6_4_2, B1=>nx10350, C0=>que_out_9_4_2, C1=>nx10324);
   ix7090 : aoi22 port map ( Y=>nx7089, A0=>que_out_5_4_2, A1=>nx10246, B0=>
      que_out_18_4_2, B1=>nx10272);
   ix7092 : aoi22 port map ( Y=>nx7091, A0=>que_out_17_4_2, A1=>nx10220, B0
      =>que_out_20_4_2, B1=>nx10194);
   ix433 : nand03 port map ( Y=>nx432, A0=>nx7095, A1=>nx7097, A2=>nx7099);
   ix7096 : aoi222 port map ( Y=>nx7095, A0=>que_out_19_4_2, A1=>nx10168, B0
      =>que_out_21_4_2, B1=>nx10142, C0=>que_out_8_4_2, C1=>nx10116);
   ix7098 : aoi22 port map ( Y=>nx7097, A0=>que_out_25_4_2, A1=>nx10064, B0
      =>que_out_16_4_2, B1=>nx10090);
   ix7100 : aoi22 port map ( Y=>nx7099, A0=>que_out_24_4_2, A1=>nx10038, B0
      =>que_out_22_4_2, B1=>nx10012);
   ix405 : nand03 port map ( Y=>nx404, A0=>nx7103, A1=>nx7105, A2=>nx7107);
   ix7104 : aoi222 port map ( Y=>nx7103, A0=>que_out_15_4_2, A1=>nx9960, B0
      =>que_out_3_4_2, B1=>nx9986, C0=>que_out_23_4_2, C1=>nx9934);
   ix7106 : aoi22 port map ( Y=>nx7105, A0=>que_out_27_4_2, A1=>nx9908, B0=>
      que_out_4_4_2, B1=>nx9882);
   ix7108 : aoi22 port map ( Y=>nx7107, A0=>que_out_0_4_2, A1=>nx9830, B0=>
      que_out_2_4_2, B1=>nx9856);
   ix379 : nand03 port map ( Y=>nx378, A0=>nx7111, A1=>nx7113, A2=>nx7115);
   ix7112 : aoi222 port map ( Y=>nx7111, A0=>que_out_26_4_2, A1=>nx9804, B0
      =>que_out_14_4_2, B1=>nx9778, C0=>que_out_11_4_2, C1=>nx9752);
   ix7114 : aoi22 port map ( Y=>nx7113, A0=>que_out_13_4_2, A1=>nx9726, B0=>
      que_out_7_4_2, B1=>nx9700);
   ix7116 : aoi22 port map ( Y=>nx7115, A0=>que_out_12_4_2, A1=>nx9674, B0=>
      que_out_1_4_2, B1=>nx9648);
   ix573 : or04 port map ( Y=>out_column_4_3, A0=>nx568, A1=>nx542, A2=>
      nx514, A3=>nx488);
   ix569 : nand03 port map ( Y=>nx568, A0=>nx7121, A1=>nx7123, A2=>nx7125);
   ix7122 : aoi222 port map ( Y=>nx7121, A0=>que_out_10_4_3, A1=>nx10298, B0
      =>que_out_6_4_3, B1=>nx10350, C0=>que_out_9_4_3, C1=>nx10324);
   ix7124 : aoi22 port map ( Y=>nx7123, A0=>que_out_5_4_3, A1=>nx10246, B0=>
      que_out_18_4_3, B1=>nx10272);
   ix7126 : aoi22 port map ( Y=>nx7125, A0=>que_out_17_4_3, A1=>nx10220, B0
      =>que_out_20_4_3, B1=>nx10194);
   ix543 : nand03 port map ( Y=>nx542, A0=>nx7129, A1=>nx7131, A2=>nx7133);
   ix7130 : aoi222 port map ( Y=>nx7129, A0=>que_out_19_4_3, A1=>nx10168, B0
      =>que_out_21_4_3, B1=>nx10142, C0=>que_out_8_4_3, C1=>nx10116);
   ix7132 : aoi22 port map ( Y=>nx7131, A0=>que_out_25_4_3, A1=>nx10064, B0
      =>que_out_16_4_3, B1=>nx10090);
   ix7134 : aoi22 port map ( Y=>nx7133, A0=>que_out_24_4_3, A1=>nx10038, B0
      =>que_out_22_4_3, B1=>nx10012);
   ix515 : nand03 port map ( Y=>nx514, A0=>nx7137, A1=>nx7139, A2=>nx7141);
   ix7138 : aoi222 port map ( Y=>nx7137, A0=>que_out_15_4_3, A1=>nx9960, B0
      =>que_out_3_4_3, B1=>nx9986, C0=>que_out_23_4_3, C1=>nx9934);
   ix7140 : aoi22 port map ( Y=>nx7139, A0=>que_out_27_4_3, A1=>nx9908, B0=>
      que_out_4_4_3, B1=>nx9882);
   ix7142 : aoi22 port map ( Y=>nx7141, A0=>que_out_0_4_3, A1=>nx9830, B0=>
      que_out_2_4_3, B1=>nx9856);
   ix489 : nand03 port map ( Y=>nx488, A0=>nx7145, A1=>nx7147, A2=>nx7149);
   ix7146 : aoi222 port map ( Y=>nx7145, A0=>que_out_26_4_3, A1=>nx9804, B0
      =>que_out_14_4_3, B1=>nx9778, C0=>que_out_11_4_3, C1=>nx9752);
   ix7148 : aoi22 port map ( Y=>nx7147, A0=>que_out_13_4_3, A1=>nx9726, B0=>
      que_out_7_4_3, B1=>nx9700);
   ix7150 : aoi22 port map ( Y=>nx7149, A0=>que_out_12_4_3, A1=>nx9674, B0=>
      que_out_1_4_3, B1=>nx9648);
   ix683 : or04 port map ( Y=>out_column_4_4, A0=>nx678, A1=>nx652, A2=>
      nx624, A3=>nx598);
   ix679 : nand03 port map ( Y=>nx678, A0=>nx7155, A1=>nx7157, A2=>nx7159);
   ix7156 : aoi222 port map ( Y=>nx7155, A0=>que_out_10_4_4, A1=>nx10298, B0
      =>que_out_6_4_4, B1=>nx10350, C0=>que_out_9_4_4, C1=>nx10324);
   ix7158 : aoi22 port map ( Y=>nx7157, A0=>que_out_5_4_4, A1=>nx10246, B0=>
      que_out_18_4_4, B1=>nx10272);
   ix7160 : aoi22 port map ( Y=>nx7159, A0=>que_out_17_4_4, A1=>nx10220, B0
      =>que_out_20_4_4, B1=>nx10194);
   ix653 : nand03 port map ( Y=>nx652, A0=>nx7163, A1=>nx7165, A2=>nx7167);
   ix7164 : aoi222 port map ( Y=>nx7163, A0=>que_out_19_4_4, A1=>nx10168, B0
      =>que_out_21_4_4, B1=>nx10142, C0=>que_out_8_4_4, C1=>nx10116);
   ix7166 : aoi22 port map ( Y=>nx7165, A0=>que_out_25_4_4, A1=>nx10064, B0
      =>que_out_16_4_4, B1=>nx10090);
   ix7168 : aoi22 port map ( Y=>nx7167, A0=>que_out_24_4_4, A1=>nx10038, B0
      =>que_out_22_4_4, B1=>nx10012);
   ix625 : nand03 port map ( Y=>nx624, A0=>nx7171, A1=>nx7173, A2=>nx7175);
   ix7172 : aoi222 port map ( Y=>nx7171, A0=>que_out_15_4_4, A1=>nx9960, B0
      =>que_out_3_4_4, B1=>nx9986, C0=>que_out_23_4_4, C1=>nx9934);
   ix7174 : aoi22 port map ( Y=>nx7173, A0=>que_out_27_4_4, A1=>nx9908, B0=>
      que_out_4_4_4, B1=>nx9882);
   ix7176 : aoi22 port map ( Y=>nx7175, A0=>que_out_0_4_4, A1=>nx9830, B0=>
      que_out_2_4_4, B1=>nx9856);
   ix599 : nand03 port map ( Y=>nx598, A0=>nx7179, A1=>nx7181, A2=>nx7183);
   ix7180 : aoi222 port map ( Y=>nx7179, A0=>que_out_26_4_4, A1=>nx9804, B0
      =>que_out_14_4_4, B1=>nx9778, C0=>que_out_11_4_4, C1=>nx9752);
   ix7182 : aoi22 port map ( Y=>nx7181, A0=>que_out_13_4_4, A1=>nx9726, B0=>
      que_out_7_4_4, B1=>nx9700);
   ix7184 : aoi22 port map ( Y=>nx7183, A0=>que_out_12_4_4, A1=>nx9674, B0=>
      que_out_1_4_4, B1=>nx9648);
   ix793 : or04 port map ( Y=>out_column_4_5, A0=>nx788, A1=>nx762, A2=>
      nx734, A3=>nx708);
   ix789 : nand03 port map ( Y=>nx788, A0=>nx7189, A1=>nx7191, A2=>nx7193);
   ix7190 : aoi222 port map ( Y=>nx7189, A0=>que_out_10_4_5, A1=>nx10298, B0
      =>que_out_6_4_5, B1=>nx10350, C0=>que_out_9_4_5, C1=>nx10324);
   ix7192 : aoi22 port map ( Y=>nx7191, A0=>que_out_5_4_5, A1=>nx10246, B0=>
      que_out_18_4_5, B1=>nx10272);
   ix7194 : aoi22 port map ( Y=>nx7193, A0=>que_out_17_4_5, A1=>nx10220, B0
      =>que_out_20_4_5, B1=>nx10194);
   ix763 : nand03 port map ( Y=>nx762, A0=>nx7197, A1=>nx7199, A2=>nx7201);
   ix7198 : aoi222 port map ( Y=>nx7197, A0=>que_out_19_4_5, A1=>nx10168, B0
      =>que_out_21_4_5, B1=>nx10142, C0=>que_out_8_4_5, C1=>nx10116);
   ix7200 : aoi22 port map ( Y=>nx7199, A0=>que_out_25_4_5, A1=>nx10064, B0
      =>que_out_16_4_5, B1=>nx10090);
   ix7202 : aoi22 port map ( Y=>nx7201, A0=>que_out_24_4_5, A1=>nx10038, B0
      =>que_out_22_4_5, B1=>nx10012);
   ix735 : nand03 port map ( Y=>nx734, A0=>nx7205, A1=>nx7207, A2=>nx7209);
   ix7206 : aoi222 port map ( Y=>nx7205, A0=>que_out_15_4_5, A1=>nx9960, B0
      =>que_out_3_4_5, B1=>nx9986, C0=>que_out_23_4_5, C1=>nx9934);
   ix7208 : aoi22 port map ( Y=>nx7207, A0=>que_out_27_4_5, A1=>nx9908, B0=>
      que_out_4_4_5, B1=>nx9882);
   ix7210 : aoi22 port map ( Y=>nx7209, A0=>que_out_0_4_5, A1=>nx9830, B0=>
      que_out_2_4_5, B1=>nx9856);
   ix709 : nand03 port map ( Y=>nx708, A0=>nx7213, A1=>nx7215, A2=>nx7217);
   ix7214 : aoi222 port map ( Y=>nx7213, A0=>que_out_26_4_5, A1=>nx9804, B0
      =>que_out_14_4_5, B1=>nx9778, C0=>que_out_11_4_5, C1=>nx9752);
   ix7216 : aoi22 port map ( Y=>nx7215, A0=>que_out_13_4_5, A1=>nx9726, B0=>
      que_out_7_4_5, B1=>nx9700);
   ix7218 : aoi22 port map ( Y=>nx7217, A0=>que_out_12_4_5, A1=>nx9674, B0=>
      que_out_1_4_5, B1=>nx9648);
   ix903 : or04 port map ( Y=>out_column_4_6, A0=>nx898, A1=>nx872, A2=>
      nx844, A3=>nx818);
   ix899 : nand03 port map ( Y=>nx898, A0=>nx7223, A1=>nx7225, A2=>nx7227);
   ix7224 : aoi222 port map ( Y=>nx7223, A0=>que_out_10_4_6, A1=>nx10298, B0
      =>que_out_6_4_6, B1=>nx10350, C0=>que_out_9_4_6, C1=>nx10324);
   ix7226 : aoi22 port map ( Y=>nx7225, A0=>que_out_5_4_6, A1=>nx10246, B0=>
      que_out_18_4_6, B1=>nx10272);
   ix7228 : aoi22 port map ( Y=>nx7227, A0=>que_out_17_4_6, A1=>nx10220, B0
      =>que_out_20_4_6, B1=>nx10194);
   ix873 : nand03 port map ( Y=>nx872, A0=>nx7231, A1=>nx7233, A2=>nx7235);
   ix7232 : aoi222 port map ( Y=>nx7231, A0=>que_out_19_4_6, A1=>nx10168, B0
      =>que_out_21_4_6, B1=>nx10142, C0=>que_out_8_4_6, C1=>nx10116);
   ix7234 : aoi22 port map ( Y=>nx7233, A0=>que_out_25_4_6, A1=>nx10064, B0
      =>que_out_16_4_6, B1=>nx10090);
   ix7236 : aoi22 port map ( Y=>nx7235, A0=>que_out_24_4_6, A1=>nx10038, B0
      =>que_out_22_4_6, B1=>nx10012);
   ix845 : nand03 port map ( Y=>nx844, A0=>nx7239, A1=>nx7241, A2=>nx7243);
   ix7240 : aoi222 port map ( Y=>nx7239, A0=>que_out_15_4_6, A1=>nx9960, B0
      =>que_out_3_4_6, B1=>nx9986, C0=>que_out_23_4_6, C1=>nx9934);
   ix7242 : aoi22 port map ( Y=>nx7241, A0=>que_out_27_4_6, A1=>nx9908, B0=>
      que_out_4_4_6, B1=>nx9882);
   ix7244 : aoi22 port map ( Y=>nx7243, A0=>que_out_0_4_6, A1=>nx9830, B0=>
      que_out_2_4_6, B1=>nx9856);
   ix819 : nand03 port map ( Y=>nx818, A0=>nx7247, A1=>nx7249, A2=>nx7251);
   ix7248 : aoi222 port map ( Y=>nx7247, A0=>que_out_26_4_6, A1=>nx9804, B0
      =>que_out_14_4_6, B1=>nx9778, C0=>que_out_11_4_6, C1=>nx9752);
   ix7250 : aoi22 port map ( Y=>nx7249, A0=>que_out_13_4_6, A1=>nx9726, B0=>
      que_out_7_4_6, B1=>nx9700);
   ix7252 : aoi22 port map ( Y=>nx7251, A0=>que_out_12_4_6, A1=>nx9674, B0=>
      que_out_1_4_6, B1=>nx9648);
   ix1013 : or04 port map ( Y=>out_column_4_7, A0=>nx1008, A1=>nx982, A2=>
      nx954, A3=>nx928);
   ix1009 : nand03 port map ( Y=>nx1008, A0=>nx7257, A1=>nx7259, A2=>nx7261
   );
   ix7258 : aoi222 port map ( Y=>nx7257, A0=>que_out_10_4_7, A1=>nx10300, B0
      =>que_out_6_4_7, B1=>nx10352, C0=>que_out_9_4_7, C1=>nx10326);
   ix7260 : aoi22 port map ( Y=>nx7259, A0=>que_out_5_4_7, A1=>nx10248, B0=>
      que_out_18_4_7, B1=>nx10274);
   ix7262 : aoi22 port map ( Y=>nx7261, A0=>que_out_17_4_7, A1=>nx10222, B0
      =>que_out_20_4_7, B1=>nx10196);
   ix983 : nand03 port map ( Y=>nx982, A0=>nx7265, A1=>nx7267, A2=>nx7269);
   ix7266 : aoi222 port map ( Y=>nx7265, A0=>que_out_19_4_7, A1=>nx10170, B0
      =>que_out_21_4_7, B1=>nx10144, C0=>que_out_8_4_7, C1=>nx10118);
   ix7268 : aoi22 port map ( Y=>nx7267, A0=>que_out_25_4_7, A1=>nx10066, B0
      =>que_out_16_4_7, B1=>nx10092);
   ix7270 : aoi22 port map ( Y=>nx7269, A0=>que_out_24_4_7, A1=>nx10040, B0
      =>que_out_22_4_7, B1=>nx10014);
   ix955 : nand03 port map ( Y=>nx954, A0=>nx7273, A1=>nx7275, A2=>nx7277);
   ix7274 : aoi222 port map ( Y=>nx7273, A0=>que_out_15_4_7, A1=>nx9962, B0
      =>que_out_3_4_7, B1=>nx9988, C0=>que_out_23_4_7, C1=>nx9936);
   ix7276 : aoi22 port map ( Y=>nx7275, A0=>que_out_27_4_7, A1=>nx9910, B0=>
      que_out_4_4_7, B1=>nx9884);
   ix7278 : aoi22 port map ( Y=>nx7277, A0=>que_out_0_4_7, A1=>nx9832, B0=>
      que_out_2_4_7, B1=>nx9858);
   ix929 : nand03 port map ( Y=>nx928, A0=>nx7281, A1=>nx7283, A2=>nx7285);
   ix7282 : aoi222 port map ( Y=>nx7281, A0=>que_out_26_4_7, A1=>nx9806, B0
      =>que_out_14_4_7, B1=>nx9780, C0=>que_out_11_4_7, C1=>nx9754);
   ix7284 : aoi22 port map ( Y=>nx7283, A0=>que_out_13_4_7, A1=>nx9728, B0=>
      que_out_7_4_7, B1=>nx9702);
   ix7286 : aoi22 port map ( Y=>nx7285, A0=>que_out_12_4_7, A1=>nx9676, B0=>
      que_out_1_4_7, B1=>nx9650);
   ix1123 : or04 port map ( Y=>out_column_4_8, A0=>nx1118, A1=>nx1092, A2=>
      nx1064, A3=>nx1038);
   ix1119 : nand03 port map ( Y=>nx1118, A0=>nx7291, A1=>nx7293, A2=>nx7295
   );
   ix7292 : aoi222 port map ( Y=>nx7291, A0=>que_out_10_4_8, A1=>nx10300, B0
      =>que_out_6_4_8, B1=>nx10352, C0=>que_out_9_4_8, C1=>nx10326);
   ix7294 : aoi22 port map ( Y=>nx7293, A0=>que_out_5_4_8, A1=>nx10248, B0=>
      que_out_18_4_8, B1=>nx10274);
   ix7296 : aoi22 port map ( Y=>nx7295, A0=>que_out_17_4_8, A1=>nx10222, B0
      =>que_out_20_4_8, B1=>nx10196);
   ix1093 : nand03 port map ( Y=>nx1092, A0=>nx7299, A1=>nx7301, A2=>nx7303
   );
   ix7300 : aoi222 port map ( Y=>nx7299, A0=>que_out_19_4_8, A1=>nx10170, B0
      =>que_out_21_4_8, B1=>nx10144, C0=>que_out_8_4_8, C1=>nx10118);
   ix7302 : aoi22 port map ( Y=>nx7301, A0=>que_out_25_4_8, A1=>nx10066, B0
      =>que_out_16_4_8, B1=>nx10092);
   ix7304 : aoi22 port map ( Y=>nx7303, A0=>que_out_24_4_8, A1=>nx10040, B0
      =>que_out_22_4_8, B1=>nx10014);
   ix1065 : nand03 port map ( Y=>nx1064, A0=>nx7307, A1=>nx7309, A2=>nx7311
   );
   ix7308 : aoi222 port map ( Y=>nx7307, A0=>que_out_15_4_8, A1=>nx9962, B0
      =>que_out_3_4_8, B1=>nx9988, C0=>que_out_23_4_8, C1=>nx9936);
   ix7310 : aoi22 port map ( Y=>nx7309, A0=>que_out_27_4_8, A1=>nx9910, B0=>
      que_out_4_4_8, B1=>nx9884);
   ix7312 : aoi22 port map ( Y=>nx7311, A0=>que_out_0_4_8, A1=>nx9832, B0=>
      que_out_2_4_8, B1=>nx9858);
   ix1039 : nand03 port map ( Y=>nx1038, A0=>nx7315, A1=>nx7317, A2=>nx7319
   );
   ix7316 : aoi222 port map ( Y=>nx7315, A0=>que_out_26_4_8, A1=>nx9806, B0
      =>que_out_14_4_8, B1=>nx9780, C0=>que_out_11_4_8, C1=>nx9754);
   ix7318 : aoi22 port map ( Y=>nx7317, A0=>que_out_13_4_8, A1=>nx9728, B0=>
      que_out_7_4_8, B1=>nx9702);
   ix7320 : aoi22 port map ( Y=>nx7319, A0=>que_out_12_4_8, A1=>nx9676, B0=>
      que_out_1_4_8, B1=>nx9650);
   ix1233 : or04 port map ( Y=>out_column_4_9, A0=>nx1228, A1=>nx1202, A2=>
      nx1174, A3=>nx1148);
   ix1229 : nand03 port map ( Y=>nx1228, A0=>nx7325, A1=>nx7327, A2=>nx7329
   );
   ix7326 : aoi222 port map ( Y=>nx7325, A0=>que_out_10_4_9, A1=>nx10300, B0
      =>que_out_6_4_9, B1=>nx10352, C0=>que_out_9_4_9, C1=>nx10326);
   ix7328 : aoi22 port map ( Y=>nx7327, A0=>que_out_5_4_9, A1=>nx10248, B0=>
      que_out_18_4_9, B1=>nx10274);
   ix7330 : aoi22 port map ( Y=>nx7329, A0=>que_out_17_4_9, A1=>nx10222, B0
      =>que_out_20_4_9, B1=>nx10196);
   ix1203 : nand03 port map ( Y=>nx1202, A0=>nx7333, A1=>nx7335, A2=>nx7337
   );
   ix7334 : aoi222 port map ( Y=>nx7333, A0=>que_out_19_4_9, A1=>nx10170, B0
      =>que_out_21_4_9, B1=>nx10144, C0=>que_out_8_4_9, C1=>nx10118);
   ix7336 : aoi22 port map ( Y=>nx7335, A0=>que_out_25_4_9, A1=>nx10066, B0
      =>que_out_16_4_9, B1=>nx10092);
   ix7338 : aoi22 port map ( Y=>nx7337, A0=>que_out_24_4_9, A1=>nx10040, B0
      =>que_out_22_4_9, B1=>nx10014);
   ix1175 : nand03 port map ( Y=>nx1174, A0=>nx7341, A1=>nx7343, A2=>nx7345
   );
   ix7342 : aoi222 port map ( Y=>nx7341, A0=>que_out_15_4_9, A1=>nx9962, B0
      =>que_out_3_4_9, B1=>nx9988, C0=>que_out_23_4_9, C1=>nx9936);
   ix7344 : aoi22 port map ( Y=>nx7343, A0=>que_out_27_4_9, A1=>nx9910, B0=>
      que_out_4_4_9, B1=>nx9884);
   ix7346 : aoi22 port map ( Y=>nx7345, A0=>que_out_0_4_9, A1=>nx9832, B0=>
      que_out_2_4_9, B1=>nx9858);
   ix1149 : nand03 port map ( Y=>nx1148, A0=>nx7349, A1=>nx7351, A2=>nx7353
   );
   ix7350 : aoi222 port map ( Y=>nx7349, A0=>que_out_26_4_9, A1=>nx9806, B0
      =>que_out_14_4_9, B1=>nx9780, C0=>que_out_11_4_9, C1=>nx9754);
   ix7352 : aoi22 port map ( Y=>nx7351, A0=>que_out_13_4_9, A1=>nx9728, B0=>
      que_out_7_4_9, B1=>nx9702);
   ix7354 : aoi22 port map ( Y=>nx7353, A0=>que_out_12_4_9, A1=>nx9676, B0=>
      que_out_1_4_9, B1=>nx9650);
   ix1343 : or04 port map ( Y=>out_column_4_10, A0=>nx1338, A1=>nx1312, A2=>
      nx1284, A3=>nx1258);
   ix1339 : nand03 port map ( Y=>nx1338, A0=>nx7359, A1=>nx7361, A2=>nx7363
   );
   ix7360 : aoi222 port map ( Y=>nx7359, A0=>que_out_10_4_10, A1=>nx10300, 
      B0=>que_out_6_4_10, B1=>nx10352, C0=>que_out_9_4_10, C1=>nx10326);
   ix7362 : aoi22 port map ( Y=>nx7361, A0=>que_out_5_4_10, A1=>nx10248, B0
      =>que_out_18_4_10, B1=>nx10274);
   ix7364 : aoi22 port map ( Y=>nx7363, A0=>que_out_17_4_10, A1=>nx10222, B0
      =>que_out_20_4_10, B1=>nx10196);
   ix1313 : nand03 port map ( Y=>nx1312, A0=>nx7367, A1=>nx7369, A2=>nx7371
   );
   ix7368 : aoi222 port map ( Y=>nx7367, A0=>que_out_19_4_10, A1=>nx10170, 
      B0=>que_out_21_4_10, B1=>nx10144, C0=>que_out_8_4_10, C1=>nx10118);
   ix7370 : aoi22 port map ( Y=>nx7369, A0=>que_out_25_4_10, A1=>nx10066, B0
      =>que_out_16_4_10, B1=>nx10092);
   ix7372 : aoi22 port map ( Y=>nx7371, A0=>que_out_24_4_10, A1=>nx10040, B0
      =>que_out_22_4_10, B1=>nx10014);
   ix1285 : nand03 port map ( Y=>nx1284, A0=>nx7375, A1=>nx7377, A2=>nx7379
   );
   ix7376 : aoi222 port map ( Y=>nx7375, A0=>que_out_15_4_10, A1=>nx9962, B0
      =>que_out_3_4_10, B1=>nx9988, C0=>que_out_23_4_10, C1=>nx9936);
   ix7378 : aoi22 port map ( Y=>nx7377, A0=>que_out_27_4_10, A1=>nx9910, B0
      =>que_out_4_4_10, B1=>nx9884);
   ix7380 : aoi22 port map ( Y=>nx7379, A0=>que_out_0_4_10, A1=>nx9832, B0=>
      que_out_2_4_10, B1=>nx9858);
   ix1259 : nand03 port map ( Y=>nx1258, A0=>nx7383, A1=>nx7385, A2=>nx7387
   );
   ix7384 : aoi222 port map ( Y=>nx7383, A0=>que_out_26_4_10, A1=>nx9806, B0
      =>que_out_14_4_10, B1=>nx9780, C0=>que_out_11_4_10, C1=>nx9754);
   ix7386 : aoi22 port map ( Y=>nx7385, A0=>que_out_13_4_10, A1=>nx9728, B0
      =>que_out_7_4_10, B1=>nx9702);
   ix7388 : aoi22 port map ( Y=>nx7387, A0=>que_out_12_4_10, A1=>nx9676, B0
      =>que_out_1_4_10, B1=>nx9650);
   ix1453 : or04 port map ( Y=>out_column_4_11, A0=>nx1448, A1=>nx1422, A2=>
      nx1394, A3=>nx1368);
   ix1449 : nand03 port map ( Y=>nx1448, A0=>nx7393, A1=>nx7395, A2=>nx7397
   );
   ix7394 : aoi222 port map ( Y=>nx7393, A0=>que_out_10_4_11, A1=>nx10300, 
      B0=>que_out_6_4_11, B1=>nx10352, C0=>que_out_9_4_11, C1=>nx10326);
   ix7396 : aoi22 port map ( Y=>nx7395, A0=>que_out_5_4_11, A1=>nx10248, B0
      =>que_out_18_4_11, B1=>nx10274);
   ix7398 : aoi22 port map ( Y=>nx7397, A0=>que_out_17_4_11, A1=>nx10222, B0
      =>que_out_20_4_11, B1=>nx10196);
   ix1423 : nand03 port map ( Y=>nx1422, A0=>nx7401, A1=>nx7403, A2=>nx7405
   );
   ix7402 : aoi222 port map ( Y=>nx7401, A0=>que_out_19_4_11, A1=>nx10170, 
      B0=>que_out_21_4_11, B1=>nx10144, C0=>que_out_8_4_11, C1=>nx10118);
   ix7404 : aoi22 port map ( Y=>nx7403, A0=>que_out_25_4_11, A1=>nx10066, B0
      =>que_out_16_4_11, B1=>nx10092);
   ix7406 : aoi22 port map ( Y=>nx7405, A0=>que_out_24_4_11, A1=>nx10040, B0
      =>que_out_22_4_11, B1=>nx10014);
   ix1395 : nand03 port map ( Y=>nx1394, A0=>nx7409, A1=>nx7411, A2=>nx7413
   );
   ix7410 : aoi222 port map ( Y=>nx7409, A0=>que_out_15_4_11, A1=>nx9962, B0
      =>que_out_3_4_11, B1=>nx9988, C0=>que_out_23_4_11, C1=>nx9936);
   ix7412 : aoi22 port map ( Y=>nx7411, A0=>que_out_27_4_11, A1=>nx9910, B0
      =>que_out_4_4_11, B1=>nx9884);
   ix7414 : aoi22 port map ( Y=>nx7413, A0=>que_out_0_4_11, A1=>nx9832, B0=>
      que_out_2_4_11, B1=>nx9858);
   ix1369 : nand03 port map ( Y=>nx1368, A0=>nx7417, A1=>nx7419, A2=>nx7421
   );
   ix7418 : aoi222 port map ( Y=>nx7417, A0=>que_out_26_4_11, A1=>nx9806, B0
      =>que_out_14_4_11, B1=>nx9780, C0=>que_out_11_4_11, C1=>nx9754);
   ix7420 : aoi22 port map ( Y=>nx7419, A0=>que_out_13_4_11, A1=>nx9728, B0
      =>que_out_7_4_11, B1=>nx9702);
   ix7422 : aoi22 port map ( Y=>nx7421, A0=>que_out_12_4_11, A1=>nx9676, B0
      =>que_out_1_4_11, B1=>nx9650);
   ix1563 : or04 port map ( Y=>out_column_4_12, A0=>nx1558, A1=>nx1532, A2=>
      nx1504, A3=>nx1478);
   ix1559 : nand03 port map ( Y=>nx1558, A0=>nx7427, A1=>nx7429, A2=>nx7431
   );
   ix7428 : aoi222 port map ( Y=>nx7427, A0=>que_out_10_4_12, A1=>nx10300, 
      B0=>que_out_6_4_12, B1=>nx10352, C0=>que_out_9_4_12, C1=>nx10326);
   ix7430 : aoi22 port map ( Y=>nx7429, A0=>que_out_5_4_12, A1=>nx10248, B0
      =>que_out_18_4_12, B1=>nx10274);
   ix7432 : aoi22 port map ( Y=>nx7431, A0=>que_out_17_4_12, A1=>nx10222, B0
      =>que_out_20_4_12, B1=>nx10196);
   ix1533 : nand03 port map ( Y=>nx1532, A0=>nx7435, A1=>nx7437, A2=>nx7439
   );
   ix7436 : aoi222 port map ( Y=>nx7435, A0=>que_out_19_4_12, A1=>nx10170, 
      B0=>que_out_21_4_12, B1=>nx10144, C0=>que_out_8_4_12, C1=>nx10118);
   ix7438 : aoi22 port map ( Y=>nx7437, A0=>que_out_25_4_12, A1=>nx10066, B0
      =>que_out_16_4_12, B1=>nx10092);
   ix7440 : aoi22 port map ( Y=>nx7439, A0=>que_out_24_4_12, A1=>nx10040, B0
      =>que_out_22_4_12, B1=>nx10014);
   ix1505 : nand03 port map ( Y=>nx1504, A0=>nx7443, A1=>nx7445, A2=>nx7447
   );
   ix7444 : aoi222 port map ( Y=>nx7443, A0=>que_out_15_4_12, A1=>nx9962, B0
      =>que_out_3_4_12, B1=>nx9988, C0=>que_out_23_4_12, C1=>nx9936);
   ix7446 : aoi22 port map ( Y=>nx7445, A0=>que_out_27_4_12, A1=>nx9910, B0
      =>que_out_4_4_12, B1=>nx9884);
   ix7448 : aoi22 port map ( Y=>nx7447, A0=>que_out_0_4_12, A1=>nx9832, B0=>
      que_out_2_4_12, B1=>nx9858);
   ix1479 : nand03 port map ( Y=>nx1478, A0=>nx7451, A1=>nx7453, A2=>nx7455
   );
   ix7452 : aoi222 port map ( Y=>nx7451, A0=>que_out_26_4_12, A1=>nx9806, B0
      =>que_out_14_4_12, B1=>nx9780, C0=>que_out_11_4_12, C1=>nx9754);
   ix7454 : aoi22 port map ( Y=>nx7453, A0=>que_out_13_4_12, A1=>nx9728, B0
      =>que_out_7_4_12, B1=>nx9702);
   ix7456 : aoi22 port map ( Y=>nx7455, A0=>que_out_12_4_12, A1=>nx9676, B0
      =>que_out_1_4_12, B1=>nx9650);
   ix1673 : or04 port map ( Y=>out_column_4_13, A0=>nx1668, A1=>nx1642, A2=>
      nx1614, A3=>nx1588);
   ix1669 : nand03 port map ( Y=>nx1668, A0=>nx7461, A1=>nx7463, A2=>nx7465
   );
   ix7462 : aoi222 port map ( Y=>nx7461, A0=>que_out_10_4_13, A1=>nx10300, 
      B0=>que_out_6_4_13, B1=>nx10352, C0=>que_out_9_4_13, C1=>nx10326);
   ix7464 : aoi22 port map ( Y=>nx7463, A0=>que_out_5_4_13, A1=>nx10248, B0
      =>que_out_18_4_13, B1=>nx10274);
   ix7466 : aoi22 port map ( Y=>nx7465, A0=>que_out_17_4_13, A1=>nx10222, B0
      =>que_out_20_4_13, B1=>nx10196);
   ix1643 : nand03 port map ( Y=>nx1642, A0=>nx7469, A1=>nx7471, A2=>nx7473
   );
   ix7470 : aoi222 port map ( Y=>nx7469, A0=>que_out_19_4_13, A1=>nx10170, 
      B0=>que_out_21_4_13, B1=>nx10144, C0=>que_out_8_4_13, C1=>nx10118);
   ix7472 : aoi22 port map ( Y=>nx7471, A0=>que_out_25_4_13, A1=>nx10066, B0
      =>que_out_16_4_13, B1=>nx10092);
   ix7474 : aoi22 port map ( Y=>nx7473, A0=>que_out_24_4_13, A1=>nx10040, B0
      =>que_out_22_4_13, B1=>nx10014);
   ix1615 : nand03 port map ( Y=>nx1614, A0=>nx7477, A1=>nx7479, A2=>nx7481
   );
   ix7478 : aoi222 port map ( Y=>nx7477, A0=>que_out_15_4_13, A1=>nx9962, B0
      =>que_out_3_4_13, B1=>nx9988, C0=>que_out_23_4_13, C1=>nx9936);
   ix7480 : aoi22 port map ( Y=>nx7479, A0=>que_out_27_4_13, A1=>nx9910, B0
      =>que_out_4_4_13, B1=>nx9884);
   ix7482 : aoi22 port map ( Y=>nx7481, A0=>que_out_0_4_13, A1=>nx9832, B0=>
      que_out_2_4_13, B1=>nx9858);
   ix1589 : nand03 port map ( Y=>nx1588, A0=>nx7485, A1=>nx7487, A2=>nx7489
   );
   ix7486 : aoi222 port map ( Y=>nx7485, A0=>que_out_26_4_13, A1=>nx9806, B0
      =>que_out_14_4_13, B1=>nx9780, C0=>que_out_11_4_13, C1=>nx9754);
   ix7488 : aoi22 port map ( Y=>nx7487, A0=>que_out_13_4_13, A1=>nx9728, B0
      =>que_out_7_4_13, B1=>nx9702);
   ix7490 : aoi22 port map ( Y=>nx7489, A0=>que_out_12_4_13, A1=>nx9676, B0
      =>que_out_1_4_13, B1=>nx9650);
   ix1783 : or04 port map ( Y=>out_column_4_14, A0=>nx1778, A1=>nx1752, A2=>
      nx1724, A3=>nx1698);
   ix1779 : nand03 port map ( Y=>nx1778, A0=>nx7495, A1=>nx7497, A2=>nx7499
   );
   ix7496 : aoi222 port map ( Y=>nx7495, A0=>que_out_10_4_14, A1=>nx10302, 
      B0=>que_out_6_4_14, B1=>nx10354, C0=>que_out_9_4_14, C1=>nx10328);
   ix7498 : aoi22 port map ( Y=>nx7497, A0=>que_out_5_4_14, A1=>nx10250, B0
      =>que_out_18_4_14, B1=>nx10276);
   ix7500 : aoi22 port map ( Y=>nx7499, A0=>que_out_17_4_14, A1=>nx10224, B0
      =>que_out_20_4_14, B1=>nx10198);
   ix1753 : nand03 port map ( Y=>nx1752, A0=>nx7503, A1=>nx7505, A2=>nx7507
   );
   ix7504 : aoi222 port map ( Y=>nx7503, A0=>que_out_19_4_14, A1=>nx10172, 
      B0=>que_out_21_4_14, B1=>nx10146, C0=>que_out_8_4_14, C1=>nx10120);
   ix7506 : aoi22 port map ( Y=>nx7505, A0=>que_out_25_4_14, A1=>nx10068, B0
      =>que_out_16_4_14, B1=>nx10094);
   ix7508 : aoi22 port map ( Y=>nx7507, A0=>que_out_24_4_14, A1=>nx10042, B0
      =>que_out_22_4_14, B1=>nx10016);
   ix1725 : nand03 port map ( Y=>nx1724, A0=>nx7511, A1=>nx7513, A2=>nx7515
   );
   ix7512 : aoi222 port map ( Y=>nx7511, A0=>que_out_15_4_14, A1=>nx9964, B0
      =>que_out_3_4_14, B1=>nx9990, C0=>que_out_23_4_14, C1=>nx9938);
   ix7514 : aoi22 port map ( Y=>nx7513, A0=>que_out_27_4_14, A1=>nx9912, B0
      =>que_out_4_4_14, B1=>nx9886);
   ix7516 : aoi22 port map ( Y=>nx7515, A0=>que_out_0_4_14, A1=>nx9834, B0=>
      que_out_2_4_14, B1=>nx9860);
   ix1699 : nand03 port map ( Y=>nx1698, A0=>nx7519, A1=>nx7521, A2=>nx7523
   );
   ix7520 : aoi222 port map ( Y=>nx7519, A0=>que_out_26_4_14, A1=>nx9808, B0
      =>que_out_14_4_14, B1=>nx9782, C0=>que_out_11_4_14, C1=>nx9756);
   ix7522 : aoi22 port map ( Y=>nx7521, A0=>que_out_13_4_14, A1=>nx9730, B0
      =>que_out_7_4_14, B1=>nx9704);
   ix7524 : aoi22 port map ( Y=>nx7523, A0=>que_out_12_4_14, A1=>nx9678, B0
      =>que_out_1_4_14, B1=>nx9652);
   ix1893 : or04 port map ( Y=>out_column_4_15, A0=>nx1888, A1=>nx1862, A2=>
      nx1834, A3=>nx1808);
   ix1889 : nand03 port map ( Y=>nx1888, A0=>nx7529, A1=>nx7531, A2=>nx7533
   );
   ix7530 : aoi222 port map ( Y=>nx7529, A0=>que_out_10_4_15, A1=>nx10302, 
      B0=>que_out_6_4_15, B1=>nx10354, C0=>que_out_9_4_15, C1=>nx10328);
   ix7532 : aoi22 port map ( Y=>nx7531, A0=>que_out_5_4_15, A1=>nx10250, B0
      =>que_out_18_4_15, B1=>nx10276);
   ix7534 : aoi22 port map ( Y=>nx7533, A0=>que_out_17_4_15, A1=>nx10224, B0
      =>que_out_20_4_15, B1=>nx10198);
   ix1863 : nand03 port map ( Y=>nx1862, A0=>nx7537, A1=>nx7539, A2=>nx7541
   );
   ix7538 : aoi222 port map ( Y=>nx7537, A0=>que_out_19_4_15, A1=>nx10172, 
      B0=>que_out_21_4_15, B1=>nx10146, C0=>que_out_8_4_15, C1=>nx10120);
   ix7540 : aoi22 port map ( Y=>nx7539, A0=>que_out_25_4_15, A1=>nx10068, B0
      =>que_out_16_4_15, B1=>nx10094);
   ix7542 : aoi22 port map ( Y=>nx7541, A0=>que_out_24_4_15, A1=>nx10042, B0
      =>que_out_22_4_15, B1=>nx10016);
   ix1835 : nand03 port map ( Y=>nx1834, A0=>nx7545, A1=>nx7547, A2=>nx7549
   );
   ix7546 : aoi222 port map ( Y=>nx7545, A0=>que_out_15_4_15, A1=>nx9964, B0
      =>que_out_3_4_15, B1=>nx9990, C0=>que_out_23_4_15, C1=>nx9938);
   ix7548 : aoi22 port map ( Y=>nx7547, A0=>que_out_27_4_15, A1=>nx9912, B0
      =>que_out_4_4_15, B1=>nx9886);
   ix7550 : aoi22 port map ( Y=>nx7549, A0=>que_out_0_4_15, A1=>nx9834, B0=>
      que_out_2_4_15, B1=>nx9860);
   ix1809 : nand03 port map ( Y=>nx1808, A0=>nx7553, A1=>nx7555, A2=>nx7557
   );
   ix7554 : aoi222 port map ( Y=>nx7553, A0=>que_out_26_4_15, A1=>nx9808, B0
      =>que_out_14_4_15, B1=>nx9782, C0=>que_out_11_4_15, C1=>nx9756);
   ix7556 : aoi22 port map ( Y=>nx7555, A0=>que_out_13_4_15, A1=>nx9730, B0
      =>que_out_7_4_15, B1=>nx9704);
   ix7558 : aoi22 port map ( Y=>nx7557, A0=>que_out_12_4_15, A1=>nx9678, B0
      =>que_out_1_4_15, B1=>nx9652);
   ix2003 : or04 port map ( Y=>out_column_3_0, A0=>nx1998, A1=>nx1972, A2=>
      nx1944, A3=>nx1918);
   ix1999 : nand03 port map ( Y=>nx1998, A0=>nx7563, A1=>nx7565, A2=>nx7567
   );
   ix7564 : aoi222 port map ( Y=>nx7563, A0=>que_out_10_3_0, A1=>nx10302, B0
      =>que_out_6_3_0, B1=>nx10354, C0=>que_out_9_3_0, C1=>nx10328);
   ix7566 : aoi22 port map ( Y=>nx7565, A0=>que_out_5_3_0, A1=>nx10250, B0=>
      que_out_18_3_0, B1=>nx10276);
   ix7568 : aoi22 port map ( Y=>nx7567, A0=>que_out_17_3_0, A1=>nx10224, B0
      =>que_out_20_3_0, B1=>nx10198);
   ix1973 : nand03 port map ( Y=>nx1972, A0=>nx7571, A1=>nx7573, A2=>nx7575
   );
   ix7572 : aoi222 port map ( Y=>nx7571, A0=>que_out_19_3_0, A1=>nx10172, B0
      =>que_out_21_3_0, B1=>nx10146, C0=>que_out_8_3_0, C1=>nx10120);
   ix7574 : aoi22 port map ( Y=>nx7573, A0=>que_out_25_3_0, A1=>nx10068, B0
      =>que_out_16_3_0, B1=>nx10094);
   ix7576 : aoi22 port map ( Y=>nx7575, A0=>que_out_24_3_0, A1=>nx10042, B0
      =>que_out_22_3_0, B1=>nx10016);
   ix1945 : nand03 port map ( Y=>nx1944, A0=>nx7579, A1=>nx7581, A2=>nx7583
   );
   ix7580 : aoi222 port map ( Y=>nx7579, A0=>que_out_15_3_0, A1=>nx9964, B0
      =>que_out_3_3_0, B1=>nx9990, C0=>que_out_23_3_0, C1=>nx9938);
   ix7582 : aoi22 port map ( Y=>nx7581, A0=>que_out_27_3_0, A1=>nx9912, B0=>
      que_out_4_3_0, B1=>nx9886);
   ix7584 : aoi22 port map ( Y=>nx7583, A0=>que_out_0_3_0, A1=>nx9834, B0=>
      que_out_2_3_0, B1=>nx9860);
   ix1919 : nand03 port map ( Y=>nx1918, A0=>nx7587, A1=>nx7589, A2=>nx7591
   );
   ix7588 : aoi222 port map ( Y=>nx7587, A0=>que_out_26_3_0, A1=>nx9808, B0
      =>que_out_14_3_0, B1=>nx9782, C0=>que_out_11_3_0, C1=>nx9756);
   ix7590 : aoi22 port map ( Y=>nx7589, A0=>que_out_13_3_0, A1=>nx9730, B0=>
      que_out_7_3_0, B1=>nx9704);
   ix7592 : aoi22 port map ( Y=>nx7591, A0=>que_out_12_3_0, A1=>nx9678, B0=>
      que_out_1_3_0, B1=>nx9652);
   ix2113 : or04 port map ( Y=>out_column_3_1, A0=>nx2108, A1=>nx2082, A2=>
      nx2054, A3=>nx2028);
   ix2109 : nand03 port map ( Y=>nx2108, A0=>nx7597, A1=>nx7599, A2=>nx7601
   );
   ix7598 : aoi222 port map ( Y=>nx7597, A0=>que_out_10_3_1, A1=>nx10302, B0
      =>que_out_6_3_1, B1=>nx10354, C0=>que_out_9_3_1, C1=>nx10328);
   ix7600 : aoi22 port map ( Y=>nx7599, A0=>que_out_5_3_1, A1=>nx10250, B0=>
      que_out_18_3_1, B1=>nx10276);
   ix7602 : aoi22 port map ( Y=>nx7601, A0=>que_out_17_3_1, A1=>nx10224, B0
      =>que_out_20_3_1, B1=>nx10198);
   ix2083 : nand03 port map ( Y=>nx2082, A0=>nx7605, A1=>nx7607, A2=>nx7609
   );
   ix7606 : aoi222 port map ( Y=>nx7605, A0=>que_out_19_3_1, A1=>nx10172, B0
      =>que_out_21_3_1, B1=>nx10146, C0=>que_out_8_3_1, C1=>nx10120);
   ix7608 : aoi22 port map ( Y=>nx7607, A0=>que_out_25_3_1, A1=>nx10068, B0
      =>que_out_16_3_1, B1=>nx10094);
   ix7610 : aoi22 port map ( Y=>nx7609, A0=>que_out_24_3_1, A1=>nx10042, B0
      =>que_out_22_3_1, B1=>nx10016);
   ix2055 : nand03 port map ( Y=>nx2054, A0=>nx7613, A1=>nx7615, A2=>nx7617
   );
   ix7614 : aoi222 port map ( Y=>nx7613, A0=>que_out_15_3_1, A1=>nx9964, B0
      =>que_out_3_3_1, B1=>nx9990, C0=>que_out_23_3_1, C1=>nx9938);
   ix7616 : aoi22 port map ( Y=>nx7615, A0=>que_out_27_3_1, A1=>nx9912, B0=>
      que_out_4_3_1, B1=>nx9886);
   ix7618 : aoi22 port map ( Y=>nx7617, A0=>que_out_0_3_1, A1=>nx9834, B0=>
      que_out_2_3_1, B1=>nx9860);
   ix2029 : nand03 port map ( Y=>nx2028, A0=>nx7621, A1=>nx7623, A2=>nx7625
   );
   ix7622 : aoi222 port map ( Y=>nx7621, A0=>que_out_26_3_1, A1=>nx9808, B0
      =>que_out_14_3_1, B1=>nx9782, C0=>que_out_11_3_1, C1=>nx9756);
   ix7624 : aoi22 port map ( Y=>nx7623, A0=>que_out_13_3_1, A1=>nx9730, B0=>
      que_out_7_3_1, B1=>nx9704);
   ix7626 : aoi22 port map ( Y=>nx7625, A0=>que_out_12_3_1, A1=>nx9678, B0=>
      que_out_1_3_1, B1=>nx9652);
   ix2223 : or04 port map ( Y=>out_column_3_2, A0=>nx2218, A1=>nx2192, A2=>
      nx2164, A3=>nx2138);
   ix2219 : nand03 port map ( Y=>nx2218, A0=>nx7631, A1=>nx7633, A2=>nx7635
   );
   ix7632 : aoi222 port map ( Y=>nx7631, A0=>que_out_10_3_2, A1=>nx10302, B0
      =>que_out_6_3_2, B1=>nx10354, C0=>que_out_9_3_2, C1=>nx10328);
   ix7634 : aoi22 port map ( Y=>nx7633, A0=>que_out_5_3_2, A1=>nx10250, B0=>
      que_out_18_3_2, B1=>nx10276);
   ix7636 : aoi22 port map ( Y=>nx7635, A0=>que_out_17_3_2, A1=>nx10224, B0
      =>que_out_20_3_2, B1=>nx10198);
   ix2193 : nand03 port map ( Y=>nx2192, A0=>nx7639, A1=>nx7641, A2=>nx7643
   );
   ix7640 : aoi222 port map ( Y=>nx7639, A0=>que_out_19_3_2, A1=>nx10172, B0
      =>que_out_21_3_2, B1=>nx10146, C0=>que_out_8_3_2, C1=>nx10120);
   ix7642 : aoi22 port map ( Y=>nx7641, A0=>que_out_25_3_2, A1=>nx10068, B0
      =>que_out_16_3_2, B1=>nx10094);
   ix7644 : aoi22 port map ( Y=>nx7643, A0=>que_out_24_3_2, A1=>nx10042, B0
      =>que_out_22_3_2, B1=>nx10016);
   ix2165 : nand03 port map ( Y=>nx2164, A0=>nx7647, A1=>nx7649, A2=>nx7651
   );
   ix7648 : aoi222 port map ( Y=>nx7647, A0=>que_out_15_3_2, A1=>nx9964, B0
      =>que_out_3_3_2, B1=>nx9990, C0=>que_out_23_3_2, C1=>nx9938);
   ix7650 : aoi22 port map ( Y=>nx7649, A0=>que_out_27_3_2, A1=>nx9912, B0=>
      que_out_4_3_2, B1=>nx9886);
   ix7652 : aoi22 port map ( Y=>nx7651, A0=>que_out_0_3_2, A1=>nx9834, B0=>
      que_out_2_3_2, B1=>nx9860);
   ix2139 : nand03 port map ( Y=>nx2138, A0=>nx7655, A1=>nx7657, A2=>nx7659
   );
   ix7656 : aoi222 port map ( Y=>nx7655, A0=>que_out_26_3_2, A1=>nx9808, B0
      =>que_out_14_3_2, B1=>nx9782, C0=>que_out_11_3_2, C1=>nx9756);
   ix7658 : aoi22 port map ( Y=>nx7657, A0=>que_out_13_3_2, A1=>nx9730, B0=>
      que_out_7_3_2, B1=>nx9704);
   ix7660 : aoi22 port map ( Y=>nx7659, A0=>que_out_12_3_2, A1=>nx9678, B0=>
      que_out_1_3_2, B1=>nx9652);
   ix2333 : or04 port map ( Y=>out_column_3_3, A0=>nx2328, A1=>nx2302, A2=>
      nx2274, A3=>nx2248);
   ix2329 : nand03 port map ( Y=>nx2328, A0=>nx7665, A1=>nx7667, A2=>nx7669
   );
   ix7666 : aoi222 port map ( Y=>nx7665, A0=>que_out_10_3_3, A1=>nx10302, B0
      =>que_out_6_3_3, B1=>nx10354, C0=>que_out_9_3_3, C1=>nx10328);
   ix7668 : aoi22 port map ( Y=>nx7667, A0=>que_out_5_3_3, A1=>nx10250, B0=>
      que_out_18_3_3, B1=>nx10276);
   ix7670 : aoi22 port map ( Y=>nx7669, A0=>que_out_17_3_3, A1=>nx10224, B0
      =>que_out_20_3_3, B1=>nx10198);
   ix2303 : nand03 port map ( Y=>nx2302, A0=>nx7673, A1=>nx7675, A2=>nx7677
   );
   ix7674 : aoi222 port map ( Y=>nx7673, A0=>que_out_19_3_3, A1=>nx10172, B0
      =>que_out_21_3_3, B1=>nx10146, C0=>que_out_8_3_3, C1=>nx10120);
   ix7676 : aoi22 port map ( Y=>nx7675, A0=>que_out_25_3_3, A1=>nx10068, B0
      =>que_out_16_3_3, B1=>nx10094);
   ix7678 : aoi22 port map ( Y=>nx7677, A0=>que_out_24_3_3, A1=>nx10042, B0
      =>que_out_22_3_3, B1=>nx10016);
   ix2275 : nand03 port map ( Y=>nx2274, A0=>nx7681, A1=>nx7683, A2=>nx7685
   );
   ix7682 : aoi222 port map ( Y=>nx7681, A0=>que_out_15_3_3, A1=>nx9964, B0
      =>que_out_3_3_3, B1=>nx9990, C0=>que_out_23_3_3, C1=>nx9938);
   ix7684 : aoi22 port map ( Y=>nx7683, A0=>que_out_27_3_3, A1=>nx9912, B0=>
      que_out_4_3_3, B1=>nx9886);
   ix7686 : aoi22 port map ( Y=>nx7685, A0=>que_out_0_3_3, A1=>nx9834, B0=>
      que_out_2_3_3, B1=>nx9860);
   ix2249 : nand03 port map ( Y=>nx2248, A0=>nx7689, A1=>nx7691, A2=>nx7693
   );
   ix7690 : aoi222 port map ( Y=>nx7689, A0=>que_out_26_3_3, A1=>nx9808, B0
      =>que_out_14_3_3, B1=>nx9782, C0=>que_out_11_3_3, C1=>nx9756);
   ix7692 : aoi22 port map ( Y=>nx7691, A0=>que_out_13_3_3, A1=>nx9730, B0=>
      que_out_7_3_3, B1=>nx9704);
   ix7694 : aoi22 port map ( Y=>nx7693, A0=>que_out_12_3_3, A1=>nx9678, B0=>
      que_out_1_3_3, B1=>nx9652);
   ix2443 : or04 port map ( Y=>out_column_3_4, A0=>nx2438, A1=>nx2412, A2=>
      nx2384, A3=>nx2358);
   ix2439 : nand03 port map ( Y=>nx2438, A0=>nx7699, A1=>nx7701, A2=>nx7703
   );
   ix7700 : aoi222 port map ( Y=>nx7699, A0=>que_out_10_3_4, A1=>nx10302, B0
      =>que_out_6_3_4, B1=>nx10354, C0=>que_out_9_3_4, C1=>nx10328);
   ix7702 : aoi22 port map ( Y=>nx7701, A0=>que_out_5_3_4, A1=>nx10250, B0=>
      que_out_18_3_4, B1=>nx10276);
   ix7704 : aoi22 port map ( Y=>nx7703, A0=>que_out_17_3_4, A1=>nx10224, B0
      =>que_out_20_3_4, B1=>nx10198);
   ix2413 : nand03 port map ( Y=>nx2412, A0=>nx7707, A1=>nx7709, A2=>nx7711
   );
   ix7708 : aoi222 port map ( Y=>nx7707, A0=>que_out_19_3_4, A1=>nx10172, B0
      =>que_out_21_3_4, B1=>nx10146, C0=>que_out_8_3_4, C1=>nx10120);
   ix7710 : aoi22 port map ( Y=>nx7709, A0=>que_out_25_3_4, A1=>nx10068, B0
      =>que_out_16_3_4, B1=>nx10094);
   ix7712 : aoi22 port map ( Y=>nx7711, A0=>que_out_24_3_4, A1=>nx10042, B0
      =>que_out_22_3_4, B1=>nx10016);
   ix2385 : nand03 port map ( Y=>nx2384, A0=>nx7715, A1=>nx7717, A2=>nx7719
   );
   ix7716 : aoi222 port map ( Y=>nx7715, A0=>que_out_15_3_4, A1=>nx9964, B0
      =>que_out_3_3_4, B1=>nx9990, C0=>que_out_23_3_4, C1=>nx9938);
   ix7718 : aoi22 port map ( Y=>nx7717, A0=>que_out_27_3_4, A1=>nx9912, B0=>
      que_out_4_3_4, B1=>nx9886);
   ix7720 : aoi22 port map ( Y=>nx7719, A0=>que_out_0_3_4, A1=>nx9834, B0=>
      que_out_2_3_4, B1=>nx9860);
   ix2359 : nand03 port map ( Y=>nx2358, A0=>nx7723, A1=>nx7725, A2=>nx7727
   );
   ix7724 : aoi222 port map ( Y=>nx7723, A0=>que_out_26_3_4, A1=>nx9808, B0
      =>que_out_14_3_4, B1=>nx9782, C0=>que_out_11_3_4, C1=>nx9756);
   ix7726 : aoi22 port map ( Y=>nx7725, A0=>que_out_13_3_4, A1=>nx9730, B0=>
      que_out_7_3_4, B1=>nx9704);
   ix7728 : aoi22 port map ( Y=>nx7727, A0=>que_out_12_3_4, A1=>nx9678, B0=>
      que_out_1_3_4, B1=>nx9652);
   ix2553 : or04 port map ( Y=>out_column_3_5, A0=>nx2548, A1=>nx2522, A2=>
      nx2494, A3=>nx2468);
   ix2549 : nand03 port map ( Y=>nx2548, A0=>nx7733, A1=>nx7735, A2=>nx7737
   );
   ix7734 : aoi222 port map ( Y=>nx7733, A0=>que_out_10_3_5, A1=>nx10304, B0
      =>que_out_6_3_5, B1=>nx10356, C0=>que_out_9_3_5, C1=>nx10330);
   ix7736 : aoi22 port map ( Y=>nx7735, A0=>que_out_5_3_5, A1=>nx10252, B0=>
      que_out_18_3_5, B1=>nx10278);
   ix7738 : aoi22 port map ( Y=>nx7737, A0=>que_out_17_3_5, A1=>nx10226, B0
      =>que_out_20_3_5, B1=>nx10200);
   ix2523 : nand03 port map ( Y=>nx2522, A0=>nx7741, A1=>nx7743, A2=>nx7745
   );
   ix7742 : aoi222 port map ( Y=>nx7741, A0=>que_out_19_3_5, A1=>nx10174, B0
      =>que_out_21_3_5, B1=>nx10148, C0=>que_out_8_3_5, C1=>nx10122);
   ix7744 : aoi22 port map ( Y=>nx7743, A0=>que_out_25_3_5, A1=>nx10070, B0
      =>que_out_16_3_5, B1=>nx10096);
   ix7746 : aoi22 port map ( Y=>nx7745, A0=>que_out_24_3_5, A1=>nx10044, B0
      =>que_out_22_3_5, B1=>nx10018);
   ix2495 : nand03 port map ( Y=>nx2494, A0=>nx7749, A1=>nx7751, A2=>nx7753
   );
   ix7750 : aoi222 port map ( Y=>nx7749, A0=>que_out_15_3_5, A1=>nx9966, B0
      =>que_out_3_3_5, B1=>nx9992, C0=>que_out_23_3_5, C1=>nx9940);
   ix7752 : aoi22 port map ( Y=>nx7751, A0=>que_out_27_3_5, A1=>nx9914, B0=>
      que_out_4_3_5, B1=>nx9888);
   ix7754 : aoi22 port map ( Y=>nx7753, A0=>que_out_0_3_5, A1=>nx9836, B0=>
      que_out_2_3_5, B1=>nx9862);
   ix2469 : nand03 port map ( Y=>nx2468, A0=>nx7757, A1=>nx7759, A2=>nx7761
   );
   ix7758 : aoi222 port map ( Y=>nx7757, A0=>que_out_26_3_5, A1=>nx9810, B0
      =>que_out_14_3_5, B1=>nx9784, C0=>que_out_11_3_5, C1=>nx9758);
   ix7760 : aoi22 port map ( Y=>nx7759, A0=>que_out_13_3_5, A1=>nx9732, B0=>
      que_out_7_3_5, B1=>nx9706);
   ix7762 : aoi22 port map ( Y=>nx7761, A0=>que_out_12_3_5, A1=>nx9680, B0=>
      que_out_1_3_5, B1=>nx9654);
   ix2663 : or04 port map ( Y=>out_column_3_6, A0=>nx2658, A1=>nx2632, A2=>
      nx2604, A3=>nx2578);
   ix2659 : nand03 port map ( Y=>nx2658, A0=>nx7767, A1=>nx7769, A2=>nx7771
   );
   ix7768 : aoi222 port map ( Y=>nx7767, A0=>que_out_10_3_6, A1=>nx10304, B0
      =>que_out_6_3_6, B1=>nx10356, C0=>que_out_9_3_6, C1=>nx10330);
   ix7770 : aoi22 port map ( Y=>nx7769, A0=>que_out_5_3_6, A1=>nx10252, B0=>
      que_out_18_3_6, B1=>nx10278);
   ix7772 : aoi22 port map ( Y=>nx7771, A0=>que_out_17_3_6, A1=>nx10226, B0
      =>que_out_20_3_6, B1=>nx10200);
   ix2633 : nand03 port map ( Y=>nx2632, A0=>nx7775, A1=>nx7777, A2=>nx7779
   );
   ix7776 : aoi222 port map ( Y=>nx7775, A0=>que_out_19_3_6, A1=>nx10174, B0
      =>que_out_21_3_6, B1=>nx10148, C0=>que_out_8_3_6, C1=>nx10122);
   ix7778 : aoi22 port map ( Y=>nx7777, A0=>que_out_25_3_6, A1=>nx10070, B0
      =>que_out_16_3_6, B1=>nx10096);
   ix7780 : aoi22 port map ( Y=>nx7779, A0=>que_out_24_3_6, A1=>nx10044, B0
      =>que_out_22_3_6, B1=>nx10018);
   ix2605 : nand03 port map ( Y=>nx2604, A0=>nx7783, A1=>nx7785, A2=>nx7787
   );
   ix7784 : aoi222 port map ( Y=>nx7783, A0=>que_out_15_3_6, A1=>nx9966, B0
      =>que_out_3_3_6, B1=>nx9992, C0=>que_out_23_3_6, C1=>nx9940);
   ix7786 : aoi22 port map ( Y=>nx7785, A0=>que_out_27_3_6, A1=>nx9914, B0=>
      que_out_4_3_6, B1=>nx9888);
   ix7788 : aoi22 port map ( Y=>nx7787, A0=>que_out_0_3_6, A1=>nx9836, B0=>
      que_out_2_3_6, B1=>nx9862);
   ix2579 : nand03 port map ( Y=>nx2578, A0=>nx7791, A1=>nx7793, A2=>nx7795
   );
   ix7792 : aoi222 port map ( Y=>nx7791, A0=>que_out_26_3_6, A1=>nx9810, B0
      =>que_out_14_3_6, B1=>nx9784, C0=>que_out_11_3_6, C1=>nx9758);
   ix7794 : aoi22 port map ( Y=>nx7793, A0=>que_out_13_3_6, A1=>nx9732, B0=>
      que_out_7_3_6, B1=>nx9706);
   ix7796 : aoi22 port map ( Y=>nx7795, A0=>que_out_12_3_6, A1=>nx9680, B0=>
      que_out_1_3_6, B1=>nx9654);
   ix2773 : or04 port map ( Y=>out_column_3_7, A0=>nx2768, A1=>nx2742, A2=>
      nx2714, A3=>nx2688);
   ix2769 : nand03 port map ( Y=>nx2768, A0=>nx7801, A1=>nx7803, A2=>nx7805
   );
   ix7802 : aoi222 port map ( Y=>nx7801, A0=>que_out_10_3_7, A1=>nx10304, B0
      =>que_out_6_3_7, B1=>nx10356, C0=>que_out_9_3_7, C1=>nx10330);
   ix7804 : aoi22 port map ( Y=>nx7803, A0=>que_out_5_3_7, A1=>nx10252, B0=>
      que_out_18_3_7, B1=>nx10278);
   ix7806 : aoi22 port map ( Y=>nx7805, A0=>que_out_17_3_7, A1=>nx10226, B0
      =>que_out_20_3_7, B1=>nx10200);
   ix2743 : nand03 port map ( Y=>nx2742, A0=>nx7809, A1=>nx7811, A2=>nx7813
   );
   ix7810 : aoi222 port map ( Y=>nx7809, A0=>que_out_19_3_7, A1=>nx10174, B0
      =>que_out_21_3_7, B1=>nx10148, C0=>que_out_8_3_7, C1=>nx10122);
   ix7812 : aoi22 port map ( Y=>nx7811, A0=>que_out_25_3_7, A1=>nx10070, B0
      =>que_out_16_3_7, B1=>nx10096);
   ix7814 : aoi22 port map ( Y=>nx7813, A0=>que_out_24_3_7, A1=>nx10044, B0
      =>que_out_22_3_7, B1=>nx10018);
   ix2715 : nand03 port map ( Y=>nx2714, A0=>nx7817, A1=>nx7819, A2=>nx7821
   );
   ix7818 : aoi222 port map ( Y=>nx7817, A0=>que_out_15_3_7, A1=>nx9966, B0
      =>que_out_3_3_7, B1=>nx9992, C0=>que_out_23_3_7, C1=>nx9940);
   ix7820 : aoi22 port map ( Y=>nx7819, A0=>que_out_27_3_7, A1=>nx9914, B0=>
      que_out_4_3_7, B1=>nx9888);
   ix7822 : aoi22 port map ( Y=>nx7821, A0=>que_out_0_3_7, A1=>nx9836, B0=>
      que_out_2_3_7, B1=>nx9862);
   ix2689 : nand03 port map ( Y=>nx2688, A0=>nx7825, A1=>nx7827, A2=>nx7829
   );
   ix7826 : aoi222 port map ( Y=>nx7825, A0=>que_out_26_3_7, A1=>nx9810, B0
      =>que_out_14_3_7, B1=>nx9784, C0=>que_out_11_3_7, C1=>nx9758);
   ix7828 : aoi22 port map ( Y=>nx7827, A0=>que_out_13_3_7, A1=>nx9732, B0=>
      que_out_7_3_7, B1=>nx9706);
   ix7830 : aoi22 port map ( Y=>nx7829, A0=>que_out_12_3_7, A1=>nx9680, B0=>
      que_out_1_3_7, B1=>nx9654);
   ix2883 : or04 port map ( Y=>out_column_3_8, A0=>nx2878, A1=>nx2852, A2=>
      nx2824, A3=>nx2798);
   ix2879 : nand03 port map ( Y=>nx2878, A0=>nx7835, A1=>nx7837, A2=>nx7839
   );
   ix7836 : aoi222 port map ( Y=>nx7835, A0=>que_out_10_3_8, A1=>nx10304, B0
      =>que_out_6_3_8, B1=>nx10356, C0=>que_out_9_3_8, C1=>nx10330);
   ix7838 : aoi22 port map ( Y=>nx7837, A0=>que_out_5_3_8, A1=>nx10252, B0=>
      que_out_18_3_8, B1=>nx10278);
   ix7840 : aoi22 port map ( Y=>nx7839, A0=>que_out_17_3_8, A1=>nx10226, B0
      =>que_out_20_3_8, B1=>nx10200);
   ix2853 : nand03 port map ( Y=>nx2852, A0=>nx7843, A1=>nx7845, A2=>nx7847
   );
   ix7844 : aoi222 port map ( Y=>nx7843, A0=>que_out_19_3_8, A1=>nx10174, B0
      =>que_out_21_3_8, B1=>nx10148, C0=>que_out_8_3_8, C1=>nx10122);
   ix7846 : aoi22 port map ( Y=>nx7845, A0=>que_out_25_3_8, A1=>nx10070, B0
      =>que_out_16_3_8, B1=>nx10096);
   ix7848 : aoi22 port map ( Y=>nx7847, A0=>que_out_24_3_8, A1=>nx10044, B0
      =>que_out_22_3_8, B1=>nx10018);
   ix2825 : nand03 port map ( Y=>nx2824, A0=>nx7851, A1=>nx7853, A2=>nx7855
   );
   ix7852 : aoi222 port map ( Y=>nx7851, A0=>que_out_15_3_8, A1=>nx9966, B0
      =>que_out_3_3_8, B1=>nx9992, C0=>que_out_23_3_8, C1=>nx9940);
   ix7854 : aoi22 port map ( Y=>nx7853, A0=>que_out_27_3_8, A1=>nx9914, B0=>
      que_out_4_3_8, B1=>nx9888);
   ix7856 : aoi22 port map ( Y=>nx7855, A0=>que_out_0_3_8, A1=>nx9836, B0=>
      que_out_2_3_8, B1=>nx9862);
   ix2799 : nand03 port map ( Y=>nx2798, A0=>nx7859, A1=>nx7861, A2=>nx7863
   );
   ix7860 : aoi222 port map ( Y=>nx7859, A0=>que_out_26_3_8, A1=>nx9810, B0
      =>que_out_14_3_8, B1=>nx9784, C0=>que_out_11_3_8, C1=>nx9758);
   ix7862 : aoi22 port map ( Y=>nx7861, A0=>que_out_13_3_8, A1=>nx9732, B0=>
      que_out_7_3_8, B1=>nx9706);
   ix7864 : aoi22 port map ( Y=>nx7863, A0=>que_out_12_3_8, A1=>nx9680, B0=>
      que_out_1_3_8, B1=>nx9654);
   ix2993 : or04 port map ( Y=>out_column_3_9, A0=>nx2988, A1=>nx2962, A2=>
      nx2934, A3=>nx2908);
   ix2989 : nand03 port map ( Y=>nx2988, A0=>nx7869, A1=>nx7871, A2=>nx7873
   );
   ix7870 : aoi222 port map ( Y=>nx7869, A0=>que_out_10_3_9, A1=>nx10304, B0
      =>que_out_6_3_9, B1=>nx10356, C0=>que_out_9_3_9, C1=>nx10330);
   ix7872 : aoi22 port map ( Y=>nx7871, A0=>que_out_5_3_9, A1=>nx10252, B0=>
      que_out_18_3_9, B1=>nx10278);
   ix7874 : aoi22 port map ( Y=>nx7873, A0=>que_out_17_3_9, A1=>nx10226, B0
      =>que_out_20_3_9, B1=>nx10200);
   ix2963 : nand03 port map ( Y=>nx2962, A0=>nx7877, A1=>nx7879, A2=>nx7881
   );
   ix7878 : aoi222 port map ( Y=>nx7877, A0=>que_out_19_3_9, A1=>nx10174, B0
      =>que_out_21_3_9, B1=>nx10148, C0=>que_out_8_3_9, C1=>nx10122);
   ix7880 : aoi22 port map ( Y=>nx7879, A0=>que_out_25_3_9, A1=>nx10070, B0
      =>que_out_16_3_9, B1=>nx10096);
   ix7882 : aoi22 port map ( Y=>nx7881, A0=>que_out_24_3_9, A1=>nx10044, B0
      =>que_out_22_3_9, B1=>nx10018);
   ix2935 : nand03 port map ( Y=>nx2934, A0=>nx7885, A1=>nx7887, A2=>nx7889
   );
   ix7886 : aoi222 port map ( Y=>nx7885, A0=>que_out_15_3_9, A1=>nx9966, B0
      =>que_out_3_3_9, B1=>nx9992, C0=>que_out_23_3_9, C1=>nx9940);
   ix7888 : aoi22 port map ( Y=>nx7887, A0=>que_out_27_3_9, A1=>nx9914, B0=>
      que_out_4_3_9, B1=>nx9888);
   ix7890 : aoi22 port map ( Y=>nx7889, A0=>que_out_0_3_9, A1=>nx9836, B0=>
      que_out_2_3_9, B1=>nx9862);
   ix2909 : nand03 port map ( Y=>nx2908, A0=>nx7893, A1=>nx7895, A2=>nx7897
   );
   ix7894 : aoi222 port map ( Y=>nx7893, A0=>que_out_26_3_9, A1=>nx9810, B0
      =>que_out_14_3_9, B1=>nx9784, C0=>que_out_11_3_9, C1=>nx9758);
   ix7896 : aoi22 port map ( Y=>nx7895, A0=>que_out_13_3_9, A1=>nx9732, B0=>
      que_out_7_3_9, B1=>nx9706);
   ix7898 : aoi22 port map ( Y=>nx7897, A0=>que_out_12_3_9, A1=>nx9680, B0=>
      que_out_1_3_9, B1=>nx9654);
   ix3103 : or04 port map ( Y=>out_column_3_10, A0=>nx3098, A1=>nx3072, A2=>
      nx3044, A3=>nx3018);
   ix3099 : nand03 port map ( Y=>nx3098, A0=>nx7903, A1=>nx7905, A2=>nx7907
   );
   ix7904 : aoi222 port map ( Y=>nx7903, A0=>que_out_10_3_10, A1=>nx10304, 
      B0=>que_out_6_3_10, B1=>nx10356, C0=>que_out_9_3_10, C1=>nx10330);
   ix7906 : aoi22 port map ( Y=>nx7905, A0=>que_out_5_3_10, A1=>nx10252, B0
      =>que_out_18_3_10, B1=>nx10278);
   ix7908 : aoi22 port map ( Y=>nx7907, A0=>que_out_17_3_10, A1=>nx10226, B0
      =>que_out_20_3_10, B1=>nx10200);
   ix3073 : nand03 port map ( Y=>nx3072, A0=>nx7911, A1=>nx7913, A2=>nx7915
   );
   ix7912 : aoi222 port map ( Y=>nx7911, A0=>que_out_19_3_10, A1=>nx10174, 
      B0=>que_out_21_3_10, B1=>nx10148, C0=>que_out_8_3_10, C1=>nx10122);
   ix7914 : aoi22 port map ( Y=>nx7913, A0=>que_out_25_3_10, A1=>nx10070, B0
      =>que_out_16_3_10, B1=>nx10096);
   ix7916 : aoi22 port map ( Y=>nx7915, A0=>que_out_24_3_10, A1=>nx10044, B0
      =>que_out_22_3_10, B1=>nx10018);
   ix3045 : nand03 port map ( Y=>nx3044, A0=>nx7919, A1=>nx7921, A2=>nx7923
   );
   ix7920 : aoi222 port map ( Y=>nx7919, A0=>que_out_15_3_10, A1=>nx9966, B0
      =>que_out_3_3_10, B1=>nx9992, C0=>que_out_23_3_10, C1=>nx9940);
   ix7922 : aoi22 port map ( Y=>nx7921, A0=>que_out_27_3_10, A1=>nx9914, B0
      =>que_out_4_3_10, B1=>nx9888);
   ix7924 : aoi22 port map ( Y=>nx7923, A0=>que_out_0_3_10, A1=>nx9836, B0=>
      que_out_2_3_10, B1=>nx9862);
   ix3019 : nand03 port map ( Y=>nx3018, A0=>nx7927, A1=>nx7929, A2=>nx7931
   );
   ix7928 : aoi222 port map ( Y=>nx7927, A0=>que_out_26_3_10, A1=>nx9810, B0
      =>que_out_14_3_10, B1=>nx9784, C0=>que_out_11_3_10, C1=>nx9758);
   ix7930 : aoi22 port map ( Y=>nx7929, A0=>que_out_13_3_10, A1=>nx9732, B0
      =>que_out_7_3_10, B1=>nx9706);
   ix7932 : aoi22 port map ( Y=>nx7931, A0=>que_out_12_3_10, A1=>nx9680, B0
      =>que_out_1_3_10, B1=>nx9654);
   ix3213 : or04 port map ( Y=>out_column_3_11, A0=>nx3208, A1=>nx3182, A2=>
      nx3154, A3=>nx3128);
   ix3209 : nand03 port map ( Y=>nx3208, A0=>nx7937, A1=>nx7939, A2=>nx7941
   );
   ix7938 : aoi222 port map ( Y=>nx7937, A0=>que_out_10_3_11, A1=>nx10304, 
      B0=>que_out_6_3_11, B1=>nx10356, C0=>que_out_9_3_11, C1=>nx10330);
   ix7940 : aoi22 port map ( Y=>nx7939, A0=>que_out_5_3_11, A1=>nx10252, B0
      =>que_out_18_3_11, B1=>nx10278);
   ix7942 : aoi22 port map ( Y=>nx7941, A0=>que_out_17_3_11, A1=>nx10226, B0
      =>que_out_20_3_11, B1=>nx10200);
   ix3183 : nand03 port map ( Y=>nx3182, A0=>nx7945, A1=>nx7947, A2=>nx7949
   );
   ix7946 : aoi222 port map ( Y=>nx7945, A0=>que_out_19_3_11, A1=>nx10174, 
      B0=>que_out_21_3_11, B1=>nx10148, C0=>que_out_8_3_11, C1=>nx10122);
   ix7948 : aoi22 port map ( Y=>nx7947, A0=>que_out_25_3_11, A1=>nx10070, B0
      =>que_out_16_3_11, B1=>nx10096);
   ix7950 : aoi22 port map ( Y=>nx7949, A0=>que_out_24_3_11, A1=>nx10044, B0
      =>que_out_22_3_11, B1=>nx10018);
   ix3155 : nand03 port map ( Y=>nx3154, A0=>nx7953, A1=>nx7955, A2=>nx7957
   );
   ix7954 : aoi222 port map ( Y=>nx7953, A0=>que_out_15_3_11, A1=>nx9966, B0
      =>que_out_3_3_11, B1=>nx9992, C0=>que_out_23_3_11, C1=>nx9940);
   ix7956 : aoi22 port map ( Y=>nx7955, A0=>que_out_27_3_11, A1=>nx9914, B0
      =>que_out_4_3_11, B1=>nx9888);
   ix7958 : aoi22 port map ( Y=>nx7957, A0=>que_out_0_3_11, A1=>nx9836, B0=>
      que_out_2_3_11, B1=>nx9862);
   ix3129 : nand03 port map ( Y=>nx3128, A0=>nx7961, A1=>nx7963, A2=>nx7965
   );
   ix7962 : aoi222 port map ( Y=>nx7961, A0=>que_out_26_3_11, A1=>nx9810, B0
      =>que_out_14_3_11, B1=>nx9784, C0=>que_out_11_3_11, C1=>nx9758);
   ix7964 : aoi22 port map ( Y=>nx7963, A0=>que_out_13_3_11, A1=>nx9732, B0
      =>que_out_7_3_11, B1=>nx9706);
   ix7966 : aoi22 port map ( Y=>nx7965, A0=>que_out_12_3_11, A1=>nx9680, B0
      =>que_out_1_3_11, B1=>nx9654);
   ix3323 : or04 port map ( Y=>out_column_3_12, A0=>nx3318, A1=>nx3292, A2=>
      nx3264, A3=>nx3238);
   ix3319 : nand03 port map ( Y=>nx3318, A0=>nx7971, A1=>nx7973, A2=>nx7975
   );
   ix7972 : aoi222 port map ( Y=>nx7971, A0=>que_out_10_3_12, A1=>nx10306, 
      B0=>que_out_6_3_12, B1=>nx10358, C0=>que_out_9_3_12, C1=>nx10332);
   ix7974 : aoi22 port map ( Y=>nx7973, A0=>que_out_5_3_12, A1=>nx10254, B0
      =>que_out_18_3_12, B1=>nx10280);
   ix7976 : aoi22 port map ( Y=>nx7975, A0=>que_out_17_3_12, A1=>nx10228, B0
      =>que_out_20_3_12, B1=>nx10202);
   ix3293 : nand03 port map ( Y=>nx3292, A0=>nx7979, A1=>nx7981, A2=>nx7983
   );
   ix7980 : aoi222 port map ( Y=>nx7979, A0=>que_out_19_3_12, A1=>nx10176, 
      B0=>que_out_21_3_12, B1=>nx10150, C0=>que_out_8_3_12, C1=>nx10124);
   ix7982 : aoi22 port map ( Y=>nx7981, A0=>que_out_25_3_12, A1=>nx10072, B0
      =>que_out_16_3_12, B1=>nx10098);
   ix7984 : aoi22 port map ( Y=>nx7983, A0=>que_out_24_3_12, A1=>nx10046, B0
      =>que_out_22_3_12, B1=>nx10020);
   ix3265 : nand03 port map ( Y=>nx3264, A0=>nx7987, A1=>nx7989, A2=>nx7991
   );
   ix7988 : aoi222 port map ( Y=>nx7987, A0=>que_out_15_3_12, A1=>nx9968, B0
      =>que_out_3_3_12, B1=>nx9994, C0=>que_out_23_3_12, C1=>nx9942);
   ix7990 : aoi22 port map ( Y=>nx7989, A0=>que_out_27_3_12, A1=>nx9916, B0
      =>que_out_4_3_12, B1=>nx9890);
   ix7992 : aoi22 port map ( Y=>nx7991, A0=>que_out_0_3_12, A1=>nx9838, B0=>
      que_out_2_3_12, B1=>nx9864);
   ix3239 : nand03 port map ( Y=>nx3238, A0=>nx7995, A1=>nx7997, A2=>nx7999
   );
   ix7996 : aoi222 port map ( Y=>nx7995, A0=>que_out_26_3_12, A1=>nx9812, B0
      =>que_out_14_3_12, B1=>nx9786, C0=>que_out_11_3_12, C1=>nx9760);
   ix7998 : aoi22 port map ( Y=>nx7997, A0=>que_out_13_3_12, A1=>nx9734, B0
      =>que_out_7_3_12, B1=>nx9708);
   ix8000 : aoi22 port map ( Y=>nx7999, A0=>que_out_12_3_12, A1=>nx9682, B0
      =>que_out_1_3_12, B1=>nx9656);
   ix3433 : or04 port map ( Y=>out_column_3_13, A0=>nx3428, A1=>nx3402, A2=>
      nx3374, A3=>nx3348);
   ix3429 : nand03 port map ( Y=>nx3428, A0=>nx8005, A1=>nx8007, A2=>nx8009
   );
   ix8006 : aoi222 port map ( Y=>nx8005, A0=>que_out_10_3_13, A1=>nx10306, 
      B0=>que_out_6_3_13, B1=>nx10358, C0=>que_out_9_3_13, C1=>nx10332);
   ix8008 : aoi22 port map ( Y=>nx8007, A0=>que_out_5_3_13, A1=>nx10254, B0
      =>que_out_18_3_13, B1=>nx10280);
   ix8010 : aoi22 port map ( Y=>nx8009, A0=>que_out_17_3_13, A1=>nx10228, B0
      =>que_out_20_3_13, B1=>nx10202);
   ix3403 : nand03 port map ( Y=>nx3402, A0=>nx8013, A1=>nx8015, A2=>nx8017
   );
   ix8014 : aoi222 port map ( Y=>nx8013, A0=>que_out_19_3_13, A1=>nx10176, 
      B0=>que_out_21_3_13, B1=>nx10150, C0=>que_out_8_3_13, C1=>nx10124);
   ix8016 : aoi22 port map ( Y=>nx8015, A0=>que_out_25_3_13, A1=>nx10072, B0
      =>que_out_16_3_13, B1=>nx10098);
   ix8018 : aoi22 port map ( Y=>nx8017, A0=>que_out_24_3_13, A1=>nx10046, B0
      =>que_out_22_3_13, B1=>nx10020);
   ix3375 : nand03 port map ( Y=>nx3374, A0=>nx8021, A1=>nx8023, A2=>nx8025
   );
   ix8022 : aoi222 port map ( Y=>nx8021, A0=>que_out_15_3_13, A1=>nx9968, B0
      =>que_out_3_3_13, B1=>nx9994, C0=>que_out_23_3_13, C1=>nx9942);
   ix8024 : aoi22 port map ( Y=>nx8023, A0=>que_out_27_3_13, A1=>nx9916, B0
      =>que_out_4_3_13, B1=>nx9890);
   ix8026 : aoi22 port map ( Y=>nx8025, A0=>que_out_0_3_13, A1=>nx9838, B0=>
      que_out_2_3_13, B1=>nx9864);
   ix3349 : nand03 port map ( Y=>nx3348, A0=>nx8029, A1=>nx8031, A2=>nx8033
   );
   ix8030 : aoi222 port map ( Y=>nx8029, A0=>que_out_26_3_13, A1=>nx9812, B0
      =>que_out_14_3_13, B1=>nx9786, C0=>que_out_11_3_13, C1=>nx9760);
   ix8032 : aoi22 port map ( Y=>nx8031, A0=>que_out_13_3_13, A1=>nx9734, B0
      =>que_out_7_3_13, B1=>nx9708);
   ix8034 : aoi22 port map ( Y=>nx8033, A0=>que_out_12_3_13, A1=>nx9682, B0
      =>que_out_1_3_13, B1=>nx9656);
   ix3543 : or04 port map ( Y=>out_column_3_14, A0=>nx3538, A1=>nx3512, A2=>
      nx3484, A3=>nx3458);
   ix3539 : nand03 port map ( Y=>nx3538, A0=>nx8039, A1=>nx8041, A2=>nx8043
   );
   ix8040 : aoi222 port map ( Y=>nx8039, A0=>que_out_10_3_14, A1=>nx10306, 
      B0=>que_out_6_3_14, B1=>nx10358, C0=>que_out_9_3_14, C1=>nx10332);
   ix8042 : aoi22 port map ( Y=>nx8041, A0=>que_out_5_3_14, A1=>nx10254, B0
      =>que_out_18_3_14, B1=>nx10280);
   ix8044 : aoi22 port map ( Y=>nx8043, A0=>que_out_17_3_14, A1=>nx10228, B0
      =>que_out_20_3_14, B1=>nx10202);
   ix3513 : nand03 port map ( Y=>nx3512, A0=>nx8047, A1=>nx8049, A2=>nx8051
   );
   ix8048 : aoi222 port map ( Y=>nx8047, A0=>que_out_19_3_14, A1=>nx10176, 
      B0=>que_out_21_3_14, B1=>nx10150, C0=>que_out_8_3_14, C1=>nx10124);
   ix8050 : aoi22 port map ( Y=>nx8049, A0=>que_out_25_3_14, A1=>nx10072, B0
      =>que_out_16_3_14, B1=>nx10098);
   ix8052 : aoi22 port map ( Y=>nx8051, A0=>que_out_24_3_14, A1=>nx10046, B0
      =>que_out_22_3_14, B1=>nx10020);
   ix3485 : nand03 port map ( Y=>nx3484, A0=>nx8055, A1=>nx8057, A2=>nx8059
   );
   ix8056 : aoi222 port map ( Y=>nx8055, A0=>que_out_15_3_14, A1=>nx9968, B0
      =>que_out_3_3_14, B1=>nx9994, C0=>que_out_23_3_14, C1=>nx9942);
   ix8058 : aoi22 port map ( Y=>nx8057, A0=>que_out_27_3_14, A1=>nx9916, B0
      =>que_out_4_3_14, B1=>nx9890);
   ix8060 : aoi22 port map ( Y=>nx8059, A0=>que_out_0_3_14, A1=>nx9838, B0=>
      que_out_2_3_14, B1=>nx9864);
   ix3459 : nand03 port map ( Y=>nx3458, A0=>nx8063, A1=>nx8065, A2=>nx8067
   );
   ix8064 : aoi222 port map ( Y=>nx8063, A0=>que_out_26_3_14, A1=>nx9812, B0
      =>que_out_14_3_14, B1=>nx9786, C0=>que_out_11_3_14, C1=>nx9760);
   ix8066 : aoi22 port map ( Y=>nx8065, A0=>que_out_13_3_14, A1=>nx9734, B0
      =>que_out_7_3_14, B1=>nx9708);
   ix8068 : aoi22 port map ( Y=>nx8067, A0=>que_out_12_3_14, A1=>nx9682, B0
      =>que_out_1_3_14, B1=>nx9656);
   ix3653 : or04 port map ( Y=>out_column_3_15, A0=>nx3648, A1=>nx3622, A2=>
      nx3594, A3=>nx3568);
   ix3649 : nand03 port map ( Y=>nx3648, A0=>nx8073, A1=>nx8075, A2=>nx8077
   );
   ix8074 : aoi222 port map ( Y=>nx8073, A0=>que_out_10_3_15, A1=>nx10306, 
      B0=>que_out_6_3_15, B1=>nx10358, C0=>que_out_9_3_15, C1=>nx10332);
   ix8076 : aoi22 port map ( Y=>nx8075, A0=>que_out_5_3_15, A1=>nx10254, B0
      =>que_out_18_3_15, B1=>nx10280);
   ix8078 : aoi22 port map ( Y=>nx8077, A0=>que_out_17_3_15, A1=>nx10228, B0
      =>que_out_20_3_15, B1=>nx10202);
   ix3623 : nand03 port map ( Y=>nx3622, A0=>nx8081, A1=>nx8083, A2=>nx8085
   );
   ix8082 : aoi222 port map ( Y=>nx8081, A0=>que_out_19_3_15, A1=>nx10176, 
      B0=>que_out_21_3_15, B1=>nx10150, C0=>que_out_8_3_15, C1=>nx10124);
   ix8084 : aoi22 port map ( Y=>nx8083, A0=>que_out_25_3_15, A1=>nx10072, B0
      =>que_out_16_3_15, B1=>nx10098);
   ix8086 : aoi22 port map ( Y=>nx8085, A0=>que_out_24_3_15, A1=>nx10046, B0
      =>que_out_22_3_15, B1=>nx10020);
   ix3595 : nand03 port map ( Y=>nx3594, A0=>nx8089, A1=>nx8091, A2=>nx8093
   );
   ix8090 : aoi222 port map ( Y=>nx8089, A0=>que_out_15_3_15, A1=>nx9968, B0
      =>que_out_3_3_15, B1=>nx9994, C0=>que_out_23_3_15, C1=>nx9942);
   ix8092 : aoi22 port map ( Y=>nx8091, A0=>que_out_27_3_15, A1=>nx9916, B0
      =>que_out_4_3_15, B1=>nx9890);
   ix8094 : aoi22 port map ( Y=>nx8093, A0=>que_out_0_3_15, A1=>nx9838, B0=>
      que_out_2_3_15, B1=>nx9864);
   ix3569 : nand03 port map ( Y=>nx3568, A0=>nx8097, A1=>nx8099, A2=>nx8101
   );
   ix8098 : aoi222 port map ( Y=>nx8097, A0=>que_out_26_3_15, A1=>nx9812, B0
      =>que_out_14_3_15, B1=>nx9786, C0=>que_out_11_3_15, C1=>nx9760);
   ix8100 : aoi22 port map ( Y=>nx8099, A0=>que_out_13_3_15, A1=>nx9734, B0
      =>que_out_7_3_15, B1=>nx9708);
   ix8102 : aoi22 port map ( Y=>nx8101, A0=>que_out_12_3_15, A1=>nx9682, B0
      =>que_out_1_3_15, B1=>nx9656);
   ix3763 : or04 port map ( Y=>out_column_2_0, A0=>nx3758, A1=>nx3732, A2=>
      nx3704, A3=>nx3678);
   ix3759 : nand03 port map ( Y=>nx3758, A0=>nx8107, A1=>nx8109, A2=>nx8111
   );
   ix8108 : aoi222 port map ( Y=>nx8107, A0=>que_out_10_2_0, A1=>nx10306, B0
      =>que_out_6_2_0, B1=>nx10358, C0=>que_out_9_2_0, C1=>nx10332);
   ix8110 : aoi22 port map ( Y=>nx8109, A0=>que_out_5_2_0, A1=>nx10254, B0=>
      que_out_18_2_0, B1=>nx10280);
   ix8112 : aoi22 port map ( Y=>nx8111, A0=>que_out_17_2_0, A1=>nx10228, B0
      =>que_out_20_2_0, B1=>nx10202);
   ix3733 : nand03 port map ( Y=>nx3732, A0=>nx8115, A1=>nx8117, A2=>nx8119
   );
   ix8116 : aoi222 port map ( Y=>nx8115, A0=>que_out_19_2_0, A1=>nx10176, B0
      =>que_out_21_2_0, B1=>nx10150, C0=>que_out_8_2_0, C1=>nx10124);
   ix8118 : aoi22 port map ( Y=>nx8117, A0=>que_out_25_2_0, A1=>nx10072, B0
      =>que_out_16_2_0, B1=>nx10098);
   ix8120 : aoi22 port map ( Y=>nx8119, A0=>que_out_24_2_0, A1=>nx10046, B0
      =>que_out_22_2_0, B1=>nx10020);
   ix3705 : nand03 port map ( Y=>nx3704, A0=>nx8123, A1=>nx8125, A2=>nx8127
   );
   ix8124 : aoi222 port map ( Y=>nx8123, A0=>que_out_15_2_0, A1=>nx9968, B0
      =>que_out_3_2_0, B1=>nx9994, C0=>que_out_23_2_0, C1=>nx9942);
   ix8126 : aoi22 port map ( Y=>nx8125, A0=>que_out_27_2_0, A1=>nx9916, B0=>
      que_out_4_2_0, B1=>nx9890);
   ix8128 : aoi22 port map ( Y=>nx8127, A0=>que_out_0_2_0, A1=>nx9838, B0=>
      que_out_2_2_0, B1=>nx9864);
   ix3679 : nand03 port map ( Y=>nx3678, A0=>nx8131, A1=>nx8133, A2=>nx8135
   );
   ix8132 : aoi222 port map ( Y=>nx8131, A0=>que_out_26_2_0, A1=>nx9812, B0
      =>que_out_14_2_0, B1=>nx9786, C0=>que_out_11_2_0, C1=>nx9760);
   ix8134 : aoi22 port map ( Y=>nx8133, A0=>que_out_13_2_0, A1=>nx9734, B0=>
      que_out_7_2_0, B1=>nx9708);
   ix8136 : aoi22 port map ( Y=>nx8135, A0=>que_out_12_2_0, A1=>nx9682, B0=>
      que_out_1_2_0, B1=>nx9656);
   ix3873 : or04 port map ( Y=>out_column_2_1, A0=>nx3868, A1=>nx3842, A2=>
      nx3814, A3=>nx3788);
   ix3869 : nand03 port map ( Y=>nx3868, A0=>nx8141, A1=>nx8143, A2=>nx8145
   );
   ix8142 : aoi222 port map ( Y=>nx8141, A0=>que_out_10_2_1, A1=>nx10306, B0
      =>que_out_6_2_1, B1=>nx10358, C0=>que_out_9_2_1, C1=>nx10332);
   ix8144 : aoi22 port map ( Y=>nx8143, A0=>que_out_5_2_1, A1=>nx10254, B0=>
      que_out_18_2_1, B1=>nx10280);
   ix8146 : aoi22 port map ( Y=>nx8145, A0=>que_out_17_2_1, A1=>nx10228, B0
      =>que_out_20_2_1, B1=>nx10202);
   ix3843 : nand03 port map ( Y=>nx3842, A0=>nx8149, A1=>nx8151, A2=>nx8153
   );
   ix8150 : aoi222 port map ( Y=>nx8149, A0=>que_out_19_2_1, A1=>nx10176, B0
      =>que_out_21_2_1, B1=>nx10150, C0=>que_out_8_2_1, C1=>nx10124);
   ix8152 : aoi22 port map ( Y=>nx8151, A0=>que_out_25_2_1, A1=>nx10072, B0
      =>que_out_16_2_1, B1=>nx10098);
   ix8154 : aoi22 port map ( Y=>nx8153, A0=>que_out_24_2_1, A1=>nx10046, B0
      =>que_out_22_2_1, B1=>nx10020);
   ix3815 : nand03 port map ( Y=>nx3814, A0=>nx8157, A1=>nx8159, A2=>nx8161
   );
   ix8158 : aoi222 port map ( Y=>nx8157, A0=>que_out_15_2_1, A1=>nx9968, B0
      =>que_out_3_2_1, B1=>nx9994, C0=>que_out_23_2_1, C1=>nx9942);
   ix8160 : aoi22 port map ( Y=>nx8159, A0=>que_out_27_2_1, A1=>nx9916, B0=>
      que_out_4_2_1, B1=>nx9890);
   ix8162 : aoi22 port map ( Y=>nx8161, A0=>que_out_0_2_1, A1=>nx9838, B0=>
      que_out_2_2_1, B1=>nx9864);
   ix3789 : nand03 port map ( Y=>nx3788, A0=>nx8165, A1=>nx8167, A2=>nx8169
   );
   ix8166 : aoi222 port map ( Y=>nx8165, A0=>que_out_26_2_1, A1=>nx9812, B0
      =>que_out_14_2_1, B1=>nx9786, C0=>que_out_11_2_1, C1=>nx9760);
   ix8168 : aoi22 port map ( Y=>nx8167, A0=>que_out_13_2_1, A1=>nx9734, B0=>
      que_out_7_2_1, B1=>nx9708);
   ix8170 : aoi22 port map ( Y=>nx8169, A0=>que_out_12_2_1, A1=>nx9682, B0=>
      que_out_1_2_1, B1=>nx9656);
   ix3983 : or04 port map ( Y=>out_column_2_2, A0=>nx3978, A1=>nx3952, A2=>
      nx3924, A3=>nx3898);
   ix3979 : nand03 port map ( Y=>nx3978, A0=>nx8175, A1=>nx8177, A2=>nx8179
   );
   ix8176 : aoi222 port map ( Y=>nx8175, A0=>que_out_10_2_2, A1=>nx10306, B0
      =>que_out_6_2_2, B1=>nx10358, C0=>que_out_9_2_2, C1=>nx10332);
   ix8178 : aoi22 port map ( Y=>nx8177, A0=>que_out_5_2_2, A1=>nx10254, B0=>
      que_out_18_2_2, B1=>nx10280);
   ix8180 : aoi22 port map ( Y=>nx8179, A0=>que_out_17_2_2, A1=>nx10228, B0
      =>que_out_20_2_2, B1=>nx10202);
   ix3953 : nand03 port map ( Y=>nx3952, A0=>nx8183, A1=>nx8185, A2=>nx8187
   );
   ix8184 : aoi222 port map ( Y=>nx8183, A0=>que_out_19_2_2, A1=>nx10176, B0
      =>que_out_21_2_2, B1=>nx10150, C0=>que_out_8_2_2, C1=>nx10124);
   ix8186 : aoi22 port map ( Y=>nx8185, A0=>que_out_25_2_2, A1=>nx10072, B0
      =>que_out_16_2_2, B1=>nx10098);
   ix8188 : aoi22 port map ( Y=>nx8187, A0=>que_out_24_2_2, A1=>nx10046, B0
      =>que_out_22_2_2, B1=>nx10020);
   ix3925 : nand03 port map ( Y=>nx3924, A0=>nx8191, A1=>nx8193, A2=>nx8195
   );
   ix8192 : aoi222 port map ( Y=>nx8191, A0=>que_out_15_2_2, A1=>nx9968, B0
      =>que_out_3_2_2, B1=>nx9994, C0=>que_out_23_2_2, C1=>nx9942);
   ix8194 : aoi22 port map ( Y=>nx8193, A0=>que_out_27_2_2, A1=>nx9916, B0=>
      que_out_4_2_2, B1=>nx9890);
   ix8196 : aoi22 port map ( Y=>nx8195, A0=>que_out_0_2_2, A1=>nx9838, B0=>
      que_out_2_2_2, B1=>nx9864);
   ix3899 : nand03 port map ( Y=>nx3898, A0=>nx8199, A1=>nx8201, A2=>nx8203
   );
   ix8200 : aoi222 port map ( Y=>nx8199, A0=>que_out_26_2_2, A1=>nx9812, B0
      =>que_out_14_2_2, B1=>nx9786, C0=>que_out_11_2_2, C1=>nx9760);
   ix8202 : aoi22 port map ( Y=>nx8201, A0=>que_out_13_2_2, A1=>nx9734, B0=>
      que_out_7_2_2, B1=>nx9708);
   ix8204 : aoi22 port map ( Y=>nx8203, A0=>que_out_12_2_2, A1=>nx9682, B0=>
      que_out_1_2_2, B1=>nx9656);
   ix4093 : or04 port map ( Y=>out_column_2_3, A0=>nx4088, A1=>nx4062, A2=>
      nx4034, A3=>nx4008);
   ix4089 : nand03 port map ( Y=>nx4088, A0=>nx8209, A1=>nx8211, A2=>nx8213
   );
   ix8210 : aoi222 port map ( Y=>nx8209, A0=>que_out_10_2_3, A1=>nx10308, B0
      =>que_out_6_2_3, B1=>nx10360, C0=>que_out_9_2_3, C1=>nx10334);
   ix8212 : aoi22 port map ( Y=>nx8211, A0=>que_out_5_2_3, A1=>nx10256, B0=>
      que_out_18_2_3, B1=>nx10282);
   ix8214 : aoi22 port map ( Y=>nx8213, A0=>que_out_17_2_3, A1=>nx10230, B0
      =>que_out_20_2_3, B1=>nx10204);
   ix4063 : nand03 port map ( Y=>nx4062, A0=>nx8217, A1=>nx8219, A2=>nx8221
   );
   ix8218 : aoi222 port map ( Y=>nx8217, A0=>que_out_19_2_3, A1=>nx10178, B0
      =>que_out_21_2_3, B1=>nx10152, C0=>que_out_8_2_3, C1=>nx10126);
   ix8220 : aoi22 port map ( Y=>nx8219, A0=>que_out_25_2_3, A1=>nx10074, B0
      =>que_out_16_2_3, B1=>nx10100);
   ix8222 : aoi22 port map ( Y=>nx8221, A0=>que_out_24_2_3, A1=>nx10048, B0
      =>que_out_22_2_3, B1=>nx10022);
   ix4035 : nand03 port map ( Y=>nx4034, A0=>nx8225, A1=>nx8227, A2=>nx8229
   );
   ix8226 : aoi222 port map ( Y=>nx8225, A0=>que_out_15_2_3, A1=>nx9970, B0
      =>que_out_3_2_3, B1=>nx9996, C0=>que_out_23_2_3, C1=>nx9944);
   ix8228 : aoi22 port map ( Y=>nx8227, A0=>que_out_27_2_3, A1=>nx9918, B0=>
      que_out_4_2_3, B1=>nx9892);
   ix8230 : aoi22 port map ( Y=>nx8229, A0=>que_out_0_2_3, A1=>nx9840, B0=>
      que_out_2_2_3, B1=>nx9866);
   ix4009 : nand03 port map ( Y=>nx4008, A0=>nx8233, A1=>nx8235, A2=>nx8237
   );
   ix8234 : aoi222 port map ( Y=>nx8233, A0=>que_out_26_2_3, A1=>nx9814, B0
      =>que_out_14_2_3, B1=>nx9788, C0=>que_out_11_2_3, C1=>nx9762);
   ix8236 : aoi22 port map ( Y=>nx8235, A0=>que_out_13_2_3, A1=>nx9736, B0=>
      que_out_7_2_3, B1=>nx9710);
   ix8238 : aoi22 port map ( Y=>nx8237, A0=>que_out_12_2_3, A1=>nx9684, B0=>
      que_out_1_2_3, B1=>nx9658);
   ix4203 : or04 port map ( Y=>out_column_2_4, A0=>nx4198, A1=>nx4172, A2=>
      nx4144, A3=>nx4118);
   ix4199 : nand03 port map ( Y=>nx4198, A0=>nx8243, A1=>nx8245, A2=>nx8247
   );
   ix8244 : aoi222 port map ( Y=>nx8243, A0=>que_out_10_2_4, A1=>nx10308, B0
      =>que_out_6_2_4, B1=>nx10360, C0=>que_out_9_2_4, C1=>nx10334);
   ix8246 : aoi22 port map ( Y=>nx8245, A0=>que_out_5_2_4, A1=>nx10256, B0=>
      que_out_18_2_4, B1=>nx10282);
   ix8248 : aoi22 port map ( Y=>nx8247, A0=>que_out_17_2_4, A1=>nx10230, B0
      =>que_out_20_2_4, B1=>nx10204);
   ix4173 : nand03 port map ( Y=>nx4172, A0=>nx8251, A1=>nx8253, A2=>nx8255
   );
   ix8252 : aoi222 port map ( Y=>nx8251, A0=>que_out_19_2_4, A1=>nx10178, B0
      =>que_out_21_2_4, B1=>nx10152, C0=>que_out_8_2_4, C1=>nx10126);
   ix8254 : aoi22 port map ( Y=>nx8253, A0=>que_out_25_2_4, A1=>nx10074, B0
      =>que_out_16_2_4, B1=>nx10100);
   ix8256 : aoi22 port map ( Y=>nx8255, A0=>que_out_24_2_4, A1=>nx10048, B0
      =>que_out_22_2_4, B1=>nx10022);
   ix4145 : nand03 port map ( Y=>nx4144, A0=>nx8259, A1=>nx8261, A2=>nx8263
   );
   ix8260 : aoi222 port map ( Y=>nx8259, A0=>que_out_15_2_4, A1=>nx9970, B0
      =>que_out_3_2_4, B1=>nx9996, C0=>que_out_23_2_4, C1=>nx9944);
   ix8262 : aoi22 port map ( Y=>nx8261, A0=>que_out_27_2_4, A1=>nx9918, B0=>
      que_out_4_2_4, B1=>nx9892);
   ix8264 : aoi22 port map ( Y=>nx8263, A0=>que_out_0_2_4, A1=>nx9840, B0=>
      que_out_2_2_4, B1=>nx9866);
   ix4119 : nand03 port map ( Y=>nx4118, A0=>nx8267, A1=>nx8269, A2=>nx8271
   );
   ix8268 : aoi222 port map ( Y=>nx8267, A0=>que_out_26_2_4, A1=>nx9814, B0
      =>que_out_14_2_4, B1=>nx9788, C0=>que_out_11_2_4, C1=>nx9762);
   ix8270 : aoi22 port map ( Y=>nx8269, A0=>que_out_13_2_4, A1=>nx9736, B0=>
      que_out_7_2_4, B1=>nx9710);
   ix8272 : aoi22 port map ( Y=>nx8271, A0=>que_out_12_2_4, A1=>nx9684, B0=>
      que_out_1_2_4, B1=>nx9658);
   ix4313 : or04 port map ( Y=>out_column_2_5, A0=>nx4308, A1=>nx4282, A2=>
      nx4254, A3=>nx4228);
   ix4309 : nand03 port map ( Y=>nx4308, A0=>nx8277, A1=>nx8279, A2=>nx8281
   );
   ix8278 : aoi222 port map ( Y=>nx8277, A0=>que_out_10_2_5, A1=>nx10308, B0
      =>que_out_6_2_5, B1=>nx10360, C0=>que_out_9_2_5, C1=>nx10334);
   ix8280 : aoi22 port map ( Y=>nx8279, A0=>que_out_5_2_5, A1=>nx10256, B0=>
      que_out_18_2_5, B1=>nx10282);
   ix8282 : aoi22 port map ( Y=>nx8281, A0=>que_out_17_2_5, A1=>nx10230, B0
      =>que_out_20_2_5, B1=>nx10204);
   ix4283 : nand03 port map ( Y=>nx4282, A0=>nx8285, A1=>nx8287, A2=>nx8289
   );
   ix8286 : aoi222 port map ( Y=>nx8285, A0=>que_out_19_2_5, A1=>nx10178, B0
      =>que_out_21_2_5, B1=>nx10152, C0=>que_out_8_2_5, C1=>nx10126);
   ix8288 : aoi22 port map ( Y=>nx8287, A0=>que_out_25_2_5, A1=>nx10074, B0
      =>que_out_16_2_5, B1=>nx10100);
   ix8290 : aoi22 port map ( Y=>nx8289, A0=>que_out_24_2_5, A1=>nx10048, B0
      =>que_out_22_2_5, B1=>nx10022);
   ix4255 : nand03 port map ( Y=>nx4254, A0=>nx8293, A1=>nx8295, A2=>nx8297
   );
   ix8294 : aoi222 port map ( Y=>nx8293, A0=>que_out_15_2_5, A1=>nx9970, B0
      =>que_out_3_2_5, B1=>nx9996, C0=>que_out_23_2_5, C1=>nx9944);
   ix8296 : aoi22 port map ( Y=>nx8295, A0=>que_out_27_2_5, A1=>nx9918, B0=>
      que_out_4_2_5, B1=>nx9892);
   ix8298 : aoi22 port map ( Y=>nx8297, A0=>que_out_0_2_5, A1=>nx9840, B0=>
      que_out_2_2_5, B1=>nx9866);
   ix4229 : nand03 port map ( Y=>nx4228, A0=>nx8301, A1=>nx8303, A2=>nx8305
   );
   ix8302 : aoi222 port map ( Y=>nx8301, A0=>que_out_26_2_5, A1=>nx9814, B0
      =>que_out_14_2_5, B1=>nx9788, C0=>que_out_11_2_5, C1=>nx9762);
   ix8304 : aoi22 port map ( Y=>nx8303, A0=>que_out_13_2_5, A1=>nx9736, B0=>
      que_out_7_2_5, B1=>nx9710);
   ix8306 : aoi22 port map ( Y=>nx8305, A0=>que_out_12_2_5, A1=>nx9684, B0=>
      que_out_1_2_5, B1=>nx9658);
   ix4423 : or04 port map ( Y=>out_column_2_6, A0=>nx4418, A1=>nx4392, A2=>
      nx4364, A3=>nx4338);
   ix4419 : nand03 port map ( Y=>nx4418, A0=>nx8311, A1=>nx8313, A2=>nx8315
   );
   ix8312 : aoi222 port map ( Y=>nx8311, A0=>que_out_10_2_6, A1=>nx10308, B0
      =>que_out_6_2_6, B1=>nx10360, C0=>que_out_9_2_6, C1=>nx10334);
   ix8314 : aoi22 port map ( Y=>nx8313, A0=>que_out_5_2_6, A1=>nx10256, B0=>
      que_out_18_2_6, B1=>nx10282);
   ix8316 : aoi22 port map ( Y=>nx8315, A0=>que_out_17_2_6, A1=>nx10230, B0
      =>que_out_20_2_6, B1=>nx10204);
   ix4393 : nand03 port map ( Y=>nx4392, A0=>nx8319, A1=>nx8321, A2=>nx8323
   );
   ix8320 : aoi222 port map ( Y=>nx8319, A0=>que_out_19_2_6, A1=>nx10178, B0
      =>que_out_21_2_6, B1=>nx10152, C0=>que_out_8_2_6, C1=>nx10126);
   ix8322 : aoi22 port map ( Y=>nx8321, A0=>que_out_25_2_6, A1=>nx10074, B0
      =>que_out_16_2_6, B1=>nx10100);
   ix8324 : aoi22 port map ( Y=>nx8323, A0=>que_out_24_2_6, A1=>nx10048, B0
      =>que_out_22_2_6, B1=>nx10022);
   ix4365 : nand03 port map ( Y=>nx4364, A0=>nx8327, A1=>nx8329, A2=>nx8331
   );
   ix8328 : aoi222 port map ( Y=>nx8327, A0=>que_out_15_2_6, A1=>nx9970, B0
      =>que_out_3_2_6, B1=>nx9996, C0=>que_out_23_2_6, C1=>nx9944);
   ix8330 : aoi22 port map ( Y=>nx8329, A0=>que_out_27_2_6, A1=>nx9918, B0=>
      que_out_4_2_6, B1=>nx9892);
   ix8332 : aoi22 port map ( Y=>nx8331, A0=>que_out_0_2_6, A1=>nx9840, B0=>
      que_out_2_2_6, B1=>nx9866);
   ix4339 : nand03 port map ( Y=>nx4338, A0=>nx8335, A1=>nx8337, A2=>nx8339
   );
   ix8336 : aoi222 port map ( Y=>nx8335, A0=>que_out_26_2_6, A1=>nx9814, B0
      =>que_out_14_2_6, B1=>nx9788, C0=>que_out_11_2_6, C1=>nx9762);
   ix8338 : aoi22 port map ( Y=>nx8337, A0=>que_out_13_2_6, A1=>nx9736, B0=>
      que_out_7_2_6, B1=>nx9710);
   ix8340 : aoi22 port map ( Y=>nx8339, A0=>que_out_12_2_6, A1=>nx9684, B0=>
      que_out_1_2_6, B1=>nx9658);
   ix4533 : or04 port map ( Y=>out_column_2_7, A0=>nx4528, A1=>nx4502, A2=>
      nx4474, A3=>nx4448);
   ix4529 : nand03 port map ( Y=>nx4528, A0=>nx8345, A1=>nx8347, A2=>nx8349
   );
   ix8346 : aoi222 port map ( Y=>nx8345, A0=>que_out_10_2_7, A1=>nx10308, B0
      =>que_out_6_2_7, B1=>nx10360, C0=>que_out_9_2_7, C1=>nx10334);
   ix8348 : aoi22 port map ( Y=>nx8347, A0=>que_out_5_2_7, A1=>nx10256, B0=>
      que_out_18_2_7, B1=>nx10282);
   ix8350 : aoi22 port map ( Y=>nx8349, A0=>que_out_17_2_7, A1=>nx10230, B0
      =>que_out_20_2_7, B1=>nx10204);
   ix4503 : nand03 port map ( Y=>nx4502, A0=>nx8353, A1=>nx8355, A2=>nx8357
   );
   ix8354 : aoi222 port map ( Y=>nx8353, A0=>que_out_19_2_7, A1=>nx10178, B0
      =>que_out_21_2_7, B1=>nx10152, C0=>que_out_8_2_7, C1=>nx10126);
   ix8356 : aoi22 port map ( Y=>nx8355, A0=>que_out_25_2_7, A1=>nx10074, B0
      =>que_out_16_2_7, B1=>nx10100);
   ix8358 : aoi22 port map ( Y=>nx8357, A0=>que_out_24_2_7, A1=>nx10048, B0
      =>que_out_22_2_7, B1=>nx10022);
   ix4475 : nand03 port map ( Y=>nx4474, A0=>nx8361, A1=>nx8363, A2=>nx8365
   );
   ix8362 : aoi222 port map ( Y=>nx8361, A0=>que_out_15_2_7, A1=>nx9970, B0
      =>que_out_3_2_7, B1=>nx9996, C0=>que_out_23_2_7, C1=>nx9944);
   ix8364 : aoi22 port map ( Y=>nx8363, A0=>que_out_27_2_7, A1=>nx9918, B0=>
      que_out_4_2_7, B1=>nx9892);
   ix8366 : aoi22 port map ( Y=>nx8365, A0=>que_out_0_2_7, A1=>nx9840, B0=>
      que_out_2_2_7, B1=>nx9866);
   ix4449 : nand03 port map ( Y=>nx4448, A0=>nx8369, A1=>nx8371, A2=>nx8373
   );
   ix8370 : aoi222 port map ( Y=>nx8369, A0=>que_out_26_2_7, A1=>nx9814, B0
      =>que_out_14_2_7, B1=>nx9788, C0=>que_out_11_2_7, C1=>nx9762);
   ix8372 : aoi22 port map ( Y=>nx8371, A0=>que_out_13_2_7, A1=>nx9736, B0=>
      que_out_7_2_7, B1=>nx9710);
   ix8374 : aoi22 port map ( Y=>nx8373, A0=>que_out_12_2_7, A1=>nx9684, B0=>
      que_out_1_2_7, B1=>nx9658);
   ix4643 : or04 port map ( Y=>out_column_2_8, A0=>nx4638, A1=>nx4612, A2=>
      nx4584, A3=>nx4558);
   ix4639 : nand03 port map ( Y=>nx4638, A0=>nx8379, A1=>nx8381, A2=>nx8383
   );
   ix8380 : aoi222 port map ( Y=>nx8379, A0=>que_out_10_2_8, A1=>nx10308, B0
      =>que_out_6_2_8, B1=>nx10360, C0=>que_out_9_2_8, C1=>nx10334);
   ix8382 : aoi22 port map ( Y=>nx8381, A0=>que_out_5_2_8, A1=>nx10256, B0=>
      que_out_18_2_8, B1=>nx10282);
   ix8384 : aoi22 port map ( Y=>nx8383, A0=>que_out_17_2_8, A1=>nx10230, B0
      =>que_out_20_2_8, B1=>nx10204);
   ix4613 : nand03 port map ( Y=>nx4612, A0=>nx8387, A1=>nx8389, A2=>nx8391
   );
   ix8388 : aoi222 port map ( Y=>nx8387, A0=>que_out_19_2_8, A1=>nx10178, B0
      =>que_out_21_2_8, B1=>nx10152, C0=>que_out_8_2_8, C1=>nx10126);
   ix8390 : aoi22 port map ( Y=>nx8389, A0=>que_out_25_2_8, A1=>nx10074, B0
      =>que_out_16_2_8, B1=>nx10100);
   ix8392 : aoi22 port map ( Y=>nx8391, A0=>que_out_24_2_8, A1=>nx10048, B0
      =>que_out_22_2_8, B1=>nx10022);
   ix4585 : nand03 port map ( Y=>nx4584, A0=>nx8395, A1=>nx8397, A2=>nx8399
   );
   ix8396 : aoi222 port map ( Y=>nx8395, A0=>que_out_15_2_8, A1=>nx9970, B0
      =>que_out_3_2_8, B1=>nx9996, C0=>que_out_23_2_8, C1=>nx9944);
   ix8398 : aoi22 port map ( Y=>nx8397, A0=>que_out_27_2_8, A1=>nx9918, B0=>
      que_out_4_2_8, B1=>nx9892);
   ix8400 : aoi22 port map ( Y=>nx8399, A0=>que_out_0_2_8, A1=>nx9840, B0=>
      que_out_2_2_8, B1=>nx9866);
   ix4559 : nand03 port map ( Y=>nx4558, A0=>nx8403, A1=>nx8405, A2=>nx8407
   );
   ix8404 : aoi222 port map ( Y=>nx8403, A0=>que_out_26_2_8, A1=>nx9814, B0
      =>que_out_14_2_8, B1=>nx9788, C0=>que_out_11_2_8, C1=>nx9762);
   ix8406 : aoi22 port map ( Y=>nx8405, A0=>que_out_13_2_8, A1=>nx9736, B0=>
      que_out_7_2_8, B1=>nx9710);
   ix8408 : aoi22 port map ( Y=>nx8407, A0=>que_out_12_2_8, A1=>nx9684, B0=>
      que_out_1_2_8, B1=>nx9658);
   ix4753 : or04 port map ( Y=>out_column_2_9, A0=>nx4748, A1=>nx4722, A2=>
      nx4694, A3=>nx4668);
   ix4749 : nand03 port map ( Y=>nx4748, A0=>nx8413, A1=>nx8415, A2=>nx8417
   );
   ix8414 : aoi222 port map ( Y=>nx8413, A0=>que_out_10_2_9, A1=>nx10308, B0
      =>que_out_6_2_9, B1=>nx10360, C0=>que_out_9_2_9, C1=>nx10334);
   ix8416 : aoi22 port map ( Y=>nx8415, A0=>que_out_5_2_9, A1=>nx10256, B0=>
      que_out_18_2_9, B1=>nx10282);
   ix8418 : aoi22 port map ( Y=>nx8417, A0=>que_out_17_2_9, A1=>nx10230, B0
      =>que_out_20_2_9, B1=>nx10204);
   ix4723 : nand03 port map ( Y=>nx4722, A0=>nx8421, A1=>nx8423, A2=>nx8425
   );
   ix8422 : aoi222 port map ( Y=>nx8421, A0=>que_out_19_2_9, A1=>nx10178, B0
      =>que_out_21_2_9, B1=>nx10152, C0=>que_out_8_2_9, C1=>nx10126);
   ix8424 : aoi22 port map ( Y=>nx8423, A0=>que_out_25_2_9, A1=>nx10074, B0
      =>que_out_16_2_9, B1=>nx10100);
   ix8426 : aoi22 port map ( Y=>nx8425, A0=>que_out_24_2_9, A1=>nx10048, B0
      =>que_out_22_2_9, B1=>nx10022);
   ix4695 : nand03 port map ( Y=>nx4694, A0=>nx8429, A1=>nx8431, A2=>nx8433
   );
   ix8430 : aoi222 port map ( Y=>nx8429, A0=>que_out_15_2_9, A1=>nx9970, B0
      =>que_out_3_2_9, B1=>nx9996, C0=>que_out_23_2_9, C1=>nx9944);
   ix8432 : aoi22 port map ( Y=>nx8431, A0=>que_out_27_2_9, A1=>nx9918, B0=>
      que_out_4_2_9, B1=>nx9892);
   ix8434 : aoi22 port map ( Y=>nx8433, A0=>que_out_0_2_9, A1=>nx9840, B0=>
      que_out_2_2_9, B1=>nx9866);
   ix4669 : nand03 port map ( Y=>nx4668, A0=>nx8437, A1=>nx8439, A2=>nx8441
   );
   ix8438 : aoi222 port map ( Y=>nx8437, A0=>que_out_26_2_9, A1=>nx9814, B0
      =>que_out_14_2_9, B1=>nx9788, C0=>que_out_11_2_9, C1=>nx9762);
   ix8440 : aoi22 port map ( Y=>nx8439, A0=>que_out_13_2_9, A1=>nx9736, B0=>
      que_out_7_2_9, B1=>nx9710);
   ix8442 : aoi22 port map ( Y=>nx8441, A0=>que_out_12_2_9, A1=>nx9684, B0=>
      que_out_1_2_9, B1=>nx9658);
   ix4863 : or04 port map ( Y=>out_column_2_10, A0=>nx4858, A1=>nx4832, A2=>
      nx4804, A3=>nx4778);
   ix4859 : nand03 port map ( Y=>nx4858, A0=>nx8447, A1=>nx8449, A2=>nx8451
   );
   ix8448 : aoi222 port map ( Y=>nx8447, A0=>que_out_10_2_10, A1=>nx10310, 
      B0=>que_out_6_2_10, B1=>nx10362, C0=>que_out_9_2_10, C1=>nx10336);
   ix8450 : aoi22 port map ( Y=>nx8449, A0=>que_out_5_2_10, A1=>nx10258, B0
      =>que_out_18_2_10, B1=>nx10284);
   ix8452 : aoi22 port map ( Y=>nx8451, A0=>que_out_17_2_10, A1=>nx10232, B0
      =>que_out_20_2_10, B1=>nx10206);
   ix4833 : nand03 port map ( Y=>nx4832, A0=>nx8455, A1=>nx8457, A2=>nx8459
   );
   ix8456 : aoi222 port map ( Y=>nx8455, A0=>que_out_19_2_10, A1=>nx10180, 
      B0=>que_out_21_2_10, B1=>nx10154, C0=>que_out_8_2_10, C1=>nx10128);
   ix8458 : aoi22 port map ( Y=>nx8457, A0=>que_out_25_2_10, A1=>nx10076, B0
      =>que_out_16_2_10, B1=>nx10102);
   ix8460 : aoi22 port map ( Y=>nx8459, A0=>que_out_24_2_10, A1=>nx10050, B0
      =>que_out_22_2_10, B1=>nx10024);
   ix4805 : nand03 port map ( Y=>nx4804, A0=>nx8463, A1=>nx8465, A2=>nx8467
   );
   ix8464 : aoi222 port map ( Y=>nx8463, A0=>que_out_15_2_10, A1=>nx9972, B0
      =>que_out_3_2_10, B1=>nx9998, C0=>que_out_23_2_10, C1=>nx9946);
   ix8466 : aoi22 port map ( Y=>nx8465, A0=>que_out_27_2_10, A1=>nx9920, B0
      =>que_out_4_2_10, B1=>nx9894);
   ix8468 : aoi22 port map ( Y=>nx8467, A0=>que_out_0_2_10, A1=>nx9842, B0=>
      que_out_2_2_10, B1=>nx9868);
   ix4779 : nand03 port map ( Y=>nx4778, A0=>nx8471, A1=>nx8473, A2=>nx8475
   );
   ix8472 : aoi222 port map ( Y=>nx8471, A0=>que_out_26_2_10, A1=>nx9816, B0
      =>que_out_14_2_10, B1=>nx9790, C0=>que_out_11_2_10, C1=>nx9764);
   ix8474 : aoi22 port map ( Y=>nx8473, A0=>que_out_13_2_10, A1=>nx9738, B0
      =>que_out_7_2_10, B1=>nx9712);
   ix8476 : aoi22 port map ( Y=>nx8475, A0=>que_out_12_2_10, A1=>nx9686, B0
      =>que_out_1_2_10, B1=>nx9660);
   ix4973 : or04 port map ( Y=>out_column_2_11, A0=>nx4968, A1=>nx4942, A2=>
      nx4914, A3=>nx4888);
   ix4969 : nand03 port map ( Y=>nx4968, A0=>nx8481, A1=>nx8483, A2=>nx8485
   );
   ix8482 : aoi222 port map ( Y=>nx8481, A0=>que_out_10_2_11, A1=>nx10310, 
      B0=>que_out_6_2_11, B1=>nx10362, C0=>que_out_9_2_11, C1=>nx10336);
   ix8484 : aoi22 port map ( Y=>nx8483, A0=>que_out_5_2_11, A1=>nx10258, B0
      =>que_out_18_2_11, B1=>nx10284);
   ix8486 : aoi22 port map ( Y=>nx8485, A0=>que_out_17_2_11, A1=>nx10232, B0
      =>que_out_20_2_11, B1=>nx10206);
   ix4943 : nand03 port map ( Y=>nx4942, A0=>nx8489, A1=>nx8491, A2=>nx8493
   );
   ix8490 : aoi222 port map ( Y=>nx8489, A0=>que_out_19_2_11, A1=>nx10180, 
      B0=>que_out_21_2_11, B1=>nx10154, C0=>que_out_8_2_11, C1=>nx10128);
   ix8492 : aoi22 port map ( Y=>nx8491, A0=>que_out_25_2_11, A1=>nx10076, B0
      =>que_out_16_2_11, B1=>nx10102);
   ix8494 : aoi22 port map ( Y=>nx8493, A0=>que_out_24_2_11, A1=>nx10050, B0
      =>que_out_22_2_11, B1=>nx10024);
   ix4915 : nand03 port map ( Y=>nx4914, A0=>nx8497, A1=>nx8499, A2=>nx8501
   );
   ix8498 : aoi222 port map ( Y=>nx8497, A0=>que_out_15_2_11, A1=>nx9972, B0
      =>que_out_3_2_11, B1=>nx9998, C0=>que_out_23_2_11, C1=>nx9946);
   ix8500 : aoi22 port map ( Y=>nx8499, A0=>que_out_27_2_11, A1=>nx9920, B0
      =>que_out_4_2_11, B1=>nx9894);
   ix8502 : aoi22 port map ( Y=>nx8501, A0=>que_out_0_2_11, A1=>nx9842, B0=>
      que_out_2_2_11, B1=>nx9868);
   ix4889 : nand03 port map ( Y=>nx4888, A0=>nx8505, A1=>nx8507, A2=>nx8509
   );
   ix8506 : aoi222 port map ( Y=>nx8505, A0=>que_out_26_2_11, A1=>nx9816, B0
      =>que_out_14_2_11, B1=>nx9790, C0=>que_out_11_2_11, C1=>nx9764);
   ix8508 : aoi22 port map ( Y=>nx8507, A0=>que_out_13_2_11, A1=>nx9738, B0
      =>que_out_7_2_11, B1=>nx9712);
   ix8510 : aoi22 port map ( Y=>nx8509, A0=>que_out_12_2_11, A1=>nx9686, B0
      =>que_out_1_2_11, B1=>nx9660);
   ix5083 : or04 port map ( Y=>out_column_2_12, A0=>nx5078, A1=>nx5052, A2=>
      nx5024, A3=>nx4998);
   ix5079 : nand03 port map ( Y=>nx5078, A0=>nx8515, A1=>nx8517, A2=>nx8519
   );
   ix8516 : aoi222 port map ( Y=>nx8515, A0=>que_out_10_2_12, A1=>nx10310, 
      B0=>que_out_6_2_12, B1=>nx10362, C0=>que_out_9_2_12, C1=>nx10336);
   ix8518 : aoi22 port map ( Y=>nx8517, A0=>que_out_5_2_12, A1=>nx10258, B0
      =>que_out_18_2_12, B1=>nx10284);
   ix8520 : aoi22 port map ( Y=>nx8519, A0=>que_out_17_2_12, A1=>nx10232, B0
      =>que_out_20_2_12, B1=>nx10206);
   ix5053 : nand03 port map ( Y=>nx5052, A0=>nx8523, A1=>nx8525, A2=>nx8527
   );
   ix8524 : aoi222 port map ( Y=>nx8523, A0=>que_out_19_2_12, A1=>nx10180, 
      B0=>que_out_21_2_12, B1=>nx10154, C0=>que_out_8_2_12, C1=>nx10128);
   ix8526 : aoi22 port map ( Y=>nx8525, A0=>que_out_25_2_12, A1=>nx10076, B0
      =>que_out_16_2_12, B1=>nx10102);
   ix8528 : aoi22 port map ( Y=>nx8527, A0=>que_out_24_2_12, A1=>nx10050, B0
      =>que_out_22_2_12, B1=>nx10024);
   ix5025 : nand03 port map ( Y=>nx5024, A0=>nx8531, A1=>nx8533, A2=>nx8535
   );
   ix8532 : aoi222 port map ( Y=>nx8531, A0=>que_out_15_2_12, A1=>nx9972, B0
      =>que_out_3_2_12, B1=>nx9998, C0=>que_out_23_2_12, C1=>nx9946);
   ix8534 : aoi22 port map ( Y=>nx8533, A0=>que_out_27_2_12, A1=>nx9920, B0
      =>que_out_4_2_12, B1=>nx9894);
   ix8536 : aoi22 port map ( Y=>nx8535, A0=>que_out_0_2_12, A1=>nx9842, B0=>
      que_out_2_2_12, B1=>nx9868);
   ix4999 : nand03 port map ( Y=>nx4998, A0=>nx8539, A1=>nx8541, A2=>nx8543
   );
   ix8540 : aoi222 port map ( Y=>nx8539, A0=>que_out_26_2_12, A1=>nx9816, B0
      =>que_out_14_2_12, B1=>nx9790, C0=>que_out_11_2_12, C1=>nx9764);
   ix8542 : aoi22 port map ( Y=>nx8541, A0=>que_out_13_2_12, A1=>nx9738, B0
      =>que_out_7_2_12, B1=>nx9712);
   ix8544 : aoi22 port map ( Y=>nx8543, A0=>que_out_12_2_12, A1=>nx9686, B0
      =>que_out_1_2_12, B1=>nx9660);
   ix5193 : or04 port map ( Y=>out_column_2_13, A0=>nx5188, A1=>nx5162, A2=>
      nx5134, A3=>nx5108);
   ix5189 : nand03 port map ( Y=>nx5188, A0=>nx8549, A1=>nx8551, A2=>nx8553
   );
   ix8550 : aoi222 port map ( Y=>nx8549, A0=>que_out_10_2_13, A1=>nx10310, 
      B0=>que_out_6_2_13, B1=>nx10362, C0=>que_out_9_2_13, C1=>nx10336);
   ix8552 : aoi22 port map ( Y=>nx8551, A0=>que_out_5_2_13, A1=>nx10258, B0
      =>que_out_18_2_13, B1=>nx10284);
   ix8554 : aoi22 port map ( Y=>nx8553, A0=>que_out_17_2_13, A1=>nx10232, B0
      =>que_out_20_2_13, B1=>nx10206);
   ix5163 : nand03 port map ( Y=>nx5162, A0=>nx8557, A1=>nx8559, A2=>nx8561
   );
   ix8558 : aoi222 port map ( Y=>nx8557, A0=>que_out_19_2_13, A1=>nx10180, 
      B0=>que_out_21_2_13, B1=>nx10154, C0=>que_out_8_2_13, C1=>nx10128);
   ix8560 : aoi22 port map ( Y=>nx8559, A0=>que_out_25_2_13, A1=>nx10076, B0
      =>que_out_16_2_13, B1=>nx10102);
   ix8562 : aoi22 port map ( Y=>nx8561, A0=>que_out_24_2_13, A1=>nx10050, B0
      =>que_out_22_2_13, B1=>nx10024);
   ix5135 : nand03 port map ( Y=>nx5134, A0=>nx8565, A1=>nx8567, A2=>nx8569
   );
   ix8566 : aoi222 port map ( Y=>nx8565, A0=>que_out_15_2_13, A1=>nx9972, B0
      =>que_out_3_2_13, B1=>nx9998, C0=>que_out_23_2_13, C1=>nx9946);
   ix8568 : aoi22 port map ( Y=>nx8567, A0=>que_out_27_2_13, A1=>nx9920, B0
      =>que_out_4_2_13, B1=>nx9894);
   ix8570 : aoi22 port map ( Y=>nx8569, A0=>que_out_0_2_13, A1=>nx9842, B0=>
      que_out_2_2_13, B1=>nx9868);
   ix5109 : nand03 port map ( Y=>nx5108, A0=>nx8573, A1=>nx8575, A2=>nx8577
   );
   ix8574 : aoi222 port map ( Y=>nx8573, A0=>que_out_26_2_13, A1=>nx9816, B0
      =>que_out_14_2_13, B1=>nx9790, C0=>que_out_11_2_13, C1=>nx9764);
   ix8576 : aoi22 port map ( Y=>nx8575, A0=>que_out_13_2_13, A1=>nx9738, B0
      =>que_out_7_2_13, B1=>nx9712);
   ix8578 : aoi22 port map ( Y=>nx8577, A0=>que_out_12_2_13, A1=>nx9686, B0
      =>que_out_1_2_13, B1=>nx9660);
   ix5303 : or04 port map ( Y=>out_column_2_14, A0=>nx5298, A1=>nx5272, A2=>
      nx5244, A3=>nx5218);
   ix5299 : nand03 port map ( Y=>nx5298, A0=>nx8583, A1=>nx8585, A2=>nx8587
   );
   ix8584 : aoi222 port map ( Y=>nx8583, A0=>que_out_10_2_14, A1=>nx10310, 
      B0=>que_out_6_2_14, B1=>nx10362, C0=>que_out_9_2_14, C1=>nx10336);
   ix8586 : aoi22 port map ( Y=>nx8585, A0=>que_out_5_2_14, A1=>nx10258, B0
      =>que_out_18_2_14, B1=>nx10284);
   ix8588 : aoi22 port map ( Y=>nx8587, A0=>que_out_17_2_14, A1=>nx10232, B0
      =>que_out_20_2_14, B1=>nx10206);
   ix5273 : nand03 port map ( Y=>nx5272, A0=>nx8591, A1=>nx8593, A2=>nx8595
   );
   ix8592 : aoi222 port map ( Y=>nx8591, A0=>que_out_19_2_14, A1=>nx10180, 
      B0=>que_out_21_2_14, B1=>nx10154, C0=>que_out_8_2_14, C1=>nx10128);
   ix8594 : aoi22 port map ( Y=>nx8593, A0=>que_out_25_2_14, A1=>nx10076, B0
      =>que_out_16_2_14, B1=>nx10102);
   ix8596 : aoi22 port map ( Y=>nx8595, A0=>que_out_24_2_14, A1=>nx10050, B0
      =>que_out_22_2_14, B1=>nx10024);
   ix5245 : nand03 port map ( Y=>nx5244, A0=>nx8599, A1=>nx8601, A2=>nx8603
   );
   ix8600 : aoi222 port map ( Y=>nx8599, A0=>que_out_15_2_14, A1=>nx9972, B0
      =>que_out_3_2_14, B1=>nx9998, C0=>que_out_23_2_14, C1=>nx9946);
   ix8602 : aoi22 port map ( Y=>nx8601, A0=>que_out_27_2_14, A1=>nx9920, B0
      =>que_out_4_2_14, B1=>nx9894);
   ix8604 : aoi22 port map ( Y=>nx8603, A0=>que_out_0_2_14, A1=>nx9842, B0=>
      que_out_2_2_14, B1=>nx9868);
   ix5219 : nand03 port map ( Y=>nx5218, A0=>nx8607, A1=>nx8609, A2=>nx8611
   );
   ix8608 : aoi222 port map ( Y=>nx8607, A0=>que_out_26_2_14, A1=>nx9816, B0
      =>que_out_14_2_14, B1=>nx9790, C0=>que_out_11_2_14, C1=>nx9764);
   ix8610 : aoi22 port map ( Y=>nx8609, A0=>que_out_13_2_14, A1=>nx9738, B0
      =>que_out_7_2_14, B1=>nx9712);
   ix8612 : aoi22 port map ( Y=>nx8611, A0=>que_out_12_2_14, A1=>nx9686, B0
      =>que_out_1_2_14, B1=>nx9660);
   ix5413 : or04 port map ( Y=>out_column_2_15, A0=>nx5408, A1=>nx5382, A2=>
      nx5354, A3=>nx5328);
   ix5409 : nand03 port map ( Y=>nx5408, A0=>nx8617, A1=>nx8619, A2=>nx8621
   );
   ix8618 : aoi222 port map ( Y=>nx8617, A0=>que_out_10_2_15, A1=>nx10310, 
      B0=>que_out_6_2_15, B1=>nx10362, C0=>que_out_9_2_15, C1=>nx10336);
   ix8620 : aoi22 port map ( Y=>nx8619, A0=>que_out_5_2_15, A1=>nx10258, B0
      =>que_out_18_2_15, B1=>nx10284);
   ix8622 : aoi22 port map ( Y=>nx8621, A0=>que_out_17_2_15, A1=>nx10232, B0
      =>que_out_20_2_15, B1=>nx10206);
   ix5383 : nand03 port map ( Y=>nx5382, A0=>nx8625, A1=>nx8627, A2=>nx8629
   );
   ix8626 : aoi222 port map ( Y=>nx8625, A0=>que_out_19_2_15, A1=>nx10180, 
      B0=>que_out_21_2_15, B1=>nx10154, C0=>que_out_8_2_15, C1=>nx10128);
   ix8628 : aoi22 port map ( Y=>nx8627, A0=>que_out_25_2_15, A1=>nx10076, B0
      =>que_out_16_2_15, B1=>nx10102);
   ix8630 : aoi22 port map ( Y=>nx8629, A0=>que_out_24_2_15, A1=>nx10050, B0
      =>que_out_22_2_15, B1=>nx10024);
   ix5355 : nand03 port map ( Y=>nx5354, A0=>nx8633, A1=>nx8635, A2=>nx8637
   );
   ix8634 : aoi222 port map ( Y=>nx8633, A0=>que_out_15_2_15, A1=>nx9972, B0
      =>que_out_3_2_15, B1=>nx9998, C0=>que_out_23_2_15, C1=>nx9946);
   ix8636 : aoi22 port map ( Y=>nx8635, A0=>que_out_27_2_15, A1=>nx9920, B0
      =>que_out_4_2_15, B1=>nx9894);
   ix8638 : aoi22 port map ( Y=>nx8637, A0=>que_out_0_2_15, A1=>nx9842, B0=>
      que_out_2_2_15, B1=>nx9868);
   ix5329 : nand03 port map ( Y=>nx5328, A0=>nx8641, A1=>nx8643, A2=>nx8645
   );
   ix8642 : aoi222 port map ( Y=>nx8641, A0=>que_out_26_2_15, A1=>nx9816, B0
      =>que_out_14_2_15, B1=>nx9790, C0=>que_out_11_2_15, C1=>nx9764);
   ix8644 : aoi22 port map ( Y=>nx8643, A0=>que_out_13_2_15, A1=>nx9738, B0
      =>que_out_7_2_15, B1=>nx9712);
   ix8646 : aoi22 port map ( Y=>nx8645, A0=>que_out_12_2_15, A1=>nx9686, B0
      =>que_out_1_2_15, B1=>nx9660);
   ix5523 : or04 port map ( Y=>out_column_1_0, A0=>nx5518, A1=>nx5492, A2=>
      nx5464, A3=>nx5438);
   ix5519 : nand03 port map ( Y=>nx5518, A0=>nx8651, A1=>nx8653, A2=>nx8655
   );
   ix8652 : aoi222 port map ( Y=>nx8651, A0=>que_out_10_1_0, A1=>nx10310, B0
      =>que_out_6_1_0, B1=>nx10362, C0=>que_out_9_1_0, C1=>nx10336);
   ix8654 : aoi22 port map ( Y=>nx8653, A0=>que_out_5_1_0, A1=>nx10258, B0=>
      que_out_18_1_0, B1=>nx10284);
   ix8656 : aoi22 port map ( Y=>nx8655, A0=>que_out_17_1_0, A1=>nx10232, B0
      =>que_out_20_1_0, B1=>nx10206);
   ix5493 : nand03 port map ( Y=>nx5492, A0=>nx8659, A1=>nx8661, A2=>nx8663
   );
   ix8660 : aoi222 port map ( Y=>nx8659, A0=>que_out_19_1_0, A1=>nx10180, B0
      =>que_out_21_1_0, B1=>nx10154, C0=>que_out_8_1_0, C1=>nx10128);
   ix8662 : aoi22 port map ( Y=>nx8661, A0=>que_out_25_1_0, A1=>nx10076, B0
      =>que_out_16_1_0, B1=>nx10102);
   ix8664 : aoi22 port map ( Y=>nx8663, A0=>que_out_24_1_0, A1=>nx10050, B0
      =>que_out_22_1_0, B1=>nx10024);
   ix5465 : nand03 port map ( Y=>nx5464, A0=>nx8667, A1=>nx8669, A2=>nx8671
   );
   ix8668 : aoi222 port map ( Y=>nx8667, A0=>que_out_15_1_0, A1=>nx9972, B0
      =>que_out_3_1_0, B1=>nx9998, C0=>que_out_23_1_0, C1=>nx9946);
   ix8670 : aoi22 port map ( Y=>nx8669, A0=>que_out_27_1_0, A1=>nx9920, B0=>
      que_out_4_1_0, B1=>nx9894);
   ix8672 : aoi22 port map ( Y=>nx8671, A0=>que_out_0_1_0, A1=>nx9842, B0=>
      que_out_2_1_0, B1=>nx9868);
   ix5439 : nand03 port map ( Y=>nx5438, A0=>nx8675, A1=>nx8677, A2=>nx8679
   );
   ix8676 : aoi222 port map ( Y=>nx8675, A0=>que_out_26_1_0, A1=>nx9816, B0
      =>que_out_14_1_0, B1=>nx9790, C0=>que_out_11_1_0, C1=>nx9764);
   ix8678 : aoi22 port map ( Y=>nx8677, A0=>que_out_13_1_0, A1=>nx9738, B0=>
      que_out_7_1_0, B1=>nx9712);
   ix8680 : aoi22 port map ( Y=>nx8679, A0=>que_out_12_1_0, A1=>nx9686, B0=>
      que_out_1_1_0, B1=>nx9660);
   ix5633 : or04 port map ( Y=>out_column_1_1, A0=>nx5628, A1=>nx5602, A2=>
      nx5574, A3=>nx5548);
   ix5629 : nand03 port map ( Y=>nx5628, A0=>nx8685, A1=>nx8687, A2=>nx8689
   );
   ix8686 : aoi222 port map ( Y=>nx8685, A0=>que_out_10_1_1, A1=>nx10312, B0
      =>que_out_6_1_1, B1=>nx10364, C0=>que_out_9_1_1, C1=>nx10338);
   ix8688 : aoi22 port map ( Y=>nx8687, A0=>que_out_5_1_1, A1=>nx10260, B0=>
      que_out_18_1_1, B1=>nx10286);
   ix8690 : aoi22 port map ( Y=>nx8689, A0=>que_out_17_1_1, A1=>nx10234, B0
      =>que_out_20_1_1, B1=>nx10208);
   ix5603 : nand03 port map ( Y=>nx5602, A0=>nx8693, A1=>nx8695, A2=>nx8697
   );
   ix8694 : aoi222 port map ( Y=>nx8693, A0=>que_out_19_1_1, A1=>nx10182, B0
      =>que_out_21_1_1, B1=>nx10156, C0=>que_out_8_1_1, C1=>nx10130);
   ix8696 : aoi22 port map ( Y=>nx8695, A0=>que_out_25_1_1, A1=>nx10078, B0
      =>que_out_16_1_1, B1=>nx10104);
   ix8698 : aoi22 port map ( Y=>nx8697, A0=>que_out_24_1_1, A1=>nx10052, B0
      =>que_out_22_1_1, B1=>nx10026);
   ix5575 : nand03 port map ( Y=>nx5574, A0=>nx8701, A1=>nx8703, A2=>nx8705
   );
   ix8702 : aoi222 port map ( Y=>nx8701, A0=>que_out_15_1_1, A1=>nx9974, B0
      =>que_out_3_1_1, B1=>nx10000, C0=>que_out_23_1_1, C1=>nx9948);
   ix8704 : aoi22 port map ( Y=>nx8703, A0=>que_out_27_1_1, A1=>nx9922, B0=>
      que_out_4_1_1, B1=>nx9896);
   ix8706 : aoi22 port map ( Y=>nx8705, A0=>que_out_0_1_1, A1=>nx9844, B0=>
      que_out_2_1_1, B1=>nx9870);
   ix5549 : nand03 port map ( Y=>nx5548, A0=>nx8709, A1=>nx8711, A2=>nx8713
   );
   ix8710 : aoi222 port map ( Y=>nx8709, A0=>que_out_26_1_1, A1=>nx9818, B0
      =>que_out_14_1_1, B1=>nx9792, C0=>que_out_11_1_1, C1=>nx9766);
   ix8712 : aoi22 port map ( Y=>nx8711, A0=>que_out_13_1_1, A1=>nx9740, B0=>
      que_out_7_1_1, B1=>nx9714);
   ix8714 : aoi22 port map ( Y=>nx8713, A0=>que_out_12_1_1, A1=>nx9688, B0=>
      que_out_1_1_1, B1=>nx9662);
   ix5743 : or04 port map ( Y=>out_column_1_2, A0=>nx5738, A1=>nx5712, A2=>
      nx5684, A3=>nx5658);
   ix5739 : nand03 port map ( Y=>nx5738, A0=>nx8719, A1=>nx8721, A2=>nx8723
   );
   ix8720 : aoi222 port map ( Y=>nx8719, A0=>que_out_10_1_2, A1=>nx10312, B0
      =>que_out_6_1_2, B1=>nx10364, C0=>que_out_9_1_2, C1=>nx10338);
   ix8722 : aoi22 port map ( Y=>nx8721, A0=>que_out_5_1_2, A1=>nx10260, B0=>
      que_out_18_1_2, B1=>nx10286);
   ix8724 : aoi22 port map ( Y=>nx8723, A0=>que_out_17_1_2, A1=>nx10234, B0
      =>que_out_20_1_2, B1=>nx10208);
   ix5713 : nand03 port map ( Y=>nx5712, A0=>nx8727, A1=>nx8729, A2=>nx8731
   );
   ix8728 : aoi222 port map ( Y=>nx8727, A0=>que_out_19_1_2, A1=>nx10182, B0
      =>que_out_21_1_2, B1=>nx10156, C0=>que_out_8_1_2, C1=>nx10130);
   ix8730 : aoi22 port map ( Y=>nx8729, A0=>que_out_25_1_2, A1=>nx10078, B0
      =>que_out_16_1_2, B1=>nx10104);
   ix8732 : aoi22 port map ( Y=>nx8731, A0=>que_out_24_1_2, A1=>nx10052, B0
      =>que_out_22_1_2, B1=>nx10026);
   ix5685 : nand03 port map ( Y=>nx5684, A0=>nx8735, A1=>nx8737, A2=>nx8739
   );
   ix8736 : aoi222 port map ( Y=>nx8735, A0=>que_out_15_1_2, A1=>nx9974, B0
      =>que_out_3_1_2, B1=>nx10000, C0=>que_out_23_1_2, C1=>nx9948);
   ix8738 : aoi22 port map ( Y=>nx8737, A0=>que_out_27_1_2, A1=>nx9922, B0=>
      que_out_4_1_2, B1=>nx9896);
   ix8740 : aoi22 port map ( Y=>nx8739, A0=>que_out_0_1_2, A1=>nx9844, B0=>
      que_out_2_1_2, B1=>nx9870);
   ix5659 : nand03 port map ( Y=>nx5658, A0=>nx8743, A1=>nx8745, A2=>nx8747
   );
   ix8744 : aoi222 port map ( Y=>nx8743, A0=>que_out_26_1_2, A1=>nx9818, B0
      =>que_out_14_1_2, B1=>nx9792, C0=>que_out_11_1_2, C1=>nx9766);
   ix8746 : aoi22 port map ( Y=>nx8745, A0=>que_out_13_1_2, A1=>nx9740, B0=>
      que_out_7_1_2, B1=>nx9714);
   ix8748 : aoi22 port map ( Y=>nx8747, A0=>que_out_12_1_2, A1=>nx9688, B0=>
      que_out_1_1_2, B1=>nx9662);
   ix5853 : or04 port map ( Y=>out_column_1_3, A0=>nx5848, A1=>nx5822, A2=>
      nx5794, A3=>nx5768);
   ix5849 : nand03 port map ( Y=>nx5848, A0=>nx8753, A1=>nx8755, A2=>nx8757
   );
   ix8754 : aoi222 port map ( Y=>nx8753, A0=>que_out_10_1_3, A1=>nx10312, B0
      =>que_out_6_1_3, B1=>nx10364, C0=>que_out_9_1_3, C1=>nx10338);
   ix8756 : aoi22 port map ( Y=>nx8755, A0=>que_out_5_1_3, A1=>nx10260, B0=>
      que_out_18_1_3, B1=>nx10286);
   ix8758 : aoi22 port map ( Y=>nx8757, A0=>que_out_17_1_3, A1=>nx10234, B0
      =>que_out_20_1_3, B1=>nx10208);
   ix5823 : nand03 port map ( Y=>nx5822, A0=>nx8761, A1=>nx8763, A2=>nx8765
   );
   ix8762 : aoi222 port map ( Y=>nx8761, A0=>que_out_19_1_3, A1=>nx10182, B0
      =>que_out_21_1_3, B1=>nx10156, C0=>que_out_8_1_3, C1=>nx10130);
   ix8764 : aoi22 port map ( Y=>nx8763, A0=>que_out_25_1_3, A1=>nx10078, B0
      =>que_out_16_1_3, B1=>nx10104);
   ix8766 : aoi22 port map ( Y=>nx8765, A0=>que_out_24_1_3, A1=>nx10052, B0
      =>que_out_22_1_3, B1=>nx10026);
   ix5795 : nand03 port map ( Y=>nx5794, A0=>nx8769, A1=>nx8771, A2=>nx8773
   );
   ix8770 : aoi222 port map ( Y=>nx8769, A0=>que_out_15_1_3, A1=>nx9974, B0
      =>que_out_3_1_3, B1=>nx10000, C0=>que_out_23_1_3, C1=>nx9948);
   ix8772 : aoi22 port map ( Y=>nx8771, A0=>que_out_27_1_3, A1=>nx9922, B0=>
      que_out_4_1_3, B1=>nx9896);
   ix8774 : aoi22 port map ( Y=>nx8773, A0=>que_out_0_1_3, A1=>nx9844, B0=>
      que_out_2_1_3, B1=>nx9870);
   ix5769 : nand03 port map ( Y=>nx5768, A0=>nx8777, A1=>nx8779, A2=>nx8781
   );
   ix8778 : aoi222 port map ( Y=>nx8777, A0=>que_out_26_1_3, A1=>nx9818, B0
      =>que_out_14_1_3, B1=>nx9792, C0=>que_out_11_1_3, C1=>nx9766);
   ix8780 : aoi22 port map ( Y=>nx8779, A0=>que_out_13_1_3, A1=>nx9740, B0=>
      que_out_7_1_3, B1=>nx9714);
   ix8782 : aoi22 port map ( Y=>nx8781, A0=>que_out_12_1_3, A1=>nx9688, B0=>
      que_out_1_1_3, B1=>nx9662);
   ix5963 : or04 port map ( Y=>out_column_1_4, A0=>nx5958, A1=>nx5932, A2=>
      nx5904, A3=>nx5878);
   ix5959 : nand03 port map ( Y=>nx5958, A0=>nx8787, A1=>nx8789, A2=>nx8791
   );
   ix8788 : aoi222 port map ( Y=>nx8787, A0=>que_out_10_1_4, A1=>nx10312, B0
      =>que_out_6_1_4, B1=>nx10364, C0=>que_out_9_1_4, C1=>nx10338);
   ix8790 : aoi22 port map ( Y=>nx8789, A0=>que_out_5_1_4, A1=>nx10260, B0=>
      que_out_18_1_4, B1=>nx10286);
   ix8792 : aoi22 port map ( Y=>nx8791, A0=>que_out_17_1_4, A1=>nx10234, B0
      =>que_out_20_1_4, B1=>nx10208);
   ix5933 : nand03 port map ( Y=>nx5932, A0=>nx8795, A1=>nx8797, A2=>nx8799
   );
   ix8796 : aoi222 port map ( Y=>nx8795, A0=>que_out_19_1_4, A1=>nx10182, B0
      =>que_out_21_1_4, B1=>nx10156, C0=>que_out_8_1_4, C1=>nx10130);
   ix8798 : aoi22 port map ( Y=>nx8797, A0=>que_out_25_1_4, A1=>nx10078, B0
      =>que_out_16_1_4, B1=>nx10104);
   ix8800 : aoi22 port map ( Y=>nx8799, A0=>que_out_24_1_4, A1=>nx10052, B0
      =>que_out_22_1_4, B1=>nx10026);
   ix5905 : nand03 port map ( Y=>nx5904, A0=>nx8803, A1=>nx8805, A2=>nx8807
   );
   ix8804 : aoi222 port map ( Y=>nx8803, A0=>que_out_15_1_4, A1=>nx9974, B0
      =>que_out_3_1_4, B1=>nx10000, C0=>que_out_23_1_4, C1=>nx9948);
   ix8806 : aoi22 port map ( Y=>nx8805, A0=>que_out_27_1_4, A1=>nx9922, B0=>
      que_out_4_1_4, B1=>nx9896);
   ix8808 : aoi22 port map ( Y=>nx8807, A0=>que_out_0_1_4, A1=>nx9844, B0=>
      que_out_2_1_4, B1=>nx9870);
   ix5879 : nand03 port map ( Y=>nx5878, A0=>nx8811, A1=>nx8813, A2=>nx8815
   );
   ix8812 : aoi222 port map ( Y=>nx8811, A0=>que_out_26_1_4, A1=>nx9818, B0
      =>que_out_14_1_4, B1=>nx9792, C0=>que_out_11_1_4, C1=>nx9766);
   ix8814 : aoi22 port map ( Y=>nx8813, A0=>que_out_13_1_4, A1=>nx9740, B0=>
      que_out_7_1_4, B1=>nx9714);
   ix8816 : aoi22 port map ( Y=>nx8815, A0=>que_out_12_1_4, A1=>nx9688, B0=>
      que_out_1_1_4, B1=>nx9662);
   ix6073 : or04 port map ( Y=>out_column_1_5, A0=>nx6068, A1=>nx6042, A2=>
      nx6014, A3=>nx5988);
   ix6069 : nand03 port map ( Y=>nx6068, A0=>nx8821, A1=>nx8823, A2=>nx8825
   );
   ix8822 : aoi222 port map ( Y=>nx8821, A0=>que_out_10_1_5, A1=>nx10312, B0
      =>que_out_6_1_5, B1=>nx10364, C0=>que_out_9_1_5, C1=>nx10338);
   ix8824 : aoi22 port map ( Y=>nx8823, A0=>que_out_5_1_5, A1=>nx10260, B0=>
      que_out_18_1_5, B1=>nx10286);
   ix8826 : aoi22 port map ( Y=>nx8825, A0=>que_out_17_1_5, A1=>nx10234, B0
      =>que_out_20_1_5, B1=>nx10208);
   ix6043 : nand03 port map ( Y=>nx6042, A0=>nx8829, A1=>nx8831, A2=>nx8833
   );
   ix8830 : aoi222 port map ( Y=>nx8829, A0=>que_out_19_1_5, A1=>nx10182, B0
      =>que_out_21_1_5, B1=>nx10156, C0=>que_out_8_1_5, C1=>nx10130);
   ix8832 : aoi22 port map ( Y=>nx8831, A0=>que_out_25_1_5, A1=>nx10078, B0
      =>que_out_16_1_5, B1=>nx10104);
   ix8834 : aoi22 port map ( Y=>nx8833, A0=>que_out_24_1_5, A1=>nx10052, B0
      =>que_out_22_1_5, B1=>nx10026);
   ix6015 : nand03 port map ( Y=>nx6014, A0=>nx8837, A1=>nx8839, A2=>nx8841
   );
   ix8838 : aoi222 port map ( Y=>nx8837, A0=>que_out_15_1_5, A1=>nx9974, B0
      =>que_out_3_1_5, B1=>nx10000, C0=>que_out_23_1_5, C1=>nx9948);
   ix8840 : aoi22 port map ( Y=>nx8839, A0=>que_out_27_1_5, A1=>nx9922, B0=>
      que_out_4_1_5, B1=>nx9896);
   ix8842 : aoi22 port map ( Y=>nx8841, A0=>que_out_0_1_5, A1=>nx9844, B0=>
      que_out_2_1_5, B1=>nx9870);
   ix5989 : nand03 port map ( Y=>nx5988, A0=>nx8845, A1=>nx8847, A2=>nx8849
   );
   ix8846 : aoi222 port map ( Y=>nx8845, A0=>que_out_26_1_5, A1=>nx9818, B0
      =>que_out_14_1_5, B1=>nx9792, C0=>que_out_11_1_5, C1=>nx9766);
   ix8848 : aoi22 port map ( Y=>nx8847, A0=>que_out_13_1_5, A1=>nx9740, B0=>
      que_out_7_1_5, B1=>nx9714);
   ix8850 : aoi22 port map ( Y=>nx8849, A0=>que_out_12_1_5, A1=>nx9688, B0=>
      que_out_1_1_5, B1=>nx9662);
   ix6183 : or04 port map ( Y=>out_column_1_6, A0=>nx6178, A1=>nx6152, A2=>
      nx6124, A3=>nx6098);
   ix6179 : nand03 port map ( Y=>nx6178, A0=>nx8855, A1=>nx8857, A2=>nx8859
   );
   ix8856 : aoi222 port map ( Y=>nx8855, A0=>que_out_10_1_6, A1=>nx10312, B0
      =>que_out_6_1_6, B1=>nx10364, C0=>que_out_9_1_6, C1=>nx10338);
   ix8858 : aoi22 port map ( Y=>nx8857, A0=>que_out_5_1_6, A1=>nx10260, B0=>
      que_out_18_1_6, B1=>nx10286);
   ix8860 : aoi22 port map ( Y=>nx8859, A0=>que_out_17_1_6, A1=>nx10234, B0
      =>que_out_20_1_6, B1=>nx10208);
   ix6153 : nand03 port map ( Y=>nx6152, A0=>nx8863, A1=>nx8865, A2=>nx8867
   );
   ix8864 : aoi222 port map ( Y=>nx8863, A0=>que_out_19_1_6, A1=>nx10182, B0
      =>que_out_21_1_6, B1=>nx10156, C0=>que_out_8_1_6, C1=>nx10130);
   ix8866 : aoi22 port map ( Y=>nx8865, A0=>que_out_25_1_6, A1=>nx10078, B0
      =>que_out_16_1_6, B1=>nx10104);
   ix8868 : aoi22 port map ( Y=>nx8867, A0=>que_out_24_1_6, A1=>nx10052, B0
      =>que_out_22_1_6, B1=>nx10026);
   ix6125 : nand03 port map ( Y=>nx6124, A0=>nx8871, A1=>nx8873, A2=>nx8875
   );
   ix8872 : aoi222 port map ( Y=>nx8871, A0=>que_out_15_1_6, A1=>nx9974, B0
      =>que_out_3_1_6, B1=>nx10000, C0=>que_out_23_1_6, C1=>nx9948);
   ix8874 : aoi22 port map ( Y=>nx8873, A0=>que_out_27_1_6, A1=>nx9922, B0=>
      que_out_4_1_6, B1=>nx9896);
   ix8876 : aoi22 port map ( Y=>nx8875, A0=>que_out_0_1_6, A1=>nx9844, B0=>
      que_out_2_1_6, B1=>nx9870);
   ix6099 : nand03 port map ( Y=>nx6098, A0=>nx8879, A1=>nx8881, A2=>nx8883
   );
   ix8880 : aoi222 port map ( Y=>nx8879, A0=>que_out_26_1_6, A1=>nx9818, B0
      =>que_out_14_1_6, B1=>nx9792, C0=>que_out_11_1_6, C1=>nx9766);
   ix8882 : aoi22 port map ( Y=>nx8881, A0=>que_out_13_1_6, A1=>nx9740, B0=>
      que_out_7_1_6, B1=>nx9714);
   ix8884 : aoi22 port map ( Y=>nx8883, A0=>que_out_12_1_6, A1=>nx9688, B0=>
      que_out_1_1_6, B1=>nx9662);
   ix6293 : or04 port map ( Y=>out_column_1_7, A0=>nx6288, A1=>nx6262, A2=>
      nx6234, A3=>nx6208);
   ix6289 : nand03 port map ( Y=>nx6288, A0=>nx8889, A1=>nx8891, A2=>nx8893
   );
   ix8890 : aoi222 port map ( Y=>nx8889, A0=>que_out_10_1_7, A1=>nx10312, B0
      =>que_out_6_1_7, B1=>nx10364, C0=>que_out_9_1_7, C1=>nx10338);
   ix8892 : aoi22 port map ( Y=>nx8891, A0=>que_out_5_1_7, A1=>nx10260, B0=>
      que_out_18_1_7, B1=>nx10286);
   ix8894 : aoi22 port map ( Y=>nx8893, A0=>que_out_17_1_7, A1=>nx10234, B0
      =>que_out_20_1_7, B1=>nx10208);
   ix6263 : nand03 port map ( Y=>nx6262, A0=>nx8897, A1=>nx8899, A2=>nx8901
   );
   ix8898 : aoi222 port map ( Y=>nx8897, A0=>que_out_19_1_7, A1=>nx10182, B0
      =>que_out_21_1_7, B1=>nx10156, C0=>que_out_8_1_7, C1=>nx10130);
   ix8900 : aoi22 port map ( Y=>nx8899, A0=>que_out_25_1_7, A1=>nx10078, B0
      =>que_out_16_1_7, B1=>nx10104);
   ix8902 : aoi22 port map ( Y=>nx8901, A0=>que_out_24_1_7, A1=>nx10052, B0
      =>que_out_22_1_7, B1=>nx10026);
   ix6235 : nand03 port map ( Y=>nx6234, A0=>nx8905, A1=>nx8907, A2=>nx8909
   );
   ix8906 : aoi222 port map ( Y=>nx8905, A0=>que_out_15_1_7, A1=>nx9974, B0
      =>que_out_3_1_7, B1=>nx10000, C0=>que_out_23_1_7, C1=>nx9948);
   ix8908 : aoi22 port map ( Y=>nx8907, A0=>que_out_27_1_7, A1=>nx9922, B0=>
      que_out_4_1_7, B1=>nx9896);
   ix8910 : aoi22 port map ( Y=>nx8909, A0=>que_out_0_1_7, A1=>nx9844, B0=>
      que_out_2_1_7, B1=>nx9870);
   ix6209 : nand03 port map ( Y=>nx6208, A0=>nx8913, A1=>nx8915, A2=>nx8917
   );
   ix8914 : aoi222 port map ( Y=>nx8913, A0=>que_out_26_1_7, A1=>nx9818, B0
      =>que_out_14_1_7, B1=>nx9792, C0=>que_out_11_1_7, C1=>nx9766);
   ix8916 : aoi22 port map ( Y=>nx8915, A0=>que_out_13_1_7, A1=>nx9740, B0=>
      que_out_7_1_7, B1=>nx9714);
   ix8918 : aoi22 port map ( Y=>nx8917, A0=>que_out_12_1_7, A1=>nx9688, B0=>
      que_out_1_1_7, B1=>nx9662);
   ix6403 : or04 port map ( Y=>out_column_1_8, A0=>nx6398, A1=>nx6372, A2=>
      nx6344, A3=>nx6318);
   ix6399 : nand03 port map ( Y=>nx6398, A0=>nx8923, A1=>nx8925, A2=>nx8927
   );
   ix8924 : aoi222 port map ( Y=>nx8923, A0=>que_out_10_1_8, A1=>nx10314, B0
      =>que_out_6_1_8, B1=>nx10366, C0=>que_out_9_1_8, C1=>nx10340);
   ix8926 : aoi22 port map ( Y=>nx8925, A0=>que_out_5_1_8, A1=>nx10262, B0=>
      que_out_18_1_8, B1=>nx10288);
   ix8928 : aoi22 port map ( Y=>nx8927, A0=>que_out_17_1_8, A1=>nx10236, B0
      =>que_out_20_1_8, B1=>nx10210);
   ix6373 : nand03 port map ( Y=>nx6372, A0=>nx8931, A1=>nx8933, A2=>nx8935
   );
   ix8932 : aoi222 port map ( Y=>nx8931, A0=>que_out_19_1_8, A1=>nx10184, B0
      =>que_out_21_1_8, B1=>nx10158, C0=>que_out_8_1_8, C1=>nx10132);
   ix8934 : aoi22 port map ( Y=>nx8933, A0=>que_out_25_1_8, A1=>nx10080, B0
      =>que_out_16_1_8, B1=>nx10106);
   ix8936 : aoi22 port map ( Y=>nx8935, A0=>que_out_24_1_8, A1=>nx10054, B0
      =>que_out_22_1_8, B1=>nx10028);
   ix6345 : nand03 port map ( Y=>nx6344, A0=>nx8939, A1=>nx8941, A2=>nx8943
   );
   ix8940 : aoi222 port map ( Y=>nx8939, A0=>que_out_15_1_8, A1=>nx9976, B0
      =>que_out_3_1_8, B1=>nx10002, C0=>que_out_23_1_8, C1=>nx9950);
   ix8942 : aoi22 port map ( Y=>nx8941, A0=>que_out_27_1_8, A1=>nx9924, B0=>
      que_out_4_1_8, B1=>nx9898);
   ix8944 : aoi22 port map ( Y=>nx8943, A0=>que_out_0_1_8, A1=>nx9846, B0=>
      que_out_2_1_8, B1=>nx9872);
   ix6319 : nand03 port map ( Y=>nx6318, A0=>nx8947, A1=>nx8949, A2=>nx8951
   );
   ix8948 : aoi222 port map ( Y=>nx8947, A0=>que_out_26_1_8, A1=>nx9820, B0
      =>que_out_14_1_8, B1=>nx9794, C0=>que_out_11_1_8, C1=>nx9768);
   ix8950 : aoi22 port map ( Y=>nx8949, A0=>que_out_13_1_8, A1=>nx9742, B0=>
      que_out_7_1_8, B1=>nx9716);
   ix8952 : aoi22 port map ( Y=>nx8951, A0=>que_out_12_1_8, A1=>nx9690, B0=>
      que_out_1_1_8, B1=>nx9664);
   ix6513 : or04 port map ( Y=>out_column_1_9, A0=>nx6508, A1=>nx6482, A2=>
      nx6454, A3=>nx6428);
   ix6509 : nand03 port map ( Y=>nx6508, A0=>nx8955, A1=>nx8957, A2=>nx8959
   );
   ix8956 : aoi222 port map ( Y=>nx8955, A0=>que_out_10_1_9, A1=>nx10314, B0
      =>que_out_6_1_9, B1=>nx10366, C0=>que_out_9_1_9, C1=>nx10340);
   ix8958 : aoi22 port map ( Y=>nx8957, A0=>que_out_5_1_9, A1=>nx10262, B0=>
      que_out_18_1_9, B1=>nx10288);
   ix8960 : aoi22 port map ( Y=>nx8959, A0=>que_out_17_1_9, A1=>nx10236, B0
      =>que_out_20_1_9, B1=>nx10210);
   ix6483 : nand03 port map ( Y=>nx6482, A0=>nx8963, A1=>nx8965, A2=>nx8967
   );
   ix8964 : aoi222 port map ( Y=>nx8963, A0=>que_out_19_1_9, A1=>nx10184, B0
      =>que_out_21_1_9, B1=>nx10158, C0=>que_out_8_1_9, C1=>nx10132);
   ix8966 : aoi22 port map ( Y=>nx8965, A0=>que_out_25_1_9, A1=>nx10080, B0
      =>que_out_16_1_9, B1=>nx10106);
   ix8968 : aoi22 port map ( Y=>nx8967, A0=>que_out_24_1_9, A1=>nx10054, B0
      =>que_out_22_1_9, B1=>nx10028);
   ix6455 : nand03 port map ( Y=>nx6454, A0=>nx8970, A1=>nx8973, A2=>nx8975
   );
   ix8972 : aoi222 port map ( Y=>nx8970, A0=>que_out_15_1_9, A1=>nx9976, B0
      =>que_out_3_1_9, B1=>nx10002, C0=>que_out_23_1_9, C1=>nx9950);
   ix8974 : aoi22 port map ( Y=>nx8973, A0=>que_out_27_1_9, A1=>nx9924, B0=>
      que_out_4_1_9, B1=>nx9898);
   ix8976 : aoi22 port map ( Y=>nx8975, A0=>que_out_0_1_9, A1=>nx9846, B0=>
      que_out_2_1_9, B1=>nx9872);
   ix6429 : nand03 port map ( Y=>nx6428, A0=>nx8978, A1=>nx8981, A2=>nx8983
   );
   ix8980 : aoi222 port map ( Y=>nx8978, A0=>que_out_26_1_9, A1=>nx9820, B0
      =>que_out_14_1_9, B1=>nx9794, C0=>que_out_11_1_9, C1=>nx9768);
   ix8982 : aoi22 port map ( Y=>nx8981, A0=>que_out_13_1_9, A1=>nx9742, B0=>
      que_out_7_1_9, B1=>nx9716);
   ix8984 : aoi22 port map ( Y=>nx8983, A0=>que_out_12_1_9, A1=>nx9690, B0=>
      que_out_1_1_9, B1=>nx9664);
   ix6623 : or04 port map ( Y=>out_column_1_10, A0=>nx6618, A1=>nx6592, A2=>
      nx6564, A3=>nx6538);
   ix6619 : nand03 port map ( Y=>nx6618, A0=>nx8989, A1=>nx8991, A2=>nx8993
   );
   ix8990 : aoi222 port map ( Y=>nx8989, A0=>que_out_10_1_10, A1=>nx10314, 
      B0=>que_out_6_1_10, B1=>nx10366, C0=>que_out_9_1_10, C1=>nx10340);
   ix8992 : aoi22 port map ( Y=>nx8991, A0=>que_out_5_1_10, A1=>nx10262, B0
      =>que_out_18_1_10, B1=>nx10288);
   ix8994 : aoi22 port map ( Y=>nx8993, A0=>que_out_17_1_10, A1=>nx10236, B0
      =>que_out_20_1_10, B1=>nx10210);
   ix6593 : nand03 port map ( Y=>nx6592, A0=>nx8997, A1=>nx8999, A2=>nx9001
   );
   ix8998 : aoi222 port map ( Y=>nx8997, A0=>que_out_19_1_10, A1=>nx10184, 
      B0=>que_out_21_1_10, B1=>nx10158, C0=>que_out_8_1_10, C1=>nx10132);
   ix9000 : aoi22 port map ( Y=>nx8999, A0=>que_out_25_1_10, A1=>nx10080, B0
      =>que_out_16_1_10, B1=>nx10106);
   ix9002 : aoi22 port map ( Y=>nx9001, A0=>que_out_24_1_10, A1=>nx10054, B0
      =>que_out_22_1_10, B1=>nx10028);
   ix6565 : nand03 port map ( Y=>nx6564, A0=>nx9005, A1=>nx9007, A2=>nx9009
   );
   ix9006 : aoi222 port map ( Y=>nx9005, A0=>que_out_15_1_10, A1=>nx9976, B0
      =>que_out_3_1_10, B1=>nx10002, C0=>que_out_23_1_10, C1=>nx9950);
   ix9008 : aoi22 port map ( Y=>nx9007, A0=>que_out_27_1_10, A1=>nx9924, B0
      =>que_out_4_1_10, B1=>nx9898);
   ix9010 : aoi22 port map ( Y=>nx9009, A0=>que_out_0_1_10, A1=>nx9846, B0=>
      que_out_2_1_10, B1=>nx9872);
   ix6539 : nand03 port map ( Y=>nx6538, A0=>nx9013, A1=>nx9015, A2=>nx9017
   );
   ix9014 : aoi222 port map ( Y=>nx9013, A0=>que_out_26_1_10, A1=>nx9820, B0
      =>que_out_14_1_10, B1=>nx9794, C0=>que_out_11_1_10, C1=>nx9768);
   ix9016 : aoi22 port map ( Y=>nx9015, A0=>que_out_13_1_10, A1=>nx9742, B0
      =>que_out_7_1_10, B1=>nx9716);
   ix9018 : aoi22 port map ( Y=>nx9017, A0=>que_out_12_1_10, A1=>nx9690, B0
      =>que_out_1_1_10, B1=>nx9664);
   ix6733 : or04 port map ( Y=>out_column_1_11, A0=>nx6728, A1=>nx6702, A2=>
      nx6674, A3=>nx6648);
   ix6729 : nand03 port map ( Y=>nx6728, A0=>nx9023, A1=>nx9025, A2=>nx9027
   );
   ix9024 : aoi222 port map ( Y=>nx9023, A0=>que_out_10_1_11, A1=>nx10314, 
      B0=>que_out_6_1_11, B1=>nx10366, C0=>que_out_9_1_11, C1=>nx10340);
   ix9026 : aoi22 port map ( Y=>nx9025, A0=>que_out_5_1_11, A1=>nx10262, B0
      =>que_out_18_1_11, B1=>nx10288);
   ix9028 : aoi22 port map ( Y=>nx9027, A0=>que_out_17_1_11, A1=>nx10236, B0
      =>que_out_20_1_11, B1=>nx10210);
   ix6703 : nand03 port map ( Y=>nx6702, A0=>nx9031, A1=>nx9033, A2=>nx9035
   );
   ix9032 : aoi222 port map ( Y=>nx9031, A0=>que_out_19_1_11, A1=>nx10184, 
      B0=>que_out_21_1_11, B1=>nx10158, C0=>que_out_8_1_11, C1=>nx10132);
   ix9034 : aoi22 port map ( Y=>nx9033, A0=>que_out_25_1_11, A1=>nx10080, B0
      =>que_out_16_1_11, B1=>nx10106);
   ix9036 : aoi22 port map ( Y=>nx9035, A0=>que_out_24_1_11, A1=>nx10054, B0
      =>que_out_22_1_11, B1=>nx10028);
   ix6675 : nand03 port map ( Y=>nx6674, A0=>nx9039, A1=>nx9041, A2=>nx9043
   );
   ix9040 : aoi222 port map ( Y=>nx9039, A0=>que_out_15_1_11, A1=>nx9976, B0
      =>que_out_3_1_11, B1=>nx10002, C0=>que_out_23_1_11, C1=>nx9950);
   ix9042 : aoi22 port map ( Y=>nx9041, A0=>que_out_27_1_11, A1=>nx9924, B0
      =>que_out_4_1_11, B1=>nx9898);
   ix9044 : aoi22 port map ( Y=>nx9043, A0=>que_out_0_1_11, A1=>nx9846, B0=>
      que_out_2_1_11, B1=>nx9872);
   ix6649 : nand03 port map ( Y=>nx6648, A0=>nx9047, A1=>nx9049, A2=>nx9051
   );
   ix9048 : aoi222 port map ( Y=>nx9047, A0=>que_out_26_1_11, A1=>nx9820, B0
      =>que_out_14_1_11, B1=>nx9794, C0=>que_out_11_1_11, C1=>nx9768);
   ix9050 : aoi22 port map ( Y=>nx9049, A0=>que_out_13_1_11, A1=>nx9742, B0
      =>que_out_7_1_11, B1=>nx9716);
   ix9052 : aoi22 port map ( Y=>nx9051, A0=>que_out_12_1_11, A1=>nx9690, B0
      =>que_out_1_1_11, B1=>nx9664);
   ix6843 : or04 port map ( Y=>out_column_1_12, A0=>nx6838, A1=>nx6812, A2=>
      nx6784, A3=>nx6758);
   ix6839 : nand03 port map ( Y=>nx6838, A0=>nx9057, A1=>nx9059, A2=>nx9061
   );
   ix9058 : aoi222 port map ( Y=>nx9057, A0=>que_out_10_1_12, A1=>nx10314, 
      B0=>que_out_6_1_12, B1=>nx10366, C0=>que_out_9_1_12, C1=>nx10340);
   ix9060 : aoi22 port map ( Y=>nx9059, A0=>que_out_5_1_12, A1=>nx10262, B0
      =>que_out_18_1_12, B1=>nx10288);
   ix9062 : aoi22 port map ( Y=>nx9061, A0=>que_out_17_1_12, A1=>nx10236, B0
      =>que_out_20_1_12, B1=>nx10210);
   ix6813 : nand03 port map ( Y=>nx6812, A0=>nx9065, A1=>nx9067, A2=>nx9069
   );
   ix9066 : aoi222 port map ( Y=>nx9065, A0=>que_out_19_1_12, A1=>nx10184, 
      B0=>que_out_21_1_12, B1=>nx10158, C0=>que_out_8_1_12, C1=>nx10132);
   ix9068 : aoi22 port map ( Y=>nx9067, A0=>que_out_25_1_12, A1=>nx10080, B0
      =>que_out_16_1_12, B1=>nx10106);
   ix9070 : aoi22 port map ( Y=>nx9069, A0=>que_out_24_1_12, A1=>nx10054, B0
      =>que_out_22_1_12, B1=>nx10028);
   ix6785 : nand03 port map ( Y=>nx6784, A0=>nx9073, A1=>nx9075, A2=>nx9077
   );
   ix9074 : aoi222 port map ( Y=>nx9073, A0=>que_out_15_1_12, A1=>nx9976, B0
      =>que_out_3_1_12, B1=>nx10002, C0=>que_out_23_1_12, C1=>nx9950);
   ix9076 : aoi22 port map ( Y=>nx9075, A0=>que_out_27_1_12, A1=>nx9924, B0
      =>que_out_4_1_12, B1=>nx9898);
   ix9078 : aoi22 port map ( Y=>nx9077, A0=>que_out_0_1_12, A1=>nx9846, B0=>
      que_out_2_1_12, B1=>nx9872);
   ix6759 : nand03 port map ( Y=>nx6758, A0=>nx9081, A1=>nx9083, A2=>nx9085
   );
   ix9082 : aoi222 port map ( Y=>nx9081, A0=>que_out_26_1_12, A1=>nx9820, B0
      =>que_out_14_1_12, B1=>nx9794, C0=>que_out_11_1_12, C1=>nx9768);
   ix9084 : aoi22 port map ( Y=>nx9083, A0=>que_out_13_1_12, A1=>nx9742, B0
      =>que_out_7_1_12, B1=>nx9716);
   ix9086 : aoi22 port map ( Y=>nx9085, A0=>que_out_12_1_12, A1=>nx9690, B0
      =>que_out_1_1_12, B1=>nx9664);
   ix6953 : or04 port map ( Y=>out_column_1_13, A0=>nx6948, A1=>nx6922, A2=>
      nx6894, A3=>nx6868);
   ix6949 : nand03 port map ( Y=>nx6948, A0=>nx9090, A1=>nx9093, A2=>nx9095
   );
   ix9092 : aoi222 port map ( Y=>nx9090, A0=>que_out_10_1_13, A1=>nx10314, 
      B0=>que_out_6_1_13, B1=>nx10366, C0=>que_out_9_1_13, C1=>nx10340);
   ix9094 : aoi22 port map ( Y=>nx9093, A0=>que_out_5_1_13, A1=>nx10262, B0
      =>que_out_18_1_13, B1=>nx10288);
   ix9096 : aoi22 port map ( Y=>nx9095, A0=>que_out_17_1_13, A1=>nx10236, B0
      =>que_out_20_1_13, B1=>nx10210);
   ix6923 : nand03 port map ( Y=>nx6922, A0=>nx9098, A1=>nx9101, A2=>nx9103
   );
   ix9100 : aoi222 port map ( Y=>nx9098, A0=>que_out_19_1_13, A1=>nx10184, 
      B0=>que_out_21_1_13, B1=>nx10158, C0=>que_out_8_1_13, C1=>nx10132);
   ix9102 : aoi22 port map ( Y=>nx9101, A0=>que_out_25_1_13, A1=>nx10080, B0
      =>que_out_16_1_13, B1=>nx10106);
   ix9104 : aoi22 port map ( Y=>nx9103, A0=>que_out_24_1_13, A1=>nx10054, B0
      =>que_out_22_1_13, B1=>nx10028);
   ix6895 : nand03 port map ( Y=>nx6894, A0=>nx9106, A1=>nx9108, A2=>nx9110
   );
   ix9107 : aoi222 port map ( Y=>nx9106, A0=>que_out_15_1_13, A1=>nx9976, B0
      =>que_out_3_1_13, B1=>nx10002, C0=>que_out_23_1_13, C1=>nx9950);
   ix9109 : aoi22 port map ( Y=>nx9108, A0=>que_out_27_1_13, A1=>nx9924, B0
      =>que_out_4_1_13, B1=>nx9898);
   ix9111 : aoi22 port map ( Y=>nx9110, A0=>que_out_0_1_13, A1=>nx9846, B0=>
      que_out_2_1_13, B1=>nx9872);
   ix6869 : nand03 port map ( Y=>nx6868, A0=>nx9113, A1=>nx9115, A2=>nx9117
   );
   ix9114 : aoi222 port map ( Y=>nx9113, A0=>que_out_26_1_13, A1=>nx9820, B0
      =>que_out_14_1_13, B1=>nx9794, C0=>que_out_11_1_13, C1=>nx9768);
   ix9116 : aoi22 port map ( Y=>nx9115, A0=>que_out_13_1_13, A1=>nx9742, B0
      =>que_out_7_1_13, B1=>nx9716);
   ix9118 : aoi22 port map ( Y=>nx9117, A0=>que_out_12_1_13, A1=>nx9690, B0
      =>que_out_1_1_13, B1=>nx9664);
   ix7063 : or04 port map ( Y=>out_column_1_14, A0=>nx7058, A1=>nx7032, A2=>
      nx7004, A3=>nx6978);
   ix7059 : nand03 port map ( Y=>nx7058, A0=>nx9121, A1=>nx9123, A2=>nx9125
   );
   ix9122 : aoi222 port map ( Y=>nx9121, A0=>que_out_10_1_14, A1=>nx10314, 
      B0=>que_out_6_1_14, B1=>nx10366, C0=>que_out_9_1_14, C1=>nx10340);
   ix9124 : aoi22 port map ( Y=>nx9123, A0=>que_out_5_1_14, A1=>nx10262, B0
      =>que_out_18_1_14, B1=>nx10288);
   ix9126 : aoi22 port map ( Y=>nx9125, A0=>que_out_17_1_14, A1=>nx10236, B0
      =>que_out_20_1_14, B1=>nx10210);
   ix7033 : nand03 port map ( Y=>nx7032, A0=>nx9128, A1=>nx9130, A2=>nx9132
   );
   ix9129 : aoi222 port map ( Y=>nx9128, A0=>que_out_19_1_14, A1=>nx10184, 
      B0=>que_out_21_1_14, B1=>nx10158, C0=>que_out_8_1_14, C1=>nx10132);
   ix9131 : aoi22 port map ( Y=>nx9130, A0=>que_out_25_1_14, A1=>nx10080, B0
      =>que_out_16_1_14, B1=>nx10106);
   ix9133 : aoi22 port map ( Y=>nx9132, A0=>que_out_24_1_14, A1=>nx10054, B0
      =>que_out_22_1_14, B1=>nx10028);
   ix7005 : nand03 port map ( Y=>nx7004, A0=>nx9135, A1=>nx9137, A2=>nx9139
   );
   ix9136 : aoi222 port map ( Y=>nx9135, A0=>que_out_15_1_14, A1=>nx9976, B0
      =>que_out_3_1_14, B1=>nx10002, C0=>que_out_23_1_14, C1=>nx9950);
   ix9138 : aoi22 port map ( Y=>nx9137, A0=>que_out_27_1_14, A1=>nx9924, B0
      =>que_out_4_1_14, B1=>nx9898);
   ix9140 : aoi22 port map ( Y=>nx9139, A0=>que_out_0_1_14, A1=>nx9846, B0=>
      que_out_2_1_14, B1=>nx9872);
   ix6979 : nand03 port map ( Y=>nx6978, A0=>nx9142, A1=>nx9144, A2=>nx9146
   );
   ix9143 : aoi222 port map ( Y=>nx9142, A0=>que_out_26_1_14, A1=>nx9820, B0
      =>que_out_14_1_14, B1=>nx9794, C0=>que_out_11_1_14, C1=>nx9768);
   ix9145 : aoi22 port map ( Y=>nx9144, A0=>que_out_13_1_14, A1=>nx9742, B0
      =>que_out_7_1_14, B1=>nx9716);
   ix9147 : aoi22 port map ( Y=>nx9146, A0=>que_out_12_1_14, A1=>nx9690, B0
      =>que_out_1_1_14, B1=>nx9664);
   ix7173 : or04 port map ( Y=>out_column_1_15, A0=>nx7168, A1=>nx7142, A2=>
      nx7114, A3=>nx7088);
   ix7169 : nand03 port map ( Y=>nx7168, A0=>nx9150, A1=>nx9152, A2=>nx9154
   );
   ix9151 : aoi222 port map ( Y=>nx9150, A0=>que_out_10_1_15, A1=>nx10316, 
      B0=>que_out_6_1_15, B1=>nx10368, C0=>que_out_9_1_15, C1=>nx10342);
   ix9153 : aoi22 port map ( Y=>nx9152, A0=>que_out_5_1_15, A1=>nx10264, B0
      =>que_out_18_1_15, B1=>nx10290);
   ix9155 : aoi22 port map ( Y=>nx9154, A0=>que_out_17_1_15, A1=>nx10238, B0
      =>que_out_20_1_15, B1=>nx10212);
   ix7143 : nand03 port map ( Y=>nx7142, A0=>nx9157, A1=>nx9159, A2=>nx9161
   );
   ix9158 : aoi222 port map ( Y=>nx9157, A0=>que_out_19_1_15, A1=>nx10186, 
      B0=>que_out_21_1_15, B1=>nx10160, C0=>que_out_8_1_15, C1=>nx10134);
   ix9160 : aoi22 port map ( Y=>nx9159, A0=>que_out_25_1_15, A1=>nx10082, B0
      =>que_out_16_1_15, B1=>nx10108);
   ix9162 : aoi22 port map ( Y=>nx9161, A0=>que_out_24_1_15, A1=>nx10056, B0
      =>que_out_22_1_15, B1=>nx10030);
   ix7115 : nand03 port map ( Y=>nx7114, A0=>nx9164, A1=>nx9166, A2=>nx9168
   );
   ix9165 : aoi222 port map ( Y=>nx9164, A0=>que_out_15_1_15, A1=>nx9978, B0
      =>que_out_3_1_15, B1=>nx10004, C0=>que_out_23_1_15, C1=>nx9952);
   ix9167 : aoi22 port map ( Y=>nx9166, A0=>que_out_27_1_15, A1=>nx9926, B0
      =>que_out_4_1_15, B1=>nx9900);
   ix9169 : aoi22 port map ( Y=>nx9168, A0=>que_out_0_1_15, A1=>nx9848, B0=>
      que_out_2_1_15, B1=>nx9874);
   ix7089 : nand03 port map ( Y=>nx7088, A0=>nx9171, A1=>nx9173, A2=>nx9175
   );
   ix9172 : aoi222 port map ( Y=>nx9171, A0=>que_out_26_1_15, A1=>nx9822, B0
      =>que_out_14_1_15, B1=>nx9796, C0=>que_out_11_1_15, C1=>nx9770);
   ix9174 : aoi22 port map ( Y=>nx9173, A0=>que_out_13_1_15, A1=>nx9744, B0
      =>que_out_7_1_15, B1=>nx9718);
   ix9176 : aoi22 port map ( Y=>nx9175, A0=>que_out_12_1_15, A1=>nx9692, B0
      =>que_out_1_1_15, B1=>nx9666);
   ix7283 : or04 port map ( Y=>out_column_0_0, A0=>nx7278, A1=>nx7252, A2=>
      nx7224, A3=>nx7198);
   ix7279 : nand03 port map ( Y=>nx7278, A0=>nx9179, A1=>nx9181, A2=>nx9183
   );
   ix9180 : aoi222 port map ( Y=>nx9179, A0=>que_out_10_0_0, A1=>nx10316, B0
      =>que_out_6_0_0, B1=>nx10368, C0=>que_out_9_0_0, C1=>nx10342);
   ix9182 : aoi22 port map ( Y=>nx9181, A0=>que_out_5_0_0, A1=>nx10264, B0=>
      que_out_18_0_0, B1=>nx10290);
   ix9184 : aoi22 port map ( Y=>nx9183, A0=>que_out_17_0_0, A1=>nx10238, B0
      =>que_out_20_0_0, B1=>nx10212);
   ix7253 : nand03 port map ( Y=>nx7252, A0=>nx9186, A1=>nx9188, A2=>nx9190
   );
   ix9187 : aoi222 port map ( Y=>nx9186, A0=>que_out_19_0_0, A1=>nx10186, B0
      =>que_out_21_0_0, B1=>nx10160, C0=>que_out_8_0_0, C1=>nx10134);
   ix9189 : aoi22 port map ( Y=>nx9188, A0=>que_out_25_0_0, A1=>nx10082, B0
      =>que_out_16_0_0, B1=>nx10108);
   ix9191 : aoi22 port map ( Y=>nx9190, A0=>que_out_24_0_0, A1=>nx10056, B0
      =>que_out_22_0_0, B1=>nx10030);
   ix7225 : nand03 port map ( Y=>nx7224, A0=>nx9193, A1=>nx9195, A2=>nx9197
   );
   ix9194 : aoi222 port map ( Y=>nx9193, A0=>que_out_15_0_0, A1=>nx9978, B0
      =>que_out_3_0_0, B1=>nx10004, C0=>que_out_23_0_0, C1=>nx9952);
   ix9196 : aoi22 port map ( Y=>nx9195, A0=>que_out_27_0_0, A1=>nx9926, B0=>
      que_out_4_0_0, B1=>nx9900);
   ix9198 : aoi22 port map ( Y=>nx9197, A0=>que_out_0_0_0, A1=>nx9848, B0=>
      que_out_2_0_0, B1=>nx9874);
   ix7199 : nand03 port map ( Y=>nx7198, A0=>nx9200, A1=>nx9202, A2=>nx9204
   );
   ix9201 : aoi222 port map ( Y=>nx9200, A0=>que_out_26_0_0, A1=>nx9822, B0
      =>que_out_14_0_0, B1=>nx9796, C0=>que_out_11_0_0, C1=>nx9770);
   ix9203 : aoi22 port map ( Y=>nx9202, A0=>que_out_13_0_0, A1=>nx9744, B0=>
      que_out_7_0_0, B1=>nx9718);
   ix9205 : aoi22 port map ( Y=>nx9204, A0=>que_out_12_0_0, A1=>nx9692, B0=>
      que_out_1_0_0, B1=>nx9666);
   ix7393 : or04 port map ( Y=>out_column_0_1, A0=>nx7388, A1=>nx7362, A2=>
      nx7334, A3=>nx7308);
   ix7389 : nand03 port map ( Y=>nx7388, A0=>nx9208, A1=>nx9210, A2=>nx9212
   );
   ix9209 : aoi222 port map ( Y=>nx9208, A0=>que_out_10_0_1, A1=>nx10316, B0
      =>que_out_6_0_1, B1=>nx10368, C0=>que_out_9_0_1, C1=>nx10342);
   ix9211 : aoi22 port map ( Y=>nx9210, A0=>que_out_5_0_1, A1=>nx10264, B0=>
      que_out_18_0_1, B1=>nx10290);
   ix9213 : aoi22 port map ( Y=>nx9212, A0=>que_out_17_0_1, A1=>nx10238, B0
      =>que_out_20_0_1, B1=>nx10212);
   ix7363 : nand03 port map ( Y=>nx7362, A0=>nx9215, A1=>nx9217, A2=>nx9219
   );
   ix9216 : aoi222 port map ( Y=>nx9215, A0=>que_out_19_0_1, A1=>nx10186, B0
      =>que_out_21_0_1, B1=>nx10160, C0=>que_out_8_0_1, C1=>nx10134);
   ix9218 : aoi22 port map ( Y=>nx9217, A0=>que_out_25_0_1, A1=>nx10082, B0
      =>que_out_16_0_1, B1=>nx10108);
   ix9220 : aoi22 port map ( Y=>nx9219, A0=>que_out_24_0_1, A1=>nx10056, B0
      =>que_out_22_0_1, B1=>nx10030);
   ix7335 : nand03 port map ( Y=>nx7334, A0=>nx9222, A1=>nx9224, A2=>nx9226
   );
   ix9223 : aoi222 port map ( Y=>nx9222, A0=>que_out_15_0_1, A1=>nx9978, B0
      =>que_out_3_0_1, B1=>nx10004, C0=>que_out_23_0_1, C1=>nx9952);
   ix9225 : aoi22 port map ( Y=>nx9224, A0=>que_out_27_0_1, A1=>nx9926, B0=>
      que_out_4_0_1, B1=>nx9900);
   ix9227 : aoi22 port map ( Y=>nx9226, A0=>que_out_0_0_1, A1=>nx9848, B0=>
      que_out_2_0_1, B1=>nx9874);
   ix7309 : nand03 port map ( Y=>nx7308, A0=>nx9229, A1=>nx9231, A2=>nx9233
   );
   ix9230 : aoi222 port map ( Y=>nx9229, A0=>que_out_26_0_1, A1=>nx9822, B0
      =>que_out_14_0_1, B1=>nx9796, C0=>que_out_11_0_1, C1=>nx9770);
   ix9232 : aoi22 port map ( Y=>nx9231, A0=>que_out_13_0_1, A1=>nx9744, B0=>
      que_out_7_0_1, B1=>nx9718);
   ix9234 : aoi22 port map ( Y=>nx9233, A0=>que_out_12_0_1, A1=>nx9692, B0=>
      que_out_1_0_1, B1=>nx9666);
   ix7503 : or04 port map ( Y=>out_column_0_2, A0=>nx7498, A1=>nx7472, A2=>
      nx7444, A3=>nx7418);
   ix7499 : nand03 port map ( Y=>nx7498, A0=>nx9237, A1=>nx9239, A2=>nx9241
   );
   ix9238 : aoi222 port map ( Y=>nx9237, A0=>que_out_10_0_2, A1=>nx10316, B0
      =>que_out_6_0_2, B1=>nx10368, C0=>que_out_9_0_2, C1=>nx10342);
   ix9240 : aoi22 port map ( Y=>nx9239, A0=>que_out_5_0_2, A1=>nx10264, B0=>
      que_out_18_0_2, B1=>nx10290);
   ix9242 : aoi22 port map ( Y=>nx9241, A0=>que_out_17_0_2, A1=>nx10238, B0
      =>que_out_20_0_2, B1=>nx10212);
   ix7473 : nand03 port map ( Y=>nx7472, A0=>nx9244, A1=>nx9246, A2=>nx9248
   );
   ix9245 : aoi222 port map ( Y=>nx9244, A0=>que_out_19_0_2, A1=>nx10186, B0
      =>que_out_21_0_2, B1=>nx10160, C0=>que_out_8_0_2, C1=>nx10134);
   ix9247 : aoi22 port map ( Y=>nx9246, A0=>que_out_25_0_2, A1=>nx10082, B0
      =>que_out_16_0_2, B1=>nx10108);
   ix9249 : aoi22 port map ( Y=>nx9248, A0=>que_out_24_0_2, A1=>nx10056, B0
      =>que_out_22_0_2, B1=>nx10030);
   ix7445 : nand03 port map ( Y=>nx7444, A0=>nx9251, A1=>nx9253, A2=>nx9255
   );
   ix9252 : aoi222 port map ( Y=>nx9251, A0=>que_out_15_0_2, A1=>nx9978, B0
      =>que_out_3_0_2, B1=>nx10004, C0=>que_out_23_0_2, C1=>nx9952);
   ix9254 : aoi22 port map ( Y=>nx9253, A0=>que_out_27_0_2, A1=>nx9926, B0=>
      que_out_4_0_2, B1=>nx9900);
   ix9256 : aoi22 port map ( Y=>nx9255, A0=>que_out_0_0_2, A1=>nx9848, B0=>
      que_out_2_0_2, B1=>nx9874);
   ix7419 : nand03 port map ( Y=>nx7418, A0=>nx9258, A1=>nx9260, A2=>nx9262
   );
   ix9259 : aoi222 port map ( Y=>nx9258, A0=>que_out_26_0_2, A1=>nx9822, B0
      =>que_out_14_0_2, B1=>nx9796, C0=>que_out_11_0_2, C1=>nx9770);
   ix9261 : aoi22 port map ( Y=>nx9260, A0=>que_out_13_0_2, A1=>nx9744, B0=>
      que_out_7_0_2, B1=>nx9718);
   ix9263 : aoi22 port map ( Y=>nx9262, A0=>que_out_12_0_2, A1=>nx9692, B0=>
      que_out_1_0_2, B1=>nx9666);
   ix7613 : or04 port map ( Y=>out_column_0_3, A0=>nx7608, A1=>nx7582, A2=>
      nx7554, A3=>nx7528);
   ix7609 : nand03 port map ( Y=>nx7608, A0=>nx9266, A1=>nx9268, A2=>nx9270
   );
   ix9267 : aoi222 port map ( Y=>nx9266, A0=>que_out_10_0_3, A1=>nx10316, B0
      =>que_out_6_0_3, B1=>nx10368, C0=>que_out_9_0_3, C1=>nx10342);
   ix9269 : aoi22 port map ( Y=>nx9268, A0=>que_out_5_0_3, A1=>nx10264, B0=>
      que_out_18_0_3, B1=>nx10290);
   ix9271 : aoi22 port map ( Y=>nx9270, A0=>que_out_17_0_3, A1=>nx10238, B0
      =>que_out_20_0_3, B1=>nx10212);
   ix7583 : nand03 port map ( Y=>nx7582, A0=>nx9273, A1=>nx9275, A2=>nx9277
   );
   ix9274 : aoi222 port map ( Y=>nx9273, A0=>que_out_19_0_3, A1=>nx10186, B0
      =>que_out_21_0_3, B1=>nx10160, C0=>que_out_8_0_3, C1=>nx10134);
   ix9276 : aoi22 port map ( Y=>nx9275, A0=>que_out_25_0_3, A1=>nx10082, B0
      =>que_out_16_0_3, B1=>nx10108);
   ix9278 : aoi22 port map ( Y=>nx9277, A0=>que_out_24_0_3, A1=>nx10056, B0
      =>que_out_22_0_3, B1=>nx10030);
   ix7555 : nand03 port map ( Y=>nx7554, A0=>nx9280, A1=>nx9282, A2=>nx9284
   );
   ix9281 : aoi222 port map ( Y=>nx9280, A0=>que_out_15_0_3, A1=>nx9978, B0
      =>que_out_3_0_3, B1=>nx10004, C0=>que_out_23_0_3, C1=>nx9952);
   ix9283 : aoi22 port map ( Y=>nx9282, A0=>que_out_27_0_3, A1=>nx9926, B0=>
      que_out_4_0_3, B1=>nx9900);
   ix9285 : aoi22 port map ( Y=>nx9284, A0=>que_out_0_0_3, A1=>nx9848, B0=>
      que_out_2_0_3, B1=>nx9874);
   ix7529 : nand03 port map ( Y=>nx7528, A0=>nx9287, A1=>nx9289, A2=>nx9291
   );
   ix9288 : aoi222 port map ( Y=>nx9287, A0=>que_out_26_0_3, A1=>nx9822, B0
      =>que_out_14_0_3, B1=>nx9796, C0=>que_out_11_0_3, C1=>nx9770);
   ix9290 : aoi22 port map ( Y=>nx9289, A0=>que_out_13_0_3, A1=>nx9744, B0=>
      que_out_7_0_3, B1=>nx9718);
   ix9292 : aoi22 port map ( Y=>nx9291, A0=>que_out_12_0_3, A1=>nx9692, B0=>
      que_out_1_0_3, B1=>nx9666);
   ix7723 : or04 port map ( Y=>out_column_0_4, A0=>nx7718, A1=>nx7692, A2=>
      nx7664, A3=>nx7638);
   ix7719 : nand03 port map ( Y=>nx7718, A0=>nx9295, A1=>nx9297, A2=>nx9299
   );
   ix9296 : aoi222 port map ( Y=>nx9295, A0=>que_out_10_0_4, A1=>nx10316, B0
      =>que_out_6_0_4, B1=>nx10368, C0=>que_out_9_0_4, C1=>nx10342);
   ix9298 : aoi22 port map ( Y=>nx9297, A0=>que_out_5_0_4, A1=>nx10264, B0=>
      que_out_18_0_4, B1=>nx10290);
   ix9300 : aoi22 port map ( Y=>nx9299, A0=>que_out_17_0_4, A1=>nx10238, B0
      =>que_out_20_0_4, B1=>nx10212);
   ix7693 : nand03 port map ( Y=>nx7692, A0=>nx9302, A1=>nx9304, A2=>nx9306
   );
   ix9303 : aoi222 port map ( Y=>nx9302, A0=>que_out_19_0_4, A1=>nx10186, B0
      =>que_out_21_0_4, B1=>nx10160, C0=>que_out_8_0_4, C1=>nx10134);
   ix9305 : aoi22 port map ( Y=>nx9304, A0=>que_out_25_0_4, A1=>nx10082, B0
      =>que_out_16_0_4, B1=>nx10108);
   ix9307 : aoi22 port map ( Y=>nx9306, A0=>que_out_24_0_4, A1=>nx10056, B0
      =>que_out_22_0_4, B1=>nx10030);
   ix7665 : nand03 port map ( Y=>nx7664, A0=>nx9309, A1=>nx9311, A2=>nx9313
   );
   ix9310 : aoi222 port map ( Y=>nx9309, A0=>que_out_15_0_4, A1=>nx9978, B0
      =>que_out_3_0_4, B1=>nx10004, C0=>que_out_23_0_4, C1=>nx9952);
   ix9312 : aoi22 port map ( Y=>nx9311, A0=>que_out_27_0_4, A1=>nx9926, B0=>
      que_out_4_0_4, B1=>nx9900);
   ix9314 : aoi22 port map ( Y=>nx9313, A0=>que_out_0_0_4, A1=>nx9848, B0=>
      que_out_2_0_4, B1=>nx9874);
   ix7639 : nand03 port map ( Y=>nx7638, A0=>nx9316, A1=>nx9318, A2=>nx9320
   );
   ix9317 : aoi222 port map ( Y=>nx9316, A0=>que_out_26_0_4, A1=>nx9822, B0
      =>que_out_14_0_4, B1=>nx9796, C0=>que_out_11_0_4, C1=>nx9770);
   ix9319 : aoi22 port map ( Y=>nx9318, A0=>que_out_13_0_4, A1=>nx9744, B0=>
      que_out_7_0_4, B1=>nx9718);
   ix9321 : aoi22 port map ( Y=>nx9320, A0=>que_out_12_0_4, A1=>nx9692, B0=>
      que_out_1_0_4, B1=>nx9666);
   ix7833 : or04 port map ( Y=>out_column_0_5, A0=>nx7828, A1=>nx7802, A2=>
      nx7774, A3=>nx7748);
   ix7829 : nand03 port map ( Y=>nx7828, A0=>nx9324, A1=>nx9326, A2=>nx9328
   );
   ix9325 : aoi222 port map ( Y=>nx9324, A0=>que_out_10_0_5, A1=>nx10316, B0
      =>que_out_6_0_5, B1=>nx10368, C0=>que_out_9_0_5, C1=>nx10342);
   ix9327 : aoi22 port map ( Y=>nx9326, A0=>que_out_5_0_5, A1=>nx10264, B0=>
      que_out_18_0_5, B1=>nx10290);
   ix9329 : aoi22 port map ( Y=>nx9328, A0=>que_out_17_0_5, A1=>nx10238, B0
      =>que_out_20_0_5, B1=>nx10212);
   ix7803 : nand03 port map ( Y=>nx7802, A0=>nx9331, A1=>nx9333, A2=>nx9335
   );
   ix9332 : aoi222 port map ( Y=>nx9331, A0=>que_out_19_0_5, A1=>nx10186, B0
      =>que_out_21_0_5, B1=>nx10160, C0=>que_out_8_0_5, C1=>nx10134);
   ix9334 : aoi22 port map ( Y=>nx9333, A0=>que_out_25_0_5, A1=>nx10082, B0
      =>que_out_16_0_5, B1=>nx10108);
   ix9336 : aoi22 port map ( Y=>nx9335, A0=>que_out_24_0_5, A1=>nx10056, B0
      =>que_out_22_0_5, B1=>nx10030);
   ix7775 : nand03 port map ( Y=>nx7774, A0=>nx9338, A1=>nx9340, A2=>nx9342
   );
   ix9339 : aoi222 port map ( Y=>nx9338, A0=>que_out_15_0_5, A1=>nx9978, B0
      =>que_out_3_0_5, B1=>nx10004, C0=>que_out_23_0_5, C1=>nx9952);
   ix9341 : aoi22 port map ( Y=>nx9340, A0=>que_out_27_0_5, A1=>nx9926, B0=>
      que_out_4_0_5, B1=>nx9900);
   ix9343 : aoi22 port map ( Y=>nx9342, A0=>que_out_0_0_5, A1=>nx9848, B0=>
      que_out_2_0_5, B1=>nx9874);
   ix7749 : nand03 port map ( Y=>nx7748, A0=>nx9345, A1=>nx9347, A2=>nx9349
   );
   ix9346 : aoi222 port map ( Y=>nx9345, A0=>que_out_26_0_5, A1=>nx9822, B0
      =>que_out_14_0_5, B1=>nx9796, C0=>que_out_11_0_5, C1=>nx9770);
   ix9348 : aoi22 port map ( Y=>nx9347, A0=>que_out_13_0_5, A1=>nx9744, B0=>
      que_out_7_0_5, B1=>nx9718);
   ix9350 : aoi22 port map ( Y=>nx9349, A0=>que_out_12_0_5, A1=>nx9692, B0=>
      que_out_1_0_5, B1=>nx9666);
   ix7943 : or04 port map ( Y=>out_column_0_6, A0=>nx7938, A1=>nx7912, A2=>
      nx7884, A3=>nx7858);
   ix7939 : nand03 port map ( Y=>nx7938, A0=>nx9353, A1=>nx9355, A2=>nx9357
   );
   ix9354 : aoi222 port map ( Y=>nx9353, A0=>que_out_10_0_6, A1=>nx10318, B0
      =>que_out_6_0_6, B1=>nx10370, C0=>que_out_9_0_6, C1=>nx10344);
   ix9356 : aoi22 port map ( Y=>nx9355, A0=>que_out_5_0_6, A1=>nx10266, B0=>
      que_out_18_0_6, B1=>nx10292);
   ix9358 : aoi22 port map ( Y=>nx9357, A0=>que_out_17_0_6, A1=>nx10240, B0
      =>que_out_20_0_6, B1=>nx10214);
   ix7913 : nand03 port map ( Y=>nx7912, A0=>nx9360, A1=>nx9362, A2=>nx9364
   );
   ix9361 : aoi222 port map ( Y=>nx9360, A0=>que_out_19_0_6, A1=>nx10188, B0
      =>que_out_21_0_6, B1=>nx10162, C0=>que_out_8_0_6, C1=>nx10136);
   ix9363 : aoi22 port map ( Y=>nx9362, A0=>que_out_25_0_6, A1=>nx10084, B0
      =>que_out_16_0_6, B1=>nx10110);
   ix9365 : aoi22 port map ( Y=>nx9364, A0=>que_out_24_0_6, A1=>nx10058, B0
      =>que_out_22_0_6, B1=>nx10032);
   ix7885 : nand03 port map ( Y=>nx7884, A0=>nx9367, A1=>nx9369, A2=>nx9371
   );
   ix9368 : aoi222 port map ( Y=>nx9367, A0=>que_out_15_0_6, A1=>nx9980, B0
      =>que_out_3_0_6, B1=>nx10006, C0=>que_out_23_0_6, C1=>nx9954);
   ix9370 : aoi22 port map ( Y=>nx9369, A0=>que_out_27_0_6, A1=>nx9928, B0=>
      que_out_4_0_6, B1=>nx9902);
   ix9372 : aoi22 port map ( Y=>nx9371, A0=>que_out_0_0_6, A1=>nx9850, B0=>
      que_out_2_0_6, B1=>nx9876);
   ix7859 : nand03 port map ( Y=>nx7858, A0=>nx9374, A1=>nx9376, A2=>nx9378
   );
   ix9375 : aoi222 port map ( Y=>nx9374, A0=>que_out_26_0_6, A1=>nx9824, B0
      =>que_out_14_0_6, B1=>nx9798, C0=>que_out_11_0_6, C1=>nx9772);
   ix9377 : aoi22 port map ( Y=>nx9376, A0=>que_out_13_0_6, A1=>nx9746, B0=>
      que_out_7_0_6, B1=>nx9720);
   ix9379 : aoi22 port map ( Y=>nx9378, A0=>que_out_12_0_6, A1=>nx9694, B0=>
      que_out_1_0_6, B1=>nx9668);
   ix8053 : or04 port map ( Y=>out_column_0_7, A0=>nx8048, A1=>nx8022, A2=>
      nx7994, A3=>nx7968);
   ix8049 : nand03 port map ( Y=>nx8048, A0=>nx9382, A1=>nx9384, A2=>nx9386
   );
   ix9383 : aoi222 port map ( Y=>nx9382, A0=>que_out_10_0_7, A1=>nx10318, B0
      =>que_out_6_0_7, B1=>nx10370, C0=>que_out_9_0_7, C1=>nx10344);
   ix9385 : aoi22 port map ( Y=>nx9384, A0=>que_out_5_0_7, A1=>nx10266, B0=>
      que_out_18_0_7, B1=>nx10292);
   ix9387 : aoi22 port map ( Y=>nx9386, A0=>que_out_17_0_7, A1=>nx10240, B0
      =>que_out_20_0_7, B1=>nx10214);
   ix8023 : nand03 port map ( Y=>nx8022, A0=>nx9389, A1=>nx9391, A2=>nx9393
   );
   ix9390 : aoi222 port map ( Y=>nx9389, A0=>que_out_19_0_7, A1=>nx10188, B0
      =>que_out_21_0_7, B1=>nx10162, C0=>que_out_8_0_7, C1=>nx10136);
   ix9392 : aoi22 port map ( Y=>nx9391, A0=>que_out_25_0_7, A1=>nx10084, B0
      =>que_out_16_0_7, B1=>nx10110);
   ix9394 : aoi22 port map ( Y=>nx9393, A0=>que_out_24_0_7, A1=>nx10058, B0
      =>que_out_22_0_7, B1=>nx10032);
   ix7995 : nand03 port map ( Y=>nx7994, A0=>nx9396, A1=>nx9398, A2=>nx9400
   );
   ix9397 : aoi222 port map ( Y=>nx9396, A0=>que_out_15_0_7, A1=>nx9980, B0
      =>que_out_3_0_7, B1=>nx10006, C0=>que_out_23_0_7, C1=>nx9954);
   ix9399 : aoi22 port map ( Y=>nx9398, A0=>que_out_27_0_7, A1=>nx9928, B0=>
      que_out_4_0_7, B1=>nx9902);
   ix9401 : aoi22 port map ( Y=>nx9400, A0=>que_out_0_0_7, A1=>nx9850, B0=>
      que_out_2_0_7, B1=>nx9876);
   ix7969 : nand03 port map ( Y=>nx7968, A0=>nx9403, A1=>nx9405, A2=>nx9407
   );
   ix9404 : aoi222 port map ( Y=>nx9403, A0=>que_out_26_0_7, A1=>nx9824, B0
      =>que_out_14_0_7, B1=>nx9798, C0=>que_out_11_0_7, C1=>nx9772);
   ix9406 : aoi22 port map ( Y=>nx9405, A0=>que_out_13_0_7, A1=>nx9746, B0=>
      que_out_7_0_7, B1=>nx9720);
   ix9408 : aoi22 port map ( Y=>nx9407, A0=>que_out_12_0_7, A1=>nx9694, B0=>
      que_out_1_0_7, B1=>nx9668);
   ix8163 : or04 port map ( Y=>out_column_0_8, A0=>nx8158, A1=>nx8132, A2=>
      nx8104, A3=>nx8078);
   ix8159 : nand03 port map ( Y=>nx8158, A0=>nx9411, A1=>nx9413, A2=>nx9415
   );
   ix9412 : aoi222 port map ( Y=>nx9411, A0=>que_out_10_0_8, A1=>nx10318, B0
      =>que_out_6_0_8, B1=>nx10370, C0=>que_out_9_0_8, C1=>nx10344);
   ix9414 : aoi22 port map ( Y=>nx9413, A0=>que_out_5_0_8, A1=>nx10266, B0=>
      que_out_18_0_8, B1=>nx10292);
   ix9416 : aoi22 port map ( Y=>nx9415, A0=>que_out_17_0_8, A1=>nx10240, B0
      =>que_out_20_0_8, B1=>nx10214);
   ix8133 : nand03 port map ( Y=>nx8132, A0=>nx9418, A1=>nx9420, A2=>nx9422
   );
   ix9419 : aoi222 port map ( Y=>nx9418, A0=>que_out_19_0_8, A1=>nx10188, B0
      =>que_out_21_0_8, B1=>nx10162, C0=>que_out_8_0_8, C1=>nx10136);
   ix9421 : aoi22 port map ( Y=>nx9420, A0=>que_out_25_0_8, A1=>nx10084, B0
      =>que_out_16_0_8, B1=>nx10110);
   ix9423 : aoi22 port map ( Y=>nx9422, A0=>que_out_24_0_8, A1=>nx10058, B0
      =>que_out_22_0_8, B1=>nx10032);
   ix8105 : nand03 port map ( Y=>nx8104, A0=>nx9425, A1=>nx9427, A2=>nx9429
   );
   ix9426 : aoi222 port map ( Y=>nx9425, A0=>que_out_15_0_8, A1=>nx9980, B0
      =>que_out_3_0_8, B1=>nx10006, C0=>que_out_23_0_8, C1=>nx9954);
   ix9428 : aoi22 port map ( Y=>nx9427, A0=>que_out_27_0_8, A1=>nx9928, B0=>
      que_out_4_0_8, B1=>nx9902);
   ix9430 : aoi22 port map ( Y=>nx9429, A0=>que_out_0_0_8, A1=>nx9850, B0=>
      que_out_2_0_8, B1=>nx9876);
   ix8079 : nand03 port map ( Y=>nx8078, A0=>nx9432, A1=>nx9434, A2=>nx9436
   );
   ix9433 : aoi222 port map ( Y=>nx9432, A0=>que_out_26_0_8, A1=>nx9824, B0
      =>que_out_14_0_8, B1=>nx9798, C0=>que_out_11_0_8, C1=>nx9772);
   ix9435 : aoi22 port map ( Y=>nx9434, A0=>que_out_13_0_8, A1=>nx9746, B0=>
      que_out_7_0_8, B1=>nx9720);
   ix9437 : aoi22 port map ( Y=>nx9436, A0=>que_out_12_0_8, A1=>nx9694, B0=>
      que_out_1_0_8, B1=>nx9668);
   ix8273 : or04 port map ( Y=>out_column_0_9, A0=>nx8268, A1=>nx8242, A2=>
      nx8214, A3=>nx8188);
   ix8269 : nand03 port map ( Y=>nx8268, A0=>nx9440, A1=>nx9442, A2=>nx9444
   );
   ix9441 : aoi222 port map ( Y=>nx9440, A0=>que_out_10_0_9, A1=>nx10318, B0
      =>que_out_6_0_9, B1=>nx10370, C0=>que_out_9_0_9, C1=>nx10344);
   ix9443 : aoi22 port map ( Y=>nx9442, A0=>que_out_5_0_9, A1=>nx10266, B0=>
      que_out_18_0_9, B1=>nx10292);
   ix9445 : aoi22 port map ( Y=>nx9444, A0=>que_out_17_0_9, A1=>nx10240, B0
      =>que_out_20_0_9, B1=>nx10214);
   ix8243 : nand03 port map ( Y=>nx8242, A0=>nx9447, A1=>nx9449, A2=>nx9451
   );
   ix9448 : aoi222 port map ( Y=>nx9447, A0=>que_out_19_0_9, A1=>nx10188, B0
      =>que_out_21_0_9, B1=>nx10162, C0=>que_out_8_0_9, C1=>nx10136);
   ix9450 : aoi22 port map ( Y=>nx9449, A0=>que_out_25_0_9, A1=>nx10084, B0
      =>que_out_16_0_9, B1=>nx10110);
   ix9452 : aoi22 port map ( Y=>nx9451, A0=>que_out_24_0_9, A1=>nx10058, B0
      =>que_out_22_0_9, B1=>nx10032);
   ix8215 : nand03 port map ( Y=>nx8214, A0=>nx9454, A1=>nx9456, A2=>nx9458
   );
   ix9455 : aoi222 port map ( Y=>nx9454, A0=>que_out_15_0_9, A1=>nx9980, B0
      =>que_out_3_0_9, B1=>nx10006, C0=>que_out_23_0_9, C1=>nx9954);
   ix9457 : aoi22 port map ( Y=>nx9456, A0=>que_out_27_0_9, A1=>nx9928, B0=>
      que_out_4_0_9, B1=>nx9902);
   ix9459 : aoi22 port map ( Y=>nx9458, A0=>que_out_0_0_9, A1=>nx9850, B0=>
      que_out_2_0_9, B1=>nx9876);
   ix8189 : nand03 port map ( Y=>nx8188, A0=>nx9461, A1=>nx9463, A2=>nx9465
   );
   ix9462 : aoi222 port map ( Y=>nx9461, A0=>que_out_26_0_9, A1=>nx9824, B0
      =>que_out_14_0_9, B1=>nx9798, C0=>que_out_11_0_9, C1=>nx9772);
   ix9464 : aoi22 port map ( Y=>nx9463, A0=>que_out_13_0_9, A1=>nx9746, B0=>
      que_out_7_0_9, B1=>nx9720);
   ix9466 : aoi22 port map ( Y=>nx9465, A0=>que_out_12_0_9, A1=>nx9694, B0=>
      que_out_1_0_9, B1=>nx9668);
   ix8383 : or04 port map ( Y=>out_column_0_10, A0=>nx8378, A1=>nx8352, A2=>
      nx8324, A3=>nx8298);
   ix8379 : nand03 port map ( Y=>nx8378, A0=>nx9469, A1=>nx9471, A2=>nx9473
   );
   ix9470 : aoi222 port map ( Y=>nx9469, A0=>que_out_10_0_10, A1=>nx10318, 
      B0=>que_out_6_0_10, B1=>nx10370, C0=>que_out_9_0_10, C1=>nx10344);
   ix9472 : aoi22 port map ( Y=>nx9471, A0=>que_out_5_0_10, A1=>nx10266, B0
      =>que_out_18_0_10, B1=>nx10292);
   ix9474 : aoi22 port map ( Y=>nx9473, A0=>que_out_17_0_10, A1=>nx10240, B0
      =>que_out_20_0_10, B1=>nx10214);
   ix8353 : nand03 port map ( Y=>nx8352, A0=>nx9476, A1=>nx9478, A2=>nx9480
   );
   ix9477 : aoi222 port map ( Y=>nx9476, A0=>que_out_19_0_10, A1=>nx10188, 
      B0=>que_out_21_0_10, B1=>nx10162, C0=>que_out_8_0_10, C1=>nx10136);
   ix9479 : aoi22 port map ( Y=>nx9478, A0=>que_out_25_0_10, A1=>nx10084, B0
      =>que_out_16_0_10, B1=>nx10110);
   ix9481 : aoi22 port map ( Y=>nx9480, A0=>que_out_24_0_10, A1=>nx10058, B0
      =>que_out_22_0_10, B1=>nx10032);
   ix8325 : nand03 port map ( Y=>nx8324, A0=>nx9483, A1=>nx9485, A2=>nx9487
   );
   ix9484 : aoi222 port map ( Y=>nx9483, A0=>que_out_15_0_10, A1=>nx9980, B0
      =>que_out_3_0_10, B1=>nx10006, C0=>que_out_23_0_10, C1=>nx9954);
   ix9486 : aoi22 port map ( Y=>nx9485, A0=>que_out_27_0_10, A1=>nx9928, B0
      =>que_out_4_0_10, B1=>nx9902);
   ix9488 : aoi22 port map ( Y=>nx9487, A0=>que_out_0_0_10, A1=>nx9850, B0=>
      que_out_2_0_10, B1=>nx9876);
   ix8299 : nand03 port map ( Y=>nx8298, A0=>nx9490, A1=>nx9492, A2=>nx9494
   );
   ix9491 : aoi222 port map ( Y=>nx9490, A0=>que_out_26_0_10, A1=>nx9824, B0
      =>que_out_14_0_10, B1=>nx9798, C0=>que_out_11_0_10, C1=>nx9772);
   ix9493 : aoi22 port map ( Y=>nx9492, A0=>que_out_13_0_10, A1=>nx9746, B0
      =>que_out_7_0_10, B1=>nx9720);
   ix9495 : aoi22 port map ( Y=>nx9494, A0=>que_out_12_0_10, A1=>nx9694, B0
      =>que_out_1_0_10, B1=>nx9668);
   ix8493 : or04 port map ( Y=>out_column_0_11, A0=>nx8488, A1=>nx8462, A2=>
      nx8434, A3=>nx8408);
   ix8489 : nand03 port map ( Y=>nx8488, A0=>nx9498, A1=>nx9500, A2=>nx9502
   );
   ix9499 : aoi222 port map ( Y=>nx9498, A0=>que_out_10_0_11, A1=>nx10318, 
      B0=>que_out_6_0_11, B1=>nx10370, C0=>que_out_9_0_11, C1=>nx10344);
   ix9501 : aoi22 port map ( Y=>nx9500, A0=>que_out_5_0_11, A1=>nx10266, B0
      =>que_out_18_0_11, B1=>nx10292);
   ix9503 : aoi22 port map ( Y=>nx9502, A0=>que_out_17_0_11, A1=>nx10240, B0
      =>que_out_20_0_11, B1=>nx10214);
   ix8463 : nand03 port map ( Y=>nx8462, A0=>nx9505, A1=>nx9507, A2=>nx9509
   );
   ix9506 : aoi222 port map ( Y=>nx9505, A0=>que_out_19_0_11, A1=>nx10188, 
      B0=>que_out_21_0_11, B1=>nx10162, C0=>que_out_8_0_11, C1=>nx10136);
   ix9508 : aoi22 port map ( Y=>nx9507, A0=>que_out_25_0_11, A1=>nx10084, B0
      =>que_out_16_0_11, B1=>nx10110);
   ix9510 : aoi22 port map ( Y=>nx9509, A0=>que_out_24_0_11, A1=>nx10058, B0
      =>que_out_22_0_11, B1=>nx10032);
   ix8435 : nand03 port map ( Y=>nx8434, A0=>nx9512, A1=>nx9514, A2=>nx9516
   );
   ix9513 : aoi222 port map ( Y=>nx9512, A0=>que_out_15_0_11, A1=>nx9980, B0
      =>que_out_3_0_11, B1=>nx10006, C0=>que_out_23_0_11, C1=>nx9954);
   ix9515 : aoi22 port map ( Y=>nx9514, A0=>que_out_27_0_11, A1=>nx9928, B0
      =>que_out_4_0_11, B1=>nx9902);
   ix9517 : aoi22 port map ( Y=>nx9516, A0=>que_out_0_0_11, A1=>nx9850, B0=>
      que_out_2_0_11, B1=>nx9876);
   ix8409 : nand03 port map ( Y=>nx8408, A0=>nx9519, A1=>nx9521, A2=>nx9523
   );
   ix9520 : aoi222 port map ( Y=>nx9519, A0=>que_out_26_0_11, A1=>nx9824, B0
      =>que_out_14_0_11, B1=>nx9798, C0=>que_out_11_0_11, C1=>nx9772);
   ix9522 : aoi22 port map ( Y=>nx9521, A0=>que_out_13_0_11, A1=>nx9746, B0
      =>que_out_7_0_11, B1=>nx9720);
   ix9524 : aoi22 port map ( Y=>nx9523, A0=>que_out_12_0_11, A1=>nx9694, B0
      =>que_out_1_0_11, B1=>nx9668);
   ix8603 : or04 port map ( Y=>out_column_0_12, A0=>nx8598, A1=>nx8572, A2=>
      nx8544, A3=>nx8518);
   ix8599 : nand03 port map ( Y=>nx8598, A0=>nx9527, A1=>nx9529, A2=>nx9531
   );
   ix9528 : aoi222 port map ( Y=>nx9527, A0=>que_out_10_0_12, A1=>nx10318, 
      B0=>que_out_6_0_12, B1=>nx10370, C0=>que_out_9_0_12, C1=>nx10344);
   ix9530 : aoi22 port map ( Y=>nx9529, A0=>que_out_5_0_12, A1=>nx10266, B0
      =>que_out_18_0_12, B1=>nx10292);
   ix9532 : aoi22 port map ( Y=>nx9531, A0=>que_out_17_0_12, A1=>nx10240, B0
      =>que_out_20_0_12, B1=>nx10214);
   ix8573 : nand03 port map ( Y=>nx8572, A0=>nx9534, A1=>nx9536, A2=>nx9538
   );
   ix9535 : aoi222 port map ( Y=>nx9534, A0=>que_out_19_0_12, A1=>nx10188, 
      B0=>que_out_21_0_12, B1=>nx10162, C0=>que_out_8_0_12, C1=>nx10136);
   ix9537 : aoi22 port map ( Y=>nx9536, A0=>que_out_25_0_12, A1=>nx10084, B0
      =>que_out_16_0_12, B1=>nx10110);
   ix9539 : aoi22 port map ( Y=>nx9538, A0=>que_out_24_0_12, A1=>nx10058, B0
      =>que_out_22_0_12, B1=>nx10032);
   ix8545 : nand03 port map ( Y=>nx8544, A0=>nx9541, A1=>nx9543, A2=>nx9545
   );
   ix9542 : aoi222 port map ( Y=>nx9541, A0=>que_out_15_0_12, A1=>nx9980, B0
      =>que_out_3_0_12, B1=>nx10006, C0=>que_out_23_0_12, C1=>nx9954);
   ix9544 : aoi22 port map ( Y=>nx9543, A0=>que_out_27_0_12, A1=>nx9928, B0
      =>que_out_4_0_12, B1=>nx9902);
   ix9546 : aoi22 port map ( Y=>nx9545, A0=>que_out_0_0_12, A1=>nx9850, B0=>
      que_out_2_0_12, B1=>nx9876);
   ix8519 : nand03 port map ( Y=>nx8518, A0=>nx9548, A1=>nx9550, A2=>nx9552
   );
   ix9549 : aoi222 port map ( Y=>nx9548, A0=>que_out_26_0_12, A1=>nx9824, B0
      =>que_out_14_0_12, B1=>nx9798, C0=>que_out_11_0_12, C1=>nx9772);
   ix9551 : aoi22 port map ( Y=>nx9550, A0=>que_out_13_0_12, A1=>nx9746, B0
      =>que_out_7_0_12, B1=>nx9720);
   ix9553 : aoi22 port map ( Y=>nx9552, A0=>que_out_12_0_12, A1=>nx9694, B0
      =>que_out_1_0_12, B1=>nx9668);
   ix8713 : or04 port map ( Y=>out_column_0_13, A0=>nx8708, A1=>nx8682, A2=>
      nx8654, A3=>nx8628);
   ix8709 : nand03 port map ( Y=>nx8708, A0=>nx9556, A1=>nx9558, A2=>nx9560
   );
   ix9557 : aoi222 port map ( Y=>nx9556, A0=>que_out_10_0_13, A1=>nx10320, 
      B0=>que_out_6_0_13, B1=>nx10372, C0=>que_out_9_0_13, C1=>nx10346);
   ix9559 : aoi22 port map ( Y=>nx9558, A0=>que_out_5_0_13, A1=>nx10268, B0
      =>que_out_18_0_13, B1=>nx10294);
   ix9561 : aoi22 port map ( Y=>nx9560, A0=>que_out_17_0_13, A1=>nx10242, B0
      =>que_out_20_0_13, B1=>nx10216);
   ix8683 : nand03 port map ( Y=>nx8682, A0=>nx9563, A1=>nx9565, A2=>nx9567
   );
   ix9564 : aoi222 port map ( Y=>nx9563, A0=>que_out_19_0_13, A1=>nx10190, 
      B0=>que_out_21_0_13, B1=>nx10164, C0=>que_out_8_0_13, C1=>nx10138);
   ix9566 : aoi22 port map ( Y=>nx9565, A0=>que_out_25_0_13, A1=>nx10086, B0
      =>que_out_16_0_13, B1=>nx10112);
   ix9568 : aoi22 port map ( Y=>nx9567, A0=>que_out_24_0_13, A1=>nx10060, B0
      =>que_out_22_0_13, B1=>nx10034);
   ix8655 : nand03 port map ( Y=>nx8654, A0=>nx9570, A1=>nx9572, A2=>nx9574
   );
   ix9571 : aoi222 port map ( Y=>nx9570, A0=>que_out_15_0_13, A1=>nx9982, B0
      =>que_out_3_0_13, B1=>nx10008, C0=>que_out_23_0_13, C1=>nx9956);
   ix9573 : aoi22 port map ( Y=>nx9572, A0=>que_out_27_0_13, A1=>nx9930, B0
      =>que_out_4_0_13, B1=>nx9904);
   ix9575 : aoi22 port map ( Y=>nx9574, A0=>que_out_0_0_13, A1=>nx9852, B0=>
      que_out_2_0_13, B1=>nx9878);
   ix8629 : nand03 port map ( Y=>nx8628, A0=>nx9577, A1=>nx9579, A2=>nx9581
   );
   ix9578 : aoi222 port map ( Y=>nx9577, A0=>que_out_26_0_13, A1=>nx9826, B0
      =>que_out_14_0_13, B1=>nx9800, C0=>que_out_11_0_13, C1=>nx9774);
   ix9580 : aoi22 port map ( Y=>nx9579, A0=>que_out_13_0_13, A1=>nx9748, B0
      =>que_out_7_0_13, B1=>nx9722);
   ix9582 : aoi22 port map ( Y=>nx9581, A0=>que_out_12_0_13, A1=>nx9696, B0
      =>que_out_1_0_13, B1=>nx9670);
   ix8823 : or04 port map ( Y=>out_column_0_14, A0=>nx8818, A1=>nx8792, A2=>
      nx8764, A3=>nx8738);
   ix8819 : nand03 port map ( Y=>nx8818, A0=>nx9585, A1=>nx9587, A2=>nx9589
   );
   ix9586 : aoi222 port map ( Y=>nx9585, A0=>que_out_10_0_14, A1=>nx10320, 
      B0=>que_out_6_0_14, B1=>nx10372, C0=>que_out_9_0_14, C1=>nx10346);
   ix9588 : aoi22 port map ( Y=>nx9587, A0=>que_out_5_0_14, A1=>nx10268, B0
      =>que_out_18_0_14, B1=>nx10294);
   ix9590 : aoi22 port map ( Y=>nx9589, A0=>que_out_17_0_14, A1=>nx10242, B0
      =>que_out_20_0_14, B1=>nx10216);
   ix8793 : nand03 port map ( Y=>nx8792, A0=>nx9592, A1=>nx9594, A2=>nx9596
   );
   ix9593 : aoi222 port map ( Y=>nx9592, A0=>que_out_19_0_14, A1=>nx10190, 
      B0=>que_out_21_0_14, B1=>nx10164, C0=>que_out_8_0_14, C1=>nx10138);
   ix9595 : aoi22 port map ( Y=>nx9594, A0=>que_out_25_0_14, A1=>nx10086, B0
      =>que_out_16_0_14, B1=>nx10112);
   ix9597 : aoi22 port map ( Y=>nx9596, A0=>que_out_24_0_14, A1=>nx10060, B0
      =>que_out_22_0_14, B1=>nx10034);
   ix8765 : nand03 port map ( Y=>nx8764, A0=>nx9599, A1=>nx9601, A2=>nx9603
   );
   ix9600 : aoi222 port map ( Y=>nx9599, A0=>que_out_15_0_14, A1=>nx9982, B0
      =>que_out_3_0_14, B1=>nx10008, C0=>que_out_23_0_14, C1=>nx9956);
   ix9602 : aoi22 port map ( Y=>nx9601, A0=>que_out_27_0_14, A1=>nx9930, B0
      =>que_out_4_0_14, B1=>nx9904);
   ix9604 : aoi22 port map ( Y=>nx9603, A0=>que_out_0_0_14, A1=>nx9852, B0=>
      que_out_2_0_14, B1=>nx9878);
   ix8739 : nand03 port map ( Y=>nx8738, A0=>nx9606, A1=>nx9608, A2=>nx9610
   );
   ix9607 : aoi222 port map ( Y=>nx9606, A0=>que_out_26_0_14, A1=>nx9826, B0
      =>que_out_14_0_14, B1=>nx9800, C0=>que_out_11_0_14, C1=>nx9774);
   ix9609 : aoi22 port map ( Y=>nx9608, A0=>que_out_13_0_14, A1=>nx9748, B0
      =>que_out_7_0_14, B1=>nx9722);
   ix9611 : aoi22 port map ( Y=>nx9610, A0=>que_out_12_0_14, A1=>nx9696, B0
      =>que_out_1_0_14, B1=>nx9670);
   ix8933 : or04 port map ( Y=>out_column_0_15, A0=>nx8928, A1=>nx8902, A2=>
      nx8874, A3=>nx8848);
   ix8929 : nand03 port map ( Y=>nx8928, A0=>nx9614, A1=>nx9616, A2=>nx9618
   );
   ix9615 : aoi222 port map ( Y=>nx9614, A0=>que_out_10_0_15, A1=>nx10320, 
      B0=>que_out_6_0_15, B1=>nx10372, C0=>que_out_9_0_15, C1=>nx10346);
   ix9617 : aoi22 port map ( Y=>nx9616, A0=>que_out_5_0_15, A1=>nx10268, B0
      =>que_out_18_0_15, B1=>nx10294);
   ix9619 : aoi22 port map ( Y=>nx9618, A0=>que_out_17_0_15, A1=>nx10242, B0
      =>que_out_20_0_15, B1=>nx10216);
   ix8903 : nand03 port map ( Y=>nx8902, A0=>nx9621, A1=>nx9623, A2=>nx9625
   );
   ix9622 : aoi222 port map ( Y=>nx9621, A0=>que_out_19_0_15, A1=>nx10190, 
      B0=>que_out_21_0_15, B1=>nx10164, C0=>que_out_8_0_15, C1=>nx10138);
   ix9624 : aoi22 port map ( Y=>nx9623, A0=>que_out_25_0_15, A1=>nx10086, B0
      =>que_out_16_0_15, B1=>nx10112);
   ix9626 : aoi22 port map ( Y=>nx9625, A0=>que_out_24_0_15, A1=>nx10060, B0
      =>que_out_22_0_15, B1=>nx10034);
   ix8875 : nand03 port map ( Y=>nx8874, A0=>nx9628, A1=>nx9630, A2=>nx9632
   );
   ix9629 : aoi222 port map ( Y=>nx9628, A0=>que_out_15_0_15, A1=>nx9982, B0
      =>que_out_3_0_15, B1=>nx10008, C0=>que_out_23_0_15, C1=>nx9956);
   ix9631 : aoi22 port map ( Y=>nx9630, A0=>que_out_27_0_15, A1=>nx9930, B0
      =>que_out_4_0_15, B1=>nx9904);
   ix9633 : aoi22 port map ( Y=>nx9632, A0=>que_out_0_0_15, A1=>nx9852, B0=>
      que_out_2_0_15, B1=>nx9878);
   ix8849 : nand03 port map ( Y=>nx8848, A0=>nx9635, A1=>nx9637, A2=>nx9639
   );
   ix9636 : aoi222 port map ( Y=>nx9635, A0=>que_out_26_0_15, A1=>nx9826, B0
      =>que_out_14_0_15, B1=>nx9800, C0=>que_out_11_0_15, C1=>nx9774);
   ix9638 : aoi22 port map ( Y=>nx9637, A0=>que_out_13_0_15, A1=>nx9748, B0
      =>que_out_7_0_15, B1=>nx9722);
   ix9640 : aoi22 port map ( Y=>nx9639, A0=>que_out_12_0_15, A1=>nx9696, B0
      =>que_out_1_0_15, B1=>nx9670);
   ix6944 : inv02 port map ( Y=>nx6943, A=>nx88);
   ix9647 : inv02 port map ( Y=>nx9648, A=>nx10378);
   ix9649 : inv02 port map ( Y=>nx9650, A=>nx10378);
   ix9651 : inv02 port map ( Y=>nx9652, A=>nx10378);
   ix9653 : inv02 port map ( Y=>nx9654, A=>nx10378);
   ix9655 : inv02 port map ( Y=>nx9656, A=>nx10378);
   ix9657 : inv02 port map ( Y=>nx9658, A=>nx10378);
   ix9659 : inv02 port map ( Y=>nx9660, A=>nx10378);
   ix9661 : inv02 port map ( Y=>nx9662, A=>nx10380);
   ix9663 : inv02 port map ( Y=>nx9664, A=>nx10380);
   ix9665 : inv02 port map ( Y=>nx9666, A=>nx10380);
   ix9667 : inv02 port map ( Y=>nx9668, A=>nx10380);
   ix9669 : inv02 port map ( Y=>nx9670, A=>nx10380);
   ix9673 : inv02 port map ( Y=>nx9674, A=>nx10382);
   ix9675 : inv02 port map ( Y=>nx9676, A=>nx10382);
   ix9677 : inv02 port map ( Y=>nx9678, A=>nx10382);
   ix9679 : inv02 port map ( Y=>nx9680, A=>nx10382);
   ix9681 : inv02 port map ( Y=>nx9682, A=>nx10382);
   ix9683 : inv02 port map ( Y=>nx9684, A=>nx10382);
   ix9685 : inv02 port map ( Y=>nx9686, A=>nx10382);
   ix9687 : inv02 port map ( Y=>nx9688, A=>nx10384);
   ix9689 : inv02 port map ( Y=>nx9690, A=>nx10384);
   ix9691 : inv02 port map ( Y=>nx9692, A=>nx10384);
   ix9693 : inv02 port map ( Y=>nx9694, A=>nx10384);
   ix9695 : inv02 port map ( Y=>nx9696, A=>nx10384);
   ix9699 : inv02 port map ( Y=>nx9700, A=>nx10386);
   ix9701 : inv02 port map ( Y=>nx9702, A=>nx10386);
   ix9703 : inv02 port map ( Y=>nx9704, A=>nx10386);
   ix9705 : inv02 port map ( Y=>nx9706, A=>nx10386);
   ix9707 : inv02 port map ( Y=>nx9708, A=>nx10386);
   ix9709 : inv02 port map ( Y=>nx9710, A=>nx10386);
   ix9711 : inv02 port map ( Y=>nx9712, A=>nx10386);
   ix9713 : inv02 port map ( Y=>nx9714, A=>nx10388);
   ix9715 : inv02 port map ( Y=>nx9716, A=>nx10388);
   ix9717 : inv02 port map ( Y=>nx9718, A=>nx10388);
   ix9719 : inv02 port map ( Y=>nx9720, A=>nx10388);
   ix9721 : inv02 port map ( Y=>nx9722, A=>nx10388);
   ix9725 : inv02 port map ( Y=>nx9726, A=>nx10390);
   ix9727 : inv02 port map ( Y=>nx9728, A=>nx10390);
   ix9729 : inv02 port map ( Y=>nx9730, A=>nx10390);
   ix9731 : inv02 port map ( Y=>nx9732, A=>nx10390);
   ix9733 : inv02 port map ( Y=>nx9734, A=>nx10390);
   ix9735 : inv02 port map ( Y=>nx9736, A=>nx10390);
   ix9737 : inv02 port map ( Y=>nx9738, A=>nx10390);
   ix9739 : inv02 port map ( Y=>nx9740, A=>nx10392);
   ix9741 : inv02 port map ( Y=>nx9742, A=>nx10392);
   ix9743 : inv02 port map ( Y=>nx9744, A=>nx10392);
   ix9745 : inv02 port map ( Y=>nx9746, A=>nx10392);
   ix9747 : inv02 port map ( Y=>nx9748, A=>nx10392);
   ix9751 : inv02 port map ( Y=>nx9752, A=>nx10394);
   ix9753 : inv02 port map ( Y=>nx9754, A=>nx10394);
   ix9755 : inv02 port map ( Y=>nx9756, A=>nx10394);
   ix9757 : inv02 port map ( Y=>nx9758, A=>nx10394);
   ix9759 : inv02 port map ( Y=>nx9760, A=>nx10394);
   ix9761 : inv02 port map ( Y=>nx9762, A=>nx10394);
   ix9763 : inv02 port map ( Y=>nx9764, A=>nx10394);
   ix9765 : inv02 port map ( Y=>nx9766, A=>nx10396);
   ix9767 : inv02 port map ( Y=>nx9768, A=>nx10396);
   ix9769 : inv02 port map ( Y=>nx9770, A=>nx10396);
   ix9771 : inv02 port map ( Y=>nx9772, A=>nx10396);
   ix9773 : inv02 port map ( Y=>nx9774, A=>nx10396);
   ix9777 : inv02 port map ( Y=>nx9778, A=>nx10398);
   ix9779 : inv02 port map ( Y=>nx9780, A=>nx10398);
   ix9781 : inv02 port map ( Y=>nx9782, A=>nx10398);
   ix9783 : inv02 port map ( Y=>nx9784, A=>nx10398);
   ix9785 : inv02 port map ( Y=>nx9786, A=>nx10398);
   ix9787 : inv02 port map ( Y=>nx9788, A=>nx10398);
   ix9789 : inv02 port map ( Y=>nx9790, A=>nx10398);
   ix9791 : inv02 port map ( Y=>nx9792, A=>nx10400);
   ix9793 : inv02 port map ( Y=>nx9794, A=>nx10400);
   ix9795 : inv02 port map ( Y=>nx9796, A=>nx10400);
   ix9797 : inv02 port map ( Y=>nx9798, A=>nx10400);
   ix9799 : inv02 port map ( Y=>nx9800, A=>nx10400);
   ix9803 : inv02 port map ( Y=>nx9804, A=>nx10402);
   ix9805 : inv02 port map ( Y=>nx9806, A=>nx10402);
   ix9807 : inv02 port map ( Y=>nx9808, A=>nx10402);
   ix9809 : inv02 port map ( Y=>nx9810, A=>nx10402);
   ix9811 : inv02 port map ( Y=>nx9812, A=>nx10402);
   ix9813 : inv02 port map ( Y=>nx9814, A=>nx10402);
   ix9815 : inv02 port map ( Y=>nx9816, A=>nx10402);
   ix9817 : inv02 port map ( Y=>nx9818, A=>nx10404);
   ix9819 : inv02 port map ( Y=>nx9820, A=>nx10404);
   ix9821 : inv02 port map ( Y=>nx9822, A=>nx10404);
   ix9823 : inv02 port map ( Y=>nx9824, A=>nx10404);
   ix9825 : inv02 port map ( Y=>nx9826, A=>nx10404);
   ix9829 : inv02 port map ( Y=>nx9830, A=>nx10406);
   ix9831 : inv02 port map ( Y=>nx9832, A=>nx10406);
   ix9833 : inv02 port map ( Y=>nx9834, A=>nx10406);
   ix9835 : inv02 port map ( Y=>nx9836, A=>nx10406);
   ix9837 : inv02 port map ( Y=>nx9838, A=>nx10406);
   ix9839 : inv02 port map ( Y=>nx9840, A=>nx10406);
   ix9841 : inv02 port map ( Y=>nx9842, A=>nx10406);
   ix9843 : inv02 port map ( Y=>nx9844, A=>nx10408);
   ix9845 : inv02 port map ( Y=>nx9846, A=>nx10408);
   ix9847 : inv02 port map ( Y=>nx9848, A=>nx10408);
   ix9849 : inv02 port map ( Y=>nx9850, A=>nx10408);
   ix9851 : inv02 port map ( Y=>nx9852, A=>nx10408);
   ix9855 : inv02 port map ( Y=>nx9856, A=>nx10410);
   ix9857 : inv02 port map ( Y=>nx9858, A=>nx10410);
   ix9859 : inv02 port map ( Y=>nx9860, A=>nx10410);
   ix9861 : inv02 port map ( Y=>nx9862, A=>nx10410);
   ix9863 : inv02 port map ( Y=>nx9864, A=>nx10410);
   ix9865 : inv02 port map ( Y=>nx9866, A=>nx10410);
   ix9867 : inv02 port map ( Y=>nx9868, A=>nx10410);
   ix9869 : inv02 port map ( Y=>nx9870, A=>nx10412);
   ix9871 : inv02 port map ( Y=>nx9872, A=>nx10412);
   ix9873 : inv02 port map ( Y=>nx9874, A=>nx10412);
   ix9875 : inv02 port map ( Y=>nx9876, A=>nx10412);
   ix9877 : inv02 port map ( Y=>nx9878, A=>nx10412);
   ix9881 : inv02 port map ( Y=>nx9882, A=>nx10414);
   ix9883 : inv02 port map ( Y=>nx9884, A=>nx10414);
   ix9885 : inv02 port map ( Y=>nx9886, A=>nx10414);
   ix9887 : inv02 port map ( Y=>nx9888, A=>nx10414);
   ix9889 : inv02 port map ( Y=>nx9890, A=>nx10414);
   ix9891 : inv02 port map ( Y=>nx9892, A=>nx10414);
   ix9893 : inv02 port map ( Y=>nx9894, A=>nx10414);
   ix9895 : inv02 port map ( Y=>nx9896, A=>nx10416);
   ix9897 : inv02 port map ( Y=>nx9898, A=>nx10416);
   ix9899 : inv02 port map ( Y=>nx9900, A=>nx10416);
   ix9901 : inv02 port map ( Y=>nx9902, A=>nx10416);
   ix9903 : inv02 port map ( Y=>nx9904, A=>nx10416);
   ix9907 : inv02 port map ( Y=>nx9908, A=>nx10418);
   ix9909 : inv02 port map ( Y=>nx9910, A=>nx10418);
   ix9911 : inv02 port map ( Y=>nx9912, A=>nx10418);
   ix9913 : inv02 port map ( Y=>nx9914, A=>nx10418);
   ix9915 : inv02 port map ( Y=>nx9916, A=>nx10418);
   ix9917 : inv02 port map ( Y=>nx9918, A=>nx10418);
   ix9919 : inv02 port map ( Y=>nx9920, A=>nx10418);
   ix9921 : inv02 port map ( Y=>nx9922, A=>nx10420);
   ix9923 : inv02 port map ( Y=>nx9924, A=>nx10420);
   ix9925 : inv02 port map ( Y=>nx9926, A=>nx10420);
   ix9927 : inv02 port map ( Y=>nx9928, A=>nx10420);
   ix9929 : inv02 port map ( Y=>nx9930, A=>nx10420);
   ix9933 : inv02 port map ( Y=>nx9934, A=>nx10422);
   ix9935 : inv02 port map ( Y=>nx9936, A=>nx10422);
   ix9937 : inv02 port map ( Y=>nx9938, A=>nx10422);
   ix9939 : inv02 port map ( Y=>nx9940, A=>nx10422);
   ix9941 : inv02 port map ( Y=>nx9942, A=>nx10422);
   ix9943 : inv02 port map ( Y=>nx9944, A=>nx10422);
   ix9945 : inv02 port map ( Y=>nx9946, A=>nx10422);
   ix9947 : inv02 port map ( Y=>nx9948, A=>nx10424);
   ix9949 : inv02 port map ( Y=>nx9950, A=>nx10424);
   ix9951 : inv02 port map ( Y=>nx9952, A=>nx10424);
   ix9953 : inv02 port map ( Y=>nx9954, A=>nx10424);
   ix9955 : inv02 port map ( Y=>nx9956, A=>nx10424);
   ix9959 : inv02 port map ( Y=>nx9960, A=>nx10426);
   ix9961 : inv02 port map ( Y=>nx9962, A=>nx10426);
   ix9963 : inv02 port map ( Y=>nx9964, A=>nx10426);
   ix9965 : inv02 port map ( Y=>nx9966, A=>nx10426);
   ix9967 : inv02 port map ( Y=>nx9968, A=>nx10426);
   ix9969 : inv02 port map ( Y=>nx9970, A=>nx10426);
   ix9971 : inv02 port map ( Y=>nx9972, A=>nx10426);
   ix9973 : inv02 port map ( Y=>nx9974, A=>nx10428);
   ix9975 : inv02 port map ( Y=>nx9976, A=>nx10428);
   ix9977 : inv02 port map ( Y=>nx9978, A=>nx10428);
   ix9979 : inv02 port map ( Y=>nx9980, A=>nx10428);
   ix9981 : inv02 port map ( Y=>nx9982, A=>nx10428);
   ix9985 : inv02 port map ( Y=>nx9986, A=>nx10430);
   ix9987 : inv02 port map ( Y=>nx9988, A=>nx10430);
   ix9989 : inv02 port map ( Y=>nx9990, A=>nx10430);
   ix9991 : inv02 port map ( Y=>nx9992, A=>nx10430);
   ix9993 : inv02 port map ( Y=>nx9994, A=>nx10430);
   ix9995 : inv02 port map ( Y=>nx9996, A=>nx10430);
   ix9997 : inv02 port map ( Y=>nx9998, A=>nx10430);
   ix9999 : inv02 port map ( Y=>nx10000, A=>nx10432);
   ix10001 : inv02 port map ( Y=>nx10002, A=>nx10432);
   ix10003 : inv02 port map ( Y=>nx10004, A=>nx10432);
   ix10005 : inv02 port map ( Y=>nx10006, A=>nx10432);
   ix10007 : inv02 port map ( Y=>nx10008, A=>nx10432);
   ix10011 : inv02 port map ( Y=>nx10012, A=>nx10434);
   ix10013 : inv02 port map ( Y=>nx10014, A=>nx10434);
   ix10015 : inv02 port map ( Y=>nx10016, A=>nx10434);
   ix10017 : inv02 port map ( Y=>nx10018, A=>nx10434);
   ix10019 : inv02 port map ( Y=>nx10020, A=>nx10434);
   ix10021 : inv02 port map ( Y=>nx10022, A=>nx10434);
   ix10023 : inv02 port map ( Y=>nx10024, A=>nx10434);
   ix10025 : inv02 port map ( Y=>nx10026, A=>nx10436);
   ix10027 : inv02 port map ( Y=>nx10028, A=>nx10436);
   ix10029 : inv02 port map ( Y=>nx10030, A=>nx10436);
   ix10031 : inv02 port map ( Y=>nx10032, A=>nx10436);
   ix10033 : inv02 port map ( Y=>nx10034, A=>nx10436);
   ix10037 : inv02 port map ( Y=>nx10038, A=>nx10438);
   ix10039 : inv02 port map ( Y=>nx10040, A=>nx10438);
   ix10041 : inv02 port map ( Y=>nx10042, A=>nx10438);
   ix10043 : inv02 port map ( Y=>nx10044, A=>nx10438);
   ix10045 : inv02 port map ( Y=>nx10046, A=>nx10438);
   ix10047 : inv02 port map ( Y=>nx10048, A=>nx10438);
   ix10049 : inv02 port map ( Y=>nx10050, A=>nx10438);
   ix10051 : inv02 port map ( Y=>nx10052, A=>nx10440);
   ix10053 : inv02 port map ( Y=>nx10054, A=>nx10440);
   ix10055 : inv02 port map ( Y=>nx10056, A=>nx10440);
   ix10057 : inv02 port map ( Y=>nx10058, A=>nx10440);
   ix10059 : inv02 port map ( Y=>nx10060, A=>nx10440);
   ix10063 : inv02 port map ( Y=>nx10064, A=>nx10442);
   ix10065 : inv02 port map ( Y=>nx10066, A=>nx10442);
   ix10067 : inv02 port map ( Y=>nx10068, A=>nx10442);
   ix10069 : inv02 port map ( Y=>nx10070, A=>nx10442);
   ix10071 : inv02 port map ( Y=>nx10072, A=>nx10442);
   ix10073 : inv02 port map ( Y=>nx10074, A=>nx10442);
   ix10075 : inv02 port map ( Y=>nx10076, A=>nx10442);
   ix10077 : inv02 port map ( Y=>nx10078, A=>nx10444);
   ix10079 : inv02 port map ( Y=>nx10080, A=>nx10444);
   ix10081 : inv02 port map ( Y=>nx10082, A=>nx10444);
   ix10083 : inv02 port map ( Y=>nx10084, A=>nx10444);
   ix10085 : inv02 port map ( Y=>nx10086, A=>nx10444);
   ix10089 : inv02 port map ( Y=>nx10090, A=>nx10446);
   ix10091 : inv02 port map ( Y=>nx10092, A=>nx10446);
   ix10093 : inv02 port map ( Y=>nx10094, A=>nx10446);
   ix10095 : inv02 port map ( Y=>nx10096, A=>nx10446);
   ix10097 : inv02 port map ( Y=>nx10098, A=>nx10446);
   ix10099 : inv02 port map ( Y=>nx10100, A=>nx10446);
   ix10101 : inv02 port map ( Y=>nx10102, A=>nx10446);
   ix10103 : inv02 port map ( Y=>nx10104, A=>nx10448);
   ix10105 : inv02 port map ( Y=>nx10106, A=>nx10448);
   ix10107 : inv02 port map ( Y=>nx10108, A=>nx10448);
   ix10109 : inv02 port map ( Y=>nx10110, A=>nx10448);
   ix10111 : inv02 port map ( Y=>nx10112, A=>nx10448);
   ix10115 : inv02 port map ( Y=>nx10116, A=>nx10450);
   ix10117 : inv02 port map ( Y=>nx10118, A=>nx10450);
   ix10119 : inv02 port map ( Y=>nx10120, A=>nx10450);
   ix10121 : inv02 port map ( Y=>nx10122, A=>nx10450);
   ix10123 : inv02 port map ( Y=>nx10124, A=>nx10450);
   ix10125 : inv02 port map ( Y=>nx10126, A=>nx10450);
   ix10127 : inv02 port map ( Y=>nx10128, A=>nx10450);
   ix10129 : inv02 port map ( Y=>nx10130, A=>nx10452);
   ix10131 : inv02 port map ( Y=>nx10132, A=>nx10452);
   ix10133 : inv02 port map ( Y=>nx10134, A=>nx10452);
   ix10135 : inv02 port map ( Y=>nx10136, A=>nx10452);
   ix10137 : inv02 port map ( Y=>nx10138, A=>nx10452);
   ix10141 : inv02 port map ( Y=>nx10142, A=>nx10454);
   ix10143 : inv02 port map ( Y=>nx10144, A=>nx10454);
   ix10145 : inv02 port map ( Y=>nx10146, A=>nx10454);
   ix10147 : inv02 port map ( Y=>nx10148, A=>nx10454);
   ix10149 : inv02 port map ( Y=>nx10150, A=>nx10454);
   ix10151 : inv02 port map ( Y=>nx10152, A=>nx10454);
   ix10153 : inv02 port map ( Y=>nx10154, A=>nx10454);
   ix10155 : inv02 port map ( Y=>nx10156, A=>nx10456);
   ix10157 : inv02 port map ( Y=>nx10158, A=>nx10456);
   ix10159 : inv02 port map ( Y=>nx10160, A=>nx10456);
   ix10161 : inv02 port map ( Y=>nx10162, A=>nx10456);
   ix10163 : inv02 port map ( Y=>nx10164, A=>nx10456);
   ix10167 : inv02 port map ( Y=>nx10168, A=>nx10458);
   ix10169 : inv02 port map ( Y=>nx10170, A=>nx10458);
   ix10171 : inv02 port map ( Y=>nx10172, A=>nx10458);
   ix10173 : inv02 port map ( Y=>nx10174, A=>nx10458);
   ix10175 : inv02 port map ( Y=>nx10176, A=>nx10458);
   ix10177 : inv02 port map ( Y=>nx10178, A=>nx10458);
   ix10179 : inv02 port map ( Y=>nx10180, A=>nx10458);
   ix10181 : inv02 port map ( Y=>nx10182, A=>nx10460);
   ix10183 : inv02 port map ( Y=>nx10184, A=>nx10460);
   ix10185 : inv02 port map ( Y=>nx10186, A=>nx10460);
   ix10187 : inv02 port map ( Y=>nx10188, A=>nx10460);
   ix10189 : inv02 port map ( Y=>nx10190, A=>nx10460);
   ix10193 : inv02 port map ( Y=>nx10194, A=>nx10462);
   ix10195 : inv02 port map ( Y=>nx10196, A=>nx10462);
   ix10197 : inv02 port map ( Y=>nx10198, A=>nx10462);
   ix10199 : inv02 port map ( Y=>nx10200, A=>nx10462);
   ix10201 : inv02 port map ( Y=>nx10202, A=>nx10462);
   ix10203 : inv02 port map ( Y=>nx10204, A=>nx10462);
   ix10205 : inv02 port map ( Y=>nx10206, A=>nx10462);
   ix10207 : inv02 port map ( Y=>nx10208, A=>nx10464);
   ix10209 : inv02 port map ( Y=>nx10210, A=>nx10464);
   ix10211 : inv02 port map ( Y=>nx10212, A=>nx10464);
   ix10213 : inv02 port map ( Y=>nx10214, A=>nx10464);
   ix10215 : inv02 port map ( Y=>nx10216, A=>nx10464);
   ix10219 : inv02 port map ( Y=>nx10220, A=>nx10466);
   ix10221 : inv02 port map ( Y=>nx10222, A=>nx10466);
   ix10223 : inv02 port map ( Y=>nx10224, A=>nx10466);
   ix10225 : inv02 port map ( Y=>nx10226, A=>nx10466);
   ix10227 : inv02 port map ( Y=>nx10228, A=>nx10466);
   ix10229 : inv02 port map ( Y=>nx10230, A=>nx10466);
   ix10231 : inv02 port map ( Y=>nx10232, A=>nx10466);
   ix10233 : inv02 port map ( Y=>nx10234, A=>nx10468);
   ix10235 : inv02 port map ( Y=>nx10236, A=>nx10468);
   ix10237 : inv02 port map ( Y=>nx10238, A=>nx10468);
   ix10239 : inv02 port map ( Y=>nx10240, A=>nx10468);
   ix10241 : inv02 port map ( Y=>nx10242, A=>nx10468);
   ix10245 : inv02 port map ( Y=>nx10246, A=>nx10470);
   ix10247 : inv02 port map ( Y=>nx10248, A=>nx10470);
   ix10249 : inv02 port map ( Y=>nx10250, A=>nx10470);
   ix10251 : inv02 port map ( Y=>nx10252, A=>nx10470);
   ix10253 : inv02 port map ( Y=>nx10254, A=>nx10470);
   ix10255 : inv02 port map ( Y=>nx10256, A=>nx10470);
   ix10257 : inv02 port map ( Y=>nx10258, A=>nx10470);
   ix10259 : inv02 port map ( Y=>nx10260, A=>nx10472);
   ix10261 : inv02 port map ( Y=>nx10262, A=>nx10472);
   ix10263 : inv02 port map ( Y=>nx10264, A=>nx10472);
   ix10265 : inv02 port map ( Y=>nx10266, A=>nx10472);
   ix10267 : inv02 port map ( Y=>nx10268, A=>nx10472);
   ix10271 : inv02 port map ( Y=>nx10272, A=>nx10474);
   ix10273 : inv02 port map ( Y=>nx10274, A=>nx10474);
   ix10275 : inv02 port map ( Y=>nx10276, A=>nx10474);
   ix10277 : inv02 port map ( Y=>nx10278, A=>nx10474);
   ix10279 : inv02 port map ( Y=>nx10280, A=>nx10474);
   ix10281 : inv02 port map ( Y=>nx10282, A=>nx10474);
   ix10283 : inv02 port map ( Y=>nx10284, A=>nx10474);
   ix10285 : inv02 port map ( Y=>nx10286, A=>nx10476);
   ix10287 : inv02 port map ( Y=>nx10288, A=>nx10476);
   ix10289 : inv02 port map ( Y=>nx10290, A=>nx10476);
   ix10291 : inv02 port map ( Y=>nx10292, A=>nx10476);
   ix10293 : inv02 port map ( Y=>nx10294, A=>nx10476);
   ix10297 : inv02 port map ( Y=>nx10298, A=>nx10478);
   ix10299 : inv02 port map ( Y=>nx10300, A=>nx10478);
   ix10301 : inv02 port map ( Y=>nx10302, A=>nx10478);
   ix10303 : inv02 port map ( Y=>nx10304, A=>nx10478);
   ix10305 : inv02 port map ( Y=>nx10306, A=>nx10478);
   ix10307 : inv02 port map ( Y=>nx10308, A=>nx10478);
   ix10309 : inv02 port map ( Y=>nx10310, A=>nx10478);
   ix10311 : inv02 port map ( Y=>nx10312, A=>nx10480);
   ix10313 : inv02 port map ( Y=>nx10314, A=>nx10480);
   ix10315 : inv02 port map ( Y=>nx10316, A=>nx10480);
   ix10317 : inv02 port map ( Y=>nx10318, A=>nx10480);
   ix10319 : inv02 port map ( Y=>nx10320, A=>nx10480);
   ix10323 : inv02 port map ( Y=>nx10324, A=>nx10482);
   ix10325 : inv02 port map ( Y=>nx10326, A=>nx10482);
   ix10327 : inv02 port map ( Y=>nx10328, A=>nx10482);
   ix10329 : inv02 port map ( Y=>nx10330, A=>nx10482);
   ix10331 : inv02 port map ( Y=>nx10332, A=>nx10482);
   ix10333 : inv02 port map ( Y=>nx10334, A=>nx10482);
   ix10335 : inv02 port map ( Y=>nx10336, A=>nx10482);
   ix10337 : inv02 port map ( Y=>nx10338, A=>nx10484);
   ix10339 : inv02 port map ( Y=>nx10340, A=>nx10484);
   ix10341 : inv02 port map ( Y=>nx10342, A=>nx10484);
   ix10343 : inv02 port map ( Y=>nx10344, A=>nx10484);
   ix10345 : inv02 port map ( Y=>nx10346, A=>nx10484);
   ix10349 : inv02 port map ( Y=>nx10350, A=>nx10486);
   ix10351 : inv02 port map ( Y=>nx10352, A=>nx10486);
   ix10353 : inv02 port map ( Y=>nx10354, A=>nx10486);
   ix10355 : inv02 port map ( Y=>nx10356, A=>nx10486);
   ix10357 : inv02 port map ( Y=>nx10358, A=>nx10486);
   ix10359 : inv02 port map ( Y=>nx10360, A=>nx10486);
   ix10361 : inv02 port map ( Y=>nx10362, A=>nx10486);
   ix10363 : inv02 port map ( Y=>nx10364, A=>nx10488);
   ix10365 : inv02 port map ( Y=>nx10366, A=>nx10488);
   ix10367 : inv02 port map ( Y=>nx10368, A=>nx10488);
   ix10369 : inv02 port map ( Y=>nx10370, A=>nx10488);
   ix10371 : inv02 port map ( Y=>nx10372, A=>nx10488);
   ix10373 : buf02 port map ( Y=>nx10374, A=>nx6955);
   ix10375 : buf02 port map ( Y=>nx10376, A=>nx6955);
   ix10377 : inv02 port map ( Y=>nx10378, A=>nx14);
   ix10379 : inv02 port map ( Y=>nx10380, A=>nx14);
   ix10381 : inv02 port map ( Y=>nx10382, A=>nx30);
   ix10383 : inv02 port map ( Y=>nx10384, A=>nx30);
   ix10385 : inv02 port map ( Y=>nx10386, A=>nx42);
   ix10387 : inv02 port map ( Y=>nx10388, A=>nx42);
   ix10389 : inv02 port map ( Y=>nx10390, A=>nx48);
   ix10391 : inv02 port map ( Y=>nx10392, A=>nx48);
   ix10393 : inv02 port map ( Y=>nx10394, A=>nx64);
   ix10395 : inv02 port map ( Y=>nx10396, A=>nx64);
   ix10397 : inv02 port map ( Y=>nx10398, A=>nx68);
   ix10399 : inv02 port map ( Y=>nx10400, A=>nx68);
   ix10401 : inv02 port map ( Y=>nx10402, A=>nx74);
   ix10403 : inv02 port map ( Y=>nx10404, A=>nx74);
   ix10405 : inv02 port map ( Y=>nx10406, A=>nx90);
   ix10407 : inv02 port map ( Y=>nx10408, A=>nx90);
   ix10409 : inv02 port map ( Y=>nx10410, A=>nx94);
   ix10411 : inv02 port map ( Y=>nx10412, A=>nx94);
   ix10413 : inv02 port map ( Y=>nx10414, A=>nx100);
   ix10415 : inv02 port map ( Y=>nx10416, A=>nx100);
   ix10417 : inv02 port map ( Y=>nx10418, A=>nx104);
   ix10419 : inv02 port map ( Y=>nx10420, A=>nx104);
   ix10421 : inv02 port map ( Y=>nx10422, A=>nx114);
   ix10423 : inv02 port map ( Y=>nx10424, A=>nx114);
   ix10425 : inv02 port map ( Y=>nx10426, A=>nx118);
   ix10427 : inv02 port map ( Y=>nx10428, A=>nx118);
   ix10429 : inv02 port map ( Y=>nx10430, A=>nx122);
   ix10431 : inv02 port map ( Y=>nx10432, A=>nx122);
   ix10433 : inv02 port map ( Y=>nx10434, A=>nx136);
   ix10435 : inv02 port map ( Y=>nx10436, A=>nx136);
   ix10437 : inv02 port map ( Y=>nx10438, A=>nx144);
   ix10439 : inv02 port map ( Y=>nx10440, A=>nx144);
   ix10441 : inv02 port map ( Y=>nx10442, A=>nx150);
   ix10443 : inv02 port map ( Y=>nx10444, A=>nx150);
   ix10445 : inv02 port map ( Y=>nx10446, A=>nx158);
   ix10447 : inv02 port map ( Y=>nx10448, A=>nx158);
   ix10449 : inv02 port map ( Y=>nx10450, A=>nx166);
   ix10451 : inv02 port map ( Y=>nx10452, A=>nx166);
   ix10453 : inv02 port map ( Y=>nx10454, A=>nx172);
   ix10455 : inv02 port map ( Y=>nx10456, A=>nx172);
   ix10457 : inv02 port map ( Y=>nx10458, A=>nx180);
   ix10459 : inv02 port map ( Y=>nx10460, A=>nx180);
   ix10461 : inv02 port map ( Y=>nx10462, A=>nx192);
   ix10463 : inv02 port map ( Y=>nx10464, A=>nx192);
   ix10465 : inv02 port map ( Y=>nx10466, A=>nx200);
   ix10467 : inv02 port map ( Y=>nx10468, A=>nx200);
   ix10469 : inv02 port map ( Y=>nx10470, A=>nx206);
   ix10471 : inv02 port map ( Y=>nx10472, A=>nx206);
   ix10473 : inv02 port map ( Y=>nx10474, A=>nx214);
   ix10475 : inv02 port map ( Y=>nx10476, A=>nx214);
   ix10477 : inv02 port map ( Y=>nx10478, A=>nx222);
   ix10479 : inv02 port map ( Y=>nx10480, A=>nx222);
   ix10481 : inv02 port map ( Y=>nx10482, A=>nx226);
   ix10483 : inv02 port map ( Y=>nx10484, A=>nx226);
   ix10485 : inv02 port map ( Y=>nx10486, A=>nx230);
   ix10487 : inv02 port map ( Y=>nx10488, A=>nx230);
   ix8951 : nor02ii port map ( Y=>sel_que_0, A0=>nx6829, A1=>nx6885);
   ix8961 : nor02ii port map ( Y=>sel_que_1, A0=>nx6839, A1=>nx6885);
   ix8971 : nor02ii port map ( Y=>sel_que_2, A0=>nx6843, A1=>nx6885);
   ix8979 : nor02ii port map ( Y=>sel_que_3, A0=>nx6847, A1=>nx6885);
   ix8987 : nor02ii port map ( Y=>sel_que_4, A0=>nx6829, A1=>nx6905);
   ix8991 : nor02ii port map ( Y=>sel_que_5, A0=>nx6839, A1=>nx6905);
   ix8995 : nor02ii port map ( Y=>sel_que_6, A0=>nx6843, A1=>nx6905);
   ix8999 : nor02ii port map ( Y=>sel_que_7, A0=>nx6847, A1=>nx6905);
   ix9007 : nor02ii port map ( Y=>sel_que_8, A0=>nx6829, A1=>nx6915);
   ix9011 : nor02ii port map ( Y=>sel_que_9, A0=>nx6839, A1=>nx6915);
   ix9015 : nor02ii port map ( Y=>sel_que_10, A0=>nx6843, A1=>nx6915);
   ix9019 : nor02ii port map ( Y=>sel_que_11, A0=>nx6847, A1=>nx6915);
   ix9053 : nor02ii port map ( Y=>sel_que_17, A0=>nx6893, A1=>nx6885);
   ix9063 : nor02ii port map ( Y=>sel_que_18, A0=>nx6897, A1=>nx6885);
   ix9071 : nor02ii port map ( Y=>sel_que_19, A0=>nx6901, A1=>nx6885);
   ix6906 : nor02ii port map ( Y=>nx6905, A0=>cache_in_sel(3), A1=>
      cache_in_sel(2));
   ix9079 : nor02ii port map ( Y=>sel_que_21, A0=>nx6893, A1=>nx6905);
   ix9083 : nor02ii port map ( Y=>sel_que_22, A0=>nx6897, A1=>nx6905);
   ix9087 : nor02ii port map ( Y=>sel_que_23, A0=>nx6901, A1=>nx6905);
   ix6916 : nor02ii port map ( Y=>nx6915, A0=>cache_in_sel(2), A1=>
      cache_in_sel(3));
   ix9095 : nor02ii port map ( Y=>sel_que_25, A0=>nx6893, A1=>nx6915);
   ix9099 : nor02ii port map ( Y=>sel_que_26, A0=>nx6897, A1=>nx6915);
   ix9103 : nor02ii port map ( Y=>sel_que_27, A0=>nx6901, A1=>nx6915);
   ix223 : nor02ii port map ( Y=>nx222, A0=>nx6931, A1=>nx62);
   ix231 : nor02ii port map ( Y=>nx230, A0=>nx6945, A1=>nx88);
   ix207 : nor02ii port map ( Y=>nx206, A0=>nx10374, A1=>nx28);
   ix123 : nor02ii port map ( Y=>nx122, A0=>nx10374, A1=>nx62);
   ix65 : nor02ii port map ( Y=>nx64, A0=>nx6949, A1=>nx62);
   ix49 : nor02ii port map ( Y=>nx48, A0=>nx6949, A1=>nx28);
   ix31 : nor02ii port map ( Y=>nx30, A0=>nx6931, A1=>nx28);
   ix10493 : inv02 port map ( Y=>nx10494, A=>nx6937);
   ix10495 : inv02 port map ( Y=>nx10496, A=>nx6937);
   ix10497 : inv02 port map ( Y=>nx10498, A=>nx6939);
   ix10499 : inv02 port map ( Y=>nx10500, A=>nx6939);
   ix10501 : inv01 port map ( Y=>nx10502, A=>nx6961);
   ix10503 : inv01 port map ( Y=>nx10504, A=>nx6961);
   ix10505 : inv02 port map ( Y=>nx10506, A=>nx6833);
   ix10507 : inv02 port map ( Y=>nx10508, A=>nx6835);
   ix10509 : inv01 port map ( Y=>nx10510, A=>in_word(15));
   ix10511 : inv01 port map ( Y=>nx10512, A=>nx10510);
   ix10513 : inv01 port map ( Y=>nx10514, A=>nx10510);
   ix10515 : inv01 port map ( Y=>nx10516, A=>nx10510);
   ix10517 : inv01 port map ( Y=>nx10518, A=>nx10510);
   ix10519 : inv01 port map ( Y=>nx10520, A=>in_word(14));
   ix10521 : inv01 port map ( Y=>nx10522, A=>nx10520);
   ix10523 : inv01 port map ( Y=>nx10524, A=>nx10520);
   ix10525 : inv01 port map ( Y=>nx10526, A=>nx10520);
   ix10527 : inv01 port map ( Y=>nx10528, A=>nx10520);
   ix10529 : inv01 port map ( Y=>nx10530, A=>in_word(13));
   ix10531 : inv01 port map ( Y=>nx10532, A=>nx10530);
   ix10533 : inv01 port map ( Y=>nx10534, A=>nx10530);
   ix10535 : inv01 port map ( Y=>nx10536, A=>nx10530);
   ix10537 : inv01 port map ( Y=>nx10538, A=>nx10530);
   ix10539 : inv01 port map ( Y=>nx10540, A=>in_word(12));
   ix10541 : inv01 port map ( Y=>nx10542, A=>nx10540);
   ix10543 : inv01 port map ( Y=>nx10544, A=>nx10540);
   ix10545 : inv01 port map ( Y=>nx10546, A=>nx10540);
   ix10547 : inv01 port map ( Y=>nx10548, A=>nx10540);
   ix10549 : inv01 port map ( Y=>nx10550, A=>in_word(11));
   ix10551 : inv01 port map ( Y=>nx10552, A=>nx10550);
   ix10553 : inv01 port map ( Y=>nx10554, A=>nx10550);
   ix10555 : inv01 port map ( Y=>nx10556, A=>nx10550);
   ix10557 : inv01 port map ( Y=>nx10558, A=>nx10550);
   ix10559 : inv01 port map ( Y=>nx10560, A=>in_word(10));
   ix10561 : inv01 port map ( Y=>nx10562, A=>nx10560);
   ix10563 : inv01 port map ( Y=>nx10564, A=>nx10560);
   ix10565 : inv01 port map ( Y=>nx10566, A=>nx10560);
   ix10567 : inv01 port map ( Y=>nx10568, A=>nx10560);
   ix10569 : inv01 port map ( Y=>nx10570, A=>in_word(9));
   ix10571 : inv01 port map ( Y=>nx10572, A=>nx10570);
   ix10573 : inv01 port map ( Y=>nx10574, A=>nx10570);
   ix10575 : inv01 port map ( Y=>nx10576, A=>nx10570);
   ix10577 : inv01 port map ( Y=>nx10578, A=>nx10570);
   ix10579 : inv01 port map ( Y=>nx10580, A=>in_word(8));
   ix10581 : inv01 port map ( Y=>nx10582, A=>nx10580);
   ix10583 : inv01 port map ( Y=>nx10584, A=>nx10580);
   ix10585 : inv01 port map ( Y=>nx10586, A=>nx10580);
   ix10587 : inv01 port map ( Y=>nx10588, A=>nx10580);
   ix10589 : inv01 port map ( Y=>nx10590, A=>in_word(7));
   ix10591 : inv01 port map ( Y=>nx10592, A=>nx10590);
   ix10593 : inv01 port map ( Y=>nx10594, A=>nx10590);
   ix10595 : inv01 port map ( Y=>nx10596, A=>nx10590);
   ix10597 : inv01 port map ( Y=>nx10598, A=>nx10590);
   ix10599 : inv01 port map ( Y=>nx10600, A=>in_word(6));
   ix10601 : inv01 port map ( Y=>nx10602, A=>nx10600);
   ix10603 : inv01 port map ( Y=>nx10604, A=>nx10600);
   ix10605 : inv01 port map ( Y=>nx10606, A=>nx10600);
   ix10607 : inv01 port map ( Y=>nx10608, A=>nx10600);
   ix10609 : inv01 port map ( Y=>nx10610, A=>in_word(5));
   ix10611 : inv01 port map ( Y=>nx10612, A=>nx10610);
   ix10613 : inv01 port map ( Y=>nx10614, A=>nx10610);
   ix10615 : inv01 port map ( Y=>nx10616, A=>nx10610);
   ix10617 : inv01 port map ( Y=>nx10618, A=>nx10610);
   ix10619 : inv01 port map ( Y=>nx10620, A=>in_word(4));
   ix10621 : inv01 port map ( Y=>nx10622, A=>nx10620);
   ix10623 : inv01 port map ( Y=>nx10624, A=>nx10620);
   ix10625 : inv01 port map ( Y=>nx10626, A=>nx10620);
   ix10627 : inv01 port map ( Y=>nx10628, A=>nx10620);
   ix10629 : inv01 port map ( Y=>nx10630, A=>in_word(3));
   ix10631 : inv01 port map ( Y=>nx10632, A=>nx10630);
   ix10633 : inv01 port map ( Y=>nx10634, A=>nx10630);
   ix10635 : inv01 port map ( Y=>nx10636, A=>nx10630);
   ix10637 : inv01 port map ( Y=>nx10638, A=>nx10630);
   ix10639 : inv01 port map ( Y=>nx10640, A=>in_word(2));
   ix10641 : inv01 port map ( Y=>nx10642, A=>nx10640);
   ix10643 : inv01 port map ( Y=>nx10644, A=>nx10640);
   ix10645 : inv01 port map ( Y=>nx10646, A=>nx10640);
   ix10647 : inv01 port map ( Y=>nx10648, A=>nx10640);
   ix10649 : inv01 port map ( Y=>nx10650, A=>in_word(1));
   ix10651 : inv01 port map ( Y=>nx10652, A=>nx10650);
   ix10653 : inv01 port map ( Y=>nx10654, A=>nx10650);
   ix10655 : inv01 port map ( Y=>nx10656, A=>nx10650);
   ix10657 : inv01 port map ( Y=>nx10658, A=>nx10650);
   ix10659 : inv01 port map ( Y=>nx10660, A=>in_word(0));
   ix10661 : inv01 port map ( Y=>nx10662, A=>nx10660);
   ix10663 : inv01 port map ( Y=>nx10664, A=>nx10660);
   ix10665 : inv01 port map ( Y=>nx10666, A=>nx10660);
   ix10667 : inv01 port map ( Y=>nx10668, A=>nx10660);
   ix10689 : inv02 port map ( Y=>nx10690, A=>nx10742);
   ix10691 : inv02 port map ( Y=>nx10692, A=>nx10742);
   ix10693 : inv02 port map ( Y=>nx10694, A=>nx10742);
   ix10695 : inv02 port map ( Y=>nx10696, A=>nx10742);
   ix10697 : inv02 port map ( Y=>nx10698, A=>nx10742);
   ix10699 : inv02 port map ( Y=>nx10700, A=>nx10742);
   ix10701 : inv02 port map ( Y=>nx10702, A=>nx10742);
   ix10703 : inv02 port map ( Y=>nx10704, A=>nx10744);
   ix10705 : inv02 port map ( Y=>nx10706, A=>nx10744);
   ix10707 : inv02 port map ( Y=>nx10708, A=>nx10744);
   ix10709 : inv02 port map ( Y=>nx10710, A=>nx10744);
   ix10711 : inv02 port map ( Y=>nx10712, A=>nx10744);
   ix10713 : inv02 port map ( Y=>nx10714, A=>nx10746);
   ix10715 : inv02 port map ( Y=>nx10716, A=>nx10746);
   ix10717 : inv02 port map ( Y=>nx10718, A=>nx10746);
   ix10719 : inv02 port map ( Y=>nx10720, A=>nx10746);
   ix10721 : inv02 port map ( Y=>nx10722, A=>nx10746);
   ix10723 : inv02 port map ( Y=>nx10724, A=>nx10746);
   ix10725 : inv02 port map ( Y=>nx10726, A=>nx10746);
   ix10727 : inv02 port map ( Y=>nx10728, A=>nx10748);
   ix10729 : inv02 port map ( Y=>nx10730, A=>nx10748);
   ix10731 : inv02 port map ( Y=>nx10732, A=>nx10748);
   ix10733 : inv02 port map ( Y=>nx10734, A=>nx10748);
   ix10735 : inv02 port map ( Y=>nx10736, A=>nx10748);
   ix10741 : inv02 port map ( Y=>nx10742, A=>reset);
   ix10743 : inv02 port map ( Y=>nx10744, A=>reset);
   ix10745 : inv02 port map ( Y=>nx10746, A=>clk);
   ix10747 : inv02 port map ( Y=>nx10748, A=>clk);
end Dataflow ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity AdvancedCounter_16 is
   port (
      clk : IN std_logic ;
      reset : IN std_logic ;
      enable : IN std_logic ;
      mode_in : IN std_logic_vector (1 DOWNTO 0) ;
      max_val_in : IN std_logic_vector (15 DOWNTO 0) ;
      max_reached_out : OUT std_logic ;
      counter_out : OUT std_logic_vector (15 DOWNTO 0)) ;
end AdvancedCounter_16 ;

architecture behavioural_unfold_2902 of AdvancedCounter_16 is
   signal counter_out_0_EXMPLR, counter_out_15_EXMPLR, counter_out_14_EXMPLR, 
      nx149, counter_out_13_EXMPLR, counter_out_12_EXMPLR, nx152, 
      counter_out_11_EXMPLR, counter_out_10_EXMPLR, nx155, 
      counter_out_9_EXMPLR, counter_out_8_EXMPLR, nx157, 
      counter_out_7_EXMPLR, counter_out_6_EXMPLR, nx159, 
      counter_out_5_EXMPLR, counter_out_4_EXMPLR, nx161, 
      counter_out_3_EXMPLR, counter_out_2_EXMPLR, counter_out_1_EXMPLR, 
      counter_out_dup0_0, nx22, nx34, nx46, nx70, nx94, nx118, nx142, nx166, 
      nx174, nx192, nx206, nx224, nx246, nx173, nx183, nx193, nx203, nx213, 
      nx223, nx233, nx243, nx253, nx263, nx273, nx283, nx293, nx303, nx313, 
      nx323, nx339, nx344, nx348, nx350, nx353, nx358, nx362, nx364, nx367, 
      nx372, nx376, nx378, nx381, nx386, nx390, nx392, nx395, nx400, nx404, 
      nx406, nx409, nx414, nx419, nx424, nx428, nx430, nx436, nx439, nx445, 
      nx447, nx449, nx451, nx458, nx460, nx462, nx464, nx466, nx468, nx470, 
      nx472, nx474: std_logic ;

begin
   counter_out(15) <= counter_out_0_EXMPLR ;
   counter_out(14) <= counter_out_0_EXMPLR ;
   counter_out(13) <= counter_out_0_EXMPLR ;
   counter_out(12) <= counter_out_0_EXMPLR ;
   counter_out(11) <= counter_out_0_EXMPLR ;
   counter_out(10) <= counter_out_0_EXMPLR ;
   counter_out(9) <= counter_out_0_EXMPLR ;
   counter_out(8) <= counter_out_0_EXMPLR ;
   counter_out(7) <= counter_out_0_EXMPLR ;
   counter_out(6) <= counter_out_0_EXMPLR ;
   counter_out(5) <= counter_out_0_EXMPLR ;
   counter_out(4) <= counter_out_0_EXMPLR ;
   counter_out(3) <= counter_out_0_EXMPLR ;
   counter_out(2) <= counter_out_0_EXMPLR ;
   counter_out(1) <= counter_out_0_EXMPLR ;
   counter_out(0) <= counter_out_0_EXMPLR ;
   ix140 : fake_gnd port map ( Y=>counter_out_0_EXMPLR);
   ix251 : and04 port map ( Y=>max_reached_out, A0=>nx192, A1=>nx206, A2=>
      nx224, A3=>nx246);
   ix324 : mux21_ni port map ( Y=>nx323, A0=>counter_out_15_EXMPLR, A1=>
      nx174, S0=>nx474);
   ix314 : mux21_ni port map ( Y=>nx313, A0=>counter_out_14_EXMPLR, A1=>
      nx166, S0=>nx472);
   reg_counter_data_14 : dffr port map ( Q=>counter_out_14_EXMPLR, QB=>nx339, 
      D=>nx313, CLK=>clk, R=>nx462);
   ix345 : nand02 port map ( Y=>nx344, A0=>counter_out_13_EXMPLR, A1=>nx152
   );
   ix304 : mux21 port map ( Y=>nx303, A0=>nx348, A1=>nx350, S0=>nx472);
   reg_counter_data_13 : dffr port map ( Q=>counter_out_13_EXMPLR, QB=>nx348, 
      D=>nx303, CLK=>clk, R=>nx462);
   ix351 : oai21 port map ( Y=>nx350, A0=>nx152, A1=>counter_out_13_EXMPLR, 
      B0=>nx344);
   ix294 : mux21_ni port map ( Y=>nx293, A0=>counter_out_12_EXMPLR, A1=>
      nx142, S0=>nx472);
   reg_counter_data_12 : dffr port map ( Q=>counter_out_12_EXMPLR, QB=>nx353, 
      D=>nx293, CLK=>clk, R=>nx462);
   ix359 : nand02 port map ( Y=>nx358, A0=>counter_out_11_EXMPLR, A1=>nx155
   );
   ix284 : mux21 port map ( Y=>nx283, A0=>nx362, A1=>nx364, S0=>nx472);
   reg_counter_data_11 : dffr port map ( Q=>counter_out_11_EXMPLR, QB=>nx362, 
      D=>nx283, CLK=>clk, R=>nx462);
   ix365 : oai21 port map ( Y=>nx364, A0=>nx155, A1=>counter_out_11_EXMPLR, 
      B0=>nx358);
   ix274 : mux21_ni port map ( Y=>nx273, A0=>counter_out_10_EXMPLR, A1=>
      nx118, S0=>nx472);
   reg_counter_data_10 : dffr port map ( Q=>counter_out_10_EXMPLR, QB=>nx367, 
      D=>nx273, CLK=>clk, R=>nx462);
   ix373 : nand02 port map ( Y=>nx372, A0=>counter_out_9_EXMPLR, A1=>nx157);
   ix264 : mux21 port map ( Y=>nx263, A0=>nx376, A1=>nx378, S0=>nx472);
   reg_counter_data_9 : dffr port map ( Q=>counter_out_9_EXMPLR, QB=>nx376, 
      D=>nx263, CLK=>clk, R=>nx462);
   ix379 : oai21 port map ( Y=>nx378, A0=>nx157, A1=>counter_out_9_EXMPLR, 
      B0=>nx372);
   ix254 : mux21_ni port map ( Y=>nx253, A0=>counter_out_8_EXMPLR, A1=>nx94, 
      S0=>nx472);
   reg_counter_data_8 : dffr port map ( Q=>counter_out_8_EXMPLR, QB=>nx381, 
      D=>nx253, CLK=>clk, R=>nx462);
   ix387 : nand02 port map ( Y=>nx386, A0=>counter_out_7_EXMPLR, A1=>nx159);
   ix244 : mux21 port map ( Y=>nx243, A0=>nx390, A1=>nx392, S0=>nx470);
   reg_counter_data_7 : dffr port map ( Q=>counter_out_7_EXMPLR, QB=>nx390, 
      D=>nx243, CLK=>clk, R=>nx464);
   ix393 : oai21 port map ( Y=>nx392, A0=>nx159, A1=>counter_out_7_EXMPLR, 
      B0=>nx386);
   ix234 : mux21_ni port map ( Y=>nx233, A0=>counter_out_6_EXMPLR, A1=>nx70, 
      S0=>nx470);
   reg_counter_data_6 : dffr port map ( Q=>counter_out_6_EXMPLR, QB=>nx395, 
      D=>nx233, CLK=>clk, R=>nx464);
   ix401 : nand02 port map ( Y=>nx400, A0=>counter_out_5_EXMPLR, A1=>nx161);
   ix224 : mux21 port map ( Y=>nx223, A0=>nx404, A1=>nx406, S0=>nx470);
   reg_counter_data_5 : dffr port map ( Q=>counter_out_5_EXMPLR, QB=>nx404, 
      D=>nx223, CLK=>clk, R=>nx464);
   ix407 : oai21 port map ( Y=>nx406, A0=>nx161, A1=>counter_out_5_EXMPLR, 
      B0=>nx400);
   ix214 : mux21_ni port map ( Y=>nx213, A0=>counter_out_4_EXMPLR, A1=>nx46, 
      S0=>nx470);
   reg_counter_data_4 : dffr port map ( Q=>counter_out_4_EXMPLR, QB=>nx409, 
      D=>nx213, CLK=>clk, R=>nx464);
   ix47 : aoi21 port map ( Y=>nx46, A0=>nx414, A1=>nx409, B0=>nx161);
   ix415 : nand04 port map ( Y=>nx414, A0=>counter_out_3_EXMPLR, A1=>
      counter_out_2_EXMPLR, A2=>counter_out_1_EXMPLR, A3=>counter_out_dup0_0
   );
   reg_counter_data_3 : dffr port map ( Q=>counter_out_3_EXMPLR, QB=>OPEN, D
      =>nx203, CLK=>clk, R=>nx466);
   ix204 : mux21_ni port map ( Y=>nx203, A0=>counter_out_3_EXMPLR, A1=>nx34, 
      S0=>nx470);
   ix35 : xnor2 port map ( Y=>nx34, A0=>counter_out_3_EXMPLR, A1=>nx419);
   ix420 : nand03 port map ( Y=>nx419, A0=>counter_out_2_EXMPLR, A1=>
      counter_out_1_EXMPLR, A2=>counter_out_dup0_0);
   reg_counter_data_2 : dffr port map ( Q=>counter_out_2_EXMPLR, QB=>OPEN, D
      =>nx193, CLK=>clk, R=>nx464);
   ix194 : mux21_ni port map ( Y=>nx193, A0=>counter_out_2_EXMPLR, A1=>nx22, 
      S0=>nx470);
   ix23 : xnor2 port map ( Y=>nx22, A0=>counter_out_2_EXMPLR, A1=>nx424);
   ix184 : mux21 port map ( Y=>nx183, A0=>nx428, A1=>nx430, S0=>nx470);
   reg_counter_data_1 : dffr port map ( Q=>counter_out_1_EXMPLR, QB=>nx428, 
      D=>nx183, CLK=>clk, R=>nx464);
   ix431 : oai21 port map ( Y=>nx430, A0=>counter_out_dup0_0, A1=>
      counter_out_1_EXMPLR, B0=>nx424);
   reg_counter_data_0 : dffr port map ( Q=>counter_out_dup0_0, QB=>nx436, D
      =>nx173, CLK=>clk, R=>nx464);
   reg_counter_data_15 : dffr port map ( Q=>counter_out_15_EXMPLR, QB=>nx439, 
      D=>nx323, CLK=>clk, R=>nx466);
   ix247 : and04 port map ( Y=>nx246, A0=>nx445, A1=>nx447, A2=>nx449, A3=>
      nx451);
   ix448 : xnor2 port map ( Y=>nx447, A0=>counter_out_2_EXMPLR, A1=>
      max_val_in(2));
   ix450 : xnor2 port map ( Y=>nx449, A0=>counter_out_3_EXMPLR, A1=>
      max_val_in(3));
   ix193 : and04 port map ( Y=>nx192, A0=>nx439, A1=>nx339, A2=>nx348, A3=>
      nx353);
   ix175 : xor2 port map ( Y=>nx174, A0=>nx149, A1=>counter_out_15_EXMPLR);
   ix173 : nor02ii port map ( Y=>nx149, A0=>nx344, A1=>counter_out_14_EXMPLR
   );
   ix167 : xor2 port map ( Y=>nx166, A0=>nx339, A1=>nx344);
   ix149 : nor02ii port map ( Y=>nx152, A0=>nx358, A1=>counter_out_12_EXMPLR
   );
   ix143 : xor2 port map ( Y=>nx142, A0=>nx353, A1=>nx358);
   ix125 : nor02ii port map ( Y=>nx155, A0=>nx372, A1=>counter_out_10_EXMPLR
   );
   ix119 : xor2 port map ( Y=>nx118, A0=>nx367, A1=>nx372);
   ix101 : nor02ii port map ( Y=>nx157, A0=>nx386, A1=>counter_out_8_EXMPLR
   );
   ix95 : xor2 port map ( Y=>nx94, A0=>nx381, A1=>nx386);
   ix77 : nor02ii port map ( Y=>nx159, A0=>nx400, A1=>counter_out_6_EXMPLR);
   ix71 : xor2 port map ( Y=>nx70, A0=>nx395, A1=>nx400);
   ix53 : nor02ii port map ( Y=>nx161, A0=>nx414, A1=>counter_out_4_EXMPLR);
   ix425 : or02 port map ( Y=>nx424, A0=>nx428, A1=>nx436);
   ix174 : xnor2 port map ( Y=>nx173, A0=>nx436, A1=>nx474);
   ix207 : and04 port map ( Y=>nx206, A0=>nx362, A1=>nx367, A2=>nx376, A3=>
      nx381);
   ix225 : and04 port map ( Y=>nx224, A0=>nx390, A1=>nx395, A2=>nx404, A3=>
      nx458);
   ix217 : xnor2 port map ( Y=>nx458, A0=>max_val_in(0), A1=>
      counter_out_dup0_0);
   ix446 : xor2 port map ( Y=>nx445, A0=>nx428, A1=>max_val_in(1));
   ix452 : xor2 port map ( Y=>nx451, A0=>nx409, A1=>max_val_in(4));
   ix459 : inv01 port map ( Y=>nx460, A=>reset);
   ix461 : inv02 port map ( Y=>nx462, A=>nx460);
   ix463 : inv02 port map ( Y=>nx464, A=>nx460);
   ix465 : inv02 port map ( Y=>nx466, A=>nx460);
   ix467 : inv01 port map ( Y=>nx468, A=>enable);
   ix469 : inv02 port map ( Y=>nx470, A=>nx468);
   ix471 : inv02 port map ( Y=>nx472, A=>nx468);
   ix473 : inv02 port map ( Y=>nx474, A=>nx468);
end behavioural_unfold_2902 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Controller_16_16_5_16 is
   port (
      clk : IN std_logic ;
      reset : IN std_logic ;
      io_ready_in : IN std_logic ;
      io_done_out : OUT std_logic ;
      mem_data_in : IN std_logic_vector (15 DOWNTO 0) ;
      mem_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
      mem_addr_out : OUT std_logic_vector (15 DOWNTO 0) ;
      mem_write_out : OUT std_logic ;
      mem_read_out : OUT std_logic ;
      wind_en : OUT std_logic ;
      wind_rst : OUT std_logic ;
      wind_col_in_4_15 : OUT std_logic ;
      wind_col_in_4_14 : OUT std_logic ;
      wind_col_in_4_13 : OUT std_logic ;
      wind_col_in_4_12 : OUT std_logic ;
      wind_col_in_4_11 : OUT std_logic ;
      wind_col_in_4_10 : OUT std_logic ;
      wind_col_in_4_9 : OUT std_logic ;
      wind_col_in_4_8 : OUT std_logic ;
      wind_col_in_4_7 : OUT std_logic ;
      wind_col_in_4_6 : OUT std_logic ;
      wind_col_in_4_5 : OUT std_logic ;
      wind_col_in_4_4 : OUT std_logic ;
      wind_col_in_4_3 : OUT std_logic ;
      wind_col_in_4_2 : OUT std_logic ;
      wind_col_in_4_1 : OUT std_logic ;
      wind_col_in_4_0 : OUT std_logic ;
      wind_col_in_3_15 : OUT std_logic ;
      wind_col_in_3_14 : OUT std_logic ;
      wind_col_in_3_13 : OUT std_logic ;
      wind_col_in_3_12 : OUT std_logic ;
      wind_col_in_3_11 : OUT std_logic ;
      wind_col_in_3_10 : OUT std_logic ;
      wind_col_in_3_9 : OUT std_logic ;
      wind_col_in_3_8 : OUT std_logic ;
      wind_col_in_3_7 : OUT std_logic ;
      wind_col_in_3_6 : OUT std_logic ;
      wind_col_in_3_5 : OUT std_logic ;
      wind_col_in_3_4 : OUT std_logic ;
      wind_col_in_3_3 : OUT std_logic ;
      wind_col_in_3_2 : OUT std_logic ;
      wind_col_in_3_1 : OUT std_logic ;
      wind_col_in_3_0 : OUT std_logic ;
      wind_col_in_2_15 : OUT std_logic ;
      wind_col_in_2_14 : OUT std_logic ;
      wind_col_in_2_13 : OUT std_logic ;
      wind_col_in_2_12 : OUT std_logic ;
      wind_col_in_2_11 : OUT std_logic ;
      wind_col_in_2_10 : OUT std_logic ;
      wind_col_in_2_9 : OUT std_logic ;
      wind_col_in_2_8 : OUT std_logic ;
      wind_col_in_2_7 : OUT std_logic ;
      wind_col_in_2_6 : OUT std_logic ;
      wind_col_in_2_5 : OUT std_logic ;
      wind_col_in_2_4 : OUT std_logic ;
      wind_col_in_2_3 : OUT std_logic ;
      wind_col_in_2_2 : OUT std_logic ;
      wind_col_in_2_1 : OUT std_logic ;
      wind_col_in_2_0 : OUT std_logic ;
      wind_col_in_1_15 : OUT std_logic ;
      wind_col_in_1_14 : OUT std_logic ;
      wind_col_in_1_13 : OUT std_logic ;
      wind_col_in_1_12 : OUT std_logic ;
      wind_col_in_1_11 : OUT std_logic ;
      wind_col_in_1_10 : OUT std_logic ;
      wind_col_in_1_9 : OUT std_logic ;
      wind_col_in_1_8 : OUT std_logic ;
      wind_col_in_1_7 : OUT std_logic ;
      wind_col_in_1_6 : OUT std_logic ;
      wind_col_in_1_5 : OUT std_logic ;
      wind_col_in_1_4 : OUT std_logic ;
      wind_col_in_1_3 : OUT std_logic ;
      wind_col_in_1_2 : OUT std_logic ;
      wind_col_in_1_1 : OUT std_logic ;
      wind_col_in_1_0 : OUT std_logic ;
      wind_col_in_0_15 : OUT std_logic ;
      wind_col_in_0_14 : OUT std_logic ;
      wind_col_in_0_13 : OUT std_logic ;
      wind_col_in_0_12 : OUT std_logic ;
      wind_col_in_0_11 : OUT std_logic ;
      wind_col_in_0_10 : OUT std_logic ;
      wind_col_in_0_9 : OUT std_logic ;
      wind_col_in_0_8 : OUT std_logic ;
      wind_col_in_0_7 : OUT std_logic ;
      wind_col_in_0_6 : OUT std_logic ;
      wind_col_in_0_5 : OUT std_logic ;
      wind_col_in_0_4 : OUT std_logic ;
      wind_col_in_0_3 : OUT std_logic ;
      wind_col_in_0_2 : OUT std_logic ;
      wind_col_in_0_1 : OUT std_logic ;
      wind_col_in_0_0 : OUT std_logic ;
      filter_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
      filter_ready_out : OUT std_logic ;
      filter_reset : OUT std_logic ;
      comp_unit_ready : OUT std_logic ;
      comp_unit_operation : OUT std_logic ;
      comp_unit_flt_size : OUT std_logic ;
      comp_unit_relu : OUT std_logic ;
      comp_unit_data1_out : OUT std_logic_vector (15 DOWNTO 0) ;
      comp_unit_data2_out : OUT std_logic_vector (15 DOWNTO 0) ;
      comp_unit_buffer_finished : IN std_logic ;
      comp_unit_finished : IN std_logic ;
      comp_unit_data1_in : IN std_logic_vector (15 DOWNTO 0) ;
      comp_unit_data2_in : IN std_logic_vector (15 DOWNTO 0) ;
      argmax_ready : OUT std_logic ;
      argmax_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
      argmax_data_in : IN std_logic_vector (15 DOWNTO 0)) ;
end Controller_16_16_5_16 ;

architecture Mixed_unfold_2045 of Controller_16_16_5_16 is
   component Cache_5_16_28_5
      port (
         in_word : IN std_logic_vector (15 DOWNTO 0) ;
         cache_in_sel : IN std_logic_vector (4 DOWNTO 0) ;
         cache_out_sel : IN std_logic_vector (4 DOWNTO 0) ;
         decoder_enable : IN std_logic ;
         out_column_0_15 : OUT std_logic ;
         out_column_0_14 : OUT std_logic ;
         out_column_0_13 : OUT std_logic ;
         out_column_0_12 : OUT std_logic ;
         out_column_0_11 : OUT std_logic ;
         out_column_0_10 : OUT std_logic ;
         out_column_0_9 : OUT std_logic ;
         out_column_0_8 : OUT std_logic ;
         out_column_0_7 : OUT std_logic ;
         out_column_0_6 : OUT std_logic ;
         out_column_0_5 : OUT std_logic ;
         out_column_0_4 : OUT std_logic ;
         out_column_0_3 : OUT std_logic ;
         out_column_0_2 : OUT std_logic ;
         out_column_0_1 : OUT std_logic ;
         out_column_0_0 : OUT std_logic ;
         out_column_1_15 : OUT std_logic ;
         out_column_1_14 : OUT std_logic ;
         out_column_1_13 : OUT std_logic ;
         out_column_1_12 : OUT std_logic ;
         out_column_1_11 : OUT std_logic ;
         out_column_1_10 : OUT std_logic ;
         out_column_1_9 : OUT std_logic ;
         out_column_1_8 : OUT std_logic ;
         out_column_1_7 : OUT std_logic ;
         out_column_1_6 : OUT std_logic ;
         out_column_1_5 : OUT std_logic ;
         out_column_1_4 : OUT std_logic ;
         out_column_1_3 : OUT std_logic ;
         out_column_1_2 : OUT std_logic ;
         out_column_1_1 : OUT std_logic ;
         out_column_1_0 : OUT std_logic ;
         out_column_2_15 : OUT std_logic ;
         out_column_2_14 : OUT std_logic ;
         out_column_2_13 : OUT std_logic ;
         out_column_2_12 : OUT std_logic ;
         out_column_2_11 : OUT std_logic ;
         out_column_2_10 : OUT std_logic ;
         out_column_2_9 : OUT std_logic ;
         out_column_2_8 : OUT std_logic ;
         out_column_2_7 : OUT std_logic ;
         out_column_2_6 : OUT std_logic ;
         out_column_2_5 : OUT std_logic ;
         out_column_2_4 : OUT std_logic ;
         out_column_2_3 : OUT std_logic ;
         out_column_2_2 : OUT std_logic ;
         out_column_2_1 : OUT std_logic ;
         out_column_2_0 : OUT std_logic ;
         out_column_3_15 : OUT std_logic ;
         out_column_3_14 : OUT std_logic ;
         out_column_3_13 : OUT std_logic ;
         out_column_3_12 : OUT std_logic ;
         out_column_3_11 : OUT std_logic ;
         out_column_3_10 : OUT std_logic ;
         out_column_3_9 : OUT std_logic ;
         out_column_3_8 : OUT std_logic ;
         out_column_3_7 : OUT std_logic ;
         out_column_3_6 : OUT std_logic ;
         out_column_3_5 : OUT std_logic ;
         out_column_3_4 : OUT std_logic ;
         out_column_3_3 : OUT std_logic ;
         out_column_3_2 : OUT std_logic ;
         out_column_3_1 : OUT std_logic ;
         out_column_3_0 : OUT std_logic ;
         out_column_4_15 : OUT std_logic ;
         out_column_4_14 : OUT std_logic ;
         out_column_4_13 : OUT std_logic ;
         out_column_4_12 : OUT std_logic ;
         out_column_4_11 : OUT std_logic ;
         out_column_4_10 : OUT std_logic ;
         out_column_4_9 : OUT std_logic ;
         out_column_4_8 : OUT std_logic ;
         out_column_4_7 : OUT std_logic ;
         out_column_4_6 : OUT std_logic ;
         out_column_4_5 : OUT std_logic ;
         out_column_4_4 : OUT std_logic ;
         out_column_4_3 : OUT std_logic ;
         out_column_4_2 : OUT std_logic ;
         out_column_4_1 : OUT std_logic ;
         out_column_4_0 : OUT std_logic ;
         clk : IN std_logic ;
         reset : IN std_logic) ;
   end component ;
   component AdvancedCounter_16
      port (
         clk : IN std_logic ;
         reset : IN std_logic ;
         enable : IN std_logic ;
         mode_in : IN std_logic_vector (1 DOWNTO 0) ;
         max_val_in : IN std_logic_vector (15 DOWNTO 0) ;
         max_reached_out : OUT std_logic ;
         counter_out : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   signal current_state_13, wind_width_count_4, wind_width_count_3, 
      wind_width_count_2, wind_width_count_1, wind_width_count_0, 
      cache_height_count_en, cache_height_ended, max_height_2, max_height_0, 
      cache_width_count_4, cache_width_count_3, cache_width_count_2, 
      cache_width_count_1, cache_width_count_0, cache_data_in_15, 
      cache_data_in_14, cache_data_in_13, cache_data_in_12, cache_data_in_11, 
      cache_data_in_10, cache_data_in_9, cache_data_in_8, cache_data_in_7, 
      cache_data_in_6, cache_data_in_5, cache_data_in_4, cache_data_in_3, 
      cache_data_in_2, cache_data_in_1, cache_data_in_0, cache_data_out_4_15, 
      cache_data_out_4_14, cache_data_out_4_13, cache_data_out_4_12, 
      cache_data_out_4_11, cache_data_out_4_10, cache_data_out_4_9, 
      cache_data_out_4_8, cache_data_out_4_7, cache_data_out_4_6, 
      cache_data_out_4_5, cache_data_out_4_4, cache_data_out_4_3, 
      cache_data_out_4_2, cache_data_out_4_1, cache_data_out_4_0, 
      cache_data_out_3_15, cache_data_out_3_14, cache_data_out_3_13, 
      cache_data_out_3_12, cache_data_out_3_11, cache_data_out_3_10, 
      cache_data_out_3_9, cache_data_out_3_8, cache_data_out_3_7, 
      cache_data_out_3_6, cache_data_out_3_5, cache_data_out_3_4, 
      cache_data_out_3_3, cache_data_out_3_2, cache_data_out_3_1, 
      cache_data_out_3_0, cache_data_out_2_15, cache_data_out_2_14, 
      cache_data_out_2_13, cache_data_out_2_12, cache_data_out_2_11, 
      cache_data_out_2_10, cache_data_out_2_9, cache_data_out_2_8, 
      cache_data_out_2_7, cache_data_out_2_6, cache_data_out_2_5, 
      cache_data_out_2_4, cache_data_out_2_3, cache_data_out_2_2, 
      cache_data_out_2_1, cache_data_out_2_0, cache_data_out_1_15, 
      cache_data_out_1_14, cache_data_out_1_13, cache_data_out_1_12, 
      cache_data_out_1_11, cache_data_out_1_10, cache_data_out_1_9, 
      cache_data_out_1_8, cache_data_out_1_7, cache_data_out_1_6, 
      cache_data_out_1_5, cache_data_out_1_4, cache_data_out_1_3, 
      cache_data_out_1_2, cache_data_out_1_1, cache_data_out_1_0, 
      cache_data_out_0_15, cache_data_out_0_14, cache_data_out_0_13, 
      cache_data_out_0_12, cache_data_out_0_11, cache_data_out_0_10, 
      cache_data_out_0_9, cache_data_out_0_8, cache_data_out_0_7, 
      cache_data_out_0_6, cache_data_out_0_5, cache_data_out_0_4, 
      cache_data_out_0_3, cache_data_out_0_2, cache_data_out_0_1, 
      cache_data_out_0_0, cache_load, cache_rst_actual, max_height_4, 
      max_height_3, max_height_1, comp_unit_operation_EXMPLR, 
      filter_reset_EXMPLR, current_state_21, current_state_20, 
      layer_type_out_1, current_state_3, nx1409, current_state_24, 
      ftc_cntrl_reg_out_12, current_state_16, ftc_cntrl_reg_out_8, nx1411, 
      nx4, nx14, ftc_cntrl_reg_out_14, current_state_12, current_state_25, 
      nflt_layer_out_3, current_state_4, nflt_layer_out_1, nflt_layer_out_0, 
      nx98, nx1419, nx112, current_state_9, current_state_8, current_state_7, 
      current_state_6, current_state_5, nx136, nx146, nx1421, nx152, 
      cntr1_inst_counter_out_1, cntr1_inst_counter_out_0, nx176, 
      cntr1_inst_counter_out_3, cntr1_inst_counter_out_2, nx200, nx214, 
      cntr1_inst_counter_out_4, nx1425, nx232, nx246, nx248, flt_size_out_0, 
      flt_size_out_2, flt_size_out_1, nx278, nx280, nx286, nx300, nx1427, 
      nx306, ftc_cntrl_reg_out_13, nx320, nx332, ftc_cntrl_reg_out_11, 
      nx1429, window_width_cntr_counter_out_14, nx1430, 
      window_width_cntr_counter_out_13, window_width_cntr_counter_out_12, 
      nx1432, window_width_cntr_counter_out_11, 
      window_width_cntr_counter_out_10, nx1434, 
      window_width_cntr_counter_out_9, window_width_cntr_counter_out_8, 
      nx1436, window_width_cntr_counter_out_7, 
      window_width_cntr_counter_out_6, nx1439, 
      window_width_cntr_counter_out_5, nx348, nx354, nx362, nx370, nx378, 
      nx398, nx422, nx446, nx470, nx494, nx520, nx534, nx546, 
      img_width_out_0, new_width_out_0, nx572, nx574, nx582, img_width_out_1, 
      new_width_out_1, nx600, nx606, nx610, img_width_out_2, new_width_out_2, 
      nx644, img_width_out_3, new_width_out_3, nx674, img_width_out_4, 
      new_width_out_4, nx692, nx702, current_state_15, 
      write_offset_data_out_0, nx730, new_size_squared_out_0, 
      write_offset_data_out_1, nx750, new_size_squared_out_1, 
      write_offset_data_out_2, new_size_squared_out_2, 
      write_offset_data_out_3, nx802, new_size_squared_out_3, nx820, 
      write_offset_data_out_4, nx822, nx828, new_size_squared_out_4, 
      write_offset_data_out_5, new_size_squared_out_5, 
      write_offset_data_out_6, nx868, nx874, new_size_squared_out_6, 
      write_offset_data_out_7, new_size_squared_out_7, nx914, 
      write_offset_data_out_8, nx918, nx924, new_size_squared_out_8, 
      write_offset_data_out_9, new_size_squared_out_9, 
      write_offset_data_out_10, nx964, nx970, new_size_squared_out_10, 
      write_offset_data_out_11, new_size_squared_out_11, nx1010, 
      write_offset_data_out_12, nx1012, nx1018, new_size_squared_out_12, 
      write_offset_data_out_13, new_size_squared_out_13, 
      write_offset_data_out_14, nx1058, nx1064, new_size_squared_out_14, 
      write_offset_data_out_15, new_size_squared_out_15, nx1098, nx1108, 
      ftc_cntrl_reg_out_9, nx1116, nx1124, nx1138, ftc_cntrl_reg_out_10, 
      nx1152, nx1166, cache_width_cntr_counter_out_14, nx1447, 
      cache_width_cntr_counter_out_13, cache_width_cntr_counter_out_12, 
      nx1449, cache_width_cntr_counter_out_11, 
      cache_width_cntr_counter_out_10, nx1451, 
      cache_width_cntr_counter_out_9, cache_width_cntr_counter_out_8, nx1454, 
      cache_width_cntr_counter_out_7, cache_width_cntr_counter_out_6, nx1456, 
      nx1192, nx1198, nx1206, nx1214, nx1222, cache_width_cntr_counter_out_5, 
      nx1228, nx1248, nx1272, nx1296, nx1320, nx1344, nx1370, nx1384, nx1402, 
      nx1404, nx1406, nx1414, nx1416, nx1424, nx1428, current_state_19, 
      current_state_18, nx1446, nx1452, nx1468, nx1459, nx1486, nx1492, 
      nx1502, nx1461, nx1516, num_channels_out_3, nflt_layer_temp_3, nx1528, 
      nx1463, num_channels_out_2, nflt_layer_temp_2, nx1464, 
      num_channels_out_1, nflt_layer_temp_1, num_channels_out_0, 
      current_state_2, nx1572, nx1578, nflt_layer_temp_0, 
      max_num_channels_data_out_0, nx1594, nx1602, nx1610, nx1620, nx1630, 
      max_num_channels_data_out_1, nx1646, nx1652, nx1664, 
      max_num_channels_data_out_2, nx1678, nx1690, 
      max_num_channels_data_out_3, nx1704, nx1716, 
      max_num_channels_data_out_4, nlayers_counter_out_0, 
      nlayers_counter_out_2, nlayers_counter_out_1, nx1768, nx1784, nx1800, 
      nx1469, nx1842, nx1880, current_state_28, current_state_27, 
      class_cntr_counter_out_3, class_cntr_counter_out_2, 
      class_cntr_counter_out_1, class_cntr_counter_out_0, nx1908, nx1916, 
      nx1942, nx1950, flt_bias_out_0, nx2084, nx2096, nx2098, flt_bias_out_1, 
      nx2124, flt_bias_out_2, nx2150, flt_bias_out_3, nx2176, flt_bias_out_4, 
      nx2202, flt_bias_out_5, nx2228, flt_bias_out_6, nx2254, flt_bias_out_7, 
      nx2280, flt_bias_out_8, nx2306, flt_bias_out_9, nx2332, 
      flt_bias_out_10, nx2358, flt_bias_out_11, nx2384, flt_bias_out_12, 
      nx2410, flt_bias_out_13, nx2436, flt_bias_out_14, nx2462, 
      flt_bias_out_15, nx2488, nx2502, ftc_cntrl_reg_out_15, nx2522, nx2536, 
      nx2580, nx2582, bias_offset_data_out_0, nx2620, nx2626, 
      img_base_addr_0, write_base_prev_data_out_0, nx2636, nx2640, 
      img_addr_offset_0, nx2680, addr1_data_0, nx2706, write_base_data_out_1, 
      nx2752, nx2760, nx2766, addr1_data_1, bias_offset_data_out_1, nx2794, 
      nx2796, img_base_addr_1, write_base_prev_data_out_1, img_addr_offset_1, 
      nx2832, nx2834, write_base_data_out_2, nx2872, nx2882, nx2884, nx2886, 
      nx2894, addr1_data_2, nx2904, bias_offset_data_out_2, nx2932, 
      img_base_addr_2, write_base_prev_data_out_2, nx2950, nx2956, 
      img_addr_offset_2, nx2970, nx2978, write_base_data_out_3, nx3004, 
      nx3006, nx3016, nx3032, nx3034, addr1_data_3, nx3048, nx3066, 
      bias_offset_data_out_3, nx3074, nx3076, nx3086, img_base_addr_3, 
      write_base_prev_data_out_3, nx3100, img_addr_offset_3, nx3114, nx3120, 
      nx3122, nx3138, write_base_data_out_4, nx3158, nx3160, nx3170, nx3186, 
      addr1_data_4, nx3190, nx3196, bias_offset_data_out_4, nx3224, 
      img_base_addr_4, nx3242, nx3248, img_addr_offset_4, nx3256, nx3262, 
      nx3270, write_base_data_out_5, nx3294, nx3296, nx3298, nx3308, nx3312, 
      nx3318, nx3326, addr1_data_5, nx3354, bias_offset_data_out_5, nx3362, 
      nx3364, nx3374, img_base_addr_5, write_base_prev_data_out_5, nx3388, 
      img_addr_offset_5, nx3408, nx3410, nx3426, write_base_data_out_6, 
      nx3446, nx3448, nx3460, nx3466, addr1_data_6, nx3470, nx3476, 
      bias_offset_data_out_6, nx3504, img_base_addr_6, nx3522, nx3528, 
      img_addr_offset_6, nx3536, nx3542, nx3550, write_base_data_out_7, 
      nx3574, nx3576, nx3578, nx3588, nx3592, nx3598, nx3606, addr1_data_7, 
      nx3634, bias_offset_data_out_7, nx3642, nx3644, nx3654, 
      img_base_addr_7, write_base_prev_data_out_7, nx3668, img_addr_offset_7, 
      nx3688, nx3690, nx3706, write_base_data_out_8, nx3726, nx3728, nx3740, 
      nx3746, addr1_data_8, nx3750, nx3756, bias_offset_data_out_8, nx3784, 
      img_base_addr_8, nx3802, nx3808, img_addr_offset_8, nx3816, nx3822, 
      nx3830, write_base_data_out_9, nx3854, nx3856, nx3858, nx3868, nx3872, 
      nx3878, nx3886, addr1_data_9, nx3914, bias_offset_data_out_9, nx3922, 
      nx3924, nx3934, img_base_addr_9, write_base_prev_data_out_9, nx3948, 
      img_addr_offset_9, nx3968, nx3970, nx3986, write_base_data_out_10, 
      nx4006, nx4008, nx4020, nx4026, addr1_data_10, nx4030, nx4036, 
      bias_offset_data_out_10, nx4064, img_base_addr_10, nx4082, nx4088, 
      img_addr_offset_10, nx4096, nx4102, nx4110, write_base_data_out_11, 
      nx4134, nx4136, nx4138, nx4148, nx4152, nx4158, nx4166, addr1_data_11, 
      nx4194, bias_offset_data_out_11, nx4202, nx4204, nx4214, 
      img_base_addr_11, write_base_prev_data_out_11, nx4228, 
      img_addr_offset_11, nx4248, nx4250, nx4266, write_base_data_out_12, 
      nx4286, nx4288, nx4300, nx4306, addr1_data_12, nx4310, nx4316, 
      bias_offset_data_out_12, nx4344, img_base_addr_12, nx4362, nx4368, 
      img_addr_offset_12, nx4376, nx4382, nx4390, write_base_data_out_13, 
      nx4418, nx4428, nx4432, nx4438, nx4446, addr1_data_13, nx4474, 
      bias_offset_data_out_13, nx4482, nx4484, nx4494, img_base_addr_13, 
      write_base_prev_data_out_13, nx4508, img_addr_offset_13, nx4528, 
      nx4530, nx4546, write_base_data_out_14, nx4566, nx4568, nx4580, nx4586, 
      addr1_data_14, nx4590, nx4596, bias_offset_data_out_14, nx4624, 
      img_base_addr_14, nx4642, nx4648, img_addr_offset_14, nx4656, nx4662, 
      nx4670, nx4686, bias_offset_data_out_15, write_base_data_out_15, 
      nx4714, addr1_data_15, nx4734, nx4736, nx4744, nx4746, nx4756, 
      img_base_addr_15, write_base_prev_data_out_15, nx4764, nx4780, nx1479, 
      nx1489, nx1499, nx1509, nx1519, nx1529, nx1539, nx1549, nx1559, nx1569, 
      nx1579, nx1589, nx1599, nx1609, nx1619, nx1629, nx1639, nx1649, nx1659, 
      nx1669, nx1679, nx1689, nx1699, nx1709, nx1719, nx1729, nx1739, nx1749, 
      nx1759, nx1769, nx1779, nx1789, nx1799, nx1809, nx1819, nx1829, nx1839, 
      nx1849, nx1859, nx1869, nx1879, nx1889, nx1899, nx1909, nx1919, nx1929, 
      nx1939, nx1949, nx1959, nx1969, nx1979, nx1989, nx1999, nx2009, nx2019, 
      nx2029, nx2039, nx2049, nx2059, nx2069, nx2079, nx2089, nx2099, nx2109, 
      nx2119, nx2129, nx2139, nx2149, nx2159, nx2169, nx2179, nx2189, nx2199, 
      nx2209, nx2219, nx2229, nx2239, nx2249, nx2259, nx2269, nx2279, nx2289, 
      nx2299, nx2309, nx2319, nx2329, nx2339, nx2349, nx2359, nx2369, nx2379, 
      nx2389, nx2399, nx2409, nx2419, nx2429, nx2439, nx2449, nx2459, nx2469, 
      nx2479, nx2489, nx2499, nx2509, nx2519, nx2529, nx2539, nx2549, nx2559, 
      nx2569, nx2579, nx2589, nx2599, nx2609, nx2619, nx2629, nx2639, nx2649, 
      nx2659, nx2669, nx2679, nx2689, nx2699, nx2709, nx2719, nx2729, nx2739, 
      nx2749, nx2759, nx2769, nx2779, nx2789, nx2799, nx2809, nx2819, nx2829, 
      nx2839, nx2849, nx2859, nx2869, nx2879, nx2889, nx2899, nx2909, nx2919, 
      nx2929, nx2939, nx2949, nx2959, nx2969, nx2979, nx2989, nx2999, nx3009, 
      nx3019, nx3029, nx3039, nx3049, nx3059, nx3069, nx3079, nx3089, nx3099, 
      nx3109, nx3119, nx3129, nx3139, nx3149, nx3159, nx3169, nx3179, nx3189, 
      nx3199, nx3209, nx3219, nx3229, nx3239, nx3249, nx3259, nx3269, nx3279, 
      nx3289, nx3299, nx3309, nx3319, nx3329, nx3339, nx3349, nx3359, nx3369, 
      nx3379, nx3389, nx3399, nx3409, nx3419, nx3429, nx3439, nx3449, nx3459, 
      nx3469, nx3479, nx3489, nx3499, nx3509, nx3519, nx3529, nx3539, nx3549, 
      nx3559, nx3569, nx3579, nx3589, nx3599, nx3609, nx3619, nx3629, nx3639, 
      nx3649, nx3659, nx3669, nx3679, nx3689, nx3699, nx3709, nx3719, nx3729, 
      nx3739, nx3749, nx3759, nx3769, nx3779, nx3789, nx3799, nx3809, nx3819, 
      nx3829, nx3839, nx3849, nx3859, nx3869, nx3879, nx3889, nx3909, nx3919, 
      nx3929, nx3939, nx3957, nx3959, nx3967, nx3975, nx3979, nx3981, nx3989, 
      nx3999, nx4004, nx4009, nx4017, nx4019, nx4027, nx4031, nx4033, nx4039, 
      nx4041, nx4043, nx4045, nx4047, nx4053, nx4055, nx4057, nx4059, nx4065, 
      nx4067, nx4069, nx4073, nx4077, nx4080, nx4087, nx4099, nx4105, nx4109, 
      nx4111, nx4115, nx4119, nx4123, nx4129, nx4143, nx4149, nx4151, nx4153, 
      nx4157, nx4163, nx4167, nx4175, nx4180, nx4183, nx4191, nx4197, nx4200, 
      nx4207, nx4213, nx4217, nx4223, nx4229, nx4235, nx4239, nx4246, nx4251, 
      nx4253, nx4257, nx4265, nx4271, nx4277, nx4281, nx4284, nx4287, nx4293, 
      nx4295, nx4299, nx4301, nx4303, nx4305, nx4307, nx4314, nx4320, nx4321, 
      nx4328, nx4335, nx4337, nx4343, nx4349, nx4351, nx4358, nx4363, nx4365, 
      nx4372, nx4377, nx4379, nx4386, nx4391, nx4393, nx4400, nx4407, nx4408, 
      nx4417, nx4423, nx4427, nx4433, nx4435, nx4441, nx4447, nx4453, nx4459, 
      nx4460, nx4465, nx4469, nx4471, nx4480, nx4485, nx4487, nx4493, nx4497, 
      nx4499, nx4503, nx4507, nx4513, nx4515, nx4519, nx4526, nx4531, nx4533, 
      nx4535, nx4543, nx4553, nx4561, nx4563, nx4565, nx4571, nx4575, nx4579, 
      nx4581, nx4583, nx4589, nx4601, nx4609, nx4617, nx4621, nx4633, nx4635, 
      nx4637, nx4638, nx4647, nx4655, nx4657, nx4663, nx4669, nx4673, nx4681, 
      nx4689, nx4692, nx4701, nx4703, nx4705, nx4711, nx4717, nx4723, nx4725, 
      nx4731, nx4735, nx4743, nx4747, nx4751, nx4759, nx4761, nx4765, nx4767, 
      nx4770, nx4776, nx4781, nx4783, nx4787, nx4795, nx4801, nx4803, nx4807, 
      nx4813, nx4819, nx4821, nx4825, nx4833, nx4839, nx4841, nx4845, nx4853, 
      nx4861, nx4879, nx4881, nx4883, nx4895, nx4903, nx4911, nx4913, nx4927, 
      nx4941, nx4957, nx4961, nx4975, nx4977, nx4981, nx4993, nx4997, nx5009, 
      nx5011, nx5013, nx5019, nx5023, nx5031, nx5037, nx5041, nx5049, nx5055, 
      nx5059, nx5067, nx5072, nx5077, nx5083, nx5089, nx5099, nx5107, nx5113, 
      nx5115, nx5122, nx5128, nx5134, nx5137, nx5140, nx5142, nx5144, nx5146, 
      nx5148, nx5155, nx5157, nx5162, nx5164, nx5168, nx5188, nx5194, nx5197, 
      nx5202, nx5204, nx5206, nx5208, nx5216, nx5218, nx5243, nx5330, nx5334, 
      nx5379, nx5383, nx5386, nx5390, nx5393, nx5396, nx5399, nx5402, nx5405, 
      nx5408, nx5411, nx5414, nx5417, nx5420, nx5423, nx5426, nx5429, nx5432, 
      nx5435, nx5438, nx5441, nx5444, nx5447, nx5450, nx5453, nx5456, nx5459, 
      nx5462, nx5465, nx5468, nx5471, nx5474, nx5477, nx5480, nx5482, nx5501, 
      nx5587, nx5593, nx5596, nx5598, nx5605, nx5607, nx5611, nx5614, nx5616, 
      nx5619, nx5621, nx5629, nx5632, nx5636, nx5647, nx5651, nx5653, nx5657, 
      nx5659, nx5662, nx5664, nx5670, nx5673, nx5677, nx5679, nx5685, nx5687, 
      nx5692, nx5696, nx5698, nx5700, nx5703, nx5707, nx5709, nx5712, nx5714, 
      nx5718, nx5720, nx5722, nx5728, nx5731, nx5734, nx5737, nx5742, nx5747, 
      nx5749, nx5758, nx5762, nx5764, nx5767, nx5771, nx5773, nx5777, nx5783, 
      nx5790, nx5794, nx5805, nx5807, nx5809, nx5815, nx5820, nx5826, nx5829, 
      nx5831, nx5834, nx5836, nx5838, nx5843, nx5850, nx5853, nx5856, nx5859, 
      nx5864, nx5869, nx5871, nx5873, nx5876, nx5879, nx5882, nx5886, nx5888, 
      nx5892, nx5895, nx5900, nx5901, nx5906, nx5908, nx5913, nx5917, nx5921, 
      nx5925, nx5936, nx5938, nx5943, nx5945, nx5947, nx5951, nx5955, nx5957, 
      nx5961, nx5963, nx5965, nx5968, nx5971, nx5974, nx5977, nx5980, nx5983, 
      nx5986, nx5991, nx5996, nx5998, nx6000, nx6003, nx6006, nx6009, nx6013, 
      nx6017, nx6020, nx6025, nx6026, nx6031, nx6034, nx6037, nx6039, nx6042, 
      nx6045, nx6049, nx6060, nx6062, nx6067, nx6069, nx6071, nx6075, nx6079, 
      nx6081, nx6085, nx6088, nx6090, nx6097, nx6100, nx6103, nx6106, nx6109, 
      nx6114, nx6119, nx6121, nx6123, nx6126, nx6129, nx6132, nx6136, nx6140, 
      nx6143, nx6148, nx6149, nx6154, nx6157, nx6160, nx6162, nx6164, nx6167, 
      nx6171, nx6182, nx6184, nx6189, nx6191, nx6193, nx6197, nx6201, nx6203, 
      nx6207, nx6210, nx6212, nx6219, nx6222, nx6225, nx6228, nx6231, nx6236, 
      nx6241, nx6243, nx6245, nx6248, nx6251, nx6254, nx6258, nx6262, nx6265, 
      nx6270, nx6271, nx6276, nx6279, nx6282, nx6284, nx6286, nx6289, nx6293, 
      nx6304, nx6306, nx6311, nx6313, nx6315, nx6319, nx6323, nx6325, nx6329, 
      nx6332, nx6334, nx6341, nx6344, nx6347, nx6350, nx6353, nx6358, nx6363, 
      nx6365, nx6367, nx6373, nx6376, nx6380, nx6384, nx6387, nx6392, nx6393, 
      nx6398, nx6400, nx6402, nx6404, nx6408, nx6411, nx6415, nx6426, nx6428, 
      nx6433, nx6435, nx6437, nx6441, nx6445, nx6447, nx6451, nx6454, nx6456, 
      nx6463, nx6466, nx6469, nx6472, nx6475, nx6484, nx6486, nx6493, nx6494, 
      nx6496, nx6500, nx6502, nx6505, nx6510, nx6511, nx6516, nx6518, nx6520, 
      nx6524, nx6527, nx6532, nx6543, nx6555, nx6558, nx6560, nx6563, nx6569, 
      nx6572, nx6576, nx6580, nx6583, nx6586, nx6589, nx6592, nx6599, nx6601, 
      nx6603, nx6605, nx6607, nx6609, nx6611, nx6613, nx6615, nx6617, nx6619, 
      nx6621, nx6623, nx6625, nx6627, nx6629, nx6631, nx6633, nx6635, nx6637, 
      nx6639, nx6641, nx6643, nx6651, nx6653, nx6655, nx6657, nx6659, nx6663, 
      nx6665, nx6667, nx6673, nx6675, nx6677, nx6679, nx6681, nx6683, nx6685, 
      nx6687, nx6689, nx6691, nx6693, nx6695, nx6699, nx6705, nx6713, nx6721, 
      nx6723, nx6725, nx6727, nx6729, nx6731, nx6733, nx6735, nx6737, nx6739, 
      nx6741, nx6743, nx6749, nx6759, nx6761, nx6763, nx6765, nx6767, nx6769, 
      nx6771, nx6773, nx6781, nx6787, nx6793, nx6795, nx6797, nx6799, nx6801, 
      nx6803, nx6805, nx6807, nx6809, nx6811, nx6813, nx6815, nx6817, nx6819, 
      nx6821, nx6823, nx6825, nx6827, nx6829, nx6831, nx6833, nx6835, nx6837, 
      nx6839, nx6851, nx6855, nx6857, nx6859, nx6871, nx6897, nx6899, nx6901, 
      nx6903, nx6905, nx6927, nx6929, nx6931, nx6933, nx6939, nx6941, nx6943, 
      nx6945, nx6947, nx6949, nx6951, nx6953, nx6955, nx6957, nx6959, nx6961, 
      nx6963, nx6965, nx6967, nx6969, nx6971, nx6973, nx6975, nx6977, nx6979, 
      nx6981, nx6983, nx6985, nx6987, nx6989, nx6991, nx6993, nx6995, nx6997, 
      nx6999, nx7001, nx7003, nx7005, nx7007, nx7009, nx7011, nx7013, nx7015, 
      nx7017, nx7019, nx7021, nx7023, nx7025, nx7027, nx7033, nx7035, nx7037, 
      nx7039, nx7041, nx7043, nx7049, nx7051, nx7053, nx7055, nx7057, nx7059, 
      nx7061, nx7065, nx7071, nx7073, nx7075, nx7077, nx7079, nx7081, nx7083, 
      nx7085, nx7087, nx7089, nx7091, nx7093, nx7095, nx7097, nx7099, nx7101, 
      nx7103, nx7105, nx7107, nx7109, nx7111, nx7113, nx7115, nx7117, nx7119, 
      nx7121, nx7123, nx7125, nx7127, nx7129, nx7131, nx7133, nx7135, nx7137, 
      nx7139, nx7145, filter_ready_out_EXMPLR, nx7029, nx4593, nx4665, 
      nx7063, comp_unit_flt_size_EXMPLR, nx7031, nx6711, nx7293, nx7294, 
      nx7295, nx7296, nx7297, nx7298, nx7299, nx7300, nx7301, nx7302, nx7303, 
      nx7304, nx7305, nx3899, nx7306, nx7307, nx6488, nx7308, nx7309, nx6491, 
      nx4414, nx7310, nx7311, nx6370, nx7312, nx7313, nx7314, nx7315, nx7316, 
      nx7317, nx7318, nx7319, nx7320, nx7321, nx7322, nx3002, nx7323, nx5751, 
      nx5754, nx5689, nx7324, nx5191, argmax_ready_dup0, nx7325, nx7326, 
      nx7327, nx7328, nx1930, nx7329, nx7330, nx7331, nx7332, nx7333, nx7334, 
      nx7335, nx5847, nx7336, nx7337, nx2850, nx5667, nx5725, nx6775, nx7047, 
      nx7338, nx7339, nx7340, argmax_ready_XX0_XREP5, nx7341, nx7342, nx7343, 
      nx7344, nx7345, nx7346, nx7347, nx7348, nx7349, nx7350, nx7351, nx7352, 
      nx7353, NOT_nx4700, nx7354, nx7355, nx7356, nx7357, nx7358, nx7359, 
      nx7360, nx7361, nx7362, nx7363, nx7364, nx7365, nx7366, 
      argmax_ready_EXMPLR, nx7367, nx7445: std_logic ;
   
   signal DANGLING : std_logic_vector (15 downto 0 );

begin
   io_done_out <= filter_reset_EXMPLR ;
   wind_rst <= filter_reset_EXMPLR ;
   filter_ready_out <= filter_ready_out_EXMPLR ;
   filter_reset <= filter_reset_EXMPLR ;
   comp_unit_operation <= comp_unit_operation_EXMPLR ;
   comp_unit_flt_size <= comp_unit_flt_size_EXMPLR ;
   argmax_ready <= argmax_ready_EXMPLR ;
   img_cache : Cache_5_16_28_5 port map ( in_word(15)=>cache_data_in_15, 
      in_word(14)=>cache_data_in_14, in_word(13)=>cache_data_in_13, 
      in_word(12)=>cache_data_in_12, in_word(11)=>cache_data_in_11, 
      in_word(10)=>cache_data_in_10, in_word(9)=>cache_data_in_9, in_word(8)
      =>cache_data_in_8, in_word(7)=>cache_data_in_7, in_word(6)=>
      cache_data_in_6, in_word(5)=>cache_data_in_5, in_word(4)=>
      cache_data_in_4, in_word(3)=>cache_data_in_3, in_word(2)=>
      cache_data_in_2, in_word(1)=>cache_data_in_1, in_word(0)=>
      cache_data_in_0, cache_in_sel(4)=>nx6611, cache_in_sel(3)=>
      cache_width_count_3, cache_in_sel(2)=>nx6615, cache_in_sel(1)=>
      cache_width_count_1, cache_in_sel(0)=>cache_width_count_0, 
      cache_out_sel(4)=>wind_width_count_4, cache_out_sel(3)=>
      wind_width_count_3, cache_out_sel(2)=>wind_width_count_2, 
      cache_out_sel(1)=>wind_width_count_1, cache_out_sel(0)=>nx6607, 
      decoder_enable=>cache_load, out_column_0_15=>cache_data_out_4_15, 
      out_column_0_14=>cache_data_out_4_14, out_column_0_13=>
      cache_data_out_4_13, out_column_0_12=>cache_data_out_4_12, 
      out_column_0_11=>cache_data_out_4_11, out_column_0_10=>
      cache_data_out_4_10, out_column_0_9=>cache_data_out_4_9, 
      out_column_0_8=>cache_data_out_4_8, out_column_0_7=>cache_data_out_4_7, 
      out_column_0_6=>cache_data_out_4_6, out_column_0_5=>cache_data_out_4_5, 
      out_column_0_4=>cache_data_out_4_4, out_column_0_3=>cache_data_out_4_3, 
      out_column_0_2=>cache_data_out_4_2, out_column_0_1=>cache_data_out_4_1, 
      out_column_0_0=>cache_data_out_4_0, out_column_1_15=>
      cache_data_out_3_15, out_column_1_14=>cache_data_out_3_14, 
      out_column_1_13=>cache_data_out_3_13, out_column_1_12=>
      cache_data_out_3_12, out_column_1_11=>cache_data_out_3_11, 
      out_column_1_10=>cache_data_out_3_10, out_column_1_9=>
      cache_data_out_3_9, out_column_1_8=>cache_data_out_3_8, out_column_1_7
      =>cache_data_out_3_7, out_column_1_6=>cache_data_out_3_6, 
      out_column_1_5=>cache_data_out_3_5, out_column_1_4=>cache_data_out_3_4, 
      out_column_1_3=>cache_data_out_3_3, out_column_1_2=>cache_data_out_3_2, 
      out_column_1_1=>cache_data_out_3_1, out_column_1_0=>cache_data_out_3_0, 
      out_column_2_15=>cache_data_out_2_15, out_column_2_14=>
      cache_data_out_2_14, out_column_2_13=>cache_data_out_2_13, 
      out_column_2_12=>cache_data_out_2_12, out_column_2_11=>
      cache_data_out_2_11, out_column_2_10=>cache_data_out_2_10, 
      out_column_2_9=>cache_data_out_2_9, out_column_2_8=>cache_data_out_2_8, 
      out_column_2_7=>cache_data_out_2_7, out_column_2_6=>cache_data_out_2_6, 
      out_column_2_5=>cache_data_out_2_5, out_column_2_4=>cache_data_out_2_4, 
      out_column_2_3=>cache_data_out_2_3, out_column_2_2=>cache_data_out_2_2, 
      out_column_2_1=>cache_data_out_2_1, out_column_2_0=>cache_data_out_2_0, 
      out_column_3_15=>cache_data_out_1_15, out_column_3_14=>
      cache_data_out_1_14, out_column_3_13=>cache_data_out_1_13, 
      out_column_3_12=>cache_data_out_1_12, out_column_3_11=>
      cache_data_out_1_11, out_column_3_10=>cache_data_out_1_10, 
      out_column_3_9=>cache_data_out_1_9, out_column_3_8=>cache_data_out_1_8, 
      out_column_3_7=>cache_data_out_1_7, out_column_3_6=>cache_data_out_1_6, 
      out_column_3_5=>cache_data_out_1_5, out_column_3_4=>cache_data_out_1_4, 
      out_column_3_3=>cache_data_out_1_3, out_column_3_2=>cache_data_out_1_2, 
      out_column_3_1=>cache_data_out_1_1, out_column_3_0=>cache_data_out_1_0, 
      out_column_4_15=>cache_data_out_0_15, out_column_4_14=>
      cache_data_out_0_14, out_column_4_13=>cache_data_out_0_13, 
      out_column_4_12=>cache_data_out_0_12, out_column_4_11=>
      cache_data_out_0_11, out_column_4_10=>cache_data_out_0_10, 
      out_column_4_9=>cache_data_out_0_9, out_column_4_8=>cache_data_out_0_8, 
      out_column_4_7=>cache_data_out_0_7, out_column_4_6=>cache_data_out_0_6, 
      out_column_4_5=>cache_data_out_0_5, out_column_4_4=>cache_data_out_0_4, 
      out_column_4_3=>cache_data_out_0_3, out_column_4_2=>cache_data_out_0_2, 
      out_column_4_1=>cache_data_out_0_1, out_column_4_0=>cache_data_out_0_0, 
      clk=>nx6619, reset=>cache_rst_actual);
   cache_height_cntr : AdvancedCounter_16 port map ( clk=>clk, reset=>nx6601, 
      enable=>cache_height_count_en, mode_in(1)=>filter_reset_EXMPLR, 
      mode_in(0)=>filter_reset_EXMPLR, max_val_in(15)=>filter_reset_EXMPLR, 
      max_val_in(14)=>filter_reset_EXMPLR, max_val_in(13)=>
      filter_reset_EXMPLR, max_val_in(12)=>filter_reset_EXMPLR, 
      max_val_in(11)=>filter_reset_EXMPLR, max_val_in(10)=>
      filter_reset_EXMPLR, max_val_in(9)=>filter_reset_EXMPLR, max_val_in(8)
      =>filter_reset_EXMPLR, max_val_in(7)=>filter_reset_EXMPLR, 
      max_val_in(6)=>filter_reset_EXMPLR, max_val_in(5)=>filter_reset_EXMPLR, 
      max_val_in(4)=>max_height_4, max_val_in(3)=>max_height_3, 
      max_val_in(2)=>max_height_2, max_val_in(1)=>max_height_1, 
      max_val_in(0)=>max_height_0, max_reached_out=>cache_height_ended, 
      counter_out(15)=>DANGLING(0), counter_out(14)=>DANGLING(1), 
      counter_out(13)=>DANGLING(2), counter_out(12)=>DANGLING(3), 
      counter_out(11)=>DANGLING(4), counter_out(10)=>DANGLING(5), 
      counter_out(9)=>DANGLING(6), counter_out(8)=>DANGLING(7), 
      counter_out(7)=>DANGLING(8), counter_out(6)=>DANGLING(9), 
      counter_out(5)=>DANGLING(10), counter_out(4)=>DANGLING(11), 
      counter_out(3)=>DANGLING(12), counter_out(2)=>DANGLING(13), 
      counter_out(1)=>DANGLING(14), counter_out(0)=>DANGLING(15));
   ix1260 : fake_gnd port map ( Y=>filter_reset_EXMPLR);
   ix2001 : ao22 port map ( Y=>mem_data_out(4), A0=>comp_unit_data2_in(4), 
      A1=>nx6673, B0=>comp_unit_data1_in(4), B1=>nx6679);
   ix1487 : nand02 port map ( Y=>nx1486, A0=>nx3957, A1=>nx5011);
   ix3958 : aoi32 port map ( Y=>nx3957, A0=>nx3959, A1=>comp_unit_finished, 
      A2=>current_state_19, B0=>nx4563, B1=>nx1459);
   layer_type_reg_q_0 : dffr port map ( Q=>comp_unit_operation_EXMPLR, QB=>
      OPEN, D=>nx1519, CLK=>clk, R=>reset);
   ix1520 : mux21_ni port map ( Y=>nx1519, A0=>nx6927, A1=>mem_data_in(0), 
      S0=>current_state_3);
   reg_current_state_3 : dffr port map ( Q=>current_state_3, QB=>OPEN, D=>
      nx1461, CLK=>nx6627, R=>reset);
   reg_current_state_2 : dffr port map ( Q=>current_state_2, QB=>nx3967, D=>
      nx1578, CLK=>nx6619, R=>reset);
   ix1573 : oai21 port map ( Y=>nx1572, A0=>io_ready_in, A1=>nx3975, B0=>
      nx3979);
   reg_current_state_1 : dffr port map ( Q=>OPEN, QB=>nx3975, D=>nx1572, CLK
      =>nx6619, R=>reset);
   reg_current_state_0 : dffs_ni port map ( Q=>OPEN, QB=>nx3979, D=>
      filter_reset_EXMPLR, CLK=>nx6619, S=>reset);
   ix1737 : nand02 port map ( Y=>nx1409, A0=>nx3989, A1=>nx4503);
   ix2470 : mux21_ni port map ( Y=>nx2469, A0=>nx1620, A1=>
      num_channels_out_0, S0=>nx4115);
   ix1611 : nand03 port map ( Y=>nx1610, A0=>nx3999, A1=>nx4105, A2=>nx3967
   );
   ix4000 : oai21 port map ( Y=>nx3999, A0=>nx1602, A1=>current_state_25, B0
      =>max_num_channels_data_out_0);
   ix2590 : mux21_ni port map ( Y=>nx2589, A0=>layer_type_out_1, A1=>
      mem_data_in(1), S0=>current_state_3);
   layer_type_reg_q_1 : dffr port map ( Q=>layer_type_out_1, QB=>nx4004, D=>
      nx2589, CLK=>clk, R=>reset);
   reg_current_state_26 : dffr port map ( Q=>OPEN, QB=>nx3981, D=>nx1800, 
      CLK=>nx6619, R=>reset);
   reg_current_state_25 : dffr port map ( Q=>current_state_25, QB=>nx4073, D
      =>nx112, CLK=>nx6619, R=>reset);
   ix1480 : oai32 port map ( Y=>nx1479, A0=>nx4019, A1=>nx6689, A2=>
      current_state_25, B0=>nx4027, B1=>nx7017);
   reg_current_state_4 : dffr port map ( Q=>current_state_4, QB=>OPEN, D=>
      current_state_3, CLK=>nx6619, R=>reset);
   reg_nflt_layer_out_0 : dffr port map ( Q=>nflt_layer_out_0, QB=>nx4019, D
      =>nx1479, CLK=>clk, R=>reset);
   ix4032 : inv01 port map ( Y=>nx4031, A=>mem_data_in(0));
   ix1490 : oai32 port map ( Y=>nx1489, A0=>nx4039, A1=>nx6689, A2=>
      current_state_25, B0=>nx4041, B1=>nx7017);
   reg_nflt_layer_out_1 : dffr port map ( Q=>nflt_layer_out_1, QB=>nx4039, D
      =>nx1489, CLK=>clk, R=>reset);
   ix4042 : mux21_ni port map ( Y=>nx4041, A0=>nx4043, A1=>nx4047, S0=>
      nx6689);
   ix4044 : aoi21 port map ( Y=>nx4043, A0=>nflt_layer_out_1, A1=>
      nflt_layer_out_0, B0=>nx4045);
   ix4048 : inv01 port map ( Y=>nx4047, A=>mem_data_in(1));
   ix1500 : oai32 port map ( Y=>nx1499, A0=>nx4053, A1=>nx6689, A2=>
      current_state_25, B0=>nx4055, B1=>nx7017);
   nflt_layer_out_2 : dffr port map ( Q=>OPEN, QB=>nx4053, D=>nx1499, CLK=>
      clk, R=>reset);
   ix4056 : mux21_ni port map ( Y=>nx4055, A0=>nx4057, A1=>nx4059, S0=>
      nx6689);
   ix4060 : inv01 port map ( Y=>nx4059, A=>mem_data_in(2));
   reg_nflt_layer_out_3 : dffr port map ( Q=>nflt_layer_out_3, QB=>OPEN, D=>
      nx1509, CLK=>clk, R=>reset);
   ix1510 : mux21_ni port map ( Y=>nx1509, A0=>nx98, A1=>nflt_layer_out_3, 
      S0=>nx7017);
   ix99 : mux21 port map ( Y=>nx98, A0=>nx4065, A1=>nx4069, S0=>nx6691);
   ix4066 : xnor2 port map ( Y=>nx4065, A0=>nflt_layer_out_3, A1=>nx4067);
   ix4070 : inv01 port map ( Y=>nx4069, A=>mem_data_in(3));
   ix2460 : oai222 port map ( Y=>nx2459, A0=>nx4077, A1=>nx1594, B0=>nx4099, 
      B1=>nx7019, C0=>nx4031, C1=>nx6821);
   max_num_channels_inst_reg_q_0 : dffs_ni port map ( Q=>
      max_num_channels_data_out_0, QB=>nx4077, D=>nx2459, CLK=>clk, S=>reset
   );
   ix1595 : nand02 port map ( Y=>nx1594, A0=>nx7019, A1=>nx6821);
   reg_current_state_9 : dffr port map ( Q=>current_state_9, QB=>OPEN, D=>
      nx136, CLK=>nx6621, R=>reset);
   ix137 : nor03_2x port map ( Y=>nx136, A0=>nx4087, A1=>nx6927, A2=>nx4004
   );
   reg_current_state_8 : dffr port map ( Q=>current_state_8, QB=>nx4087, D=>
      nx6699, CLK=>nx6621, R=>reset);
   reg_current_state_7 : dffr port map ( Q=>current_state_7, QB=>OPEN, D=>
      current_state_6, CLK=>nx6621, R=>reset);
   reg_current_state_6 : dffr port map ( Q=>current_state_6, QB=>OPEN, D=>
      current_state_5, CLK=>nx6621, R=>reset);
   reg_current_state_5 : dffr port map ( Q=>current_state_5, QB=>OPEN, D=>
      nx6691, CLK=>nx6621, R=>reset);
   ix2450 : mux21_ni port map ( Y=>nx2449, A0=>nflt_layer_temp_0, A1=>
      mem_data_in(0), S0=>nx6691);
   nflt_layer_total_reg_q_0 : dffr port map ( Q=>nflt_layer_temp_0, QB=>
      nx4099, D=>nx2449, CLK=>clk, R=>reset);
   ix4106 : aoi22 port map ( Y=>nx4105, A0=>mem_data_in(0), A1=>nx6693, B0=>
      nflt_layer_temp_0, B1=>nx1528);
   reg_num_channels_out_0 : dffr port map ( Q=>num_channels_out_0, QB=>
      nx4111, D=>nx2469, CLK=>clk, R=>reset);
   ix4116 : nor02_2x port map ( Y=>nx4115, A0=>nx1516, A1=>nx1421);
   ix1513 : nor02ii port map ( Y=>nx1421, A0=>nx4123, A1=>nx1409);
   ix4124 : nand02 port map ( Y=>nx4123, A0=>current_state_24, A1=>nx4153);
   reg_current_state_24 : dffr port map ( Q=>current_state_24, QB=>nx4151, D
      =>nx1502, CLK=>nx6623, R=>reset);
   ix1503 : oai21 port map ( Y=>nx1502, A0=>nx4129, A1=>nx6641, B0=>nx4149);
   reg_current_state_22 : dffr port map ( Q=>OPEN, QB=>nx4129, D=>nx1486, 
      CLK=>nx6621, R=>reset);
   ix1590 : mux21_ni port map ( Y=>nx1589, A0=>flt_size_out_0, A1=>
      mem_data_in(0), S0=>current_state_5);
   flt_size_reg_q_0 : dffr port map ( Q=>flt_size_out_0, QB=>OPEN, D=>nx1589, 
      CLK=>clk, R=>reset);
   flt_size_reg_q_2 : dffr port map ( Q=>flt_size_out_2, QB=>nx4143, D=>
      nx1599, CLK=>clk, R=>reset);
   ix1600 : mux21_ni port map ( Y=>nx1599, A0=>flt_size_out_2, A1=>
      mem_data_in(2), S0=>current_state_5);
   ix1610 : mux21_ni port map ( Y=>nx1609, A0=>flt_size_out_1, A1=>
      mem_data_in(1), S0=>current_state_5);
   flt_size_reg_q_1 : dffr port map ( Q=>flt_size_out_1, QB=>OPEN, D=>nx1609, 
      CLK=>clk, R=>reset);
   reg_current_state_23 : dffr port map ( Q=>OPEN, QB=>nx4149, D=>nx1492, 
      CLK=>nx6621, R=>reset);
   ix4154 : nor04 port map ( Y=>nx4153, A0=>nx1098, A1=>nx1010, A2=>nx914, 
      A3=>nx820);
   ix1099 : nand04 port map ( Y=>nx1098, A0=>nx4157, A1=>nx4314, A2=>nx4321, 
      A3=>nx4328);
   ix2210 : oai22 port map ( Y=>nx2209, A0=>nx4163, A1=>nx6833, B0=>nx4307, 
      B1=>nx6735);
   reg_write_offset_reg_q_14 : dffr port map ( Q=>write_offset_data_out_14, 
      QB=>nx4167, D=>nx2189, CLK=>nx6623, R=>reset);
   ix4176 : nand02 port map ( Y=>nx4175, A0=>write_offset_data_out_13, A1=>
      nx1012);
   ix2170 : oai22 port map ( Y=>nx2169, A0=>nx4180, A1=>nx6833, B0=>nx4305, 
      B1=>nx6733);
   ix4181 : oai21 port map ( Y=>nx4180, A0=>nx1012, A1=>
      write_offset_data_out_13, B0=>nx4175);
   reg_write_offset_reg_q_12 : dffr port map ( Q=>write_offset_data_out_12, 
      QB=>nx4183, D=>nx2149, CLK=>nx6623, R=>reset);
   ix4192 : nand02 port map ( Y=>nx4191, A0=>write_offset_data_out_11, A1=>
      nx964);
   ix2130 : oai22 port map ( Y=>nx2129, A0=>nx4197, A1=>nx6831, B0=>nx4303, 
      B1=>nx6733);
   ix4198 : oai21 port map ( Y=>nx4197, A0=>nx964, A1=>
      write_offset_data_out_11, B0=>nx4191);
   reg_write_offset_reg_q_10 : dffr port map ( Q=>write_offset_data_out_10, 
      QB=>nx4200, D=>nx2109, CLK=>nx6623, R=>reset);
   ix4208 : nand02 port map ( Y=>nx4207, A0=>write_offset_data_out_9, A1=>
      nx918);
   ix2090 : oai22 port map ( Y=>nx2089, A0=>nx4213, A1=>nx6831, B0=>nx4301, 
      B1=>nx6733);
   ix4214 : oai21 port map ( Y=>nx4213, A0=>nx918, A1=>
      write_offset_data_out_9, B0=>nx4207);
   reg_write_offset_reg_q_8 : dffr port map ( Q=>write_offset_data_out_8, QB
      =>nx4217, D=>nx2069, CLK=>nx6623, R=>reset);
   ix4224 : nand02 port map ( Y=>nx4223, A0=>write_offset_data_out_7, A1=>
      nx868);
   ix2050 : oai22 port map ( Y=>nx2049, A0=>nx4229, A1=>nx6731, B0=>nx4235, 
      B1=>nx6831);
   reg_write_offset_reg_q_7 : dffr port map ( Q=>write_offset_data_out_7, QB
      =>nx4229, D=>nx2049, CLK=>nx6623, R=>reset);
   ix4236 : oai21 port map ( Y=>nx4235, A0=>nx868, A1=>
      write_offset_data_out_7, B0=>nx4223);
   reg_write_offset_reg_q_6 : dffr port map ( Q=>write_offset_data_out_6, QB
      =>nx4239, D=>nx2029, CLK=>nx6623, R=>reset);
   ix4247 : nand02 port map ( Y=>nx4246, A0=>write_offset_data_out_5, A1=>
      nx822);
   ix2010 : oai22 port map ( Y=>nx2009, A0=>nx4251, A1=>nx6731, B0=>nx4253, 
      B1=>nx6829);
   reg_write_offset_reg_q_5 : dffr port map ( Q=>write_offset_data_out_5, QB
      =>nx4251, D=>nx2009, CLK=>nx6625, R=>reset);
   ix4254 : oai21 port map ( Y=>nx4253, A0=>nx822, A1=>
      write_offset_data_out_5, B0=>nx4246);
   reg_write_offset_reg_q_4 : dffr port map ( Q=>write_offset_data_out_4, QB
      =>nx4257, D=>nx1989, CLK=>nx6625, R=>reset);
   reg_write_offset_reg_q_3 : dffr port map ( Q=>write_offset_data_out_3, QB
      =>nx4271, D=>nx1969, CLK=>nx6625, R=>reset);
   ix1950 : oai22 port map ( Y=>nx1949, A0=>nx4277, A1=>nx6731, B0=>nx4281, 
      B1=>nx6829);
   ix4282 : oai21 port map ( Y=>nx4281, A0=>nx750, A1=>
      write_offset_data_out_2, B0=>nx4299);
   ix1930 : oai22 port map ( Y=>nx1929, A0=>nx7355, A1=>nx6731, B0=>nx4287, 
      B1=>nx6829);
   ix4288 : oai21 port map ( Y=>nx4287, A0=>write_offset_data_out_0, A1=>
      write_offset_data_out_1, B0=>nx4295);
   reg_write_offset_reg_q_0 : dffr port map ( Q=>write_offset_data_out_0, QB
      =>nx4293, D=>nx1909, CLK=>nx6625, R=>reset);
   reg_write_offset_reg_q_1 : dffr port map ( Q=>write_offset_data_out_1, QB
      =>nx4284, D=>nx1929, CLK=>nx6625, R=>reset);
   reg_write_offset_reg_q_2 : dffr port map ( Q=>write_offset_data_out_2, QB
      =>nx4277, D=>nx1949, CLK=>nx6625, R=>reset);
   reg_write_offset_reg_q_9 : dffr port map ( Q=>write_offset_data_out_9, QB
      =>nx4301, D=>nx2089, CLK=>nx6625, R=>reset);
   reg_write_offset_reg_q_11 : dffr port map ( Q=>write_offset_data_out_11, 
      QB=>nx4303, D=>nx2129, CLK=>nx6627, R=>reset);
   reg_write_offset_reg_q_13 : dffr port map ( Q=>write_offset_data_out_13, 
      QB=>nx4305, D=>nx2169, CLK=>nx6627, R=>reset);
   reg_write_offset_reg_q_15 : dffr port map ( Q=>write_offset_data_out_15, 
      QB=>nx4307, D=>nx2209, CLK=>nx6627, R=>reset);
   new_size_squared_reg_q_15 : dffr port map ( Q=>new_size_squared_out_15, 
      QB=>OPEN, D=>nx2219, CLK=>clk, R=>reset);
   new_size_squared_reg_q_14 : dffr port map ( Q=>new_size_squared_out_14, 
      QB=>nx4320, D=>nx2199, CLK=>clk, R=>reset);
   new_size_squared_reg_q_13 : dffr port map ( Q=>new_size_squared_out_13, 
      QB=>OPEN, D=>nx2179, CLK=>clk, R=>reset);
   new_size_squared_reg_q_12 : dffr port map ( Q=>new_size_squared_out_12, 
      QB=>nx4335, D=>nx2159, CLK=>clk, R=>reset);
   ix1011 : nand04 port map ( Y=>nx1010, A0=>nx4337, A1=>nx4343, A2=>nx4351, 
      A3=>nx4358);
   new_size_squared_reg_q_11 : dffr port map ( Q=>new_size_squared_out_11, 
      QB=>OPEN, D=>nx2139, CLK=>clk, R=>reset);
   new_size_squared_reg_q_10 : dffr port map ( Q=>new_size_squared_out_10, 
      QB=>nx4349, D=>nx2119, CLK=>clk, R=>reset);
   new_size_squared_reg_q_9 : dffr port map ( Q=>new_size_squared_out_9, QB
      =>OPEN, D=>nx2099, CLK=>clk, R=>reset);
   new_size_squared_reg_q_8 : dffr port map ( Q=>new_size_squared_out_8, QB
      =>nx4363, D=>nx2079, CLK=>clk, R=>reset);
   ix915 : nand04 port map ( Y=>nx914, A0=>nx4365, A1=>nx4372, A2=>nx4379, 
      A3=>nx4386);
   new_size_squared_reg_q_7 : dffr port map ( Q=>new_size_squared_out_7, QB
      =>OPEN, D=>nx2059, CLK=>clk, R=>reset);
   new_size_squared_reg_q_6 : dffr port map ( Q=>new_size_squared_out_6, QB
      =>nx4377, D=>nx2039, CLK=>clk, R=>reset);
   new_size_squared_reg_q_5 : dffr port map ( Q=>new_size_squared_out_5, QB
      =>OPEN, D=>nx2019, CLK=>clk, R=>reset);
   new_size_squared_reg_q_4 : dffr port map ( Q=>new_size_squared_out_4, QB
      =>nx4391, D=>nx1999, CLK=>clk, R=>reset);
   ix821 : nand04 port map ( Y=>nx820, A0=>nx4393, A1=>nx4400, A2=>nx4408, 
      A3=>nx4417);
   new_size_squared_reg_q_3 : dffr port map ( Q=>new_size_squared_out_3, QB
      =>OPEN, D=>nx1979, CLK=>clk, R=>reset);
   new_size_squared_reg_q_2 : dffr port map ( Q=>new_size_squared_out_2, QB
      =>nx4407, D=>nx1959, CLK=>clk, R=>reset);
   new_size_squared_reg_q_1 : dffr port map ( Q=>new_size_squared_out_1, QB
      =>OPEN, D=>nx1939, CLK=>clk, R=>reset);
   new_size_squared_reg_q_0 : dffr port map ( Q=>new_size_squared_out_0, QB
      =>nx4423, D=>nx1919, CLK=>clk, R=>reset);
   reg_num_channels_out_1 : dffr port map ( Q=>num_channels_out_1, QB=>
      nx4447, D=>nx2489, CLK=>clk, R=>reset);
   ix2490 : mux21_ni port map ( Y=>nx2489, A0=>nx1652, A1=>
      num_channels_out_1, S0=>nx4115);
   ix1653 : oai21 port map ( Y=>nx1652, A0=>nx4427, A1=>nx6825, B0=>nx4435);
   ix4428 : aoi22 port map ( Y=>nx4427, A0=>mem_data_in(1), A1=>nx6693, B0=>
      nflt_layer_temp_1, B1=>nx1528);
   nflt_layer_total_reg_q_1 : dffr port map ( Q=>nflt_layer_temp_1, QB=>
      nx4433, D=>nx2439, CLK=>clk, R=>reset);
   ix2440 : mux21_ni port map ( Y=>nx2439, A0=>nflt_layer_temp_1, A1=>
      mem_data_in(1), S0=>nx6691);
   ix4436 : aoi22 port map ( Y=>nx4435, A0=>max_num_channels_data_out_1, A1
      =>nx1646, B0=>nx6825, B1=>nx1630);
   ix2480 : oai222 port map ( Y=>nx2479, A0=>nx4441, A1=>nx1594, B0=>nx4433, 
      B1=>nx7019, C0=>nx4047, C1=>nx6821);
   max_num_channels_inst_reg_q_1 : dffr port map ( Q=>
      max_num_channels_data_out_1, QB=>nx4441, D=>nx2479, CLK=>clk, R=>reset
   );
   ix1647 : oai21 port map ( Y=>nx1646, A0=>nx7009, A1=>nx6705, B0=>nx4073);
   ix2510 : mux21_ni port map ( Y=>nx2509, A0=>nx1678, A1=>
      num_channels_out_2, S0=>nx4115);
   ix1679 : oai21 port map ( Y=>nx1678, A0=>nx4453, A1=>nx6825, B0=>nx4460);
   ix4454 : aoi22 port map ( Y=>nx4453, A0=>mem_data_in(2), A1=>nx6693, B0=>
      nflt_layer_temp_2, B1=>nx1528);
   nflt_layer_total_reg_q_2 : dffr port map ( Q=>nflt_layer_temp_2, QB=>
      nx4459, D=>nx2429, CLK=>clk, R=>reset);
   ix2430 : mux21_ni port map ( Y=>nx2429, A0=>nflt_layer_temp_2, A1=>
      mem_data_in(2), S0=>nx6691);
   ix4461 : aoi22 port map ( Y=>nx4460, A0=>max_num_channels_data_out_2, A1
      =>nx1646, B0=>nx6825, B1=>nx1664);
   ix2500 : oai222 port map ( Y=>nx2499, A0=>nx4465, A1=>nx1594, B0=>nx4459, 
      B1=>nx7019, C0=>nx4059, C1=>nx6821);
   max_num_channels_inst_reg_q_2 : dffr port map ( Q=>
      max_num_channels_data_out_2, QB=>nx4465, D=>nx2499, CLK=>clk, R=>reset
   );
   ix1665 : oai21 port map ( Y=>nx1664, A0=>nx4469, A1=>nx4471, B0=>nx1464);
   reg_num_channels_out_2 : dffr port map ( Q=>num_channels_out_2, QB=>
      nx4469, D=>nx2509, CLK=>clk, R=>reset);
   ix2530 : mux21_ni port map ( Y=>nx2529, A0=>nx1704, A1=>
      num_channels_out_3, S0=>nx4115);
   ix1705 : oai21 port map ( Y=>nx1704, A0=>nx4480, A1=>nx6825, B0=>nx4487);
   ix4481 : aoi22 port map ( Y=>nx4480, A0=>mem_data_in(3), A1=>nx6693, B0=>
      nflt_layer_temp_3, B1=>nx1528);
   nflt_layer_total_reg_q_3 : dffr port map ( Q=>nflt_layer_temp_3, QB=>
      nx4485, D=>nx2419, CLK=>clk, R=>reset);
   ix2420 : mux21_ni port map ( Y=>nx2419, A0=>nflt_layer_temp_3, A1=>
      mem_data_in(3), S0=>nx6691);
   ix4488 : aoi22 port map ( Y=>nx4487, A0=>max_num_channels_data_out_3, A1
      =>nx1646, B0=>nx6825, B1=>nx1690);
   ix2520 : oai222 port map ( Y=>nx2519, A0=>nx4493, A1=>nx1594, B0=>nx4485, 
      B1=>nx7019, C0=>nx4069, C1=>nx6821);
   max_num_channels_inst_reg_q_3 : dffr port map ( Q=>
      max_num_channels_data_out_3, QB=>nx4493, D=>nx2519, CLK=>clk, R=>reset
   );
   ix1691 : oai21 port map ( Y=>nx1690, A0=>nx4497, A1=>nx4499, B0=>nx1463);
   reg_num_channels_out_3 : dffr port map ( Q=>num_channels_out_3, QB=>
      nx4497, D=>nx2529, CLK=>clk, R=>reset);
   num_channels_out_4 : dffr port map ( Q=>OPEN, QB=>nx4503, D=>nx2549, CLK
      =>clk, R=>reset);
   ix2550 : mux21 port map ( Y=>nx2549, A0=>nx4507, A1=>nx4503, S0=>nx4115);
   ix4508 : aoi222 port map ( Y=>nx4507, A0=>max_num_channels_data_out_4, A1
      =>nx1646, B0=>mem_data_in(4), B1=>nx6693, C0=>nx6827, C1=>nx1716);
   ix2540 : oai22 port map ( Y=>nx2539, A0=>nx4513, A1=>nx1594, B0=>nx4515, 
      B1=>nx6821);
   max_num_channels_inst_reg_q_4 : dffr port map ( Q=>
      max_num_channels_data_out_4, QB=>nx4513, D=>nx2539, CLK=>clk, R=>reset
   );
   ix4516 : inv01 port map ( Y=>nx4515, A=>mem_data_in(4));
   ix1717 : oai21 port map ( Y=>nx1716, A0=>nx4503, A1=>nx3989, B0=>nx1409);
   ix4520 : nor03_2x port map ( Y=>nx4519, A0=>nlayers_counter_out_1, A1=>
      nlayers_counter_out_2, A2=>nx4531);
   reg_nlayers_counter_out_1 : dffr port map ( Q=>nlayers_counter_out_1, QB
      =>OPEN, D=>nx2569, CLK=>clk, R=>reset);
   ix2570 : mux21_ni port map ( Y=>nx2569, A0=>nx1768, A1=>
      nlayers_counter_out_1, S0=>nx4009);
   ix4527 : aoi21 port map ( Y=>nx4526, A0=>nlayers_counter_out_1, A1=>
      nlayers_counter_out_0, B0=>nx4535);
   ix2560 : oai32 port map ( Y=>nx2559, A0=>nx4531, A1=>current_state_2, A2
      =>nx6665, B0=>nx4533, B1=>nx4009);
   reg_nlayers_counter_out_0 : dffr port map ( Q=>nlayers_counter_out_0, QB
      =>nx4531, D=>nx2559, CLK=>clk, R=>reset);
   reg_nlayers_counter_out_2 : dffr port map ( Q=>nlayers_counter_out_2, QB
      =>OPEN, D=>nx2579, CLK=>clk, R=>reset);
   ix2580 : mux21_ni port map ( Y=>nx2579, A0=>nx1784, A1=>
      nlayers_counter_out_2, S0=>nx4009);
   ix4544 : xnor2 port map ( Y=>nx4543, A0=>nlayers_counter_out_2, A1=>
      nx4535);
   ix1469 : oai221 port map ( Y=>nx1468, A0=>nx7023, A1=>nx6643, B0=>
      comp_unit_finished, B1=>nx4581, C0=>nx6851);
   reg_current_state_17 : dffr port map ( Q=>OPEN, QB=>nx4553, D=>nx1446, 
      CLK=>nx6633, R=>reset);
   ix1900 : mux21 port map ( Y=>nx1899, A0=>nx4561, A1=>nx4583, S0=>nx6835);
   ix4562 : aoi32 port map ( Y=>nx4561, A0=>nx4563, A1=>ftc_cntrl_reg_out_11, 
      A2=>current_state_21, B0=>ftc_cntrl_reg_out_8, B1=>nx14);
   ix1630 : mux21_ni port map ( Y=>nx1629, A0=>nx332, A1=>
      ftc_cntrl_reg_out_14, S0=>nx6835);
   ix333 : oai22 port map ( Y=>nx332, A0=>nx4563, A1=>nx4571, B0=>nx4565, B1
      =>nx5164);
   ix1843 : oai321 port map ( Y=>nx1842, A0=>nx3959, A1=>nx4579, A2=>nx4581, 
      B0=>nx4583, B1=>nx4673, C0=>nx5162);
   ix4580 : inv01 port map ( Y=>nx4579, A=>comp_unit_finished);
   reg_current_state_19 : dffr port map ( Q=>current_state_19, QB=>nx4581, D
      =>nx1468, CLK=>nx6627, R=>reset);
   ftc_cntrl_reg_reg_q_8 : dffr port map ( Q=>ftc_cntrl_reg_out_8, QB=>
      nx4583, D=>nx1899, CLK=>nx6627, R=>nx6601);
   reg_current_state_13 : dffr port map ( Q=>current_state_13, QB=>OPEN, D=>
      nx300, CLK=>nx6629, R=>reset);
   ix301 : oai22 port map ( Y=>nx300, A0=>nx7029, A1=>nx286, B0=>nx4637, B1
      =>nx6705);
   reg_cntr1_inst_counter_out_4 : dffr port map ( Q=>
      cntr1_inst_counter_out_4, QB=>nx4647, D=>nx1569, CLK=>clk, R=>nx6713);
   ix4602 : nand04 port map ( Y=>nx4601, A0=>cntr1_inst_counter_out_3, A1=>
      cntr1_inst_counter_out_2, A2=>cntr1_inst_counter_out_1, A3=>
      cntr1_inst_counter_out_0);
   reg_cntr1_inst_counter_out_3 : dffr port map ( Q=>
      cntr1_inst_counter_out_3, QB=>OPEN, D=>nx1559, CLK=>clk, R=>nx6713);
   ix215 : xnor2 port map ( Y=>nx214, A0=>cntr1_inst_counter_out_3, A1=>
      nx4609);
   ix4610 : nand03 port map ( Y=>nx4609, A0=>cntr1_inst_counter_out_2, A1=>
      cntr1_inst_counter_out_1, A2=>cntr1_inst_counter_out_0);
   reg_cntr1_inst_counter_out_2 : dffr port map ( Q=>
      cntr1_inst_counter_out_2, QB=>OPEN, D=>nx1549, CLK=>clk, R=>nx6713);
   ix201 : xnor2 port map ( Y=>nx200, A0=>cntr1_inst_counter_out_2, A1=>
      nx4617);
   ix4618 : nand02 port map ( Y=>nx4617, A0=>cntr1_inst_counter_out_1, A1=>
      cntr1_inst_counter_out_0);
   reg_cntr1_inst_counter_out_1 : dffr port map ( Q=>
      cntr1_inst_counter_out_1, QB=>nx4621, D=>nx1539, CLK=>clk, R=>nx6713);
   reg_current_state_10 : dffr port map ( Q=>OPEN, QB=>nx4637, D=>nx152, CLK
      =>nx6629, R=>reset);
   ix153 : or02 port map ( Y=>nx152, A0=>nx1421, A1=>current_state_12);
   reg_current_state_12 : dffr port map ( Q=>current_state_12, QB=>nx4635, D
      =>nx146, CLK=>nx6627, R=>reset);
   ix147 : nand03 port map ( Y=>nx146, A0=>nx4633, A1=>nx6821, A2=>nx4073);
   ix4634 : oai21 port map ( Y=>nx4633, A0=>nx6927, A1=>nx4004, B0=>
      current_state_8);
   ix4639 : oai21 port map ( Y=>nx4638, A0=>cntr1_inst_counter_out_0, A1=>
      cntr1_inst_counter_out_1, B0=>nx4617);
   reg_cntr1_inst_counter_out_0 : dffr port map ( Q=>
      cntr1_inst_counter_out_0, QB=>OPEN, D=>nx1529, CLK=>clk, R=>nx6713);
   ix1530 : xnor2 port map ( Y=>nx1529, A0=>cntr1_inst_counter_out_0, A1=>
      nx7029);
   reg_current_state_11 : dffr port map ( Q=>OPEN, QB=>nx4589, D=>nx6659, 
      CLK=>nx6629, R=>reset);
   cntr1_inst_counter_out_5 : dffr port map ( Q=>OPEN, QB=>nx4655, D=>nx1579, 
      CLK=>clk, R=>nx6713);
   ix287 : nand04 port map ( Y=>nx286, A0=>nx4669, A1=>
      cntr1_inst_counter_out_0, A2=>cntr1_inst_counter_out_3, A3=>nx4663);
   ix4670 : nor03_2x port map ( Y=>nx4669, A0=>nx280, A1=>nx248, A2=>nx246);
   ix2410 : mux21 port map ( Y=>nx2409, A0=>nx4681, A1=>nx4705, S0=>nx6835);
   ix4682 : nand04 port map ( Y=>nx4681, A0=>nx1370, A1=>nx1384, A2=>nx1402, 
      A3=>nx1424);
   reg_cache_width_cntr_counter_out_14 : dffr port map ( Q=>
      cache_width_cntr_counter_out_14, QB=>nx4692, D=>nx2389, CLK=>clk, R=>
      nx6739);
   ix1193 : nand02 port map ( Y=>nx1192, A0=>nx4701, A1=>nx5011);
   ix4702 : aoi21 port map ( Y=>nx4701, A0=>nx4703, A1=>nx6685, B0=>nx6603);
   ftc_cntrl_reg_reg_q_12 : dffr port map ( Q=>ftc_cntrl_reg_out_12, QB=>
      nx4705, D=>nx2409, CLK=>nx6629, R=>nx6601);
   ix307 : or02 port map ( Y=>nx306, A0=>nx1427, A1=>nx6603);
   reg_current_state_14 : dffr port map ( Q=>OPEN, QB=>nx4711, D=>nx306, CLK
      =>nx6629, R=>reset);
   ix1620 : mux21_ni port map ( Y=>nx1619, A0=>cache_height_ended, A1=>
      ftc_cntrl_reg_out_13, S0=>nx6835);
   reg_current_state_15 : dffr port map ( Q=>current_state_15, QB=>nx4725, D
      =>nx1108, CLK=>nx6629, R=>reset);
   ix1109 : oai22 port map ( Y=>nx1108, A0=>nx4151, A1=>nx4153, B0=>nx7033, 
      B1=>nx4723);
   ftc_cntrl_reg_reg_q_13 : dffr port map ( Q=>ftc_cntrl_reg_out_13, QB=>
      nx4723, D=>nx1619, CLK=>nx6629, R=>nx6601);
   ix1139 : nand02 port map ( Y=>nx1138, A0=>nx6977, A1=>nx4751);
   ix1890 : mux21 port map ( Y=>nx1889, A0=>nx4735, A1=>nx4731, S0=>nx6835);
   ix4736 : nand04 port map ( Y=>nx4735, A0=>nx520, A1=>nx534, A2=>nx582, A3
      =>nx702);
   window_width_cntr_counter_out_15 : dffr port map ( Q=>OPEN, QB=>nx4743, D
      =>nx1779, CLK=>clk, R=>nx6723);
   ix349 : nand02 port map ( Y=>nx348, A0=>nx4747, A1=>nx4751);
   ix4748 : aoi22 port map ( Y=>nx4747, A0=>nx6685, A1=>ftc_cntrl_reg_out_13, 
      B0=>current_state_20, B1=>ftc_cntrl_reg_out_12);
   reg_current_state_20 : dffr port map ( Q=>current_state_20, QB=>nx4575, D
      =>nx1842, CLK=>nx6631, R=>reset);
   ix2230 : mux21_ni port map ( Y=>nx2229, A0=>nx1124, A1=>
      ftc_cntrl_reg_out_9, S0=>nx6835);
   ix1125 : oai21 port map ( Y=>nx1124, A0=>nx4759, A1=>nx4761, B0=>nx4747);
   ftc_cntrl_reg_reg_q_9 : dffr port map ( Q=>ftc_cntrl_reg_out_9, QB=>
      nx4759, D=>nx2229, CLK=>nx6631, R=>nx6601);
   ix4762 : aoi21 port map ( Y=>nx4761, A0=>nx6977, A1=>nx1116, B0=>nx6685);
   reg_current_state_16 : dffr port map ( Q=>current_state_16, QB=>nx4765, D
      =>nx1138, CLK=>nx6631, R=>reset);
   reg_window_width_cntr_counter_out_14 : dffr port map ( Q=>
      window_width_cntr_counter_out_14, QB=>nx4770, D=>nx1769, CLK=>clk, R=>
      nx6723);
   ix4777 : nand02 port map ( Y=>nx4776, A0=>
      window_width_cntr_counter_out_13, A1=>nx1432);
   reg_window_width_cntr_counter_out_13 : dffr port map ( Q=>
      window_width_cntr_counter_out_13, QB=>nx4781, D=>nx1759, CLK=>clk, R=>
      nx6723);
   ix4784 : oai21 port map ( Y=>nx4783, A0=>nx1432, A1=>
      window_width_cntr_counter_out_13, B0=>nx4776);
   reg_window_width_cntr_counter_out_12 : dffr port map ( Q=>
      window_width_cntr_counter_out_12, QB=>nx4787, D=>nx1749, CLK=>clk, R=>
      nx6723);
   ix4796 : nand02 port map ( Y=>nx4795, A0=>
      window_width_cntr_counter_out_11, A1=>nx1434);
   reg_window_width_cntr_counter_out_11 : dffr port map ( Q=>
      window_width_cntr_counter_out_11, QB=>nx4801, D=>nx1739, CLK=>clk, R=>
      nx6723);
   ix4804 : oai21 port map ( Y=>nx4803, A0=>nx1434, A1=>
      window_width_cntr_counter_out_11, B0=>nx4795);
   reg_window_width_cntr_counter_out_10 : dffr port map ( Q=>
      window_width_cntr_counter_out_10, QB=>nx4807, D=>nx1729, CLK=>clk, R=>
      nx6723);
   ix4814 : nand02 port map ( Y=>nx4813, A0=>window_width_cntr_counter_out_9, 
      A1=>nx1436);
   reg_window_width_cntr_counter_out_9 : dffr port map ( Q=>
      window_width_cntr_counter_out_9, QB=>nx4819, D=>nx1719, CLK=>clk, R=>
      nx6723);
   ix4822 : oai21 port map ( Y=>nx4821, A0=>nx1436, A1=>
      window_width_cntr_counter_out_9, B0=>nx4813);
   reg_window_width_cntr_counter_out_8 : dffr port map ( Q=>
      window_width_cntr_counter_out_8, QB=>nx4825, D=>nx1709, CLK=>clk, R=>
      nx6725);
   ix4834 : nand02 port map ( Y=>nx4833, A0=>window_width_cntr_counter_out_7, 
      A1=>nx1439);
   reg_window_width_cntr_counter_out_7 : dffr port map ( Q=>
      window_width_cntr_counter_out_7, QB=>nx4839, D=>nx1699, CLK=>clk, R=>
      nx6725);
   ix4842 : oai21 port map ( Y=>nx4841, A0=>nx1439, A1=>
      window_width_cntr_counter_out_7, B0=>nx4833);
   reg_window_width_cntr_counter_out_6 : dffr port map ( Q=>
      window_width_cntr_counter_out_6, QB=>nx4845, D=>nx1689, CLK=>clk, R=>
      nx6725);
   reg_wind_width_count_4 : dffr port map ( Q=>wind_width_count_4, QB=>OPEN, 
      D=>nx2599, CLK=>clk, R=>nx6727);
   ix1881 : xnor2 port map ( Y=>nx1880, A0=>wind_width_count_4, A1=>nx4861);
   ix4862 : nand04 port map ( Y=>nx4861, A0=>wind_width_count_1, A1=>nx6607, 
      A2=>wind_width_count_2, A3=>wind_width_count_3);
   reg_wind_width_count_1 : dffr port map ( Q=>wind_width_count_1, QB=>OPEN, 
      D=>nx1649, CLK=>clk, R=>nx6725);
   ix355 : xor2 port map ( Y=>nx354, A0=>wind_width_count_1, A1=>nx6607);
   reg_wind_width_count_0 : dffr port map ( Q=>wind_width_count_0, QB=>OPEN, 
      D=>nx1639, CLK=>clk, R=>nx6725);
   ix1863 : oai21 port map ( Y=>nx1411, A0=>nx4879, A1=>nx4563, B0=>nx4881);
   reg_current_state_21 : dffr port map ( Q=>current_state_21, QB=>nx4879, D
      =>nx1411, CLK=>nx6631, R=>reset);
   ix4882 : nand03 port map ( Y=>nx4881, A0=>nx1469, A1=>nx4583, A2=>nx4563
   );
   ftc_cntrl_reg_reg_q_11 : dffr port map ( Q=>ftc_cntrl_reg_out_11, QB=>
      nx4731, D=>nx1889, CLK=>nx6631, R=>nx6601);
   ix1879 : oai22 port map ( Y=>nx1429, A0=>ftc_cntrl_reg_out_9, A1=>nx6977, 
      B0=>nx4879, B1=>ftc_cntrl_reg_out_11);
   reg_wind_width_count_2 : dffr port map ( Q=>wind_width_count_2, QB=>OPEN, 
      D=>nx1659, CLK=>clk, R=>nx6725);
   ix363 : xnor2 port map ( Y=>nx362, A0=>wind_width_count_2, A1=>nx4895);
   ix4896 : nand02 port map ( Y=>nx4895, A0=>wind_width_count_1, A1=>nx6609
   );
   reg_wind_width_count_3 : dffr port map ( Q=>wind_width_count_3, QB=>OPEN, 
      D=>nx1669, CLK=>clk, R=>nx6725);
   ix371 : xnor2 port map ( Y=>nx370, A0=>wind_width_count_3, A1=>nx4903);
   ix4904 : nand03 port map ( Y=>nx4903, A0=>wind_width_count_1, A1=>nx6609, 
      A2=>wind_width_count_2);
   reg_window_width_cntr_counter_out_5 : dffr port map ( Q=>
      window_width_cntr_counter_out_5, QB=>nx4911, D=>nx1679, CLK=>clk, R=>
      nx6727);
   ix4914 : oai21 port map ( Y=>nx4913, A0=>nx378, A1=>
      window_width_cntr_counter_out_5, B0=>nx4853);
   ix379 : nor02ii port map ( Y=>nx378, A0=>nx4861, A1=>wind_width_count_4);
   ix575 : xor2 port map ( Y=>nx574, A0=>nx572, A1=>nx6609);
   img_width_reg_q_0 : dffr port map ( Q=>img_width_out_0, QB=>nx4927, D=>
      nx1799, CLK=>clk, R=>reset);
   ix1790 : mux21_ni port map ( Y=>nx1789, A0=>new_width_out_0, A1=>
      mem_data_in(0), S0=>current_state_6);
   new_width_reg_q_0 : dffr port map ( Q=>new_width_out_0, QB=>OPEN, D=>
      nx1789, CLK=>clk, R=>reset);
   ix703 : and04 port map ( Y=>nx702, A0=>nx4941, A1=>nx4957, A2=>nx4977, A3
      =>nx4993);
   ix4942 : xnor2 port map ( Y=>nx4941, A0=>wind_width_count_1, A1=>nx610);
   img_width_reg_q_1 : dffr port map ( Q=>img_width_out_1, QB=>OPEN, D=>
      nx1819, CLK=>clk, R=>reset);
   ix1820 : ao22 port map ( Y=>nx1819, A0=>nx6665, A1=>new_width_out_1, B0=>
      img_width_out_1, B1=>nx4119);
   new_width_reg_q_1 : dffr port map ( Q=>new_width_out_1, QB=>OPEN, D=>
      nx1809, CLK=>clk, R=>reset);
   ix1810 : mux21_ni port map ( Y=>nx1809, A0=>new_width_out_1, A1=>
      mem_data_in(1), S0=>current_state_6);
   ix4958 : xnor2 port map ( Y=>nx4957, A0=>wind_width_count_2, A1=>nx644);
   ix645 : mux21 port map ( Y=>nx644, A0=>nx6641, A1=>nx6839, S0=>nx6977);
   ix4962 : aoi21 port map ( Y=>nx4961, A0=>img_width_out_2, A1=>nx600, B0=>
      nx4975);
   img_width_reg_q_2 : dffs_ni port map ( Q=>img_width_out_2, QB=>OPEN, D=>
      nx1839, CLK=>clk, S=>reset);
   ix1840 : ao221 port map ( Y=>nx1839, A0=>nx6665, A1=>new_width_out_2, B0
      =>img_width_out_2, B1=>nx4119, C0=>nx6695);
   new_width_reg_q_2 : dffr port map ( Q=>new_width_out_2, QB=>OPEN, D=>
      nx1829, CLK=>clk, R=>reset);
   ix1830 : mux21_ni port map ( Y=>nx1829, A0=>new_width_out_2, A1=>
      mem_data_in(2), S0=>current_state_6);
   ix4976 : nor03_2x port map ( Y=>nx4975, A0=>img_width_out_0, A1=>
      img_width_out_1, A2=>img_width_out_2);
   ix4978 : xnor2 port map ( Y=>nx4977, A0=>wind_width_count_3, A1=>nx674);
   ix4982 : xnor2 port map ( Y=>nx4981, A0=>img_width_out_3, A1=>nx4975);
   img_width_reg_q_3 : dffs_ni port map ( Q=>img_width_out_3, QB=>OPEN, D=>
      nx1859, CLK=>clk, S=>reset);
   ix1860 : ao22 port map ( Y=>nx1859, A0=>nx6667, A1=>new_width_out_3, B0=>
      img_width_out_3, B1=>nx4119);
   new_width_reg_q_3 : dffr port map ( Q=>new_width_out_3, QB=>OPEN, D=>
      nx1849, CLK=>clk, R=>reset);
   ix1850 : mux21_ni port map ( Y=>nx1849, A0=>new_width_out_3, A1=>
      mem_data_in(3), S0=>current_state_6);
   ix4994 : xnor2 port map ( Y=>nx4993, A0=>wind_width_count_4, A1=>nx692);
   ix4998 : xnor2 port map ( Y=>nx4997, A0=>img_width_out_4, A1=>nx5009);
   img_width_reg_q_4 : dffs_ni port map ( Q=>img_width_out_4, QB=>OPEN, D=>
      nx1879, CLK=>clk, S=>reset);
   ix1880 : ao22 port map ( Y=>nx1879, A0=>nx6667, A1=>new_width_out_4, B0=>
      img_width_out_4, B1=>nx4119);
   new_width_reg_q_4 : dffr port map ( Q=>new_width_out_4, QB=>OPEN, D=>
      nx1869, CLK=>clk, R=>reset);
   ix1870 : mux21_ni port map ( Y=>nx1869, A0=>new_width_out_4, A1=>
      mem_data_in(4), S0=>current_state_6);
   ix5010 : nor04 port map ( Y=>nx5009, A0=>img_width_out_0, A1=>
      img_width_out_1, A2=>img_width_out_2, A3=>img_width_out_3);
   ix5014 : nand02 port map ( Y=>nx5013, A0=>cache_width_cntr_counter_out_13, 
      A1=>nx1449);
   ix5020 : oai21 port map ( Y=>nx5019, A0=>nx1449, A1=>
      cache_width_cntr_counter_out_13, B0=>nx5013);
   reg_cache_width_cntr_counter_out_12 : dffr port map ( Q=>
      cache_width_cntr_counter_out_12, QB=>nx5023, D=>nx2369, CLK=>clk, R=>
      nx6739);
   ix5032 : nand02 port map ( Y=>nx5031, A0=>cache_width_cntr_counter_out_11, 
      A1=>nx1451);
   ix5038 : oai21 port map ( Y=>nx5037, A0=>nx1451, A1=>
      cache_width_cntr_counter_out_11, B0=>nx5031);
   reg_cache_width_cntr_counter_out_10 : dffr port map ( Q=>
      cache_width_cntr_counter_out_10, QB=>nx5041, D=>nx2349, CLK=>clk, R=>
      nx6739);
   ix5050 : nand02 port map ( Y=>nx5049, A0=>cache_width_cntr_counter_out_9, 
      A1=>nx1454);
   ix5056 : oai21 port map ( Y=>nx5055, A0=>nx1454, A1=>
      cache_width_cntr_counter_out_9, B0=>nx5049);
   reg_cache_width_cntr_counter_out_8 : dffr port map ( Q=>
      cache_width_cntr_counter_out_8, QB=>nx5059, D=>nx2329, CLK=>clk, R=>
      nx6739);
   ix5068 : nand02 port map ( Y=>nx5067, A0=>cache_width_cntr_counter_out_7, 
      A1=>nx1456);
   ix5074 : oai21 port map ( Y=>nx5072, A0=>nx1456, A1=>
      cache_width_cntr_counter_out_7, B0=>nx5067);
   reg_cache_width_cntr_counter_out_6 : dffr port map ( Q=>
      cache_width_cntr_counter_out_6, QB=>nx5077, D=>nx2309, CLK=>clk, R=>
      nx6739);
   reg_cache_width_count_4 : dffr port map ( Q=>cache_width_count_4, QB=>
      OPEN, D=>nx2289, CLK=>clk, R=>nx6741);
   ix1223 : xnor2 port map ( Y=>nx1222, A0=>nx6611, A1=>nx5089);
   ix5090 : nand04 port map ( Y=>nx5089, A0=>cache_width_count_1, A1=>
      cache_width_count_0, A2=>nx6615, A3=>cache_width_count_3);
   reg_cache_width_count_1 : dffr port map ( Q=>cache_width_count_1, QB=>
      OPEN, D=>nx2259, CLK=>clk, R=>nx6739);
   ix1199 : xor2 port map ( Y=>nx1198, A0=>cache_width_count_1, A1=>
      cache_width_count_0);
   reg_cache_width_count_0 : dffr port map ( Q=>cache_width_count_0, QB=>
      OPEN, D=>nx2249, CLK=>clk, R=>nx6739);
   ix5100 : oai21 port map ( Y=>nx5099, A0=>nx4, A1=>nx1152, B0=>
      ftc_cntrl_reg_out_10);
   ix1153 : nor03_2x port map ( Y=>nx1152, A0=>ftc_cntrl_reg_out_12, A1=>
      nx7033, A2=>ftc_cntrl_reg_out_13);
   ix2240 : mux21 port map ( Y=>nx2239, A0=>nx5107, A1=>nx5115, S0=>nx6835);
   ix5108 : aoi221 port map ( Y=>nx5107, A0=>current_state_20, A1=>nx4705, 
      B0=>ftc_cntrl_reg_out_10, B1=>nx1166, C0=>nx1152);
   ix1167 : oai21 port map ( Y=>nx1166, A0=>nx7033, A1=>
      cache_height_count_en, B0=>nx320);
   ix1159 : nor03_2x port map ( Y=>cache_height_count_en, A0=>nx5113, A1=>
      ftc_cntrl_reg_out_13, A2=>nx4705);
   ftc_cntrl_reg_reg_q_10 : dffr port map ( Q=>ftc_cntrl_reg_out_10, QB=>
      nx5115, D=>nx2239, CLK=>nx6631, R=>nx6603);
   reg_cache_width_count_2 : dffr port map ( Q=>cache_width_count_2, QB=>
      OPEN, D=>nx2269, CLK=>clk, R=>nx6741);
   ix1207 : xnor2 port map ( Y=>nx1206, A0=>nx6615, A1=>nx5122);
   ix5123 : nand02 port map ( Y=>nx5122, A0=>cache_width_count_1, A1=>
      cache_width_count_0);
   reg_cache_width_count_3 : dffr port map ( Q=>cache_width_count_3, QB=>
      OPEN, D=>nx2279, CLK=>clk, R=>nx6741);
   ix1215 : xnor2 port map ( Y=>nx1214, A0=>cache_width_count_3, A1=>nx5128
   );
   ix5129 : nand03 port map ( Y=>nx5128, A0=>cache_width_count_1, A1=>
      cache_width_count_0, A2=>nx6617);
   ix5135 : oai21 port map ( Y=>nx5134, A0=>nx1228, A1=>
      cache_width_cntr_counter_out_5, B0=>nx5083);
   ix1229 : nor02ii port map ( Y=>nx1228, A0=>nx5089, A1=>nx6613);
   reg_cache_width_cntr_counter_out_5 : dffr port map ( Q=>
      cache_width_cntr_counter_out_5, QB=>nx5137, D=>nx2299, CLK=>clk, R=>
      nx6741);
   reg_cache_width_cntr_counter_out_7 : dffr port map ( Q=>
      cache_width_cntr_counter_out_7, QB=>nx5140, D=>nx2319, CLK=>clk, R=>
      nx6741);
   reg_cache_width_cntr_counter_out_9 : dffr port map ( Q=>
      cache_width_cntr_counter_out_9, QB=>nx5142, D=>nx2339, CLK=>clk, R=>
      nx6741);
   reg_cache_width_cntr_counter_out_11 : dffr port map ( Q=>
      cache_width_cntr_counter_out_11, QB=>nx5144, D=>nx2359, CLK=>clk, R=>
      nx6741);
   reg_cache_width_cntr_counter_out_13 : dffr port map ( Q=>
      cache_width_cntr_counter_out_13, QB=>nx5146, D=>nx2379, CLK=>clk, R=>
      nx6743);
   cache_width_cntr_counter_out_15 : dffr port map ( Q=>OPEN, QB=>nx5148, D
      =>nx2399, CLK=>clk, R=>nx6743);
   ix1425 : nor04 port map ( Y=>nx1424, A0=>nx1404, A1=>nx1406, A2=>nx1414, 
      A3=>nx1416);
   ix5156 : aoi21 port map ( Y=>nx5155, A0=>img_width_out_1, A1=>
      img_width_out_0, B0=>nx5157);
   ix1407 : xnor2 port map ( Y=>nx1406, A0=>nx6617, A1=>nx6839);
   ix1415 : xnor2 port map ( Y=>nx1414, A0=>cache_width_count_3, A1=>nx4981
   );
   ix1417 : xnor2 port map ( Y=>nx1416, A0=>nx6613, A1=>nx4997);
   ix5163 : aoi43 port map ( Y=>nx5162, A0=>nx4565, A1=>nx6641, A2=>
      current_state_20, A3=>nx4705, B0=>nx4563, B1=>ftc_cntrl_reg_out_11, B2
      =>current_state_21);
   ix5165 : aoi22 port map ( Y=>nx5164, A0=>nx6685, A1=>nx4723, B0=>nx4879, 
      B1=>nx5113);
   ftc_cntrl_reg_reg_q_14 : dffr port map ( Q=>ftc_cntrl_reg_out_14, QB=>
      nx4565, D=>nx1629, CLK=>nx6631, R=>nx6603);
   ix15 : oai221 port map ( Y=>nx14, A0=>nx4575, A1=>ftc_cntrl_reg_out_12, 
      B0=>nx4879, B1=>nx4563, C0=>nx5168);
   ix5169 : nand02 port map ( Y=>nx5168, A0=>nx4879, A1=>nx5011);
   reg_current_state_18 : dffr port map ( Q=>current_state_18, QB=>OPEN, D=>
      nx1452, CLK=>nx6633, R=>reset);
   ix2007 : ao22 port map ( Y=>mem_data_out(5), A0=>comp_unit_data2_in(5), 
      A1=>nx6673, B0=>comp_unit_data1_in(5), B1=>nx6679);
   ix2013 : ao22 port map ( Y=>mem_data_out(6), A0=>comp_unit_data2_in(6), 
      A1=>nx6673, B0=>comp_unit_data1_in(6), B1=>nx6679);
   ix2019 : ao22 port map ( Y=>mem_data_out(7), A0=>comp_unit_data2_in(7), 
      A1=>nx6673, B0=>comp_unit_data1_in(7), B1=>nx6679);
   ix2025 : ao22 port map ( Y=>mem_data_out(8), A0=>comp_unit_data2_in(8), 
      A1=>nx6673, B0=>comp_unit_data1_in(8), B1=>nx6679);
   ix2031 : ao22 port map ( Y=>mem_data_out(9), A0=>comp_unit_data2_in(9), 
      A1=>nx6673, B0=>comp_unit_data1_in(9), B1=>nx6681);
   ix2037 : ao22 port map ( Y=>mem_data_out(10), A0=>comp_unit_data2_in(10), 
      A1=>nx6675, B0=>comp_unit_data1_in(10), B1=>nx6681);
   ix2043 : ao22 port map ( Y=>mem_data_out(11), A0=>comp_unit_data2_in(11), 
      A1=>nx6675, B0=>comp_unit_data1_in(11), B1=>nx6681);
   ix2049 : ao22 port map ( Y=>mem_data_out(12), A0=>comp_unit_data2_in(12), 
      A1=>nx6675, B0=>comp_unit_data1_in(12), B1=>nx6681);
   ix2055 : ao22 port map ( Y=>mem_data_out(13), A0=>comp_unit_data2_in(13), 
      A1=>nx6675, B0=>comp_unit_data1_in(13), B1=>nx6681);
   ix2061 : ao22 port map ( Y=>mem_data_out(14), A0=>comp_unit_data2_in(14), 
      A1=>nx6675, B0=>comp_unit_data1_in(14), B1=>nx6681);
   ix2067 : ao22 port map ( Y=>mem_data_out(15), A0=>comp_unit_data2_in(15), 
      A1=>nx6675, B0=>comp_unit_data1_in(15), B1=>nx6681);
   ix1943 : nand02 port map ( Y=>nx1942, A0=>nx5188, A1=>nx7043);
   ix5189 : nand03 port map ( Y=>nx5188, A0=>nx1419, A1=>nx4519, A2=>nx4017
   );
   ix1741 : nor02_2x port map ( Y=>nx1419, A0=>nx1409, A1=>nx4123);
   reg_current_state_27 : dffr port map ( Q=>current_state_27, QB=>nx5197, D
      =>nx1942, CLK=>nx6633, R=>reset);
   reg_class_cntr_counter_out_0 : dffr port map ( Q=>
      class_cntr_counter_out_0, QB=>nx5194, D=>nx2609, CLK=>nx6633, R=>reset
   );
   reg_class_cntr_counter_out_1 : dffr port map ( Q=>
      class_cntr_counter_out_1, QB=>nx5202, D=>nx2619, CLK=>nx6633, R=>reset
   );
   ix5205 : oai21 port map ( Y=>nx5204, A0=>class_cntr_counter_out_0, A1=>
      class_cntr_counter_out_1, B0=>nx5206);
   reg_class_cntr_counter_out_2 : dffr port map ( Q=>
      class_cntr_counter_out_2, QB=>nx5208, D=>nx2629, CLK=>nx6633, R=>reset
   );
   reg_class_cntr_counter_out_3 : dffr port map ( Q=>
      class_cntr_counter_out_3, QB=>nx5218, D=>nx2639, CLK=>nx6633, R=>reset
   );
   reg_flt_bias1_reg_q_0 : dff port map ( Q=>flt_bias_out_0, QB=>OPEN, D=>
      nx2659, CLK=>clk);
   ix2660 : mux21_ni port map ( Y=>nx2659, A0=>flt_bias_out_0, A1=>
      mem_data_in(0), S0=>nx7091);
   ix2650 : oai21 port map ( Y=>nx2649, A0=>nx7053, A1=>nx152, B0=>nx4635);
   channel_zero_reg_q_0 : dffr port map ( Q=>OPEN, QB=>nx5243, D=>nx2649, 
      CLK=>clk, R=>reset);
   reg_flt_bias1_reg_q_1 : dff port map ( Q=>flt_bias_out_1, QB=>OPEN, D=>
      nx2679, CLK=>clk);
   ix2680 : mux21_ni port map ( Y=>nx2679, A0=>flt_bias_out_1, A1=>
      mem_data_in(1), S0=>nx7091);
   reg_flt_bias1_reg_q_2 : dff port map ( Q=>flt_bias_out_2, QB=>OPEN, D=>
      nx2699, CLK=>clk);
   ix2700 : mux21_ni port map ( Y=>nx2699, A0=>flt_bias_out_2, A1=>
      mem_data_in(2), S0=>nx7091);
   reg_flt_bias1_reg_q_3 : dff port map ( Q=>flt_bias_out_3, QB=>OPEN, D=>
      nx2719, CLK=>clk);
   ix2720 : mux21_ni port map ( Y=>nx2719, A0=>flt_bias_out_3, A1=>
      mem_data_in(3), S0=>nx7091);
   reg_flt_bias1_reg_q_4 : dff port map ( Q=>flt_bias_out_4, QB=>OPEN, D=>
      nx2739, CLK=>clk);
   ix2740 : mux21_ni port map ( Y=>nx2739, A0=>flt_bias_out_4, A1=>
      mem_data_in(4), S0=>nx7091);
   reg_flt_bias1_reg_q_5 : dff port map ( Q=>flt_bias_out_5, QB=>OPEN, D=>
      nx2759, CLK=>clk);
   ix2760 : mux21_ni port map ( Y=>nx2759, A0=>flt_bias_out_5, A1=>
      mem_data_in(5), S0=>nx7091);
   reg_flt_bias1_reg_q_6 : dff port map ( Q=>flt_bias_out_6, QB=>OPEN, D=>
      nx2779, CLK=>clk);
   ix2780 : mux21_ni port map ( Y=>nx2779, A0=>flt_bias_out_6, A1=>
      mem_data_in(6), S0=>nx7093);
   reg_flt_bias1_reg_q_7 : dff port map ( Q=>flt_bias_out_7, QB=>OPEN, D=>
      nx2799, CLK=>clk);
   ix2800 : mux21_ni port map ( Y=>nx2799, A0=>flt_bias_out_7, A1=>
      mem_data_in(7), S0=>nx7093);
   reg_flt_bias1_reg_q_8 : dff port map ( Q=>flt_bias_out_8, QB=>OPEN, D=>
      nx2819, CLK=>clk);
   ix2820 : mux21_ni port map ( Y=>nx2819, A0=>flt_bias_out_8, A1=>
      mem_data_in(8), S0=>nx7093);
   reg_flt_bias1_reg_q_9 : dff port map ( Q=>flt_bias_out_9, QB=>OPEN, D=>
      nx2839, CLK=>clk);
   ix2840 : mux21_ni port map ( Y=>nx2839, A0=>flt_bias_out_9, A1=>
      mem_data_in(9), S0=>nx7093);
   reg_flt_bias1_reg_q_10 : dff port map ( Q=>flt_bias_out_10, QB=>OPEN, D=>
      nx2859, CLK=>clk);
   ix2860 : mux21_ni port map ( Y=>nx2859, A0=>flt_bias_out_10, A1=>
      mem_data_in(10), S0=>nx7093);
   reg_flt_bias1_reg_q_11 : dff port map ( Q=>flt_bias_out_11, QB=>OPEN, D=>
      nx2879, CLK=>clk);
   ix2880 : mux21_ni port map ( Y=>nx2879, A0=>flt_bias_out_11, A1=>
      mem_data_in(11), S0=>nx7093);
   reg_flt_bias1_reg_q_12 : dff port map ( Q=>flt_bias_out_12, QB=>OPEN, D=>
      nx2899, CLK=>clk);
   ix2900 : mux21_ni port map ( Y=>nx2899, A0=>flt_bias_out_12, A1=>
      mem_data_in(12), S0=>nx6993);
   reg_flt_bias1_reg_q_13 : dff port map ( Q=>flt_bias_out_13, QB=>OPEN, D=>
      nx2919, CLK=>clk);
   ix2920 : mux21_ni port map ( Y=>nx2919, A0=>flt_bias_out_13, A1=>
      mem_data_in(13), S0=>nx6993);
   reg_flt_bias1_reg_q_14 : dff port map ( Q=>flt_bias_out_14, QB=>OPEN, D=>
      nx2939, CLK=>clk);
   ix2940 : mux21_ni port map ( Y=>nx2939, A0=>flt_bias_out_14, A1=>
      mem_data_in(14), S0=>nx6993);
   reg_flt_bias1_reg_q_15 : dff port map ( Q=>flt_bias_out_15, QB=>OPEN, D=>
      nx2959, CLK=>clk);
   ix2960 : mux21_ni port map ( Y=>nx2959, A0=>flt_bias_out_15, A1=>
      mem_data_in(15), S0=>nx6993);
   ix5083 : nor03_2x port map ( Y=>max_height_3, A0=>nx4981, A1=>nx6603, A2
      =>nx6687);
   ix5087 : nor03_2x port map ( Y=>max_height_4, A0=>nx4997, A1=>nx6603, A2
      =>nx6687);
   ix4791 : or02 port map ( Y=>cache_rst_actual, A0=>nx6605, A1=>reset);
   ix2980 : mux21 port map ( Y=>nx2979, A0=>nx5330, A1=>nx5334, S0=>nx6837);
   ix5331 : aoi32 port map ( Y=>nx5330, A0=>nx1428, A1=>cache_height_ended, 
      A2=>current_state_20, B0=>ftc_cntrl_reg_out_15, B1=>nx2522);
   ftc_cntrl_reg_reg_q_15 : dffr port map ( Q=>ftc_cntrl_reg_out_15, QB=>
      nx5334, D=>nx2979, CLK=>nx6635, R=>nx6605);
   ix5073 : nand02 port map ( Y=>max_height_0, A0=>nx5379, A1=>
      img_width_out_0);
   ix5079 : nand02 port map ( Y=>max_height_2, A0=>nx5379, A1=>nx6839);
   ix2109 : oai21 port map ( Y=>comp_unit_data1_out(0), A0=>nx6855, A1=>
      nx5383, B0=>nx5386);
   bias1_reg_reg_q_0 : dffr port map ( Q=>OPEN, QB=>nx5383, D=>nx2669, CLK=>
      clk, R=>reset);
   ix5387 : nand02 port map ( Y=>nx5386, A0=>nx2096, A1=>nx6763);
   ix2135 : oai21 port map ( Y=>comp_unit_data1_out(1), A0=>nx6855, A1=>
      nx5390, B0=>nx5393);
   bias1_reg_reg_q_1 : dffr port map ( Q=>OPEN, QB=>nx5390, D=>nx2689, CLK=>
      clk, R=>reset);
   ix5394 : nand02 port map ( Y=>nx5393, A0=>nx2124, A1=>nx6763);
   ix2161 : oai21 port map ( Y=>comp_unit_data1_out(2), A0=>nx6855, A1=>
      nx5396, B0=>nx5399);
   bias1_reg_reg_q_2 : dffr port map ( Q=>OPEN, QB=>nx5396, D=>nx2709, CLK=>
      clk, R=>reset);
   ix5400 : nand02 port map ( Y=>nx5399, A0=>nx2150, A1=>nx6763);
   ix2187 : oai21 port map ( Y=>comp_unit_data1_out(3), A0=>nx6855, A1=>
      nx5402, B0=>nx5405);
   bias1_reg_reg_q_3 : dffr port map ( Q=>OPEN, QB=>nx5402, D=>nx2729, CLK=>
      clk, R=>reset);
   ix5406 : nand02 port map ( Y=>nx5405, A0=>nx2176, A1=>nx6763);
   ix2213 : oai21 port map ( Y=>comp_unit_data1_out(4), A0=>nx6857, A1=>
      nx5408, B0=>nx5411);
   bias1_reg_reg_q_4 : dffr port map ( Q=>OPEN, QB=>nx5408, D=>nx2749, CLK=>
      clk, R=>reset);
   ix5412 : nand02 port map ( Y=>nx5411, A0=>nx2202, A1=>nx6763);
   ix2239 : oai21 port map ( Y=>comp_unit_data1_out(5), A0=>nx6857, A1=>
      nx5414, B0=>nx5417);
   bias1_reg_reg_q_5 : dffr port map ( Q=>OPEN, QB=>nx5414, D=>nx2769, CLK=>
      clk, R=>reset);
   ix5418 : nand02 port map ( Y=>nx5417, A0=>nx2228, A1=>nx6763);
   ix2265 : oai21 port map ( Y=>comp_unit_data1_out(6), A0=>nx6857, A1=>
      nx5420, B0=>nx5423);
   bias1_reg_reg_q_6 : dffr port map ( Q=>OPEN, QB=>nx5420, D=>nx2789, CLK=>
      clk, R=>reset);
   ix5424 : nand02 port map ( Y=>nx5423, A0=>nx2254, A1=>nx6763);
   ix2291 : oai21 port map ( Y=>comp_unit_data1_out(7), A0=>nx6857, A1=>
      nx5426, B0=>nx5429);
   bias1_reg_reg_q_7 : dffr port map ( Q=>OPEN, QB=>nx5426, D=>nx2809, CLK=>
      clk, R=>reset);
   ix5430 : nand02 port map ( Y=>nx5429, A0=>nx2280, A1=>nx6765);
   ix2317 : oai21 port map ( Y=>comp_unit_data1_out(8), A0=>nx6857, A1=>
      nx5432, B0=>nx5435);
   bias1_reg_reg_q_8 : dffr port map ( Q=>OPEN, QB=>nx5432, D=>nx2829, CLK=>
      clk, R=>reset);
   ix5436 : nand02 port map ( Y=>nx5435, A0=>nx2306, A1=>nx6765);
   ix2343 : oai21 port map ( Y=>comp_unit_data1_out(9), A0=>nx6857, A1=>
      nx5438, B0=>nx5441);
   bias1_reg_reg_q_9 : dffr port map ( Q=>OPEN, QB=>nx5438, D=>nx2849, CLK=>
      clk, R=>reset);
   ix5442 : nand02 port map ( Y=>nx5441, A0=>nx2332, A1=>nx6765);
   ix2369 : oai21 port map ( Y=>comp_unit_data1_out(10), A0=>nx6857, A1=>
      nx5444, B0=>nx5447);
   bias1_reg_reg_q_10 : dffr port map ( Q=>OPEN, QB=>nx5444, D=>nx2869, CLK
      =>clk, R=>reset);
   ix5448 : nand02 port map ( Y=>nx5447, A0=>nx2358, A1=>nx6765);
   ix2395 : oai21 port map ( Y=>comp_unit_data1_out(11), A0=>nx6859, A1=>
      nx5450, B0=>nx5453);
   bias1_reg_reg_q_11 : dffr port map ( Q=>OPEN, QB=>nx5450, D=>nx2889, CLK
      =>clk, R=>reset);
   ix5454 : nand02 port map ( Y=>nx5453, A0=>nx2384, A1=>nx6765);
   ix2421 : oai21 port map ( Y=>comp_unit_data1_out(12), A0=>nx6859, A1=>
      nx5456, B0=>nx5459);
   bias1_reg_reg_q_12 : dffr port map ( Q=>OPEN, QB=>nx5456, D=>nx2909, CLK
      =>clk, R=>reset);
   ix5460 : nand02 port map ( Y=>nx5459, A0=>nx2410, A1=>nx6765);
   ix2447 : oai21 port map ( Y=>comp_unit_data1_out(13), A0=>nx6859, A1=>
      nx5462, B0=>nx5465);
   bias1_reg_reg_q_13 : dffr port map ( Q=>OPEN, QB=>nx5462, D=>nx2929, CLK
      =>clk, R=>reset);
   ix5466 : nand02 port map ( Y=>nx5465, A0=>nx2436, A1=>nx6765);
   ix2473 : oai21 port map ( Y=>comp_unit_data1_out(14), A0=>nx6859, A1=>
      nx5468, B0=>nx5471);
   bias1_reg_reg_q_14 : dffr port map ( Q=>OPEN, QB=>nx5468, D=>nx2949, CLK
      =>clk, R=>reset);
   ix5472 : nand02 port map ( Y=>nx5471, A0=>nx2462, A1=>nx6767);
   ix2499 : oai21 port map ( Y=>comp_unit_data1_out(15), A0=>nx6859, A1=>
      nx5474, B0=>nx5477);
   bias1_reg_reg_q_15 : dffr port map ( Q=>OPEN, QB=>nx5474, D=>nx2969, CLK
      =>clk, R=>reset);
   ix5478 : nand02 port map ( Y=>nx5477, A0=>nx2488, A1=>nx6767);
   ix2073 : oai21 port map ( Y=>comp_unit_ready, A0=>nx7023, A1=>nx6705, B0
      =>nx5480);
   ix5481 : aoi21 port map ( Y=>nx5480, A0=>nx6749, A1=>nx7063, B0=>nx6985);
   ix5483 : nand03 port map ( Y=>nx5482, A0=>flt_size_out_0, A1=>nx4143, A2
      =>flt_size_out_1);
   ix4813 : aoi21 port map ( Y=>mem_read_out, A0=>nx5587, A1=>nx5593, B0=>
      reset);
   ix5594 : nor04 port map ( Y=>nx5593, A0=>nx6769, A1=>nx6663, A2=>nx2706, 
      A3=>nx6993);
   ix2707 : nand02 port map ( Y=>nx2706, A0=>nx5596, A1=>nx5598);
   ix5597 : nor04 port map ( Y=>nx5596, A0=>current_state_2, A1=>
      current_state_3, A2=>nx6691, A3=>current_state_5);
   ix4797 : aoi21 port map ( Y=>mem_write_out, A0=>nx6833, A1=>nx6899, B0=>
      reset);
   reg_current_state_28 : dffr port map ( Q=>current_state_28, QB=>OPEN, D=>
      nx1950, CLK=>nx6635, R=>reset);
   ix2739 : nand04 port map ( Y=>mem_addr_out(0), A0=>nx5605, A1=>nx6899, A2
      =>nx5629, A3=>nx5664);
   ix5606 : aoi22 port map ( Y=>nx5605, A0=>nx5607, A1=>nx6651, B0=>
      addr1_data_0, B1=>nx6815);
   ix5608 : oai21 port map ( Y=>nx5607, A0=>class_cntr_counter_out_0, A1=>
      nx6775, B0=>nx5621);
   ix2990 : oai21 port map ( Y=>nx2989, A0=>nx7357, A1=>nx6781, B0=>nx5616);
   reg_write_base_reg_q_0 : dffr port map ( Q=>OPEN, QB=>nx5611, D=>nx2989, 
      CLK=>nx6635, R=>reset);
   ix2581 : nand02 port map ( Y=>nx2580, A0=>nx5614, A1=>nx7009);
   ix5615 : aoi21 port map ( Y=>nx5614, A0=>nx7021, A1=>nx1421, B0=>
      current_state_25);
   ix5617 : nand03 port map ( Y=>nx5616, A0=>nx2582, A1=>nx5619, A2=>nx6781
   );
   ix2583 : nand02 port map ( Y=>nx2582, A0=>nx7357, A1=>nx4423);
   reg_addr1_data_0 : dffr port map ( Q=>addr1_data_0, QB=>OPEN, D=>nx3039, 
      CLK=>clk, R=>reset);
   ix5630 : aoi43 port map ( Y=>nx5629, A0=>nx2620, A1=>nx5636, A2=>nx6985, 
      A3=>nx7053, B0=>nx2680, B1=>nx5662, B2=>nx6769);
   ix2621 : nand02 port map ( Y=>nx2620, A0=>nx7357, A1=>nx5632);
   reg_bias_offset_reg_q_0 : dffr port map ( Q=>bias_offset_data_out_0, QB=>
      nx5632, D=>nx2999, CLK=>clk, R=>reset);
   ix2681 : or02 port map ( Y=>nx2680, A0=>img_addr_offset_0, A1=>
      img_base_addr_0);
   reg_img_addr_offset_0 : dffr port map ( Q=>img_addr_offset_0, QB=>OPEN, D
      =>nx3029, CLK=>clk, R=>nx6807);
   img_base_addr_inst_reg_q_0 : dffs_ni port map ( Q=>img_base_addr_0, QB=>
      OPEN, D=>nx3019, CLK=>clk, S=>reset);
   reg_write_base_prev_reg_q_0 : dffr port map ( Q=>
      write_base_prev_data_out_0, QB=>nx5647, D=>nx3009, CLK=>clk, R=>reset
   );
   ix5652 : nand04 port map ( Y=>nx5651, A0=>nx5653, A1=>nx2640, A2=>nx5657, 
      A3=>nx5659);
   ix5663 : nand02 port map ( Y=>nx5662, A0=>img_base_addr_0, A1=>
      img_addr_offset_0);
   ix5665 : oai221 port map ( Y=>nx5664, A0=>nx6787, A1=>nx6981, B0=>
      write_offset_data_out_0, B1=>nx6775, C0=>nx5667);
   ix2843 : nand03 port map ( Y=>mem_addr_out(1), A0=>nx5670, A1=>nx6899, A2
      =>nx5709);
   ix5671 : aoi22 port map ( Y=>nx5670, A0=>nx2834, A1=>nx6769, B0=>nx2796, 
      B1=>nx6801);
   ix2835 : xor2 port map ( Y=>nx2834, A0=>nx5662, A1=>nx5673);
   img_base_addr_inst_reg_q_1 : dffs_ni port map ( Q=>img_base_addr_1, QB=>
      nx5677, D=>nx3089, CLK=>clk, S=>reset);
   ix5680 : aoi21 port map ( Y=>nx5679, A0=>write_base_prev_data_out_1, A1=>
      write_base_prev_data_out_0, B0=>nx5692);
   reg_write_base_prev_reg_q_1 : dffr port map ( Q=>
      write_base_prev_data_out_1, QB=>OPEN, D=>nx3079, CLK=>clk, R=>reset);
   reg_write_base_reg_q_1 : dffr port map ( Q=>write_base_data_out_1, QB=>
      nx5685, D=>nx3049, CLK=>nx6635, R=>reset);
   ix5688 : xnor2 port map ( Y=>nx5687, A0=>nx5619, A1=>nx5689);
   ix5697 : oai21 port map ( Y=>nx5696, A0=>img_addr_offset_0, A1=>
      img_addr_offset_1, B0=>nx5698);
   ix5699 : nand02 port map ( Y=>nx5698, A0=>img_addr_offset_1, A1=>
      img_addr_offset_0);
   reg_img_addr_offset_1 : dffr port map ( Q=>img_addr_offset_1, QB=>nx5700, 
      D=>nx3099, CLK=>clk, R=>nx6807);
   ix2797 : xor2 port map ( Y=>nx2796, A0=>nx5636, A1=>nx5703);
   reg_bias_offset_reg_q_1 : dffr port map ( Q=>bias_offset_data_out_1, QB=>
      nx5707, D=>nx3069, CLK=>clk, R=>reset);
   ix5710 : aoi222 port map ( Y=>nx5709, A0=>nx6651, A1=>nx2766, B0=>
      addr1_data_1, B1=>nx6815, C0=>nx2752, C1=>nx6795);
   ix2767 : xnor2 port map ( Y=>nx2766, A0=>nx5607, A1=>nx5712);
   ix5713 : xnor2 port map ( Y=>nx5712, A0=>nx5621, A1=>nx5714);
   ix5719 : oai21 port map ( Y=>nx5718, A0=>addr1_data_0, A1=>addr1_data_1, 
      B0=>nx5720);
   ix5721 : nand02 port map ( Y=>nx5720, A0=>addr1_data_1, A1=>addr1_data_0
   );
   reg_addr1_data_1 : dffr port map ( Q=>addr1_data_1, QB=>nx5722, D=>nx3059, 
      CLK=>clk, R=>reset);
   ix2753 : xor2 port map ( Y=>nx2752, A0=>nx5667, A1=>nx5725);
   ix2987 : nand03 port map ( Y=>mem_addr_out(2), A0=>nx5731, A1=>nx6899, A2
      =>nx5773);
   ix5732 : aoi22 port map ( Y=>nx5731, A0=>nx2978, A1=>nx6769, B0=>nx2932, 
      B1=>nx6801);
   ix2979 : xor2 port map ( Y=>nx2978, A0=>nx5734, A1=>nx5737);
   ix5735 : aoi32 port map ( Y=>nx5734, A0=>img_base_addr_0, A1=>
      img_addr_offset_0, A2=>nx2832, B0=>img_addr_offset_1, B1=>
      img_base_addr_1);
   img_base_addr_inst_reg_q_2 : dffs_ni port map ( Q=>img_base_addr_2, QB=>
      nx5758, D=>nx3149, CLK=>clk, S=>reset);
   ix2957 : oai21 port map ( Y=>nx2956, A0=>nx5742, A1=>nx5692, B0=>nx2950);
   reg_write_base_reg_q_2 : dffr port map ( Q=>write_base_data_out_2, QB=>
      nx5747, D=>nx3109, CLK=>nx6635, R=>reset);
   ix5750 : xnor2 port map ( Y=>nx5749, A0=>nx5751, A1=>nx5754);
   reg_write_base_prev_reg_q_2 : dffr port map ( Q=>
      write_base_prev_data_out_2, QB=>nx5742, D=>nx3139, CLK=>clk, R=>reset
   );
   reg_img_addr_offset_2 : dffr port map ( Q=>img_addr_offset_2, QB=>nx5762, 
      D=>nx3159, CLK=>clk, R=>nx6807);
   ix2933 : xor2 port map ( Y=>nx2932, A0=>nx5764, A1=>nx5767);
   ix5765 : aoi32 port map ( Y=>nx5764, A0=>bias_offset_data_out_0, A1=>
      nx6775, A2=>nx2794, B0=>write_base_data_out_1, B1=>
      bias_offset_data_out_1);
   reg_bias_offset_reg_q_2 : dffr port map ( Q=>bias_offset_data_out_2, QB=>
      nx5771, D=>nx3129, CLK=>clk, R=>reset);
   ix5774 : aoi222 port map ( Y=>nx5773, A0=>nx2872, A1=>nx6795, B0=>nx6651, 
      B1=>nx2894, C0=>addr1_data_2, C1=>nx6815);
   ix2873 : xnor2 port map ( Y=>nx2872, A0=>nx2850, A1=>nx5777);
   ix2895 : xnor2 port map ( Y=>nx2894, A0=>nx2760, A1=>nx2886);
   ix2761 : nand02 port map ( Y=>nx2760, A0=>nx5712, A1=>nx5607);
   ix2887 : xnor2 port map ( Y=>nx2886, A0=>nx2882, A1=>nx5783);
   ix2883 : oai22 port map ( Y=>nx2882, A0=>nx5621, A1=>nx5714, B0=>nx5202, 
      B1=>nx7359);
   reg_addr1_data_2 : dffr port map ( Q=>addr1_data_2, QB=>OPEN, D=>nx3119, 
      CLK=>clk, R=>reset);
   ix2905 : xnor2 port map ( Y=>nx2904, A0=>addr1_data_2, A1=>nx5720);
   ix3131 : nand03 port map ( Y=>mem_addr_out(3), A0=>nx5790, A1=>nx6899, A2
      =>nx5826);
   ix5791 : aoi22 port map ( Y=>nx5790, A0=>nx3122, A1=>nx6769, B0=>nx3076, 
      B1=>nx6801);
   ix3123 : xnor2 port map ( Y=>nx3122, A0=>nx3086, A1=>nx5794);
   ix3087 : oai22 port map ( Y=>nx3086, A0=>nx5734, A1=>nx5737, B0=>nx5762, 
      B1=>nx5758);
   ix5795 : xnor2 port map ( Y=>nx5794, A0=>img_base_addr_3, A1=>
      img_addr_offset_3);
   img_base_addr_inst_reg_q_3 : dffr port map ( Q=>img_base_addr_3, QB=>OPEN, 
      D=>nx3209, CLK=>clk, R=>reset);
   ix3101 : xor2 port map ( Y=>nx3100, A0=>write_base_prev_data_out_3, A1=>
      nx5809);
   reg_write_base_prev_reg_q_3 : dffr port map ( Q=>
      write_base_prev_data_out_3, QB=>OPEN, D=>nx3199, CLK=>clk, R=>reset);
   reg_write_base_reg_q_3 : dffs_ni port map ( Q=>write_base_data_out_3, QB
      =>nx5807, D=>nx3169, CLK=>nx6635, S=>reset);
   ix3007 : xnor2 port map ( Y=>nx3006, A0=>nx3002, A1=>nx5805);
   ix5810 : nor03_2x port map ( Y=>nx5809, A0=>write_base_prev_data_out_0, 
      A1=>write_base_prev_data_out_1, A2=>write_base_prev_data_out_2);
   reg_img_addr_offset_3 : dffr port map ( Q=>img_addr_offset_3, QB=>OPEN, D
      =>nx3219, CLK=>clk, R=>nx6807);
   ix3115 : xnor2 port map ( Y=>nx3114, A0=>img_addr_offset_3, A1=>nx5815);
   ix5816 : nand03 port map ( Y=>nx5815, A0=>img_addr_offset_2, A1=>
      img_addr_offset_1, A2=>img_addr_offset_0);
   ix3077 : xnor2 port map ( Y=>nx3076, A0=>nx3066, A1=>nx5820);
   ix3067 : oai22 port map ( Y=>nx3066, A0=>nx5764, A1=>nx5767, B0=>nx7361, 
      B1=>nx5771);
   reg_bias_offset_reg_q_3 : dffr port map ( Q=>bias_offset_data_out_3, QB=>
      OPEN, D=>nx3189, CLK=>clk, R=>reset);
   ix5827 : aoi322 port map ( Y=>nx5826, A0=>nx3032, A1=>nx5838, A2=>nx6651, 
      B0=>addr1_data_3, B1=>nx6815, C0=>nx3016, C1=>nx6795);
   ix3033 : nand02 port map ( Y=>nx3032, A0=>nx5829, A1=>nx5836);
   ix5830 : xnor2 port map ( Y=>nx5829, A0=>nx5831, A1=>nx5834);
   ix5832 : aoi22 port map ( Y=>nx5831, A0=>class_cntr_counter_out_2, A1=>
      write_base_data_out_2, B0=>nx2882, B1=>nx2884);
   ix5837 : nor02_2x port map ( Y=>nx5836, A0=>nx2886, A1=>nx2760);
   reg_addr1_data_3 : dffr port map ( Q=>addr1_data_3, QB=>OPEN, D=>nx3179, 
      CLK=>clk, R=>reset);
   ix3049 : xnor2 port map ( Y=>nx3048, A0=>addr1_data_3, A1=>nx5843);
   ix5844 : nand03 port map ( Y=>nx5843, A0=>addr1_data_2, A1=>addr1_data_1, 
      A2=>addr1_data_0);
   ix3017 : xor2 port map ( Y=>nx3016, A0=>nx5847, A1=>nx5850);
   ix3279 : nand03 port map ( Y=>mem_addr_out(4), A0=>nx5853, A1=>nx6899, A2
      =>nx5901);
   ix5854 : aoi22 port map ( Y=>nx5853, A0=>nx3270, A1=>nx6769, B0=>nx3224, 
      B1=>nx6801);
   ix3271 : xor2 port map ( Y=>nx3270, A0=>nx5856, A1=>nx5859);
   ix5857 : aoi22 port map ( Y=>nx5856, A0=>img_addr_offset_3, A1=>
      img_base_addr_3, B0=>nx3086, B1=>nx3120);
   img_base_addr_inst_reg_q_4 : dffs_ni port map ( Q=>img_base_addr_4, QB=>
      nx5882, D=>nx3269, CLK=>clk, S=>reset);
   ix3249 : oai21 port map ( Y=>nx3248, A0=>nx5864, A1=>nx5879, B0=>nx3242);
   reg_write_base_reg_q_4 : dffr port map ( Q=>write_base_data_out_4, QB=>
      nx5869, D=>nx3229, CLK=>nx6635, R=>reset);
   ix5872 : xnor2 port map ( Y=>nx5871, A0=>nx5873, A1=>nx5876);
   ix5874 : aoi22 port map ( Y=>nx5873, A0=>write_base_data_out_3, A1=>
      new_size_squared_out_3, B0=>nx7323, B1=>nx3004);
   reg_write_base_prev_reg_q_4 : dffr port map ( Q=>OPEN, QB=>nx5864, D=>
      nx3259, CLK=>clk, R=>reset);
   ix5880 : nor04 port map ( Y=>nx5879, A0=>write_base_prev_data_out_0, A1=>
      write_base_prev_data_out_1, A2=>write_base_prev_data_out_2, A3=>
      write_base_prev_data_out_3);
   ix3243 : nand02 port map ( Y=>nx3242, A0=>nx5879, A1=>nx5864);
   ix3263 : aoi21 port map ( Y=>nx3262, A0=>nx5886, A1=>nx5888, B0=>nx3256);
   ix5887 : nand04 port map ( Y=>nx5886, A0=>img_addr_offset_3, A1=>
      img_addr_offset_2, A2=>img_addr_offset_1, A3=>img_addr_offset_0);
   reg_img_addr_offset_4 : dffr port map ( Q=>img_addr_offset_4, QB=>nx5888, 
      D=>nx3279, CLK=>clk, R=>nx6807);
   ix3225 : xor2 port map ( Y=>nx3224, A0=>nx5892, A1=>nx5895);
   ix5893 : aoi22 port map ( Y=>nx5892, A0=>write_base_data_out_3, A1=>
      bias_offset_data_out_3, B0=>nx3066, B1=>nx3074);
   reg_bias_offset_reg_q_4 : dffr port map ( Q=>bias_offset_data_out_4, QB=>
      nx5900, D=>nx3249, CLK=>clk, R=>reset);
   ix829 : aoi21 port map ( Y=>nx828, A0=>nx4265, A1=>nx4257, B0=>nx822);
   ix5902 : aoi222 port map ( Y=>nx5901, A0=>addr1_data_4, A1=>nx6815, B0=>
      nx3160, B1=>nx6795, C0=>nx6651, C1=>nx3186);
   ix3197 : aoi21 port map ( Y=>nx3196, A0=>nx5906, A1=>nx5908, B0=>nx3190);
   ix5907 : nand04 port map ( Y=>nx5906, A0=>addr1_data_3, A1=>addr1_data_2, 
      A2=>addr1_data_1, A3=>addr1_data_0);
   reg_addr1_data_4 : dffr port map ( Q=>addr1_data_4, QB=>nx5908, D=>nx3239, 
      CLK=>clk, R=>reset);
   ix3161 : xnor2 port map ( Y=>nx3160, A0=>nx3138, A1=>nx5913);
   ix3139 : oai22 port map ( Y=>nx3138, A0=>nx7336, A1=>nx5850, B0=>nx4271, 
      B1=>nx5807);
   ix3187 : xor2 port map ( Y=>nx3186, A0=>nx3034, A1=>nx5917);
   ix3035 : nor02_2x port map ( Y=>nx3034, A0=>nx5836, A1=>nx5829);
   ix3171 : oai22 port map ( Y=>nx3170, A0=>nx5831, A1=>nx5834, B0=>nx5218, 
      B1=>nx5807);
   ix3419 : nand03 port map ( Y=>mem_addr_out(5), A0=>nx5921, A1=>nx6899, A2
      =>nx5957);
   ix5922 : aoi22 port map ( Y=>nx5921, A0=>nx3410, A1=>nx6771, B0=>nx3364, 
      B1=>nx6801);
   ix3411 : xnor2 port map ( Y=>nx3410, A0=>nx3374, A1=>nx5925);
   ix3375 : oai22 port map ( Y=>nx3374, A0=>nx5856, A1=>nx5859, B0=>nx5888, 
      B1=>nx5882);
   img_base_addr_inst_reg_q_5 : dffr port map ( Q=>img_base_addr_5, QB=>OPEN, 
      D=>nx3329, CLK=>clk, R=>reset);
   ix3389 : xnor2 port map ( Y=>nx3388, A0=>write_base_prev_data_out_5, A1=>
      nx3242);
   reg_write_base_prev_reg_q_5 : dffr port map ( Q=>
      write_base_prev_data_out_5, QB=>OPEN, D=>nx3319, CLK=>clk, R=>reset);
   reg_write_base_reg_q_5 : dffs_ni port map ( Q=>write_base_data_out_5, QB
      =>nx5938, D=>nx3289, CLK=>nx6637, S=>reset);
   ix3299 : xnor2 port map ( Y=>nx3298, A0=>nx3294, A1=>nx5936);
   ix3295 : oai22 port map ( Y=>nx3294, A0=>nx5873, A1=>nx5876, B0=>nx5869, 
      B1=>nx4391);
   ix5944 : oai21 port map ( Y=>nx5943, A0=>nx3256, A1=>img_addr_offset_5, 
      B0=>nx5945);
   ix5946 : nand02 port map ( Y=>nx5945, A0=>img_addr_offset_5, A1=>nx3256);
   reg_img_addr_offset_5 : dffr port map ( Q=>img_addr_offset_5, QB=>nx5947, 
      D=>nx3339, CLK=>clk, R=>nx6807);
   ix3365 : xnor2 port map ( Y=>nx3364, A0=>nx3354, A1=>nx5951);
   ix3355 : oai22 port map ( Y=>nx3354, A0=>nx5892, A1=>nx5895, B0=>nx5869, 
      B1=>nx5900);
   reg_bias_offset_reg_q_5 : dffr port map ( Q=>bias_offset_data_out_5, QB=>
      nx5955, D=>nx3309, CLK=>clk, R=>reset);
   ix5958 : aoi222 port map ( Y=>nx5957, A0=>addr1_data_5, A1=>nx6815, B0=>
      nx3308, B1=>nx6795, C0=>nx6651, C1=>nx3326);
   ix5962 : oai21 port map ( Y=>nx5961, A0=>nx3190, A1=>addr1_data_5, B0=>
      nx5963);
   ix5964 : nand02 port map ( Y=>nx5963, A0=>addr1_data_5, A1=>nx3190);
   reg_addr1_data_5 : dffr port map ( Q=>addr1_data_5, QB=>nx5965, D=>nx3299, 
      CLK=>clk, R=>reset);
   ix3309 : xor2 port map ( Y=>nx3308, A0=>nx5968, A1=>nx5971);
   ix5969 : aoi22 port map ( Y=>nx5968, A0=>write_offset_data_out_4, A1=>
      write_base_data_out_4, B0=>nx3138, B1=>nx3158);
   ix3327 : xor2 port map ( Y=>nx3326, A0=>nx5974, A1=>nx3318);
   ix5975 : nor02ii port map ( Y=>nx5974, A0=>nx3034, A1=>nx5917);
   ix5978 : nand02 port map ( Y=>nx5977, A0=>write_base_data_out_4, A1=>
      nx3170);
   ix3559 : nand03 port map ( Y=>mem_addr_out(6), A0=>nx5980, A1=>nx6901, A2
      =>nx6026);
   ix5981 : aoi22 port map ( Y=>nx5980, A0=>nx3550, A1=>nx6771, B0=>nx3504, 
      B1=>nx6801);
   ix3551 : xor2 port map ( Y=>nx3550, A0=>nx5983, A1=>nx5986);
   ix5984 : aoi22 port map ( Y=>nx5983, A0=>img_addr_offset_5, A1=>
      img_base_addr_5, B0=>nx3374, B1=>nx3408);
   img_base_addr_inst_reg_q_6 : dffs_ni port map ( Q=>img_base_addr_6, QB=>
      nx6009, D=>nx3389, CLK=>clk, S=>reset);
   ix3529 : oai21 port map ( Y=>nx3528, A0=>nx5991, A1=>nx6006, B0=>nx3522);
   reg_write_base_reg_q_6 : dffs_ni port map ( Q=>write_base_data_out_6, QB
      =>nx5996, D=>nx3349, CLK=>nx6637, S=>reset);
   ix5999 : xnor2 port map ( Y=>nx5998, A0=>nx6000, A1=>nx6003);
   ix6001 : aoi22 port map ( Y=>nx6000, A0=>write_base_data_out_5, A1=>
      new_size_squared_out_5, B0=>nx3294, B1=>nx3296);
   reg_write_base_prev_reg_q_6 : dffr port map ( Q=>OPEN, QB=>nx5991, D=>
      nx3379, CLK=>clk, R=>reset);
   ix6007 : nor02_2x port map ( Y=>nx6006, A0=>nx3242, A1=>
      write_base_prev_data_out_5);
   ix3523 : nand02 port map ( Y=>nx3522, A0=>nx6006, A1=>nx5991);
   ix3543 : aoi21 port map ( Y=>nx3542, A0=>nx5945, A1=>nx6013, B0=>nx3536);
   reg_img_addr_offset_6 : dffr port map ( Q=>img_addr_offset_6, QB=>nx6013, 
      D=>nx3399, CLK=>clk, R=>nx6807);
   ix3505 : xor2 port map ( Y=>nx3504, A0=>nx6017, A1=>nx6020);
   ix6018 : aoi22 port map ( Y=>nx6017, A0=>write_base_data_out_5, A1=>
      bias_offset_data_out_5, B0=>nx3354, B1=>nx3362);
   reg_bias_offset_reg_q_6 : dffr port map ( Q=>bias_offset_data_out_6, QB=>
      nx6025, D=>nx3369, CLK=>clk, R=>reset);
   ix875 : aoi21 port map ( Y=>nx874, A0=>nx4246, A1=>nx4239, B0=>nx868);
   ix6027 : aoi222 port map ( Y=>nx6026, A0=>addr1_data_6, A1=>nx6815, B0=>
      nx3448, B1=>nx6795, C0=>nx6651, C1=>nx3466);
   reg_addr1_data_6 : dffr port map ( Q=>addr1_data_6, QB=>nx6031, D=>nx3359, 
      CLK=>clk, R=>reset);
   ix3449 : xnor2 port map ( Y=>nx3448, A0=>nx3426, A1=>nx6034);
   ix3427 : oai22 port map ( Y=>nx3426, A0=>nx5968, A1=>nx5971, B0=>nx4251, 
      B1=>nx5938);
   ix3467 : xnor2 port map ( Y=>nx3466, A0=>nx6037, A1=>nx6039);
   ix6038 : nor02ii port map ( Y=>nx6037, A0=>nx3318, A1=>nx5974);
   ix6040 : oai21 port map ( Y=>nx6039, A0=>nx3312, A1=>
      write_base_data_out_6, B0=>nx6042);
   ix6043 : nand02 port map ( Y=>nx6042, A0=>write_base_data_out_6, A1=>
      nx3312);
   ix3699 : nand03 port map ( Y=>mem_addr_out(7), A0=>nx6045, A1=>nx6901, A2
      =>nx6081);
   ix6046 : aoi22 port map ( Y=>nx6045, A0=>nx3690, A1=>nx6771, B0=>nx3644, 
      B1=>nx6803);
   ix3691 : xnor2 port map ( Y=>nx3690, A0=>nx3654, A1=>nx6049);
   ix3655 : oai22 port map ( Y=>nx3654, A0=>nx5983, A1=>nx5986, B0=>nx6013, 
      B1=>nx6009);
   img_base_addr_inst_reg_q_7 : dffr port map ( Q=>img_base_addr_7, QB=>OPEN, 
      D=>nx3449, CLK=>clk, R=>reset);
   ix3669 : xnor2 port map ( Y=>nx3668, A0=>write_base_prev_data_out_7, A1=>
      nx3522);
   reg_write_base_prev_reg_q_7 : dffr port map ( Q=>
      write_base_prev_data_out_7, QB=>OPEN, D=>nx3439, CLK=>clk, R=>reset);
   reg_write_base_reg_q_7 : dffr port map ( Q=>write_base_data_out_7, QB=>
      nx6062, D=>nx3409, CLK=>nx6637, R=>reset);
   ix3579 : xnor2 port map ( Y=>nx3578, A0=>nx3574, A1=>nx6060);
   ix3575 : oai22 port map ( Y=>nx3574, A0=>nx6000, A1=>nx6003, B0=>nx5996, 
      B1=>nx4377);
   ix6068 : oai21 port map ( Y=>nx6067, A0=>nx3536, A1=>img_addr_offset_7, 
      B0=>nx6069);
   ix6070 : nand02 port map ( Y=>nx6069, A0=>img_addr_offset_7, A1=>nx3536);
   reg_img_addr_offset_7 : dffr port map ( Q=>img_addr_offset_7, QB=>nx6071, 
      D=>nx3459, CLK=>clk, R=>nx6809);
   ix3645 : xnor2 port map ( Y=>nx3644, A0=>nx3634, A1=>nx6075);
   ix3635 : oai22 port map ( Y=>nx3634, A0=>nx6017, A1=>nx6020, B0=>nx5996, 
      B1=>nx6025);
   reg_bias_offset_reg_q_7 : dffr port map ( Q=>bias_offset_data_out_7, QB=>
      nx6079, D=>nx3429, CLK=>clk, R=>reset);
   ix6082 : aoi222 port map ( Y=>nx6081, A0=>addr1_data_7, A1=>nx6817, B0=>
      nx6653, B1=>nx3606, C0=>nx3588, C1=>nx6795);
   ix6086 : oai21 port map ( Y=>nx6085, A0=>nx3470, A1=>addr1_data_7, B0=>
      nx6088);
   ix6089 : nand02 port map ( Y=>nx6088, A0=>addr1_data_7, A1=>nx3470);
   reg_addr1_data_7 : dffr port map ( Q=>addr1_data_7, QB=>nx6090, D=>nx3419, 
      CLK=>clk, R=>reset);
   ix3607 : xnor2 port map ( Y=>nx3606, A0=>nx3460, A1=>nx3598);
   ix3461 : nand02 port map ( Y=>nx3460, A0=>nx6039, A1=>nx6037);
   ix3599 : aoi21 port map ( Y=>nx3598, A0=>nx6042, A1=>nx6062, B0=>nx3592);
   ix3589 : xor2 port map ( Y=>nx3588, A0=>nx6097, A1=>nx6100);
   ix6098 : aoi22 port map ( Y=>nx6097, A0=>write_offset_data_out_6, A1=>
      write_base_data_out_6, B0=>nx3426, B1=>nx3446);
   ix3839 : nand03 port map ( Y=>mem_addr_out(8), A0=>nx6103, A1=>nx6901, A2
      =>nx6149);
   ix6104 : aoi22 port map ( Y=>nx6103, A0=>nx3830, A1=>nx6771, B0=>nx3784, 
      B1=>nx6803);
   ix3831 : xor2 port map ( Y=>nx3830, A0=>nx6106, A1=>nx6109);
   ix6107 : aoi22 port map ( Y=>nx6106, A0=>img_addr_offset_7, A1=>
      img_base_addr_7, B0=>nx3654, B1=>nx3688);
   img_base_addr_inst_reg_q_8 : dffr port map ( Q=>img_base_addr_8, QB=>
      nx6132, D=>nx3509, CLK=>clk, R=>reset);
   ix3809 : oai21 port map ( Y=>nx3808, A0=>nx6114, A1=>nx6129, B0=>nx3802);
   reg_write_base_reg_q_8 : dffs_ni port map ( Q=>write_base_data_out_8, QB
      =>nx6119, D=>nx3469, CLK=>nx6637, S=>reset);
   ix6122 : xnor2 port map ( Y=>nx6121, A0=>nx6123, A1=>nx6126);
   ix6124 : aoi22 port map ( Y=>nx6123, A0=>write_base_data_out_7, A1=>
      new_size_squared_out_7, B0=>nx3574, B1=>nx3576);
   reg_write_base_prev_reg_q_8 : dffr port map ( Q=>OPEN, QB=>nx6114, D=>
      nx3499, CLK=>clk, R=>reset);
   ix6130 : nor02_2x port map ( Y=>nx6129, A0=>nx3522, A1=>
      write_base_prev_data_out_7);
   ix3803 : nand02 port map ( Y=>nx3802, A0=>nx6129, A1=>nx6114);
   ix3823 : aoi21 port map ( Y=>nx3822, A0=>nx6069, A1=>nx6136, B0=>nx3816);
   reg_img_addr_offset_8 : dffr port map ( Q=>img_addr_offset_8, QB=>nx6136, 
      D=>nx3519, CLK=>clk, R=>nx6809);
   ix3785 : xor2 port map ( Y=>nx3784, A0=>nx6140, A1=>nx6143);
   ix6141 : aoi22 port map ( Y=>nx6140, A0=>write_base_data_out_7, A1=>
      bias_offset_data_out_7, B0=>nx3634, B1=>nx3642);
   reg_bias_offset_reg_q_8 : dffr port map ( Q=>bias_offset_data_out_8, QB=>
      nx6148, D=>nx3489, CLK=>clk, R=>reset);
   ix925 : aoi21 port map ( Y=>nx924, A0=>nx4223, A1=>nx4217, B0=>nx918);
   ix6150 : aoi222 port map ( Y=>nx6149, A0=>addr1_data_8, A1=>nx6817, B0=>
      nx3728, B1=>nx6797, C0=>nx6653, C1=>nx3746);
   reg_addr1_data_8 : dffr port map ( Q=>addr1_data_8, QB=>nx6154, D=>nx3479, 
      CLK=>clk, R=>reset);
   ix3729 : xnor2 port map ( Y=>nx3728, A0=>nx3706, A1=>nx6157);
   ix3707 : oai22 port map ( Y=>nx3706, A0=>nx6097, A1=>nx6100, B0=>nx4229, 
      B1=>nx6062);
   ix3747 : xnor2 port map ( Y=>nx3746, A0=>nx6160, A1=>nx6162);
   ix6161 : nor02_2x port map ( Y=>nx6160, A0=>nx3598, A1=>nx3460);
   ix6163 : oai21 port map ( Y=>nx6162, A0=>nx3592, A1=>
      write_base_data_out_8, B0=>nx6164);
   ix6165 : nand02 port map ( Y=>nx6164, A0=>write_base_data_out_8, A1=>
      nx3592);
   ix3979 : nand03 port map ( Y=>mem_addr_out(9), A0=>nx6167, A1=>nx6901, A2
      =>nx6203);
   ix6168 : aoi22 port map ( Y=>nx6167, A0=>nx3970, A1=>nx6771, B0=>nx3924, 
      B1=>nx6803);
   ix3971 : xnor2 port map ( Y=>nx3970, A0=>nx3934, A1=>nx6171);
   ix3935 : oai22 port map ( Y=>nx3934, A0=>nx6106, A1=>nx6109, B0=>nx6136, 
      B1=>nx6132);
   img_base_addr_inst_reg_q_9 : dffr port map ( Q=>img_base_addr_9, QB=>OPEN, 
      D=>nx3569, CLK=>clk, R=>reset);
   ix3949 : xnor2 port map ( Y=>nx3948, A0=>write_base_prev_data_out_9, A1=>
      nx3802);
   reg_write_base_prev_reg_q_9 : dffr port map ( Q=>
      write_base_prev_data_out_9, QB=>OPEN, D=>nx3559, CLK=>clk, R=>reset);
   reg_write_base_reg_q_9 : dffs_ni port map ( Q=>write_base_data_out_9, QB
      =>nx6184, D=>nx3529, CLK=>nx6637, S=>reset);
   ix3859 : xnor2 port map ( Y=>nx3858, A0=>nx3854, A1=>nx6182);
   ix3855 : oai22 port map ( Y=>nx3854, A0=>nx6123, A1=>nx6126, B0=>nx6119, 
      B1=>nx4363);
   ix6190 : oai21 port map ( Y=>nx6189, A0=>nx3816, A1=>img_addr_offset_9, 
      B0=>nx6191);
   ix6192 : nand02 port map ( Y=>nx6191, A0=>img_addr_offset_9, A1=>nx3816);
   reg_img_addr_offset_9 : dffr port map ( Q=>img_addr_offset_9, QB=>nx6193, 
      D=>nx3579, CLK=>clk, R=>nx6809);
   ix3925 : xnor2 port map ( Y=>nx3924, A0=>nx3914, A1=>nx6197);
   ix3915 : oai22 port map ( Y=>nx3914, A0=>nx6140, A1=>nx6143, B0=>nx6119, 
      B1=>nx6148);
   reg_bias_offset_reg_q_9 : dffr port map ( Q=>bias_offset_data_out_9, QB=>
      nx6201, D=>nx3549, CLK=>clk, R=>reset);
   ix6204 : aoi222 port map ( Y=>nx6203, A0=>addr1_data_9, A1=>nx6817, B0=>
      nx6653, B1=>nx3886, C0=>nx3868, C1=>nx6797);
   ix6208 : oai21 port map ( Y=>nx6207, A0=>nx3750, A1=>addr1_data_9, B0=>
      nx6210);
   ix6211 : nand02 port map ( Y=>nx6210, A0=>addr1_data_9, A1=>nx3750);
   reg_addr1_data_9 : dffr port map ( Q=>addr1_data_9, QB=>nx6212, D=>nx3539, 
      CLK=>clk, R=>reset);
   ix3887 : xnor2 port map ( Y=>nx3886, A0=>nx3740, A1=>nx3878);
   ix3741 : nand02 port map ( Y=>nx3740, A0=>nx6162, A1=>nx6160);
   ix3879 : aoi21 port map ( Y=>nx3878, A0=>nx6164, A1=>nx6184, B0=>nx3872);
   ix3869 : xor2 port map ( Y=>nx3868, A0=>nx6219, A1=>nx6222);
   ix6220 : aoi22 port map ( Y=>nx6219, A0=>write_offset_data_out_8, A1=>
      write_base_data_out_8, B0=>nx3706, B1=>nx3726);
   ix4119 : nand03 port map ( Y=>mem_addr_out(10), A0=>nx6225, A1=>nx6901, 
      A2=>nx6271);
   ix6226 : aoi22 port map ( Y=>nx6225, A0=>nx4110, A1=>nx6771, B0=>nx4064, 
      B1=>nx6803);
   ix4111 : xor2 port map ( Y=>nx4110, A0=>nx6228, A1=>nx6231);
   ix6229 : aoi22 port map ( Y=>nx6228, A0=>img_addr_offset_9, A1=>
      img_base_addr_9, B0=>nx3934, B1=>nx3968);
   img_base_addr_inst_reg_q_10 : dffr port map ( Q=>img_base_addr_10, QB=>
      nx6254, D=>nx3629, CLK=>clk, R=>reset);
   ix4089 : oai21 port map ( Y=>nx4088, A0=>nx6236, A1=>nx6251, B0=>nx4082);
   reg_write_base_reg_q_10 : dffr port map ( Q=>write_base_data_out_10, QB=>
      nx6241, D=>nx3589, CLK=>nx6637, R=>reset);
   ix6244 : xnor2 port map ( Y=>nx6243, A0=>nx6245, A1=>nx6248);
   ix6246 : aoi22 port map ( Y=>nx6245, A0=>write_base_data_out_9, A1=>
      new_size_squared_out_9, B0=>nx3854, B1=>nx3856);
   reg_write_base_prev_reg_q_10 : dffr port map ( Q=>OPEN, QB=>nx6236, D=>
      nx3619, CLK=>clk, R=>reset);
   ix6252 : nor02_2x port map ( Y=>nx6251, A0=>nx3802, A1=>
      write_base_prev_data_out_9);
   ix4083 : nand02 port map ( Y=>nx4082, A0=>nx6251, A1=>nx6236);
   ix4103 : aoi21 port map ( Y=>nx4102, A0=>nx6191, A1=>nx6258, B0=>nx4096);
   reg_img_addr_offset_10 : dffr port map ( Q=>img_addr_offset_10, QB=>
      nx6258, D=>nx3639, CLK=>clk, R=>nx6809);
   ix4065 : xor2 port map ( Y=>nx4064, A0=>nx6262, A1=>nx6265);
   ix6263 : aoi22 port map ( Y=>nx6262, A0=>write_base_data_out_9, A1=>
      bias_offset_data_out_9, B0=>nx3914, B1=>nx3922);
   reg_bias_offset_reg_q_10 : dffr port map ( Q=>bias_offset_data_out_10, QB
      =>nx6270, D=>nx3609, CLK=>clk, R=>reset);
   ix971 : aoi21 port map ( Y=>nx970, A0=>nx4207, A1=>nx4200, B0=>nx964);
   ix6272 : aoi222 port map ( Y=>nx6271, A0=>addr1_data_10, A1=>nx6817, B0=>
      nx4008, B1=>nx6797, C0=>nx6653, C1=>nx4026);
   reg_addr1_data_10 : dffr port map ( Q=>addr1_data_10, QB=>nx6276, D=>
      nx3599, CLK=>clk, R=>reset);
   ix4009 : xnor2 port map ( Y=>nx4008, A0=>nx3986, A1=>nx6279);
   ix3987 : oai22 port map ( Y=>nx3986, A0=>nx6219, A1=>nx6222, B0=>nx4301, 
      B1=>nx6184);
   ix4027 : xnor2 port map ( Y=>nx4026, A0=>nx6282, A1=>nx6284);
   ix6283 : nor02_2x port map ( Y=>nx6282, A0=>nx3878, A1=>nx3740);
   ix6285 : oai21 port map ( Y=>nx6284, A0=>nx3872, A1=>
      write_base_data_out_10, B0=>nx6286);
   ix6287 : nand02 port map ( Y=>nx6286, A0=>write_base_data_out_10, A1=>
      nx3872);
   ix4259 : nand03 port map ( Y=>mem_addr_out(11), A0=>nx6289, A1=>nx6901, 
      A2=>nx6325);
   ix6290 : aoi22 port map ( Y=>nx6289, A0=>nx4250, A1=>nx6771, B0=>nx4204, 
      B1=>nx6803);
   ix4251 : xnor2 port map ( Y=>nx4250, A0=>nx4214, A1=>nx6293);
   ix4215 : oai22 port map ( Y=>nx4214, A0=>nx6228, A1=>nx6231, B0=>nx6258, 
      B1=>nx6254);
   img_base_addr_inst_reg_q_11 : dffs_ni port map ( Q=>img_base_addr_11, QB
      =>OPEN, D=>nx3689, CLK=>clk, S=>reset);
   ix4229 : xnor2 port map ( Y=>nx4228, A0=>write_base_prev_data_out_11, A1
      =>nx4082);
   reg_write_base_prev_reg_q_11 : dffr port map ( Q=>
      write_base_prev_data_out_11, QB=>OPEN, D=>nx3679, CLK=>clk, R=>reset);
   reg_write_base_reg_q_11 : dffs_ni port map ( Q=>write_base_data_out_11, 
      QB=>nx6306, D=>nx3649, CLK=>nx6637, S=>reset);
   ix4139 : xnor2 port map ( Y=>nx4138, A0=>nx4134, A1=>nx6304);
   ix4135 : oai22 port map ( Y=>nx4134, A0=>nx6245, A1=>nx6248, B0=>nx6241, 
      B1=>nx4349);
   ix6312 : oai21 port map ( Y=>nx6311, A0=>nx4096, A1=>img_addr_offset_11, 
      B0=>nx6313);
   ix6314 : nand02 port map ( Y=>nx6313, A0=>img_addr_offset_11, A1=>nx4096
   );
   reg_img_addr_offset_11 : dffr port map ( Q=>img_addr_offset_11, QB=>
      nx6315, D=>nx3699, CLK=>clk, R=>nx6809);
   ix4205 : xnor2 port map ( Y=>nx4204, A0=>nx4194, A1=>nx6319);
   ix4195 : oai22 port map ( Y=>nx4194, A0=>nx6262, A1=>nx6265, B0=>nx6241, 
      B1=>nx6270);
   reg_bias_offset_reg_q_11 : dffr port map ( Q=>bias_offset_data_out_11, QB
      =>nx6323, D=>nx3669, CLK=>clk, R=>reset);
   ix6326 : aoi222 port map ( Y=>nx6325, A0=>addr1_data_11, A1=>nx6817, B0=>
      nx6653, B1=>nx4166, C0=>nx4148, C1=>nx6797);
   ix6330 : oai21 port map ( Y=>nx6329, A0=>nx4030, A1=>addr1_data_11, B0=>
      nx6332);
   ix6333 : nand02 port map ( Y=>nx6332, A0=>addr1_data_11, A1=>nx4030);
   reg_addr1_data_11 : dffr port map ( Q=>addr1_data_11, QB=>nx6334, D=>
      nx3659, CLK=>clk, R=>reset);
   ix4167 : xnor2 port map ( Y=>nx4166, A0=>nx4020, A1=>nx4158);
   ix4021 : nand02 port map ( Y=>nx4020, A0=>nx6284, A1=>nx6282);
   ix4159 : aoi21 port map ( Y=>nx4158, A0=>nx6286, A1=>nx6306, B0=>nx4152);
   ix4149 : xor2 port map ( Y=>nx4148, A0=>nx6341, A1=>nx6344);
   ix6342 : aoi22 port map ( Y=>nx6341, A0=>write_offset_data_out_10, A1=>
      write_base_data_out_10, B0=>nx3986, B1=>nx4006);
   ix4399 : nand03 port map ( Y=>mem_addr_out(12), A0=>nx6347, A1=>nx6901, 
      A2=>nx6393);
   ix6348 : aoi22 port map ( Y=>nx6347, A0=>nx4390, A1=>nx6773, B0=>nx4344, 
      B1=>nx6803);
   ix4391 : xor2 port map ( Y=>nx4390, A0=>nx6350, A1=>nx6353);
   ix6351 : aoi22 port map ( Y=>nx6350, A0=>img_addr_offset_11, A1=>
      img_base_addr_11, B0=>nx4214, B1=>nx4248);
   img_base_addr_inst_reg_q_12 : dffs_ni port map ( Q=>img_base_addr_12, QB
      =>nx6376, D=>nx3749, CLK=>clk, S=>reset);
   ix4369 : oai21 port map ( Y=>nx4368, A0=>nx6358, A1=>nx6373, B0=>nx4362);
   reg_write_base_reg_q_12 : dffs_ni port map ( Q=>write_base_data_out_12, 
      QB=>nx6363, D=>nx3709, CLK=>nx6639, S=>reset);
   ix6366 : xnor2 port map ( Y=>nx6365, A0=>nx7445, A1=>nx6370);
   ix6368 : aoi22 port map ( Y=>nx6367, A0=>write_base_data_out_11, A1=>
      new_size_squared_out_11, B0=>nx4134, B1=>nx4136);
   reg_write_base_prev_reg_q_12 : dffr port map ( Q=>OPEN, QB=>nx6358, D=>
      nx3739, CLK=>clk, R=>reset);
   ix6374 : nor02_2x port map ( Y=>nx6373, A0=>nx4082, A1=>
      write_base_prev_data_out_11);
   ix4363 : nand02 port map ( Y=>nx4362, A0=>nx6373, A1=>nx6358);
   ix4383 : aoi21 port map ( Y=>nx4382, A0=>nx6313, A1=>nx6380, B0=>nx4376);
   reg_img_addr_offset_12 : dffr port map ( Q=>img_addr_offset_12, QB=>
      nx6380, D=>nx3759, CLK=>clk, R=>nx6809);
   ix4345 : xor2 port map ( Y=>nx4344, A0=>nx6384, A1=>nx6387);
   ix6385 : aoi22 port map ( Y=>nx6384, A0=>write_base_data_out_11, A1=>
      bias_offset_data_out_11, B0=>nx4194, B1=>nx4202);
   reg_bias_offset_reg_q_12 : dffr port map ( Q=>bias_offset_data_out_12, QB
      =>nx6392, D=>nx3729, CLK=>clk, R=>reset);
   ix1019 : aoi21 port map ( Y=>nx1018, A0=>nx4191, A1=>nx4183, B0=>nx1012);
   ix6394 : aoi222 port map ( Y=>nx6393, A0=>addr1_data_12, A1=>nx6817, B0=>
      nx6653, B1=>nx4306, C0=>nx4288, C1=>nx6797);
   reg_addr1_data_12 : dffr port map ( Q=>addr1_data_12, QB=>nx6398, D=>
      nx3719, CLK=>clk, R=>reset);
   ix4307 : xnor2 port map ( Y=>nx4306, A0=>nx6400, A1=>nx6402);
   ix6401 : nor02_2x port map ( Y=>nx6400, A0=>nx4158, A1=>nx4020);
   ix6403 : oai21 port map ( Y=>nx6402, A0=>nx4152, A1=>
      write_base_data_out_12, B0=>nx6404);
   ix6405 : nand02 port map ( Y=>nx6404, A0=>write_base_data_out_12, A1=>
      nx4152);
   ix4289 : xnor2 port map ( Y=>nx4288, A0=>nx4266, A1=>nx6408);
   ix4267 : oai22 port map ( Y=>nx4266, A0=>nx6341, A1=>nx6344, B0=>nx4303, 
      B1=>nx6306);
   ix4539 : nand03 port map ( Y=>mem_addr_out(13), A0=>nx6411, A1=>nx6903, 
      A2=>nx6447);
   ix6412 : aoi22 port map ( Y=>nx6411, A0=>nx4530, A1=>nx6773, B0=>nx4484, 
      B1=>nx6803);
   ix4531 : xnor2 port map ( Y=>nx4530, A0=>nx4494, A1=>nx6415);
   ix4495 : oai22 port map ( Y=>nx4494, A0=>nx6350, A1=>nx6353, B0=>nx6380, 
      B1=>nx6376);
   img_base_addr_inst_reg_q_13 : dffr port map ( Q=>img_base_addr_13, QB=>
      OPEN, D=>nx3809, CLK=>clk, R=>reset);
   ix4509 : xnor2 port map ( Y=>nx4508, A0=>write_base_prev_data_out_13, A1
      =>nx4362);
   reg_write_base_prev_reg_q_13 : dffr port map ( Q=>
      write_base_prev_data_out_13, QB=>OPEN, D=>nx3799, CLK=>clk, R=>reset);
   reg_write_base_reg_q_13 : dffr port map ( Q=>write_base_data_out_13, QB=>
      nx6428, D=>nx3769, CLK=>nx6639, R=>reset);
   ix4419 : xnor2 port map ( Y=>nx4418, A0=>nx4414, A1=>nx6426);
   ix6434 : oai21 port map ( Y=>nx6433, A0=>nx4376, A1=>img_addr_offset_13, 
      B0=>nx6435);
   ix6436 : nand02 port map ( Y=>nx6435, A0=>img_addr_offset_13, A1=>nx4376
   );
   reg_img_addr_offset_13 : dffr port map ( Q=>img_addr_offset_13, QB=>
      nx6437, D=>nx3819, CLK=>clk, R=>nx6809);
   ix4485 : xnor2 port map ( Y=>nx4484, A0=>nx4474, A1=>nx6441);
   ix4475 : oai22 port map ( Y=>nx4474, A0=>nx6384, A1=>nx6387, B0=>nx7363, 
      B1=>nx6392);
   reg_bias_offset_reg_q_13 : dffr port map ( Q=>bias_offset_data_out_13, QB
      =>nx6445, D=>nx3789, CLK=>clk, R=>reset);
   ix6448 : aoi222 port map ( Y=>nx6447, A0=>addr1_data_13, A1=>nx6817, B0=>
      nx6653, B1=>nx4446, C0=>nx4428, C1=>nx6797);
   ix6452 : oai21 port map ( Y=>nx6451, A0=>nx4310, A1=>addr1_data_13, B0=>
      nx6454);
   ix6455 : nand02 port map ( Y=>nx6454, A0=>addr1_data_13, A1=>nx4310);
   reg_addr1_data_13 : dffr port map ( Q=>addr1_data_13, QB=>nx6456, D=>
      nx3779, CLK=>clk, R=>reset);
   ix4447 : xnor2 port map ( Y=>nx4446, A0=>nx4300, A1=>nx4438);
   ix4301 : nand02 port map ( Y=>nx4300, A0=>nx6402, A1=>nx6400);
   ix4439 : aoi21 port map ( Y=>nx4438, A0=>nx6404, A1=>nx6428, B0=>nx4432);
   ix4429 : xor2 port map ( Y=>nx4428, A0=>nx6463, A1=>nx6466);
   ix6464 : aoi22 port map ( Y=>nx6463, A0=>write_offset_data_out_12, A1=>
      write_base_data_out_12, B0=>nx4266, B1=>nx4286);
   ix4679 : nand03 port map ( Y=>mem_addr_out(14), A0=>nx6469, A1=>nx6903, 
      A2=>nx6511);
   ix6470 : aoi22 port map ( Y=>nx6469, A0=>nx4670, A1=>nx6773, B0=>nx4624, 
      B1=>nx2626);
   ix4671 : xor2 port map ( Y=>nx4670, A0=>nx6472, A1=>nx6475);
   ix6473 : aoi22 port map ( Y=>nx6472, A0=>img_addr_offset_13, A1=>
      img_base_addr_13, B0=>nx4494, B1=>nx4528);
   img_base_addr_inst_reg_q_14 : dffr port map ( Q=>img_base_addr_14, QB=>
      nx6496, D=>nx3869, CLK=>clk, R=>reset);
   reg_write_base_prev_reg_q_14 : dffr port map ( Q=>OPEN, QB=>nx6493, D=>
      nx3859, CLK=>clk, R=>reset);
   reg_write_base_reg_q_14 : dffr port map ( Q=>write_base_data_out_14, QB=>
      nx6484, D=>nx3829, CLK=>nx6639, R=>reset);
   ix6487 : xnor2 port map ( Y=>nx6486, A0=>nx6488, A1=>nx6491);
   ix6495 : nor02_2x port map ( Y=>nx6494, A0=>nx4362, A1=>
      write_base_prev_data_out_13);
   reg_img_addr_offset_14 : dffr port map ( Q=>img_addr_offset_14, QB=>
      nx6500, D=>nx3879, CLK=>clk, R=>nx6811);
   ix4625 : xor2 port map ( Y=>nx4624, A0=>nx6502, A1=>nx6505);
   ix6503 : aoi22 port map ( Y=>nx6502, A0=>write_base_data_out_13, A1=>
      bias_offset_data_out_13, B0=>nx4474, B1=>nx4482);
   reg_bias_offset_reg_q_14 : dffr port map ( Q=>bias_offset_data_out_14, QB
      =>nx6510, D=>nx3849, CLK=>clk, R=>reset);
   ix6512 : aoi222 port map ( Y=>nx6511, A0=>addr1_data_14, A1=>nx6819, B0=>
      nx6655, B1=>nx4586, C0=>nx4568, C1=>nx6797);
   reg_addr1_data_14 : dffr port map ( Q=>addr1_data_14, QB=>nx6516, D=>
      nx3839, CLK=>clk, R=>reset);
   ix4587 : xnor2 port map ( Y=>nx4586, A0=>nx6518, A1=>nx6520);
   ix6519 : nor02_2x port map ( Y=>nx6518, A0=>nx4438, A1=>nx4300);
   ix4569 : xnor2 port map ( Y=>nx4568, A0=>nx4546, A1=>nx6524);
   ix4547 : oai22 port map ( Y=>nx4546, A0=>nx6463, A1=>nx6466, B0=>nx4305, 
      B1=>nx6428);
   ix4789 : nand03 port map ( Y=>mem_addr_out(15), A0=>nx6527, A1=>nx6903, 
      A2=>nx6560);
   ix6528 : aoi22 port map ( Y=>nx6527, A0=>nx4746, A1=>nx6655, B0=>nx4780, 
      B1=>nx6773);
   ix4747 : xnor2 port map ( Y=>nx4746, A0=>nx4580, A1=>nx4744);
   ix4581 : nand02 port map ( Y=>nx4580, A0=>nx6520, A1=>nx6518);
   ix4745 : xnor2 port map ( Y=>nx4744, A0=>nx6532, A1=>
      write_base_data_out_15);
   ix6533 : nand02 port map ( Y=>nx6532, A0=>write_base_data_out_14, A1=>
      nx4432);
   reg_write_base_reg_q_15 : dffs_ni port map ( Q=>write_base_data_out_15, 
      QB=>OPEN, D=>nx3899, CLK=>nx6639, S=>reset);
   ix4781 : xnor2 port map ( Y=>nx4780, A0=>nx4756, A1=>nx6543);
   ix4757 : oai22 port map ( Y=>nx4756, A0=>nx6472, A1=>nx6475, B0=>nx6500, 
      B1=>nx6496);
   img_base_addr_inst_reg_q_15 : dffs_ni port map ( Q=>img_base_addr_15, QB
      =>OPEN, D=>nx3929, CLK=>clk, S=>reset);
   ix4765 : xnor2 port map ( Y=>nx4764, A0=>write_base_prev_data_out_15, A1
      =>nx4642);
   reg_write_base_prev_reg_q_15 : dffr port map ( Q=>
      write_base_prev_data_out_15, QB=>OPEN, D=>nx3919, CLK=>clk, R=>reset);
   ix4643 : nand02 port map ( Y=>nx4642, A0=>nx6494, A1=>nx6493);
   img_addr_offset_15 : dffr port map ( Q=>OPEN, QB=>nx6558, D=>nx3939, CLK
      =>clk, R=>nx6811);
   ix6561 : aoi222 port map ( Y=>nx6560, A0=>nx4736, A1=>nx6799, B0=>
      addr1_data_15, B1=>nx6819, C0=>nx4714, C1=>nx2626);
   ix4737 : xnor2 port map ( Y=>nx4736, A0=>nx6563, A1=>nx4734);
   ix6564 : aoi22 port map ( Y=>nx6563, A0=>write_offset_data_out_14, A1=>
      write_base_data_out_14, B0=>nx4546, B1=>nx4566);
   reg_addr1_data_15 : dffr port map ( Q=>addr1_data_15, QB=>nx6572, D=>
      nx3909, CLK=>clk, R=>reset);
   ix4715 : xnor2 port map ( Y=>nx4714, A0=>nx4686, A1=>nx6576);
   ix4687 : oai22 port map ( Y=>nx4686, A0=>nx6502, A1=>nx6505, B0=>nx7365, 
      B1=>nx6510);
   reg_bias_offset_reg_q_15 : dffr port map ( Q=>bias_offset_data_out_15, QB
      =>nx6580, D=>nx3889, CLK=>clk, R=>reset);
   ix1965 : inv01 port map ( Y=>mem_data_out(0), A=>nx6583);
   ix6584 : aoi222 port map ( Y=>nx6583, A0=>comp_unit_data2_in(0), A1=>
      nx6675, B0=>comp_unit_data1_in(0), B1=>nx6683, C0=>argmax_data_in(0), 
      C1=>current_state_28);
   ix1975 : inv01 port map ( Y=>mem_data_out(1), A=>nx6586);
   ix6587 : aoi222 port map ( Y=>nx6586, A0=>comp_unit_data2_in(1), A1=>
      nx6677, B0=>comp_unit_data1_in(1), B1=>nx6683, C0=>argmax_data_in(1), 
      C1=>current_state_28);
   ix1985 : inv01 port map ( Y=>mem_data_out(2), A=>nx6589);
   ix6590 : aoi222 port map ( Y=>nx6589, A0=>comp_unit_data2_in(2), A1=>
      nx6677, B0=>comp_unit_data1_in(2), B1=>nx6683, C0=>argmax_data_in(2), 
      C1=>current_state_28);
   ix1995 : inv01 port map ( Y=>mem_data_out(3), A=>nx6592);
   ix6593 : aoi222 port map ( Y=>nx6592, A0=>comp_unit_data2_in(3), A1=>
      nx6677, B0=>comp_unit_data1_in(3), B1=>nx6683, C0=>argmax_data_in(3), 
      C1=>current_state_28);
   ix4567 : inv01 port map ( Y=>nx4566, A=>nx6524);
   ix4529 : inv01 port map ( Y=>nx4528, A=>nx6415);
   ix4483 : inv01 port map ( Y=>nx4482, A=>nx6441);
   ix4287 : inv01 port map ( Y=>nx4286, A=>nx6408);
   ix4249 : inv01 port map ( Y=>nx4248, A=>nx6293);
   ix4203 : inv01 port map ( Y=>nx4202, A=>nx6319);
   ix4137 : inv01 port map ( Y=>nx4136, A=>nx6304);
   ix4007 : inv01 port map ( Y=>nx4006, A=>nx6279);
   ix3969 : inv01 port map ( Y=>nx3968, A=>nx6171);
   ix3923 : inv01 port map ( Y=>nx3922, A=>nx6197);
   ix3857 : inv01 port map ( Y=>nx3856, A=>nx6182);
   ix3727 : inv01 port map ( Y=>nx3726, A=>nx6157);
   ix3689 : inv01 port map ( Y=>nx3688, A=>nx6049);
   ix3643 : inv01 port map ( Y=>nx3642, A=>nx6075);
   ix3577 : inv01 port map ( Y=>nx3576, A=>nx6060);
   ix3447 : inv01 port map ( Y=>nx3446, A=>nx6034);
   ix3409 : inv01 port map ( Y=>nx3408, A=>nx5925);
   ix3363 : inv01 port map ( Y=>nx3362, A=>nx5951);
   ix3297 : inv01 port map ( Y=>nx3296, A=>nx5936);
   ix3159 : inv01 port map ( Y=>nx3158, A=>nx5913);
   ix3121 : inv01 port map ( Y=>nx3120, A=>nx5794);
   ix3075 : inv01 port map ( Y=>nx3074, A=>nx5820);
   ix5839 : inv01 port map ( Y=>nx5838, A=>nx3034);
   ix3005 : inv01 port map ( Y=>nx3004, A=>nx5805);
   ix2951 : inv01 port map ( Y=>nx2950, A=>nx5809);
   ix2885 : inv01 port map ( Y=>nx2884, A=>nx5783);
   ix2833 : inv01 port map ( Y=>nx2832, A=>nx5673);
   ix2795 : inv01 port map ( Y=>nx2794, A=>nx5703);
   ix5502 : inv01 port map ( Y=>nx5501, A=>nx2502);
   ix1685 : inv01 port map ( Y=>nx1464, A=>nx4499);
   ix1711 : inv01 port map ( Y=>nx1463, A=>nx3989);
   ix1529 : inv01 port map ( Y=>nx1528, A=>nx4080);
   ix1807 : inv01 port map ( Y=>nx1461, A=>nx4009);
   ix1429 : inv01 port map ( Y=>nx1428, A=>nx4681);
   ix4704 : inv01 port map ( Y=>nx4703, A=>nx1152);
   ix751 : inv01 port map ( Y=>nx750, A=>nx4295);
   ix607 : inv01 port map ( Y=>nx606, A=>nx5155);
   ix601 : inv01 port map ( Y=>nx600, A=>nx5157);
   ix4884 : inv01 port map ( Y=>nx4883, A=>nx546);
   ix321 : inv01 port map ( Y=>nx320, A=>nx5113);
   ix6598 : inv01 port map ( Y=>nx6599, A=>current_state_13);
   ix6600 : inv02 port map ( Y=>nx6601, A=>nx6599);
   ix6602 : inv02 port map ( Y=>nx6603, A=>nx6599);
   ix6604 : inv02 port map ( Y=>nx6605, A=>nx6599);
   ix6606 : buf02 port map ( Y=>nx6607, A=>wind_width_count_0);
   ix6608 : buf02 port map ( Y=>nx6609, A=>wind_width_count_0);
   ix6610 : buf02 port map ( Y=>nx6611, A=>cache_width_count_4);
   ix6612 : buf02 port map ( Y=>nx6613, A=>cache_width_count_4);
   ix6614 : buf02 port map ( Y=>nx6615, A=>cache_width_count_2);
   ix6616 : buf02 port map ( Y=>nx6617, A=>cache_width_count_2);
   ix6618 : inv02 port map ( Y=>nx6619, A=>clk);
   ix6620 : inv02 port map ( Y=>nx6621, A=>clk);
   ix6622 : inv02 port map ( Y=>nx6623, A=>clk);
   ix6624 : inv02 port map ( Y=>nx6625, A=>clk);
   ix6626 : inv02 port map ( Y=>nx6627, A=>clk);
   ix6628 : inv02 port map ( Y=>nx6629, A=>clk);
   ix6630 : inv02 port map ( Y=>nx6631, A=>clk);
   ix6632 : inv02 port map ( Y=>nx6633, A=>clk);
   ix6634 : inv02 port map ( Y=>nx6635, A=>clk);
   ix6636 : inv02 port map ( Y=>nx6637, A=>clk);
   ix6638 : inv02 port map ( Y=>nx6639, A=>clk);
   ix6640 : inv02 port map ( Y=>nx6641, A=>nx7294);
   ix6642 : inv02 port map ( Y=>nx6643, A=>nx7294);
   ix6650 : inv02 port map ( Y=>nx6651, A=>nx7043);
   ix6652 : inv02 port map ( Y=>nx6653, A=>nx7043);
   ix6654 : inv02 port map ( Y=>nx6655, A=>nx7043);
   ix6656 : inv01 port map ( Y=>nx6657, A=>nx7293);
   ix6658 : inv02 port map ( Y=>nx6659, A=>nx7077);
   ix6662 : inv02 port map ( Y=>nx6663, A=>nx7077);
   ix6664 : inv02 port map ( Y=>nx6665, A=>nx3981);
   ix6666 : inv02 port map ( Y=>nx6667, A=>nx7009);
   ix6672 : inv02 port map ( Y=>nx6673, A=>nx4149);
   ix6674 : inv02 port map ( Y=>nx6675, A=>nx4149);
   ix6676 : inv02 port map ( Y=>nx6677, A=>nx4149);
   ix6678 : inv02 port map ( Y=>nx6679, A=>nx4129);
   ix6680 : inv02 port map ( Y=>nx6681, A=>nx4129);
   ix6682 : inv02 port map ( Y=>nx6683, A=>nx4129);
   ix6684 : inv02 port map ( Y=>nx6685, A=>nx4711);
   ix6686 : inv02 port map ( Y=>nx6687, A=>nx7033);
   ix6688 : buf02 port map ( Y=>nx6689, A=>current_state_4);
   ix6690 : buf02 port map ( Y=>nx6691, A=>current_state_4);
   ix6692 : inv02 port map ( Y=>nx6693, A=>nx6823);
   ix6694 : inv02 port map ( Y=>nx6695, A=>nx6823);
   ix6698 : inv02 port map ( Y=>nx6699, A=>nx7081);
   ix6704 : inv02 port map ( Y=>nx6705, A=>nx4109);
   ix6712 : buf02 port map ( Y=>nx6713, A=>nx176);
   ix6720 : inv01 port map ( Y=>nx6721, A=>nx348);
   ix6722 : inv02 port map ( Y=>nx6723, A=>nx6721);
   ix6724 : inv02 port map ( Y=>nx6725, A=>nx6721);
   ix6726 : inv02 port map ( Y=>nx6727, A=>nx6721);
   ix6730 : inv02 port map ( Y=>nx6731, A=>nx6729);
   ix6732 : inv02 port map ( Y=>nx6733, A=>nx7087);
   ix6734 : inv02 port map ( Y=>nx6735, A=>nx7087);
   ix6736 : inv01 port map ( Y=>nx6737, A=>nx1192);
   ix6738 : inv02 port map ( Y=>nx6739, A=>nx6737);
   ix6740 : inv02 port map ( Y=>nx6741, A=>nx6737);
   ix6742 : inv02 port map ( Y=>nx6743, A=>nx6737);
   ix6748 : inv02 port map ( Y=>nx6749, A=>nx4553);
   ix6762 : inv02 port map ( Y=>nx6763, A=>nx6897);
   ix6764 : inv02 port map ( Y=>nx6765, A=>nx6897);
   ix6766 : inv02 port map ( Y=>nx6767, A=>nx6897);
   ix6768 : inv02 port map ( Y=>nx6769, A=>nx7107);
   ix6770 : inv02 port map ( Y=>nx6771, A=>nx7107);
   ix6772 : inv02 port map ( Y=>nx6773, A=>nx7107);
   ix6780 : inv02 port map ( Y=>nx6781, A=>nx7095);
   ix6786 : inv02 port map ( Y=>nx6787, A=>nx5728);
   ix6794 : inv02 port map ( Y=>nx6795, A=>nx6793);
   ix6796 : inv02 port map ( Y=>nx6797, A=>nx6793);
   ix6798 : inv02 port map ( Y=>nx6799, A=>nx6793);
   ix6806 : inv02 port map ( Y=>nx6807, A=>nx6805);
   ix6808 : inv02 port map ( Y=>nx6809, A=>nx6805);
   ix6810 : inv02 port map ( Y=>nx6811, A=>nx6805);
   ix6814 : inv02 port map ( Y=>nx6815, A=>nx6813);
   ix6816 : inv02 port map ( Y=>nx6817, A=>nx6813);
   ix6818 : inv02 port map ( Y=>nx6819, A=>nx6813);
   ix6820 : inv02 port map ( Y=>nx6821, A=>current_state_9);
   ix6822 : inv02 port map ( Y=>nx6823, A=>current_state_9);
   ix6824 : inv02 port map ( Y=>nx6825, A=>nx1516);
   ix6826 : inv02 port map ( Y=>nx6827, A=>nx1516);
   ix6828 : inv02 port map ( Y=>nx6829, A=>nx730);
   ix6830 : inv02 port map ( Y=>nx6831, A=>nx6981);
   ix6832 : inv02 port map ( Y=>nx6833, A=>nx6981);
   ix6834 : buf02 port map ( Y=>nx6835, A=>nx4717);
   ix6836 : buf02 port map ( Y=>nx6837, A=>nx4717);
   ix6838 : buf02 port map ( Y=>nx6839, A=>nx4961);
   ix6850 : inv02 port map ( Y=>nx6851, A=>current_state_18);
   ix6854 : inv02 port map ( Y=>nx6855, A=>nx6985);
   ix6856 : inv02 port map ( Y=>nx6857, A=>nx6985);
   ix6858 : inv02 port map ( Y=>nx6859, A=>nx6985);
   ix6870 : inv02 port map ( Y=>nx6871, A=>nx2536);
   ix6896 : inv02 port map ( Y=>nx6897, A=>nx2098);
   ix6898 : inv02 port map ( Y=>nx6899, A=>current_state_28);
   ix6900 : inv02 port map ( Y=>nx6901, A=>current_state_28);
   ix6902 : inv02 port map ( Y=>nx6903, A=>current_state_28);
   ix6926 : buf02 port map ( Y=>nx6927, A=>comp_unit_operation_EXMPLR);
   ix6928 : buf02 port map ( Y=>nx6929, A=>comp_unit_operation_EXMPLR);
   ix6930 : inv01 port map ( Y=>nx6931, A=>nx7145);
   ix6932 : inv01 port map ( Y=>nx6933, A=>nx7145);
   ix1493 : nor02_2x port map ( Y=>nx1492, A0=>nx4129, A1=>nx7294);
   ix3960 : nor02ii port map ( Y=>nx3959, A0=>nx6927, A1=>layer_type_out_1);
   ix1579 : nor02ii port map ( Y=>nx1578, A0=>nx3975, A1=>io_ready_in);
   ix1801 : and03 port map ( Y=>nx1800, A0=>nx1419, A1=>nx6939, A2=>nx4017);
   ix6938 : inv01 port map ( Y=>nx6939, A=>nx4519);
   ix3990 : and04 port map ( Y=>nx3989, A0=>nx4111, A1=>nx4447, A2=>nx4469, 
      A3=>nx4497);
   ix1621 : mux21_ni port map ( Y=>nx1620, A0=>nx4111, A1=>nx1610, S0=>
      nx1516);
   ix1603 : nor02ii port map ( Y=>nx1602, A0=>nx4009, A1=>nx7021);
   ix167 : nor02ii port map ( Y=>nx4109, A0=>layer_type_out_1, A1=>nx6927);
   ix4010 : and02 port map ( Y=>nx4009, A0=>nx3967, A1=>nx7009);
   ix113 : nor02ii port map ( Y=>nx112, A0=>nx4017, A1=>nx1419);
   ix4018 : and04 port map ( Y=>nx4017, A0=>nflt_layer_out_0, A1=>nx4039, A2
      =>nx4053, A3=>nx6941);
   ix6940 : inv01 port map ( Y=>nx6941, A=>nflt_layer_out_3);
   ix4028 : mux21 port map ( Y=>nx4027, A0=>nx4019, A1=>mem_data_in(0), S0=>
      nx6689);
   ix4034 : nor02ii port map ( Y=>nx4033, A0=>nx6689, A1=>nx4073);
   ix4046 : and02 port map ( Y=>nx4045, A0=>nx4019, A1=>nx4039);
   ix4058 : xor2 port map ( Y=>nx4057, A0=>nx4053, A1=>nx4045);
   ix4068 : and03 port map ( Y=>nx4067, A0=>nx4019, A1=>nx4039, A2=>nx4053);
   ix4081 : or02 port map ( Y=>nx4080, A0=>nx7009, A1=>nx7021);
   ix4114 : nand04 port map ( Y=>nx1516, A0=>nx3967, A1=>nx7009, A2=>nx4073, 
      A3=>nx6823);
   ix4120 : and02 port map ( Y=>nx4119, A0=>nx6823, A1=>nx7009);
   ix4158 : xor2 port map ( Y=>nx4157, A0=>nx4307, A1=>
      new_size_squared_out_15);
   ix4164 : xor2 port map ( Y=>nx4163, A0=>nx4307, A1=>nx1058);
   ix1059 : nor02ii port map ( Y=>nx1058, A0=>nx4175, A1=>
      write_offset_data_out_14);
   ix2190 : ao22 port map ( Y=>nx2189, A0=>nx1064, A1=>nx6981, B0=>
      write_offset_data_out_14, B1=>nx7087);
   ix1013 : nor02ii port map ( Y=>nx1012, A0=>nx4191, A1=>
      write_offset_data_out_12);
   ix2150 : ao22 port map ( Y=>nx2149, A0=>nx1018, A1=>nx6981, B0=>
      write_offset_data_out_12, B1=>nx7087);
   ix965 : nor02ii port map ( Y=>nx964, A0=>nx4207, A1=>
      write_offset_data_out_10);
   ix2110 : ao22 port map ( Y=>nx2109, A0=>nx970, A1=>nx6981, B0=>
      write_offset_data_out_10, B1=>nx7087);
   ix919 : nor02ii port map ( Y=>nx918, A0=>nx4223, A1=>
      write_offset_data_out_8);
   ix2070 : ao22 port map ( Y=>nx2069, A0=>nx924, A1=>nx6983, B0=>
      write_offset_data_out_8, B1=>nx7087);
   ix733 : nor02ii port map ( Y=>nx6729, A0=>nx6983, A1=>nx4123);
   ix4234 : nand02 port map ( Y=>nx730, A0=>nx4129, A1=>nx4149);
   ix869 : nor02ii port map ( Y=>nx868, A0=>nx4246, A1=>
      write_offset_data_out_6);
   ix2030 : ao22 port map ( Y=>nx2029, A0=>nx874, A1=>nx6983, B0=>
      write_offset_data_out_6, B1=>nx7087);
   ix823 : nor02ii port map ( Y=>nx822, A0=>nx4265, A1=>
      write_offset_data_out_4);
   ix1990 : ao22 port map ( Y=>nx1989, A0=>write_offset_data_out_4, A1=>
      nx7089, B0=>nx828, B1=>nx6983);
   ix4266 : or04 port map ( Y=>nx4265, A0=>nx4271, A1=>nx4277, A2=>nx7355, 
      A3=>nx4293);
   ix1970 : ao22 port map ( Y=>nx1969, A0=>write_offset_data_out_3, A1=>
      nx7089, B0=>nx802, B1=>nx6983);
   ix1910 : mux21_ni port map ( Y=>nx1909, A0=>nx7089, A1=>nx6983, S0=>
      nx4293);
   ix4296 : or02 port map ( Y=>nx4295, A0=>nx7355, A1=>nx4293);
   ix4300 : or03 port map ( Y=>nx4299, A0=>nx4277, A1=>nx7355, A2=>nx4293);
   ix2220 : mux21_ni port map ( Y=>nx2219, A0=>mem_data_in(15), A1=>
      new_size_squared_out_15, S0=>nx7081);
   ix4316 : xnor2 port map ( Y=>nx4314, A0=>nx4167, A1=>nx4320);
   ix2200 : mux21_ni port map ( Y=>nx2199, A0=>mem_data_in(14), A1=>
      new_size_squared_out_14, S0=>nx7081);
   ix4322 : xor2 port map ( Y=>nx4321, A0=>nx4305, A1=>
      new_size_squared_out_13);
   ix2180 : mux21_ni port map ( Y=>nx2179, A0=>mem_data_in(13), A1=>
      new_size_squared_out_13, S0=>nx7081);
   ix4330 : xnor2 port map ( Y=>nx4328, A0=>nx4183, A1=>nx4335);
   ix2160 : mux21_ni port map ( Y=>nx2159, A0=>mem_data_in(12), A1=>
      new_size_squared_out_12, S0=>nx7081);
   ix4338 : xor2 port map ( Y=>nx4337, A0=>nx4303, A1=>
      new_size_squared_out_11);
   ix2140 : mux21_ni port map ( Y=>nx2139, A0=>mem_data_in(11), A1=>
      new_size_squared_out_11, S0=>nx7081);
   ix4344 : xnor2 port map ( Y=>nx4343, A0=>nx4200, A1=>nx4349);
   ix2120 : mux21_ni port map ( Y=>nx2119, A0=>mem_data_in(10), A1=>
      new_size_squared_out_10, S0=>nx7081);
   ix4352 : xor2 port map ( Y=>nx4351, A0=>nx4301, A1=>
      new_size_squared_out_9);
   ix2100 : mux21_ni port map ( Y=>nx2099, A0=>mem_data_in(9), A1=>
      new_size_squared_out_9, S0=>nx7083);
   ix4359 : xnor2 port map ( Y=>nx4358, A0=>nx4217, A1=>nx4363);
   ix2080 : mux21_ni port map ( Y=>nx2079, A0=>mem_data_in(8), A1=>
      new_size_squared_out_8, S0=>nx7083);
   ix4366 : xor2 port map ( Y=>nx4365, A0=>nx4229, A1=>
      new_size_squared_out_7);
   ix2060 : mux21_ni port map ( Y=>nx2059, A0=>mem_data_in(7), A1=>
      new_size_squared_out_7, S0=>nx7083);
   ix4373 : xnor2 port map ( Y=>nx4372, A0=>nx4239, A1=>nx4377);
   ix2040 : mux21_ni port map ( Y=>nx2039, A0=>mem_data_in(6), A1=>
      new_size_squared_out_6, S0=>nx7083);
   ix4380 : xor2 port map ( Y=>nx4379, A0=>nx4251, A1=>
      new_size_squared_out_5);
   ix2020 : mux21_ni port map ( Y=>nx2019, A0=>mem_data_in(5), A1=>
      new_size_squared_out_5, S0=>nx7083);
   ix4387 : xnor2 port map ( Y=>nx4386, A0=>nx4257, A1=>nx4391);
   ix2000 : mux21_ni port map ( Y=>nx1999, A0=>mem_data_in(4), A1=>
      new_size_squared_out_4, S0=>nx7083);
   ix4394 : xor2 port map ( Y=>nx4393, A0=>nx4271, A1=>
      new_size_squared_out_3);
   ix1980 : mux21_ni port map ( Y=>nx1979, A0=>mem_data_in(3), A1=>
      new_size_squared_out_3, S0=>nx7083);
   ix4402 : xnor2 port map ( Y=>nx4400, A0=>nx4277, A1=>nx4407);
   ix1960 : mux21_ni port map ( Y=>nx1959, A0=>mem_data_in(2), A1=>
      new_size_squared_out_2, S0=>nx7085);
   ix4410 : xor2 port map ( Y=>nx4408, A0=>nx7355, A1=>
      new_size_squared_out_1);
   ix1940 : mux21_ni port map ( Y=>nx1939, A0=>mem_data_in(1), A1=>
      new_size_squared_out_1, S0=>nx7085);
   ix4418 : xnor2 port map ( Y=>nx4417, A0=>nx4293, A1=>nx4423);
   ix1920 : mux21_ni port map ( Y=>nx1919, A0=>mem_data_in(0), A1=>
      new_size_squared_out_0, S0=>nx7085);
   ix1631 : xnor2 port map ( Y=>nx1630, A0=>nx4447, A1=>nx4111);
   ix4472 : and02 port map ( Y=>nx4471, A0=>nx4111, A1=>nx4447);
   ix4500 : and03 port map ( Y=>nx4499, A0=>nx4111, A1=>nx4447, A2=>nx4469);
   ix1769 : mux21 port map ( Y=>nx1768, A0=>nx4047, A1=>nx4526, S0=>nx3967);
   ix4534 : mux21 port map ( Y=>nx4533, A0=>mem_data_in(0), A1=>nx4531, S0=>
      nx3967);
   ix4536 : nor02ii port map ( Y=>nx4535, A0=>nlayers_counter_out_1, A1=>
      nx4531);
   ix1785 : mux21 port map ( Y=>nx1784, A0=>nx4059, A1=>nx4543, S0=>nx3967);
   ix1447 : ao32 port map ( Y=>nx1446, A0=>nx4583, A1=>current_state_15, A2
      =>nx4759, B0=>current_state_16, B1=>ftc_cntrl_reg_out_11);
   ix4564 : or02 port map ( Y=>nx4563, A0=>ftc_cntrl_reg_out_14, A1=>nx7294
   );
   ix4572 : nor02ii port map ( Y=>nx4571, A0=>nx4, A1=>nx4879);
   ix5 : and02 port map ( Y=>nx4, A0=>current_state_20, A1=>nx4705);
   ix281 : xnor2 port map ( Y=>nx280, A0=>nx4647, A1=>nx278);
   ix1570 : mux21_ni port map ( Y=>nx1569, A0=>nx232, A1=>
      cntr1_inst_counter_out_4, S0=>nx7029);
   ix233 : xor2 port map ( Y=>nx232, A0=>nx4647, A1=>nx4601);
   ix1560 : mux21_ni port map ( Y=>nx1559, A0=>nx214, A1=>
      cntr1_inst_counter_out_3, S0=>nx7029);
   ix1550 : mux21_ni port map ( Y=>nx1549, A0=>nx200, A1=>
      cntr1_inst_counter_out_2, S0=>nx7029);
   ix1540 : mux21 port map ( Y=>nx1539, A0=>nx4638, A1=>nx4621, S0=>nx7029);
   ix177 : oai21 port map ( Y=>nx176, A0=>nx4637, A1=>nx7021, B0=>nx6599);
   ix279 : or02 port map ( Y=>nx278, A0=>nx7063, A1=>nx7031);
   ix249 : xor2 port map ( Y=>nx248, A0=>nx7295, A1=>
      cntr1_inst_counter_out_2);
   ix247 : xnor2 port map ( Y=>nx246, A0=>nx7295, A1=>nx4655);
   ix1580 : mux21 port map ( Y=>nx1579, A0=>nx4657, A1=>nx4655, S0=>nx7295);
   ix4658 : xor2 port map ( Y=>nx4657, A0=>nx4655, A1=>nx1425);
   ix239 : nor02ii port map ( Y=>nx1425, A0=>nx4601, A1=>
      cntr1_inst_counter_out_4);
   ix4664 : xnor2 port map ( Y=>nx4663, A0=>nx7295, A1=>
      cntr1_inst_counter_out_1);
   ix4674 : nor02ii port map ( Y=>nx4673, A0=>nx1469, A1=>nx4725);
   ix1851 : and02 port map ( Y=>nx1469, A0=>current_state_20, A1=>nx4705);
   ix1371 : and04 port map ( Y=>nx1370, A0=>nx5148, A1=>nx4692, A2=>nx5146, 
      A3=>nx5023);
   ix2400 : mux21 port map ( Y=>nx2399, A0=>nx5148, A1=>nx4689, S0=>nx7101);
   ix4690 : xor2 port map ( Y=>nx4689, A0=>nx5148, A1=>nx1447);
   ix1351 : nor02ii port map ( Y=>nx1447, A0=>nx5013, A1=>
      cache_width_cntr_counter_out_14);
   ix2390 : mux21_ni port map ( Y=>nx2389, A0=>
      cache_width_cntr_counter_out_14, A1=>nx1344, S0=>nx7101);
   ix1345 : xor2 port map ( Y=>nx1344, A0=>nx4692, A1=>nx5013);
   ix319 : nor02ii port map ( Y=>nx1427, A0=>nx7033, A1=>nx4723);
   ix4718 : and04 port map ( Y=>nx4717, A0=>nx5113, A1=>nx4725, A2=>nx4765, 
      A3=>nx4879);
   ix547 : or02 port map ( Y=>nx546, A0=>ftc_cntrl_reg_out_11, A1=>nx4765);
   ix521 : and04 port map ( Y=>nx520, A0=>nx4743, A1=>nx4770, A2=>nx4781, A3
      =>nx4787);
   ix1780 : mux21 port map ( Y=>nx1779, A0=>nx4767, A1=>nx4743, S0=>nx7037);
   ix4752 : or03 port map ( Y=>nx4751, A0=>ftc_cntrl_reg_out_8, A1=>nx4725, 
      A2=>nx4759);
   ix1117 : ao21 port map ( Y=>nx1116, A0=>nx7033, A1=>nx4575, B0=>
      current_state_16);
   ix4768 : xor2 port map ( Y=>nx4767, A0=>nx4743, A1=>nx1430);
   ix501 : nor02ii port map ( Y=>nx1430, A0=>nx4776, A1=>
      window_width_cntr_counter_out_14);
   ix1770 : mux21_ni port map ( Y=>nx1769, A0=>nx494, A1=>
      window_width_cntr_counter_out_14, S0=>nx7037);
   ix495 : xor2 port map ( Y=>nx494, A0=>nx4770, A1=>nx4776);
   ix1760 : mux21 port map ( Y=>nx1759, A0=>nx4783, A1=>nx4781, S0=>nx7037);
   ix477 : nor02ii port map ( Y=>nx1432, A0=>nx4795, A1=>
      window_width_cntr_counter_out_12);
   ix1750 : mux21_ni port map ( Y=>nx1749, A0=>nx470, A1=>
      window_width_cntr_counter_out_12, S0=>nx7037);
   ix471 : xor2 port map ( Y=>nx470, A0=>nx4787, A1=>nx4795);
   ix1740 : mux21 port map ( Y=>nx1739, A0=>nx4803, A1=>nx4801, S0=>nx7037);
   ix453 : nor02ii port map ( Y=>nx1434, A0=>nx4813, A1=>
      window_width_cntr_counter_out_10);
   ix1730 : mux21_ni port map ( Y=>nx1729, A0=>nx446, A1=>
      window_width_cntr_counter_out_10, S0=>nx7037);
   ix447 : xor2 port map ( Y=>nx446, A0=>nx4807, A1=>nx4813);
   ix1720 : mux21 port map ( Y=>nx1719, A0=>nx4821, A1=>nx4819, S0=>nx7037);
   ix429 : nor02ii port map ( Y=>nx1436, A0=>nx4833, A1=>
      window_width_cntr_counter_out_8);
   ix1710 : mux21_ni port map ( Y=>nx1709, A0=>nx422, A1=>
      window_width_cntr_counter_out_8, S0=>nx7039);
   ix423 : xor2 port map ( Y=>nx422, A0=>nx4825, A1=>nx4833);
   ix1700 : mux21 port map ( Y=>nx1699, A0=>nx4841, A1=>nx4839, S0=>nx7039);
   ix405 : nor02ii port map ( Y=>nx1439, A0=>nx4853, A1=>
      window_width_cntr_counter_out_6);
   ix1690 : mux21_ni port map ( Y=>nx1689, A0=>nx398, A1=>
      window_width_cntr_counter_out_6, S0=>nx7039);
   ix399 : xor2 port map ( Y=>nx398, A0=>nx4845, A1=>nx4853);
   ix4854 : or03 port map ( Y=>nx4853, A0=>nx6943, A1=>nx4911, A2=>nx4861);
   ix6942 : inv01 port map ( Y=>nx6943, A=>wind_width_count_4);
   ix2600 : mux21_ni port map ( Y=>nx2599, A0=>nx1880, A1=>
      wind_width_count_4, S0=>nx7039);
   ix1650 : mux21_ni port map ( Y=>nx1649, A0=>nx354, A1=>wind_width_count_1, 
      S0=>nx7039);
   ix1640 : xor2 port map ( Y=>nx1639, A0=>nx6607, A1=>nx1429);
   ix1660 : mux21_ni port map ( Y=>nx1659, A0=>nx362, A1=>wind_width_count_2, 
      S0=>nx7039);
   ix1670 : mux21_ni port map ( Y=>nx1669, A0=>nx370, A1=>wind_width_count_3, 
      S0=>nx7039);
   ix1680 : mux21 port map ( Y=>nx1679, A0=>nx4913, A1=>nx4911, S0=>nx7041);
   ix535 : and04 port map ( Y=>nx534, A0=>nx4801, A1=>nx4807, A2=>nx4819, A3
      =>nx4825);
   ix583 : and04 port map ( Y=>nx582, A0=>nx4839, A1=>nx4845, A2=>nx4911, A3
      =>nx6945);
   ix6944 : inv01 port map ( Y=>nx6945, A=>nx574);
   ix573 : mux21 port map ( Y=>nx572, A0=>nx7063, A1=>img_width_out_0, S0=>
      nx6977);
   ix1800 : ao221 port map ( Y=>nx1799, A0=>img_width_out_0, A1=>nx4119, B0
      =>nx6665, B1=>new_width_out_0, C0=>current_state_9);
   ix611 : mux21 port map ( Y=>nx610, A0=>nx7065, A1=>nx5155, S0=>nx6977);
   ix675 : nor02ii port map ( Y=>nx674, A0=>nx4981, A1=>nx6977);
   ix693 : nor02ii port map ( Y=>nx692, A0=>nx4997, A1=>nx6979);
   ix5012 : or02 port map ( Y=>nx5011, A0=>nx4575, A1=>nx4705);
   ix2380 : mux21 port map ( Y=>nx2379, A0=>nx5146, A1=>nx5019, S0=>nx7101);
   ix1327 : nor02ii port map ( Y=>nx1449, A0=>nx5031, A1=>
      cache_width_cntr_counter_out_12);
   ix2370 : mux21_ni port map ( Y=>nx2369, A0=>
      cache_width_cntr_counter_out_12, A1=>nx1320, S0=>nx7101);
   ix1321 : xor2 port map ( Y=>nx1320, A0=>nx5023, A1=>nx5031);
   ix2360 : mux21 port map ( Y=>nx2359, A0=>nx5144, A1=>nx5037, S0=>nx7101);
   ix1303 : nor02ii port map ( Y=>nx1451, A0=>nx5049, A1=>
      cache_width_cntr_counter_out_10);
   ix2350 : mux21_ni port map ( Y=>nx2349, A0=>
      cache_width_cntr_counter_out_10, A1=>nx1296, S0=>nx7101);
   ix1297 : xor2 port map ( Y=>nx1296, A0=>nx5041, A1=>nx5049);
   ix2340 : mux21 port map ( Y=>nx2339, A0=>nx5142, A1=>nx5055, S0=>nx7101);
   ix1279 : nor02ii port map ( Y=>nx1454, A0=>nx5067, A1=>
      cache_width_cntr_counter_out_8);
   ix2330 : mux21_ni port map ( Y=>nx2329, A0=>
      cache_width_cntr_counter_out_8, A1=>nx1272, S0=>nx7103);
   ix1273 : xor2 port map ( Y=>nx1272, A0=>nx5059, A1=>nx5067);
   ix2320 : mux21 port map ( Y=>nx2319, A0=>nx5140, A1=>nx5072, S0=>nx7103);
   ix1255 : nor02ii port map ( Y=>nx1456, A0=>nx5083, A1=>
      cache_width_cntr_counter_out_6);
   ix2310 : mux21_ni port map ( Y=>nx2309, A0=>
      cache_width_cntr_counter_out_6, A1=>nx1248, S0=>nx7103);
   ix1249 : xor2 port map ( Y=>nx1248, A0=>nx5077, A1=>nx5083);
   ix5084 : or03 port map ( Y=>nx5083, A0=>nx6947, A1=>nx5137, A2=>nx5089);
   ix6946 : inv01 port map ( Y=>nx6947, A=>nx6613);
   ix2290 : mux21_ni port map ( Y=>nx2289, A0=>nx6611, A1=>nx1222, S0=>
      nx7103);
   ix2260 : mux21_ni port map ( Y=>nx2259, A0=>cache_width_count_1, A1=>
      nx1198, S0=>nx7103);
   ix2250 : xor2 port map ( Y=>nx2249, A0=>cache_width_count_0, A1=>nx7103);
   ix5114 : and02 port map ( Y=>nx5113, A0=>nx7033, A1=>nx4575);
   ix2270 : mux21_ni port map ( Y=>nx2269, A0=>nx6615, A1=>nx1206, S0=>
      nx7103);
   ix2280 : mux21_ni port map ( Y=>nx2279, A0=>cache_width_count_3, A1=>
      nx1214, S0=>nx7105);
   ix2300 : mux21 port map ( Y=>nx2299, A0=>nx5137, A1=>nx5134, S0=>nx7105);
   ix1385 : and04 port map ( Y=>nx1384, A0=>nx5144, A1=>nx5041, A2=>nx5142, 
      A3=>nx5059);
   ix1403 : and04 port map ( Y=>nx1402, A0=>nx5140, A1=>nx5077, A2=>nx5137, 
      A3=>nx6949);
   ix1395 : xnor2 port map ( Y=>nx6949, A0=>nx4927, A1=>cache_width_count_0
   );
   ix1405 : xor2 port map ( Y=>nx1404, A0=>cache_width_count_1, A1=>nx606);
   ix5158 : nor02ii port map ( Y=>nx5157, A0=>img_width_out_1, A1=>nx4927);
   ix1453 : nor02_2x port map ( Y=>nx1452, A0=>nx7023, A1=>nx7065);
   ix1871 : and02 port map ( Y=>nx1459, A0=>current_state_21, A1=>nx4731);
   ix2610 : mux21 port map ( Y=>nx2609, A0=>current_state_27, A1=>nx7043, S0
      =>nx5194);
   ix2620 : mux21 port map ( Y=>nx2619, A0=>nx5204, A1=>nx5202, S0=>nx7043);
   ix5207 : or02 port map ( Y=>nx5206, A0=>nx5202, A1=>nx5194);
   ix2630 : mux21_ni port map ( Y=>nx2629, A0=>nx1908, A1=>
      class_cntr_counter_out_2, S0=>nx7043);
   ix1909 : xor2 port map ( Y=>nx1908, A0=>nx5208, A1=>nx5206);
   ix2640 : mux21_ni port map ( Y=>nx2639, A0=>nx1916, A1=>
      class_cntr_counter_out_3, S0=>nx5191);
   ix1917 : xor2 port map ( Y=>nx1916, A0=>nx5218, A1=>nx5216);
   ix5217 : or03 port map ( Y=>nx5216, A0=>nx5208, A1=>nx5202, A2=>nx5194);
   ix4847 : nor02ii port map ( Y=>argmax_data_out(0), A0=>argmax_ready_dup0, 
      A1=>mem_data_in(0));
   ix4849 : nor02ii port map ( Y=>argmax_data_out(1), A0=>nx7325, A1=>
      mem_data_in(1));
   ix4851 : nor02ii port map ( Y=>argmax_data_out(2), A0=>nx7326, A1=>
      mem_data_in(2));
   ix4855 : nor02ii port map ( Y=>argmax_data_out(4), A0=>nx7327, A1=>
      mem_data_in(4));
   ix4857 : nor02ii port map ( Y=>argmax_data_out(5), A0=>nx7328, A1=>
      mem_data_in(5));
   ix4861 : nor02ii port map ( Y=>argmax_data_out(7), A0=>nx7047, A1=>
      mem_data_in(7));
   ix4863 : nor02ii port map ( Y=>argmax_data_out(8), A0=>nx7047, A1=>
      mem_data_in(8));
   ix4865 : nor02ii port map ( Y=>argmax_data_out(9), A0=>nx7047, A1=>
      mem_data_in(9));
   ix4867 : nor02ii port map ( Y=>argmax_data_out(10), A0=>nx7047, A1=>
      mem_data_in(10));
   ix4869 : nor02ii port map ( Y=>argmax_data_out(11), A0=>nx7047, A1=>
      mem_data_in(11));
   ix4871 : nor02ii port map ( Y=>argmax_data_out(12), A0=>nx7047, A1=>
      mem_data_in(12));
   ix4873 : nor02ii port map ( Y=>argmax_data_out(13), A0=>nx7049, A1=>
      mem_data_in(13));
   ix4875 : nor02ii port map ( Y=>argmax_data_out(14), A0=>nx7049, A1=>
      mem_data_in(14));
   ix4877 : nor02ii port map ( Y=>argmax_data_out(15), A0=>nx7049, A1=>
      mem_data_in(15));
   ix4879 : and02 port map ( Y=>comp_unit_data2_out(0), A0=>nx6985, A1=>
      nx2096);
   ix2097 : mux21_ni port map ( Y=>nx2096, A0=>flt_bias_out_0, A1=>
      mem_data_in(0), S0=>nx7053);
   ix2085 : nor02ii port map ( Y=>nx2084, A0=>nx6927, A1=>current_state_12);
   ix4881 : and02 port map ( Y=>comp_unit_data2_out(1), A0=>nx6987, A1=>
      nx2124);
   ix2125 : mux21_ni port map ( Y=>nx2124, A0=>flt_bias_out_1, A1=>
      mem_data_in(1), S0=>nx7053);
   ix4883 : and02 port map ( Y=>comp_unit_data2_out(2), A0=>nx6987, A1=>
      nx2150);
   ix2151 : mux21_ni port map ( Y=>nx2150, A0=>flt_bias_out_2, A1=>
      mem_data_in(2), S0=>nx7053);
   ix4885 : and02 port map ( Y=>comp_unit_data2_out(3), A0=>nx6987, A1=>
      nx2176);
   ix2177 : mux21_ni port map ( Y=>nx2176, A0=>flt_bias_out_3, A1=>
      mem_data_in(3), S0=>nx7053);
   ix4887 : and02 port map ( Y=>comp_unit_data2_out(4), A0=>nx6987, A1=>
      nx2202);
   ix2203 : mux21_ni port map ( Y=>nx2202, A0=>flt_bias_out_4, A1=>
      mem_data_in(4), S0=>nx7053);
   ix4889 : and02 port map ( Y=>comp_unit_data2_out(5), A0=>nx6987, A1=>
      nx2228);
   ix2229 : mux21_ni port map ( Y=>nx2228, A0=>flt_bias_out_5, A1=>
      mem_data_in(5), S0=>nx7055);
   ix4891 : and02 port map ( Y=>comp_unit_data2_out(6), A0=>nx6987, A1=>
      nx2254);
   ix2255 : mux21_ni port map ( Y=>nx2254, A0=>flt_bias_out_6, A1=>
      mem_data_in(6), S0=>nx7055);
   ix4893 : and02 port map ( Y=>comp_unit_data2_out(7), A0=>nx6987, A1=>
      nx2280);
   ix2281 : mux21_ni port map ( Y=>nx2280, A0=>flt_bias_out_7, A1=>
      mem_data_in(7), S0=>nx7055);
   ix4895 : and02 port map ( Y=>comp_unit_data2_out(8), A0=>nx6989, A1=>
      nx2306);
   ix2307 : mux21_ni port map ( Y=>nx2306, A0=>flt_bias_out_8, A1=>
      mem_data_in(8), S0=>nx7055);
   ix4897 : and02 port map ( Y=>comp_unit_data2_out(9), A0=>nx6989, A1=>
      nx2332);
   ix2333 : mux21_ni port map ( Y=>nx2332, A0=>flt_bias_out_9, A1=>
      mem_data_in(9), S0=>nx7055);
   ix4899 : and02 port map ( Y=>comp_unit_data2_out(10), A0=>nx6989, A1=>
      nx2358);
   ix2359 : mux21_ni port map ( Y=>nx2358, A0=>flt_bias_out_10, A1=>
      mem_data_in(10), S0=>nx7055);
   ix4901 : and02 port map ( Y=>comp_unit_data2_out(11), A0=>nx6989, A1=>
      nx2384);
   ix2385 : mux21_ni port map ( Y=>nx2384, A0=>flt_bias_out_11, A1=>
      mem_data_in(11), S0=>nx7055);
   ix4903 : and02 port map ( Y=>comp_unit_data2_out(12), A0=>nx6989, A1=>
      nx2410);
   ix2411 : mux21_ni port map ( Y=>nx2410, A0=>flt_bias_out_12, A1=>
      mem_data_in(12), S0=>nx7057);
   ix4905 : and02 port map ( Y=>comp_unit_data2_out(13), A0=>nx6989, A1=>
      nx2436);
   ix2437 : mux21_ni port map ( Y=>nx2436, A0=>flt_bias_out_13, A1=>
      mem_data_in(13), S0=>nx7057);
   ix4907 : and02 port map ( Y=>comp_unit_data2_out(14), A0=>nx6989, A1=>
      nx2462);
   ix2463 : mux21_ni port map ( Y=>nx2462, A0=>flt_bias_out_14, A1=>
      mem_data_in(14), S0=>nx7057);
   ix4909 : and02 port map ( Y=>comp_unit_data2_out(15), A0=>nx6991, A1=>
      nx2488);
   ix2489 : mux21_ni port map ( Y=>nx2488, A0=>flt_bias_out_15, A1=>
      mem_data_in(15), S0=>nx7057);
   ix5077 : and03 port map ( Y=>max_height_1, A0=>nx606, A1=>nx6599, A2=>
      nx7035);
   ix5111 : nor04 port map ( Y=>comp_unit_relu, A0=>nx6951, A1=>nx4111, A2=>
      num_channels_out_2, A3=>num_channels_out_1);
   ix5101 : nand04 port map ( Y=>nx6951, A0=>nx4004, A1=>nx6953, A2=>nx4503, 
      A3=>nx4497);
   ix6952 : inv01 port map ( Y=>nx6953, A=>nx6927);
   ix2573 : oai21 port map ( Y=>cache_load, A0=>nx7065, A1=>nx6955, B0=>
      nx7107);
   ix6954 : inv01 port map ( Y=>nx6955, A=>nx4);
   ix2523 : or03 port map ( Y=>nx2522, A0=>nx4723, A1=>current_state_20, A2
      =>nx7035);
   ix2539 : and02 port map ( Y=>cache_data_in_0, A0=>mem_data_in(0), A1=>
      nx6999);
   ix5340 : ao21 port map ( Y=>nx2536, A0=>nx5334, A1=>nx1469, B0=>nx1152);
   ix2541 : and02 port map ( Y=>cache_data_in_1, A0=>mem_data_in(1), A1=>
      nx6999);
   ix2543 : and02 port map ( Y=>cache_data_in_2, A0=>mem_data_in(2), A1=>
      nx6999);
   ix2545 : and02 port map ( Y=>cache_data_in_3, A0=>mem_data_in(3), A1=>
      nx6999);
   ix2547 : and02 port map ( Y=>cache_data_in_4, A0=>mem_data_in(4), A1=>
      nx6999);
   ix2549 : and02 port map ( Y=>cache_data_in_5, A0=>mem_data_in(5), A1=>
      nx6999);
   ix2551 : and02 port map ( Y=>cache_data_in_6, A0=>mem_data_in(6), A1=>
      nx6999);
   ix2553 : and02 port map ( Y=>cache_data_in_7, A0=>mem_data_in(7), A1=>
      nx7001);
   ix2555 : and02 port map ( Y=>cache_data_in_8, A0=>mem_data_in(8), A1=>
      nx7001);
   ix2557 : and02 port map ( Y=>cache_data_in_9, A0=>mem_data_in(9), A1=>
      nx7001);
   ix2559 : and02 port map ( Y=>cache_data_in_10, A0=>mem_data_in(10), A1=>
      nx7001);
   ix2561 : and02 port map ( Y=>cache_data_in_11, A0=>mem_data_in(11), A1=>
      nx7001);
   ix2563 : and02 port map ( Y=>cache_data_in_12, A0=>mem_data_in(12), A1=>
      nx7001);
   ix2565 : and02 port map ( Y=>cache_data_in_13, A0=>mem_data_in(13), A1=>
      nx7001);
   ix2567 : and02 port map ( Y=>cache_data_in_14, A0=>mem_data_in(14), A1=>
      nx7003);
   ix2569 : and02 port map ( Y=>cache_data_in_15, A0=>mem_data_in(15), A1=>
      nx7003);
   ix5380 : and02 port map ( Y=>nx5379, A0=>nx6599, A1=>nx7035);
   ix2670 : mux21 port map ( Y=>nx2669, A0=>nx5386, A1=>nx5383, S0=>nx7023);
   ix2690 : mux21 port map ( Y=>nx2689, A0=>nx5393, A1=>nx5390, S0=>nx7023);
   ix2710 : mux21 port map ( Y=>nx2709, A0=>nx5399, A1=>nx5396, S0=>nx7023);
   ix2730 : mux21 port map ( Y=>nx2729, A0=>nx5405, A1=>nx5402, S0=>nx7023);
   ix2750 : mux21 port map ( Y=>nx2749, A0=>nx5411, A1=>nx5408, S0=>nx7025);
   ix2770 : mux21 port map ( Y=>nx2769, A0=>nx5417, A1=>nx5414, S0=>nx7025);
   ix2790 : mux21 port map ( Y=>nx2789, A0=>nx5423, A1=>nx5420, S0=>nx7025);
   ix2810 : mux21 port map ( Y=>nx2809, A0=>nx5429, A1=>nx5426, S0=>nx7025);
   ix2830 : mux21 port map ( Y=>nx2829, A0=>nx5435, A1=>nx5432, S0=>nx7025);
   ix2850 : mux21 port map ( Y=>nx2849, A0=>nx5441, A1=>nx5438, S0=>nx7025);
   ix2870 : mux21 port map ( Y=>nx2869, A0=>nx5447, A1=>nx5444, S0=>nx7025);
   ix2890 : mux21 port map ( Y=>nx2889, A0=>nx5453, A1=>nx5450, S0=>nx7027);
   ix2910 : mux21 port map ( Y=>nx2909, A0=>nx5459, A1=>nx5456, S0=>nx7027);
   ix2930 : mux21 port map ( Y=>nx2929, A0=>nx5465, A1=>nx5462, S0=>nx7027);
   ix2950 : mux21 port map ( Y=>nx2949, A0=>nx5471, A1=>nx5468, S0=>nx7027);
   ix2970 : mux21 port map ( Y=>nx2969, A0=>nx5477, A1=>nx5474, S0=>nx7027);
   ix4815 : nor02ii port map ( Y=>filter_data_out(0), A0=>nx7077, A1=>
      mem_data_in(0));
   ix4817 : nor02ii port map ( Y=>filter_data_out(1), A0=>nx7077, A1=>
      mem_data_in(1));
   ix4819 : nor02ii port map ( Y=>filter_data_out(2), A0=>nx7077, A1=>
      mem_data_in(2));
   ix4821 : nor02ii port map ( Y=>filter_data_out(3), A0=>nx7077, A1=>
      mem_data_in(3));
   ix4823 : nor02ii port map ( Y=>filter_data_out(4), A0=>nx7077, A1=>
      mem_data_in(4));
   ix4825 : nor02ii port map ( Y=>filter_data_out(5), A0=>nx7079, A1=>
      mem_data_in(5));
   ix4827 : nor02ii port map ( Y=>filter_data_out(6), A0=>nx7079, A1=>
      mem_data_in(6));
   ix4829 : nor02ii port map ( Y=>filter_data_out(7), A0=>nx7079, A1=>
      mem_data_in(7));
   ix4831 : nor02ii port map ( Y=>filter_data_out(8), A0=>nx7079, A1=>
      mem_data_in(8));
   ix4833 : nor02ii port map ( Y=>filter_data_out(9), A0=>nx7079, A1=>
      mem_data_in(9));
   ix4835 : nor02ii port map ( Y=>filter_data_out(10), A0=>nx7079, A1=>
      mem_data_in(10));
   ix4837 : nor02ii port map ( Y=>filter_data_out(11), A0=>nx7079, A1=>
      mem_data_in(11));
   ix4839 : nor02ii port map ( Y=>filter_data_out(12), A0=>nx6657, A1=>
      mem_data_in(12));
   ix4841 : nor02ii port map ( Y=>filter_data_out(13), A0=>nx6657, A1=>
      mem_data_in(13));
   ix4843 : nor02ii port map ( Y=>filter_data_out(14), A0=>nx6657, A1=>
      mem_data_in(14));
   ix4845 : nor02ii port map ( Y=>filter_data_out(15), A0=>nx6657, A1=>
      mem_data_in(15));
   ix4911 : and02 port map ( Y=>wind_col_in_0_0, A0=>nx7123, A1=>
      cache_data_out_0_0);
   ix4913 : and02 port map ( Y=>wind_col_in_0_1, A0=>nx7123, A1=>
      cache_data_out_0_1);
   ix4915 : and02 port map ( Y=>wind_col_in_0_2, A0=>nx7123, A1=>
      cache_data_out_0_2);
   ix4917 : and02 port map ( Y=>wind_col_in_0_3, A0=>nx7123, A1=>
      cache_data_out_0_3);
   ix4919 : and02 port map ( Y=>wind_col_in_0_4, A0=>nx7123, A1=>
      cache_data_out_0_4);
   ix4921 : and02 port map ( Y=>wind_col_in_0_5, A0=>nx7123, A1=>
      cache_data_out_0_5);
   ix4923 : and02 port map ( Y=>wind_col_in_0_6, A0=>nx7123, A1=>
      cache_data_out_0_6);
   ix4925 : and02 port map ( Y=>wind_col_in_0_7, A0=>nx7125, A1=>
      cache_data_out_0_7);
   ix4927 : and02 port map ( Y=>wind_col_in_0_8, A0=>nx7125, A1=>
      cache_data_out_0_8);
   ix4929 : and02 port map ( Y=>wind_col_in_0_9, A0=>nx7125, A1=>
      cache_data_out_0_9);
   ix4931 : and02 port map ( Y=>wind_col_in_0_10, A0=>nx7125, A1=>
      cache_data_out_0_10);
   ix4933 : and02 port map ( Y=>wind_col_in_0_11, A0=>nx7125, A1=>
      cache_data_out_0_11);
   ix4935 : and02 port map ( Y=>wind_col_in_0_12, A0=>nx7125, A1=>
      cache_data_out_0_12);
   ix4937 : and02 port map ( Y=>wind_col_in_0_13, A0=>nx7125, A1=>
      cache_data_out_0_13);
   ix4939 : and02 port map ( Y=>wind_col_in_0_14, A0=>nx7127, A1=>
      cache_data_out_0_14);
   ix4941 : and02 port map ( Y=>wind_col_in_0_15, A0=>nx7127, A1=>
      cache_data_out_0_15);
   ix4943 : and02 port map ( Y=>wind_col_in_1_0, A0=>nx7127, A1=>
      cache_data_out_1_0);
   ix4945 : and02 port map ( Y=>wind_col_in_1_1, A0=>nx7127, A1=>
      cache_data_out_1_1);
   ix4947 : and02 port map ( Y=>wind_col_in_1_2, A0=>nx7127, A1=>
      cache_data_out_1_2);
   ix4949 : and02 port map ( Y=>wind_col_in_1_3, A0=>nx7127, A1=>
      cache_data_out_1_3);
   ix4951 : and02 port map ( Y=>wind_col_in_1_4, A0=>nx7127, A1=>
      cache_data_out_1_4);
   ix4953 : and02 port map ( Y=>wind_col_in_1_5, A0=>nx7129, A1=>
      cache_data_out_1_5);
   ix4955 : and02 port map ( Y=>wind_col_in_1_6, A0=>nx7129, A1=>
      cache_data_out_1_6);
   ix4957 : and02 port map ( Y=>wind_col_in_1_7, A0=>nx7129, A1=>
      cache_data_out_1_7);
   ix4959 : and02 port map ( Y=>wind_col_in_1_8, A0=>nx7129, A1=>
      cache_data_out_1_8);
   ix4961 : and02 port map ( Y=>wind_col_in_1_9, A0=>nx7129, A1=>
      cache_data_out_1_9);
   ix4963 : and02 port map ( Y=>wind_col_in_1_10, A0=>nx7129, A1=>
      cache_data_out_1_10);
   ix4965 : and02 port map ( Y=>wind_col_in_1_11, A0=>nx7129, A1=>
      cache_data_out_1_11);
   ix4967 : and02 port map ( Y=>wind_col_in_1_12, A0=>nx7131, A1=>
      cache_data_out_1_12);
   ix4969 : and02 port map ( Y=>wind_col_in_1_13, A0=>nx7131, A1=>
      cache_data_out_1_13);
   ix4971 : and02 port map ( Y=>wind_col_in_1_14, A0=>nx7131, A1=>
      cache_data_out_1_14);
   ix4973 : and02 port map ( Y=>wind_col_in_1_15, A0=>nx7131, A1=>
      cache_data_out_1_15);
   ix4975 : and02 port map ( Y=>wind_col_in_2_0, A0=>nx7131, A1=>
      cache_data_out_2_0);
   ix4977 : and02 port map ( Y=>wind_col_in_2_1, A0=>nx7131, A1=>
      cache_data_out_2_1);
   ix4979 : and02 port map ( Y=>wind_col_in_2_2, A0=>nx7131, A1=>
      cache_data_out_2_2);
   ix4981 : and02 port map ( Y=>wind_col_in_2_3, A0=>nx6931, A1=>
      cache_data_out_2_3);
   ix4983 : and02 port map ( Y=>wind_col_in_2_4, A0=>nx6931, A1=>
      cache_data_out_2_4);
   ix4985 : and02 port map ( Y=>wind_col_in_2_5, A0=>nx6931, A1=>
      cache_data_out_2_5);
   ix4987 : and02 port map ( Y=>wind_col_in_2_6, A0=>nx6931, A1=>
      cache_data_out_2_6);
   ix4989 : and02 port map ( Y=>wind_col_in_2_7, A0=>nx6931, A1=>
      cache_data_out_2_7);
   ix4991 : and02 port map ( Y=>wind_col_in_2_8, A0=>nx6931, A1=>
      cache_data_out_2_8);
   ix4993 : and02 port map ( Y=>wind_col_in_2_9, A0=>nx6931, A1=>
      cache_data_out_2_9);
   ix4995 : and02 port map ( Y=>wind_col_in_2_10, A0=>nx7133, A1=>
      cache_data_out_2_10);
   ix4997 : and02 port map ( Y=>wind_col_in_2_11, A0=>nx7133, A1=>
      cache_data_out_2_11);
   ix4999 : and02 port map ( Y=>wind_col_in_2_12, A0=>nx7133, A1=>
      cache_data_out_2_12);
   ix5001 : and02 port map ( Y=>wind_col_in_2_13, A0=>nx7133, A1=>
      cache_data_out_2_13);
   ix5003 : and02 port map ( Y=>wind_col_in_2_14, A0=>nx7133, A1=>
      cache_data_out_2_14);
   ix5005 : and02 port map ( Y=>wind_col_in_2_15, A0=>nx7133, A1=>
      cache_data_out_2_15);
   ix5007 : and02 port map ( Y=>wind_col_in_3_0, A0=>nx7133, A1=>
      cache_data_out_3_0);
   ix5009 : and02 port map ( Y=>wind_col_in_3_1, A0=>nx7135, A1=>
      cache_data_out_3_1);
   ix5011 : and02 port map ( Y=>wind_col_in_3_2, A0=>nx7135, A1=>
      cache_data_out_3_2);
   ix5013 : and02 port map ( Y=>wind_col_in_3_3, A0=>nx7135, A1=>
      cache_data_out_3_3);
   ix5015 : and02 port map ( Y=>wind_col_in_3_4, A0=>nx7135, A1=>
      cache_data_out_3_4);
   ix5017 : and02 port map ( Y=>wind_col_in_3_5, A0=>nx7135, A1=>
      cache_data_out_3_5);
   ix5019 : and02 port map ( Y=>wind_col_in_3_6, A0=>nx7135, A1=>
      cache_data_out_3_6);
   ix5021 : and02 port map ( Y=>wind_col_in_3_7, A0=>nx7135, A1=>
      cache_data_out_3_7);
   ix5023 : and02 port map ( Y=>wind_col_in_3_8, A0=>nx7137, A1=>
      cache_data_out_3_8);
   ix5025 : and02 port map ( Y=>wind_col_in_3_9, A0=>nx7137, A1=>
      cache_data_out_3_9);
   ix5027 : and02 port map ( Y=>wind_col_in_3_10, A0=>nx7137, A1=>
      cache_data_out_3_10);
   ix5029 : and02 port map ( Y=>wind_col_in_3_11, A0=>nx7137, A1=>
      cache_data_out_3_11);
   ix5031 : and02 port map ( Y=>wind_col_in_3_12, A0=>nx7137, A1=>
      cache_data_out_3_12);
   ix5033 : and02 port map ( Y=>wind_col_in_3_13, A0=>nx7137, A1=>
      cache_data_out_3_13);
   ix5035 : and02 port map ( Y=>wind_col_in_3_14, A0=>nx7137, A1=>
      cache_data_out_3_14);
   ix5037 : and02 port map ( Y=>wind_col_in_3_15, A0=>nx7139, A1=>
      cache_data_out_3_15);
   ix5039 : and02 port map ( Y=>wind_col_in_4_0, A0=>nx7139, A1=>
      cache_data_out_4_0);
   ix5041 : and02 port map ( Y=>wind_col_in_4_1, A0=>nx7139, A1=>
      cache_data_out_4_1);
   ix5043 : and02 port map ( Y=>wind_col_in_4_2, A0=>nx7139, A1=>
      cache_data_out_4_2);
   ix5045 : and02 port map ( Y=>wind_col_in_4_3, A0=>nx7139, A1=>
      cache_data_out_4_3);
   ix5047 : and02 port map ( Y=>wind_col_in_4_4, A0=>nx7139, A1=>
      cache_data_out_4_4);
   ix5049 : and02 port map ( Y=>wind_col_in_4_5, A0=>nx7139, A1=>
      cache_data_out_4_5);
   ix5051 : and02 port map ( Y=>wind_col_in_4_6, A0=>nx6933, A1=>
      cache_data_out_4_6);
   ix5053 : and02 port map ( Y=>wind_col_in_4_7, A0=>nx6933, A1=>
      cache_data_out_4_7);
   ix5055 : and02 port map ( Y=>wind_col_in_4_8, A0=>nx6933, A1=>
      cache_data_out_4_8);
   ix5057 : and02 port map ( Y=>wind_col_in_4_9, A0=>nx6933, A1=>
      cache_data_out_4_9);
   ix5059 : and02 port map ( Y=>wind_col_in_4_10, A0=>nx6933, A1=>
      cache_data_out_4_10);
   ix5061 : and02 port map ( Y=>wind_col_in_4_11, A0=>nx6933, A1=>
      cache_data_out_4_11);
   ix5063 : and02 port map ( Y=>wind_col_in_4_12, A0=>nx6933, A1=>
      cache_data_out_4_12);
   ix5065 : and02 port map ( Y=>wind_col_in_4_13, A0=>nx2502, A1=>
      cache_data_out_4_13);
   ix5067 : and02 port map ( Y=>wind_col_in_4_14, A0=>nx2502, A1=>
      cache_data_out_4_14);
   ix5069 : and02 port map ( Y=>wind_col_in_4_15, A0=>nx2502, A1=>
      cache_data_out_4_15);
   ix2511 : or03 port map ( Y=>wind_en, A0=>nx4883, A1=>nx7145, A2=>nx1459);
   ix2503 : or03 port map ( Y=>nx2502, A0=>nx4731, A1=>nx4879, A2=>nx7065);
   ix5588 : and03 port map ( Y=>nx5587, A0=>nx6957, A1=>nx7049, A2=>nx7071);
   ix6956 : inv01 port map ( Y=>nx6957, A=>nx6801);
   ix2627 : and02 port map ( Y=>nx2626, A0=>nx6991, A1=>nx7057);
   ix2603 : nand02 port map ( Y=>nx5728, A0=>nx7057, A1=>nx6995);
   ix5592 : nor02_2x port map ( Y=>nx2098, A0=>nx7027, A1=>nx7021);
   ix5599 : and04 port map ( Y=>nx5598, A0=>nx6959, A1=>nx7085, A2=>nx4087, 
      A3=>nx6823);
   ix6958 : inv01 port map ( Y=>nx6959, A=>current_state_6);
   ix1951 : nor02_2x port map ( Y=>nx1950, A0=>nx1930, A1=>nx5197);
   ix5620 : or02 port map ( Y=>nx5619, A0=>nx4423, A1=>nx7357);
   ix5622 : or02 port map ( Y=>nx5621, A0=>nx7357, A1=>nx5194);
   ix3040 : xor2 port map ( Y=>nx3039, A0=>addr1_data_0, A1=>nx7111);
   ix5626 : or03 port map ( Y=>nx6905, A0=>nx6993, A1=>nx6711, A2=>nx2706);
   ix2719 : nor02ii port map ( Y=>nx6813, A0=>nx7111, A1=>nx4665);
   ix3000 : mux21 port map ( Y=>nx2999, A0=>write_offset_data_out_0, A1=>
      nx5632, S0=>nx7071);
   ix5637 : or02 port map ( Y=>nx5636, A0=>nx5632, A1=>nx7358);
   ix3030 : xor2 port map ( Y=>nx3029, A0=>img_addr_offset_0, A1=>nx7003);
   ix2675 : nor02_2x port map ( Y=>nx6805, A0=>nx1419, A1=>reset);
   ix3020 : mux21_ni port map ( Y=>nx3019, A0=>nx5647, A1=>img_base_addr_0, 
      S0=>nx7011);
   ix3010 : mux21 port map ( Y=>nx3009, A0=>nx5647, A1=>nx7358, S0=>nx7117);
   ix5654 : xnor2 port map ( Y=>nx5653, A0=>nx4433, A1=>nx4039);
   ix2641 : nor02ii port map ( Y=>nx2640, A0=>nx2636, A1=>current_state_12);
   ix2637 : xnor2 port map ( Y=>nx2636, A0=>nx4099, A1=>nflt_layer_out_0);
   ix5658 : xnor2 port map ( Y=>nx5657, A0=>nx4459, A1=>nx4053);
   ix5660 : xor2 port map ( Y=>nx5659, A0=>nx4485, A1=>nflt_layer_out_3);
   ix5674 : xnor2 port map ( Y=>nx5673, A0=>nx5677, A1=>nx5700);
   ix3090 : mux21 port map ( Y=>nx3089, A0=>nx5679, A1=>nx5677, S0=>nx7011);
   ix3080 : mux21_ni port map ( Y=>nx3079, A0=>write_base_prev_data_out_1, 
      A1=>write_base_data_out_1, S0=>nx7117);
   ix3050 : mux21 port map ( Y=>nx3049, A0=>nx5687, A1=>nx7359, S0=>nx7095);
   ix5693 : nor02ii port map ( Y=>nx5692, A0=>write_base_prev_data_out_1, A1
      =>nx5647);
   ix3100 : mux21 port map ( Y=>nx3099, A0=>nx5700, A1=>nx5696, S0=>nx7003);
   ix5704 : xnor2 port map ( Y=>nx5703, A0=>nx5707, A1=>nx7359);
   ix3070 : ao32 port map ( Y=>nx3069, A0=>nx6961, A1=>nx7057, A2=>nx6995, 
      B0=>bias_offset_data_out_1, B1=>nx7071);
   ix6960 : inv01 port map ( Y=>nx6961, A=>nx4287);
   ix5715 : xnor2 port map ( Y=>nx5714, A0=>nx7359, A1=>nx5202);
   ix3060 : mux21 port map ( Y=>nx3059, A0=>nx5722, A1=>nx5718, S0=>nx7111);
   ix2605 : nor02ii port map ( Y=>nx6793, A0=>nx6983, A1=>nx7071);
   ix5738 : xnor2 port map ( Y=>nx5737, A0=>nx5758, A1=>nx5762);
   ix3150 : mux21_ni port map ( Y=>nx3149, A0=>nx2956, A1=>img_base_addr_2, 
      S0=>nx7011);
   ix3140 : mux21 port map ( Y=>nx3139, A0=>nx5742, A1=>nx7361, S0=>nx7117);
   ix3110 : mux21 port map ( Y=>nx3109, A0=>nx5749, A1=>nx7361, S0=>nx7095);
   ix3160 : mux21_ni port map ( Y=>nx3159, A0=>img_addr_offset_2, A1=>nx2970, 
      S0=>nx7003);
   ix2971 : xor2 port map ( Y=>nx2970, A0=>nx5762, A1=>nx5698);
   ix5768 : xnor2 port map ( Y=>nx5767, A0=>nx5771, A1=>nx7361);
   ix3130 : ao32 port map ( Y=>nx3129, A0=>nx6963, A1=>nx7059, A2=>nx6995, 
      B0=>bias_offset_data_out_2, B1=>nx7071);
   ix6962 : inv01 port map ( Y=>nx6963, A=>nx4281);
   ix5778 : xnor2 port map ( Y=>nx5777, A0=>nx7362, A1=>nx4277);
   ix5784 : xnor2 port map ( Y=>nx5783, A0=>nx7362, A1=>nx5208);
   ix3120 : mux21_ni port map ( Y=>nx3119, A0=>addr1_data_2, A1=>nx2904, S0
      =>nx7111);
   ix3210 : mux21_ni port map ( Y=>nx3209, A0=>nx3100, A1=>img_base_addr_3, 
      S0=>nx7011);
   ix3200 : mux21_ni port map ( Y=>nx3199, A0=>write_base_prev_data_out_3, 
      A1=>write_base_data_out_3, S0=>nx7117);
   ix3170 : mux21_ni port map ( Y=>nx3169, A0=>nx3006, A1=>
      write_base_data_out_3, S0=>nx7095);
   ix5806 : xor2 port map ( Y=>nx5805, A0=>new_size_squared_out_3, A1=>
      nx5807);
   ix3220 : mux21_ni port map ( Y=>nx3219, A0=>img_addr_offset_3, A1=>nx3114, 
      S0=>nx7003);
   ix5821 : xor2 port map ( Y=>nx5820, A0=>bias_offset_data_out_3, A1=>
      nx5807);
   ix3190 : mux21_ni port map ( Y=>nx3189, A0=>nx802, A1=>
      bias_offset_data_out_3, S0=>nx7071);
   ix803 : xor2 port map ( Y=>nx802, A0=>nx4271, A1=>nx4299);
   ix5835 : xnor2 port map ( Y=>nx5834, A0=>nx5807, A1=>nx5218);
   ix3180 : mux21_ni port map ( Y=>nx3179, A0=>addr1_data_3, A1=>nx3048, S0
      =>nx7111);
   ix5851 : xnor2 port map ( Y=>nx5850, A0=>nx5807, A1=>nx4271);
   ix5860 : xnor2 port map ( Y=>nx5859, A0=>nx5882, A1=>nx5888);
   ix3270 : mux21_ni port map ( Y=>nx3269, A0=>nx3248, A1=>img_base_addr_4, 
      S0=>nx7011);
   ix3260 : mux21 port map ( Y=>nx3259, A0=>nx5864, A1=>nx5869, S0=>nx7117);
   ix3230 : mux21 port map ( Y=>nx3229, A0=>nx5871, A1=>nx5869, S0=>nx7095);
   ix5877 : xnor2 port map ( Y=>nx5876, A0=>nx4391, A1=>nx5869);
   ix3280 : mux21_ni port map ( Y=>nx3279, A0=>img_addr_offset_4, A1=>nx3262, 
      S0=>nx7003);
   ix3257 : nor02ii port map ( Y=>nx3256, A0=>nx5886, A1=>img_addr_offset_4
   );
   ix5896 : xnor2 port map ( Y=>nx5895, A0=>nx5900, A1=>nx5869);
   ix3250 : mux21_ni port map ( Y=>nx3249, A0=>nx828, A1=>
      bias_offset_data_out_4, S0=>nx7071);
   ix3240 : mux21_ni port map ( Y=>nx3239, A0=>addr1_data_4, A1=>nx3196, S0
      =>nx7111);
   ix3191 : nor02ii port map ( Y=>nx3190, A0=>nx5906, A1=>addr1_data_4);
   ix5914 : xnor2 port map ( Y=>nx5913, A0=>nx5869, A1=>nx4257);
   ix5918 : xor2 port map ( Y=>nx5917, A0=>nx5869, A1=>nx3170);
   ix5926 : xor2 port map ( Y=>nx5925, A0=>img_base_addr_5, A1=>nx5947);
   ix3330 : mux21_ni port map ( Y=>nx3329, A0=>nx3388, A1=>img_base_addr_5, 
      S0=>nx7011);
   ix3320 : mux21_ni port map ( Y=>nx3319, A0=>write_base_prev_data_out_5, 
      A1=>write_base_data_out_5, S0=>nx7117);
   ix3290 : mux21_ni port map ( Y=>nx3289, A0=>nx3298, A1=>
      write_base_data_out_5, S0=>nx7095);
   ix5937 : xor2 port map ( Y=>nx5936, A0=>new_size_squared_out_5, A1=>
      nx5938);
   ix3340 : mux21 port map ( Y=>nx3339, A0=>nx5947, A1=>nx5943, S0=>nx7005);
   ix5952 : xnor2 port map ( Y=>nx5951, A0=>nx5955, A1=>nx5938);
   ix3310 : ao32 port map ( Y=>nx3309, A0=>nx6965, A1=>nx7059, A2=>nx6995, 
      B0=>bias_offset_data_out_5, B1=>nx7073);
   ix6964 : inv01 port map ( Y=>nx6965, A=>nx4253);
   ix3300 : mux21 port map ( Y=>nx3299, A0=>nx5965, A1=>nx5961, S0=>nx7111);
   ix5972 : xnor2 port map ( Y=>nx5971, A0=>nx5938, A1=>nx4251);
   ix3319 : xor2 port map ( Y=>nx3318, A0=>nx5938, A1=>nx5977);
   ix5987 : xnor2 port map ( Y=>nx5986, A0=>nx6009, A1=>nx6013);
   ix3390 : mux21_ni port map ( Y=>nx3389, A0=>nx3528, A1=>img_base_addr_6, 
      S0=>nx7011);
   ix3380 : mux21 port map ( Y=>nx3379, A0=>nx5991, A1=>nx5996, S0=>nx7117);
   ix3350 : mux21 port map ( Y=>nx3349, A0=>nx5998, A1=>nx5996, S0=>nx7095);
   ix6004 : xnor2 port map ( Y=>nx6003, A0=>nx4377, A1=>nx5996);
   ix3400 : mux21_ni port map ( Y=>nx3399, A0=>img_addr_offset_6, A1=>nx3542, 
      S0=>nx7005);
   ix3537 : nor02ii port map ( Y=>nx3536, A0=>nx5945, A1=>img_addr_offset_6
   );
   ix6021 : xnor2 port map ( Y=>nx6020, A0=>nx6025, A1=>nx5996);
   ix3370 : mux21_ni port map ( Y=>nx3369, A0=>nx874, A1=>
      bias_offset_data_out_6, S0=>nx7073);
   ix3360 : mux21_ni port map ( Y=>nx3359, A0=>addr1_data_6, A1=>nx3476, S0
      =>nx7113);
   ix3477 : xor2 port map ( Y=>nx3476, A0=>nx6031, A1=>nx5963);
   ix6035 : xnor2 port map ( Y=>nx6034, A0=>nx5996, A1=>nx4239);
   ix3313 : nor02ii port map ( Y=>nx3312, A0=>nx5977, A1=>
      write_base_data_out_5);
   ix6050 : xor2 port map ( Y=>nx6049, A0=>img_base_addr_7, A1=>nx6071);
   ix3450 : mux21_ni port map ( Y=>nx3449, A0=>nx3668, A1=>img_base_addr_7, 
      S0=>nx7013);
   ix3440 : mux21_ni port map ( Y=>nx3439, A0=>write_base_prev_data_out_7, 
      A1=>write_base_data_out_7, S0=>nx7119);
   ix3410 : mux21_ni port map ( Y=>nx3409, A0=>nx3578, A1=>
      write_base_data_out_7, S0=>nx7097);
   ix6061 : xor2 port map ( Y=>nx6060, A0=>new_size_squared_out_7, A1=>
      nx6062);
   ix3460 : mux21 port map ( Y=>nx3459, A0=>nx6071, A1=>nx6067, S0=>nx7005);
   ix6076 : xnor2 port map ( Y=>nx6075, A0=>nx6079, A1=>nx6062);
   ix3430 : ao32 port map ( Y=>nx3429, A0=>nx6967, A1=>nx7059, A2=>nx6995, 
      B0=>bias_offset_data_out_7, B1=>nx7073);
   ix6966 : inv01 port map ( Y=>nx6967, A=>nx4235);
   ix3420 : mux21 port map ( Y=>nx3419, A0=>nx6090, A1=>nx6085, S0=>nx7113);
   ix3471 : nor02ii port map ( Y=>nx3470, A0=>nx5963, A1=>addr1_data_6);
   ix3593 : nor02ii port map ( Y=>nx3592, A0=>nx6042, A1=>
      write_base_data_out_7);
   ix6101 : xnor2 port map ( Y=>nx6100, A0=>nx6062, A1=>nx4229);
   ix6110 : xnor2 port map ( Y=>nx6109, A0=>nx6132, A1=>nx6136);
   ix3510 : mux21_ni port map ( Y=>nx3509, A0=>nx3808, A1=>img_base_addr_8, 
      S0=>nx7013);
   ix3500 : mux21 port map ( Y=>nx3499, A0=>nx6114, A1=>nx6119, S0=>nx7119);
   ix3470 : mux21 port map ( Y=>nx3469, A0=>nx6121, A1=>nx6119, S0=>nx7097);
   ix6127 : xnor2 port map ( Y=>nx6126, A0=>nx4363, A1=>nx6119);
   ix3520 : mux21_ni port map ( Y=>nx3519, A0=>img_addr_offset_8, A1=>nx3822, 
      S0=>nx7005);
   ix3817 : nor02ii port map ( Y=>nx3816, A0=>nx6069, A1=>img_addr_offset_8
   );
   ix6144 : xnor2 port map ( Y=>nx6143, A0=>nx6148, A1=>nx6119);
   ix3490 : mux21_ni port map ( Y=>nx3489, A0=>nx924, A1=>
      bias_offset_data_out_8, S0=>nx7073);
   ix3480 : mux21_ni port map ( Y=>nx3479, A0=>addr1_data_8, A1=>nx3756, S0
      =>nx7113);
   ix3757 : xor2 port map ( Y=>nx3756, A0=>nx6154, A1=>nx6088);
   ix6158 : xnor2 port map ( Y=>nx6157, A0=>nx6119, A1=>nx4217);
   ix6172 : xor2 port map ( Y=>nx6171, A0=>img_base_addr_9, A1=>nx6193);
   ix3570 : mux21_ni port map ( Y=>nx3569, A0=>nx3948, A1=>img_base_addr_9, 
      S0=>nx7013);
   ix3560 : mux21_ni port map ( Y=>nx3559, A0=>write_base_prev_data_out_9, 
      A1=>write_base_data_out_9, S0=>nx7119);
   ix3530 : mux21_ni port map ( Y=>nx3529, A0=>nx3858, A1=>
      write_base_data_out_9, S0=>nx7097);
   ix6183 : xor2 port map ( Y=>nx6182, A0=>new_size_squared_out_9, A1=>
      nx6184);
   ix3580 : mux21 port map ( Y=>nx3579, A0=>nx6193, A1=>nx6189, S0=>nx7005);
   ix6198 : xnor2 port map ( Y=>nx6197, A0=>nx6201, A1=>nx6184);
   ix3550 : ao32 port map ( Y=>nx3549, A0=>nx6969, A1=>nx7059, A2=>nx6995, 
      B0=>bias_offset_data_out_9, B1=>nx7073);
   ix6968 : inv01 port map ( Y=>nx6969, A=>nx4213);
   ix3540 : mux21 port map ( Y=>nx3539, A0=>nx6212, A1=>nx6207, S0=>nx7113);
   ix3751 : nor02ii port map ( Y=>nx3750, A0=>nx6088, A1=>addr1_data_8);
   ix3873 : nor02ii port map ( Y=>nx3872, A0=>nx6164, A1=>
      write_base_data_out_9);
   ix6223 : xnor2 port map ( Y=>nx6222, A0=>nx6184, A1=>nx4301);
   ix6232 : xnor2 port map ( Y=>nx6231, A0=>nx6254, A1=>nx6258);
   ix3630 : mux21_ni port map ( Y=>nx3629, A0=>nx4088, A1=>img_base_addr_10, 
      S0=>nx7013);
   ix3620 : mux21 port map ( Y=>nx3619, A0=>nx6236, A1=>nx6241, S0=>nx7119);
   ix3590 : mux21 port map ( Y=>nx3589, A0=>nx6243, A1=>nx6241, S0=>nx7097);
   ix6249 : xnor2 port map ( Y=>nx6248, A0=>nx4349, A1=>nx6241);
   ix3640 : mux21_ni port map ( Y=>nx3639, A0=>img_addr_offset_10, A1=>
      nx4102, S0=>nx7005);
   ix4097 : nor02ii port map ( Y=>nx4096, A0=>nx6191, A1=>img_addr_offset_10
   );
   ix6266 : xnor2 port map ( Y=>nx6265, A0=>nx6270, A1=>nx6241);
   ix3610 : mux21_ni port map ( Y=>nx3609, A0=>nx970, A1=>
      bias_offset_data_out_10, S0=>nx7073);
   ix3600 : mux21_ni port map ( Y=>nx3599, A0=>addr1_data_10, A1=>nx4036, S0
      =>nx7113);
   ix4037 : xor2 port map ( Y=>nx4036, A0=>nx6276, A1=>nx6210);
   ix6280 : xnor2 port map ( Y=>nx6279, A0=>nx6241, A1=>nx4200);
   ix6294 : xor2 port map ( Y=>nx6293, A0=>img_base_addr_11, A1=>nx6315);
   ix3690 : mux21_ni port map ( Y=>nx3689, A0=>nx4228, A1=>img_base_addr_11, 
      S0=>nx7013);
   ix3680 : mux21_ni port map ( Y=>nx3679, A0=>write_base_prev_data_out_11, 
      A1=>write_base_data_out_11, S0=>nx7119);
   ix3650 : mux21_ni port map ( Y=>nx3649, A0=>nx4138, A1=>
      write_base_data_out_11, S0=>nx7097);
   ix6305 : xor2 port map ( Y=>nx6304, A0=>new_size_squared_out_11, A1=>
      nx6306);
   ix3700 : mux21 port map ( Y=>nx3699, A0=>nx6315, A1=>nx6311, S0=>nx7005);
   ix6320 : xnor2 port map ( Y=>nx6319, A0=>nx6323, A1=>nx6306);
   ix3670 : ao32 port map ( Y=>nx3669, A0=>nx6971, A1=>nx7059, A2=>nx6995, 
      B0=>bias_offset_data_out_11, B1=>nx7073);
   ix6970 : inv01 port map ( Y=>nx6971, A=>nx4197);
   ix3660 : mux21 port map ( Y=>nx3659, A0=>nx6334, A1=>nx6329, S0=>nx7113);
   ix4031 : nor02ii port map ( Y=>nx4030, A0=>nx6210, A1=>addr1_data_10);
   ix4153 : nor02ii port map ( Y=>nx4152, A0=>nx6286, A1=>
      write_base_data_out_11);
   ix6345 : xnor2 port map ( Y=>nx6344, A0=>nx6306, A1=>nx4303);
   ix6354 : xnor2 port map ( Y=>nx6353, A0=>nx6376, A1=>nx6380);
   ix3750 : mux21_ni port map ( Y=>nx3749, A0=>nx4368, A1=>img_base_addr_12, 
      S0=>nx7013);
   ix3740 : mux21 port map ( Y=>nx3739, A0=>nx6358, A1=>nx7363, S0=>nx7119);
   ix3710 : mux21 port map ( Y=>nx3709, A0=>nx6365, A1=>nx7363, S0=>nx7097);
   ix3760 : mux21_ni port map ( Y=>nx3759, A0=>img_addr_offset_12, A1=>
      nx4382, S0=>nx7007);
   ix4377 : nor02ii port map ( Y=>nx4376, A0=>nx6313, A1=>img_addr_offset_12
   );
   ix6388 : xnor2 port map ( Y=>nx6387, A0=>nx6392, A1=>nx7363);
   ix3730 : mux21_ni port map ( Y=>nx3729, A0=>nx1018, A1=>
      bias_offset_data_out_12, S0=>nx7075);
   ix3720 : mux21_ni port map ( Y=>nx3719, A0=>addr1_data_12, A1=>nx4316, S0
      =>nx7113);
   ix4317 : xor2 port map ( Y=>nx4316, A0=>nx6398, A1=>nx6332);
   ix6409 : xnor2 port map ( Y=>nx6408, A0=>nx7363, A1=>nx4183);
   ix6416 : xor2 port map ( Y=>nx6415, A0=>img_base_addr_13, A1=>nx6437);
   ix3810 : mux21_ni port map ( Y=>nx3809, A0=>nx4508, A1=>img_base_addr_13, 
      S0=>nx7013);
   ix3800 : mux21_ni port map ( Y=>nx3799, A0=>write_base_prev_data_out_13, 
      A1=>write_base_data_out_13, S0=>nx7119);
   ix3770 : mux21_ni port map ( Y=>nx3769, A0=>nx4418, A1=>
      write_base_data_out_13, S0=>nx7097);
   ix6427 : xor2_2x port map ( Y=>nx6426, A0=>new_size_squared_out_13, A1=>
      nx6428);
   ix3820 : mux21 port map ( Y=>nx3819, A0=>nx6437, A1=>nx6433, S0=>nx7007);
   ix6442 : xnor2 port map ( Y=>nx6441, A0=>nx6445, A1=>nx6428);
   ix3790 : ao32 port map ( Y=>nx3789, A0=>nx6973, A1=>nx7059, A2=>nx6997, 
      B0=>bias_offset_data_out_13, B1=>nx7075);
   ix6972 : inv01 port map ( Y=>nx6973, A=>nx4180);
   ix3780 : mux21 port map ( Y=>nx3779, A0=>nx6456, A1=>nx6451, S0=>nx7115);
   ix4311 : nor02ii port map ( Y=>nx4310, A0=>nx6332, A1=>addr1_data_12);
   ix4433 : nor02ii port map ( Y=>nx4432, A0=>nx6404, A1=>
      write_base_data_out_13);
   ix6467 : xnor2 port map ( Y=>nx6466, A0=>nx6428, A1=>nx4305);
   ix6476 : xnor2 port map ( Y=>nx6475, A0=>nx6496, A1=>nx6500);
   ix3870 : mux21_ni port map ( Y=>nx3869, A0=>nx4648, A1=>img_base_addr_14, 
      S0=>nx7015);
   ix4649 : xnor2 port map ( Y=>nx4648, A0=>nx6493, A1=>nx6494);
   ix3860 : mux21 port map ( Y=>nx3859, A0=>nx6493, A1=>nx7365, S0=>nx7121);
   ix3830 : mux21 port map ( Y=>nx3829, A0=>nx6486, A1=>nx7365, S0=>nx7099);
   ix3880 : mux21_ni port map ( Y=>nx3879, A0=>img_addr_offset_14, A1=>
      nx4662, S0=>nx7007);
   ix4663 : xor2 port map ( Y=>nx4662, A0=>nx6500, A1=>nx6435);
   ix6506 : xnor2 port map ( Y=>nx6505, A0=>nx6510, A1=>nx7365);
   ix3850 : mux21_ni port map ( Y=>nx3849, A0=>nx1064, A1=>
      bias_offset_data_out_14, S0=>nx7075);
   ix1065 : xor2 port map ( Y=>nx1064, A0=>nx4167, A1=>nx4175);
   ix3840 : mux21_ni port map ( Y=>nx3839, A0=>addr1_data_14, A1=>nx4596, S0
      =>nx7115);
   ix4597 : xor2 port map ( Y=>nx4596, A0=>nx6516, A1=>nx6454);
   ix6521 : xor2 port map ( Y=>nx6520, A0=>nx7365, A1=>nx4432);
   ix6525 : xnor2 port map ( Y=>nx6524, A0=>nx7366, A1=>nx4167);
   ix6544 : xor2 port map ( Y=>nx6543, A0=>img_base_addr_15, A1=>nx6558);
   ix3930 : mux21_ni port map ( Y=>nx3929, A0=>nx4764, A1=>img_base_addr_15, 
      S0=>nx7015);
   ix3920 : mux21_ni port map ( Y=>nx3919, A0=>write_base_prev_data_out_15, 
      A1=>write_base_data_out_15, S0=>nx7121);
   ix3940 : mux21 port map ( Y=>nx3939, A0=>nx6558, A1=>nx6555, S0=>nx7007);
   ix6556 : xor2 port map ( Y=>nx6555, A0=>nx6558, A1=>nx4656);
   ix4657 : nor02ii port map ( Y=>nx4656, A0=>nx6435, A1=>img_addr_offset_14
   );
   ix4735 : xor2 port map ( Y=>nx4734, A0=>write_base_data_out_15, A1=>
      write_offset_data_out_15);
   ix3910 : mux21 port map ( Y=>nx3909, A0=>nx6572, A1=>nx6569, S0=>nx7115);
   ix6570 : xor2 port map ( Y=>nx6569, A0=>nx6572, A1=>nx4590);
   ix4591 : nor02ii port map ( Y=>nx4590, A0=>nx6454, A1=>addr1_data_14);
   ix6577 : xor2 port map ( Y=>nx6576, A0=>nx6580, A1=>
      write_base_data_out_15);
   ix3890 : ao32 port map ( Y=>nx3889, A0=>nx6975, A1=>nx7059, A2=>nx6997, 
      B0=>bias_offset_data_out_15, B1=>nx7075);
   ix6974 : inv01 port map ( Y=>nx6975, A=>nx4163);
   ix6758 : nor02ii port map ( Y=>nx6759, A0=>nx6929, A1=>current_state_12);
   ix6760 : nor02ii port map ( Y=>nx6761, A0=>nx6929, A1=>current_state_12);
   ix6800 : and02 port map ( Y=>nx6801, A0=>nx6991, A1=>nx7061);
   ix6802 : and02 port map ( Y=>nx6803, A0=>nx6991, A1=>nx7061);
   ix6976 : inv02 port map ( Y=>nx6977, A=>nx4883);
   ix6978 : inv02 port map ( Y=>nx6979, A=>nx4883);
   ix6980 : inv01 port map ( Y=>nx6981, A=>nx6829);
   ix6982 : inv01 port map ( Y=>nx6983, A=>nx6829);
   ix6984 : inv01 port map ( Y=>nx6985, A=>nx6851);
   ix6986 : inv01 port map ( Y=>nx6987, A=>nx6851);
   ix6988 : inv01 port map ( Y=>nx6989, A=>nx6851);
   ix6990 : inv01 port map ( Y=>nx6991, A=>nx6851);
   ix6992 : buf02 port map ( Y=>nx6993, A=>nx2084);
   ix6994 : inv02 port map ( Y=>nx6995, A=>nx6897);
   ix6996 : inv02 port map ( Y=>nx6997, A=>nx6897);
   ix6998 : inv02 port map ( Y=>nx6999, A=>nx7107);
   ix7000 : inv02 port map ( Y=>nx7001, A=>nx7107);
   ix7002 : inv02 port map ( Y=>nx7003, A=>nx7107);
   ix7004 : inv02 port map ( Y=>nx7005, A=>nx6871);
   ix7006 : inv02 port map ( Y=>nx7007, A=>nx6871);
   ix7008 : inv02 port map ( Y=>nx7009, A=>nx6665);
   ix7010 : inv02 port map ( Y=>nx7011, A=>nx6665);
   ix7012 : inv02 port map ( Y=>nx7013, A=>nx6665);
   ix7014 : inv02 port map ( Y=>nx7015, A=>nx6665);
   ix7016 : buf02 port map ( Y=>nx7017, A=>nx4033);
   ix7018 : inv02 port map ( Y=>nx7019, A=>nx1528);
   ix7020 : inv01 port map ( Y=>nx7021, A=>nx6705);
   ix7022 : inv02 port map ( Y=>nx7023, A=>nx6749);
   ix7024 : inv02 port map ( Y=>nx7025, A=>nx6749);
   ix7026 : inv02 port map ( Y=>nx7027, A=>nx6749);
   ix7032 : inv02 port map ( Y=>nx7033, A=>nx6685);
   ix7034 : inv02 port map ( Y=>nx7035, A=>nx6685);
   ix7036 : inv02 port map ( Y=>nx7037, A=>nx1429);
   ix7038 : inv02 port map ( Y=>nx7039, A=>nx1429);
   ix7040 : inv02 port map ( Y=>nx7041, A=>nx1429);
   ix7042 : inv02 port map ( Y=>nx7043, A=>argmax_ready_EXMPLR);
   ix7048 : inv02 port map ( Y=>nx7049, A=>argmax_ready_EXMPLR);
   ix7050 : inv01 port map ( Y=>nx7051, A=>nx5243);
   ix7052 : inv02 port map ( Y=>nx7053, A=>nx7051);
   ix7054 : inv02 port map ( Y=>nx7055, A=>nx7051);
   ix7056 : inv02 port map ( Y=>nx7057, A=>nx7051);
   ix7058 : inv02 port map ( Y=>nx7059, A=>nx7051);
   ix7060 : inv02 port map ( Y=>nx7061, A=>nx7051);
   ix7064 : inv02 port map ( Y=>nx7065, A=>comp_unit_flt_size_EXMPLR);
   ix7070 : inv02 port map ( Y=>nx7071, A=>nx6787);
   ix7072 : inv02 port map ( Y=>nx7073, A=>nx6787);
   ix7074 : inv02 port map ( Y=>nx7075, A=>nx6787);
   ix7076 : inv01 port map ( Y=>nx7077, A=>nx7293);
   ix7078 : inv01 port map ( Y=>nx7079, A=>nx7293);
   ix7080 : inv02 port map ( Y=>nx7081, A=>current_state_7);
   ix7082 : inv02 port map ( Y=>nx7083, A=>current_state_7);
   ix7084 : inv02 port map ( Y=>nx7085, A=>current_state_7);
   ix7086 : inv02 port map ( Y=>nx7087, A=>nx6731);
   ix7088 : inv02 port map ( Y=>nx7089, A=>nx6731);
   ix7090 : buf02 port map ( Y=>nx7091, A=>nx6759);
   ix7092 : buf02 port map ( Y=>nx7093, A=>nx6761);
   ix7094 : inv02 port map ( Y=>nx7095, A=>nx2580);
   ix7096 : inv02 port map ( Y=>nx7097, A=>nx2580);
   ix7098 : inv02 port map ( Y=>nx7099, A=>nx2580);
   ix7100 : inv02 port map ( Y=>nx7101, A=>nx5099);
   ix7102 : inv02 port map ( Y=>nx7103, A=>nx5099);
   ix7104 : inv02 port map ( Y=>nx7105, A=>nx5099);
   ix7106 : inv02 port map ( Y=>nx7107, A=>nx2536);
   ix7108 : inv01 port map ( Y=>nx7109, A=>nx6905);
   ix7110 : inv02 port map ( Y=>nx7111, A=>nx7109);
   ix7112 : inv02 port map ( Y=>nx7113, A=>nx7109);
   ix7114 : inv02 port map ( Y=>nx7115, A=>nx7109);
   ix7116 : inv02 port map ( Y=>nx7117, A=>nx5651);
   ix7118 : inv02 port map ( Y=>nx7119, A=>nx5651);
   ix7120 : inv02 port map ( Y=>nx7121, A=>nx5651);
   ix7122 : inv01 port map ( Y=>nx7123, A=>nx7145);
   ix7124 : inv01 port map ( Y=>nx7125, A=>nx7145);
   ix7126 : inv01 port map ( Y=>nx7127, A=>nx7145);
   ix7128 : inv01 port map ( Y=>nx7129, A=>nx7145);
   ix7130 : inv01 port map ( Y=>nx7131, A=>nx5501);
   ix7132 : inv01 port map ( Y=>nx7133, A=>nx5501);
   ix7134 : inv01 port map ( Y=>nx7135, A=>nx5501);
   ix7136 : inv01 port map ( Y=>nx7137, A=>nx5501);
   ix7138 : inv01 port map ( Y=>nx7139, A=>nx5501);
   ix7144 : inv01 port map ( Y=>nx7145, A=>nx2502);
   ix291 : oai21 port map ( Y=>filter_ready_out_EXMPLR, A0=>nx7029, A1=>
      nx4593, B0=>nx4665);
   ix7028 : inv02 port map ( Y=>nx7029, A=>nx6711);
   ix4594 : inv01 port map ( Y=>nx4593, A=>nx286);
   ix4666 : or02 port map ( Y=>nx4665, A0=>nx4637, A1=>nx7021);
   ix7062 : inv02 port map ( Y=>nx7063, A=>comp_unit_flt_size_EXMPLR);
   ix273 : inv01 port map ( Y=>comp_unit_flt_size_EXMPLR, A=>nx5482);
   ix7030 : inv02 port map ( Y=>nx7031, A=>nx6711);
   ix6710 : inv02 port map ( Y=>nx6711, A=>nx4589);
   ix7368 : buf04 port map ( Y=>nx7293, A=>filter_ready_out_EXMPLR);
   ix7369 : buf04 port map ( Y=>nx7294, A=>nx7063);
   ix7370 : buf04 port map ( Y=>nx7295, A=>nx7031);
   ix7371 : inv02 port map ( Y=>nx7296, A=>new_size_squared_out_15);
   ix7372 : inv02 port map ( Y=>nx7297, A=>write_base_data_out_15);
   ix7373 : oai32 port map ( Y=>nx7298, A0=>nx7099, A1=>nx7296, A2=>
      write_base_data_out_15, B0=>nx7297, B1=>new_size_squared_out_15);
   ix7374 : and02 port map ( Y=>nx7299, A0=>nx7364, A1=>nx4335);
   ix7375 : nor02_2x port map ( Y=>nx7300, A0=>nx7364, A1=>nx4335);
   ix7376 : and02 port map ( Y=>nx7301, A0=>nx7366, A1=>nx4320);
   ix7377 : inv02 port map ( Y=>nx7302, A=>write_base_data_out_13);
   ix7378 : inv02 port map ( Y=>nx7303, A=>new_size_squared_out_13);
   ix7379 : inv02 port map ( Y=>nx7304, A=>nx7099);
   ix7380 : aoi32 port map ( Y=>nx7305, A0=>nx7304, A1=>nx7297, A2=>nx7296, 
      B0=>write_base_data_out_15, B1=>new_size_squared_out_15);
   reg_nx3899 : ao221 port map ( Y=>nx3899, A0=>nx7298, A1=>NOT_nx4700, B0=>
      write_base_data_out_15, B1=>nx7099, C0=>nx7350);
   ix7381 : and02 port map ( Y=>nx7306, A0=>write_base_data_out_13, A1=>
      new_size_squared_out_13);
   ix7382 : inv02 port map ( Y=>nx7307, A=>nx6426);
   reg_nx6488 : oai32 port map ( Y=>nx6488, A0=>nx7306, A1=>nx7354, A2=>
      nx7300, B0=>nx7307, B1=>nx7306);
   ix7383 : inv01 port map ( Y=>nx7308, A=>nx7366);
   ix7384 : inv02 port map ( Y=>nx7309, A=>nx4320);
   reg_nx6491 : oai22 port map ( Y=>nx6491, A0=>nx7308, A1=>nx7309, B0=>
      nx7366, B1=>nx4320);
   reg_nx4414 : oai22 port map ( Y=>nx4414, A0=>nx7364, A1=>nx4335, B0=>
      nx7299, B1=>nx7445);
   ix7385 : inv02 port map ( Y=>nx7310, A=>nx7364);
   ix7386 : inv02 port map ( Y=>nx7311, A=>nx4335);
   reg_nx6370 : oai22 port map ( Y=>nx6370, A0=>nx7310, A1=>nx7311, B0=>
      nx7364, B1=>nx4335);
   ix7387 : inv01 port map ( Y=>nx7312, A=>nx7362);
   ix7388 : inv01 port map ( Y=>nx7313, A=>nx4407);
   ix7389 : nand02_2x port map ( Y=>nx7314, A0=>nx7362, A1=>nx4407);
   ix7390 : inv01 port map ( Y=>nx7315, A=>nx7359);
   ix7391 : nand03_2x port map ( Y=>nx7316, A0=>new_size_squared_out_0, A1=>
      nx6775, A2=>nx7315);
   ix7392 : inv01 port map ( Y=>nx7317, A=>new_size_squared_out_1);
   ix7393 : nand02_2x port map ( Y=>nx7318, A0=>new_size_squared_out_1, A1=>
      nx7315);
   ix7394 : nand03_2x port map ( Y=>nx7319, A0=>nx7318, A1=>
      new_size_squared_out_0, A2=>nx6775);
   ix7395 : inv01 port map ( Y=>nx7320, A=>write_base_data_out_1);
   ix7396 : aoi22 port map ( Y=>nx7321, A0=>nx7316, A1=>nx7317, B0=>nx7319, 
      B1=>nx7320);
   ix7397 : aoi22 port map ( Y=>nx7322, A0=>nx7312, A1=>nx7313, B0=>nx7314, 
      B1=>nx7321);
   reg_nx3002 : inv01 port map ( Y=>nx3002, A=>nx7322);
   ix7398 : inv01 port map ( Y=>nx7323, A=>nx7322);
   reg_nx5751 : inv01 port map ( Y=>nx5751, A=>nx7321);
   reg_nx5754 : oai22 port map ( Y=>nx5754, A0=>nx7312, A1=>nx7313, B0=>
      nx7362, B1=>nx4407);
   reg_nx5689 : oai22 port map ( Y=>nx5689, A0=>nx7315, A1=>
      new_size_squared_out_1, B0=>nx7317, B1=>nx7360);
   ix7399 : inv01 port map ( Y=>nx7324, A=>mem_data_in(3));
   reg_argmax_data_out_3 : nor03_2x port map ( Y=>argmax_data_out(3), A0=>
      nx7338, A1=>nx7324, A2=>nx7340);
   reg_nx5191 : inv02 port map ( Y=>nx5191, A=>argmax_ready_EXMPLR);
   reg_argmax_ready : inv01 port map ( Y=>argmax_ready_dup0, A=>
      argmax_ready_EXMPLR);
   ix7400 : inv01 port map ( Y=>nx7325, A=>nx7367);
   ix7401 : inv01 port map ( Y=>nx7326, A=>nx7367);
   ix7402 : inv01 port map ( Y=>nx7327, A=>nx7367);
   ix7403 : inv01 port map ( Y=>nx7328, A=>nx7367);
   reg_nx1930 : inv01 port map ( Y=>nx1930, A=>nx7338);
   ix7404 : nand02_2x port map ( Y=>nx7329, A0=>write_offset_data_out_2, A1
      =>write_base_data_out_2);
   ix7405 : inv01 port map ( Y=>nx7330, A=>nx7356);
   ix7406 : inv01 port map ( Y=>nx7331, A=>nx7360);
   ix7407 : nand02_2x port map ( Y=>nx7332, A0=>nx7356, A1=>nx7360);
   ix7408 : nor02_2x port map ( Y=>nx7333, A0=>nx7358, A1=>nx4293);
   ix7409 : aoi22 port map ( Y=>nx7334, A0=>nx7330, A1=>nx7331, B0=>nx7332, 
      B1=>nx7333);
   ix7410 : aoi22 port map ( Y=>nx7335, A0=>nx7329, A1=>nx7334, B0=>nx5777, 
      B1=>nx7329);
   reg_nx5847 : inv02 port map ( Y=>nx5847, A=>nx7335);
   ix7411 : inv01 port map ( Y=>nx7336, A=>nx7335);
   ix7412 : and02 port map ( Y=>nx7337, A0=>nx7356, A1=>nx7360);
   reg_nx2850 : oai32 port map ( Y=>nx2850, A0=>nx7337, A1=>nx7358, A2=>
      nx4293, B0=>nx7356, B1=>nx7360);
   reg_nx5667 : or02 port map ( Y=>nx5667, A0=>nx7358, A1=>nx4293);
   reg_nx5725 : oai22 port map ( Y=>nx5725, A0=>nx7330, A1=>nx7331, B0=>
      nx7356, B1=>nx7360);
   reg_nx6775 : inv01 port map ( Y=>nx6775, A=>nx7358);
   reg_nx7047 : inv01 port map ( Y=>nx7047, A=>nx7367);
   ix7413 : nor04_2x port map ( Y=>nx7338, A0=>class_cntr_counter_out_0, A1
      =>class_cntr_counter_out_2, A2=>nx5202, A3=>nx5218);
   ix7414 : inv01 port map ( Y=>nx7339, A=>mem_data_in(6));
   ix7415 : inv01 port map ( Y=>nx7340, A=>current_state_27);
   reg_argmax_data_out_6 : nor03_2x port map ( Y=>argmax_data_out(6), A0=>
      nx7338, A1=>nx7339, A2=>nx7340);
   reg_argmax_ready_XX0_XREP5 : nor02_2x port map ( Y=>
      argmax_ready_XX0_XREP5, A0=>nx7340, A1=>nx7338);
   ix7416 : inv02 port map ( Y=>nx7341, A=>nx6426);
   ix7417 : inv01 port map ( Y=>nx7342, A=>nx7301);
   ix7418 : inv01 port map ( Y=>nx7343, A=>nx7299);
   ix7419 : nand03_2x port map ( Y=>nx7344, A0=>nx7341, A1=>nx7342, A2=>
      nx7343);
   ix7420 : inv01 port map ( Y=>nx7345, A=>nx7366);
   ix7421 : inv02 port map ( Y=>nx7346, A=>nx4320);
   ix7422 : nor02_2x port map ( Y=>nx7347, A0=>nx7302, A1=>nx7303);
   ix7423 : nor02ii port map ( Y=>nx7348, A0=>nx6426, A1=>nx7300);
   ix7424 : aoi222 port map ( Y=>nx7349, A0=>nx7345, A1=>nx7346, B0=>nx7342, 
      B1=>nx7347, C0=>nx7342, C1=>nx7348);
   ix7425 : oai32 port map ( Y=>nx7350, A0=>nx7305, A1=>nx7445, A2=>nx7344, 
      B0=>nx7349, B1=>nx7305);
   ix7426 : inv02 port map ( Y=>nx7351, A=>nx7300);
   ix7427 : oai22 port map ( Y=>nx7352, A0=>nx7351, A1=>nx6426, B0=>nx7302, 
      B1=>nx7303);
   ix7428 : nor04_2x port map ( Y=>nx7353, A0=>nx7445, A1=>nx6426, A2=>
      nx7301, A3=>nx7299);
   reg_NOT_nx4700 : aoi221 port map ( Y=>NOT_nx4700, A0=>nx7345, A1=>nx7346, 
      B0=>nx7352, B1=>nx7342, C0=>nx7353);
   ix7429 : nor02_2x port map ( Y=>nx7354, A0=>nx7445, A1=>nx7299);
   ix7430 : buf16 port map ( Y=>nx7355, A=>nx4284);
   ix7431 : buf16 port map ( Y=>nx7356, A=>nx4284);
   ix7432 : buf16 port map ( Y=>nx7357, A=>nx5611);
   ix7433 : buf16 port map ( Y=>nx7358, A=>nx5611);
   ix7434 : buf16 port map ( Y=>nx7359, A=>nx5685);
   ix7435 : buf16 port map ( Y=>nx7360, A=>nx5685);
   ix7436 : buf16 port map ( Y=>nx7361, A=>nx5747);
   ix7437 : buf16 port map ( Y=>nx7362, A=>nx5747);
   ix7438 : buf16 port map ( Y=>nx7363, A=>nx6363);
   ix7439 : buf16 port map ( Y=>nx7364, A=>nx6363);
   ix7440 : buf16 port map ( Y=>nx7365, A=>nx6484);
   ix7441 : buf16 port map ( Y=>nx7366, A=>nx6484);
   ix7442 : buf16 port map ( Y=>argmax_ready_EXMPLR, A=>
      argmax_ready_XX0_XREP5);
   ix7443 : buf16 port map ( Y=>nx7367, A=>argmax_ready_XX0_XREP5);
   ix7444 : buf02 port map ( Y=>nx7445, A=>nx6367);
end Mixed_unfold_2045 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity CacheMuxer is
   port (
      d_arr_mux_0_31 : IN std_logic ;
      d_arr_mux_0_30 : IN std_logic ;
      d_arr_mux_0_29 : IN std_logic ;
      d_arr_mux_0_28 : IN std_logic ;
      d_arr_mux_0_27 : IN std_logic ;
      d_arr_mux_0_26 : IN std_logic ;
      d_arr_mux_0_25 : IN std_logic ;
      d_arr_mux_0_24 : IN std_logic ;
      d_arr_mux_0_23 : IN std_logic ;
      d_arr_mux_0_22 : IN std_logic ;
      d_arr_mux_0_21 : IN std_logic ;
      d_arr_mux_0_20 : IN std_logic ;
      d_arr_mux_0_19 : IN std_logic ;
      d_arr_mux_0_18 : IN std_logic ;
      d_arr_mux_0_17 : IN std_logic ;
      d_arr_mux_0_16 : IN std_logic ;
      d_arr_mux_0_15 : IN std_logic ;
      d_arr_mux_0_14 : IN std_logic ;
      d_arr_mux_0_13 : IN std_logic ;
      d_arr_mux_0_12 : IN std_logic ;
      d_arr_mux_0_11 : IN std_logic ;
      d_arr_mux_0_10 : IN std_logic ;
      d_arr_mux_0_9 : IN std_logic ;
      d_arr_mux_0_8 : IN std_logic ;
      d_arr_mux_0_7 : IN std_logic ;
      d_arr_mux_0_6 : IN std_logic ;
      d_arr_mux_0_5 : IN std_logic ;
      d_arr_mux_0_4 : IN std_logic ;
      d_arr_mux_0_3 : IN std_logic ;
      d_arr_mux_0_2 : IN std_logic ;
      d_arr_mux_0_1 : IN std_logic ;
      d_arr_mux_0_0 : IN std_logic ;
      d_arr_mux_1_31 : IN std_logic ;
      d_arr_mux_1_30 : IN std_logic ;
      d_arr_mux_1_29 : IN std_logic ;
      d_arr_mux_1_28 : IN std_logic ;
      d_arr_mux_1_27 : IN std_logic ;
      d_arr_mux_1_26 : IN std_logic ;
      d_arr_mux_1_25 : IN std_logic ;
      d_arr_mux_1_24 : IN std_logic ;
      d_arr_mux_1_23 : IN std_logic ;
      d_arr_mux_1_22 : IN std_logic ;
      d_arr_mux_1_21 : IN std_logic ;
      d_arr_mux_1_20 : IN std_logic ;
      d_arr_mux_1_19 : IN std_logic ;
      d_arr_mux_1_18 : IN std_logic ;
      d_arr_mux_1_17 : IN std_logic ;
      d_arr_mux_1_16 : IN std_logic ;
      d_arr_mux_1_15 : IN std_logic ;
      d_arr_mux_1_14 : IN std_logic ;
      d_arr_mux_1_13 : IN std_logic ;
      d_arr_mux_1_12 : IN std_logic ;
      d_arr_mux_1_11 : IN std_logic ;
      d_arr_mux_1_10 : IN std_logic ;
      d_arr_mux_1_9 : IN std_logic ;
      d_arr_mux_1_8 : IN std_logic ;
      d_arr_mux_1_7 : IN std_logic ;
      d_arr_mux_1_6 : IN std_logic ;
      d_arr_mux_1_5 : IN std_logic ;
      d_arr_mux_1_4 : IN std_logic ;
      d_arr_mux_1_3 : IN std_logic ;
      d_arr_mux_1_2 : IN std_logic ;
      d_arr_mux_1_1 : IN std_logic ;
      d_arr_mux_1_0 : IN std_logic ;
      d_arr_mux_2_31 : IN std_logic ;
      d_arr_mux_2_30 : IN std_logic ;
      d_arr_mux_2_29 : IN std_logic ;
      d_arr_mux_2_28 : IN std_logic ;
      d_arr_mux_2_27 : IN std_logic ;
      d_arr_mux_2_26 : IN std_logic ;
      d_arr_mux_2_25 : IN std_logic ;
      d_arr_mux_2_24 : IN std_logic ;
      d_arr_mux_2_23 : IN std_logic ;
      d_arr_mux_2_22 : IN std_logic ;
      d_arr_mux_2_21 : IN std_logic ;
      d_arr_mux_2_20 : IN std_logic ;
      d_arr_mux_2_19 : IN std_logic ;
      d_arr_mux_2_18 : IN std_logic ;
      d_arr_mux_2_17 : IN std_logic ;
      d_arr_mux_2_16 : IN std_logic ;
      d_arr_mux_2_15 : IN std_logic ;
      d_arr_mux_2_14 : IN std_logic ;
      d_arr_mux_2_13 : IN std_logic ;
      d_arr_mux_2_12 : IN std_logic ;
      d_arr_mux_2_11 : IN std_logic ;
      d_arr_mux_2_10 : IN std_logic ;
      d_arr_mux_2_9 : IN std_logic ;
      d_arr_mux_2_8 : IN std_logic ;
      d_arr_mux_2_7 : IN std_logic ;
      d_arr_mux_2_6 : IN std_logic ;
      d_arr_mux_2_5 : IN std_logic ;
      d_arr_mux_2_4 : IN std_logic ;
      d_arr_mux_2_3 : IN std_logic ;
      d_arr_mux_2_2 : IN std_logic ;
      d_arr_mux_2_1 : IN std_logic ;
      d_arr_mux_2_0 : IN std_logic ;
      d_arr_mux_3_31 : IN std_logic ;
      d_arr_mux_3_30 : IN std_logic ;
      d_arr_mux_3_29 : IN std_logic ;
      d_arr_mux_3_28 : IN std_logic ;
      d_arr_mux_3_27 : IN std_logic ;
      d_arr_mux_3_26 : IN std_logic ;
      d_arr_mux_3_25 : IN std_logic ;
      d_arr_mux_3_24 : IN std_logic ;
      d_arr_mux_3_23 : IN std_logic ;
      d_arr_mux_3_22 : IN std_logic ;
      d_arr_mux_3_21 : IN std_logic ;
      d_arr_mux_3_20 : IN std_logic ;
      d_arr_mux_3_19 : IN std_logic ;
      d_arr_mux_3_18 : IN std_logic ;
      d_arr_mux_3_17 : IN std_logic ;
      d_arr_mux_3_16 : IN std_logic ;
      d_arr_mux_3_15 : IN std_logic ;
      d_arr_mux_3_14 : IN std_logic ;
      d_arr_mux_3_13 : IN std_logic ;
      d_arr_mux_3_12 : IN std_logic ;
      d_arr_mux_3_11 : IN std_logic ;
      d_arr_mux_3_10 : IN std_logic ;
      d_arr_mux_3_9 : IN std_logic ;
      d_arr_mux_3_8 : IN std_logic ;
      d_arr_mux_3_7 : IN std_logic ;
      d_arr_mux_3_6 : IN std_logic ;
      d_arr_mux_3_5 : IN std_logic ;
      d_arr_mux_3_4 : IN std_logic ;
      d_arr_mux_3_3 : IN std_logic ;
      d_arr_mux_3_2 : IN std_logic ;
      d_arr_mux_3_1 : IN std_logic ;
      d_arr_mux_3_0 : IN std_logic ;
      d_arr_mux_4_31 : IN std_logic ;
      d_arr_mux_4_30 : IN std_logic ;
      d_arr_mux_4_29 : IN std_logic ;
      d_arr_mux_4_28 : IN std_logic ;
      d_arr_mux_4_27 : IN std_logic ;
      d_arr_mux_4_26 : IN std_logic ;
      d_arr_mux_4_25 : IN std_logic ;
      d_arr_mux_4_24 : IN std_logic ;
      d_arr_mux_4_23 : IN std_logic ;
      d_arr_mux_4_22 : IN std_logic ;
      d_arr_mux_4_21 : IN std_logic ;
      d_arr_mux_4_20 : IN std_logic ;
      d_arr_mux_4_19 : IN std_logic ;
      d_arr_mux_4_18 : IN std_logic ;
      d_arr_mux_4_17 : IN std_logic ;
      d_arr_mux_4_16 : IN std_logic ;
      d_arr_mux_4_15 : IN std_logic ;
      d_arr_mux_4_14 : IN std_logic ;
      d_arr_mux_4_13 : IN std_logic ;
      d_arr_mux_4_12 : IN std_logic ;
      d_arr_mux_4_11 : IN std_logic ;
      d_arr_mux_4_10 : IN std_logic ;
      d_arr_mux_4_9 : IN std_logic ;
      d_arr_mux_4_8 : IN std_logic ;
      d_arr_mux_4_7 : IN std_logic ;
      d_arr_mux_4_6 : IN std_logic ;
      d_arr_mux_4_5 : IN std_logic ;
      d_arr_mux_4_4 : IN std_logic ;
      d_arr_mux_4_3 : IN std_logic ;
      d_arr_mux_4_2 : IN std_logic ;
      d_arr_mux_4_1 : IN std_logic ;
      d_arr_mux_4_0 : IN std_logic ;
      d_arr_mux_5_31 : IN std_logic ;
      d_arr_mux_5_30 : IN std_logic ;
      d_arr_mux_5_29 : IN std_logic ;
      d_arr_mux_5_28 : IN std_logic ;
      d_arr_mux_5_27 : IN std_logic ;
      d_arr_mux_5_26 : IN std_logic ;
      d_arr_mux_5_25 : IN std_logic ;
      d_arr_mux_5_24 : IN std_logic ;
      d_arr_mux_5_23 : IN std_logic ;
      d_arr_mux_5_22 : IN std_logic ;
      d_arr_mux_5_21 : IN std_logic ;
      d_arr_mux_5_20 : IN std_logic ;
      d_arr_mux_5_19 : IN std_logic ;
      d_arr_mux_5_18 : IN std_logic ;
      d_arr_mux_5_17 : IN std_logic ;
      d_arr_mux_5_16 : IN std_logic ;
      d_arr_mux_5_15 : IN std_logic ;
      d_arr_mux_5_14 : IN std_logic ;
      d_arr_mux_5_13 : IN std_logic ;
      d_arr_mux_5_12 : IN std_logic ;
      d_arr_mux_5_11 : IN std_logic ;
      d_arr_mux_5_10 : IN std_logic ;
      d_arr_mux_5_9 : IN std_logic ;
      d_arr_mux_5_8 : IN std_logic ;
      d_arr_mux_5_7 : IN std_logic ;
      d_arr_mux_5_6 : IN std_logic ;
      d_arr_mux_5_5 : IN std_logic ;
      d_arr_mux_5_4 : IN std_logic ;
      d_arr_mux_5_3 : IN std_logic ;
      d_arr_mux_5_2 : IN std_logic ;
      d_arr_mux_5_1 : IN std_logic ;
      d_arr_mux_5_0 : IN std_logic ;
      d_arr_mux_6_31 : IN std_logic ;
      d_arr_mux_6_30 : IN std_logic ;
      d_arr_mux_6_29 : IN std_logic ;
      d_arr_mux_6_28 : IN std_logic ;
      d_arr_mux_6_27 : IN std_logic ;
      d_arr_mux_6_26 : IN std_logic ;
      d_arr_mux_6_25 : IN std_logic ;
      d_arr_mux_6_24 : IN std_logic ;
      d_arr_mux_6_23 : IN std_logic ;
      d_arr_mux_6_22 : IN std_logic ;
      d_arr_mux_6_21 : IN std_logic ;
      d_arr_mux_6_20 : IN std_logic ;
      d_arr_mux_6_19 : IN std_logic ;
      d_arr_mux_6_18 : IN std_logic ;
      d_arr_mux_6_17 : IN std_logic ;
      d_arr_mux_6_16 : IN std_logic ;
      d_arr_mux_6_15 : IN std_logic ;
      d_arr_mux_6_14 : IN std_logic ;
      d_arr_mux_6_13 : IN std_logic ;
      d_arr_mux_6_12 : IN std_logic ;
      d_arr_mux_6_11 : IN std_logic ;
      d_arr_mux_6_10 : IN std_logic ;
      d_arr_mux_6_9 : IN std_logic ;
      d_arr_mux_6_8 : IN std_logic ;
      d_arr_mux_6_7 : IN std_logic ;
      d_arr_mux_6_6 : IN std_logic ;
      d_arr_mux_6_5 : IN std_logic ;
      d_arr_mux_6_4 : IN std_logic ;
      d_arr_mux_6_3 : IN std_logic ;
      d_arr_mux_6_2 : IN std_logic ;
      d_arr_mux_6_1 : IN std_logic ;
      d_arr_mux_6_0 : IN std_logic ;
      d_arr_mux_7_31 : IN std_logic ;
      d_arr_mux_7_30 : IN std_logic ;
      d_arr_mux_7_29 : IN std_logic ;
      d_arr_mux_7_28 : IN std_logic ;
      d_arr_mux_7_27 : IN std_logic ;
      d_arr_mux_7_26 : IN std_logic ;
      d_arr_mux_7_25 : IN std_logic ;
      d_arr_mux_7_24 : IN std_logic ;
      d_arr_mux_7_23 : IN std_logic ;
      d_arr_mux_7_22 : IN std_logic ;
      d_arr_mux_7_21 : IN std_logic ;
      d_arr_mux_7_20 : IN std_logic ;
      d_arr_mux_7_19 : IN std_logic ;
      d_arr_mux_7_18 : IN std_logic ;
      d_arr_mux_7_17 : IN std_logic ;
      d_arr_mux_7_16 : IN std_logic ;
      d_arr_mux_7_15 : IN std_logic ;
      d_arr_mux_7_14 : IN std_logic ;
      d_arr_mux_7_13 : IN std_logic ;
      d_arr_mux_7_12 : IN std_logic ;
      d_arr_mux_7_11 : IN std_logic ;
      d_arr_mux_7_10 : IN std_logic ;
      d_arr_mux_7_9 : IN std_logic ;
      d_arr_mux_7_8 : IN std_logic ;
      d_arr_mux_7_7 : IN std_logic ;
      d_arr_mux_7_6 : IN std_logic ;
      d_arr_mux_7_5 : IN std_logic ;
      d_arr_mux_7_4 : IN std_logic ;
      d_arr_mux_7_3 : IN std_logic ;
      d_arr_mux_7_2 : IN std_logic ;
      d_arr_mux_7_1 : IN std_logic ;
      d_arr_mux_7_0 : IN std_logic ;
      d_arr_mux_8_31 : IN std_logic ;
      d_arr_mux_8_30 : IN std_logic ;
      d_arr_mux_8_29 : IN std_logic ;
      d_arr_mux_8_28 : IN std_logic ;
      d_arr_mux_8_27 : IN std_logic ;
      d_arr_mux_8_26 : IN std_logic ;
      d_arr_mux_8_25 : IN std_logic ;
      d_arr_mux_8_24 : IN std_logic ;
      d_arr_mux_8_23 : IN std_logic ;
      d_arr_mux_8_22 : IN std_logic ;
      d_arr_mux_8_21 : IN std_logic ;
      d_arr_mux_8_20 : IN std_logic ;
      d_arr_mux_8_19 : IN std_logic ;
      d_arr_mux_8_18 : IN std_logic ;
      d_arr_mux_8_17 : IN std_logic ;
      d_arr_mux_8_16 : IN std_logic ;
      d_arr_mux_8_15 : IN std_logic ;
      d_arr_mux_8_14 : IN std_logic ;
      d_arr_mux_8_13 : IN std_logic ;
      d_arr_mux_8_12 : IN std_logic ;
      d_arr_mux_8_11 : IN std_logic ;
      d_arr_mux_8_10 : IN std_logic ;
      d_arr_mux_8_9 : IN std_logic ;
      d_arr_mux_8_8 : IN std_logic ;
      d_arr_mux_8_7 : IN std_logic ;
      d_arr_mux_8_6 : IN std_logic ;
      d_arr_mux_8_5 : IN std_logic ;
      d_arr_mux_8_4 : IN std_logic ;
      d_arr_mux_8_3 : IN std_logic ;
      d_arr_mux_8_2 : IN std_logic ;
      d_arr_mux_8_1 : IN std_logic ;
      d_arr_mux_8_0 : IN std_logic ;
      d_arr_mux_9_31 : IN std_logic ;
      d_arr_mux_9_30 : IN std_logic ;
      d_arr_mux_9_29 : IN std_logic ;
      d_arr_mux_9_28 : IN std_logic ;
      d_arr_mux_9_27 : IN std_logic ;
      d_arr_mux_9_26 : IN std_logic ;
      d_arr_mux_9_25 : IN std_logic ;
      d_arr_mux_9_24 : IN std_logic ;
      d_arr_mux_9_23 : IN std_logic ;
      d_arr_mux_9_22 : IN std_logic ;
      d_arr_mux_9_21 : IN std_logic ;
      d_arr_mux_9_20 : IN std_logic ;
      d_arr_mux_9_19 : IN std_logic ;
      d_arr_mux_9_18 : IN std_logic ;
      d_arr_mux_9_17 : IN std_logic ;
      d_arr_mux_9_16 : IN std_logic ;
      d_arr_mux_9_15 : IN std_logic ;
      d_arr_mux_9_14 : IN std_logic ;
      d_arr_mux_9_13 : IN std_logic ;
      d_arr_mux_9_12 : IN std_logic ;
      d_arr_mux_9_11 : IN std_logic ;
      d_arr_mux_9_10 : IN std_logic ;
      d_arr_mux_9_9 : IN std_logic ;
      d_arr_mux_9_8 : IN std_logic ;
      d_arr_mux_9_7 : IN std_logic ;
      d_arr_mux_9_6 : IN std_logic ;
      d_arr_mux_9_5 : IN std_logic ;
      d_arr_mux_9_4 : IN std_logic ;
      d_arr_mux_9_3 : IN std_logic ;
      d_arr_mux_9_2 : IN std_logic ;
      d_arr_mux_9_1 : IN std_logic ;
      d_arr_mux_9_0 : IN std_logic ;
      d_arr_mux_10_31 : IN std_logic ;
      d_arr_mux_10_30 : IN std_logic ;
      d_arr_mux_10_29 : IN std_logic ;
      d_arr_mux_10_28 : IN std_logic ;
      d_arr_mux_10_27 : IN std_logic ;
      d_arr_mux_10_26 : IN std_logic ;
      d_arr_mux_10_25 : IN std_logic ;
      d_arr_mux_10_24 : IN std_logic ;
      d_arr_mux_10_23 : IN std_logic ;
      d_arr_mux_10_22 : IN std_logic ;
      d_arr_mux_10_21 : IN std_logic ;
      d_arr_mux_10_20 : IN std_logic ;
      d_arr_mux_10_19 : IN std_logic ;
      d_arr_mux_10_18 : IN std_logic ;
      d_arr_mux_10_17 : IN std_logic ;
      d_arr_mux_10_16 : IN std_logic ;
      d_arr_mux_10_15 : IN std_logic ;
      d_arr_mux_10_14 : IN std_logic ;
      d_arr_mux_10_13 : IN std_logic ;
      d_arr_mux_10_12 : IN std_logic ;
      d_arr_mux_10_11 : IN std_logic ;
      d_arr_mux_10_10 : IN std_logic ;
      d_arr_mux_10_9 : IN std_logic ;
      d_arr_mux_10_8 : IN std_logic ;
      d_arr_mux_10_7 : IN std_logic ;
      d_arr_mux_10_6 : IN std_logic ;
      d_arr_mux_10_5 : IN std_logic ;
      d_arr_mux_10_4 : IN std_logic ;
      d_arr_mux_10_3 : IN std_logic ;
      d_arr_mux_10_2 : IN std_logic ;
      d_arr_mux_10_1 : IN std_logic ;
      d_arr_mux_10_0 : IN std_logic ;
      d_arr_mux_11_31 : IN std_logic ;
      d_arr_mux_11_30 : IN std_logic ;
      d_arr_mux_11_29 : IN std_logic ;
      d_arr_mux_11_28 : IN std_logic ;
      d_arr_mux_11_27 : IN std_logic ;
      d_arr_mux_11_26 : IN std_logic ;
      d_arr_mux_11_25 : IN std_logic ;
      d_arr_mux_11_24 : IN std_logic ;
      d_arr_mux_11_23 : IN std_logic ;
      d_arr_mux_11_22 : IN std_logic ;
      d_arr_mux_11_21 : IN std_logic ;
      d_arr_mux_11_20 : IN std_logic ;
      d_arr_mux_11_19 : IN std_logic ;
      d_arr_mux_11_18 : IN std_logic ;
      d_arr_mux_11_17 : IN std_logic ;
      d_arr_mux_11_16 : IN std_logic ;
      d_arr_mux_11_15 : IN std_logic ;
      d_arr_mux_11_14 : IN std_logic ;
      d_arr_mux_11_13 : IN std_logic ;
      d_arr_mux_11_12 : IN std_logic ;
      d_arr_mux_11_11 : IN std_logic ;
      d_arr_mux_11_10 : IN std_logic ;
      d_arr_mux_11_9 : IN std_logic ;
      d_arr_mux_11_8 : IN std_logic ;
      d_arr_mux_11_7 : IN std_logic ;
      d_arr_mux_11_6 : IN std_logic ;
      d_arr_mux_11_5 : IN std_logic ;
      d_arr_mux_11_4 : IN std_logic ;
      d_arr_mux_11_3 : IN std_logic ;
      d_arr_mux_11_2 : IN std_logic ;
      d_arr_mux_11_1 : IN std_logic ;
      d_arr_mux_11_0 : IN std_logic ;
      d_arr_mux_12_31 : IN std_logic ;
      d_arr_mux_12_30 : IN std_logic ;
      d_arr_mux_12_29 : IN std_logic ;
      d_arr_mux_12_28 : IN std_logic ;
      d_arr_mux_12_27 : IN std_logic ;
      d_arr_mux_12_26 : IN std_logic ;
      d_arr_mux_12_25 : IN std_logic ;
      d_arr_mux_12_24 : IN std_logic ;
      d_arr_mux_12_23 : IN std_logic ;
      d_arr_mux_12_22 : IN std_logic ;
      d_arr_mux_12_21 : IN std_logic ;
      d_arr_mux_12_20 : IN std_logic ;
      d_arr_mux_12_19 : IN std_logic ;
      d_arr_mux_12_18 : IN std_logic ;
      d_arr_mux_12_17 : IN std_logic ;
      d_arr_mux_12_16 : IN std_logic ;
      d_arr_mux_12_15 : IN std_logic ;
      d_arr_mux_12_14 : IN std_logic ;
      d_arr_mux_12_13 : IN std_logic ;
      d_arr_mux_12_12 : IN std_logic ;
      d_arr_mux_12_11 : IN std_logic ;
      d_arr_mux_12_10 : IN std_logic ;
      d_arr_mux_12_9 : IN std_logic ;
      d_arr_mux_12_8 : IN std_logic ;
      d_arr_mux_12_7 : IN std_logic ;
      d_arr_mux_12_6 : IN std_logic ;
      d_arr_mux_12_5 : IN std_logic ;
      d_arr_mux_12_4 : IN std_logic ;
      d_arr_mux_12_3 : IN std_logic ;
      d_arr_mux_12_2 : IN std_logic ;
      d_arr_mux_12_1 : IN std_logic ;
      d_arr_mux_12_0 : IN std_logic ;
      d_arr_mux_13_31 : IN std_logic ;
      d_arr_mux_13_30 : IN std_logic ;
      d_arr_mux_13_29 : IN std_logic ;
      d_arr_mux_13_28 : IN std_logic ;
      d_arr_mux_13_27 : IN std_logic ;
      d_arr_mux_13_26 : IN std_logic ;
      d_arr_mux_13_25 : IN std_logic ;
      d_arr_mux_13_24 : IN std_logic ;
      d_arr_mux_13_23 : IN std_logic ;
      d_arr_mux_13_22 : IN std_logic ;
      d_arr_mux_13_21 : IN std_logic ;
      d_arr_mux_13_20 : IN std_logic ;
      d_arr_mux_13_19 : IN std_logic ;
      d_arr_mux_13_18 : IN std_logic ;
      d_arr_mux_13_17 : IN std_logic ;
      d_arr_mux_13_16 : IN std_logic ;
      d_arr_mux_13_15 : IN std_logic ;
      d_arr_mux_13_14 : IN std_logic ;
      d_arr_mux_13_13 : IN std_logic ;
      d_arr_mux_13_12 : IN std_logic ;
      d_arr_mux_13_11 : IN std_logic ;
      d_arr_mux_13_10 : IN std_logic ;
      d_arr_mux_13_9 : IN std_logic ;
      d_arr_mux_13_8 : IN std_logic ;
      d_arr_mux_13_7 : IN std_logic ;
      d_arr_mux_13_6 : IN std_logic ;
      d_arr_mux_13_5 : IN std_logic ;
      d_arr_mux_13_4 : IN std_logic ;
      d_arr_mux_13_3 : IN std_logic ;
      d_arr_mux_13_2 : IN std_logic ;
      d_arr_mux_13_1 : IN std_logic ;
      d_arr_mux_13_0 : IN std_logic ;
      d_arr_mux_14_31 : IN std_logic ;
      d_arr_mux_14_30 : IN std_logic ;
      d_arr_mux_14_29 : IN std_logic ;
      d_arr_mux_14_28 : IN std_logic ;
      d_arr_mux_14_27 : IN std_logic ;
      d_arr_mux_14_26 : IN std_logic ;
      d_arr_mux_14_25 : IN std_logic ;
      d_arr_mux_14_24 : IN std_logic ;
      d_arr_mux_14_23 : IN std_logic ;
      d_arr_mux_14_22 : IN std_logic ;
      d_arr_mux_14_21 : IN std_logic ;
      d_arr_mux_14_20 : IN std_logic ;
      d_arr_mux_14_19 : IN std_logic ;
      d_arr_mux_14_18 : IN std_logic ;
      d_arr_mux_14_17 : IN std_logic ;
      d_arr_mux_14_16 : IN std_logic ;
      d_arr_mux_14_15 : IN std_logic ;
      d_arr_mux_14_14 : IN std_logic ;
      d_arr_mux_14_13 : IN std_logic ;
      d_arr_mux_14_12 : IN std_logic ;
      d_arr_mux_14_11 : IN std_logic ;
      d_arr_mux_14_10 : IN std_logic ;
      d_arr_mux_14_9 : IN std_logic ;
      d_arr_mux_14_8 : IN std_logic ;
      d_arr_mux_14_7 : IN std_logic ;
      d_arr_mux_14_6 : IN std_logic ;
      d_arr_mux_14_5 : IN std_logic ;
      d_arr_mux_14_4 : IN std_logic ;
      d_arr_mux_14_3 : IN std_logic ;
      d_arr_mux_14_2 : IN std_logic ;
      d_arr_mux_14_1 : IN std_logic ;
      d_arr_mux_14_0 : IN std_logic ;
      d_arr_mux_15_31 : IN std_logic ;
      d_arr_mux_15_30 : IN std_logic ;
      d_arr_mux_15_29 : IN std_logic ;
      d_arr_mux_15_28 : IN std_logic ;
      d_arr_mux_15_27 : IN std_logic ;
      d_arr_mux_15_26 : IN std_logic ;
      d_arr_mux_15_25 : IN std_logic ;
      d_arr_mux_15_24 : IN std_logic ;
      d_arr_mux_15_23 : IN std_logic ;
      d_arr_mux_15_22 : IN std_logic ;
      d_arr_mux_15_21 : IN std_logic ;
      d_arr_mux_15_20 : IN std_logic ;
      d_arr_mux_15_19 : IN std_logic ;
      d_arr_mux_15_18 : IN std_logic ;
      d_arr_mux_15_17 : IN std_logic ;
      d_arr_mux_15_16 : IN std_logic ;
      d_arr_mux_15_15 : IN std_logic ;
      d_arr_mux_15_14 : IN std_logic ;
      d_arr_mux_15_13 : IN std_logic ;
      d_arr_mux_15_12 : IN std_logic ;
      d_arr_mux_15_11 : IN std_logic ;
      d_arr_mux_15_10 : IN std_logic ;
      d_arr_mux_15_9 : IN std_logic ;
      d_arr_mux_15_8 : IN std_logic ;
      d_arr_mux_15_7 : IN std_logic ;
      d_arr_mux_15_6 : IN std_logic ;
      d_arr_mux_15_5 : IN std_logic ;
      d_arr_mux_15_4 : IN std_logic ;
      d_arr_mux_15_3 : IN std_logic ;
      d_arr_mux_15_2 : IN std_logic ;
      d_arr_mux_15_1 : IN std_logic ;
      d_arr_mux_15_0 : IN std_logic ;
      d_arr_mux_16_31 : IN std_logic ;
      d_arr_mux_16_30 : IN std_logic ;
      d_arr_mux_16_29 : IN std_logic ;
      d_arr_mux_16_28 : IN std_logic ;
      d_arr_mux_16_27 : IN std_logic ;
      d_arr_mux_16_26 : IN std_logic ;
      d_arr_mux_16_25 : IN std_logic ;
      d_arr_mux_16_24 : IN std_logic ;
      d_arr_mux_16_23 : IN std_logic ;
      d_arr_mux_16_22 : IN std_logic ;
      d_arr_mux_16_21 : IN std_logic ;
      d_arr_mux_16_20 : IN std_logic ;
      d_arr_mux_16_19 : IN std_logic ;
      d_arr_mux_16_18 : IN std_logic ;
      d_arr_mux_16_17 : IN std_logic ;
      d_arr_mux_16_16 : IN std_logic ;
      d_arr_mux_16_15 : IN std_logic ;
      d_arr_mux_16_14 : IN std_logic ;
      d_arr_mux_16_13 : IN std_logic ;
      d_arr_mux_16_12 : IN std_logic ;
      d_arr_mux_16_11 : IN std_logic ;
      d_arr_mux_16_10 : IN std_logic ;
      d_arr_mux_16_9 : IN std_logic ;
      d_arr_mux_16_8 : IN std_logic ;
      d_arr_mux_16_7 : IN std_logic ;
      d_arr_mux_16_6 : IN std_logic ;
      d_arr_mux_16_5 : IN std_logic ;
      d_arr_mux_16_4 : IN std_logic ;
      d_arr_mux_16_3 : IN std_logic ;
      d_arr_mux_16_2 : IN std_logic ;
      d_arr_mux_16_1 : IN std_logic ;
      d_arr_mux_16_0 : IN std_logic ;
      d_arr_mux_17_31 : IN std_logic ;
      d_arr_mux_17_30 : IN std_logic ;
      d_arr_mux_17_29 : IN std_logic ;
      d_arr_mux_17_28 : IN std_logic ;
      d_arr_mux_17_27 : IN std_logic ;
      d_arr_mux_17_26 : IN std_logic ;
      d_arr_mux_17_25 : IN std_logic ;
      d_arr_mux_17_24 : IN std_logic ;
      d_arr_mux_17_23 : IN std_logic ;
      d_arr_mux_17_22 : IN std_logic ;
      d_arr_mux_17_21 : IN std_logic ;
      d_arr_mux_17_20 : IN std_logic ;
      d_arr_mux_17_19 : IN std_logic ;
      d_arr_mux_17_18 : IN std_logic ;
      d_arr_mux_17_17 : IN std_logic ;
      d_arr_mux_17_16 : IN std_logic ;
      d_arr_mux_17_15 : IN std_logic ;
      d_arr_mux_17_14 : IN std_logic ;
      d_arr_mux_17_13 : IN std_logic ;
      d_arr_mux_17_12 : IN std_logic ;
      d_arr_mux_17_11 : IN std_logic ;
      d_arr_mux_17_10 : IN std_logic ;
      d_arr_mux_17_9 : IN std_logic ;
      d_arr_mux_17_8 : IN std_logic ;
      d_arr_mux_17_7 : IN std_logic ;
      d_arr_mux_17_6 : IN std_logic ;
      d_arr_mux_17_5 : IN std_logic ;
      d_arr_mux_17_4 : IN std_logic ;
      d_arr_mux_17_3 : IN std_logic ;
      d_arr_mux_17_2 : IN std_logic ;
      d_arr_mux_17_1 : IN std_logic ;
      d_arr_mux_17_0 : IN std_logic ;
      d_arr_mux_18_31 : IN std_logic ;
      d_arr_mux_18_30 : IN std_logic ;
      d_arr_mux_18_29 : IN std_logic ;
      d_arr_mux_18_28 : IN std_logic ;
      d_arr_mux_18_27 : IN std_logic ;
      d_arr_mux_18_26 : IN std_logic ;
      d_arr_mux_18_25 : IN std_logic ;
      d_arr_mux_18_24 : IN std_logic ;
      d_arr_mux_18_23 : IN std_logic ;
      d_arr_mux_18_22 : IN std_logic ;
      d_arr_mux_18_21 : IN std_logic ;
      d_arr_mux_18_20 : IN std_logic ;
      d_arr_mux_18_19 : IN std_logic ;
      d_arr_mux_18_18 : IN std_logic ;
      d_arr_mux_18_17 : IN std_logic ;
      d_arr_mux_18_16 : IN std_logic ;
      d_arr_mux_18_15 : IN std_logic ;
      d_arr_mux_18_14 : IN std_logic ;
      d_arr_mux_18_13 : IN std_logic ;
      d_arr_mux_18_12 : IN std_logic ;
      d_arr_mux_18_11 : IN std_logic ;
      d_arr_mux_18_10 : IN std_logic ;
      d_arr_mux_18_9 : IN std_logic ;
      d_arr_mux_18_8 : IN std_logic ;
      d_arr_mux_18_7 : IN std_logic ;
      d_arr_mux_18_6 : IN std_logic ;
      d_arr_mux_18_5 : IN std_logic ;
      d_arr_mux_18_4 : IN std_logic ;
      d_arr_mux_18_3 : IN std_logic ;
      d_arr_mux_18_2 : IN std_logic ;
      d_arr_mux_18_1 : IN std_logic ;
      d_arr_mux_18_0 : IN std_logic ;
      d_arr_mux_19_31 : IN std_logic ;
      d_arr_mux_19_30 : IN std_logic ;
      d_arr_mux_19_29 : IN std_logic ;
      d_arr_mux_19_28 : IN std_logic ;
      d_arr_mux_19_27 : IN std_logic ;
      d_arr_mux_19_26 : IN std_logic ;
      d_arr_mux_19_25 : IN std_logic ;
      d_arr_mux_19_24 : IN std_logic ;
      d_arr_mux_19_23 : IN std_logic ;
      d_arr_mux_19_22 : IN std_logic ;
      d_arr_mux_19_21 : IN std_logic ;
      d_arr_mux_19_20 : IN std_logic ;
      d_arr_mux_19_19 : IN std_logic ;
      d_arr_mux_19_18 : IN std_logic ;
      d_arr_mux_19_17 : IN std_logic ;
      d_arr_mux_19_16 : IN std_logic ;
      d_arr_mux_19_15 : IN std_logic ;
      d_arr_mux_19_14 : IN std_logic ;
      d_arr_mux_19_13 : IN std_logic ;
      d_arr_mux_19_12 : IN std_logic ;
      d_arr_mux_19_11 : IN std_logic ;
      d_arr_mux_19_10 : IN std_logic ;
      d_arr_mux_19_9 : IN std_logic ;
      d_arr_mux_19_8 : IN std_logic ;
      d_arr_mux_19_7 : IN std_logic ;
      d_arr_mux_19_6 : IN std_logic ;
      d_arr_mux_19_5 : IN std_logic ;
      d_arr_mux_19_4 : IN std_logic ;
      d_arr_mux_19_3 : IN std_logic ;
      d_arr_mux_19_2 : IN std_logic ;
      d_arr_mux_19_1 : IN std_logic ;
      d_arr_mux_19_0 : IN std_logic ;
      d_arr_mux_20_31 : IN std_logic ;
      d_arr_mux_20_30 : IN std_logic ;
      d_arr_mux_20_29 : IN std_logic ;
      d_arr_mux_20_28 : IN std_logic ;
      d_arr_mux_20_27 : IN std_logic ;
      d_arr_mux_20_26 : IN std_logic ;
      d_arr_mux_20_25 : IN std_logic ;
      d_arr_mux_20_24 : IN std_logic ;
      d_arr_mux_20_23 : IN std_logic ;
      d_arr_mux_20_22 : IN std_logic ;
      d_arr_mux_20_21 : IN std_logic ;
      d_arr_mux_20_20 : IN std_logic ;
      d_arr_mux_20_19 : IN std_logic ;
      d_arr_mux_20_18 : IN std_logic ;
      d_arr_mux_20_17 : IN std_logic ;
      d_arr_mux_20_16 : IN std_logic ;
      d_arr_mux_20_15 : IN std_logic ;
      d_arr_mux_20_14 : IN std_logic ;
      d_arr_mux_20_13 : IN std_logic ;
      d_arr_mux_20_12 : IN std_logic ;
      d_arr_mux_20_11 : IN std_logic ;
      d_arr_mux_20_10 : IN std_logic ;
      d_arr_mux_20_9 : IN std_logic ;
      d_arr_mux_20_8 : IN std_logic ;
      d_arr_mux_20_7 : IN std_logic ;
      d_arr_mux_20_6 : IN std_logic ;
      d_arr_mux_20_5 : IN std_logic ;
      d_arr_mux_20_4 : IN std_logic ;
      d_arr_mux_20_3 : IN std_logic ;
      d_arr_mux_20_2 : IN std_logic ;
      d_arr_mux_20_1 : IN std_logic ;
      d_arr_mux_20_0 : IN std_logic ;
      d_arr_mux_21_31 : IN std_logic ;
      d_arr_mux_21_30 : IN std_logic ;
      d_arr_mux_21_29 : IN std_logic ;
      d_arr_mux_21_28 : IN std_logic ;
      d_arr_mux_21_27 : IN std_logic ;
      d_arr_mux_21_26 : IN std_logic ;
      d_arr_mux_21_25 : IN std_logic ;
      d_arr_mux_21_24 : IN std_logic ;
      d_arr_mux_21_23 : IN std_logic ;
      d_arr_mux_21_22 : IN std_logic ;
      d_arr_mux_21_21 : IN std_logic ;
      d_arr_mux_21_20 : IN std_logic ;
      d_arr_mux_21_19 : IN std_logic ;
      d_arr_mux_21_18 : IN std_logic ;
      d_arr_mux_21_17 : IN std_logic ;
      d_arr_mux_21_16 : IN std_logic ;
      d_arr_mux_21_15 : IN std_logic ;
      d_arr_mux_21_14 : IN std_logic ;
      d_arr_mux_21_13 : IN std_logic ;
      d_arr_mux_21_12 : IN std_logic ;
      d_arr_mux_21_11 : IN std_logic ;
      d_arr_mux_21_10 : IN std_logic ;
      d_arr_mux_21_9 : IN std_logic ;
      d_arr_mux_21_8 : IN std_logic ;
      d_arr_mux_21_7 : IN std_logic ;
      d_arr_mux_21_6 : IN std_logic ;
      d_arr_mux_21_5 : IN std_logic ;
      d_arr_mux_21_4 : IN std_logic ;
      d_arr_mux_21_3 : IN std_logic ;
      d_arr_mux_21_2 : IN std_logic ;
      d_arr_mux_21_1 : IN std_logic ;
      d_arr_mux_21_0 : IN std_logic ;
      d_arr_mux_22_31 : IN std_logic ;
      d_arr_mux_22_30 : IN std_logic ;
      d_arr_mux_22_29 : IN std_logic ;
      d_arr_mux_22_28 : IN std_logic ;
      d_arr_mux_22_27 : IN std_logic ;
      d_arr_mux_22_26 : IN std_logic ;
      d_arr_mux_22_25 : IN std_logic ;
      d_arr_mux_22_24 : IN std_logic ;
      d_arr_mux_22_23 : IN std_logic ;
      d_arr_mux_22_22 : IN std_logic ;
      d_arr_mux_22_21 : IN std_logic ;
      d_arr_mux_22_20 : IN std_logic ;
      d_arr_mux_22_19 : IN std_logic ;
      d_arr_mux_22_18 : IN std_logic ;
      d_arr_mux_22_17 : IN std_logic ;
      d_arr_mux_22_16 : IN std_logic ;
      d_arr_mux_22_15 : IN std_logic ;
      d_arr_mux_22_14 : IN std_logic ;
      d_arr_mux_22_13 : IN std_logic ;
      d_arr_mux_22_12 : IN std_logic ;
      d_arr_mux_22_11 : IN std_logic ;
      d_arr_mux_22_10 : IN std_logic ;
      d_arr_mux_22_9 : IN std_logic ;
      d_arr_mux_22_8 : IN std_logic ;
      d_arr_mux_22_7 : IN std_logic ;
      d_arr_mux_22_6 : IN std_logic ;
      d_arr_mux_22_5 : IN std_logic ;
      d_arr_mux_22_4 : IN std_logic ;
      d_arr_mux_22_3 : IN std_logic ;
      d_arr_mux_22_2 : IN std_logic ;
      d_arr_mux_22_1 : IN std_logic ;
      d_arr_mux_22_0 : IN std_logic ;
      d_arr_mux_23_31 : IN std_logic ;
      d_arr_mux_23_30 : IN std_logic ;
      d_arr_mux_23_29 : IN std_logic ;
      d_arr_mux_23_28 : IN std_logic ;
      d_arr_mux_23_27 : IN std_logic ;
      d_arr_mux_23_26 : IN std_logic ;
      d_arr_mux_23_25 : IN std_logic ;
      d_arr_mux_23_24 : IN std_logic ;
      d_arr_mux_23_23 : IN std_logic ;
      d_arr_mux_23_22 : IN std_logic ;
      d_arr_mux_23_21 : IN std_logic ;
      d_arr_mux_23_20 : IN std_logic ;
      d_arr_mux_23_19 : IN std_logic ;
      d_arr_mux_23_18 : IN std_logic ;
      d_arr_mux_23_17 : IN std_logic ;
      d_arr_mux_23_16 : IN std_logic ;
      d_arr_mux_23_15 : IN std_logic ;
      d_arr_mux_23_14 : IN std_logic ;
      d_arr_mux_23_13 : IN std_logic ;
      d_arr_mux_23_12 : IN std_logic ;
      d_arr_mux_23_11 : IN std_logic ;
      d_arr_mux_23_10 : IN std_logic ;
      d_arr_mux_23_9 : IN std_logic ;
      d_arr_mux_23_8 : IN std_logic ;
      d_arr_mux_23_7 : IN std_logic ;
      d_arr_mux_23_6 : IN std_logic ;
      d_arr_mux_23_5 : IN std_logic ;
      d_arr_mux_23_4 : IN std_logic ;
      d_arr_mux_23_3 : IN std_logic ;
      d_arr_mux_23_2 : IN std_logic ;
      d_arr_mux_23_1 : IN std_logic ;
      d_arr_mux_23_0 : IN std_logic ;
      d_arr_mux_24_31 : IN std_logic ;
      d_arr_mux_24_30 : IN std_logic ;
      d_arr_mux_24_29 : IN std_logic ;
      d_arr_mux_24_28 : IN std_logic ;
      d_arr_mux_24_27 : IN std_logic ;
      d_arr_mux_24_26 : IN std_logic ;
      d_arr_mux_24_25 : IN std_logic ;
      d_arr_mux_24_24 : IN std_logic ;
      d_arr_mux_24_23 : IN std_logic ;
      d_arr_mux_24_22 : IN std_logic ;
      d_arr_mux_24_21 : IN std_logic ;
      d_arr_mux_24_20 : IN std_logic ;
      d_arr_mux_24_19 : IN std_logic ;
      d_arr_mux_24_18 : IN std_logic ;
      d_arr_mux_24_17 : IN std_logic ;
      d_arr_mux_24_16 : IN std_logic ;
      d_arr_mux_24_15 : IN std_logic ;
      d_arr_mux_24_14 : IN std_logic ;
      d_arr_mux_24_13 : IN std_logic ;
      d_arr_mux_24_12 : IN std_logic ;
      d_arr_mux_24_11 : IN std_logic ;
      d_arr_mux_24_10 : IN std_logic ;
      d_arr_mux_24_9 : IN std_logic ;
      d_arr_mux_24_8 : IN std_logic ;
      d_arr_mux_24_7 : IN std_logic ;
      d_arr_mux_24_6 : IN std_logic ;
      d_arr_mux_24_5 : IN std_logic ;
      d_arr_mux_24_4 : IN std_logic ;
      d_arr_mux_24_3 : IN std_logic ;
      d_arr_mux_24_2 : IN std_logic ;
      d_arr_mux_24_1 : IN std_logic ;
      d_arr_mux_24_0 : IN std_logic ;
      d_arr_mul_0_31 : IN std_logic ;
      d_arr_mul_0_30 : IN std_logic ;
      d_arr_mul_0_29 : IN std_logic ;
      d_arr_mul_0_28 : IN std_logic ;
      d_arr_mul_0_27 : IN std_logic ;
      d_arr_mul_0_26 : IN std_logic ;
      d_arr_mul_0_25 : IN std_logic ;
      d_arr_mul_0_24 : IN std_logic ;
      d_arr_mul_0_23 : IN std_logic ;
      d_arr_mul_0_22 : IN std_logic ;
      d_arr_mul_0_21 : IN std_logic ;
      d_arr_mul_0_20 : IN std_logic ;
      d_arr_mul_0_19 : IN std_logic ;
      d_arr_mul_0_18 : IN std_logic ;
      d_arr_mul_0_17 : IN std_logic ;
      d_arr_mul_0_16 : IN std_logic ;
      d_arr_mul_0_15 : IN std_logic ;
      d_arr_mul_0_14 : IN std_logic ;
      d_arr_mul_0_13 : IN std_logic ;
      d_arr_mul_0_12 : IN std_logic ;
      d_arr_mul_0_11 : IN std_logic ;
      d_arr_mul_0_10 : IN std_logic ;
      d_arr_mul_0_9 : IN std_logic ;
      d_arr_mul_0_8 : IN std_logic ;
      d_arr_mul_0_7 : IN std_logic ;
      d_arr_mul_0_6 : IN std_logic ;
      d_arr_mul_0_5 : IN std_logic ;
      d_arr_mul_0_4 : IN std_logic ;
      d_arr_mul_0_3 : IN std_logic ;
      d_arr_mul_0_2 : IN std_logic ;
      d_arr_mul_0_1 : IN std_logic ;
      d_arr_mul_0_0 : IN std_logic ;
      d_arr_mul_1_31 : IN std_logic ;
      d_arr_mul_1_30 : IN std_logic ;
      d_arr_mul_1_29 : IN std_logic ;
      d_arr_mul_1_28 : IN std_logic ;
      d_arr_mul_1_27 : IN std_logic ;
      d_arr_mul_1_26 : IN std_logic ;
      d_arr_mul_1_25 : IN std_logic ;
      d_arr_mul_1_24 : IN std_logic ;
      d_arr_mul_1_23 : IN std_logic ;
      d_arr_mul_1_22 : IN std_logic ;
      d_arr_mul_1_21 : IN std_logic ;
      d_arr_mul_1_20 : IN std_logic ;
      d_arr_mul_1_19 : IN std_logic ;
      d_arr_mul_1_18 : IN std_logic ;
      d_arr_mul_1_17 : IN std_logic ;
      d_arr_mul_1_16 : IN std_logic ;
      d_arr_mul_1_15 : IN std_logic ;
      d_arr_mul_1_14 : IN std_logic ;
      d_arr_mul_1_13 : IN std_logic ;
      d_arr_mul_1_12 : IN std_logic ;
      d_arr_mul_1_11 : IN std_logic ;
      d_arr_mul_1_10 : IN std_logic ;
      d_arr_mul_1_9 : IN std_logic ;
      d_arr_mul_1_8 : IN std_logic ;
      d_arr_mul_1_7 : IN std_logic ;
      d_arr_mul_1_6 : IN std_logic ;
      d_arr_mul_1_5 : IN std_logic ;
      d_arr_mul_1_4 : IN std_logic ;
      d_arr_mul_1_3 : IN std_logic ;
      d_arr_mul_1_2 : IN std_logic ;
      d_arr_mul_1_1 : IN std_logic ;
      d_arr_mul_1_0 : IN std_logic ;
      d_arr_mul_2_31 : IN std_logic ;
      d_arr_mul_2_30 : IN std_logic ;
      d_arr_mul_2_29 : IN std_logic ;
      d_arr_mul_2_28 : IN std_logic ;
      d_arr_mul_2_27 : IN std_logic ;
      d_arr_mul_2_26 : IN std_logic ;
      d_arr_mul_2_25 : IN std_logic ;
      d_arr_mul_2_24 : IN std_logic ;
      d_arr_mul_2_23 : IN std_logic ;
      d_arr_mul_2_22 : IN std_logic ;
      d_arr_mul_2_21 : IN std_logic ;
      d_arr_mul_2_20 : IN std_logic ;
      d_arr_mul_2_19 : IN std_logic ;
      d_arr_mul_2_18 : IN std_logic ;
      d_arr_mul_2_17 : IN std_logic ;
      d_arr_mul_2_16 : IN std_logic ;
      d_arr_mul_2_15 : IN std_logic ;
      d_arr_mul_2_14 : IN std_logic ;
      d_arr_mul_2_13 : IN std_logic ;
      d_arr_mul_2_12 : IN std_logic ;
      d_arr_mul_2_11 : IN std_logic ;
      d_arr_mul_2_10 : IN std_logic ;
      d_arr_mul_2_9 : IN std_logic ;
      d_arr_mul_2_8 : IN std_logic ;
      d_arr_mul_2_7 : IN std_logic ;
      d_arr_mul_2_6 : IN std_logic ;
      d_arr_mul_2_5 : IN std_logic ;
      d_arr_mul_2_4 : IN std_logic ;
      d_arr_mul_2_3 : IN std_logic ;
      d_arr_mul_2_2 : IN std_logic ;
      d_arr_mul_2_1 : IN std_logic ;
      d_arr_mul_2_0 : IN std_logic ;
      d_arr_mul_3_31 : IN std_logic ;
      d_arr_mul_3_30 : IN std_logic ;
      d_arr_mul_3_29 : IN std_logic ;
      d_arr_mul_3_28 : IN std_logic ;
      d_arr_mul_3_27 : IN std_logic ;
      d_arr_mul_3_26 : IN std_logic ;
      d_arr_mul_3_25 : IN std_logic ;
      d_arr_mul_3_24 : IN std_logic ;
      d_arr_mul_3_23 : IN std_logic ;
      d_arr_mul_3_22 : IN std_logic ;
      d_arr_mul_3_21 : IN std_logic ;
      d_arr_mul_3_20 : IN std_logic ;
      d_arr_mul_3_19 : IN std_logic ;
      d_arr_mul_3_18 : IN std_logic ;
      d_arr_mul_3_17 : IN std_logic ;
      d_arr_mul_3_16 : IN std_logic ;
      d_arr_mul_3_15 : IN std_logic ;
      d_arr_mul_3_14 : IN std_logic ;
      d_arr_mul_3_13 : IN std_logic ;
      d_arr_mul_3_12 : IN std_logic ;
      d_arr_mul_3_11 : IN std_logic ;
      d_arr_mul_3_10 : IN std_logic ;
      d_arr_mul_3_9 : IN std_logic ;
      d_arr_mul_3_8 : IN std_logic ;
      d_arr_mul_3_7 : IN std_logic ;
      d_arr_mul_3_6 : IN std_logic ;
      d_arr_mul_3_5 : IN std_logic ;
      d_arr_mul_3_4 : IN std_logic ;
      d_arr_mul_3_3 : IN std_logic ;
      d_arr_mul_3_2 : IN std_logic ;
      d_arr_mul_3_1 : IN std_logic ;
      d_arr_mul_3_0 : IN std_logic ;
      d_arr_mul_4_31 : IN std_logic ;
      d_arr_mul_4_30 : IN std_logic ;
      d_arr_mul_4_29 : IN std_logic ;
      d_arr_mul_4_28 : IN std_logic ;
      d_arr_mul_4_27 : IN std_logic ;
      d_arr_mul_4_26 : IN std_logic ;
      d_arr_mul_4_25 : IN std_logic ;
      d_arr_mul_4_24 : IN std_logic ;
      d_arr_mul_4_23 : IN std_logic ;
      d_arr_mul_4_22 : IN std_logic ;
      d_arr_mul_4_21 : IN std_logic ;
      d_arr_mul_4_20 : IN std_logic ;
      d_arr_mul_4_19 : IN std_logic ;
      d_arr_mul_4_18 : IN std_logic ;
      d_arr_mul_4_17 : IN std_logic ;
      d_arr_mul_4_16 : IN std_logic ;
      d_arr_mul_4_15 : IN std_logic ;
      d_arr_mul_4_14 : IN std_logic ;
      d_arr_mul_4_13 : IN std_logic ;
      d_arr_mul_4_12 : IN std_logic ;
      d_arr_mul_4_11 : IN std_logic ;
      d_arr_mul_4_10 : IN std_logic ;
      d_arr_mul_4_9 : IN std_logic ;
      d_arr_mul_4_8 : IN std_logic ;
      d_arr_mul_4_7 : IN std_logic ;
      d_arr_mul_4_6 : IN std_logic ;
      d_arr_mul_4_5 : IN std_logic ;
      d_arr_mul_4_4 : IN std_logic ;
      d_arr_mul_4_3 : IN std_logic ;
      d_arr_mul_4_2 : IN std_logic ;
      d_arr_mul_4_1 : IN std_logic ;
      d_arr_mul_4_0 : IN std_logic ;
      d_arr_mul_5_31 : IN std_logic ;
      d_arr_mul_5_30 : IN std_logic ;
      d_arr_mul_5_29 : IN std_logic ;
      d_arr_mul_5_28 : IN std_logic ;
      d_arr_mul_5_27 : IN std_logic ;
      d_arr_mul_5_26 : IN std_logic ;
      d_arr_mul_5_25 : IN std_logic ;
      d_arr_mul_5_24 : IN std_logic ;
      d_arr_mul_5_23 : IN std_logic ;
      d_arr_mul_5_22 : IN std_logic ;
      d_arr_mul_5_21 : IN std_logic ;
      d_arr_mul_5_20 : IN std_logic ;
      d_arr_mul_5_19 : IN std_logic ;
      d_arr_mul_5_18 : IN std_logic ;
      d_arr_mul_5_17 : IN std_logic ;
      d_arr_mul_5_16 : IN std_logic ;
      d_arr_mul_5_15 : IN std_logic ;
      d_arr_mul_5_14 : IN std_logic ;
      d_arr_mul_5_13 : IN std_logic ;
      d_arr_mul_5_12 : IN std_logic ;
      d_arr_mul_5_11 : IN std_logic ;
      d_arr_mul_5_10 : IN std_logic ;
      d_arr_mul_5_9 : IN std_logic ;
      d_arr_mul_5_8 : IN std_logic ;
      d_arr_mul_5_7 : IN std_logic ;
      d_arr_mul_5_6 : IN std_logic ;
      d_arr_mul_5_5 : IN std_logic ;
      d_arr_mul_5_4 : IN std_logic ;
      d_arr_mul_5_3 : IN std_logic ;
      d_arr_mul_5_2 : IN std_logic ;
      d_arr_mul_5_1 : IN std_logic ;
      d_arr_mul_5_0 : IN std_logic ;
      d_arr_mul_6_31 : IN std_logic ;
      d_arr_mul_6_30 : IN std_logic ;
      d_arr_mul_6_29 : IN std_logic ;
      d_arr_mul_6_28 : IN std_logic ;
      d_arr_mul_6_27 : IN std_logic ;
      d_arr_mul_6_26 : IN std_logic ;
      d_arr_mul_6_25 : IN std_logic ;
      d_arr_mul_6_24 : IN std_logic ;
      d_arr_mul_6_23 : IN std_logic ;
      d_arr_mul_6_22 : IN std_logic ;
      d_arr_mul_6_21 : IN std_logic ;
      d_arr_mul_6_20 : IN std_logic ;
      d_arr_mul_6_19 : IN std_logic ;
      d_arr_mul_6_18 : IN std_logic ;
      d_arr_mul_6_17 : IN std_logic ;
      d_arr_mul_6_16 : IN std_logic ;
      d_arr_mul_6_15 : IN std_logic ;
      d_arr_mul_6_14 : IN std_logic ;
      d_arr_mul_6_13 : IN std_logic ;
      d_arr_mul_6_12 : IN std_logic ;
      d_arr_mul_6_11 : IN std_logic ;
      d_arr_mul_6_10 : IN std_logic ;
      d_arr_mul_6_9 : IN std_logic ;
      d_arr_mul_6_8 : IN std_logic ;
      d_arr_mul_6_7 : IN std_logic ;
      d_arr_mul_6_6 : IN std_logic ;
      d_arr_mul_6_5 : IN std_logic ;
      d_arr_mul_6_4 : IN std_logic ;
      d_arr_mul_6_3 : IN std_logic ;
      d_arr_mul_6_2 : IN std_logic ;
      d_arr_mul_6_1 : IN std_logic ;
      d_arr_mul_6_0 : IN std_logic ;
      d_arr_mul_7_31 : IN std_logic ;
      d_arr_mul_7_30 : IN std_logic ;
      d_arr_mul_7_29 : IN std_logic ;
      d_arr_mul_7_28 : IN std_logic ;
      d_arr_mul_7_27 : IN std_logic ;
      d_arr_mul_7_26 : IN std_logic ;
      d_arr_mul_7_25 : IN std_logic ;
      d_arr_mul_7_24 : IN std_logic ;
      d_arr_mul_7_23 : IN std_logic ;
      d_arr_mul_7_22 : IN std_logic ;
      d_arr_mul_7_21 : IN std_logic ;
      d_arr_mul_7_20 : IN std_logic ;
      d_arr_mul_7_19 : IN std_logic ;
      d_arr_mul_7_18 : IN std_logic ;
      d_arr_mul_7_17 : IN std_logic ;
      d_arr_mul_7_16 : IN std_logic ;
      d_arr_mul_7_15 : IN std_logic ;
      d_arr_mul_7_14 : IN std_logic ;
      d_arr_mul_7_13 : IN std_logic ;
      d_arr_mul_7_12 : IN std_logic ;
      d_arr_mul_7_11 : IN std_logic ;
      d_arr_mul_7_10 : IN std_logic ;
      d_arr_mul_7_9 : IN std_logic ;
      d_arr_mul_7_8 : IN std_logic ;
      d_arr_mul_7_7 : IN std_logic ;
      d_arr_mul_7_6 : IN std_logic ;
      d_arr_mul_7_5 : IN std_logic ;
      d_arr_mul_7_4 : IN std_logic ;
      d_arr_mul_7_3 : IN std_logic ;
      d_arr_mul_7_2 : IN std_logic ;
      d_arr_mul_7_1 : IN std_logic ;
      d_arr_mul_7_0 : IN std_logic ;
      d_arr_mul_8_31 : IN std_logic ;
      d_arr_mul_8_30 : IN std_logic ;
      d_arr_mul_8_29 : IN std_logic ;
      d_arr_mul_8_28 : IN std_logic ;
      d_arr_mul_8_27 : IN std_logic ;
      d_arr_mul_8_26 : IN std_logic ;
      d_arr_mul_8_25 : IN std_logic ;
      d_arr_mul_8_24 : IN std_logic ;
      d_arr_mul_8_23 : IN std_logic ;
      d_arr_mul_8_22 : IN std_logic ;
      d_arr_mul_8_21 : IN std_logic ;
      d_arr_mul_8_20 : IN std_logic ;
      d_arr_mul_8_19 : IN std_logic ;
      d_arr_mul_8_18 : IN std_logic ;
      d_arr_mul_8_17 : IN std_logic ;
      d_arr_mul_8_16 : IN std_logic ;
      d_arr_mul_8_15 : IN std_logic ;
      d_arr_mul_8_14 : IN std_logic ;
      d_arr_mul_8_13 : IN std_logic ;
      d_arr_mul_8_12 : IN std_logic ;
      d_arr_mul_8_11 : IN std_logic ;
      d_arr_mul_8_10 : IN std_logic ;
      d_arr_mul_8_9 : IN std_logic ;
      d_arr_mul_8_8 : IN std_logic ;
      d_arr_mul_8_7 : IN std_logic ;
      d_arr_mul_8_6 : IN std_logic ;
      d_arr_mul_8_5 : IN std_logic ;
      d_arr_mul_8_4 : IN std_logic ;
      d_arr_mul_8_3 : IN std_logic ;
      d_arr_mul_8_2 : IN std_logic ;
      d_arr_mul_8_1 : IN std_logic ;
      d_arr_mul_8_0 : IN std_logic ;
      d_arr_mul_9_31 : IN std_logic ;
      d_arr_mul_9_30 : IN std_logic ;
      d_arr_mul_9_29 : IN std_logic ;
      d_arr_mul_9_28 : IN std_logic ;
      d_arr_mul_9_27 : IN std_logic ;
      d_arr_mul_9_26 : IN std_logic ;
      d_arr_mul_9_25 : IN std_logic ;
      d_arr_mul_9_24 : IN std_logic ;
      d_arr_mul_9_23 : IN std_logic ;
      d_arr_mul_9_22 : IN std_logic ;
      d_arr_mul_9_21 : IN std_logic ;
      d_arr_mul_9_20 : IN std_logic ;
      d_arr_mul_9_19 : IN std_logic ;
      d_arr_mul_9_18 : IN std_logic ;
      d_arr_mul_9_17 : IN std_logic ;
      d_arr_mul_9_16 : IN std_logic ;
      d_arr_mul_9_15 : IN std_logic ;
      d_arr_mul_9_14 : IN std_logic ;
      d_arr_mul_9_13 : IN std_logic ;
      d_arr_mul_9_12 : IN std_logic ;
      d_arr_mul_9_11 : IN std_logic ;
      d_arr_mul_9_10 : IN std_logic ;
      d_arr_mul_9_9 : IN std_logic ;
      d_arr_mul_9_8 : IN std_logic ;
      d_arr_mul_9_7 : IN std_logic ;
      d_arr_mul_9_6 : IN std_logic ;
      d_arr_mul_9_5 : IN std_logic ;
      d_arr_mul_9_4 : IN std_logic ;
      d_arr_mul_9_3 : IN std_logic ;
      d_arr_mul_9_2 : IN std_logic ;
      d_arr_mul_9_1 : IN std_logic ;
      d_arr_mul_9_0 : IN std_logic ;
      d_arr_mul_10_31 : IN std_logic ;
      d_arr_mul_10_30 : IN std_logic ;
      d_arr_mul_10_29 : IN std_logic ;
      d_arr_mul_10_28 : IN std_logic ;
      d_arr_mul_10_27 : IN std_logic ;
      d_arr_mul_10_26 : IN std_logic ;
      d_arr_mul_10_25 : IN std_logic ;
      d_arr_mul_10_24 : IN std_logic ;
      d_arr_mul_10_23 : IN std_logic ;
      d_arr_mul_10_22 : IN std_logic ;
      d_arr_mul_10_21 : IN std_logic ;
      d_arr_mul_10_20 : IN std_logic ;
      d_arr_mul_10_19 : IN std_logic ;
      d_arr_mul_10_18 : IN std_logic ;
      d_arr_mul_10_17 : IN std_logic ;
      d_arr_mul_10_16 : IN std_logic ;
      d_arr_mul_10_15 : IN std_logic ;
      d_arr_mul_10_14 : IN std_logic ;
      d_arr_mul_10_13 : IN std_logic ;
      d_arr_mul_10_12 : IN std_logic ;
      d_arr_mul_10_11 : IN std_logic ;
      d_arr_mul_10_10 : IN std_logic ;
      d_arr_mul_10_9 : IN std_logic ;
      d_arr_mul_10_8 : IN std_logic ;
      d_arr_mul_10_7 : IN std_logic ;
      d_arr_mul_10_6 : IN std_logic ;
      d_arr_mul_10_5 : IN std_logic ;
      d_arr_mul_10_4 : IN std_logic ;
      d_arr_mul_10_3 : IN std_logic ;
      d_arr_mul_10_2 : IN std_logic ;
      d_arr_mul_10_1 : IN std_logic ;
      d_arr_mul_10_0 : IN std_logic ;
      d_arr_mul_11_31 : IN std_logic ;
      d_arr_mul_11_30 : IN std_logic ;
      d_arr_mul_11_29 : IN std_logic ;
      d_arr_mul_11_28 : IN std_logic ;
      d_arr_mul_11_27 : IN std_logic ;
      d_arr_mul_11_26 : IN std_logic ;
      d_arr_mul_11_25 : IN std_logic ;
      d_arr_mul_11_24 : IN std_logic ;
      d_arr_mul_11_23 : IN std_logic ;
      d_arr_mul_11_22 : IN std_logic ;
      d_arr_mul_11_21 : IN std_logic ;
      d_arr_mul_11_20 : IN std_logic ;
      d_arr_mul_11_19 : IN std_logic ;
      d_arr_mul_11_18 : IN std_logic ;
      d_arr_mul_11_17 : IN std_logic ;
      d_arr_mul_11_16 : IN std_logic ;
      d_arr_mul_11_15 : IN std_logic ;
      d_arr_mul_11_14 : IN std_logic ;
      d_arr_mul_11_13 : IN std_logic ;
      d_arr_mul_11_12 : IN std_logic ;
      d_arr_mul_11_11 : IN std_logic ;
      d_arr_mul_11_10 : IN std_logic ;
      d_arr_mul_11_9 : IN std_logic ;
      d_arr_mul_11_8 : IN std_logic ;
      d_arr_mul_11_7 : IN std_logic ;
      d_arr_mul_11_6 : IN std_logic ;
      d_arr_mul_11_5 : IN std_logic ;
      d_arr_mul_11_4 : IN std_logic ;
      d_arr_mul_11_3 : IN std_logic ;
      d_arr_mul_11_2 : IN std_logic ;
      d_arr_mul_11_1 : IN std_logic ;
      d_arr_mul_11_0 : IN std_logic ;
      d_arr_mul_12_31 : IN std_logic ;
      d_arr_mul_12_30 : IN std_logic ;
      d_arr_mul_12_29 : IN std_logic ;
      d_arr_mul_12_28 : IN std_logic ;
      d_arr_mul_12_27 : IN std_logic ;
      d_arr_mul_12_26 : IN std_logic ;
      d_arr_mul_12_25 : IN std_logic ;
      d_arr_mul_12_24 : IN std_logic ;
      d_arr_mul_12_23 : IN std_logic ;
      d_arr_mul_12_22 : IN std_logic ;
      d_arr_mul_12_21 : IN std_logic ;
      d_arr_mul_12_20 : IN std_logic ;
      d_arr_mul_12_19 : IN std_logic ;
      d_arr_mul_12_18 : IN std_logic ;
      d_arr_mul_12_17 : IN std_logic ;
      d_arr_mul_12_16 : IN std_logic ;
      d_arr_mul_12_15 : IN std_logic ;
      d_arr_mul_12_14 : IN std_logic ;
      d_arr_mul_12_13 : IN std_logic ;
      d_arr_mul_12_12 : IN std_logic ;
      d_arr_mul_12_11 : IN std_logic ;
      d_arr_mul_12_10 : IN std_logic ;
      d_arr_mul_12_9 : IN std_logic ;
      d_arr_mul_12_8 : IN std_logic ;
      d_arr_mul_12_7 : IN std_logic ;
      d_arr_mul_12_6 : IN std_logic ;
      d_arr_mul_12_5 : IN std_logic ;
      d_arr_mul_12_4 : IN std_logic ;
      d_arr_mul_12_3 : IN std_logic ;
      d_arr_mul_12_2 : IN std_logic ;
      d_arr_mul_12_1 : IN std_logic ;
      d_arr_mul_12_0 : IN std_logic ;
      d_arr_mul_13_31 : IN std_logic ;
      d_arr_mul_13_30 : IN std_logic ;
      d_arr_mul_13_29 : IN std_logic ;
      d_arr_mul_13_28 : IN std_logic ;
      d_arr_mul_13_27 : IN std_logic ;
      d_arr_mul_13_26 : IN std_logic ;
      d_arr_mul_13_25 : IN std_logic ;
      d_arr_mul_13_24 : IN std_logic ;
      d_arr_mul_13_23 : IN std_logic ;
      d_arr_mul_13_22 : IN std_logic ;
      d_arr_mul_13_21 : IN std_logic ;
      d_arr_mul_13_20 : IN std_logic ;
      d_arr_mul_13_19 : IN std_logic ;
      d_arr_mul_13_18 : IN std_logic ;
      d_arr_mul_13_17 : IN std_logic ;
      d_arr_mul_13_16 : IN std_logic ;
      d_arr_mul_13_15 : IN std_logic ;
      d_arr_mul_13_14 : IN std_logic ;
      d_arr_mul_13_13 : IN std_logic ;
      d_arr_mul_13_12 : IN std_logic ;
      d_arr_mul_13_11 : IN std_logic ;
      d_arr_mul_13_10 : IN std_logic ;
      d_arr_mul_13_9 : IN std_logic ;
      d_arr_mul_13_8 : IN std_logic ;
      d_arr_mul_13_7 : IN std_logic ;
      d_arr_mul_13_6 : IN std_logic ;
      d_arr_mul_13_5 : IN std_logic ;
      d_arr_mul_13_4 : IN std_logic ;
      d_arr_mul_13_3 : IN std_logic ;
      d_arr_mul_13_2 : IN std_logic ;
      d_arr_mul_13_1 : IN std_logic ;
      d_arr_mul_13_0 : IN std_logic ;
      d_arr_mul_14_31 : IN std_logic ;
      d_arr_mul_14_30 : IN std_logic ;
      d_arr_mul_14_29 : IN std_logic ;
      d_arr_mul_14_28 : IN std_logic ;
      d_arr_mul_14_27 : IN std_logic ;
      d_arr_mul_14_26 : IN std_logic ;
      d_arr_mul_14_25 : IN std_logic ;
      d_arr_mul_14_24 : IN std_logic ;
      d_arr_mul_14_23 : IN std_logic ;
      d_arr_mul_14_22 : IN std_logic ;
      d_arr_mul_14_21 : IN std_logic ;
      d_arr_mul_14_20 : IN std_logic ;
      d_arr_mul_14_19 : IN std_logic ;
      d_arr_mul_14_18 : IN std_logic ;
      d_arr_mul_14_17 : IN std_logic ;
      d_arr_mul_14_16 : IN std_logic ;
      d_arr_mul_14_15 : IN std_logic ;
      d_arr_mul_14_14 : IN std_logic ;
      d_arr_mul_14_13 : IN std_logic ;
      d_arr_mul_14_12 : IN std_logic ;
      d_arr_mul_14_11 : IN std_logic ;
      d_arr_mul_14_10 : IN std_logic ;
      d_arr_mul_14_9 : IN std_logic ;
      d_arr_mul_14_8 : IN std_logic ;
      d_arr_mul_14_7 : IN std_logic ;
      d_arr_mul_14_6 : IN std_logic ;
      d_arr_mul_14_5 : IN std_logic ;
      d_arr_mul_14_4 : IN std_logic ;
      d_arr_mul_14_3 : IN std_logic ;
      d_arr_mul_14_2 : IN std_logic ;
      d_arr_mul_14_1 : IN std_logic ;
      d_arr_mul_14_0 : IN std_logic ;
      d_arr_mul_15_31 : IN std_logic ;
      d_arr_mul_15_30 : IN std_logic ;
      d_arr_mul_15_29 : IN std_logic ;
      d_arr_mul_15_28 : IN std_logic ;
      d_arr_mul_15_27 : IN std_logic ;
      d_arr_mul_15_26 : IN std_logic ;
      d_arr_mul_15_25 : IN std_logic ;
      d_arr_mul_15_24 : IN std_logic ;
      d_arr_mul_15_23 : IN std_logic ;
      d_arr_mul_15_22 : IN std_logic ;
      d_arr_mul_15_21 : IN std_logic ;
      d_arr_mul_15_20 : IN std_logic ;
      d_arr_mul_15_19 : IN std_logic ;
      d_arr_mul_15_18 : IN std_logic ;
      d_arr_mul_15_17 : IN std_logic ;
      d_arr_mul_15_16 : IN std_logic ;
      d_arr_mul_15_15 : IN std_logic ;
      d_arr_mul_15_14 : IN std_logic ;
      d_arr_mul_15_13 : IN std_logic ;
      d_arr_mul_15_12 : IN std_logic ;
      d_arr_mul_15_11 : IN std_logic ;
      d_arr_mul_15_10 : IN std_logic ;
      d_arr_mul_15_9 : IN std_logic ;
      d_arr_mul_15_8 : IN std_logic ;
      d_arr_mul_15_7 : IN std_logic ;
      d_arr_mul_15_6 : IN std_logic ;
      d_arr_mul_15_5 : IN std_logic ;
      d_arr_mul_15_4 : IN std_logic ;
      d_arr_mul_15_3 : IN std_logic ;
      d_arr_mul_15_2 : IN std_logic ;
      d_arr_mul_15_1 : IN std_logic ;
      d_arr_mul_15_0 : IN std_logic ;
      d_arr_mul_16_31 : IN std_logic ;
      d_arr_mul_16_30 : IN std_logic ;
      d_arr_mul_16_29 : IN std_logic ;
      d_arr_mul_16_28 : IN std_logic ;
      d_arr_mul_16_27 : IN std_logic ;
      d_arr_mul_16_26 : IN std_logic ;
      d_arr_mul_16_25 : IN std_logic ;
      d_arr_mul_16_24 : IN std_logic ;
      d_arr_mul_16_23 : IN std_logic ;
      d_arr_mul_16_22 : IN std_logic ;
      d_arr_mul_16_21 : IN std_logic ;
      d_arr_mul_16_20 : IN std_logic ;
      d_arr_mul_16_19 : IN std_logic ;
      d_arr_mul_16_18 : IN std_logic ;
      d_arr_mul_16_17 : IN std_logic ;
      d_arr_mul_16_16 : IN std_logic ;
      d_arr_mul_16_15 : IN std_logic ;
      d_arr_mul_16_14 : IN std_logic ;
      d_arr_mul_16_13 : IN std_logic ;
      d_arr_mul_16_12 : IN std_logic ;
      d_arr_mul_16_11 : IN std_logic ;
      d_arr_mul_16_10 : IN std_logic ;
      d_arr_mul_16_9 : IN std_logic ;
      d_arr_mul_16_8 : IN std_logic ;
      d_arr_mul_16_7 : IN std_logic ;
      d_arr_mul_16_6 : IN std_logic ;
      d_arr_mul_16_5 : IN std_logic ;
      d_arr_mul_16_4 : IN std_logic ;
      d_arr_mul_16_3 : IN std_logic ;
      d_arr_mul_16_2 : IN std_logic ;
      d_arr_mul_16_1 : IN std_logic ;
      d_arr_mul_16_0 : IN std_logic ;
      d_arr_mul_17_31 : IN std_logic ;
      d_arr_mul_17_30 : IN std_logic ;
      d_arr_mul_17_29 : IN std_logic ;
      d_arr_mul_17_28 : IN std_logic ;
      d_arr_mul_17_27 : IN std_logic ;
      d_arr_mul_17_26 : IN std_logic ;
      d_arr_mul_17_25 : IN std_logic ;
      d_arr_mul_17_24 : IN std_logic ;
      d_arr_mul_17_23 : IN std_logic ;
      d_arr_mul_17_22 : IN std_logic ;
      d_arr_mul_17_21 : IN std_logic ;
      d_arr_mul_17_20 : IN std_logic ;
      d_arr_mul_17_19 : IN std_logic ;
      d_arr_mul_17_18 : IN std_logic ;
      d_arr_mul_17_17 : IN std_logic ;
      d_arr_mul_17_16 : IN std_logic ;
      d_arr_mul_17_15 : IN std_logic ;
      d_arr_mul_17_14 : IN std_logic ;
      d_arr_mul_17_13 : IN std_logic ;
      d_arr_mul_17_12 : IN std_logic ;
      d_arr_mul_17_11 : IN std_logic ;
      d_arr_mul_17_10 : IN std_logic ;
      d_arr_mul_17_9 : IN std_logic ;
      d_arr_mul_17_8 : IN std_logic ;
      d_arr_mul_17_7 : IN std_logic ;
      d_arr_mul_17_6 : IN std_logic ;
      d_arr_mul_17_5 : IN std_logic ;
      d_arr_mul_17_4 : IN std_logic ;
      d_arr_mul_17_3 : IN std_logic ;
      d_arr_mul_17_2 : IN std_logic ;
      d_arr_mul_17_1 : IN std_logic ;
      d_arr_mul_17_0 : IN std_logic ;
      d_arr_mul_18_31 : IN std_logic ;
      d_arr_mul_18_30 : IN std_logic ;
      d_arr_mul_18_29 : IN std_logic ;
      d_arr_mul_18_28 : IN std_logic ;
      d_arr_mul_18_27 : IN std_logic ;
      d_arr_mul_18_26 : IN std_logic ;
      d_arr_mul_18_25 : IN std_logic ;
      d_arr_mul_18_24 : IN std_logic ;
      d_arr_mul_18_23 : IN std_logic ;
      d_arr_mul_18_22 : IN std_logic ;
      d_arr_mul_18_21 : IN std_logic ;
      d_arr_mul_18_20 : IN std_logic ;
      d_arr_mul_18_19 : IN std_logic ;
      d_arr_mul_18_18 : IN std_logic ;
      d_arr_mul_18_17 : IN std_logic ;
      d_arr_mul_18_16 : IN std_logic ;
      d_arr_mul_18_15 : IN std_logic ;
      d_arr_mul_18_14 : IN std_logic ;
      d_arr_mul_18_13 : IN std_logic ;
      d_arr_mul_18_12 : IN std_logic ;
      d_arr_mul_18_11 : IN std_logic ;
      d_arr_mul_18_10 : IN std_logic ;
      d_arr_mul_18_9 : IN std_logic ;
      d_arr_mul_18_8 : IN std_logic ;
      d_arr_mul_18_7 : IN std_logic ;
      d_arr_mul_18_6 : IN std_logic ;
      d_arr_mul_18_5 : IN std_logic ;
      d_arr_mul_18_4 : IN std_logic ;
      d_arr_mul_18_3 : IN std_logic ;
      d_arr_mul_18_2 : IN std_logic ;
      d_arr_mul_18_1 : IN std_logic ;
      d_arr_mul_18_0 : IN std_logic ;
      d_arr_mul_19_31 : IN std_logic ;
      d_arr_mul_19_30 : IN std_logic ;
      d_arr_mul_19_29 : IN std_logic ;
      d_arr_mul_19_28 : IN std_logic ;
      d_arr_mul_19_27 : IN std_logic ;
      d_arr_mul_19_26 : IN std_logic ;
      d_arr_mul_19_25 : IN std_logic ;
      d_arr_mul_19_24 : IN std_logic ;
      d_arr_mul_19_23 : IN std_logic ;
      d_arr_mul_19_22 : IN std_logic ;
      d_arr_mul_19_21 : IN std_logic ;
      d_arr_mul_19_20 : IN std_logic ;
      d_arr_mul_19_19 : IN std_logic ;
      d_arr_mul_19_18 : IN std_logic ;
      d_arr_mul_19_17 : IN std_logic ;
      d_arr_mul_19_16 : IN std_logic ;
      d_arr_mul_19_15 : IN std_logic ;
      d_arr_mul_19_14 : IN std_logic ;
      d_arr_mul_19_13 : IN std_logic ;
      d_arr_mul_19_12 : IN std_logic ;
      d_arr_mul_19_11 : IN std_logic ;
      d_arr_mul_19_10 : IN std_logic ;
      d_arr_mul_19_9 : IN std_logic ;
      d_arr_mul_19_8 : IN std_logic ;
      d_arr_mul_19_7 : IN std_logic ;
      d_arr_mul_19_6 : IN std_logic ;
      d_arr_mul_19_5 : IN std_logic ;
      d_arr_mul_19_4 : IN std_logic ;
      d_arr_mul_19_3 : IN std_logic ;
      d_arr_mul_19_2 : IN std_logic ;
      d_arr_mul_19_1 : IN std_logic ;
      d_arr_mul_19_0 : IN std_logic ;
      d_arr_mul_20_31 : IN std_logic ;
      d_arr_mul_20_30 : IN std_logic ;
      d_arr_mul_20_29 : IN std_logic ;
      d_arr_mul_20_28 : IN std_logic ;
      d_arr_mul_20_27 : IN std_logic ;
      d_arr_mul_20_26 : IN std_logic ;
      d_arr_mul_20_25 : IN std_logic ;
      d_arr_mul_20_24 : IN std_logic ;
      d_arr_mul_20_23 : IN std_logic ;
      d_arr_mul_20_22 : IN std_logic ;
      d_arr_mul_20_21 : IN std_logic ;
      d_arr_mul_20_20 : IN std_logic ;
      d_arr_mul_20_19 : IN std_logic ;
      d_arr_mul_20_18 : IN std_logic ;
      d_arr_mul_20_17 : IN std_logic ;
      d_arr_mul_20_16 : IN std_logic ;
      d_arr_mul_20_15 : IN std_logic ;
      d_arr_mul_20_14 : IN std_logic ;
      d_arr_mul_20_13 : IN std_logic ;
      d_arr_mul_20_12 : IN std_logic ;
      d_arr_mul_20_11 : IN std_logic ;
      d_arr_mul_20_10 : IN std_logic ;
      d_arr_mul_20_9 : IN std_logic ;
      d_arr_mul_20_8 : IN std_logic ;
      d_arr_mul_20_7 : IN std_logic ;
      d_arr_mul_20_6 : IN std_logic ;
      d_arr_mul_20_5 : IN std_logic ;
      d_arr_mul_20_4 : IN std_logic ;
      d_arr_mul_20_3 : IN std_logic ;
      d_arr_mul_20_2 : IN std_logic ;
      d_arr_mul_20_1 : IN std_logic ;
      d_arr_mul_20_0 : IN std_logic ;
      d_arr_mul_21_31 : IN std_logic ;
      d_arr_mul_21_30 : IN std_logic ;
      d_arr_mul_21_29 : IN std_logic ;
      d_arr_mul_21_28 : IN std_logic ;
      d_arr_mul_21_27 : IN std_logic ;
      d_arr_mul_21_26 : IN std_logic ;
      d_arr_mul_21_25 : IN std_logic ;
      d_arr_mul_21_24 : IN std_logic ;
      d_arr_mul_21_23 : IN std_logic ;
      d_arr_mul_21_22 : IN std_logic ;
      d_arr_mul_21_21 : IN std_logic ;
      d_arr_mul_21_20 : IN std_logic ;
      d_arr_mul_21_19 : IN std_logic ;
      d_arr_mul_21_18 : IN std_logic ;
      d_arr_mul_21_17 : IN std_logic ;
      d_arr_mul_21_16 : IN std_logic ;
      d_arr_mul_21_15 : IN std_logic ;
      d_arr_mul_21_14 : IN std_logic ;
      d_arr_mul_21_13 : IN std_logic ;
      d_arr_mul_21_12 : IN std_logic ;
      d_arr_mul_21_11 : IN std_logic ;
      d_arr_mul_21_10 : IN std_logic ;
      d_arr_mul_21_9 : IN std_logic ;
      d_arr_mul_21_8 : IN std_logic ;
      d_arr_mul_21_7 : IN std_logic ;
      d_arr_mul_21_6 : IN std_logic ;
      d_arr_mul_21_5 : IN std_logic ;
      d_arr_mul_21_4 : IN std_logic ;
      d_arr_mul_21_3 : IN std_logic ;
      d_arr_mul_21_2 : IN std_logic ;
      d_arr_mul_21_1 : IN std_logic ;
      d_arr_mul_21_0 : IN std_logic ;
      d_arr_mul_22_31 : IN std_logic ;
      d_arr_mul_22_30 : IN std_logic ;
      d_arr_mul_22_29 : IN std_logic ;
      d_arr_mul_22_28 : IN std_logic ;
      d_arr_mul_22_27 : IN std_logic ;
      d_arr_mul_22_26 : IN std_logic ;
      d_arr_mul_22_25 : IN std_logic ;
      d_arr_mul_22_24 : IN std_logic ;
      d_arr_mul_22_23 : IN std_logic ;
      d_arr_mul_22_22 : IN std_logic ;
      d_arr_mul_22_21 : IN std_logic ;
      d_arr_mul_22_20 : IN std_logic ;
      d_arr_mul_22_19 : IN std_logic ;
      d_arr_mul_22_18 : IN std_logic ;
      d_arr_mul_22_17 : IN std_logic ;
      d_arr_mul_22_16 : IN std_logic ;
      d_arr_mul_22_15 : IN std_logic ;
      d_arr_mul_22_14 : IN std_logic ;
      d_arr_mul_22_13 : IN std_logic ;
      d_arr_mul_22_12 : IN std_logic ;
      d_arr_mul_22_11 : IN std_logic ;
      d_arr_mul_22_10 : IN std_logic ;
      d_arr_mul_22_9 : IN std_logic ;
      d_arr_mul_22_8 : IN std_logic ;
      d_arr_mul_22_7 : IN std_logic ;
      d_arr_mul_22_6 : IN std_logic ;
      d_arr_mul_22_5 : IN std_logic ;
      d_arr_mul_22_4 : IN std_logic ;
      d_arr_mul_22_3 : IN std_logic ;
      d_arr_mul_22_2 : IN std_logic ;
      d_arr_mul_22_1 : IN std_logic ;
      d_arr_mul_22_0 : IN std_logic ;
      d_arr_mul_23_31 : IN std_logic ;
      d_arr_mul_23_30 : IN std_logic ;
      d_arr_mul_23_29 : IN std_logic ;
      d_arr_mul_23_28 : IN std_logic ;
      d_arr_mul_23_27 : IN std_logic ;
      d_arr_mul_23_26 : IN std_logic ;
      d_arr_mul_23_25 : IN std_logic ;
      d_arr_mul_23_24 : IN std_logic ;
      d_arr_mul_23_23 : IN std_logic ;
      d_arr_mul_23_22 : IN std_logic ;
      d_arr_mul_23_21 : IN std_logic ;
      d_arr_mul_23_20 : IN std_logic ;
      d_arr_mul_23_19 : IN std_logic ;
      d_arr_mul_23_18 : IN std_logic ;
      d_arr_mul_23_17 : IN std_logic ;
      d_arr_mul_23_16 : IN std_logic ;
      d_arr_mul_23_15 : IN std_logic ;
      d_arr_mul_23_14 : IN std_logic ;
      d_arr_mul_23_13 : IN std_logic ;
      d_arr_mul_23_12 : IN std_logic ;
      d_arr_mul_23_11 : IN std_logic ;
      d_arr_mul_23_10 : IN std_logic ;
      d_arr_mul_23_9 : IN std_logic ;
      d_arr_mul_23_8 : IN std_logic ;
      d_arr_mul_23_7 : IN std_logic ;
      d_arr_mul_23_6 : IN std_logic ;
      d_arr_mul_23_5 : IN std_logic ;
      d_arr_mul_23_4 : IN std_logic ;
      d_arr_mul_23_3 : IN std_logic ;
      d_arr_mul_23_2 : IN std_logic ;
      d_arr_mul_23_1 : IN std_logic ;
      d_arr_mul_23_0 : IN std_logic ;
      d_arr_mul_24_31 : IN std_logic ;
      d_arr_mul_24_30 : IN std_logic ;
      d_arr_mul_24_29 : IN std_logic ;
      d_arr_mul_24_28 : IN std_logic ;
      d_arr_mul_24_27 : IN std_logic ;
      d_arr_mul_24_26 : IN std_logic ;
      d_arr_mul_24_25 : IN std_logic ;
      d_arr_mul_24_24 : IN std_logic ;
      d_arr_mul_24_23 : IN std_logic ;
      d_arr_mul_24_22 : IN std_logic ;
      d_arr_mul_24_21 : IN std_logic ;
      d_arr_mul_24_20 : IN std_logic ;
      d_arr_mul_24_19 : IN std_logic ;
      d_arr_mul_24_18 : IN std_logic ;
      d_arr_mul_24_17 : IN std_logic ;
      d_arr_mul_24_16 : IN std_logic ;
      d_arr_mul_24_15 : IN std_logic ;
      d_arr_mul_24_14 : IN std_logic ;
      d_arr_mul_24_13 : IN std_logic ;
      d_arr_mul_24_12 : IN std_logic ;
      d_arr_mul_24_11 : IN std_logic ;
      d_arr_mul_24_10 : IN std_logic ;
      d_arr_mul_24_9 : IN std_logic ;
      d_arr_mul_24_8 : IN std_logic ;
      d_arr_mul_24_7 : IN std_logic ;
      d_arr_mul_24_6 : IN std_logic ;
      d_arr_mul_24_5 : IN std_logic ;
      d_arr_mul_24_4 : IN std_logic ;
      d_arr_mul_24_3 : IN std_logic ;
      d_arr_mul_24_2 : IN std_logic ;
      d_arr_mul_24_1 : IN std_logic ;
      d_arr_mul_24_0 : IN std_logic ;
      d_arr_add_0_31 : IN std_logic ;
      d_arr_add_0_30 : IN std_logic ;
      d_arr_add_0_29 : IN std_logic ;
      d_arr_add_0_28 : IN std_logic ;
      d_arr_add_0_27 : IN std_logic ;
      d_arr_add_0_26 : IN std_logic ;
      d_arr_add_0_25 : IN std_logic ;
      d_arr_add_0_24 : IN std_logic ;
      d_arr_add_0_23 : IN std_logic ;
      d_arr_add_0_22 : IN std_logic ;
      d_arr_add_0_21 : IN std_logic ;
      d_arr_add_0_20 : IN std_logic ;
      d_arr_add_0_19 : IN std_logic ;
      d_arr_add_0_18 : IN std_logic ;
      d_arr_add_0_17 : IN std_logic ;
      d_arr_add_0_16 : IN std_logic ;
      d_arr_add_0_15 : IN std_logic ;
      d_arr_add_0_14 : IN std_logic ;
      d_arr_add_0_13 : IN std_logic ;
      d_arr_add_0_12 : IN std_logic ;
      d_arr_add_0_11 : IN std_logic ;
      d_arr_add_0_10 : IN std_logic ;
      d_arr_add_0_9 : IN std_logic ;
      d_arr_add_0_8 : IN std_logic ;
      d_arr_add_0_7 : IN std_logic ;
      d_arr_add_0_6 : IN std_logic ;
      d_arr_add_0_5 : IN std_logic ;
      d_arr_add_0_4 : IN std_logic ;
      d_arr_add_0_3 : IN std_logic ;
      d_arr_add_0_2 : IN std_logic ;
      d_arr_add_0_1 : IN std_logic ;
      d_arr_add_0_0 : IN std_logic ;
      d_arr_add_1_31 : IN std_logic ;
      d_arr_add_1_30 : IN std_logic ;
      d_arr_add_1_29 : IN std_logic ;
      d_arr_add_1_28 : IN std_logic ;
      d_arr_add_1_27 : IN std_logic ;
      d_arr_add_1_26 : IN std_logic ;
      d_arr_add_1_25 : IN std_logic ;
      d_arr_add_1_24 : IN std_logic ;
      d_arr_add_1_23 : IN std_logic ;
      d_arr_add_1_22 : IN std_logic ;
      d_arr_add_1_21 : IN std_logic ;
      d_arr_add_1_20 : IN std_logic ;
      d_arr_add_1_19 : IN std_logic ;
      d_arr_add_1_18 : IN std_logic ;
      d_arr_add_1_17 : IN std_logic ;
      d_arr_add_1_16 : IN std_logic ;
      d_arr_add_1_15 : IN std_logic ;
      d_arr_add_1_14 : IN std_logic ;
      d_arr_add_1_13 : IN std_logic ;
      d_arr_add_1_12 : IN std_logic ;
      d_arr_add_1_11 : IN std_logic ;
      d_arr_add_1_10 : IN std_logic ;
      d_arr_add_1_9 : IN std_logic ;
      d_arr_add_1_8 : IN std_logic ;
      d_arr_add_1_7 : IN std_logic ;
      d_arr_add_1_6 : IN std_logic ;
      d_arr_add_1_5 : IN std_logic ;
      d_arr_add_1_4 : IN std_logic ;
      d_arr_add_1_3 : IN std_logic ;
      d_arr_add_1_2 : IN std_logic ;
      d_arr_add_1_1 : IN std_logic ;
      d_arr_add_1_0 : IN std_logic ;
      d_arr_add_2_31 : IN std_logic ;
      d_arr_add_2_30 : IN std_logic ;
      d_arr_add_2_29 : IN std_logic ;
      d_arr_add_2_28 : IN std_logic ;
      d_arr_add_2_27 : IN std_logic ;
      d_arr_add_2_26 : IN std_logic ;
      d_arr_add_2_25 : IN std_logic ;
      d_arr_add_2_24 : IN std_logic ;
      d_arr_add_2_23 : IN std_logic ;
      d_arr_add_2_22 : IN std_logic ;
      d_arr_add_2_21 : IN std_logic ;
      d_arr_add_2_20 : IN std_logic ;
      d_arr_add_2_19 : IN std_logic ;
      d_arr_add_2_18 : IN std_logic ;
      d_arr_add_2_17 : IN std_logic ;
      d_arr_add_2_16 : IN std_logic ;
      d_arr_add_2_15 : IN std_logic ;
      d_arr_add_2_14 : IN std_logic ;
      d_arr_add_2_13 : IN std_logic ;
      d_arr_add_2_12 : IN std_logic ;
      d_arr_add_2_11 : IN std_logic ;
      d_arr_add_2_10 : IN std_logic ;
      d_arr_add_2_9 : IN std_logic ;
      d_arr_add_2_8 : IN std_logic ;
      d_arr_add_2_7 : IN std_logic ;
      d_arr_add_2_6 : IN std_logic ;
      d_arr_add_2_5 : IN std_logic ;
      d_arr_add_2_4 : IN std_logic ;
      d_arr_add_2_3 : IN std_logic ;
      d_arr_add_2_2 : IN std_logic ;
      d_arr_add_2_1 : IN std_logic ;
      d_arr_add_2_0 : IN std_logic ;
      d_arr_add_3_31 : IN std_logic ;
      d_arr_add_3_30 : IN std_logic ;
      d_arr_add_3_29 : IN std_logic ;
      d_arr_add_3_28 : IN std_logic ;
      d_arr_add_3_27 : IN std_logic ;
      d_arr_add_3_26 : IN std_logic ;
      d_arr_add_3_25 : IN std_logic ;
      d_arr_add_3_24 : IN std_logic ;
      d_arr_add_3_23 : IN std_logic ;
      d_arr_add_3_22 : IN std_logic ;
      d_arr_add_3_21 : IN std_logic ;
      d_arr_add_3_20 : IN std_logic ;
      d_arr_add_3_19 : IN std_logic ;
      d_arr_add_3_18 : IN std_logic ;
      d_arr_add_3_17 : IN std_logic ;
      d_arr_add_3_16 : IN std_logic ;
      d_arr_add_3_15 : IN std_logic ;
      d_arr_add_3_14 : IN std_logic ;
      d_arr_add_3_13 : IN std_logic ;
      d_arr_add_3_12 : IN std_logic ;
      d_arr_add_3_11 : IN std_logic ;
      d_arr_add_3_10 : IN std_logic ;
      d_arr_add_3_9 : IN std_logic ;
      d_arr_add_3_8 : IN std_logic ;
      d_arr_add_3_7 : IN std_logic ;
      d_arr_add_3_6 : IN std_logic ;
      d_arr_add_3_5 : IN std_logic ;
      d_arr_add_3_4 : IN std_logic ;
      d_arr_add_3_3 : IN std_logic ;
      d_arr_add_3_2 : IN std_logic ;
      d_arr_add_3_1 : IN std_logic ;
      d_arr_add_3_0 : IN std_logic ;
      d_arr_add_4_31 : IN std_logic ;
      d_arr_add_4_30 : IN std_logic ;
      d_arr_add_4_29 : IN std_logic ;
      d_arr_add_4_28 : IN std_logic ;
      d_arr_add_4_27 : IN std_logic ;
      d_arr_add_4_26 : IN std_logic ;
      d_arr_add_4_25 : IN std_logic ;
      d_arr_add_4_24 : IN std_logic ;
      d_arr_add_4_23 : IN std_logic ;
      d_arr_add_4_22 : IN std_logic ;
      d_arr_add_4_21 : IN std_logic ;
      d_arr_add_4_20 : IN std_logic ;
      d_arr_add_4_19 : IN std_logic ;
      d_arr_add_4_18 : IN std_logic ;
      d_arr_add_4_17 : IN std_logic ;
      d_arr_add_4_16 : IN std_logic ;
      d_arr_add_4_15 : IN std_logic ;
      d_arr_add_4_14 : IN std_logic ;
      d_arr_add_4_13 : IN std_logic ;
      d_arr_add_4_12 : IN std_logic ;
      d_arr_add_4_11 : IN std_logic ;
      d_arr_add_4_10 : IN std_logic ;
      d_arr_add_4_9 : IN std_logic ;
      d_arr_add_4_8 : IN std_logic ;
      d_arr_add_4_7 : IN std_logic ;
      d_arr_add_4_6 : IN std_logic ;
      d_arr_add_4_5 : IN std_logic ;
      d_arr_add_4_4 : IN std_logic ;
      d_arr_add_4_3 : IN std_logic ;
      d_arr_add_4_2 : IN std_logic ;
      d_arr_add_4_1 : IN std_logic ;
      d_arr_add_4_0 : IN std_logic ;
      d_arr_add_5_31 : IN std_logic ;
      d_arr_add_5_30 : IN std_logic ;
      d_arr_add_5_29 : IN std_logic ;
      d_arr_add_5_28 : IN std_logic ;
      d_arr_add_5_27 : IN std_logic ;
      d_arr_add_5_26 : IN std_logic ;
      d_arr_add_5_25 : IN std_logic ;
      d_arr_add_5_24 : IN std_logic ;
      d_arr_add_5_23 : IN std_logic ;
      d_arr_add_5_22 : IN std_logic ;
      d_arr_add_5_21 : IN std_logic ;
      d_arr_add_5_20 : IN std_logic ;
      d_arr_add_5_19 : IN std_logic ;
      d_arr_add_5_18 : IN std_logic ;
      d_arr_add_5_17 : IN std_logic ;
      d_arr_add_5_16 : IN std_logic ;
      d_arr_add_5_15 : IN std_logic ;
      d_arr_add_5_14 : IN std_logic ;
      d_arr_add_5_13 : IN std_logic ;
      d_arr_add_5_12 : IN std_logic ;
      d_arr_add_5_11 : IN std_logic ;
      d_arr_add_5_10 : IN std_logic ;
      d_arr_add_5_9 : IN std_logic ;
      d_arr_add_5_8 : IN std_logic ;
      d_arr_add_5_7 : IN std_logic ;
      d_arr_add_5_6 : IN std_logic ;
      d_arr_add_5_5 : IN std_logic ;
      d_arr_add_5_4 : IN std_logic ;
      d_arr_add_5_3 : IN std_logic ;
      d_arr_add_5_2 : IN std_logic ;
      d_arr_add_5_1 : IN std_logic ;
      d_arr_add_5_0 : IN std_logic ;
      d_arr_add_6_31 : IN std_logic ;
      d_arr_add_6_30 : IN std_logic ;
      d_arr_add_6_29 : IN std_logic ;
      d_arr_add_6_28 : IN std_logic ;
      d_arr_add_6_27 : IN std_logic ;
      d_arr_add_6_26 : IN std_logic ;
      d_arr_add_6_25 : IN std_logic ;
      d_arr_add_6_24 : IN std_logic ;
      d_arr_add_6_23 : IN std_logic ;
      d_arr_add_6_22 : IN std_logic ;
      d_arr_add_6_21 : IN std_logic ;
      d_arr_add_6_20 : IN std_logic ;
      d_arr_add_6_19 : IN std_logic ;
      d_arr_add_6_18 : IN std_logic ;
      d_arr_add_6_17 : IN std_logic ;
      d_arr_add_6_16 : IN std_logic ;
      d_arr_add_6_15 : IN std_logic ;
      d_arr_add_6_14 : IN std_logic ;
      d_arr_add_6_13 : IN std_logic ;
      d_arr_add_6_12 : IN std_logic ;
      d_arr_add_6_11 : IN std_logic ;
      d_arr_add_6_10 : IN std_logic ;
      d_arr_add_6_9 : IN std_logic ;
      d_arr_add_6_8 : IN std_logic ;
      d_arr_add_6_7 : IN std_logic ;
      d_arr_add_6_6 : IN std_logic ;
      d_arr_add_6_5 : IN std_logic ;
      d_arr_add_6_4 : IN std_logic ;
      d_arr_add_6_3 : IN std_logic ;
      d_arr_add_6_2 : IN std_logic ;
      d_arr_add_6_1 : IN std_logic ;
      d_arr_add_6_0 : IN std_logic ;
      d_arr_add_7_31 : IN std_logic ;
      d_arr_add_7_30 : IN std_logic ;
      d_arr_add_7_29 : IN std_logic ;
      d_arr_add_7_28 : IN std_logic ;
      d_arr_add_7_27 : IN std_logic ;
      d_arr_add_7_26 : IN std_logic ;
      d_arr_add_7_25 : IN std_logic ;
      d_arr_add_7_24 : IN std_logic ;
      d_arr_add_7_23 : IN std_logic ;
      d_arr_add_7_22 : IN std_logic ;
      d_arr_add_7_21 : IN std_logic ;
      d_arr_add_7_20 : IN std_logic ;
      d_arr_add_7_19 : IN std_logic ;
      d_arr_add_7_18 : IN std_logic ;
      d_arr_add_7_17 : IN std_logic ;
      d_arr_add_7_16 : IN std_logic ;
      d_arr_add_7_15 : IN std_logic ;
      d_arr_add_7_14 : IN std_logic ;
      d_arr_add_7_13 : IN std_logic ;
      d_arr_add_7_12 : IN std_logic ;
      d_arr_add_7_11 : IN std_logic ;
      d_arr_add_7_10 : IN std_logic ;
      d_arr_add_7_9 : IN std_logic ;
      d_arr_add_7_8 : IN std_logic ;
      d_arr_add_7_7 : IN std_logic ;
      d_arr_add_7_6 : IN std_logic ;
      d_arr_add_7_5 : IN std_logic ;
      d_arr_add_7_4 : IN std_logic ;
      d_arr_add_7_3 : IN std_logic ;
      d_arr_add_7_2 : IN std_logic ;
      d_arr_add_7_1 : IN std_logic ;
      d_arr_add_7_0 : IN std_logic ;
      d_arr_add_8_31 : IN std_logic ;
      d_arr_add_8_30 : IN std_logic ;
      d_arr_add_8_29 : IN std_logic ;
      d_arr_add_8_28 : IN std_logic ;
      d_arr_add_8_27 : IN std_logic ;
      d_arr_add_8_26 : IN std_logic ;
      d_arr_add_8_25 : IN std_logic ;
      d_arr_add_8_24 : IN std_logic ;
      d_arr_add_8_23 : IN std_logic ;
      d_arr_add_8_22 : IN std_logic ;
      d_arr_add_8_21 : IN std_logic ;
      d_arr_add_8_20 : IN std_logic ;
      d_arr_add_8_19 : IN std_logic ;
      d_arr_add_8_18 : IN std_logic ;
      d_arr_add_8_17 : IN std_logic ;
      d_arr_add_8_16 : IN std_logic ;
      d_arr_add_8_15 : IN std_logic ;
      d_arr_add_8_14 : IN std_logic ;
      d_arr_add_8_13 : IN std_logic ;
      d_arr_add_8_12 : IN std_logic ;
      d_arr_add_8_11 : IN std_logic ;
      d_arr_add_8_10 : IN std_logic ;
      d_arr_add_8_9 : IN std_logic ;
      d_arr_add_8_8 : IN std_logic ;
      d_arr_add_8_7 : IN std_logic ;
      d_arr_add_8_6 : IN std_logic ;
      d_arr_add_8_5 : IN std_logic ;
      d_arr_add_8_4 : IN std_logic ;
      d_arr_add_8_3 : IN std_logic ;
      d_arr_add_8_2 : IN std_logic ;
      d_arr_add_8_1 : IN std_logic ;
      d_arr_add_8_0 : IN std_logic ;
      d_arr_add_9_31 : IN std_logic ;
      d_arr_add_9_30 : IN std_logic ;
      d_arr_add_9_29 : IN std_logic ;
      d_arr_add_9_28 : IN std_logic ;
      d_arr_add_9_27 : IN std_logic ;
      d_arr_add_9_26 : IN std_logic ;
      d_arr_add_9_25 : IN std_logic ;
      d_arr_add_9_24 : IN std_logic ;
      d_arr_add_9_23 : IN std_logic ;
      d_arr_add_9_22 : IN std_logic ;
      d_arr_add_9_21 : IN std_logic ;
      d_arr_add_9_20 : IN std_logic ;
      d_arr_add_9_19 : IN std_logic ;
      d_arr_add_9_18 : IN std_logic ;
      d_arr_add_9_17 : IN std_logic ;
      d_arr_add_9_16 : IN std_logic ;
      d_arr_add_9_15 : IN std_logic ;
      d_arr_add_9_14 : IN std_logic ;
      d_arr_add_9_13 : IN std_logic ;
      d_arr_add_9_12 : IN std_logic ;
      d_arr_add_9_11 : IN std_logic ;
      d_arr_add_9_10 : IN std_logic ;
      d_arr_add_9_9 : IN std_logic ;
      d_arr_add_9_8 : IN std_logic ;
      d_arr_add_9_7 : IN std_logic ;
      d_arr_add_9_6 : IN std_logic ;
      d_arr_add_9_5 : IN std_logic ;
      d_arr_add_9_4 : IN std_logic ;
      d_arr_add_9_3 : IN std_logic ;
      d_arr_add_9_2 : IN std_logic ;
      d_arr_add_9_1 : IN std_logic ;
      d_arr_add_9_0 : IN std_logic ;
      d_arr_add_10_31 : IN std_logic ;
      d_arr_add_10_30 : IN std_logic ;
      d_arr_add_10_29 : IN std_logic ;
      d_arr_add_10_28 : IN std_logic ;
      d_arr_add_10_27 : IN std_logic ;
      d_arr_add_10_26 : IN std_logic ;
      d_arr_add_10_25 : IN std_logic ;
      d_arr_add_10_24 : IN std_logic ;
      d_arr_add_10_23 : IN std_logic ;
      d_arr_add_10_22 : IN std_logic ;
      d_arr_add_10_21 : IN std_logic ;
      d_arr_add_10_20 : IN std_logic ;
      d_arr_add_10_19 : IN std_logic ;
      d_arr_add_10_18 : IN std_logic ;
      d_arr_add_10_17 : IN std_logic ;
      d_arr_add_10_16 : IN std_logic ;
      d_arr_add_10_15 : IN std_logic ;
      d_arr_add_10_14 : IN std_logic ;
      d_arr_add_10_13 : IN std_logic ;
      d_arr_add_10_12 : IN std_logic ;
      d_arr_add_10_11 : IN std_logic ;
      d_arr_add_10_10 : IN std_logic ;
      d_arr_add_10_9 : IN std_logic ;
      d_arr_add_10_8 : IN std_logic ;
      d_arr_add_10_7 : IN std_logic ;
      d_arr_add_10_6 : IN std_logic ;
      d_arr_add_10_5 : IN std_logic ;
      d_arr_add_10_4 : IN std_logic ;
      d_arr_add_10_3 : IN std_logic ;
      d_arr_add_10_2 : IN std_logic ;
      d_arr_add_10_1 : IN std_logic ;
      d_arr_add_10_0 : IN std_logic ;
      d_arr_add_11_31 : IN std_logic ;
      d_arr_add_11_30 : IN std_logic ;
      d_arr_add_11_29 : IN std_logic ;
      d_arr_add_11_28 : IN std_logic ;
      d_arr_add_11_27 : IN std_logic ;
      d_arr_add_11_26 : IN std_logic ;
      d_arr_add_11_25 : IN std_logic ;
      d_arr_add_11_24 : IN std_logic ;
      d_arr_add_11_23 : IN std_logic ;
      d_arr_add_11_22 : IN std_logic ;
      d_arr_add_11_21 : IN std_logic ;
      d_arr_add_11_20 : IN std_logic ;
      d_arr_add_11_19 : IN std_logic ;
      d_arr_add_11_18 : IN std_logic ;
      d_arr_add_11_17 : IN std_logic ;
      d_arr_add_11_16 : IN std_logic ;
      d_arr_add_11_15 : IN std_logic ;
      d_arr_add_11_14 : IN std_logic ;
      d_arr_add_11_13 : IN std_logic ;
      d_arr_add_11_12 : IN std_logic ;
      d_arr_add_11_11 : IN std_logic ;
      d_arr_add_11_10 : IN std_logic ;
      d_arr_add_11_9 : IN std_logic ;
      d_arr_add_11_8 : IN std_logic ;
      d_arr_add_11_7 : IN std_logic ;
      d_arr_add_11_6 : IN std_logic ;
      d_arr_add_11_5 : IN std_logic ;
      d_arr_add_11_4 : IN std_logic ;
      d_arr_add_11_3 : IN std_logic ;
      d_arr_add_11_2 : IN std_logic ;
      d_arr_add_11_1 : IN std_logic ;
      d_arr_add_11_0 : IN std_logic ;
      d_arr_add_12_31 : IN std_logic ;
      d_arr_add_12_30 : IN std_logic ;
      d_arr_add_12_29 : IN std_logic ;
      d_arr_add_12_28 : IN std_logic ;
      d_arr_add_12_27 : IN std_logic ;
      d_arr_add_12_26 : IN std_logic ;
      d_arr_add_12_25 : IN std_logic ;
      d_arr_add_12_24 : IN std_logic ;
      d_arr_add_12_23 : IN std_logic ;
      d_arr_add_12_22 : IN std_logic ;
      d_arr_add_12_21 : IN std_logic ;
      d_arr_add_12_20 : IN std_logic ;
      d_arr_add_12_19 : IN std_logic ;
      d_arr_add_12_18 : IN std_logic ;
      d_arr_add_12_17 : IN std_logic ;
      d_arr_add_12_16 : IN std_logic ;
      d_arr_add_12_15 : IN std_logic ;
      d_arr_add_12_14 : IN std_logic ;
      d_arr_add_12_13 : IN std_logic ;
      d_arr_add_12_12 : IN std_logic ;
      d_arr_add_12_11 : IN std_logic ;
      d_arr_add_12_10 : IN std_logic ;
      d_arr_add_12_9 : IN std_logic ;
      d_arr_add_12_8 : IN std_logic ;
      d_arr_add_12_7 : IN std_logic ;
      d_arr_add_12_6 : IN std_logic ;
      d_arr_add_12_5 : IN std_logic ;
      d_arr_add_12_4 : IN std_logic ;
      d_arr_add_12_3 : IN std_logic ;
      d_arr_add_12_2 : IN std_logic ;
      d_arr_add_12_1 : IN std_logic ;
      d_arr_add_12_0 : IN std_logic ;
      d_arr_add_13_31 : IN std_logic ;
      d_arr_add_13_30 : IN std_logic ;
      d_arr_add_13_29 : IN std_logic ;
      d_arr_add_13_28 : IN std_logic ;
      d_arr_add_13_27 : IN std_logic ;
      d_arr_add_13_26 : IN std_logic ;
      d_arr_add_13_25 : IN std_logic ;
      d_arr_add_13_24 : IN std_logic ;
      d_arr_add_13_23 : IN std_logic ;
      d_arr_add_13_22 : IN std_logic ;
      d_arr_add_13_21 : IN std_logic ;
      d_arr_add_13_20 : IN std_logic ;
      d_arr_add_13_19 : IN std_logic ;
      d_arr_add_13_18 : IN std_logic ;
      d_arr_add_13_17 : IN std_logic ;
      d_arr_add_13_16 : IN std_logic ;
      d_arr_add_13_15 : IN std_logic ;
      d_arr_add_13_14 : IN std_logic ;
      d_arr_add_13_13 : IN std_logic ;
      d_arr_add_13_12 : IN std_logic ;
      d_arr_add_13_11 : IN std_logic ;
      d_arr_add_13_10 : IN std_logic ;
      d_arr_add_13_9 : IN std_logic ;
      d_arr_add_13_8 : IN std_logic ;
      d_arr_add_13_7 : IN std_logic ;
      d_arr_add_13_6 : IN std_logic ;
      d_arr_add_13_5 : IN std_logic ;
      d_arr_add_13_4 : IN std_logic ;
      d_arr_add_13_3 : IN std_logic ;
      d_arr_add_13_2 : IN std_logic ;
      d_arr_add_13_1 : IN std_logic ;
      d_arr_add_13_0 : IN std_logic ;
      d_arr_add_14_31 : IN std_logic ;
      d_arr_add_14_30 : IN std_logic ;
      d_arr_add_14_29 : IN std_logic ;
      d_arr_add_14_28 : IN std_logic ;
      d_arr_add_14_27 : IN std_logic ;
      d_arr_add_14_26 : IN std_logic ;
      d_arr_add_14_25 : IN std_logic ;
      d_arr_add_14_24 : IN std_logic ;
      d_arr_add_14_23 : IN std_logic ;
      d_arr_add_14_22 : IN std_logic ;
      d_arr_add_14_21 : IN std_logic ;
      d_arr_add_14_20 : IN std_logic ;
      d_arr_add_14_19 : IN std_logic ;
      d_arr_add_14_18 : IN std_logic ;
      d_arr_add_14_17 : IN std_logic ;
      d_arr_add_14_16 : IN std_logic ;
      d_arr_add_14_15 : IN std_logic ;
      d_arr_add_14_14 : IN std_logic ;
      d_arr_add_14_13 : IN std_logic ;
      d_arr_add_14_12 : IN std_logic ;
      d_arr_add_14_11 : IN std_logic ;
      d_arr_add_14_10 : IN std_logic ;
      d_arr_add_14_9 : IN std_logic ;
      d_arr_add_14_8 : IN std_logic ;
      d_arr_add_14_7 : IN std_logic ;
      d_arr_add_14_6 : IN std_logic ;
      d_arr_add_14_5 : IN std_logic ;
      d_arr_add_14_4 : IN std_logic ;
      d_arr_add_14_3 : IN std_logic ;
      d_arr_add_14_2 : IN std_logic ;
      d_arr_add_14_1 : IN std_logic ;
      d_arr_add_14_0 : IN std_logic ;
      d_arr_add_15_31 : IN std_logic ;
      d_arr_add_15_30 : IN std_logic ;
      d_arr_add_15_29 : IN std_logic ;
      d_arr_add_15_28 : IN std_logic ;
      d_arr_add_15_27 : IN std_logic ;
      d_arr_add_15_26 : IN std_logic ;
      d_arr_add_15_25 : IN std_logic ;
      d_arr_add_15_24 : IN std_logic ;
      d_arr_add_15_23 : IN std_logic ;
      d_arr_add_15_22 : IN std_logic ;
      d_arr_add_15_21 : IN std_logic ;
      d_arr_add_15_20 : IN std_logic ;
      d_arr_add_15_19 : IN std_logic ;
      d_arr_add_15_18 : IN std_logic ;
      d_arr_add_15_17 : IN std_logic ;
      d_arr_add_15_16 : IN std_logic ;
      d_arr_add_15_15 : IN std_logic ;
      d_arr_add_15_14 : IN std_logic ;
      d_arr_add_15_13 : IN std_logic ;
      d_arr_add_15_12 : IN std_logic ;
      d_arr_add_15_11 : IN std_logic ;
      d_arr_add_15_10 : IN std_logic ;
      d_arr_add_15_9 : IN std_logic ;
      d_arr_add_15_8 : IN std_logic ;
      d_arr_add_15_7 : IN std_logic ;
      d_arr_add_15_6 : IN std_logic ;
      d_arr_add_15_5 : IN std_logic ;
      d_arr_add_15_4 : IN std_logic ;
      d_arr_add_15_3 : IN std_logic ;
      d_arr_add_15_2 : IN std_logic ;
      d_arr_add_15_1 : IN std_logic ;
      d_arr_add_15_0 : IN std_logic ;
      d_arr_add_16_31 : IN std_logic ;
      d_arr_add_16_30 : IN std_logic ;
      d_arr_add_16_29 : IN std_logic ;
      d_arr_add_16_28 : IN std_logic ;
      d_arr_add_16_27 : IN std_logic ;
      d_arr_add_16_26 : IN std_logic ;
      d_arr_add_16_25 : IN std_logic ;
      d_arr_add_16_24 : IN std_logic ;
      d_arr_add_16_23 : IN std_logic ;
      d_arr_add_16_22 : IN std_logic ;
      d_arr_add_16_21 : IN std_logic ;
      d_arr_add_16_20 : IN std_logic ;
      d_arr_add_16_19 : IN std_logic ;
      d_arr_add_16_18 : IN std_logic ;
      d_arr_add_16_17 : IN std_logic ;
      d_arr_add_16_16 : IN std_logic ;
      d_arr_add_16_15 : IN std_logic ;
      d_arr_add_16_14 : IN std_logic ;
      d_arr_add_16_13 : IN std_logic ;
      d_arr_add_16_12 : IN std_logic ;
      d_arr_add_16_11 : IN std_logic ;
      d_arr_add_16_10 : IN std_logic ;
      d_arr_add_16_9 : IN std_logic ;
      d_arr_add_16_8 : IN std_logic ;
      d_arr_add_16_7 : IN std_logic ;
      d_arr_add_16_6 : IN std_logic ;
      d_arr_add_16_5 : IN std_logic ;
      d_arr_add_16_4 : IN std_logic ;
      d_arr_add_16_3 : IN std_logic ;
      d_arr_add_16_2 : IN std_logic ;
      d_arr_add_16_1 : IN std_logic ;
      d_arr_add_16_0 : IN std_logic ;
      d_arr_add_17_31 : IN std_logic ;
      d_arr_add_17_30 : IN std_logic ;
      d_arr_add_17_29 : IN std_logic ;
      d_arr_add_17_28 : IN std_logic ;
      d_arr_add_17_27 : IN std_logic ;
      d_arr_add_17_26 : IN std_logic ;
      d_arr_add_17_25 : IN std_logic ;
      d_arr_add_17_24 : IN std_logic ;
      d_arr_add_17_23 : IN std_logic ;
      d_arr_add_17_22 : IN std_logic ;
      d_arr_add_17_21 : IN std_logic ;
      d_arr_add_17_20 : IN std_logic ;
      d_arr_add_17_19 : IN std_logic ;
      d_arr_add_17_18 : IN std_logic ;
      d_arr_add_17_17 : IN std_logic ;
      d_arr_add_17_16 : IN std_logic ;
      d_arr_add_17_15 : IN std_logic ;
      d_arr_add_17_14 : IN std_logic ;
      d_arr_add_17_13 : IN std_logic ;
      d_arr_add_17_12 : IN std_logic ;
      d_arr_add_17_11 : IN std_logic ;
      d_arr_add_17_10 : IN std_logic ;
      d_arr_add_17_9 : IN std_logic ;
      d_arr_add_17_8 : IN std_logic ;
      d_arr_add_17_7 : IN std_logic ;
      d_arr_add_17_6 : IN std_logic ;
      d_arr_add_17_5 : IN std_logic ;
      d_arr_add_17_4 : IN std_logic ;
      d_arr_add_17_3 : IN std_logic ;
      d_arr_add_17_2 : IN std_logic ;
      d_arr_add_17_1 : IN std_logic ;
      d_arr_add_17_0 : IN std_logic ;
      d_arr_add_18_31 : IN std_logic ;
      d_arr_add_18_30 : IN std_logic ;
      d_arr_add_18_29 : IN std_logic ;
      d_arr_add_18_28 : IN std_logic ;
      d_arr_add_18_27 : IN std_logic ;
      d_arr_add_18_26 : IN std_logic ;
      d_arr_add_18_25 : IN std_logic ;
      d_arr_add_18_24 : IN std_logic ;
      d_arr_add_18_23 : IN std_logic ;
      d_arr_add_18_22 : IN std_logic ;
      d_arr_add_18_21 : IN std_logic ;
      d_arr_add_18_20 : IN std_logic ;
      d_arr_add_18_19 : IN std_logic ;
      d_arr_add_18_18 : IN std_logic ;
      d_arr_add_18_17 : IN std_logic ;
      d_arr_add_18_16 : IN std_logic ;
      d_arr_add_18_15 : IN std_logic ;
      d_arr_add_18_14 : IN std_logic ;
      d_arr_add_18_13 : IN std_logic ;
      d_arr_add_18_12 : IN std_logic ;
      d_arr_add_18_11 : IN std_logic ;
      d_arr_add_18_10 : IN std_logic ;
      d_arr_add_18_9 : IN std_logic ;
      d_arr_add_18_8 : IN std_logic ;
      d_arr_add_18_7 : IN std_logic ;
      d_arr_add_18_6 : IN std_logic ;
      d_arr_add_18_5 : IN std_logic ;
      d_arr_add_18_4 : IN std_logic ;
      d_arr_add_18_3 : IN std_logic ;
      d_arr_add_18_2 : IN std_logic ;
      d_arr_add_18_1 : IN std_logic ;
      d_arr_add_18_0 : IN std_logic ;
      d_arr_add_19_31 : IN std_logic ;
      d_arr_add_19_30 : IN std_logic ;
      d_arr_add_19_29 : IN std_logic ;
      d_arr_add_19_28 : IN std_logic ;
      d_arr_add_19_27 : IN std_logic ;
      d_arr_add_19_26 : IN std_logic ;
      d_arr_add_19_25 : IN std_logic ;
      d_arr_add_19_24 : IN std_logic ;
      d_arr_add_19_23 : IN std_logic ;
      d_arr_add_19_22 : IN std_logic ;
      d_arr_add_19_21 : IN std_logic ;
      d_arr_add_19_20 : IN std_logic ;
      d_arr_add_19_19 : IN std_logic ;
      d_arr_add_19_18 : IN std_logic ;
      d_arr_add_19_17 : IN std_logic ;
      d_arr_add_19_16 : IN std_logic ;
      d_arr_add_19_15 : IN std_logic ;
      d_arr_add_19_14 : IN std_logic ;
      d_arr_add_19_13 : IN std_logic ;
      d_arr_add_19_12 : IN std_logic ;
      d_arr_add_19_11 : IN std_logic ;
      d_arr_add_19_10 : IN std_logic ;
      d_arr_add_19_9 : IN std_logic ;
      d_arr_add_19_8 : IN std_logic ;
      d_arr_add_19_7 : IN std_logic ;
      d_arr_add_19_6 : IN std_logic ;
      d_arr_add_19_5 : IN std_logic ;
      d_arr_add_19_4 : IN std_logic ;
      d_arr_add_19_3 : IN std_logic ;
      d_arr_add_19_2 : IN std_logic ;
      d_arr_add_19_1 : IN std_logic ;
      d_arr_add_19_0 : IN std_logic ;
      d_arr_add_20_31 : IN std_logic ;
      d_arr_add_20_30 : IN std_logic ;
      d_arr_add_20_29 : IN std_logic ;
      d_arr_add_20_28 : IN std_logic ;
      d_arr_add_20_27 : IN std_logic ;
      d_arr_add_20_26 : IN std_logic ;
      d_arr_add_20_25 : IN std_logic ;
      d_arr_add_20_24 : IN std_logic ;
      d_arr_add_20_23 : IN std_logic ;
      d_arr_add_20_22 : IN std_logic ;
      d_arr_add_20_21 : IN std_logic ;
      d_arr_add_20_20 : IN std_logic ;
      d_arr_add_20_19 : IN std_logic ;
      d_arr_add_20_18 : IN std_logic ;
      d_arr_add_20_17 : IN std_logic ;
      d_arr_add_20_16 : IN std_logic ;
      d_arr_add_20_15 : IN std_logic ;
      d_arr_add_20_14 : IN std_logic ;
      d_arr_add_20_13 : IN std_logic ;
      d_arr_add_20_12 : IN std_logic ;
      d_arr_add_20_11 : IN std_logic ;
      d_arr_add_20_10 : IN std_logic ;
      d_arr_add_20_9 : IN std_logic ;
      d_arr_add_20_8 : IN std_logic ;
      d_arr_add_20_7 : IN std_logic ;
      d_arr_add_20_6 : IN std_logic ;
      d_arr_add_20_5 : IN std_logic ;
      d_arr_add_20_4 : IN std_logic ;
      d_arr_add_20_3 : IN std_logic ;
      d_arr_add_20_2 : IN std_logic ;
      d_arr_add_20_1 : IN std_logic ;
      d_arr_add_20_0 : IN std_logic ;
      d_arr_add_21_31 : IN std_logic ;
      d_arr_add_21_30 : IN std_logic ;
      d_arr_add_21_29 : IN std_logic ;
      d_arr_add_21_28 : IN std_logic ;
      d_arr_add_21_27 : IN std_logic ;
      d_arr_add_21_26 : IN std_logic ;
      d_arr_add_21_25 : IN std_logic ;
      d_arr_add_21_24 : IN std_logic ;
      d_arr_add_21_23 : IN std_logic ;
      d_arr_add_21_22 : IN std_logic ;
      d_arr_add_21_21 : IN std_logic ;
      d_arr_add_21_20 : IN std_logic ;
      d_arr_add_21_19 : IN std_logic ;
      d_arr_add_21_18 : IN std_logic ;
      d_arr_add_21_17 : IN std_logic ;
      d_arr_add_21_16 : IN std_logic ;
      d_arr_add_21_15 : IN std_logic ;
      d_arr_add_21_14 : IN std_logic ;
      d_arr_add_21_13 : IN std_logic ;
      d_arr_add_21_12 : IN std_logic ;
      d_arr_add_21_11 : IN std_logic ;
      d_arr_add_21_10 : IN std_logic ;
      d_arr_add_21_9 : IN std_logic ;
      d_arr_add_21_8 : IN std_logic ;
      d_arr_add_21_7 : IN std_logic ;
      d_arr_add_21_6 : IN std_logic ;
      d_arr_add_21_5 : IN std_logic ;
      d_arr_add_21_4 : IN std_logic ;
      d_arr_add_21_3 : IN std_logic ;
      d_arr_add_21_2 : IN std_logic ;
      d_arr_add_21_1 : IN std_logic ;
      d_arr_add_21_0 : IN std_logic ;
      d_arr_add_22_31 : IN std_logic ;
      d_arr_add_22_30 : IN std_logic ;
      d_arr_add_22_29 : IN std_logic ;
      d_arr_add_22_28 : IN std_logic ;
      d_arr_add_22_27 : IN std_logic ;
      d_arr_add_22_26 : IN std_logic ;
      d_arr_add_22_25 : IN std_logic ;
      d_arr_add_22_24 : IN std_logic ;
      d_arr_add_22_23 : IN std_logic ;
      d_arr_add_22_22 : IN std_logic ;
      d_arr_add_22_21 : IN std_logic ;
      d_arr_add_22_20 : IN std_logic ;
      d_arr_add_22_19 : IN std_logic ;
      d_arr_add_22_18 : IN std_logic ;
      d_arr_add_22_17 : IN std_logic ;
      d_arr_add_22_16 : IN std_logic ;
      d_arr_add_22_15 : IN std_logic ;
      d_arr_add_22_14 : IN std_logic ;
      d_arr_add_22_13 : IN std_logic ;
      d_arr_add_22_12 : IN std_logic ;
      d_arr_add_22_11 : IN std_logic ;
      d_arr_add_22_10 : IN std_logic ;
      d_arr_add_22_9 : IN std_logic ;
      d_arr_add_22_8 : IN std_logic ;
      d_arr_add_22_7 : IN std_logic ;
      d_arr_add_22_6 : IN std_logic ;
      d_arr_add_22_5 : IN std_logic ;
      d_arr_add_22_4 : IN std_logic ;
      d_arr_add_22_3 : IN std_logic ;
      d_arr_add_22_2 : IN std_logic ;
      d_arr_add_22_1 : IN std_logic ;
      d_arr_add_22_0 : IN std_logic ;
      d_arr_add_23_31 : IN std_logic ;
      d_arr_add_23_30 : IN std_logic ;
      d_arr_add_23_29 : IN std_logic ;
      d_arr_add_23_28 : IN std_logic ;
      d_arr_add_23_27 : IN std_logic ;
      d_arr_add_23_26 : IN std_logic ;
      d_arr_add_23_25 : IN std_logic ;
      d_arr_add_23_24 : IN std_logic ;
      d_arr_add_23_23 : IN std_logic ;
      d_arr_add_23_22 : IN std_logic ;
      d_arr_add_23_21 : IN std_logic ;
      d_arr_add_23_20 : IN std_logic ;
      d_arr_add_23_19 : IN std_logic ;
      d_arr_add_23_18 : IN std_logic ;
      d_arr_add_23_17 : IN std_logic ;
      d_arr_add_23_16 : IN std_logic ;
      d_arr_add_23_15 : IN std_logic ;
      d_arr_add_23_14 : IN std_logic ;
      d_arr_add_23_13 : IN std_logic ;
      d_arr_add_23_12 : IN std_logic ;
      d_arr_add_23_11 : IN std_logic ;
      d_arr_add_23_10 : IN std_logic ;
      d_arr_add_23_9 : IN std_logic ;
      d_arr_add_23_8 : IN std_logic ;
      d_arr_add_23_7 : IN std_logic ;
      d_arr_add_23_6 : IN std_logic ;
      d_arr_add_23_5 : IN std_logic ;
      d_arr_add_23_4 : IN std_logic ;
      d_arr_add_23_3 : IN std_logic ;
      d_arr_add_23_2 : IN std_logic ;
      d_arr_add_23_1 : IN std_logic ;
      d_arr_add_23_0 : IN std_logic ;
      d_arr_add_24_31 : IN std_logic ;
      d_arr_add_24_30 : IN std_logic ;
      d_arr_add_24_29 : IN std_logic ;
      d_arr_add_24_28 : IN std_logic ;
      d_arr_add_24_27 : IN std_logic ;
      d_arr_add_24_26 : IN std_logic ;
      d_arr_add_24_25 : IN std_logic ;
      d_arr_add_24_24 : IN std_logic ;
      d_arr_add_24_23 : IN std_logic ;
      d_arr_add_24_22 : IN std_logic ;
      d_arr_add_24_21 : IN std_logic ;
      d_arr_add_24_20 : IN std_logic ;
      d_arr_add_24_19 : IN std_logic ;
      d_arr_add_24_18 : IN std_logic ;
      d_arr_add_24_17 : IN std_logic ;
      d_arr_add_24_16 : IN std_logic ;
      d_arr_add_24_15 : IN std_logic ;
      d_arr_add_24_14 : IN std_logic ;
      d_arr_add_24_13 : IN std_logic ;
      d_arr_add_24_12 : IN std_logic ;
      d_arr_add_24_11 : IN std_logic ;
      d_arr_add_24_10 : IN std_logic ;
      d_arr_add_24_9 : IN std_logic ;
      d_arr_add_24_8 : IN std_logic ;
      d_arr_add_24_7 : IN std_logic ;
      d_arr_add_24_6 : IN std_logic ;
      d_arr_add_24_5 : IN std_logic ;
      d_arr_add_24_4 : IN std_logic ;
      d_arr_add_24_3 : IN std_logic ;
      d_arr_add_24_2 : IN std_logic ;
      d_arr_add_24_1 : IN std_logic ;
      d_arr_add_24_0 : IN std_logic ;
      d_arr_merge1_0_31 : IN std_logic ;
      d_arr_merge1_0_30 : IN std_logic ;
      d_arr_merge1_0_29 : IN std_logic ;
      d_arr_merge1_0_28 : IN std_logic ;
      d_arr_merge1_0_27 : IN std_logic ;
      d_arr_merge1_0_26 : IN std_logic ;
      d_arr_merge1_0_25 : IN std_logic ;
      d_arr_merge1_0_24 : IN std_logic ;
      d_arr_merge1_0_23 : IN std_logic ;
      d_arr_merge1_0_22 : IN std_logic ;
      d_arr_merge1_0_21 : IN std_logic ;
      d_arr_merge1_0_20 : IN std_logic ;
      d_arr_merge1_0_19 : IN std_logic ;
      d_arr_merge1_0_18 : IN std_logic ;
      d_arr_merge1_0_17 : IN std_logic ;
      d_arr_merge1_0_16 : IN std_logic ;
      d_arr_merge1_0_15 : IN std_logic ;
      d_arr_merge1_0_14 : IN std_logic ;
      d_arr_merge1_0_13 : IN std_logic ;
      d_arr_merge1_0_12 : IN std_logic ;
      d_arr_merge1_0_11 : IN std_logic ;
      d_arr_merge1_0_10 : IN std_logic ;
      d_arr_merge1_0_9 : IN std_logic ;
      d_arr_merge1_0_8 : IN std_logic ;
      d_arr_merge1_0_7 : IN std_logic ;
      d_arr_merge1_0_6 : IN std_logic ;
      d_arr_merge1_0_5 : IN std_logic ;
      d_arr_merge1_0_4 : IN std_logic ;
      d_arr_merge1_0_3 : IN std_logic ;
      d_arr_merge1_0_2 : IN std_logic ;
      d_arr_merge1_0_1 : IN std_logic ;
      d_arr_merge1_0_0 : IN std_logic ;
      d_arr_merge1_1_31 : IN std_logic ;
      d_arr_merge1_1_30 : IN std_logic ;
      d_arr_merge1_1_29 : IN std_logic ;
      d_arr_merge1_1_28 : IN std_logic ;
      d_arr_merge1_1_27 : IN std_logic ;
      d_arr_merge1_1_26 : IN std_logic ;
      d_arr_merge1_1_25 : IN std_logic ;
      d_arr_merge1_1_24 : IN std_logic ;
      d_arr_merge1_1_23 : IN std_logic ;
      d_arr_merge1_1_22 : IN std_logic ;
      d_arr_merge1_1_21 : IN std_logic ;
      d_arr_merge1_1_20 : IN std_logic ;
      d_arr_merge1_1_19 : IN std_logic ;
      d_arr_merge1_1_18 : IN std_logic ;
      d_arr_merge1_1_17 : IN std_logic ;
      d_arr_merge1_1_16 : IN std_logic ;
      d_arr_merge1_1_15 : IN std_logic ;
      d_arr_merge1_1_14 : IN std_logic ;
      d_arr_merge1_1_13 : IN std_logic ;
      d_arr_merge1_1_12 : IN std_logic ;
      d_arr_merge1_1_11 : IN std_logic ;
      d_arr_merge1_1_10 : IN std_logic ;
      d_arr_merge1_1_9 : IN std_logic ;
      d_arr_merge1_1_8 : IN std_logic ;
      d_arr_merge1_1_7 : IN std_logic ;
      d_arr_merge1_1_6 : IN std_logic ;
      d_arr_merge1_1_5 : IN std_logic ;
      d_arr_merge1_1_4 : IN std_logic ;
      d_arr_merge1_1_3 : IN std_logic ;
      d_arr_merge1_1_2 : IN std_logic ;
      d_arr_merge1_1_1 : IN std_logic ;
      d_arr_merge1_1_0 : IN std_logic ;
      d_arr_merge1_2_31 : IN std_logic ;
      d_arr_merge1_2_30 : IN std_logic ;
      d_arr_merge1_2_29 : IN std_logic ;
      d_arr_merge1_2_28 : IN std_logic ;
      d_arr_merge1_2_27 : IN std_logic ;
      d_arr_merge1_2_26 : IN std_logic ;
      d_arr_merge1_2_25 : IN std_logic ;
      d_arr_merge1_2_24 : IN std_logic ;
      d_arr_merge1_2_23 : IN std_logic ;
      d_arr_merge1_2_22 : IN std_logic ;
      d_arr_merge1_2_21 : IN std_logic ;
      d_arr_merge1_2_20 : IN std_logic ;
      d_arr_merge1_2_19 : IN std_logic ;
      d_arr_merge1_2_18 : IN std_logic ;
      d_arr_merge1_2_17 : IN std_logic ;
      d_arr_merge1_2_16 : IN std_logic ;
      d_arr_merge1_2_15 : IN std_logic ;
      d_arr_merge1_2_14 : IN std_logic ;
      d_arr_merge1_2_13 : IN std_logic ;
      d_arr_merge1_2_12 : IN std_logic ;
      d_arr_merge1_2_11 : IN std_logic ;
      d_arr_merge1_2_10 : IN std_logic ;
      d_arr_merge1_2_9 : IN std_logic ;
      d_arr_merge1_2_8 : IN std_logic ;
      d_arr_merge1_2_7 : IN std_logic ;
      d_arr_merge1_2_6 : IN std_logic ;
      d_arr_merge1_2_5 : IN std_logic ;
      d_arr_merge1_2_4 : IN std_logic ;
      d_arr_merge1_2_3 : IN std_logic ;
      d_arr_merge1_2_2 : IN std_logic ;
      d_arr_merge1_2_1 : IN std_logic ;
      d_arr_merge1_2_0 : IN std_logic ;
      d_arr_merge1_3_31 : IN std_logic ;
      d_arr_merge1_3_30 : IN std_logic ;
      d_arr_merge1_3_29 : IN std_logic ;
      d_arr_merge1_3_28 : IN std_logic ;
      d_arr_merge1_3_27 : IN std_logic ;
      d_arr_merge1_3_26 : IN std_logic ;
      d_arr_merge1_3_25 : IN std_logic ;
      d_arr_merge1_3_24 : IN std_logic ;
      d_arr_merge1_3_23 : IN std_logic ;
      d_arr_merge1_3_22 : IN std_logic ;
      d_arr_merge1_3_21 : IN std_logic ;
      d_arr_merge1_3_20 : IN std_logic ;
      d_arr_merge1_3_19 : IN std_logic ;
      d_arr_merge1_3_18 : IN std_logic ;
      d_arr_merge1_3_17 : IN std_logic ;
      d_arr_merge1_3_16 : IN std_logic ;
      d_arr_merge1_3_15 : IN std_logic ;
      d_arr_merge1_3_14 : IN std_logic ;
      d_arr_merge1_3_13 : IN std_logic ;
      d_arr_merge1_3_12 : IN std_logic ;
      d_arr_merge1_3_11 : IN std_logic ;
      d_arr_merge1_3_10 : IN std_logic ;
      d_arr_merge1_3_9 : IN std_logic ;
      d_arr_merge1_3_8 : IN std_logic ;
      d_arr_merge1_3_7 : IN std_logic ;
      d_arr_merge1_3_6 : IN std_logic ;
      d_arr_merge1_3_5 : IN std_logic ;
      d_arr_merge1_3_4 : IN std_logic ;
      d_arr_merge1_3_3 : IN std_logic ;
      d_arr_merge1_3_2 : IN std_logic ;
      d_arr_merge1_3_1 : IN std_logic ;
      d_arr_merge1_3_0 : IN std_logic ;
      d_arr_merge1_4_31 : IN std_logic ;
      d_arr_merge1_4_30 : IN std_logic ;
      d_arr_merge1_4_29 : IN std_logic ;
      d_arr_merge1_4_28 : IN std_logic ;
      d_arr_merge1_4_27 : IN std_logic ;
      d_arr_merge1_4_26 : IN std_logic ;
      d_arr_merge1_4_25 : IN std_logic ;
      d_arr_merge1_4_24 : IN std_logic ;
      d_arr_merge1_4_23 : IN std_logic ;
      d_arr_merge1_4_22 : IN std_logic ;
      d_arr_merge1_4_21 : IN std_logic ;
      d_arr_merge1_4_20 : IN std_logic ;
      d_arr_merge1_4_19 : IN std_logic ;
      d_arr_merge1_4_18 : IN std_logic ;
      d_arr_merge1_4_17 : IN std_logic ;
      d_arr_merge1_4_16 : IN std_logic ;
      d_arr_merge1_4_15 : IN std_logic ;
      d_arr_merge1_4_14 : IN std_logic ;
      d_arr_merge1_4_13 : IN std_logic ;
      d_arr_merge1_4_12 : IN std_logic ;
      d_arr_merge1_4_11 : IN std_logic ;
      d_arr_merge1_4_10 : IN std_logic ;
      d_arr_merge1_4_9 : IN std_logic ;
      d_arr_merge1_4_8 : IN std_logic ;
      d_arr_merge1_4_7 : IN std_logic ;
      d_arr_merge1_4_6 : IN std_logic ;
      d_arr_merge1_4_5 : IN std_logic ;
      d_arr_merge1_4_4 : IN std_logic ;
      d_arr_merge1_4_3 : IN std_logic ;
      d_arr_merge1_4_2 : IN std_logic ;
      d_arr_merge1_4_1 : IN std_logic ;
      d_arr_merge1_4_0 : IN std_logic ;
      d_arr_merge1_5_31 : IN std_logic ;
      d_arr_merge1_5_30 : IN std_logic ;
      d_arr_merge1_5_29 : IN std_logic ;
      d_arr_merge1_5_28 : IN std_logic ;
      d_arr_merge1_5_27 : IN std_logic ;
      d_arr_merge1_5_26 : IN std_logic ;
      d_arr_merge1_5_25 : IN std_logic ;
      d_arr_merge1_5_24 : IN std_logic ;
      d_arr_merge1_5_23 : IN std_logic ;
      d_arr_merge1_5_22 : IN std_logic ;
      d_arr_merge1_5_21 : IN std_logic ;
      d_arr_merge1_5_20 : IN std_logic ;
      d_arr_merge1_5_19 : IN std_logic ;
      d_arr_merge1_5_18 : IN std_logic ;
      d_arr_merge1_5_17 : IN std_logic ;
      d_arr_merge1_5_16 : IN std_logic ;
      d_arr_merge1_5_15 : IN std_logic ;
      d_arr_merge1_5_14 : IN std_logic ;
      d_arr_merge1_5_13 : IN std_logic ;
      d_arr_merge1_5_12 : IN std_logic ;
      d_arr_merge1_5_11 : IN std_logic ;
      d_arr_merge1_5_10 : IN std_logic ;
      d_arr_merge1_5_9 : IN std_logic ;
      d_arr_merge1_5_8 : IN std_logic ;
      d_arr_merge1_5_7 : IN std_logic ;
      d_arr_merge1_5_6 : IN std_logic ;
      d_arr_merge1_5_5 : IN std_logic ;
      d_arr_merge1_5_4 : IN std_logic ;
      d_arr_merge1_5_3 : IN std_logic ;
      d_arr_merge1_5_2 : IN std_logic ;
      d_arr_merge1_5_1 : IN std_logic ;
      d_arr_merge1_5_0 : IN std_logic ;
      d_arr_merge1_6_31 : IN std_logic ;
      d_arr_merge1_6_30 : IN std_logic ;
      d_arr_merge1_6_29 : IN std_logic ;
      d_arr_merge1_6_28 : IN std_logic ;
      d_arr_merge1_6_27 : IN std_logic ;
      d_arr_merge1_6_26 : IN std_logic ;
      d_arr_merge1_6_25 : IN std_logic ;
      d_arr_merge1_6_24 : IN std_logic ;
      d_arr_merge1_6_23 : IN std_logic ;
      d_arr_merge1_6_22 : IN std_logic ;
      d_arr_merge1_6_21 : IN std_logic ;
      d_arr_merge1_6_20 : IN std_logic ;
      d_arr_merge1_6_19 : IN std_logic ;
      d_arr_merge1_6_18 : IN std_logic ;
      d_arr_merge1_6_17 : IN std_logic ;
      d_arr_merge1_6_16 : IN std_logic ;
      d_arr_merge1_6_15 : IN std_logic ;
      d_arr_merge1_6_14 : IN std_logic ;
      d_arr_merge1_6_13 : IN std_logic ;
      d_arr_merge1_6_12 : IN std_logic ;
      d_arr_merge1_6_11 : IN std_logic ;
      d_arr_merge1_6_10 : IN std_logic ;
      d_arr_merge1_6_9 : IN std_logic ;
      d_arr_merge1_6_8 : IN std_logic ;
      d_arr_merge1_6_7 : IN std_logic ;
      d_arr_merge1_6_6 : IN std_logic ;
      d_arr_merge1_6_5 : IN std_logic ;
      d_arr_merge1_6_4 : IN std_logic ;
      d_arr_merge1_6_3 : IN std_logic ;
      d_arr_merge1_6_2 : IN std_logic ;
      d_arr_merge1_6_1 : IN std_logic ;
      d_arr_merge1_6_0 : IN std_logic ;
      d_arr_merge1_7_31 : IN std_logic ;
      d_arr_merge1_7_30 : IN std_logic ;
      d_arr_merge1_7_29 : IN std_logic ;
      d_arr_merge1_7_28 : IN std_logic ;
      d_arr_merge1_7_27 : IN std_logic ;
      d_arr_merge1_7_26 : IN std_logic ;
      d_arr_merge1_7_25 : IN std_logic ;
      d_arr_merge1_7_24 : IN std_logic ;
      d_arr_merge1_7_23 : IN std_logic ;
      d_arr_merge1_7_22 : IN std_logic ;
      d_arr_merge1_7_21 : IN std_logic ;
      d_arr_merge1_7_20 : IN std_logic ;
      d_arr_merge1_7_19 : IN std_logic ;
      d_arr_merge1_7_18 : IN std_logic ;
      d_arr_merge1_7_17 : IN std_logic ;
      d_arr_merge1_7_16 : IN std_logic ;
      d_arr_merge1_7_15 : IN std_logic ;
      d_arr_merge1_7_14 : IN std_logic ;
      d_arr_merge1_7_13 : IN std_logic ;
      d_arr_merge1_7_12 : IN std_logic ;
      d_arr_merge1_7_11 : IN std_logic ;
      d_arr_merge1_7_10 : IN std_logic ;
      d_arr_merge1_7_9 : IN std_logic ;
      d_arr_merge1_7_8 : IN std_logic ;
      d_arr_merge1_7_7 : IN std_logic ;
      d_arr_merge1_7_6 : IN std_logic ;
      d_arr_merge1_7_5 : IN std_logic ;
      d_arr_merge1_7_4 : IN std_logic ;
      d_arr_merge1_7_3 : IN std_logic ;
      d_arr_merge1_7_2 : IN std_logic ;
      d_arr_merge1_7_1 : IN std_logic ;
      d_arr_merge1_7_0 : IN std_logic ;
      d_arr_merge1_8_31 : IN std_logic ;
      d_arr_merge1_8_30 : IN std_logic ;
      d_arr_merge1_8_29 : IN std_logic ;
      d_arr_merge1_8_28 : IN std_logic ;
      d_arr_merge1_8_27 : IN std_logic ;
      d_arr_merge1_8_26 : IN std_logic ;
      d_arr_merge1_8_25 : IN std_logic ;
      d_arr_merge1_8_24 : IN std_logic ;
      d_arr_merge1_8_23 : IN std_logic ;
      d_arr_merge1_8_22 : IN std_logic ;
      d_arr_merge1_8_21 : IN std_logic ;
      d_arr_merge1_8_20 : IN std_logic ;
      d_arr_merge1_8_19 : IN std_logic ;
      d_arr_merge1_8_18 : IN std_logic ;
      d_arr_merge1_8_17 : IN std_logic ;
      d_arr_merge1_8_16 : IN std_logic ;
      d_arr_merge1_8_15 : IN std_logic ;
      d_arr_merge1_8_14 : IN std_logic ;
      d_arr_merge1_8_13 : IN std_logic ;
      d_arr_merge1_8_12 : IN std_logic ;
      d_arr_merge1_8_11 : IN std_logic ;
      d_arr_merge1_8_10 : IN std_logic ;
      d_arr_merge1_8_9 : IN std_logic ;
      d_arr_merge1_8_8 : IN std_logic ;
      d_arr_merge1_8_7 : IN std_logic ;
      d_arr_merge1_8_6 : IN std_logic ;
      d_arr_merge1_8_5 : IN std_logic ;
      d_arr_merge1_8_4 : IN std_logic ;
      d_arr_merge1_8_3 : IN std_logic ;
      d_arr_merge1_8_2 : IN std_logic ;
      d_arr_merge1_8_1 : IN std_logic ;
      d_arr_merge1_8_0 : IN std_logic ;
      d_arr_merge1_9_31 : IN std_logic ;
      d_arr_merge1_9_30 : IN std_logic ;
      d_arr_merge1_9_29 : IN std_logic ;
      d_arr_merge1_9_28 : IN std_logic ;
      d_arr_merge1_9_27 : IN std_logic ;
      d_arr_merge1_9_26 : IN std_logic ;
      d_arr_merge1_9_25 : IN std_logic ;
      d_arr_merge1_9_24 : IN std_logic ;
      d_arr_merge1_9_23 : IN std_logic ;
      d_arr_merge1_9_22 : IN std_logic ;
      d_arr_merge1_9_21 : IN std_logic ;
      d_arr_merge1_9_20 : IN std_logic ;
      d_arr_merge1_9_19 : IN std_logic ;
      d_arr_merge1_9_18 : IN std_logic ;
      d_arr_merge1_9_17 : IN std_logic ;
      d_arr_merge1_9_16 : IN std_logic ;
      d_arr_merge1_9_15 : IN std_logic ;
      d_arr_merge1_9_14 : IN std_logic ;
      d_arr_merge1_9_13 : IN std_logic ;
      d_arr_merge1_9_12 : IN std_logic ;
      d_arr_merge1_9_11 : IN std_logic ;
      d_arr_merge1_9_10 : IN std_logic ;
      d_arr_merge1_9_9 : IN std_logic ;
      d_arr_merge1_9_8 : IN std_logic ;
      d_arr_merge1_9_7 : IN std_logic ;
      d_arr_merge1_9_6 : IN std_logic ;
      d_arr_merge1_9_5 : IN std_logic ;
      d_arr_merge1_9_4 : IN std_logic ;
      d_arr_merge1_9_3 : IN std_logic ;
      d_arr_merge1_9_2 : IN std_logic ;
      d_arr_merge1_9_1 : IN std_logic ;
      d_arr_merge1_9_0 : IN std_logic ;
      d_arr_merge1_10_31 : IN std_logic ;
      d_arr_merge1_10_30 : IN std_logic ;
      d_arr_merge1_10_29 : IN std_logic ;
      d_arr_merge1_10_28 : IN std_logic ;
      d_arr_merge1_10_27 : IN std_logic ;
      d_arr_merge1_10_26 : IN std_logic ;
      d_arr_merge1_10_25 : IN std_logic ;
      d_arr_merge1_10_24 : IN std_logic ;
      d_arr_merge1_10_23 : IN std_logic ;
      d_arr_merge1_10_22 : IN std_logic ;
      d_arr_merge1_10_21 : IN std_logic ;
      d_arr_merge1_10_20 : IN std_logic ;
      d_arr_merge1_10_19 : IN std_logic ;
      d_arr_merge1_10_18 : IN std_logic ;
      d_arr_merge1_10_17 : IN std_logic ;
      d_arr_merge1_10_16 : IN std_logic ;
      d_arr_merge1_10_15 : IN std_logic ;
      d_arr_merge1_10_14 : IN std_logic ;
      d_arr_merge1_10_13 : IN std_logic ;
      d_arr_merge1_10_12 : IN std_logic ;
      d_arr_merge1_10_11 : IN std_logic ;
      d_arr_merge1_10_10 : IN std_logic ;
      d_arr_merge1_10_9 : IN std_logic ;
      d_arr_merge1_10_8 : IN std_logic ;
      d_arr_merge1_10_7 : IN std_logic ;
      d_arr_merge1_10_6 : IN std_logic ;
      d_arr_merge1_10_5 : IN std_logic ;
      d_arr_merge1_10_4 : IN std_logic ;
      d_arr_merge1_10_3 : IN std_logic ;
      d_arr_merge1_10_2 : IN std_logic ;
      d_arr_merge1_10_1 : IN std_logic ;
      d_arr_merge1_10_0 : IN std_logic ;
      d_arr_merge1_11_31 : IN std_logic ;
      d_arr_merge1_11_30 : IN std_logic ;
      d_arr_merge1_11_29 : IN std_logic ;
      d_arr_merge1_11_28 : IN std_logic ;
      d_arr_merge1_11_27 : IN std_logic ;
      d_arr_merge1_11_26 : IN std_logic ;
      d_arr_merge1_11_25 : IN std_logic ;
      d_arr_merge1_11_24 : IN std_logic ;
      d_arr_merge1_11_23 : IN std_logic ;
      d_arr_merge1_11_22 : IN std_logic ;
      d_arr_merge1_11_21 : IN std_logic ;
      d_arr_merge1_11_20 : IN std_logic ;
      d_arr_merge1_11_19 : IN std_logic ;
      d_arr_merge1_11_18 : IN std_logic ;
      d_arr_merge1_11_17 : IN std_logic ;
      d_arr_merge1_11_16 : IN std_logic ;
      d_arr_merge1_11_15 : IN std_logic ;
      d_arr_merge1_11_14 : IN std_logic ;
      d_arr_merge1_11_13 : IN std_logic ;
      d_arr_merge1_11_12 : IN std_logic ;
      d_arr_merge1_11_11 : IN std_logic ;
      d_arr_merge1_11_10 : IN std_logic ;
      d_arr_merge1_11_9 : IN std_logic ;
      d_arr_merge1_11_8 : IN std_logic ;
      d_arr_merge1_11_7 : IN std_logic ;
      d_arr_merge1_11_6 : IN std_logic ;
      d_arr_merge1_11_5 : IN std_logic ;
      d_arr_merge1_11_4 : IN std_logic ;
      d_arr_merge1_11_3 : IN std_logic ;
      d_arr_merge1_11_2 : IN std_logic ;
      d_arr_merge1_11_1 : IN std_logic ;
      d_arr_merge1_11_0 : IN std_logic ;
      d_arr_merge1_12_31 : IN std_logic ;
      d_arr_merge1_12_30 : IN std_logic ;
      d_arr_merge1_12_29 : IN std_logic ;
      d_arr_merge1_12_28 : IN std_logic ;
      d_arr_merge1_12_27 : IN std_logic ;
      d_arr_merge1_12_26 : IN std_logic ;
      d_arr_merge1_12_25 : IN std_logic ;
      d_arr_merge1_12_24 : IN std_logic ;
      d_arr_merge1_12_23 : IN std_logic ;
      d_arr_merge1_12_22 : IN std_logic ;
      d_arr_merge1_12_21 : IN std_logic ;
      d_arr_merge1_12_20 : IN std_logic ;
      d_arr_merge1_12_19 : IN std_logic ;
      d_arr_merge1_12_18 : IN std_logic ;
      d_arr_merge1_12_17 : IN std_logic ;
      d_arr_merge1_12_16 : IN std_logic ;
      d_arr_merge1_12_15 : IN std_logic ;
      d_arr_merge1_12_14 : IN std_logic ;
      d_arr_merge1_12_13 : IN std_logic ;
      d_arr_merge1_12_12 : IN std_logic ;
      d_arr_merge1_12_11 : IN std_logic ;
      d_arr_merge1_12_10 : IN std_logic ;
      d_arr_merge1_12_9 : IN std_logic ;
      d_arr_merge1_12_8 : IN std_logic ;
      d_arr_merge1_12_7 : IN std_logic ;
      d_arr_merge1_12_6 : IN std_logic ;
      d_arr_merge1_12_5 : IN std_logic ;
      d_arr_merge1_12_4 : IN std_logic ;
      d_arr_merge1_12_3 : IN std_logic ;
      d_arr_merge1_12_2 : IN std_logic ;
      d_arr_merge1_12_1 : IN std_logic ;
      d_arr_merge1_12_0 : IN std_logic ;
      d_arr_merge1_13_31 : IN std_logic ;
      d_arr_merge1_13_30 : IN std_logic ;
      d_arr_merge1_13_29 : IN std_logic ;
      d_arr_merge1_13_28 : IN std_logic ;
      d_arr_merge1_13_27 : IN std_logic ;
      d_arr_merge1_13_26 : IN std_logic ;
      d_arr_merge1_13_25 : IN std_logic ;
      d_arr_merge1_13_24 : IN std_logic ;
      d_arr_merge1_13_23 : IN std_logic ;
      d_arr_merge1_13_22 : IN std_logic ;
      d_arr_merge1_13_21 : IN std_logic ;
      d_arr_merge1_13_20 : IN std_logic ;
      d_arr_merge1_13_19 : IN std_logic ;
      d_arr_merge1_13_18 : IN std_logic ;
      d_arr_merge1_13_17 : IN std_logic ;
      d_arr_merge1_13_16 : IN std_logic ;
      d_arr_merge1_13_15 : IN std_logic ;
      d_arr_merge1_13_14 : IN std_logic ;
      d_arr_merge1_13_13 : IN std_logic ;
      d_arr_merge1_13_12 : IN std_logic ;
      d_arr_merge1_13_11 : IN std_logic ;
      d_arr_merge1_13_10 : IN std_logic ;
      d_arr_merge1_13_9 : IN std_logic ;
      d_arr_merge1_13_8 : IN std_logic ;
      d_arr_merge1_13_7 : IN std_logic ;
      d_arr_merge1_13_6 : IN std_logic ;
      d_arr_merge1_13_5 : IN std_logic ;
      d_arr_merge1_13_4 : IN std_logic ;
      d_arr_merge1_13_3 : IN std_logic ;
      d_arr_merge1_13_2 : IN std_logic ;
      d_arr_merge1_13_1 : IN std_logic ;
      d_arr_merge1_13_0 : IN std_logic ;
      d_arr_merge1_14_31 : IN std_logic ;
      d_arr_merge1_14_30 : IN std_logic ;
      d_arr_merge1_14_29 : IN std_logic ;
      d_arr_merge1_14_28 : IN std_logic ;
      d_arr_merge1_14_27 : IN std_logic ;
      d_arr_merge1_14_26 : IN std_logic ;
      d_arr_merge1_14_25 : IN std_logic ;
      d_arr_merge1_14_24 : IN std_logic ;
      d_arr_merge1_14_23 : IN std_logic ;
      d_arr_merge1_14_22 : IN std_logic ;
      d_arr_merge1_14_21 : IN std_logic ;
      d_arr_merge1_14_20 : IN std_logic ;
      d_arr_merge1_14_19 : IN std_logic ;
      d_arr_merge1_14_18 : IN std_logic ;
      d_arr_merge1_14_17 : IN std_logic ;
      d_arr_merge1_14_16 : IN std_logic ;
      d_arr_merge1_14_15 : IN std_logic ;
      d_arr_merge1_14_14 : IN std_logic ;
      d_arr_merge1_14_13 : IN std_logic ;
      d_arr_merge1_14_12 : IN std_logic ;
      d_arr_merge1_14_11 : IN std_logic ;
      d_arr_merge1_14_10 : IN std_logic ;
      d_arr_merge1_14_9 : IN std_logic ;
      d_arr_merge1_14_8 : IN std_logic ;
      d_arr_merge1_14_7 : IN std_logic ;
      d_arr_merge1_14_6 : IN std_logic ;
      d_arr_merge1_14_5 : IN std_logic ;
      d_arr_merge1_14_4 : IN std_logic ;
      d_arr_merge1_14_3 : IN std_logic ;
      d_arr_merge1_14_2 : IN std_logic ;
      d_arr_merge1_14_1 : IN std_logic ;
      d_arr_merge1_14_0 : IN std_logic ;
      d_arr_merge1_15_31 : IN std_logic ;
      d_arr_merge1_15_30 : IN std_logic ;
      d_arr_merge1_15_29 : IN std_logic ;
      d_arr_merge1_15_28 : IN std_logic ;
      d_arr_merge1_15_27 : IN std_logic ;
      d_arr_merge1_15_26 : IN std_logic ;
      d_arr_merge1_15_25 : IN std_logic ;
      d_arr_merge1_15_24 : IN std_logic ;
      d_arr_merge1_15_23 : IN std_logic ;
      d_arr_merge1_15_22 : IN std_logic ;
      d_arr_merge1_15_21 : IN std_logic ;
      d_arr_merge1_15_20 : IN std_logic ;
      d_arr_merge1_15_19 : IN std_logic ;
      d_arr_merge1_15_18 : IN std_logic ;
      d_arr_merge1_15_17 : IN std_logic ;
      d_arr_merge1_15_16 : IN std_logic ;
      d_arr_merge1_15_15 : IN std_logic ;
      d_arr_merge1_15_14 : IN std_logic ;
      d_arr_merge1_15_13 : IN std_logic ;
      d_arr_merge1_15_12 : IN std_logic ;
      d_arr_merge1_15_11 : IN std_logic ;
      d_arr_merge1_15_10 : IN std_logic ;
      d_arr_merge1_15_9 : IN std_logic ;
      d_arr_merge1_15_8 : IN std_logic ;
      d_arr_merge1_15_7 : IN std_logic ;
      d_arr_merge1_15_6 : IN std_logic ;
      d_arr_merge1_15_5 : IN std_logic ;
      d_arr_merge1_15_4 : IN std_logic ;
      d_arr_merge1_15_3 : IN std_logic ;
      d_arr_merge1_15_2 : IN std_logic ;
      d_arr_merge1_15_1 : IN std_logic ;
      d_arr_merge1_15_0 : IN std_logic ;
      d_arr_merge1_16_31 : IN std_logic ;
      d_arr_merge1_16_30 : IN std_logic ;
      d_arr_merge1_16_29 : IN std_logic ;
      d_arr_merge1_16_28 : IN std_logic ;
      d_arr_merge1_16_27 : IN std_logic ;
      d_arr_merge1_16_26 : IN std_logic ;
      d_arr_merge1_16_25 : IN std_logic ;
      d_arr_merge1_16_24 : IN std_logic ;
      d_arr_merge1_16_23 : IN std_logic ;
      d_arr_merge1_16_22 : IN std_logic ;
      d_arr_merge1_16_21 : IN std_logic ;
      d_arr_merge1_16_20 : IN std_logic ;
      d_arr_merge1_16_19 : IN std_logic ;
      d_arr_merge1_16_18 : IN std_logic ;
      d_arr_merge1_16_17 : IN std_logic ;
      d_arr_merge1_16_16 : IN std_logic ;
      d_arr_merge1_16_15 : IN std_logic ;
      d_arr_merge1_16_14 : IN std_logic ;
      d_arr_merge1_16_13 : IN std_logic ;
      d_arr_merge1_16_12 : IN std_logic ;
      d_arr_merge1_16_11 : IN std_logic ;
      d_arr_merge1_16_10 : IN std_logic ;
      d_arr_merge1_16_9 : IN std_logic ;
      d_arr_merge1_16_8 : IN std_logic ;
      d_arr_merge1_16_7 : IN std_logic ;
      d_arr_merge1_16_6 : IN std_logic ;
      d_arr_merge1_16_5 : IN std_logic ;
      d_arr_merge1_16_4 : IN std_logic ;
      d_arr_merge1_16_3 : IN std_logic ;
      d_arr_merge1_16_2 : IN std_logic ;
      d_arr_merge1_16_1 : IN std_logic ;
      d_arr_merge1_16_0 : IN std_logic ;
      d_arr_merge1_17_31 : IN std_logic ;
      d_arr_merge1_17_30 : IN std_logic ;
      d_arr_merge1_17_29 : IN std_logic ;
      d_arr_merge1_17_28 : IN std_logic ;
      d_arr_merge1_17_27 : IN std_logic ;
      d_arr_merge1_17_26 : IN std_logic ;
      d_arr_merge1_17_25 : IN std_logic ;
      d_arr_merge1_17_24 : IN std_logic ;
      d_arr_merge1_17_23 : IN std_logic ;
      d_arr_merge1_17_22 : IN std_logic ;
      d_arr_merge1_17_21 : IN std_logic ;
      d_arr_merge1_17_20 : IN std_logic ;
      d_arr_merge1_17_19 : IN std_logic ;
      d_arr_merge1_17_18 : IN std_logic ;
      d_arr_merge1_17_17 : IN std_logic ;
      d_arr_merge1_17_16 : IN std_logic ;
      d_arr_merge1_17_15 : IN std_logic ;
      d_arr_merge1_17_14 : IN std_logic ;
      d_arr_merge1_17_13 : IN std_logic ;
      d_arr_merge1_17_12 : IN std_logic ;
      d_arr_merge1_17_11 : IN std_logic ;
      d_arr_merge1_17_10 : IN std_logic ;
      d_arr_merge1_17_9 : IN std_logic ;
      d_arr_merge1_17_8 : IN std_logic ;
      d_arr_merge1_17_7 : IN std_logic ;
      d_arr_merge1_17_6 : IN std_logic ;
      d_arr_merge1_17_5 : IN std_logic ;
      d_arr_merge1_17_4 : IN std_logic ;
      d_arr_merge1_17_3 : IN std_logic ;
      d_arr_merge1_17_2 : IN std_logic ;
      d_arr_merge1_17_1 : IN std_logic ;
      d_arr_merge1_17_0 : IN std_logic ;
      d_arr_merge1_18_31 : IN std_logic ;
      d_arr_merge1_18_30 : IN std_logic ;
      d_arr_merge1_18_29 : IN std_logic ;
      d_arr_merge1_18_28 : IN std_logic ;
      d_arr_merge1_18_27 : IN std_logic ;
      d_arr_merge1_18_26 : IN std_logic ;
      d_arr_merge1_18_25 : IN std_logic ;
      d_arr_merge1_18_24 : IN std_logic ;
      d_arr_merge1_18_23 : IN std_logic ;
      d_arr_merge1_18_22 : IN std_logic ;
      d_arr_merge1_18_21 : IN std_logic ;
      d_arr_merge1_18_20 : IN std_logic ;
      d_arr_merge1_18_19 : IN std_logic ;
      d_arr_merge1_18_18 : IN std_logic ;
      d_arr_merge1_18_17 : IN std_logic ;
      d_arr_merge1_18_16 : IN std_logic ;
      d_arr_merge1_18_15 : IN std_logic ;
      d_arr_merge1_18_14 : IN std_logic ;
      d_arr_merge1_18_13 : IN std_logic ;
      d_arr_merge1_18_12 : IN std_logic ;
      d_arr_merge1_18_11 : IN std_logic ;
      d_arr_merge1_18_10 : IN std_logic ;
      d_arr_merge1_18_9 : IN std_logic ;
      d_arr_merge1_18_8 : IN std_logic ;
      d_arr_merge1_18_7 : IN std_logic ;
      d_arr_merge1_18_6 : IN std_logic ;
      d_arr_merge1_18_5 : IN std_logic ;
      d_arr_merge1_18_4 : IN std_logic ;
      d_arr_merge1_18_3 : IN std_logic ;
      d_arr_merge1_18_2 : IN std_logic ;
      d_arr_merge1_18_1 : IN std_logic ;
      d_arr_merge1_18_0 : IN std_logic ;
      d_arr_merge1_19_31 : IN std_logic ;
      d_arr_merge1_19_30 : IN std_logic ;
      d_arr_merge1_19_29 : IN std_logic ;
      d_arr_merge1_19_28 : IN std_logic ;
      d_arr_merge1_19_27 : IN std_logic ;
      d_arr_merge1_19_26 : IN std_logic ;
      d_arr_merge1_19_25 : IN std_logic ;
      d_arr_merge1_19_24 : IN std_logic ;
      d_arr_merge1_19_23 : IN std_logic ;
      d_arr_merge1_19_22 : IN std_logic ;
      d_arr_merge1_19_21 : IN std_logic ;
      d_arr_merge1_19_20 : IN std_logic ;
      d_arr_merge1_19_19 : IN std_logic ;
      d_arr_merge1_19_18 : IN std_logic ;
      d_arr_merge1_19_17 : IN std_logic ;
      d_arr_merge1_19_16 : IN std_logic ;
      d_arr_merge1_19_15 : IN std_logic ;
      d_arr_merge1_19_14 : IN std_logic ;
      d_arr_merge1_19_13 : IN std_logic ;
      d_arr_merge1_19_12 : IN std_logic ;
      d_arr_merge1_19_11 : IN std_logic ;
      d_arr_merge1_19_10 : IN std_logic ;
      d_arr_merge1_19_9 : IN std_logic ;
      d_arr_merge1_19_8 : IN std_logic ;
      d_arr_merge1_19_7 : IN std_logic ;
      d_arr_merge1_19_6 : IN std_logic ;
      d_arr_merge1_19_5 : IN std_logic ;
      d_arr_merge1_19_4 : IN std_logic ;
      d_arr_merge1_19_3 : IN std_logic ;
      d_arr_merge1_19_2 : IN std_logic ;
      d_arr_merge1_19_1 : IN std_logic ;
      d_arr_merge1_19_0 : IN std_logic ;
      d_arr_merge1_20_31 : IN std_logic ;
      d_arr_merge1_20_30 : IN std_logic ;
      d_arr_merge1_20_29 : IN std_logic ;
      d_arr_merge1_20_28 : IN std_logic ;
      d_arr_merge1_20_27 : IN std_logic ;
      d_arr_merge1_20_26 : IN std_logic ;
      d_arr_merge1_20_25 : IN std_logic ;
      d_arr_merge1_20_24 : IN std_logic ;
      d_arr_merge1_20_23 : IN std_logic ;
      d_arr_merge1_20_22 : IN std_logic ;
      d_arr_merge1_20_21 : IN std_logic ;
      d_arr_merge1_20_20 : IN std_logic ;
      d_arr_merge1_20_19 : IN std_logic ;
      d_arr_merge1_20_18 : IN std_logic ;
      d_arr_merge1_20_17 : IN std_logic ;
      d_arr_merge1_20_16 : IN std_logic ;
      d_arr_merge1_20_15 : IN std_logic ;
      d_arr_merge1_20_14 : IN std_logic ;
      d_arr_merge1_20_13 : IN std_logic ;
      d_arr_merge1_20_12 : IN std_logic ;
      d_arr_merge1_20_11 : IN std_logic ;
      d_arr_merge1_20_10 : IN std_logic ;
      d_arr_merge1_20_9 : IN std_logic ;
      d_arr_merge1_20_8 : IN std_logic ;
      d_arr_merge1_20_7 : IN std_logic ;
      d_arr_merge1_20_6 : IN std_logic ;
      d_arr_merge1_20_5 : IN std_logic ;
      d_arr_merge1_20_4 : IN std_logic ;
      d_arr_merge1_20_3 : IN std_logic ;
      d_arr_merge1_20_2 : IN std_logic ;
      d_arr_merge1_20_1 : IN std_logic ;
      d_arr_merge1_20_0 : IN std_logic ;
      d_arr_merge1_21_31 : IN std_logic ;
      d_arr_merge1_21_30 : IN std_logic ;
      d_arr_merge1_21_29 : IN std_logic ;
      d_arr_merge1_21_28 : IN std_logic ;
      d_arr_merge1_21_27 : IN std_logic ;
      d_arr_merge1_21_26 : IN std_logic ;
      d_arr_merge1_21_25 : IN std_logic ;
      d_arr_merge1_21_24 : IN std_logic ;
      d_arr_merge1_21_23 : IN std_logic ;
      d_arr_merge1_21_22 : IN std_logic ;
      d_arr_merge1_21_21 : IN std_logic ;
      d_arr_merge1_21_20 : IN std_logic ;
      d_arr_merge1_21_19 : IN std_logic ;
      d_arr_merge1_21_18 : IN std_logic ;
      d_arr_merge1_21_17 : IN std_logic ;
      d_arr_merge1_21_16 : IN std_logic ;
      d_arr_merge1_21_15 : IN std_logic ;
      d_arr_merge1_21_14 : IN std_logic ;
      d_arr_merge1_21_13 : IN std_logic ;
      d_arr_merge1_21_12 : IN std_logic ;
      d_arr_merge1_21_11 : IN std_logic ;
      d_arr_merge1_21_10 : IN std_logic ;
      d_arr_merge1_21_9 : IN std_logic ;
      d_arr_merge1_21_8 : IN std_logic ;
      d_arr_merge1_21_7 : IN std_logic ;
      d_arr_merge1_21_6 : IN std_logic ;
      d_arr_merge1_21_5 : IN std_logic ;
      d_arr_merge1_21_4 : IN std_logic ;
      d_arr_merge1_21_3 : IN std_logic ;
      d_arr_merge1_21_2 : IN std_logic ;
      d_arr_merge1_21_1 : IN std_logic ;
      d_arr_merge1_21_0 : IN std_logic ;
      d_arr_merge1_22_31 : IN std_logic ;
      d_arr_merge1_22_30 : IN std_logic ;
      d_arr_merge1_22_29 : IN std_logic ;
      d_arr_merge1_22_28 : IN std_logic ;
      d_arr_merge1_22_27 : IN std_logic ;
      d_arr_merge1_22_26 : IN std_logic ;
      d_arr_merge1_22_25 : IN std_logic ;
      d_arr_merge1_22_24 : IN std_logic ;
      d_arr_merge1_22_23 : IN std_logic ;
      d_arr_merge1_22_22 : IN std_logic ;
      d_arr_merge1_22_21 : IN std_logic ;
      d_arr_merge1_22_20 : IN std_logic ;
      d_arr_merge1_22_19 : IN std_logic ;
      d_arr_merge1_22_18 : IN std_logic ;
      d_arr_merge1_22_17 : IN std_logic ;
      d_arr_merge1_22_16 : IN std_logic ;
      d_arr_merge1_22_15 : IN std_logic ;
      d_arr_merge1_22_14 : IN std_logic ;
      d_arr_merge1_22_13 : IN std_logic ;
      d_arr_merge1_22_12 : IN std_logic ;
      d_arr_merge1_22_11 : IN std_logic ;
      d_arr_merge1_22_10 : IN std_logic ;
      d_arr_merge1_22_9 : IN std_logic ;
      d_arr_merge1_22_8 : IN std_logic ;
      d_arr_merge1_22_7 : IN std_logic ;
      d_arr_merge1_22_6 : IN std_logic ;
      d_arr_merge1_22_5 : IN std_logic ;
      d_arr_merge1_22_4 : IN std_logic ;
      d_arr_merge1_22_3 : IN std_logic ;
      d_arr_merge1_22_2 : IN std_logic ;
      d_arr_merge1_22_1 : IN std_logic ;
      d_arr_merge1_22_0 : IN std_logic ;
      d_arr_merge1_23_31 : IN std_logic ;
      d_arr_merge1_23_30 : IN std_logic ;
      d_arr_merge1_23_29 : IN std_logic ;
      d_arr_merge1_23_28 : IN std_logic ;
      d_arr_merge1_23_27 : IN std_logic ;
      d_arr_merge1_23_26 : IN std_logic ;
      d_arr_merge1_23_25 : IN std_logic ;
      d_arr_merge1_23_24 : IN std_logic ;
      d_arr_merge1_23_23 : IN std_logic ;
      d_arr_merge1_23_22 : IN std_logic ;
      d_arr_merge1_23_21 : IN std_logic ;
      d_arr_merge1_23_20 : IN std_logic ;
      d_arr_merge1_23_19 : IN std_logic ;
      d_arr_merge1_23_18 : IN std_logic ;
      d_arr_merge1_23_17 : IN std_logic ;
      d_arr_merge1_23_16 : IN std_logic ;
      d_arr_merge1_23_15 : IN std_logic ;
      d_arr_merge1_23_14 : IN std_logic ;
      d_arr_merge1_23_13 : IN std_logic ;
      d_arr_merge1_23_12 : IN std_logic ;
      d_arr_merge1_23_11 : IN std_logic ;
      d_arr_merge1_23_10 : IN std_logic ;
      d_arr_merge1_23_9 : IN std_logic ;
      d_arr_merge1_23_8 : IN std_logic ;
      d_arr_merge1_23_7 : IN std_logic ;
      d_arr_merge1_23_6 : IN std_logic ;
      d_arr_merge1_23_5 : IN std_logic ;
      d_arr_merge1_23_4 : IN std_logic ;
      d_arr_merge1_23_3 : IN std_logic ;
      d_arr_merge1_23_2 : IN std_logic ;
      d_arr_merge1_23_1 : IN std_logic ;
      d_arr_merge1_23_0 : IN std_logic ;
      d_arr_merge1_24_31 : IN std_logic ;
      d_arr_merge1_24_30 : IN std_logic ;
      d_arr_merge1_24_29 : IN std_logic ;
      d_arr_merge1_24_28 : IN std_logic ;
      d_arr_merge1_24_27 : IN std_logic ;
      d_arr_merge1_24_26 : IN std_logic ;
      d_arr_merge1_24_25 : IN std_logic ;
      d_arr_merge1_24_24 : IN std_logic ;
      d_arr_merge1_24_23 : IN std_logic ;
      d_arr_merge1_24_22 : IN std_logic ;
      d_arr_merge1_24_21 : IN std_logic ;
      d_arr_merge1_24_20 : IN std_logic ;
      d_arr_merge1_24_19 : IN std_logic ;
      d_arr_merge1_24_18 : IN std_logic ;
      d_arr_merge1_24_17 : IN std_logic ;
      d_arr_merge1_24_16 : IN std_logic ;
      d_arr_merge1_24_15 : IN std_logic ;
      d_arr_merge1_24_14 : IN std_logic ;
      d_arr_merge1_24_13 : IN std_logic ;
      d_arr_merge1_24_12 : IN std_logic ;
      d_arr_merge1_24_11 : IN std_logic ;
      d_arr_merge1_24_10 : IN std_logic ;
      d_arr_merge1_24_9 : IN std_logic ;
      d_arr_merge1_24_8 : IN std_logic ;
      d_arr_merge1_24_7 : IN std_logic ;
      d_arr_merge1_24_6 : IN std_logic ;
      d_arr_merge1_24_5 : IN std_logic ;
      d_arr_merge1_24_4 : IN std_logic ;
      d_arr_merge1_24_3 : IN std_logic ;
      d_arr_merge1_24_2 : IN std_logic ;
      d_arr_merge1_24_1 : IN std_logic ;
      d_arr_merge1_24_0 : IN std_logic ;
      d_arr_merge2_0_31 : IN std_logic ;
      d_arr_merge2_0_30 : IN std_logic ;
      d_arr_merge2_0_29 : IN std_logic ;
      d_arr_merge2_0_28 : IN std_logic ;
      d_arr_merge2_0_27 : IN std_logic ;
      d_arr_merge2_0_26 : IN std_logic ;
      d_arr_merge2_0_25 : IN std_logic ;
      d_arr_merge2_0_24 : IN std_logic ;
      d_arr_merge2_0_23 : IN std_logic ;
      d_arr_merge2_0_22 : IN std_logic ;
      d_arr_merge2_0_21 : IN std_logic ;
      d_arr_merge2_0_20 : IN std_logic ;
      d_arr_merge2_0_19 : IN std_logic ;
      d_arr_merge2_0_18 : IN std_logic ;
      d_arr_merge2_0_17 : IN std_logic ;
      d_arr_merge2_0_16 : IN std_logic ;
      d_arr_merge2_0_15 : IN std_logic ;
      d_arr_merge2_0_14 : IN std_logic ;
      d_arr_merge2_0_13 : IN std_logic ;
      d_arr_merge2_0_12 : IN std_logic ;
      d_arr_merge2_0_11 : IN std_logic ;
      d_arr_merge2_0_10 : IN std_logic ;
      d_arr_merge2_0_9 : IN std_logic ;
      d_arr_merge2_0_8 : IN std_logic ;
      d_arr_merge2_0_7 : IN std_logic ;
      d_arr_merge2_0_6 : IN std_logic ;
      d_arr_merge2_0_5 : IN std_logic ;
      d_arr_merge2_0_4 : IN std_logic ;
      d_arr_merge2_0_3 : IN std_logic ;
      d_arr_merge2_0_2 : IN std_logic ;
      d_arr_merge2_0_1 : IN std_logic ;
      d_arr_merge2_0_0 : IN std_logic ;
      d_arr_merge2_1_31 : IN std_logic ;
      d_arr_merge2_1_30 : IN std_logic ;
      d_arr_merge2_1_29 : IN std_logic ;
      d_arr_merge2_1_28 : IN std_logic ;
      d_arr_merge2_1_27 : IN std_logic ;
      d_arr_merge2_1_26 : IN std_logic ;
      d_arr_merge2_1_25 : IN std_logic ;
      d_arr_merge2_1_24 : IN std_logic ;
      d_arr_merge2_1_23 : IN std_logic ;
      d_arr_merge2_1_22 : IN std_logic ;
      d_arr_merge2_1_21 : IN std_logic ;
      d_arr_merge2_1_20 : IN std_logic ;
      d_arr_merge2_1_19 : IN std_logic ;
      d_arr_merge2_1_18 : IN std_logic ;
      d_arr_merge2_1_17 : IN std_logic ;
      d_arr_merge2_1_16 : IN std_logic ;
      d_arr_merge2_1_15 : IN std_logic ;
      d_arr_merge2_1_14 : IN std_logic ;
      d_arr_merge2_1_13 : IN std_logic ;
      d_arr_merge2_1_12 : IN std_logic ;
      d_arr_merge2_1_11 : IN std_logic ;
      d_arr_merge2_1_10 : IN std_logic ;
      d_arr_merge2_1_9 : IN std_logic ;
      d_arr_merge2_1_8 : IN std_logic ;
      d_arr_merge2_1_7 : IN std_logic ;
      d_arr_merge2_1_6 : IN std_logic ;
      d_arr_merge2_1_5 : IN std_logic ;
      d_arr_merge2_1_4 : IN std_logic ;
      d_arr_merge2_1_3 : IN std_logic ;
      d_arr_merge2_1_2 : IN std_logic ;
      d_arr_merge2_1_1 : IN std_logic ;
      d_arr_merge2_1_0 : IN std_logic ;
      d_arr_merge2_2_31 : IN std_logic ;
      d_arr_merge2_2_30 : IN std_logic ;
      d_arr_merge2_2_29 : IN std_logic ;
      d_arr_merge2_2_28 : IN std_logic ;
      d_arr_merge2_2_27 : IN std_logic ;
      d_arr_merge2_2_26 : IN std_logic ;
      d_arr_merge2_2_25 : IN std_logic ;
      d_arr_merge2_2_24 : IN std_logic ;
      d_arr_merge2_2_23 : IN std_logic ;
      d_arr_merge2_2_22 : IN std_logic ;
      d_arr_merge2_2_21 : IN std_logic ;
      d_arr_merge2_2_20 : IN std_logic ;
      d_arr_merge2_2_19 : IN std_logic ;
      d_arr_merge2_2_18 : IN std_logic ;
      d_arr_merge2_2_17 : IN std_logic ;
      d_arr_merge2_2_16 : IN std_logic ;
      d_arr_merge2_2_15 : IN std_logic ;
      d_arr_merge2_2_14 : IN std_logic ;
      d_arr_merge2_2_13 : IN std_logic ;
      d_arr_merge2_2_12 : IN std_logic ;
      d_arr_merge2_2_11 : IN std_logic ;
      d_arr_merge2_2_10 : IN std_logic ;
      d_arr_merge2_2_9 : IN std_logic ;
      d_arr_merge2_2_8 : IN std_logic ;
      d_arr_merge2_2_7 : IN std_logic ;
      d_arr_merge2_2_6 : IN std_logic ;
      d_arr_merge2_2_5 : IN std_logic ;
      d_arr_merge2_2_4 : IN std_logic ;
      d_arr_merge2_2_3 : IN std_logic ;
      d_arr_merge2_2_2 : IN std_logic ;
      d_arr_merge2_2_1 : IN std_logic ;
      d_arr_merge2_2_0 : IN std_logic ;
      d_arr_merge2_3_31 : IN std_logic ;
      d_arr_merge2_3_30 : IN std_logic ;
      d_arr_merge2_3_29 : IN std_logic ;
      d_arr_merge2_3_28 : IN std_logic ;
      d_arr_merge2_3_27 : IN std_logic ;
      d_arr_merge2_3_26 : IN std_logic ;
      d_arr_merge2_3_25 : IN std_logic ;
      d_arr_merge2_3_24 : IN std_logic ;
      d_arr_merge2_3_23 : IN std_logic ;
      d_arr_merge2_3_22 : IN std_logic ;
      d_arr_merge2_3_21 : IN std_logic ;
      d_arr_merge2_3_20 : IN std_logic ;
      d_arr_merge2_3_19 : IN std_logic ;
      d_arr_merge2_3_18 : IN std_logic ;
      d_arr_merge2_3_17 : IN std_logic ;
      d_arr_merge2_3_16 : IN std_logic ;
      d_arr_merge2_3_15 : IN std_logic ;
      d_arr_merge2_3_14 : IN std_logic ;
      d_arr_merge2_3_13 : IN std_logic ;
      d_arr_merge2_3_12 : IN std_logic ;
      d_arr_merge2_3_11 : IN std_logic ;
      d_arr_merge2_3_10 : IN std_logic ;
      d_arr_merge2_3_9 : IN std_logic ;
      d_arr_merge2_3_8 : IN std_logic ;
      d_arr_merge2_3_7 : IN std_logic ;
      d_arr_merge2_3_6 : IN std_logic ;
      d_arr_merge2_3_5 : IN std_logic ;
      d_arr_merge2_3_4 : IN std_logic ;
      d_arr_merge2_3_3 : IN std_logic ;
      d_arr_merge2_3_2 : IN std_logic ;
      d_arr_merge2_3_1 : IN std_logic ;
      d_arr_merge2_3_0 : IN std_logic ;
      d_arr_merge2_4_31 : IN std_logic ;
      d_arr_merge2_4_30 : IN std_logic ;
      d_arr_merge2_4_29 : IN std_logic ;
      d_arr_merge2_4_28 : IN std_logic ;
      d_arr_merge2_4_27 : IN std_logic ;
      d_arr_merge2_4_26 : IN std_logic ;
      d_arr_merge2_4_25 : IN std_logic ;
      d_arr_merge2_4_24 : IN std_logic ;
      d_arr_merge2_4_23 : IN std_logic ;
      d_arr_merge2_4_22 : IN std_logic ;
      d_arr_merge2_4_21 : IN std_logic ;
      d_arr_merge2_4_20 : IN std_logic ;
      d_arr_merge2_4_19 : IN std_logic ;
      d_arr_merge2_4_18 : IN std_logic ;
      d_arr_merge2_4_17 : IN std_logic ;
      d_arr_merge2_4_16 : IN std_logic ;
      d_arr_merge2_4_15 : IN std_logic ;
      d_arr_merge2_4_14 : IN std_logic ;
      d_arr_merge2_4_13 : IN std_logic ;
      d_arr_merge2_4_12 : IN std_logic ;
      d_arr_merge2_4_11 : IN std_logic ;
      d_arr_merge2_4_10 : IN std_logic ;
      d_arr_merge2_4_9 : IN std_logic ;
      d_arr_merge2_4_8 : IN std_logic ;
      d_arr_merge2_4_7 : IN std_logic ;
      d_arr_merge2_4_6 : IN std_logic ;
      d_arr_merge2_4_5 : IN std_logic ;
      d_arr_merge2_4_4 : IN std_logic ;
      d_arr_merge2_4_3 : IN std_logic ;
      d_arr_merge2_4_2 : IN std_logic ;
      d_arr_merge2_4_1 : IN std_logic ;
      d_arr_merge2_4_0 : IN std_logic ;
      d_arr_merge2_5_31 : IN std_logic ;
      d_arr_merge2_5_30 : IN std_logic ;
      d_arr_merge2_5_29 : IN std_logic ;
      d_arr_merge2_5_28 : IN std_logic ;
      d_arr_merge2_5_27 : IN std_logic ;
      d_arr_merge2_5_26 : IN std_logic ;
      d_arr_merge2_5_25 : IN std_logic ;
      d_arr_merge2_5_24 : IN std_logic ;
      d_arr_merge2_5_23 : IN std_logic ;
      d_arr_merge2_5_22 : IN std_logic ;
      d_arr_merge2_5_21 : IN std_logic ;
      d_arr_merge2_5_20 : IN std_logic ;
      d_arr_merge2_5_19 : IN std_logic ;
      d_arr_merge2_5_18 : IN std_logic ;
      d_arr_merge2_5_17 : IN std_logic ;
      d_arr_merge2_5_16 : IN std_logic ;
      d_arr_merge2_5_15 : IN std_logic ;
      d_arr_merge2_5_14 : IN std_logic ;
      d_arr_merge2_5_13 : IN std_logic ;
      d_arr_merge2_5_12 : IN std_logic ;
      d_arr_merge2_5_11 : IN std_logic ;
      d_arr_merge2_5_10 : IN std_logic ;
      d_arr_merge2_5_9 : IN std_logic ;
      d_arr_merge2_5_8 : IN std_logic ;
      d_arr_merge2_5_7 : IN std_logic ;
      d_arr_merge2_5_6 : IN std_logic ;
      d_arr_merge2_5_5 : IN std_logic ;
      d_arr_merge2_5_4 : IN std_logic ;
      d_arr_merge2_5_3 : IN std_logic ;
      d_arr_merge2_5_2 : IN std_logic ;
      d_arr_merge2_5_1 : IN std_logic ;
      d_arr_merge2_5_0 : IN std_logic ;
      d_arr_merge2_6_31 : IN std_logic ;
      d_arr_merge2_6_30 : IN std_logic ;
      d_arr_merge2_6_29 : IN std_logic ;
      d_arr_merge2_6_28 : IN std_logic ;
      d_arr_merge2_6_27 : IN std_logic ;
      d_arr_merge2_6_26 : IN std_logic ;
      d_arr_merge2_6_25 : IN std_logic ;
      d_arr_merge2_6_24 : IN std_logic ;
      d_arr_merge2_6_23 : IN std_logic ;
      d_arr_merge2_6_22 : IN std_logic ;
      d_arr_merge2_6_21 : IN std_logic ;
      d_arr_merge2_6_20 : IN std_logic ;
      d_arr_merge2_6_19 : IN std_logic ;
      d_arr_merge2_6_18 : IN std_logic ;
      d_arr_merge2_6_17 : IN std_logic ;
      d_arr_merge2_6_16 : IN std_logic ;
      d_arr_merge2_6_15 : IN std_logic ;
      d_arr_merge2_6_14 : IN std_logic ;
      d_arr_merge2_6_13 : IN std_logic ;
      d_arr_merge2_6_12 : IN std_logic ;
      d_arr_merge2_6_11 : IN std_logic ;
      d_arr_merge2_6_10 : IN std_logic ;
      d_arr_merge2_6_9 : IN std_logic ;
      d_arr_merge2_6_8 : IN std_logic ;
      d_arr_merge2_6_7 : IN std_logic ;
      d_arr_merge2_6_6 : IN std_logic ;
      d_arr_merge2_6_5 : IN std_logic ;
      d_arr_merge2_6_4 : IN std_logic ;
      d_arr_merge2_6_3 : IN std_logic ;
      d_arr_merge2_6_2 : IN std_logic ;
      d_arr_merge2_6_1 : IN std_logic ;
      d_arr_merge2_6_0 : IN std_logic ;
      d_arr_merge2_7_31 : IN std_logic ;
      d_arr_merge2_7_30 : IN std_logic ;
      d_arr_merge2_7_29 : IN std_logic ;
      d_arr_merge2_7_28 : IN std_logic ;
      d_arr_merge2_7_27 : IN std_logic ;
      d_arr_merge2_7_26 : IN std_logic ;
      d_arr_merge2_7_25 : IN std_logic ;
      d_arr_merge2_7_24 : IN std_logic ;
      d_arr_merge2_7_23 : IN std_logic ;
      d_arr_merge2_7_22 : IN std_logic ;
      d_arr_merge2_7_21 : IN std_logic ;
      d_arr_merge2_7_20 : IN std_logic ;
      d_arr_merge2_7_19 : IN std_logic ;
      d_arr_merge2_7_18 : IN std_logic ;
      d_arr_merge2_7_17 : IN std_logic ;
      d_arr_merge2_7_16 : IN std_logic ;
      d_arr_merge2_7_15 : IN std_logic ;
      d_arr_merge2_7_14 : IN std_logic ;
      d_arr_merge2_7_13 : IN std_logic ;
      d_arr_merge2_7_12 : IN std_logic ;
      d_arr_merge2_7_11 : IN std_logic ;
      d_arr_merge2_7_10 : IN std_logic ;
      d_arr_merge2_7_9 : IN std_logic ;
      d_arr_merge2_7_8 : IN std_logic ;
      d_arr_merge2_7_7 : IN std_logic ;
      d_arr_merge2_7_6 : IN std_logic ;
      d_arr_merge2_7_5 : IN std_logic ;
      d_arr_merge2_7_4 : IN std_logic ;
      d_arr_merge2_7_3 : IN std_logic ;
      d_arr_merge2_7_2 : IN std_logic ;
      d_arr_merge2_7_1 : IN std_logic ;
      d_arr_merge2_7_0 : IN std_logic ;
      d_arr_merge2_8_31 : IN std_logic ;
      d_arr_merge2_8_30 : IN std_logic ;
      d_arr_merge2_8_29 : IN std_logic ;
      d_arr_merge2_8_28 : IN std_logic ;
      d_arr_merge2_8_27 : IN std_logic ;
      d_arr_merge2_8_26 : IN std_logic ;
      d_arr_merge2_8_25 : IN std_logic ;
      d_arr_merge2_8_24 : IN std_logic ;
      d_arr_merge2_8_23 : IN std_logic ;
      d_arr_merge2_8_22 : IN std_logic ;
      d_arr_merge2_8_21 : IN std_logic ;
      d_arr_merge2_8_20 : IN std_logic ;
      d_arr_merge2_8_19 : IN std_logic ;
      d_arr_merge2_8_18 : IN std_logic ;
      d_arr_merge2_8_17 : IN std_logic ;
      d_arr_merge2_8_16 : IN std_logic ;
      d_arr_merge2_8_15 : IN std_logic ;
      d_arr_merge2_8_14 : IN std_logic ;
      d_arr_merge2_8_13 : IN std_logic ;
      d_arr_merge2_8_12 : IN std_logic ;
      d_arr_merge2_8_11 : IN std_logic ;
      d_arr_merge2_8_10 : IN std_logic ;
      d_arr_merge2_8_9 : IN std_logic ;
      d_arr_merge2_8_8 : IN std_logic ;
      d_arr_merge2_8_7 : IN std_logic ;
      d_arr_merge2_8_6 : IN std_logic ;
      d_arr_merge2_8_5 : IN std_logic ;
      d_arr_merge2_8_4 : IN std_logic ;
      d_arr_merge2_8_3 : IN std_logic ;
      d_arr_merge2_8_2 : IN std_logic ;
      d_arr_merge2_8_1 : IN std_logic ;
      d_arr_merge2_8_0 : IN std_logic ;
      d_arr_merge2_9_31 : IN std_logic ;
      d_arr_merge2_9_30 : IN std_logic ;
      d_arr_merge2_9_29 : IN std_logic ;
      d_arr_merge2_9_28 : IN std_logic ;
      d_arr_merge2_9_27 : IN std_logic ;
      d_arr_merge2_9_26 : IN std_logic ;
      d_arr_merge2_9_25 : IN std_logic ;
      d_arr_merge2_9_24 : IN std_logic ;
      d_arr_merge2_9_23 : IN std_logic ;
      d_arr_merge2_9_22 : IN std_logic ;
      d_arr_merge2_9_21 : IN std_logic ;
      d_arr_merge2_9_20 : IN std_logic ;
      d_arr_merge2_9_19 : IN std_logic ;
      d_arr_merge2_9_18 : IN std_logic ;
      d_arr_merge2_9_17 : IN std_logic ;
      d_arr_merge2_9_16 : IN std_logic ;
      d_arr_merge2_9_15 : IN std_logic ;
      d_arr_merge2_9_14 : IN std_logic ;
      d_arr_merge2_9_13 : IN std_logic ;
      d_arr_merge2_9_12 : IN std_logic ;
      d_arr_merge2_9_11 : IN std_logic ;
      d_arr_merge2_9_10 : IN std_logic ;
      d_arr_merge2_9_9 : IN std_logic ;
      d_arr_merge2_9_8 : IN std_logic ;
      d_arr_merge2_9_7 : IN std_logic ;
      d_arr_merge2_9_6 : IN std_logic ;
      d_arr_merge2_9_5 : IN std_logic ;
      d_arr_merge2_9_4 : IN std_logic ;
      d_arr_merge2_9_3 : IN std_logic ;
      d_arr_merge2_9_2 : IN std_logic ;
      d_arr_merge2_9_1 : IN std_logic ;
      d_arr_merge2_9_0 : IN std_logic ;
      d_arr_merge2_10_31 : IN std_logic ;
      d_arr_merge2_10_30 : IN std_logic ;
      d_arr_merge2_10_29 : IN std_logic ;
      d_arr_merge2_10_28 : IN std_logic ;
      d_arr_merge2_10_27 : IN std_logic ;
      d_arr_merge2_10_26 : IN std_logic ;
      d_arr_merge2_10_25 : IN std_logic ;
      d_arr_merge2_10_24 : IN std_logic ;
      d_arr_merge2_10_23 : IN std_logic ;
      d_arr_merge2_10_22 : IN std_logic ;
      d_arr_merge2_10_21 : IN std_logic ;
      d_arr_merge2_10_20 : IN std_logic ;
      d_arr_merge2_10_19 : IN std_logic ;
      d_arr_merge2_10_18 : IN std_logic ;
      d_arr_merge2_10_17 : IN std_logic ;
      d_arr_merge2_10_16 : IN std_logic ;
      d_arr_merge2_10_15 : IN std_logic ;
      d_arr_merge2_10_14 : IN std_logic ;
      d_arr_merge2_10_13 : IN std_logic ;
      d_arr_merge2_10_12 : IN std_logic ;
      d_arr_merge2_10_11 : IN std_logic ;
      d_arr_merge2_10_10 : IN std_logic ;
      d_arr_merge2_10_9 : IN std_logic ;
      d_arr_merge2_10_8 : IN std_logic ;
      d_arr_merge2_10_7 : IN std_logic ;
      d_arr_merge2_10_6 : IN std_logic ;
      d_arr_merge2_10_5 : IN std_logic ;
      d_arr_merge2_10_4 : IN std_logic ;
      d_arr_merge2_10_3 : IN std_logic ;
      d_arr_merge2_10_2 : IN std_logic ;
      d_arr_merge2_10_1 : IN std_logic ;
      d_arr_merge2_10_0 : IN std_logic ;
      d_arr_merge2_11_31 : IN std_logic ;
      d_arr_merge2_11_30 : IN std_logic ;
      d_arr_merge2_11_29 : IN std_logic ;
      d_arr_merge2_11_28 : IN std_logic ;
      d_arr_merge2_11_27 : IN std_logic ;
      d_arr_merge2_11_26 : IN std_logic ;
      d_arr_merge2_11_25 : IN std_logic ;
      d_arr_merge2_11_24 : IN std_logic ;
      d_arr_merge2_11_23 : IN std_logic ;
      d_arr_merge2_11_22 : IN std_logic ;
      d_arr_merge2_11_21 : IN std_logic ;
      d_arr_merge2_11_20 : IN std_logic ;
      d_arr_merge2_11_19 : IN std_logic ;
      d_arr_merge2_11_18 : IN std_logic ;
      d_arr_merge2_11_17 : IN std_logic ;
      d_arr_merge2_11_16 : IN std_logic ;
      d_arr_merge2_11_15 : IN std_logic ;
      d_arr_merge2_11_14 : IN std_logic ;
      d_arr_merge2_11_13 : IN std_logic ;
      d_arr_merge2_11_12 : IN std_logic ;
      d_arr_merge2_11_11 : IN std_logic ;
      d_arr_merge2_11_10 : IN std_logic ;
      d_arr_merge2_11_9 : IN std_logic ;
      d_arr_merge2_11_8 : IN std_logic ;
      d_arr_merge2_11_7 : IN std_logic ;
      d_arr_merge2_11_6 : IN std_logic ;
      d_arr_merge2_11_5 : IN std_logic ;
      d_arr_merge2_11_4 : IN std_logic ;
      d_arr_merge2_11_3 : IN std_logic ;
      d_arr_merge2_11_2 : IN std_logic ;
      d_arr_merge2_11_1 : IN std_logic ;
      d_arr_merge2_11_0 : IN std_logic ;
      d_arr_merge2_12_31 : IN std_logic ;
      d_arr_merge2_12_30 : IN std_logic ;
      d_arr_merge2_12_29 : IN std_logic ;
      d_arr_merge2_12_28 : IN std_logic ;
      d_arr_merge2_12_27 : IN std_logic ;
      d_arr_merge2_12_26 : IN std_logic ;
      d_arr_merge2_12_25 : IN std_logic ;
      d_arr_merge2_12_24 : IN std_logic ;
      d_arr_merge2_12_23 : IN std_logic ;
      d_arr_merge2_12_22 : IN std_logic ;
      d_arr_merge2_12_21 : IN std_logic ;
      d_arr_merge2_12_20 : IN std_logic ;
      d_arr_merge2_12_19 : IN std_logic ;
      d_arr_merge2_12_18 : IN std_logic ;
      d_arr_merge2_12_17 : IN std_logic ;
      d_arr_merge2_12_16 : IN std_logic ;
      d_arr_merge2_12_15 : IN std_logic ;
      d_arr_merge2_12_14 : IN std_logic ;
      d_arr_merge2_12_13 : IN std_logic ;
      d_arr_merge2_12_12 : IN std_logic ;
      d_arr_merge2_12_11 : IN std_logic ;
      d_arr_merge2_12_10 : IN std_logic ;
      d_arr_merge2_12_9 : IN std_logic ;
      d_arr_merge2_12_8 : IN std_logic ;
      d_arr_merge2_12_7 : IN std_logic ;
      d_arr_merge2_12_6 : IN std_logic ;
      d_arr_merge2_12_5 : IN std_logic ;
      d_arr_merge2_12_4 : IN std_logic ;
      d_arr_merge2_12_3 : IN std_logic ;
      d_arr_merge2_12_2 : IN std_logic ;
      d_arr_merge2_12_1 : IN std_logic ;
      d_arr_merge2_12_0 : IN std_logic ;
      d_arr_merge2_13_31 : IN std_logic ;
      d_arr_merge2_13_30 : IN std_logic ;
      d_arr_merge2_13_29 : IN std_logic ;
      d_arr_merge2_13_28 : IN std_logic ;
      d_arr_merge2_13_27 : IN std_logic ;
      d_arr_merge2_13_26 : IN std_logic ;
      d_arr_merge2_13_25 : IN std_logic ;
      d_arr_merge2_13_24 : IN std_logic ;
      d_arr_merge2_13_23 : IN std_logic ;
      d_arr_merge2_13_22 : IN std_logic ;
      d_arr_merge2_13_21 : IN std_logic ;
      d_arr_merge2_13_20 : IN std_logic ;
      d_arr_merge2_13_19 : IN std_logic ;
      d_arr_merge2_13_18 : IN std_logic ;
      d_arr_merge2_13_17 : IN std_logic ;
      d_arr_merge2_13_16 : IN std_logic ;
      d_arr_merge2_13_15 : IN std_logic ;
      d_arr_merge2_13_14 : IN std_logic ;
      d_arr_merge2_13_13 : IN std_logic ;
      d_arr_merge2_13_12 : IN std_logic ;
      d_arr_merge2_13_11 : IN std_logic ;
      d_arr_merge2_13_10 : IN std_logic ;
      d_arr_merge2_13_9 : IN std_logic ;
      d_arr_merge2_13_8 : IN std_logic ;
      d_arr_merge2_13_7 : IN std_logic ;
      d_arr_merge2_13_6 : IN std_logic ;
      d_arr_merge2_13_5 : IN std_logic ;
      d_arr_merge2_13_4 : IN std_logic ;
      d_arr_merge2_13_3 : IN std_logic ;
      d_arr_merge2_13_2 : IN std_logic ;
      d_arr_merge2_13_1 : IN std_logic ;
      d_arr_merge2_13_0 : IN std_logic ;
      d_arr_merge2_14_31 : IN std_logic ;
      d_arr_merge2_14_30 : IN std_logic ;
      d_arr_merge2_14_29 : IN std_logic ;
      d_arr_merge2_14_28 : IN std_logic ;
      d_arr_merge2_14_27 : IN std_logic ;
      d_arr_merge2_14_26 : IN std_logic ;
      d_arr_merge2_14_25 : IN std_logic ;
      d_arr_merge2_14_24 : IN std_logic ;
      d_arr_merge2_14_23 : IN std_logic ;
      d_arr_merge2_14_22 : IN std_logic ;
      d_arr_merge2_14_21 : IN std_logic ;
      d_arr_merge2_14_20 : IN std_logic ;
      d_arr_merge2_14_19 : IN std_logic ;
      d_arr_merge2_14_18 : IN std_logic ;
      d_arr_merge2_14_17 : IN std_logic ;
      d_arr_merge2_14_16 : IN std_logic ;
      d_arr_merge2_14_15 : IN std_logic ;
      d_arr_merge2_14_14 : IN std_logic ;
      d_arr_merge2_14_13 : IN std_logic ;
      d_arr_merge2_14_12 : IN std_logic ;
      d_arr_merge2_14_11 : IN std_logic ;
      d_arr_merge2_14_10 : IN std_logic ;
      d_arr_merge2_14_9 : IN std_logic ;
      d_arr_merge2_14_8 : IN std_logic ;
      d_arr_merge2_14_7 : IN std_logic ;
      d_arr_merge2_14_6 : IN std_logic ;
      d_arr_merge2_14_5 : IN std_logic ;
      d_arr_merge2_14_4 : IN std_logic ;
      d_arr_merge2_14_3 : IN std_logic ;
      d_arr_merge2_14_2 : IN std_logic ;
      d_arr_merge2_14_1 : IN std_logic ;
      d_arr_merge2_14_0 : IN std_logic ;
      d_arr_merge2_15_31 : IN std_logic ;
      d_arr_merge2_15_30 : IN std_logic ;
      d_arr_merge2_15_29 : IN std_logic ;
      d_arr_merge2_15_28 : IN std_logic ;
      d_arr_merge2_15_27 : IN std_logic ;
      d_arr_merge2_15_26 : IN std_logic ;
      d_arr_merge2_15_25 : IN std_logic ;
      d_arr_merge2_15_24 : IN std_logic ;
      d_arr_merge2_15_23 : IN std_logic ;
      d_arr_merge2_15_22 : IN std_logic ;
      d_arr_merge2_15_21 : IN std_logic ;
      d_arr_merge2_15_20 : IN std_logic ;
      d_arr_merge2_15_19 : IN std_logic ;
      d_arr_merge2_15_18 : IN std_logic ;
      d_arr_merge2_15_17 : IN std_logic ;
      d_arr_merge2_15_16 : IN std_logic ;
      d_arr_merge2_15_15 : IN std_logic ;
      d_arr_merge2_15_14 : IN std_logic ;
      d_arr_merge2_15_13 : IN std_logic ;
      d_arr_merge2_15_12 : IN std_logic ;
      d_arr_merge2_15_11 : IN std_logic ;
      d_arr_merge2_15_10 : IN std_logic ;
      d_arr_merge2_15_9 : IN std_logic ;
      d_arr_merge2_15_8 : IN std_logic ;
      d_arr_merge2_15_7 : IN std_logic ;
      d_arr_merge2_15_6 : IN std_logic ;
      d_arr_merge2_15_5 : IN std_logic ;
      d_arr_merge2_15_4 : IN std_logic ;
      d_arr_merge2_15_3 : IN std_logic ;
      d_arr_merge2_15_2 : IN std_logic ;
      d_arr_merge2_15_1 : IN std_logic ;
      d_arr_merge2_15_0 : IN std_logic ;
      d_arr_merge2_16_31 : IN std_logic ;
      d_arr_merge2_16_30 : IN std_logic ;
      d_arr_merge2_16_29 : IN std_logic ;
      d_arr_merge2_16_28 : IN std_logic ;
      d_arr_merge2_16_27 : IN std_logic ;
      d_arr_merge2_16_26 : IN std_logic ;
      d_arr_merge2_16_25 : IN std_logic ;
      d_arr_merge2_16_24 : IN std_logic ;
      d_arr_merge2_16_23 : IN std_logic ;
      d_arr_merge2_16_22 : IN std_logic ;
      d_arr_merge2_16_21 : IN std_logic ;
      d_arr_merge2_16_20 : IN std_logic ;
      d_arr_merge2_16_19 : IN std_logic ;
      d_arr_merge2_16_18 : IN std_logic ;
      d_arr_merge2_16_17 : IN std_logic ;
      d_arr_merge2_16_16 : IN std_logic ;
      d_arr_merge2_16_15 : IN std_logic ;
      d_arr_merge2_16_14 : IN std_logic ;
      d_arr_merge2_16_13 : IN std_logic ;
      d_arr_merge2_16_12 : IN std_logic ;
      d_arr_merge2_16_11 : IN std_logic ;
      d_arr_merge2_16_10 : IN std_logic ;
      d_arr_merge2_16_9 : IN std_logic ;
      d_arr_merge2_16_8 : IN std_logic ;
      d_arr_merge2_16_7 : IN std_logic ;
      d_arr_merge2_16_6 : IN std_logic ;
      d_arr_merge2_16_5 : IN std_logic ;
      d_arr_merge2_16_4 : IN std_logic ;
      d_arr_merge2_16_3 : IN std_logic ;
      d_arr_merge2_16_2 : IN std_logic ;
      d_arr_merge2_16_1 : IN std_logic ;
      d_arr_merge2_16_0 : IN std_logic ;
      d_arr_merge2_17_31 : IN std_logic ;
      d_arr_merge2_17_30 : IN std_logic ;
      d_arr_merge2_17_29 : IN std_logic ;
      d_arr_merge2_17_28 : IN std_logic ;
      d_arr_merge2_17_27 : IN std_logic ;
      d_arr_merge2_17_26 : IN std_logic ;
      d_arr_merge2_17_25 : IN std_logic ;
      d_arr_merge2_17_24 : IN std_logic ;
      d_arr_merge2_17_23 : IN std_logic ;
      d_arr_merge2_17_22 : IN std_logic ;
      d_arr_merge2_17_21 : IN std_logic ;
      d_arr_merge2_17_20 : IN std_logic ;
      d_arr_merge2_17_19 : IN std_logic ;
      d_arr_merge2_17_18 : IN std_logic ;
      d_arr_merge2_17_17 : IN std_logic ;
      d_arr_merge2_17_16 : IN std_logic ;
      d_arr_merge2_17_15 : IN std_logic ;
      d_arr_merge2_17_14 : IN std_logic ;
      d_arr_merge2_17_13 : IN std_logic ;
      d_arr_merge2_17_12 : IN std_logic ;
      d_arr_merge2_17_11 : IN std_logic ;
      d_arr_merge2_17_10 : IN std_logic ;
      d_arr_merge2_17_9 : IN std_logic ;
      d_arr_merge2_17_8 : IN std_logic ;
      d_arr_merge2_17_7 : IN std_logic ;
      d_arr_merge2_17_6 : IN std_logic ;
      d_arr_merge2_17_5 : IN std_logic ;
      d_arr_merge2_17_4 : IN std_logic ;
      d_arr_merge2_17_3 : IN std_logic ;
      d_arr_merge2_17_2 : IN std_logic ;
      d_arr_merge2_17_1 : IN std_logic ;
      d_arr_merge2_17_0 : IN std_logic ;
      d_arr_merge2_18_31 : IN std_logic ;
      d_arr_merge2_18_30 : IN std_logic ;
      d_arr_merge2_18_29 : IN std_logic ;
      d_arr_merge2_18_28 : IN std_logic ;
      d_arr_merge2_18_27 : IN std_logic ;
      d_arr_merge2_18_26 : IN std_logic ;
      d_arr_merge2_18_25 : IN std_logic ;
      d_arr_merge2_18_24 : IN std_logic ;
      d_arr_merge2_18_23 : IN std_logic ;
      d_arr_merge2_18_22 : IN std_logic ;
      d_arr_merge2_18_21 : IN std_logic ;
      d_arr_merge2_18_20 : IN std_logic ;
      d_arr_merge2_18_19 : IN std_logic ;
      d_arr_merge2_18_18 : IN std_logic ;
      d_arr_merge2_18_17 : IN std_logic ;
      d_arr_merge2_18_16 : IN std_logic ;
      d_arr_merge2_18_15 : IN std_logic ;
      d_arr_merge2_18_14 : IN std_logic ;
      d_arr_merge2_18_13 : IN std_logic ;
      d_arr_merge2_18_12 : IN std_logic ;
      d_arr_merge2_18_11 : IN std_logic ;
      d_arr_merge2_18_10 : IN std_logic ;
      d_arr_merge2_18_9 : IN std_logic ;
      d_arr_merge2_18_8 : IN std_logic ;
      d_arr_merge2_18_7 : IN std_logic ;
      d_arr_merge2_18_6 : IN std_logic ;
      d_arr_merge2_18_5 : IN std_logic ;
      d_arr_merge2_18_4 : IN std_logic ;
      d_arr_merge2_18_3 : IN std_logic ;
      d_arr_merge2_18_2 : IN std_logic ;
      d_arr_merge2_18_1 : IN std_logic ;
      d_arr_merge2_18_0 : IN std_logic ;
      d_arr_merge2_19_31 : IN std_logic ;
      d_arr_merge2_19_30 : IN std_logic ;
      d_arr_merge2_19_29 : IN std_logic ;
      d_arr_merge2_19_28 : IN std_logic ;
      d_arr_merge2_19_27 : IN std_logic ;
      d_arr_merge2_19_26 : IN std_logic ;
      d_arr_merge2_19_25 : IN std_logic ;
      d_arr_merge2_19_24 : IN std_logic ;
      d_arr_merge2_19_23 : IN std_logic ;
      d_arr_merge2_19_22 : IN std_logic ;
      d_arr_merge2_19_21 : IN std_logic ;
      d_arr_merge2_19_20 : IN std_logic ;
      d_arr_merge2_19_19 : IN std_logic ;
      d_arr_merge2_19_18 : IN std_logic ;
      d_arr_merge2_19_17 : IN std_logic ;
      d_arr_merge2_19_16 : IN std_logic ;
      d_arr_merge2_19_15 : IN std_logic ;
      d_arr_merge2_19_14 : IN std_logic ;
      d_arr_merge2_19_13 : IN std_logic ;
      d_arr_merge2_19_12 : IN std_logic ;
      d_arr_merge2_19_11 : IN std_logic ;
      d_arr_merge2_19_10 : IN std_logic ;
      d_arr_merge2_19_9 : IN std_logic ;
      d_arr_merge2_19_8 : IN std_logic ;
      d_arr_merge2_19_7 : IN std_logic ;
      d_arr_merge2_19_6 : IN std_logic ;
      d_arr_merge2_19_5 : IN std_logic ;
      d_arr_merge2_19_4 : IN std_logic ;
      d_arr_merge2_19_3 : IN std_logic ;
      d_arr_merge2_19_2 : IN std_logic ;
      d_arr_merge2_19_1 : IN std_logic ;
      d_arr_merge2_19_0 : IN std_logic ;
      d_arr_merge2_20_31 : IN std_logic ;
      d_arr_merge2_20_30 : IN std_logic ;
      d_arr_merge2_20_29 : IN std_logic ;
      d_arr_merge2_20_28 : IN std_logic ;
      d_arr_merge2_20_27 : IN std_logic ;
      d_arr_merge2_20_26 : IN std_logic ;
      d_arr_merge2_20_25 : IN std_logic ;
      d_arr_merge2_20_24 : IN std_logic ;
      d_arr_merge2_20_23 : IN std_logic ;
      d_arr_merge2_20_22 : IN std_logic ;
      d_arr_merge2_20_21 : IN std_logic ;
      d_arr_merge2_20_20 : IN std_logic ;
      d_arr_merge2_20_19 : IN std_logic ;
      d_arr_merge2_20_18 : IN std_logic ;
      d_arr_merge2_20_17 : IN std_logic ;
      d_arr_merge2_20_16 : IN std_logic ;
      d_arr_merge2_20_15 : IN std_logic ;
      d_arr_merge2_20_14 : IN std_logic ;
      d_arr_merge2_20_13 : IN std_logic ;
      d_arr_merge2_20_12 : IN std_logic ;
      d_arr_merge2_20_11 : IN std_logic ;
      d_arr_merge2_20_10 : IN std_logic ;
      d_arr_merge2_20_9 : IN std_logic ;
      d_arr_merge2_20_8 : IN std_logic ;
      d_arr_merge2_20_7 : IN std_logic ;
      d_arr_merge2_20_6 : IN std_logic ;
      d_arr_merge2_20_5 : IN std_logic ;
      d_arr_merge2_20_4 : IN std_logic ;
      d_arr_merge2_20_3 : IN std_logic ;
      d_arr_merge2_20_2 : IN std_logic ;
      d_arr_merge2_20_1 : IN std_logic ;
      d_arr_merge2_20_0 : IN std_logic ;
      d_arr_merge2_21_31 : IN std_logic ;
      d_arr_merge2_21_30 : IN std_logic ;
      d_arr_merge2_21_29 : IN std_logic ;
      d_arr_merge2_21_28 : IN std_logic ;
      d_arr_merge2_21_27 : IN std_logic ;
      d_arr_merge2_21_26 : IN std_logic ;
      d_arr_merge2_21_25 : IN std_logic ;
      d_arr_merge2_21_24 : IN std_logic ;
      d_arr_merge2_21_23 : IN std_logic ;
      d_arr_merge2_21_22 : IN std_logic ;
      d_arr_merge2_21_21 : IN std_logic ;
      d_arr_merge2_21_20 : IN std_logic ;
      d_arr_merge2_21_19 : IN std_logic ;
      d_arr_merge2_21_18 : IN std_logic ;
      d_arr_merge2_21_17 : IN std_logic ;
      d_arr_merge2_21_16 : IN std_logic ;
      d_arr_merge2_21_15 : IN std_logic ;
      d_arr_merge2_21_14 : IN std_logic ;
      d_arr_merge2_21_13 : IN std_logic ;
      d_arr_merge2_21_12 : IN std_logic ;
      d_arr_merge2_21_11 : IN std_logic ;
      d_arr_merge2_21_10 : IN std_logic ;
      d_arr_merge2_21_9 : IN std_logic ;
      d_arr_merge2_21_8 : IN std_logic ;
      d_arr_merge2_21_7 : IN std_logic ;
      d_arr_merge2_21_6 : IN std_logic ;
      d_arr_merge2_21_5 : IN std_logic ;
      d_arr_merge2_21_4 : IN std_logic ;
      d_arr_merge2_21_3 : IN std_logic ;
      d_arr_merge2_21_2 : IN std_logic ;
      d_arr_merge2_21_1 : IN std_logic ;
      d_arr_merge2_21_0 : IN std_logic ;
      d_arr_merge2_22_31 : IN std_logic ;
      d_arr_merge2_22_30 : IN std_logic ;
      d_arr_merge2_22_29 : IN std_logic ;
      d_arr_merge2_22_28 : IN std_logic ;
      d_arr_merge2_22_27 : IN std_logic ;
      d_arr_merge2_22_26 : IN std_logic ;
      d_arr_merge2_22_25 : IN std_logic ;
      d_arr_merge2_22_24 : IN std_logic ;
      d_arr_merge2_22_23 : IN std_logic ;
      d_arr_merge2_22_22 : IN std_logic ;
      d_arr_merge2_22_21 : IN std_logic ;
      d_arr_merge2_22_20 : IN std_logic ;
      d_arr_merge2_22_19 : IN std_logic ;
      d_arr_merge2_22_18 : IN std_logic ;
      d_arr_merge2_22_17 : IN std_logic ;
      d_arr_merge2_22_16 : IN std_logic ;
      d_arr_merge2_22_15 : IN std_logic ;
      d_arr_merge2_22_14 : IN std_logic ;
      d_arr_merge2_22_13 : IN std_logic ;
      d_arr_merge2_22_12 : IN std_logic ;
      d_arr_merge2_22_11 : IN std_logic ;
      d_arr_merge2_22_10 : IN std_logic ;
      d_arr_merge2_22_9 : IN std_logic ;
      d_arr_merge2_22_8 : IN std_logic ;
      d_arr_merge2_22_7 : IN std_logic ;
      d_arr_merge2_22_6 : IN std_logic ;
      d_arr_merge2_22_5 : IN std_logic ;
      d_arr_merge2_22_4 : IN std_logic ;
      d_arr_merge2_22_3 : IN std_logic ;
      d_arr_merge2_22_2 : IN std_logic ;
      d_arr_merge2_22_1 : IN std_logic ;
      d_arr_merge2_22_0 : IN std_logic ;
      d_arr_merge2_23_31 : IN std_logic ;
      d_arr_merge2_23_30 : IN std_logic ;
      d_arr_merge2_23_29 : IN std_logic ;
      d_arr_merge2_23_28 : IN std_logic ;
      d_arr_merge2_23_27 : IN std_logic ;
      d_arr_merge2_23_26 : IN std_logic ;
      d_arr_merge2_23_25 : IN std_logic ;
      d_arr_merge2_23_24 : IN std_logic ;
      d_arr_merge2_23_23 : IN std_logic ;
      d_arr_merge2_23_22 : IN std_logic ;
      d_arr_merge2_23_21 : IN std_logic ;
      d_arr_merge2_23_20 : IN std_logic ;
      d_arr_merge2_23_19 : IN std_logic ;
      d_arr_merge2_23_18 : IN std_logic ;
      d_arr_merge2_23_17 : IN std_logic ;
      d_arr_merge2_23_16 : IN std_logic ;
      d_arr_merge2_23_15 : IN std_logic ;
      d_arr_merge2_23_14 : IN std_logic ;
      d_arr_merge2_23_13 : IN std_logic ;
      d_arr_merge2_23_12 : IN std_logic ;
      d_arr_merge2_23_11 : IN std_logic ;
      d_arr_merge2_23_10 : IN std_logic ;
      d_arr_merge2_23_9 : IN std_logic ;
      d_arr_merge2_23_8 : IN std_logic ;
      d_arr_merge2_23_7 : IN std_logic ;
      d_arr_merge2_23_6 : IN std_logic ;
      d_arr_merge2_23_5 : IN std_logic ;
      d_arr_merge2_23_4 : IN std_logic ;
      d_arr_merge2_23_3 : IN std_logic ;
      d_arr_merge2_23_2 : IN std_logic ;
      d_arr_merge2_23_1 : IN std_logic ;
      d_arr_merge2_23_0 : IN std_logic ;
      d_arr_merge2_24_31 : IN std_logic ;
      d_arr_merge2_24_30 : IN std_logic ;
      d_arr_merge2_24_29 : IN std_logic ;
      d_arr_merge2_24_28 : IN std_logic ;
      d_arr_merge2_24_27 : IN std_logic ;
      d_arr_merge2_24_26 : IN std_logic ;
      d_arr_merge2_24_25 : IN std_logic ;
      d_arr_merge2_24_24 : IN std_logic ;
      d_arr_merge2_24_23 : IN std_logic ;
      d_arr_merge2_24_22 : IN std_logic ;
      d_arr_merge2_24_21 : IN std_logic ;
      d_arr_merge2_24_20 : IN std_logic ;
      d_arr_merge2_24_19 : IN std_logic ;
      d_arr_merge2_24_18 : IN std_logic ;
      d_arr_merge2_24_17 : IN std_logic ;
      d_arr_merge2_24_16 : IN std_logic ;
      d_arr_merge2_24_15 : IN std_logic ;
      d_arr_merge2_24_14 : IN std_logic ;
      d_arr_merge2_24_13 : IN std_logic ;
      d_arr_merge2_24_12 : IN std_logic ;
      d_arr_merge2_24_11 : IN std_logic ;
      d_arr_merge2_24_10 : IN std_logic ;
      d_arr_merge2_24_9 : IN std_logic ;
      d_arr_merge2_24_8 : IN std_logic ;
      d_arr_merge2_24_7 : IN std_logic ;
      d_arr_merge2_24_6 : IN std_logic ;
      d_arr_merge2_24_5 : IN std_logic ;
      d_arr_merge2_24_4 : IN std_logic ;
      d_arr_merge2_24_3 : IN std_logic ;
      d_arr_merge2_24_2 : IN std_logic ;
      d_arr_merge2_24_1 : IN std_logic ;
      d_arr_merge2_24_0 : IN std_logic ;
      d_arr_relu_0_31 : IN std_logic ;
      d_arr_relu_0_30 : IN std_logic ;
      d_arr_relu_0_29 : IN std_logic ;
      d_arr_relu_0_28 : IN std_logic ;
      d_arr_relu_0_27 : IN std_logic ;
      d_arr_relu_0_26 : IN std_logic ;
      d_arr_relu_0_25 : IN std_logic ;
      d_arr_relu_0_24 : IN std_logic ;
      d_arr_relu_0_23 : IN std_logic ;
      d_arr_relu_0_22 : IN std_logic ;
      d_arr_relu_0_21 : IN std_logic ;
      d_arr_relu_0_20 : IN std_logic ;
      d_arr_relu_0_19 : IN std_logic ;
      d_arr_relu_0_18 : IN std_logic ;
      d_arr_relu_0_17 : IN std_logic ;
      d_arr_relu_0_16 : IN std_logic ;
      d_arr_relu_0_15 : IN std_logic ;
      d_arr_relu_0_14 : IN std_logic ;
      d_arr_relu_0_13 : IN std_logic ;
      d_arr_relu_0_12 : IN std_logic ;
      d_arr_relu_0_11 : IN std_logic ;
      d_arr_relu_0_10 : IN std_logic ;
      d_arr_relu_0_9 : IN std_logic ;
      d_arr_relu_0_8 : IN std_logic ;
      d_arr_relu_0_7 : IN std_logic ;
      d_arr_relu_0_6 : IN std_logic ;
      d_arr_relu_0_5 : IN std_logic ;
      d_arr_relu_0_4 : IN std_logic ;
      d_arr_relu_0_3 : IN std_logic ;
      d_arr_relu_0_2 : IN std_logic ;
      d_arr_relu_0_1 : IN std_logic ;
      d_arr_relu_0_0 : IN std_logic ;
      d_arr_relu_1_31 : IN std_logic ;
      d_arr_relu_1_30 : IN std_logic ;
      d_arr_relu_1_29 : IN std_logic ;
      d_arr_relu_1_28 : IN std_logic ;
      d_arr_relu_1_27 : IN std_logic ;
      d_arr_relu_1_26 : IN std_logic ;
      d_arr_relu_1_25 : IN std_logic ;
      d_arr_relu_1_24 : IN std_logic ;
      d_arr_relu_1_23 : IN std_logic ;
      d_arr_relu_1_22 : IN std_logic ;
      d_arr_relu_1_21 : IN std_logic ;
      d_arr_relu_1_20 : IN std_logic ;
      d_arr_relu_1_19 : IN std_logic ;
      d_arr_relu_1_18 : IN std_logic ;
      d_arr_relu_1_17 : IN std_logic ;
      d_arr_relu_1_16 : IN std_logic ;
      d_arr_relu_1_15 : IN std_logic ;
      d_arr_relu_1_14 : IN std_logic ;
      d_arr_relu_1_13 : IN std_logic ;
      d_arr_relu_1_12 : IN std_logic ;
      d_arr_relu_1_11 : IN std_logic ;
      d_arr_relu_1_10 : IN std_logic ;
      d_arr_relu_1_9 : IN std_logic ;
      d_arr_relu_1_8 : IN std_logic ;
      d_arr_relu_1_7 : IN std_logic ;
      d_arr_relu_1_6 : IN std_logic ;
      d_arr_relu_1_5 : IN std_logic ;
      d_arr_relu_1_4 : IN std_logic ;
      d_arr_relu_1_3 : IN std_logic ;
      d_arr_relu_1_2 : IN std_logic ;
      d_arr_relu_1_1 : IN std_logic ;
      d_arr_relu_1_0 : IN std_logic ;
      d_arr_relu_2_31 : IN std_logic ;
      d_arr_relu_2_30 : IN std_logic ;
      d_arr_relu_2_29 : IN std_logic ;
      d_arr_relu_2_28 : IN std_logic ;
      d_arr_relu_2_27 : IN std_logic ;
      d_arr_relu_2_26 : IN std_logic ;
      d_arr_relu_2_25 : IN std_logic ;
      d_arr_relu_2_24 : IN std_logic ;
      d_arr_relu_2_23 : IN std_logic ;
      d_arr_relu_2_22 : IN std_logic ;
      d_arr_relu_2_21 : IN std_logic ;
      d_arr_relu_2_20 : IN std_logic ;
      d_arr_relu_2_19 : IN std_logic ;
      d_arr_relu_2_18 : IN std_logic ;
      d_arr_relu_2_17 : IN std_logic ;
      d_arr_relu_2_16 : IN std_logic ;
      d_arr_relu_2_15 : IN std_logic ;
      d_arr_relu_2_14 : IN std_logic ;
      d_arr_relu_2_13 : IN std_logic ;
      d_arr_relu_2_12 : IN std_logic ;
      d_arr_relu_2_11 : IN std_logic ;
      d_arr_relu_2_10 : IN std_logic ;
      d_arr_relu_2_9 : IN std_logic ;
      d_arr_relu_2_8 : IN std_logic ;
      d_arr_relu_2_7 : IN std_logic ;
      d_arr_relu_2_6 : IN std_logic ;
      d_arr_relu_2_5 : IN std_logic ;
      d_arr_relu_2_4 : IN std_logic ;
      d_arr_relu_2_3 : IN std_logic ;
      d_arr_relu_2_2 : IN std_logic ;
      d_arr_relu_2_1 : IN std_logic ;
      d_arr_relu_2_0 : IN std_logic ;
      d_arr_relu_3_31 : IN std_logic ;
      d_arr_relu_3_30 : IN std_logic ;
      d_arr_relu_3_29 : IN std_logic ;
      d_arr_relu_3_28 : IN std_logic ;
      d_arr_relu_3_27 : IN std_logic ;
      d_arr_relu_3_26 : IN std_logic ;
      d_arr_relu_3_25 : IN std_logic ;
      d_arr_relu_3_24 : IN std_logic ;
      d_arr_relu_3_23 : IN std_logic ;
      d_arr_relu_3_22 : IN std_logic ;
      d_arr_relu_3_21 : IN std_logic ;
      d_arr_relu_3_20 : IN std_logic ;
      d_arr_relu_3_19 : IN std_logic ;
      d_arr_relu_3_18 : IN std_logic ;
      d_arr_relu_3_17 : IN std_logic ;
      d_arr_relu_3_16 : IN std_logic ;
      d_arr_relu_3_15 : IN std_logic ;
      d_arr_relu_3_14 : IN std_logic ;
      d_arr_relu_3_13 : IN std_logic ;
      d_arr_relu_3_12 : IN std_logic ;
      d_arr_relu_3_11 : IN std_logic ;
      d_arr_relu_3_10 : IN std_logic ;
      d_arr_relu_3_9 : IN std_logic ;
      d_arr_relu_3_8 : IN std_logic ;
      d_arr_relu_3_7 : IN std_logic ;
      d_arr_relu_3_6 : IN std_logic ;
      d_arr_relu_3_5 : IN std_logic ;
      d_arr_relu_3_4 : IN std_logic ;
      d_arr_relu_3_3 : IN std_logic ;
      d_arr_relu_3_2 : IN std_logic ;
      d_arr_relu_3_1 : IN std_logic ;
      d_arr_relu_3_0 : IN std_logic ;
      d_arr_relu_4_31 : IN std_logic ;
      d_arr_relu_4_30 : IN std_logic ;
      d_arr_relu_4_29 : IN std_logic ;
      d_arr_relu_4_28 : IN std_logic ;
      d_arr_relu_4_27 : IN std_logic ;
      d_arr_relu_4_26 : IN std_logic ;
      d_arr_relu_4_25 : IN std_logic ;
      d_arr_relu_4_24 : IN std_logic ;
      d_arr_relu_4_23 : IN std_logic ;
      d_arr_relu_4_22 : IN std_logic ;
      d_arr_relu_4_21 : IN std_logic ;
      d_arr_relu_4_20 : IN std_logic ;
      d_arr_relu_4_19 : IN std_logic ;
      d_arr_relu_4_18 : IN std_logic ;
      d_arr_relu_4_17 : IN std_logic ;
      d_arr_relu_4_16 : IN std_logic ;
      d_arr_relu_4_15 : IN std_logic ;
      d_arr_relu_4_14 : IN std_logic ;
      d_arr_relu_4_13 : IN std_logic ;
      d_arr_relu_4_12 : IN std_logic ;
      d_arr_relu_4_11 : IN std_logic ;
      d_arr_relu_4_10 : IN std_logic ;
      d_arr_relu_4_9 : IN std_logic ;
      d_arr_relu_4_8 : IN std_logic ;
      d_arr_relu_4_7 : IN std_logic ;
      d_arr_relu_4_6 : IN std_logic ;
      d_arr_relu_4_5 : IN std_logic ;
      d_arr_relu_4_4 : IN std_logic ;
      d_arr_relu_4_3 : IN std_logic ;
      d_arr_relu_4_2 : IN std_logic ;
      d_arr_relu_4_1 : IN std_logic ;
      d_arr_relu_4_0 : IN std_logic ;
      d_arr_relu_5_31 : IN std_logic ;
      d_arr_relu_5_30 : IN std_logic ;
      d_arr_relu_5_29 : IN std_logic ;
      d_arr_relu_5_28 : IN std_logic ;
      d_arr_relu_5_27 : IN std_logic ;
      d_arr_relu_5_26 : IN std_logic ;
      d_arr_relu_5_25 : IN std_logic ;
      d_arr_relu_5_24 : IN std_logic ;
      d_arr_relu_5_23 : IN std_logic ;
      d_arr_relu_5_22 : IN std_logic ;
      d_arr_relu_5_21 : IN std_logic ;
      d_arr_relu_5_20 : IN std_logic ;
      d_arr_relu_5_19 : IN std_logic ;
      d_arr_relu_5_18 : IN std_logic ;
      d_arr_relu_5_17 : IN std_logic ;
      d_arr_relu_5_16 : IN std_logic ;
      d_arr_relu_5_15 : IN std_logic ;
      d_arr_relu_5_14 : IN std_logic ;
      d_arr_relu_5_13 : IN std_logic ;
      d_arr_relu_5_12 : IN std_logic ;
      d_arr_relu_5_11 : IN std_logic ;
      d_arr_relu_5_10 : IN std_logic ;
      d_arr_relu_5_9 : IN std_logic ;
      d_arr_relu_5_8 : IN std_logic ;
      d_arr_relu_5_7 : IN std_logic ;
      d_arr_relu_5_6 : IN std_logic ;
      d_arr_relu_5_5 : IN std_logic ;
      d_arr_relu_5_4 : IN std_logic ;
      d_arr_relu_5_3 : IN std_logic ;
      d_arr_relu_5_2 : IN std_logic ;
      d_arr_relu_5_1 : IN std_logic ;
      d_arr_relu_5_0 : IN std_logic ;
      d_arr_relu_6_31 : IN std_logic ;
      d_arr_relu_6_30 : IN std_logic ;
      d_arr_relu_6_29 : IN std_logic ;
      d_arr_relu_6_28 : IN std_logic ;
      d_arr_relu_6_27 : IN std_logic ;
      d_arr_relu_6_26 : IN std_logic ;
      d_arr_relu_6_25 : IN std_logic ;
      d_arr_relu_6_24 : IN std_logic ;
      d_arr_relu_6_23 : IN std_logic ;
      d_arr_relu_6_22 : IN std_logic ;
      d_arr_relu_6_21 : IN std_logic ;
      d_arr_relu_6_20 : IN std_logic ;
      d_arr_relu_6_19 : IN std_logic ;
      d_arr_relu_6_18 : IN std_logic ;
      d_arr_relu_6_17 : IN std_logic ;
      d_arr_relu_6_16 : IN std_logic ;
      d_arr_relu_6_15 : IN std_logic ;
      d_arr_relu_6_14 : IN std_logic ;
      d_arr_relu_6_13 : IN std_logic ;
      d_arr_relu_6_12 : IN std_logic ;
      d_arr_relu_6_11 : IN std_logic ;
      d_arr_relu_6_10 : IN std_logic ;
      d_arr_relu_6_9 : IN std_logic ;
      d_arr_relu_6_8 : IN std_logic ;
      d_arr_relu_6_7 : IN std_logic ;
      d_arr_relu_6_6 : IN std_logic ;
      d_arr_relu_6_5 : IN std_logic ;
      d_arr_relu_6_4 : IN std_logic ;
      d_arr_relu_6_3 : IN std_logic ;
      d_arr_relu_6_2 : IN std_logic ;
      d_arr_relu_6_1 : IN std_logic ;
      d_arr_relu_6_0 : IN std_logic ;
      d_arr_relu_7_31 : IN std_logic ;
      d_arr_relu_7_30 : IN std_logic ;
      d_arr_relu_7_29 : IN std_logic ;
      d_arr_relu_7_28 : IN std_logic ;
      d_arr_relu_7_27 : IN std_logic ;
      d_arr_relu_7_26 : IN std_logic ;
      d_arr_relu_7_25 : IN std_logic ;
      d_arr_relu_7_24 : IN std_logic ;
      d_arr_relu_7_23 : IN std_logic ;
      d_arr_relu_7_22 : IN std_logic ;
      d_arr_relu_7_21 : IN std_logic ;
      d_arr_relu_7_20 : IN std_logic ;
      d_arr_relu_7_19 : IN std_logic ;
      d_arr_relu_7_18 : IN std_logic ;
      d_arr_relu_7_17 : IN std_logic ;
      d_arr_relu_7_16 : IN std_logic ;
      d_arr_relu_7_15 : IN std_logic ;
      d_arr_relu_7_14 : IN std_logic ;
      d_arr_relu_7_13 : IN std_logic ;
      d_arr_relu_7_12 : IN std_logic ;
      d_arr_relu_7_11 : IN std_logic ;
      d_arr_relu_7_10 : IN std_logic ;
      d_arr_relu_7_9 : IN std_logic ;
      d_arr_relu_7_8 : IN std_logic ;
      d_arr_relu_7_7 : IN std_logic ;
      d_arr_relu_7_6 : IN std_logic ;
      d_arr_relu_7_5 : IN std_logic ;
      d_arr_relu_7_4 : IN std_logic ;
      d_arr_relu_7_3 : IN std_logic ;
      d_arr_relu_7_2 : IN std_logic ;
      d_arr_relu_7_1 : IN std_logic ;
      d_arr_relu_7_0 : IN std_logic ;
      d_arr_relu_8_31 : IN std_logic ;
      d_arr_relu_8_30 : IN std_logic ;
      d_arr_relu_8_29 : IN std_logic ;
      d_arr_relu_8_28 : IN std_logic ;
      d_arr_relu_8_27 : IN std_logic ;
      d_arr_relu_8_26 : IN std_logic ;
      d_arr_relu_8_25 : IN std_logic ;
      d_arr_relu_8_24 : IN std_logic ;
      d_arr_relu_8_23 : IN std_logic ;
      d_arr_relu_8_22 : IN std_logic ;
      d_arr_relu_8_21 : IN std_logic ;
      d_arr_relu_8_20 : IN std_logic ;
      d_arr_relu_8_19 : IN std_logic ;
      d_arr_relu_8_18 : IN std_logic ;
      d_arr_relu_8_17 : IN std_logic ;
      d_arr_relu_8_16 : IN std_logic ;
      d_arr_relu_8_15 : IN std_logic ;
      d_arr_relu_8_14 : IN std_logic ;
      d_arr_relu_8_13 : IN std_logic ;
      d_arr_relu_8_12 : IN std_logic ;
      d_arr_relu_8_11 : IN std_logic ;
      d_arr_relu_8_10 : IN std_logic ;
      d_arr_relu_8_9 : IN std_logic ;
      d_arr_relu_8_8 : IN std_logic ;
      d_arr_relu_8_7 : IN std_logic ;
      d_arr_relu_8_6 : IN std_logic ;
      d_arr_relu_8_5 : IN std_logic ;
      d_arr_relu_8_4 : IN std_logic ;
      d_arr_relu_8_3 : IN std_logic ;
      d_arr_relu_8_2 : IN std_logic ;
      d_arr_relu_8_1 : IN std_logic ;
      d_arr_relu_8_0 : IN std_logic ;
      d_arr_relu_9_31 : IN std_logic ;
      d_arr_relu_9_30 : IN std_logic ;
      d_arr_relu_9_29 : IN std_logic ;
      d_arr_relu_9_28 : IN std_logic ;
      d_arr_relu_9_27 : IN std_logic ;
      d_arr_relu_9_26 : IN std_logic ;
      d_arr_relu_9_25 : IN std_logic ;
      d_arr_relu_9_24 : IN std_logic ;
      d_arr_relu_9_23 : IN std_logic ;
      d_arr_relu_9_22 : IN std_logic ;
      d_arr_relu_9_21 : IN std_logic ;
      d_arr_relu_9_20 : IN std_logic ;
      d_arr_relu_9_19 : IN std_logic ;
      d_arr_relu_9_18 : IN std_logic ;
      d_arr_relu_9_17 : IN std_logic ;
      d_arr_relu_9_16 : IN std_logic ;
      d_arr_relu_9_15 : IN std_logic ;
      d_arr_relu_9_14 : IN std_logic ;
      d_arr_relu_9_13 : IN std_logic ;
      d_arr_relu_9_12 : IN std_logic ;
      d_arr_relu_9_11 : IN std_logic ;
      d_arr_relu_9_10 : IN std_logic ;
      d_arr_relu_9_9 : IN std_logic ;
      d_arr_relu_9_8 : IN std_logic ;
      d_arr_relu_9_7 : IN std_logic ;
      d_arr_relu_9_6 : IN std_logic ;
      d_arr_relu_9_5 : IN std_logic ;
      d_arr_relu_9_4 : IN std_logic ;
      d_arr_relu_9_3 : IN std_logic ;
      d_arr_relu_9_2 : IN std_logic ;
      d_arr_relu_9_1 : IN std_logic ;
      d_arr_relu_9_0 : IN std_logic ;
      d_arr_relu_10_31 : IN std_logic ;
      d_arr_relu_10_30 : IN std_logic ;
      d_arr_relu_10_29 : IN std_logic ;
      d_arr_relu_10_28 : IN std_logic ;
      d_arr_relu_10_27 : IN std_logic ;
      d_arr_relu_10_26 : IN std_logic ;
      d_arr_relu_10_25 : IN std_logic ;
      d_arr_relu_10_24 : IN std_logic ;
      d_arr_relu_10_23 : IN std_logic ;
      d_arr_relu_10_22 : IN std_logic ;
      d_arr_relu_10_21 : IN std_logic ;
      d_arr_relu_10_20 : IN std_logic ;
      d_arr_relu_10_19 : IN std_logic ;
      d_arr_relu_10_18 : IN std_logic ;
      d_arr_relu_10_17 : IN std_logic ;
      d_arr_relu_10_16 : IN std_logic ;
      d_arr_relu_10_15 : IN std_logic ;
      d_arr_relu_10_14 : IN std_logic ;
      d_arr_relu_10_13 : IN std_logic ;
      d_arr_relu_10_12 : IN std_logic ;
      d_arr_relu_10_11 : IN std_logic ;
      d_arr_relu_10_10 : IN std_logic ;
      d_arr_relu_10_9 : IN std_logic ;
      d_arr_relu_10_8 : IN std_logic ;
      d_arr_relu_10_7 : IN std_logic ;
      d_arr_relu_10_6 : IN std_logic ;
      d_arr_relu_10_5 : IN std_logic ;
      d_arr_relu_10_4 : IN std_logic ;
      d_arr_relu_10_3 : IN std_logic ;
      d_arr_relu_10_2 : IN std_logic ;
      d_arr_relu_10_1 : IN std_logic ;
      d_arr_relu_10_0 : IN std_logic ;
      d_arr_relu_11_31 : IN std_logic ;
      d_arr_relu_11_30 : IN std_logic ;
      d_arr_relu_11_29 : IN std_logic ;
      d_arr_relu_11_28 : IN std_logic ;
      d_arr_relu_11_27 : IN std_logic ;
      d_arr_relu_11_26 : IN std_logic ;
      d_arr_relu_11_25 : IN std_logic ;
      d_arr_relu_11_24 : IN std_logic ;
      d_arr_relu_11_23 : IN std_logic ;
      d_arr_relu_11_22 : IN std_logic ;
      d_arr_relu_11_21 : IN std_logic ;
      d_arr_relu_11_20 : IN std_logic ;
      d_arr_relu_11_19 : IN std_logic ;
      d_arr_relu_11_18 : IN std_logic ;
      d_arr_relu_11_17 : IN std_logic ;
      d_arr_relu_11_16 : IN std_logic ;
      d_arr_relu_11_15 : IN std_logic ;
      d_arr_relu_11_14 : IN std_logic ;
      d_arr_relu_11_13 : IN std_logic ;
      d_arr_relu_11_12 : IN std_logic ;
      d_arr_relu_11_11 : IN std_logic ;
      d_arr_relu_11_10 : IN std_logic ;
      d_arr_relu_11_9 : IN std_logic ;
      d_arr_relu_11_8 : IN std_logic ;
      d_arr_relu_11_7 : IN std_logic ;
      d_arr_relu_11_6 : IN std_logic ;
      d_arr_relu_11_5 : IN std_logic ;
      d_arr_relu_11_4 : IN std_logic ;
      d_arr_relu_11_3 : IN std_logic ;
      d_arr_relu_11_2 : IN std_logic ;
      d_arr_relu_11_1 : IN std_logic ;
      d_arr_relu_11_0 : IN std_logic ;
      d_arr_relu_12_31 : IN std_logic ;
      d_arr_relu_12_30 : IN std_logic ;
      d_arr_relu_12_29 : IN std_logic ;
      d_arr_relu_12_28 : IN std_logic ;
      d_arr_relu_12_27 : IN std_logic ;
      d_arr_relu_12_26 : IN std_logic ;
      d_arr_relu_12_25 : IN std_logic ;
      d_arr_relu_12_24 : IN std_logic ;
      d_arr_relu_12_23 : IN std_logic ;
      d_arr_relu_12_22 : IN std_logic ;
      d_arr_relu_12_21 : IN std_logic ;
      d_arr_relu_12_20 : IN std_logic ;
      d_arr_relu_12_19 : IN std_logic ;
      d_arr_relu_12_18 : IN std_logic ;
      d_arr_relu_12_17 : IN std_logic ;
      d_arr_relu_12_16 : IN std_logic ;
      d_arr_relu_12_15 : IN std_logic ;
      d_arr_relu_12_14 : IN std_logic ;
      d_arr_relu_12_13 : IN std_logic ;
      d_arr_relu_12_12 : IN std_logic ;
      d_arr_relu_12_11 : IN std_logic ;
      d_arr_relu_12_10 : IN std_logic ;
      d_arr_relu_12_9 : IN std_logic ;
      d_arr_relu_12_8 : IN std_logic ;
      d_arr_relu_12_7 : IN std_logic ;
      d_arr_relu_12_6 : IN std_logic ;
      d_arr_relu_12_5 : IN std_logic ;
      d_arr_relu_12_4 : IN std_logic ;
      d_arr_relu_12_3 : IN std_logic ;
      d_arr_relu_12_2 : IN std_logic ;
      d_arr_relu_12_1 : IN std_logic ;
      d_arr_relu_12_0 : IN std_logic ;
      d_arr_relu_13_31 : IN std_logic ;
      d_arr_relu_13_30 : IN std_logic ;
      d_arr_relu_13_29 : IN std_logic ;
      d_arr_relu_13_28 : IN std_logic ;
      d_arr_relu_13_27 : IN std_logic ;
      d_arr_relu_13_26 : IN std_logic ;
      d_arr_relu_13_25 : IN std_logic ;
      d_arr_relu_13_24 : IN std_logic ;
      d_arr_relu_13_23 : IN std_logic ;
      d_arr_relu_13_22 : IN std_logic ;
      d_arr_relu_13_21 : IN std_logic ;
      d_arr_relu_13_20 : IN std_logic ;
      d_arr_relu_13_19 : IN std_logic ;
      d_arr_relu_13_18 : IN std_logic ;
      d_arr_relu_13_17 : IN std_logic ;
      d_arr_relu_13_16 : IN std_logic ;
      d_arr_relu_13_15 : IN std_logic ;
      d_arr_relu_13_14 : IN std_logic ;
      d_arr_relu_13_13 : IN std_logic ;
      d_arr_relu_13_12 : IN std_logic ;
      d_arr_relu_13_11 : IN std_logic ;
      d_arr_relu_13_10 : IN std_logic ;
      d_arr_relu_13_9 : IN std_logic ;
      d_arr_relu_13_8 : IN std_logic ;
      d_arr_relu_13_7 : IN std_logic ;
      d_arr_relu_13_6 : IN std_logic ;
      d_arr_relu_13_5 : IN std_logic ;
      d_arr_relu_13_4 : IN std_logic ;
      d_arr_relu_13_3 : IN std_logic ;
      d_arr_relu_13_2 : IN std_logic ;
      d_arr_relu_13_1 : IN std_logic ;
      d_arr_relu_13_0 : IN std_logic ;
      d_arr_relu_14_31 : IN std_logic ;
      d_arr_relu_14_30 : IN std_logic ;
      d_arr_relu_14_29 : IN std_logic ;
      d_arr_relu_14_28 : IN std_logic ;
      d_arr_relu_14_27 : IN std_logic ;
      d_arr_relu_14_26 : IN std_logic ;
      d_arr_relu_14_25 : IN std_logic ;
      d_arr_relu_14_24 : IN std_logic ;
      d_arr_relu_14_23 : IN std_logic ;
      d_arr_relu_14_22 : IN std_logic ;
      d_arr_relu_14_21 : IN std_logic ;
      d_arr_relu_14_20 : IN std_logic ;
      d_arr_relu_14_19 : IN std_logic ;
      d_arr_relu_14_18 : IN std_logic ;
      d_arr_relu_14_17 : IN std_logic ;
      d_arr_relu_14_16 : IN std_logic ;
      d_arr_relu_14_15 : IN std_logic ;
      d_arr_relu_14_14 : IN std_logic ;
      d_arr_relu_14_13 : IN std_logic ;
      d_arr_relu_14_12 : IN std_logic ;
      d_arr_relu_14_11 : IN std_logic ;
      d_arr_relu_14_10 : IN std_logic ;
      d_arr_relu_14_9 : IN std_logic ;
      d_arr_relu_14_8 : IN std_logic ;
      d_arr_relu_14_7 : IN std_logic ;
      d_arr_relu_14_6 : IN std_logic ;
      d_arr_relu_14_5 : IN std_logic ;
      d_arr_relu_14_4 : IN std_logic ;
      d_arr_relu_14_3 : IN std_logic ;
      d_arr_relu_14_2 : IN std_logic ;
      d_arr_relu_14_1 : IN std_logic ;
      d_arr_relu_14_0 : IN std_logic ;
      d_arr_relu_15_31 : IN std_logic ;
      d_arr_relu_15_30 : IN std_logic ;
      d_arr_relu_15_29 : IN std_logic ;
      d_arr_relu_15_28 : IN std_logic ;
      d_arr_relu_15_27 : IN std_logic ;
      d_arr_relu_15_26 : IN std_logic ;
      d_arr_relu_15_25 : IN std_logic ;
      d_arr_relu_15_24 : IN std_logic ;
      d_arr_relu_15_23 : IN std_logic ;
      d_arr_relu_15_22 : IN std_logic ;
      d_arr_relu_15_21 : IN std_logic ;
      d_arr_relu_15_20 : IN std_logic ;
      d_arr_relu_15_19 : IN std_logic ;
      d_arr_relu_15_18 : IN std_logic ;
      d_arr_relu_15_17 : IN std_logic ;
      d_arr_relu_15_16 : IN std_logic ;
      d_arr_relu_15_15 : IN std_logic ;
      d_arr_relu_15_14 : IN std_logic ;
      d_arr_relu_15_13 : IN std_logic ;
      d_arr_relu_15_12 : IN std_logic ;
      d_arr_relu_15_11 : IN std_logic ;
      d_arr_relu_15_10 : IN std_logic ;
      d_arr_relu_15_9 : IN std_logic ;
      d_arr_relu_15_8 : IN std_logic ;
      d_arr_relu_15_7 : IN std_logic ;
      d_arr_relu_15_6 : IN std_logic ;
      d_arr_relu_15_5 : IN std_logic ;
      d_arr_relu_15_4 : IN std_logic ;
      d_arr_relu_15_3 : IN std_logic ;
      d_arr_relu_15_2 : IN std_logic ;
      d_arr_relu_15_1 : IN std_logic ;
      d_arr_relu_15_0 : IN std_logic ;
      d_arr_relu_16_31 : IN std_logic ;
      d_arr_relu_16_30 : IN std_logic ;
      d_arr_relu_16_29 : IN std_logic ;
      d_arr_relu_16_28 : IN std_logic ;
      d_arr_relu_16_27 : IN std_logic ;
      d_arr_relu_16_26 : IN std_logic ;
      d_arr_relu_16_25 : IN std_logic ;
      d_arr_relu_16_24 : IN std_logic ;
      d_arr_relu_16_23 : IN std_logic ;
      d_arr_relu_16_22 : IN std_logic ;
      d_arr_relu_16_21 : IN std_logic ;
      d_arr_relu_16_20 : IN std_logic ;
      d_arr_relu_16_19 : IN std_logic ;
      d_arr_relu_16_18 : IN std_logic ;
      d_arr_relu_16_17 : IN std_logic ;
      d_arr_relu_16_16 : IN std_logic ;
      d_arr_relu_16_15 : IN std_logic ;
      d_arr_relu_16_14 : IN std_logic ;
      d_arr_relu_16_13 : IN std_logic ;
      d_arr_relu_16_12 : IN std_logic ;
      d_arr_relu_16_11 : IN std_logic ;
      d_arr_relu_16_10 : IN std_logic ;
      d_arr_relu_16_9 : IN std_logic ;
      d_arr_relu_16_8 : IN std_logic ;
      d_arr_relu_16_7 : IN std_logic ;
      d_arr_relu_16_6 : IN std_logic ;
      d_arr_relu_16_5 : IN std_logic ;
      d_arr_relu_16_4 : IN std_logic ;
      d_arr_relu_16_3 : IN std_logic ;
      d_arr_relu_16_2 : IN std_logic ;
      d_arr_relu_16_1 : IN std_logic ;
      d_arr_relu_16_0 : IN std_logic ;
      d_arr_relu_17_31 : IN std_logic ;
      d_arr_relu_17_30 : IN std_logic ;
      d_arr_relu_17_29 : IN std_logic ;
      d_arr_relu_17_28 : IN std_logic ;
      d_arr_relu_17_27 : IN std_logic ;
      d_arr_relu_17_26 : IN std_logic ;
      d_arr_relu_17_25 : IN std_logic ;
      d_arr_relu_17_24 : IN std_logic ;
      d_arr_relu_17_23 : IN std_logic ;
      d_arr_relu_17_22 : IN std_logic ;
      d_arr_relu_17_21 : IN std_logic ;
      d_arr_relu_17_20 : IN std_logic ;
      d_arr_relu_17_19 : IN std_logic ;
      d_arr_relu_17_18 : IN std_logic ;
      d_arr_relu_17_17 : IN std_logic ;
      d_arr_relu_17_16 : IN std_logic ;
      d_arr_relu_17_15 : IN std_logic ;
      d_arr_relu_17_14 : IN std_logic ;
      d_arr_relu_17_13 : IN std_logic ;
      d_arr_relu_17_12 : IN std_logic ;
      d_arr_relu_17_11 : IN std_logic ;
      d_arr_relu_17_10 : IN std_logic ;
      d_arr_relu_17_9 : IN std_logic ;
      d_arr_relu_17_8 : IN std_logic ;
      d_arr_relu_17_7 : IN std_logic ;
      d_arr_relu_17_6 : IN std_logic ;
      d_arr_relu_17_5 : IN std_logic ;
      d_arr_relu_17_4 : IN std_logic ;
      d_arr_relu_17_3 : IN std_logic ;
      d_arr_relu_17_2 : IN std_logic ;
      d_arr_relu_17_1 : IN std_logic ;
      d_arr_relu_17_0 : IN std_logic ;
      d_arr_relu_18_31 : IN std_logic ;
      d_arr_relu_18_30 : IN std_logic ;
      d_arr_relu_18_29 : IN std_logic ;
      d_arr_relu_18_28 : IN std_logic ;
      d_arr_relu_18_27 : IN std_logic ;
      d_arr_relu_18_26 : IN std_logic ;
      d_arr_relu_18_25 : IN std_logic ;
      d_arr_relu_18_24 : IN std_logic ;
      d_arr_relu_18_23 : IN std_logic ;
      d_arr_relu_18_22 : IN std_logic ;
      d_arr_relu_18_21 : IN std_logic ;
      d_arr_relu_18_20 : IN std_logic ;
      d_arr_relu_18_19 : IN std_logic ;
      d_arr_relu_18_18 : IN std_logic ;
      d_arr_relu_18_17 : IN std_logic ;
      d_arr_relu_18_16 : IN std_logic ;
      d_arr_relu_18_15 : IN std_logic ;
      d_arr_relu_18_14 : IN std_logic ;
      d_arr_relu_18_13 : IN std_logic ;
      d_arr_relu_18_12 : IN std_logic ;
      d_arr_relu_18_11 : IN std_logic ;
      d_arr_relu_18_10 : IN std_logic ;
      d_arr_relu_18_9 : IN std_logic ;
      d_arr_relu_18_8 : IN std_logic ;
      d_arr_relu_18_7 : IN std_logic ;
      d_arr_relu_18_6 : IN std_logic ;
      d_arr_relu_18_5 : IN std_logic ;
      d_arr_relu_18_4 : IN std_logic ;
      d_arr_relu_18_3 : IN std_logic ;
      d_arr_relu_18_2 : IN std_logic ;
      d_arr_relu_18_1 : IN std_logic ;
      d_arr_relu_18_0 : IN std_logic ;
      d_arr_relu_19_31 : IN std_logic ;
      d_arr_relu_19_30 : IN std_logic ;
      d_arr_relu_19_29 : IN std_logic ;
      d_arr_relu_19_28 : IN std_logic ;
      d_arr_relu_19_27 : IN std_logic ;
      d_arr_relu_19_26 : IN std_logic ;
      d_arr_relu_19_25 : IN std_logic ;
      d_arr_relu_19_24 : IN std_logic ;
      d_arr_relu_19_23 : IN std_logic ;
      d_arr_relu_19_22 : IN std_logic ;
      d_arr_relu_19_21 : IN std_logic ;
      d_arr_relu_19_20 : IN std_logic ;
      d_arr_relu_19_19 : IN std_logic ;
      d_arr_relu_19_18 : IN std_logic ;
      d_arr_relu_19_17 : IN std_logic ;
      d_arr_relu_19_16 : IN std_logic ;
      d_arr_relu_19_15 : IN std_logic ;
      d_arr_relu_19_14 : IN std_logic ;
      d_arr_relu_19_13 : IN std_logic ;
      d_arr_relu_19_12 : IN std_logic ;
      d_arr_relu_19_11 : IN std_logic ;
      d_arr_relu_19_10 : IN std_logic ;
      d_arr_relu_19_9 : IN std_logic ;
      d_arr_relu_19_8 : IN std_logic ;
      d_arr_relu_19_7 : IN std_logic ;
      d_arr_relu_19_6 : IN std_logic ;
      d_arr_relu_19_5 : IN std_logic ;
      d_arr_relu_19_4 : IN std_logic ;
      d_arr_relu_19_3 : IN std_logic ;
      d_arr_relu_19_2 : IN std_logic ;
      d_arr_relu_19_1 : IN std_logic ;
      d_arr_relu_19_0 : IN std_logic ;
      d_arr_relu_20_31 : IN std_logic ;
      d_arr_relu_20_30 : IN std_logic ;
      d_arr_relu_20_29 : IN std_logic ;
      d_arr_relu_20_28 : IN std_logic ;
      d_arr_relu_20_27 : IN std_logic ;
      d_arr_relu_20_26 : IN std_logic ;
      d_arr_relu_20_25 : IN std_logic ;
      d_arr_relu_20_24 : IN std_logic ;
      d_arr_relu_20_23 : IN std_logic ;
      d_arr_relu_20_22 : IN std_logic ;
      d_arr_relu_20_21 : IN std_logic ;
      d_arr_relu_20_20 : IN std_logic ;
      d_arr_relu_20_19 : IN std_logic ;
      d_arr_relu_20_18 : IN std_logic ;
      d_arr_relu_20_17 : IN std_logic ;
      d_arr_relu_20_16 : IN std_logic ;
      d_arr_relu_20_15 : IN std_logic ;
      d_arr_relu_20_14 : IN std_logic ;
      d_arr_relu_20_13 : IN std_logic ;
      d_arr_relu_20_12 : IN std_logic ;
      d_arr_relu_20_11 : IN std_logic ;
      d_arr_relu_20_10 : IN std_logic ;
      d_arr_relu_20_9 : IN std_logic ;
      d_arr_relu_20_8 : IN std_logic ;
      d_arr_relu_20_7 : IN std_logic ;
      d_arr_relu_20_6 : IN std_logic ;
      d_arr_relu_20_5 : IN std_logic ;
      d_arr_relu_20_4 : IN std_logic ;
      d_arr_relu_20_3 : IN std_logic ;
      d_arr_relu_20_2 : IN std_logic ;
      d_arr_relu_20_1 : IN std_logic ;
      d_arr_relu_20_0 : IN std_logic ;
      d_arr_relu_21_31 : IN std_logic ;
      d_arr_relu_21_30 : IN std_logic ;
      d_arr_relu_21_29 : IN std_logic ;
      d_arr_relu_21_28 : IN std_logic ;
      d_arr_relu_21_27 : IN std_logic ;
      d_arr_relu_21_26 : IN std_logic ;
      d_arr_relu_21_25 : IN std_logic ;
      d_arr_relu_21_24 : IN std_logic ;
      d_arr_relu_21_23 : IN std_logic ;
      d_arr_relu_21_22 : IN std_logic ;
      d_arr_relu_21_21 : IN std_logic ;
      d_arr_relu_21_20 : IN std_logic ;
      d_arr_relu_21_19 : IN std_logic ;
      d_arr_relu_21_18 : IN std_logic ;
      d_arr_relu_21_17 : IN std_logic ;
      d_arr_relu_21_16 : IN std_logic ;
      d_arr_relu_21_15 : IN std_logic ;
      d_arr_relu_21_14 : IN std_logic ;
      d_arr_relu_21_13 : IN std_logic ;
      d_arr_relu_21_12 : IN std_logic ;
      d_arr_relu_21_11 : IN std_logic ;
      d_arr_relu_21_10 : IN std_logic ;
      d_arr_relu_21_9 : IN std_logic ;
      d_arr_relu_21_8 : IN std_logic ;
      d_arr_relu_21_7 : IN std_logic ;
      d_arr_relu_21_6 : IN std_logic ;
      d_arr_relu_21_5 : IN std_logic ;
      d_arr_relu_21_4 : IN std_logic ;
      d_arr_relu_21_3 : IN std_logic ;
      d_arr_relu_21_2 : IN std_logic ;
      d_arr_relu_21_1 : IN std_logic ;
      d_arr_relu_21_0 : IN std_logic ;
      d_arr_relu_22_31 : IN std_logic ;
      d_arr_relu_22_30 : IN std_logic ;
      d_arr_relu_22_29 : IN std_logic ;
      d_arr_relu_22_28 : IN std_logic ;
      d_arr_relu_22_27 : IN std_logic ;
      d_arr_relu_22_26 : IN std_logic ;
      d_arr_relu_22_25 : IN std_logic ;
      d_arr_relu_22_24 : IN std_logic ;
      d_arr_relu_22_23 : IN std_logic ;
      d_arr_relu_22_22 : IN std_logic ;
      d_arr_relu_22_21 : IN std_logic ;
      d_arr_relu_22_20 : IN std_logic ;
      d_arr_relu_22_19 : IN std_logic ;
      d_arr_relu_22_18 : IN std_logic ;
      d_arr_relu_22_17 : IN std_logic ;
      d_arr_relu_22_16 : IN std_logic ;
      d_arr_relu_22_15 : IN std_logic ;
      d_arr_relu_22_14 : IN std_logic ;
      d_arr_relu_22_13 : IN std_logic ;
      d_arr_relu_22_12 : IN std_logic ;
      d_arr_relu_22_11 : IN std_logic ;
      d_arr_relu_22_10 : IN std_logic ;
      d_arr_relu_22_9 : IN std_logic ;
      d_arr_relu_22_8 : IN std_logic ;
      d_arr_relu_22_7 : IN std_logic ;
      d_arr_relu_22_6 : IN std_logic ;
      d_arr_relu_22_5 : IN std_logic ;
      d_arr_relu_22_4 : IN std_logic ;
      d_arr_relu_22_3 : IN std_logic ;
      d_arr_relu_22_2 : IN std_logic ;
      d_arr_relu_22_1 : IN std_logic ;
      d_arr_relu_22_0 : IN std_logic ;
      d_arr_relu_23_31 : IN std_logic ;
      d_arr_relu_23_30 : IN std_logic ;
      d_arr_relu_23_29 : IN std_logic ;
      d_arr_relu_23_28 : IN std_logic ;
      d_arr_relu_23_27 : IN std_logic ;
      d_arr_relu_23_26 : IN std_logic ;
      d_arr_relu_23_25 : IN std_logic ;
      d_arr_relu_23_24 : IN std_logic ;
      d_arr_relu_23_23 : IN std_logic ;
      d_arr_relu_23_22 : IN std_logic ;
      d_arr_relu_23_21 : IN std_logic ;
      d_arr_relu_23_20 : IN std_logic ;
      d_arr_relu_23_19 : IN std_logic ;
      d_arr_relu_23_18 : IN std_logic ;
      d_arr_relu_23_17 : IN std_logic ;
      d_arr_relu_23_16 : IN std_logic ;
      d_arr_relu_23_15 : IN std_logic ;
      d_arr_relu_23_14 : IN std_logic ;
      d_arr_relu_23_13 : IN std_logic ;
      d_arr_relu_23_12 : IN std_logic ;
      d_arr_relu_23_11 : IN std_logic ;
      d_arr_relu_23_10 : IN std_logic ;
      d_arr_relu_23_9 : IN std_logic ;
      d_arr_relu_23_8 : IN std_logic ;
      d_arr_relu_23_7 : IN std_logic ;
      d_arr_relu_23_6 : IN std_logic ;
      d_arr_relu_23_5 : IN std_logic ;
      d_arr_relu_23_4 : IN std_logic ;
      d_arr_relu_23_3 : IN std_logic ;
      d_arr_relu_23_2 : IN std_logic ;
      d_arr_relu_23_1 : IN std_logic ;
      d_arr_relu_23_0 : IN std_logic ;
      d_arr_relu_24_31 : IN std_logic ;
      d_arr_relu_24_30 : IN std_logic ;
      d_arr_relu_24_29 : IN std_logic ;
      d_arr_relu_24_28 : IN std_logic ;
      d_arr_relu_24_27 : IN std_logic ;
      d_arr_relu_24_26 : IN std_logic ;
      d_arr_relu_24_25 : IN std_logic ;
      d_arr_relu_24_24 : IN std_logic ;
      d_arr_relu_24_23 : IN std_logic ;
      d_arr_relu_24_22 : IN std_logic ;
      d_arr_relu_24_21 : IN std_logic ;
      d_arr_relu_24_20 : IN std_logic ;
      d_arr_relu_24_19 : IN std_logic ;
      d_arr_relu_24_18 : IN std_logic ;
      d_arr_relu_24_17 : IN std_logic ;
      d_arr_relu_24_16 : IN std_logic ;
      d_arr_relu_24_15 : IN std_logic ;
      d_arr_relu_24_14 : IN std_logic ;
      d_arr_relu_24_13 : IN std_logic ;
      d_arr_relu_24_12 : IN std_logic ;
      d_arr_relu_24_11 : IN std_logic ;
      d_arr_relu_24_10 : IN std_logic ;
      d_arr_relu_24_9 : IN std_logic ;
      d_arr_relu_24_8 : IN std_logic ;
      d_arr_relu_24_7 : IN std_logic ;
      d_arr_relu_24_6 : IN std_logic ;
      d_arr_relu_24_5 : IN std_logic ;
      d_arr_relu_24_4 : IN std_logic ;
      d_arr_relu_24_3 : IN std_logic ;
      d_arr_relu_24_2 : IN std_logic ;
      d_arr_relu_24_1 : IN std_logic ;
      d_arr_relu_24_0 : IN std_logic ;
      sel_mux : IN std_logic ;
      sel_mul : IN std_logic ;
      sel_add : IN std_logic ;
      sel_merge1 : IN std_logic ;
      sel_merge2 : IN std_logic ;
      sel_relu : IN std_logic ;
      d_arr_0_31 : OUT std_logic ;
      d_arr_0_30 : OUT std_logic ;
      d_arr_0_29 : OUT std_logic ;
      d_arr_0_28 : OUT std_logic ;
      d_arr_0_27 : OUT std_logic ;
      d_arr_0_26 : OUT std_logic ;
      d_arr_0_25 : OUT std_logic ;
      d_arr_0_24 : OUT std_logic ;
      d_arr_0_23 : OUT std_logic ;
      d_arr_0_22 : OUT std_logic ;
      d_arr_0_21 : OUT std_logic ;
      d_arr_0_20 : OUT std_logic ;
      d_arr_0_19 : OUT std_logic ;
      d_arr_0_18 : OUT std_logic ;
      d_arr_0_17 : OUT std_logic ;
      d_arr_0_16 : OUT std_logic ;
      d_arr_0_15 : OUT std_logic ;
      d_arr_0_14 : OUT std_logic ;
      d_arr_0_13 : OUT std_logic ;
      d_arr_0_12 : OUT std_logic ;
      d_arr_0_11 : OUT std_logic ;
      d_arr_0_10 : OUT std_logic ;
      d_arr_0_9 : OUT std_logic ;
      d_arr_0_8 : OUT std_logic ;
      d_arr_0_7 : OUT std_logic ;
      d_arr_0_6 : OUT std_logic ;
      d_arr_0_5 : OUT std_logic ;
      d_arr_0_4 : OUT std_logic ;
      d_arr_0_3 : OUT std_logic ;
      d_arr_0_2 : OUT std_logic ;
      d_arr_0_1 : OUT std_logic ;
      d_arr_0_0 : OUT std_logic ;
      d_arr_1_31 : OUT std_logic ;
      d_arr_1_30 : OUT std_logic ;
      d_arr_1_29 : OUT std_logic ;
      d_arr_1_28 : OUT std_logic ;
      d_arr_1_27 : OUT std_logic ;
      d_arr_1_26 : OUT std_logic ;
      d_arr_1_25 : OUT std_logic ;
      d_arr_1_24 : OUT std_logic ;
      d_arr_1_23 : OUT std_logic ;
      d_arr_1_22 : OUT std_logic ;
      d_arr_1_21 : OUT std_logic ;
      d_arr_1_20 : OUT std_logic ;
      d_arr_1_19 : OUT std_logic ;
      d_arr_1_18 : OUT std_logic ;
      d_arr_1_17 : OUT std_logic ;
      d_arr_1_16 : OUT std_logic ;
      d_arr_1_15 : OUT std_logic ;
      d_arr_1_14 : OUT std_logic ;
      d_arr_1_13 : OUT std_logic ;
      d_arr_1_12 : OUT std_logic ;
      d_arr_1_11 : OUT std_logic ;
      d_arr_1_10 : OUT std_logic ;
      d_arr_1_9 : OUT std_logic ;
      d_arr_1_8 : OUT std_logic ;
      d_arr_1_7 : OUT std_logic ;
      d_arr_1_6 : OUT std_logic ;
      d_arr_1_5 : OUT std_logic ;
      d_arr_1_4 : OUT std_logic ;
      d_arr_1_3 : OUT std_logic ;
      d_arr_1_2 : OUT std_logic ;
      d_arr_1_1 : OUT std_logic ;
      d_arr_1_0 : OUT std_logic ;
      d_arr_2_31 : OUT std_logic ;
      d_arr_2_30 : OUT std_logic ;
      d_arr_2_29 : OUT std_logic ;
      d_arr_2_28 : OUT std_logic ;
      d_arr_2_27 : OUT std_logic ;
      d_arr_2_26 : OUT std_logic ;
      d_arr_2_25 : OUT std_logic ;
      d_arr_2_24 : OUT std_logic ;
      d_arr_2_23 : OUT std_logic ;
      d_arr_2_22 : OUT std_logic ;
      d_arr_2_21 : OUT std_logic ;
      d_arr_2_20 : OUT std_logic ;
      d_arr_2_19 : OUT std_logic ;
      d_arr_2_18 : OUT std_logic ;
      d_arr_2_17 : OUT std_logic ;
      d_arr_2_16 : OUT std_logic ;
      d_arr_2_15 : OUT std_logic ;
      d_arr_2_14 : OUT std_logic ;
      d_arr_2_13 : OUT std_logic ;
      d_arr_2_12 : OUT std_logic ;
      d_arr_2_11 : OUT std_logic ;
      d_arr_2_10 : OUT std_logic ;
      d_arr_2_9 : OUT std_logic ;
      d_arr_2_8 : OUT std_logic ;
      d_arr_2_7 : OUT std_logic ;
      d_arr_2_6 : OUT std_logic ;
      d_arr_2_5 : OUT std_logic ;
      d_arr_2_4 : OUT std_logic ;
      d_arr_2_3 : OUT std_logic ;
      d_arr_2_2 : OUT std_logic ;
      d_arr_2_1 : OUT std_logic ;
      d_arr_2_0 : OUT std_logic ;
      d_arr_3_31 : OUT std_logic ;
      d_arr_3_30 : OUT std_logic ;
      d_arr_3_29 : OUT std_logic ;
      d_arr_3_28 : OUT std_logic ;
      d_arr_3_27 : OUT std_logic ;
      d_arr_3_26 : OUT std_logic ;
      d_arr_3_25 : OUT std_logic ;
      d_arr_3_24 : OUT std_logic ;
      d_arr_3_23 : OUT std_logic ;
      d_arr_3_22 : OUT std_logic ;
      d_arr_3_21 : OUT std_logic ;
      d_arr_3_20 : OUT std_logic ;
      d_arr_3_19 : OUT std_logic ;
      d_arr_3_18 : OUT std_logic ;
      d_arr_3_17 : OUT std_logic ;
      d_arr_3_16 : OUT std_logic ;
      d_arr_3_15 : OUT std_logic ;
      d_arr_3_14 : OUT std_logic ;
      d_arr_3_13 : OUT std_logic ;
      d_arr_3_12 : OUT std_logic ;
      d_arr_3_11 : OUT std_logic ;
      d_arr_3_10 : OUT std_logic ;
      d_arr_3_9 : OUT std_logic ;
      d_arr_3_8 : OUT std_logic ;
      d_arr_3_7 : OUT std_logic ;
      d_arr_3_6 : OUT std_logic ;
      d_arr_3_5 : OUT std_logic ;
      d_arr_3_4 : OUT std_logic ;
      d_arr_3_3 : OUT std_logic ;
      d_arr_3_2 : OUT std_logic ;
      d_arr_3_1 : OUT std_logic ;
      d_arr_3_0 : OUT std_logic ;
      d_arr_4_31 : OUT std_logic ;
      d_arr_4_30 : OUT std_logic ;
      d_arr_4_29 : OUT std_logic ;
      d_arr_4_28 : OUT std_logic ;
      d_arr_4_27 : OUT std_logic ;
      d_arr_4_26 : OUT std_logic ;
      d_arr_4_25 : OUT std_logic ;
      d_arr_4_24 : OUT std_logic ;
      d_arr_4_23 : OUT std_logic ;
      d_arr_4_22 : OUT std_logic ;
      d_arr_4_21 : OUT std_logic ;
      d_arr_4_20 : OUT std_logic ;
      d_arr_4_19 : OUT std_logic ;
      d_arr_4_18 : OUT std_logic ;
      d_arr_4_17 : OUT std_logic ;
      d_arr_4_16 : OUT std_logic ;
      d_arr_4_15 : OUT std_logic ;
      d_arr_4_14 : OUT std_logic ;
      d_arr_4_13 : OUT std_logic ;
      d_arr_4_12 : OUT std_logic ;
      d_arr_4_11 : OUT std_logic ;
      d_arr_4_10 : OUT std_logic ;
      d_arr_4_9 : OUT std_logic ;
      d_arr_4_8 : OUT std_logic ;
      d_arr_4_7 : OUT std_logic ;
      d_arr_4_6 : OUT std_logic ;
      d_arr_4_5 : OUT std_logic ;
      d_arr_4_4 : OUT std_logic ;
      d_arr_4_3 : OUT std_logic ;
      d_arr_4_2 : OUT std_logic ;
      d_arr_4_1 : OUT std_logic ;
      d_arr_4_0 : OUT std_logic ;
      d_arr_5_31 : OUT std_logic ;
      d_arr_5_30 : OUT std_logic ;
      d_arr_5_29 : OUT std_logic ;
      d_arr_5_28 : OUT std_logic ;
      d_arr_5_27 : OUT std_logic ;
      d_arr_5_26 : OUT std_logic ;
      d_arr_5_25 : OUT std_logic ;
      d_arr_5_24 : OUT std_logic ;
      d_arr_5_23 : OUT std_logic ;
      d_arr_5_22 : OUT std_logic ;
      d_arr_5_21 : OUT std_logic ;
      d_arr_5_20 : OUT std_logic ;
      d_arr_5_19 : OUT std_logic ;
      d_arr_5_18 : OUT std_logic ;
      d_arr_5_17 : OUT std_logic ;
      d_arr_5_16 : OUT std_logic ;
      d_arr_5_15 : OUT std_logic ;
      d_arr_5_14 : OUT std_logic ;
      d_arr_5_13 : OUT std_logic ;
      d_arr_5_12 : OUT std_logic ;
      d_arr_5_11 : OUT std_logic ;
      d_arr_5_10 : OUT std_logic ;
      d_arr_5_9 : OUT std_logic ;
      d_arr_5_8 : OUT std_logic ;
      d_arr_5_7 : OUT std_logic ;
      d_arr_5_6 : OUT std_logic ;
      d_arr_5_5 : OUT std_logic ;
      d_arr_5_4 : OUT std_logic ;
      d_arr_5_3 : OUT std_logic ;
      d_arr_5_2 : OUT std_logic ;
      d_arr_5_1 : OUT std_logic ;
      d_arr_5_0 : OUT std_logic ;
      d_arr_6_31 : OUT std_logic ;
      d_arr_6_30 : OUT std_logic ;
      d_arr_6_29 : OUT std_logic ;
      d_arr_6_28 : OUT std_logic ;
      d_arr_6_27 : OUT std_logic ;
      d_arr_6_26 : OUT std_logic ;
      d_arr_6_25 : OUT std_logic ;
      d_arr_6_24 : OUT std_logic ;
      d_arr_6_23 : OUT std_logic ;
      d_arr_6_22 : OUT std_logic ;
      d_arr_6_21 : OUT std_logic ;
      d_arr_6_20 : OUT std_logic ;
      d_arr_6_19 : OUT std_logic ;
      d_arr_6_18 : OUT std_logic ;
      d_arr_6_17 : OUT std_logic ;
      d_arr_6_16 : OUT std_logic ;
      d_arr_6_15 : OUT std_logic ;
      d_arr_6_14 : OUT std_logic ;
      d_arr_6_13 : OUT std_logic ;
      d_arr_6_12 : OUT std_logic ;
      d_arr_6_11 : OUT std_logic ;
      d_arr_6_10 : OUT std_logic ;
      d_arr_6_9 : OUT std_logic ;
      d_arr_6_8 : OUT std_logic ;
      d_arr_6_7 : OUT std_logic ;
      d_arr_6_6 : OUT std_logic ;
      d_arr_6_5 : OUT std_logic ;
      d_arr_6_4 : OUT std_logic ;
      d_arr_6_3 : OUT std_logic ;
      d_arr_6_2 : OUT std_logic ;
      d_arr_6_1 : OUT std_logic ;
      d_arr_6_0 : OUT std_logic ;
      d_arr_7_31 : OUT std_logic ;
      d_arr_7_30 : OUT std_logic ;
      d_arr_7_29 : OUT std_logic ;
      d_arr_7_28 : OUT std_logic ;
      d_arr_7_27 : OUT std_logic ;
      d_arr_7_26 : OUT std_logic ;
      d_arr_7_25 : OUT std_logic ;
      d_arr_7_24 : OUT std_logic ;
      d_arr_7_23 : OUT std_logic ;
      d_arr_7_22 : OUT std_logic ;
      d_arr_7_21 : OUT std_logic ;
      d_arr_7_20 : OUT std_logic ;
      d_arr_7_19 : OUT std_logic ;
      d_arr_7_18 : OUT std_logic ;
      d_arr_7_17 : OUT std_logic ;
      d_arr_7_16 : OUT std_logic ;
      d_arr_7_15 : OUT std_logic ;
      d_arr_7_14 : OUT std_logic ;
      d_arr_7_13 : OUT std_logic ;
      d_arr_7_12 : OUT std_logic ;
      d_arr_7_11 : OUT std_logic ;
      d_arr_7_10 : OUT std_logic ;
      d_arr_7_9 : OUT std_logic ;
      d_arr_7_8 : OUT std_logic ;
      d_arr_7_7 : OUT std_logic ;
      d_arr_7_6 : OUT std_logic ;
      d_arr_7_5 : OUT std_logic ;
      d_arr_7_4 : OUT std_logic ;
      d_arr_7_3 : OUT std_logic ;
      d_arr_7_2 : OUT std_logic ;
      d_arr_7_1 : OUT std_logic ;
      d_arr_7_0 : OUT std_logic ;
      d_arr_8_31 : OUT std_logic ;
      d_arr_8_30 : OUT std_logic ;
      d_arr_8_29 : OUT std_logic ;
      d_arr_8_28 : OUT std_logic ;
      d_arr_8_27 : OUT std_logic ;
      d_arr_8_26 : OUT std_logic ;
      d_arr_8_25 : OUT std_logic ;
      d_arr_8_24 : OUT std_logic ;
      d_arr_8_23 : OUT std_logic ;
      d_arr_8_22 : OUT std_logic ;
      d_arr_8_21 : OUT std_logic ;
      d_arr_8_20 : OUT std_logic ;
      d_arr_8_19 : OUT std_logic ;
      d_arr_8_18 : OUT std_logic ;
      d_arr_8_17 : OUT std_logic ;
      d_arr_8_16 : OUT std_logic ;
      d_arr_8_15 : OUT std_logic ;
      d_arr_8_14 : OUT std_logic ;
      d_arr_8_13 : OUT std_logic ;
      d_arr_8_12 : OUT std_logic ;
      d_arr_8_11 : OUT std_logic ;
      d_arr_8_10 : OUT std_logic ;
      d_arr_8_9 : OUT std_logic ;
      d_arr_8_8 : OUT std_logic ;
      d_arr_8_7 : OUT std_logic ;
      d_arr_8_6 : OUT std_logic ;
      d_arr_8_5 : OUT std_logic ;
      d_arr_8_4 : OUT std_logic ;
      d_arr_8_3 : OUT std_logic ;
      d_arr_8_2 : OUT std_logic ;
      d_arr_8_1 : OUT std_logic ;
      d_arr_8_0 : OUT std_logic ;
      d_arr_9_31 : OUT std_logic ;
      d_arr_9_30 : OUT std_logic ;
      d_arr_9_29 : OUT std_logic ;
      d_arr_9_28 : OUT std_logic ;
      d_arr_9_27 : OUT std_logic ;
      d_arr_9_26 : OUT std_logic ;
      d_arr_9_25 : OUT std_logic ;
      d_arr_9_24 : OUT std_logic ;
      d_arr_9_23 : OUT std_logic ;
      d_arr_9_22 : OUT std_logic ;
      d_arr_9_21 : OUT std_logic ;
      d_arr_9_20 : OUT std_logic ;
      d_arr_9_19 : OUT std_logic ;
      d_arr_9_18 : OUT std_logic ;
      d_arr_9_17 : OUT std_logic ;
      d_arr_9_16 : OUT std_logic ;
      d_arr_9_15 : OUT std_logic ;
      d_arr_9_14 : OUT std_logic ;
      d_arr_9_13 : OUT std_logic ;
      d_arr_9_12 : OUT std_logic ;
      d_arr_9_11 : OUT std_logic ;
      d_arr_9_10 : OUT std_logic ;
      d_arr_9_9 : OUT std_logic ;
      d_arr_9_8 : OUT std_logic ;
      d_arr_9_7 : OUT std_logic ;
      d_arr_9_6 : OUT std_logic ;
      d_arr_9_5 : OUT std_logic ;
      d_arr_9_4 : OUT std_logic ;
      d_arr_9_3 : OUT std_logic ;
      d_arr_9_2 : OUT std_logic ;
      d_arr_9_1 : OUT std_logic ;
      d_arr_9_0 : OUT std_logic ;
      d_arr_10_31 : OUT std_logic ;
      d_arr_10_30 : OUT std_logic ;
      d_arr_10_29 : OUT std_logic ;
      d_arr_10_28 : OUT std_logic ;
      d_arr_10_27 : OUT std_logic ;
      d_arr_10_26 : OUT std_logic ;
      d_arr_10_25 : OUT std_logic ;
      d_arr_10_24 : OUT std_logic ;
      d_arr_10_23 : OUT std_logic ;
      d_arr_10_22 : OUT std_logic ;
      d_arr_10_21 : OUT std_logic ;
      d_arr_10_20 : OUT std_logic ;
      d_arr_10_19 : OUT std_logic ;
      d_arr_10_18 : OUT std_logic ;
      d_arr_10_17 : OUT std_logic ;
      d_arr_10_16 : OUT std_logic ;
      d_arr_10_15 : OUT std_logic ;
      d_arr_10_14 : OUT std_logic ;
      d_arr_10_13 : OUT std_logic ;
      d_arr_10_12 : OUT std_logic ;
      d_arr_10_11 : OUT std_logic ;
      d_arr_10_10 : OUT std_logic ;
      d_arr_10_9 : OUT std_logic ;
      d_arr_10_8 : OUT std_logic ;
      d_arr_10_7 : OUT std_logic ;
      d_arr_10_6 : OUT std_logic ;
      d_arr_10_5 : OUT std_logic ;
      d_arr_10_4 : OUT std_logic ;
      d_arr_10_3 : OUT std_logic ;
      d_arr_10_2 : OUT std_logic ;
      d_arr_10_1 : OUT std_logic ;
      d_arr_10_0 : OUT std_logic ;
      d_arr_11_31 : OUT std_logic ;
      d_arr_11_30 : OUT std_logic ;
      d_arr_11_29 : OUT std_logic ;
      d_arr_11_28 : OUT std_logic ;
      d_arr_11_27 : OUT std_logic ;
      d_arr_11_26 : OUT std_logic ;
      d_arr_11_25 : OUT std_logic ;
      d_arr_11_24 : OUT std_logic ;
      d_arr_11_23 : OUT std_logic ;
      d_arr_11_22 : OUT std_logic ;
      d_arr_11_21 : OUT std_logic ;
      d_arr_11_20 : OUT std_logic ;
      d_arr_11_19 : OUT std_logic ;
      d_arr_11_18 : OUT std_logic ;
      d_arr_11_17 : OUT std_logic ;
      d_arr_11_16 : OUT std_logic ;
      d_arr_11_15 : OUT std_logic ;
      d_arr_11_14 : OUT std_logic ;
      d_arr_11_13 : OUT std_logic ;
      d_arr_11_12 : OUT std_logic ;
      d_arr_11_11 : OUT std_logic ;
      d_arr_11_10 : OUT std_logic ;
      d_arr_11_9 : OUT std_logic ;
      d_arr_11_8 : OUT std_logic ;
      d_arr_11_7 : OUT std_logic ;
      d_arr_11_6 : OUT std_logic ;
      d_arr_11_5 : OUT std_logic ;
      d_arr_11_4 : OUT std_logic ;
      d_arr_11_3 : OUT std_logic ;
      d_arr_11_2 : OUT std_logic ;
      d_arr_11_1 : OUT std_logic ;
      d_arr_11_0 : OUT std_logic ;
      d_arr_12_31 : OUT std_logic ;
      d_arr_12_30 : OUT std_logic ;
      d_arr_12_29 : OUT std_logic ;
      d_arr_12_28 : OUT std_logic ;
      d_arr_12_27 : OUT std_logic ;
      d_arr_12_26 : OUT std_logic ;
      d_arr_12_25 : OUT std_logic ;
      d_arr_12_24 : OUT std_logic ;
      d_arr_12_23 : OUT std_logic ;
      d_arr_12_22 : OUT std_logic ;
      d_arr_12_21 : OUT std_logic ;
      d_arr_12_20 : OUT std_logic ;
      d_arr_12_19 : OUT std_logic ;
      d_arr_12_18 : OUT std_logic ;
      d_arr_12_17 : OUT std_logic ;
      d_arr_12_16 : OUT std_logic ;
      d_arr_12_15 : OUT std_logic ;
      d_arr_12_14 : OUT std_logic ;
      d_arr_12_13 : OUT std_logic ;
      d_arr_12_12 : OUT std_logic ;
      d_arr_12_11 : OUT std_logic ;
      d_arr_12_10 : OUT std_logic ;
      d_arr_12_9 : OUT std_logic ;
      d_arr_12_8 : OUT std_logic ;
      d_arr_12_7 : OUT std_logic ;
      d_arr_12_6 : OUT std_logic ;
      d_arr_12_5 : OUT std_logic ;
      d_arr_12_4 : OUT std_logic ;
      d_arr_12_3 : OUT std_logic ;
      d_arr_12_2 : OUT std_logic ;
      d_arr_12_1 : OUT std_logic ;
      d_arr_12_0 : OUT std_logic ;
      d_arr_13_31 : OUT std_logic ;
      d_arr_13_30 : OUT std_logic ;
      d_arr_13_29 : OUT std_logic ;
      d_arr_13_28 : OUT std_logic ;
      d_arr_13_27 : OUT std_logic ;
      d_arr_13_26 : OUT std_logic ;
      d_arr_13_25 : OUT std_logic ;
      d_arr_13_24 : OUT std_logic ;
      d_arr_13_23 : OUT std_logic ;
      d_arr_13_22 : OUT std_logic ;
      d_arr_13_21 : OUT std_logic ;
      d_arr_13_20 : OUT std_logic ;
      d_arr_13_19 : OUT std_logic ;
      d_arr_13_18 : OUT std_logic ;
      d_arr_13_17 : OUT std_logic ;
      d_arr_13_16 : OUT std_logic ;
      d_arr_13_15 : OUT std_logic ;
      d_arr_13_14 : OUT std_logic ;
      d_arr_13_13 : OUT std_logic ;
      d_arr_13_12 : OUT std_logic ;
      d_arr_13_11 : OUT std_logic ;
      d_arr_13_10 : OUT std_logic ;
      d_arr_13_9 : OUT std_logic ;
      d_arr_13_8 : OUT std_logic ;
      d_arr_13_7 : OUT std_logic ;
      d_arr_13_6 : OUT std_logic ;
      d_arr_13_5 : OUT std_logic ;
      d_arr_13_4 : OUT std_logic ;
      d_arr_13_3 : OUT std_logic ;
      d_arr_13_2 : OUT std_logic ;
      d_arr_13_1 : OUT std_logic ;
      d_arr_13_0 : OUT std_logic ;
      d_arr_14_31 : OUT std_logic ;
      d_arr_14_30 : OUT std_logic ;
      d_arr_14_29 : OUT std_logic ;
      d_arr_14_28 : OUT std_logic ;
      d_arr_14_27 : OUT std_logic ;
      d_arr_14_26 : OUT std_logic ;
      d_arr_14_25 : OUT std_logic ;
      d_arr_14_24 : OUT std_logic ;
      d_arr_14_23 : OUT std_logic ;
      d_arr_14_22 : OUT std_logic ;
      d_arr_14_21 : OUT std_logic ;
      d_arr_14_20 : OUT std_logic ;
      d_arr_14_19 : OUT std_logic ;
      d_arr_14_18 : OUT std_logic ;
      d_arr_14_17 : OUT std_logic ;
      d_arr_14_16 : OUT std_logic ;
      d_arr_14_15 : OUT std_logic ;
      d_arr_14_14 : OUT std_logic ;
      d_arr_14_13 : OUT std_logic ;
      d_arr_14_12 : OUT std_logic ;
      d_arr_14_11 : OUT std_logic ;
      d_arr_14_10 : OUT std_logic ;
      d_arr_14_9 : OUT std_logic ;
      d_arr_14_8 : OUT std_logic ;
      d_arr_14_7 : OUT std_logic ;
      d_arr_14_6 : OUT std_logic ;
      d_arr_14_5 : OUT std_logic ;
      d_arr_14_4 : OUT std_logic ;
      d_arr_14_3 : OUT std_logic ;
      d_arr_14_2 : OUT std_logic ;
      d_arr_14_1 : OUT std_logic ;
      d_arr_14_0 : OUT std_logic ;
      d_arr_15_31 : OUT std_logic ;
      d_arr_15_30 : OUT std_logic ;
      d_arr_15_29 : OUT std_logic ;
      d_arr_15_28 : OUT std_logic ;
      d_arr_15_27 : OUT std_logic ;
      d_arr_15_26 : OUT std_logic ;
      d_arr_15_25 : OUT std_logic ;
      d_arr_15_24 : OUT std_logic ;
      d_arr_15_23 : OUT std_logic ;
      d_arr_15_22 : OUT std_logic ;
      d_arr_15_21 : OUT std_logic ;
      d_arr_15_20 : OUT std_logic ;
      d_arr_15_19 : OUT std_logic ;
      d_arr_15_18 : OUT std_logic ;
      d_arr_15_17 : OUT std_logic ;
      d_arr_15_16 : OUT std_logic ;
      d_arr_15_15 : OUT std_logic ;
      d_arr_15_14 : OUT std_logic ;
      d_arr_15_13 : OUT std_logic ;
      d_arr_15_12 : OUT std_logic ;
      d_arr_15_11 : OUT std_logic ;
      d_arr_15_10 : OUT std_logic ;
      d_arr_15_9 : OUT std_logic ;
      d_arr_15_8 : OUT std_logic ;
      d_arr_15_7 : OUT std_logic ;
      d_arr_15_6 : OUT std_logic ;
      d_arr_15_5 : OUT std_logic ;
      d_arr_15_4 : OUT std_logic ;
      d_arr_15_3 : OUT std_logic ;
      d_arr_15_2 : OUT std_logic ;
      d_arr_15_1 : OUT std_logic ;
      d_arr_15_0 : OUT std_logic ;
      d_arr_16_31 : OUT std_logic ;
      d_arr_16_30 : OUT std_logic ;
      d_arr_16_29 : OUT std_logic ;
      d_arr_16_28 : OUT std_logic ;
      d_arr_16_27 : OUT std_logic ;
      d_arr_16_26 : OUT std_logic ;
      d_arr_16_25 : OUT std_logic ;
      d_arr_16_24 : OUT std_logic ;
      d_arr_16_23 : OUT std_logic ;
      d_arr_16_22 : OUT std_logic ;
      d_arr_16_21 : OUT std_logic ;
      d_arr_16_20 : OUT std_logic ;
      d_arr_16_19 : OUT std_logic ;
      d_arr_16_18 : OUT std_logic ;
      d_arr_16_17 : OUT std_logic ;
      d_arr_16_16 : OUT std_logic ;
      d_arr_16_15 : OUT std_logic ;
      d_arr_16_14 : OUT std_logic ;
      d_arr_16_13 : OUT std_logic ;
      d_arr_16_12 : OUT std_logic ;
      d_arr_16_11 : OUT std_logic ;
      d_arr_16_10 : OUT std_logic ;
      d_arr_16_9 : OUT std_logic ;
      d_arr_16_8 : OUT std_logic ;
      d_arr_16_7 : OUT std_logic ;
      d_arr_16_6 : OUT std_logic ;
      d_arr_16_5 : OUT std_logic ;
      d_arr_16_4 : OUT std_logic ;
      d_arr_16_3 : OUT std_logic ;
      d_arr_16_2 : OUT std_logic ;
      d_arr_16_1 : OUT std_logic ;
      d_arr_16_0 : OUT std_logic ;
      d_arr_17_31 : OUT std_logic ;
      d_arr_17_30 : OUT std_logic ;
      d_arr_17_29 : OUT std_logic ;
      d_arr_17_28 : OUT std_logic ;
      d_arr_17_27 : OUT std_logic ;
      d_arr_17_26 : OUT std_logic ;
      d_arr_17_25 : OUT std_logic ;
      d_arr_17_24 : OUT std_logic ;
      d_arr_17_23 : OUT std_logic ;
      d_arr_17_22 : OUT std_logic ;
      d_arr_17_21 : OUT std_logic ;
      d_arr_17_20 : OUT std_logic ;
      d_arr_17_19 : OUT std_logic ;
      d_arr_17_18 : OUT std_logic ;
      d_arr_17_17 : OUT std_logic ;
      d_arr_17_16 : OUT std_logic ;
      d_arr_17_15 : OUT std_logic ;
      d_arr_17_14 : OUT std_logic ;
      d_arr_17_13 : OUT std_logic ;
      d_arr_17_12 : OUT std_logic ;
      d_arr_17_11 : OUT std_logic ;
      d_arr_17_10 : OUT std_logic ;
      d_arr_17_9 : OUT std_logic ;
      d_arr_17_8 : OUT std_logic ;
      d_arr_17_7 : OUT std_logic ;
      d_arr_17_6 : OUT std_logic ;
      d_arr_17_5 : OUT std_logic ;
      d_arr_17_4 : OUT std_logic ;
      d_arr_17_3 : OUT std_logic ;
      d_arr_17_2 : OUT std_logic ;
      d_arr_17_1 : OUT std_logic ;
      d_arr_17_0 : OUT std_logic ;
      d_arr_18_31 : OUT std_logic ;
      d_arr_18_30 : OUT std_logic ;
      d_arr_18_29 : OUT std_logic ;
      d_arr_18_28 : OUT std_logic ;
      d_arr_18_27 : OUT std_logic ;
      d_arr_18_26 : OUT std_logic ;
      d_arr_18_25 : OUT std_logic ;
      d_arr_18_24 : OUT std_logic ;
      d_arr_18_23 : OUT std_logic ;
      d_arr_18_22 : OUT std_logic ;
      d_arr_18_21 : OUT std_logic ;
      d_arr_18_20 : OUT std_logic ;
      d_arr_18_19 : OUT std_logic ;
      d_arr_18_18 : OUT std_logic ;
      d_arr_18_17 : OUT std_logic ;
      d_arr_18_16 : OUT std_logic ;
      d_arr_18_15 : OUT std_logic ;
      d_arr_18_14 : OUT std_logic ;
      d_arr_18_13 : OUT std_logic ;
      d_arr_18_12 : OUT std_logic ;
      d_arr_18_11 : OUT std_logic ;
      d_arr_18_10 : OUT std_logic ;
      d_arr_18_9 : OUT std_logic ;
      d_arr_18_8 : OUT std_logic ;
      d_arr_18_7 : OUT std_logic ;
      d_arr_18_6 : OUT std_logic ;
      d_arr_18_5 : OUT std_logic ;
      d_arr_18_4 : OUT std_logic ;
      d_arr_18_3 : OUT std_logic ;
      d_arr_18_2 : OUT std_logic ;
      d_arr_18_1 : OUT std_logic ;
      d_arr_18_0 : OUT std_logic ;
      d_arr_19_31 : OUT std_logic ;
      d_arr_19_30 : OUT std_logic ;
      d_arr_19_29 : OUT std_logic ;
      d_arr_19_28 : OUT std_logic ;
      d_arr_19_27 : OUT std_logic ;
      d_arr_19_26 : OUT std_logic ;
      d_arr_19_25 : OUT std_logic ;
      d_arr_19_24 : OUT std_logic ;
      d_arr_19_23 : OUT std_logic ;
      d_arr_19_22 : OUT std_logic ;
      d_arr_19_21 : OUT std_logic ;
      d_arr_19_20 : OUT std_logic ;
      d_arr_19_19 : OUT std_logic ;
      d_arr_19_18 : OUT std_logic ;
      d_arr_19_17 : OUT std_logic ;
      d_arr_19_16 : OUT std_logic ;
      d_arr_19_15 : OUT std_logic ;
      d_arr_19_14 : OUT std_logic ;
      d_arr_19_13 : OUT std_logic ;
      d_arr_19_12 : OUT std_logic ;
      d_arr_19_11 : OUT std_logic ;
      d_arr_19_10 : OUT std_logic ;
      d_arr_19_9 : OUT std_logic ;
      d_arr_19_8 : OUT std_logic ;
      d_arr_19_7 : OUT std_logic ;
      d_arr_19_6 : OUT std_logic ;
      d_arr_19_5 : OUT std_logic ;
      d_arr_19_4 : OUT std_logic ;
      d_arr_19_3 : OUT std_logic ;
      d_arr_19_2 : OUT std_logic ;
      d_arr_19_1 : OUT std_logic ;
      d_arr_19_0 : OUT std_logic ;
      d_arr_20_31 : OUT std_logic ;
      d_arr_20_30 : OUT std_logic ;
      d_arr_20_29 : OUT std_logic ;
      d_arr_20_28 : OUT std_logic ;
      d_arr_20_27 : OUT std_logic ;
      d_arr_20_26 : OUT std_logic ;
      d_arr_20_25 : OUT std_logic ;
      d_arr_20_24 : OUT std_logic ;
      d_arr_20_23 : OUT std_logic ;
      d_arr_20_22 : OUT std_logic ;
      d_arr_20_21 : OUT std_logic ;
      d_arr_20_20 : OUT std_logic ;
      d_arr_20_19 : OUT std_logic ;
      d_arr_20_18 : OUT std_logic ;
      d_arr_20_17 : OUT std_logic ;
      d_arr_20_16 : OUT std_logic ;
      d_arr_20_15 : OUT std_logic ;
      d_arr_20_14 : OUT std_logic ;
      d_arr_20_13 : OUT std_logic ;
      d_arr_20_12 : OUT std_logic ;
      d_arr_20_11 : OUT std_logic ;
      d_arr_20_10 : OUT std_logic ;
      d_arr_20_9 : OUT std_logic ;
      d_arr_20_8 : OUT std_logic ;
      d_arr_20_7 : OUT std_logic ;
      d_arr_20_6 : OUT std_logic ;
      d_arr_20_5 : OUT std_logic ;
      d_arr_20_4 : OUT std_logic ;
      d_arr_20_3 : OUT std_logic ;
      d_arr_20_2 : OUT std_logic ;
      d_arr_20_1 : OUT std_logic ;
      d_arr_20_0 : OUT std_logic ;
      d_arr_21_31 : OUT std_logic ;
      d_arr_21_30 : OUT std_logic ;
      d_arr_21_29 : OUT std_logic ;
      d_arr_21_28 : OUT std_logic ;
      d_arr_21_27 : OUT std_logic ;
      d_arr_21_26 : OUT std_logic ;
      d_arr_21_25 : OUT std_logic ;
      d_arr_21_24 : OUT std_logic ;
      d_arr_21_23 : OUT std_logic ;
      d_arr_21_22 : OUT std_logic ;
      d_arr_21_21 : OUT std_logic ;
      d_arr_21_20 : OUT std_logic ;
      d_arr_21_19 : OUT std_logic ;
      d_arr_21_18 : OUT std_logic ;
      d_arr_21_17 : OUT std_logic ;
      d_arr_21_16 : OUT std_logic ;
      d_arr_21_15 : OUT std_logic ;
      d_arr_21_14 : OUT std_logic ;
      d_arr_21_13 : OUT std_logic ;
      d_arr_21_12 : OUT std_logic ;
      d_arr_21_11 : OUT std_logic ;
      d_arr_21_10 : OUT std_logic ;
      d_arr_21_9 : OUT std_logic ;
      d_arr_21_8 : OUT std_logic ;
      d_arr_21_7 : OUT std_logic ;
      d_arr_21_6 : OUT std_logic ;
      d_arr_21_5 : OUT std_logic ;
      d_arr_21_4 : OUT std_logic ;
      d_arr_21_3 : OUT std_logic ;
      d_arr_21_2 : OUT std_logic ;
      d_arr_21_1 : OUT std_logic ;
      d_arr_21_0 : OUT std_logic ;
      d_arr_22_31 : OUT std_logic ;
      d_arr_22_30 : OUT std_logic ;
      d_arr_22_29 : OUT std_logic ;
      d_arr_22_28 : OUT std_logic ;
      d_arr_22_27 : OUT std_logic ;
      d_arr_22_26 : OUT std_logic ;
      d_arr_22_25 : OUT std_logic ;
      d_arr_22_24 : OUT std_logic ;
      d_arr_22_23 : OUT std_logic ;
      d_arr_22_22 : OUT std_logic ;
      d_arr_22_21 : OUT std_logic ;
      d_arr_22_20 : OUT std_logic ;
      d_arr_22_19 : OUT std_logic ;
      d_arr_22_18 : OUT std_logic ;
      d_arr_22_17 : OUT std_logic ;
      d_arr_22_16 : OUT std_logic ;
      d_arr_22_15 : OUT std_logic ;
      d_arr_22_14 : OUT std_logic ;
      d_arr_22_13 : OUT std_logic ;
      d_arr_22_12 : OUT std_logic ;
      d_arr_22_11 : OUT std_logic ;
      d_arr_22_10 : OUT std_logic ;
      d_arr_22_9 : OUT std_logic ;
      d_arr_22_8 : OUT std_logic ;
      d_arr_22_7 : OUT std_logic ;
      d_arr_22_6 : OUT std_logic ;
      d_arr_22_5 : OUT std_logic ;
      d_arr_22_4 : OUT std_logic ;
      d_arr_22_3 : OUT std_logic ;
      d_arr_22_2 : OUT std_logic ;
      d_arr_22_1 : OUT std_logic ;
      d_arr_22_0 : OUT std_logic ;
      d_arr_23_31 : OUT std_logic ;
      d_arr_23_30 : OUT std_logic ;
      d_arr_23_29 : OUT std_logic ;
      d_arr_23_28 : OUT std_logic ;
      d_arr_23_27 : OUT std_logic ;
      d_arr_23_26 : OUT std_logic ;
      d_arr_23_25 : OUT std_logic ;
      d_arr_23_24 : OUT std_logic ;
      d_arr_23_23 : OUT std_logic ;
      d_arr_23_22 : OUT std_logic ;
      d_arr_23_21 : OUT std_logic ;
      d_arr_23_20 : OUT std_logic ;
      d_arr_23_19 : OUT std_logic ;
      d_arr_23_18 : OUT std_logic ;
      d_arr_23_17 : OUT std_logic ;
      d_arr_23_16 : OUT std_logic ;
      d_arr_23_15 : OUT std_logic ;
      d_arr_23_14 : OUT std_logic ;
      d_arr_23_13 : OUT std_logic ;
      d_arr_23_12 : OUT std_logic ;
      d_arr_23_11 : OUT std_logic ;
      d_arr_23_10 : OUT std_logic ;
      d_arr_23_9 : OUT std_logic ;
      d_arr_23_8 : OUT std_logic ;
      d_arr_23_7 : OUT std_logic ;
      d_arr_23_6 : OUT std_logic ;
      d_arr_23_5 : OUT std_logic ;
      d_arr_23_4 : OUT std_logic ;
      d_arr_23_3 : OUT std_logic ;
      d_arr_23_2 : OUT std_logic ;
      d_arr_23_1 : OUT std_logic ;
      d_arr_23_0 : OUT std_logic ;
      d_arr_24_31 : OUT std_logic ;
      d_arr_24_30 : OUT std_logic ;
      d_arr_24_29 : OUT std_logic ;
      d_arr_24_28 : OUT std_logic ;
      d_arr_24_27 : OUT std_logic ;
      d_arr_24_26 : OUT std_logic ;
      d_arr_24_25 : OUT std_logic ;
      d_arr_24_24 : OUT std_logic ;
      d_arr_24_23 : OUT std_logic ;
      d_arr_24_22 : OUT std_logic ;
      d_arr_24_21 : OUT std_logic ;
      d_arr_24_20 : OUT std_logic ;
      d_arr_24_19 : OUT std_logic ;
      d_arr_24_18 : OUT std_logic ;
      d_arr_24_17 : OUT std_logic ;
      d_arr_24_16 : OUT std_logic ;
      d_arr_24_15 : OUT std_logic ;
      d_arr_24_14 : OUT std_logic ;
      d_arr_24_13 : OUT std_logic ;
      d_arr_24_12 : OUT std_logic ;
      d_arr_24_11 : OUT std_logic ;
      d_arr_24_10 : OUT std_logic ;
      d_arr_24_9 : OUT std_logic ;
      d_arr_24_8 : OUT std_logic ;
      d_arr_24_7 : OUT std_logic ;
      d_arr_24_6 : OUT std_logic ;
      d_arr_24_5 : OUT std_logic ;
      d_arr_24_4 : OUT std_logic ;
      d_arr_24_3 : OUT std_logic ;
      d_arr_24_2 : OUT std_logic ;
      d_arr_24_1 : OUT std_logic ;
      d_arr_24_0 : OUT std_logic) ;
end CacheMuxer ;

architecture Behavioral_unfold_3297_0 of CacheMuxer is
   signal nx4, nx8, nx12, nx18, nx28, nx36, nx44, nx52, nx60, nx68, nx76, 
      nx84, nx92, nx100, nx108, nx116, nx124, nx132, nx140, nx146, nx152, 
      nx158, nx164, nx170, nx176, nx182, nx188, nx194, nx200, nx206, nx212, 
      nx218, nx224, nx230, nx236, nx244, nx252, nx260, nx268, nx276, nx284, 
      nx292, nx300, nx308, nx316, nx324, nx332, nx340, nx348, nx356, nx364, 
      nx370, nx376, nx382, nx388, nx394, nx400, nx406, nx412, nx418, nx424, 
      nx430, nx436, nx442, nx448, nx454, nx460, nx468, nx476, nx484, nx492, 
      nx500, nx508, nx516, nx524, nx532, nx540, nx548, nx556, nx564, nx572, 
      nx580, nx588, nx594, nx600, nx606, nx612, nx618, nx624, nx630, nx636, 
      nx642, nx648, nx654, nx660, nx666, nx672, nx678, nx684, nx694, nx700, 
      nx712, nx724, nx736, nx748, nx760, nx772, nx784, nx796, nx808, nx820, 
      nx832, nx844, nx856, nx868, nx880, nx890, nx900, nx910, nx920, nx930, 
      nx940, nx950, nx960, nx970, nx980, nx990, nx1000, nx1010, nx1020, 
      nx1030, nx1040, nx1052, nx1064, nx1076, nx1088, nx1100, nx1112, nx1124, 
      nx1136, nx1148, nx1160, nx1172, nx1184, nx1196, nx1208, nx1220, nx1232, 
      nx1242, nx1252, nx1262, nx1272, nx1282, nx1292, nx1302, nx1312, nx1322, 
      nx1332, nx1342, nx1352, nx1362, nx1372, nx1382, nx1392, nx1404, nx1416, 
      nx1428, nx1440, nx1452, nx1464, nx1476, nx1488, nx1500, nx1512, nx1524, 
      nx1536, nx1548, nx1560, nx1572, nx1584, nx1594, nx1604, nx1614, nx1624, 
      nx1634, nx1644, nx1654, nx1664, nx1674, nx1684, nx1694, nx1704, nx1714, 
      nx1724, nx1734, nx1744, nx1756, nx1768, nx1780, nx1792, nx1804, nx1816, 
      nx1828, nx1840, nx1852, nx1864, nx1876, nx1888, nx1900, nx1912, nx1924, 
      nx1936, nx1946, nx1956, nx1966, nx1976, nx1986, nx1996, nx2006, nx2016, 
      nx2026, nx2036, nx2046, nx2056, nx2066, nx2076, nx2086, nx2096, nx2104, 
      nx2112, nx2120, nx2128, nx2136, nx2144, nx2152, nx2160, nx2168, nx2176, 
      nx2184, nx2192, nx2200, nx2208, nx2216, nx2224, nx2232, nx2240, nx2248, 
      nx2256, nx2264, nx2272, nx2280, nx2288, nx2296, nx2304, nx2312, nx2320, 
      nx2328, nx2336, nx2344, nx2352, nx2360, nx2368, nx2376, nx2384, nx2392, 
      nx2400, nx2408, nx2416, nx2424, nx2432, nx2440, nx2448, nx2456, nx2464, 
      nx2472, nx2480, nx2488, nx2496, nx2504, nx2512, nx2520, nx2528, nx2536, 
      nx2544, nx2552, nx2560, nx2568, nx2576, nx2584, nx2592, nx2600, nx2608, 
      nx2616, nx2624, nx2632, nx2640, nx2648, nx2656, nx2664, nx2672, nx2680, 
      nx2688, nx2696, nx2704, nx2712, nx2720, nx2728, nx2736, nx2744, nx2752, 
      nx2760, nx2768, nx2776, nx2784, nx2792, nx2800, nx2808, nx2816, nx2824, 
      nx2832, nx2840, nx2848, nx2856, nx2864, nx2872, nx2880, nx2888, nx2896, 
      nx2904, nx2912, nx2920, nx2928, nx2936, nx2944, nx2952, nx2960, nx2968, 
      nx2976, nx2984, nx2992, nx3000, nx3008, nx3016, nx3024, nx3032, nx3040, 
      nx3048, nx3056, nx3064, nx3072, nx3080, nx3088, nx3096, nx3104, nx3112, 
      nx3120, nx3132, nx3144, nx3156, nx3168, nx3180, nx3192, nx3204, nx3216, 
      nx3228, nx3240, nx3252, nx3264, nx3276, nx3288, nx3300, nx3312, nx3324, 
      nx3336, nx3348, nx3360, nx3372, nx3384, nx3396, nx3408, nx3420, nx3432, 
      nx3444, nx3456, nx3468, nx3480, nx3492, nx3504, nx3516, nx3528, nx3540, 
      nx3552, nx3564, nx3576, nx3588, nx3600, nx3612, nx3624, nx3636, nx3648, 
      nx3660, nx3672, nx3684, nx3696, nx3708, nx3720, nx3732, nx3744, nx3756, 
      nx3768, nx3780, nx3792, nx3804, nx3816, nx3828, nx3840, nx3852, nx3864, 
      nx3876, nx3888, nx3900, nx3912, nx3924, nx3936, nx3948, nx3960, nx3972, 
      nx3984, nx3996, nx4008, nx4020, nx4032, nx4044, nx4056, nx4068, nx4080, 
      nx4092, nx4104, nx4116, nx4128, nx4140, nx4152, nx4164, nx4176, nx4188, 
      nx4200, nx4212, nx4224, nx4236, nx4248, nx4260, nx4272, nx4284, nx4296, 
      nx4308, nx4320, nx4332, nx4344, nx4356, nx4368, nx4380, nx4392, nx4404, 
      nx4416, nx4428, nx4440, nx4452, nx4464, nx4476, nx4488, nx4500, nx4512, 
      nx4524, nx4536, nx4548, nx4560, nx4572, nx4584, nx4596, nx4608, nx4620, 
      nx4632, nx4644, nx4656, nx4668, nx4680, nx4692, nx4704, nx4716, nx4728, 
      nx4740, nx4752, nx4764, nx4776, nx4788, nx4800, nx4812, nx4824, nx4836, 
      nx4848, nx4860, nx4872, nx4884, nx4896, nx4908, nx4920, nx4932, nx4944, 
      nx4956, nx4968, nx4980, nx4992, nx5004, nx5016, nx5028, nx5040, nx5048, 
      nx5056, nx5064, nx5072, nx5080, nx5088, nx5096, nx5104, nx5112, nx5120, 
      nx5128, nx5136, nx5144, nx5152, nx5160, nx5168, nx5174, nx5180, nx5186, 
      nx5192, nx5198, nx5204, nx5210, nx5216, nx5222, nx5228, nx5234, nx5240, 
      nx5246, nx5252, nx5258, nx5264, nx5272, nx5280, nx5288, nx5296, nx5304, 
      nx5312, nx5320, nx5328, nx5336, nx5344, nx5352, nx5360, nx5368, nx5376, 
      nx5384, nx5392, nx5398, nx5404, nx5410, nx5416, nx5422, nx5428, nx5434, 
      nx5440, nx5446, nx5452, nx5458, nx5464, nx5470, nx5476, nx5482, nx5488, 
      nx5496, nx5504, nx5512, nx5520, nx5528, nx5536, nx5544, nx5552, nx5560, 
      nx5568, nx5576, nx5584, nx5592, nx5600, nx5608, nx5616, nx5622, nx5628, 
      nx5634, nx5640, nx5646, nx5652, nx5658, nx5664, nx5670, nx5676, nx5682, 
      nx5688, nx5694, nx5700, nx5706, nx5712, nx5720, nx5728, nx5736, nx5744, 
      nx5752, nx5760, nx5768, nx5776, nx5784, nx5792, nx5800, nx5808, nx5816, 
      nx5824, nx5832, nx5840, nx5846, nx5852, nx5858, nx5864, nx5870, nx5876, 
      nx5882, nx5888, nx5894, nx5900, nx5906, nx5912, nx5918, nx5924, nx5930, 
      nx5936, nx5948, nx5960, nx5972, nx5984, nx5996, nx6008, nx6020, nx6032, 
      nx6044, nx6056, nx6068, nx6080, nx6092, nx6104, nx6116, nx6128, nx6138, 
      nx6148, nx6158, nx6168, nx6178, nx6188, nx6198, nx6208, nx6218, nx6228, 
      nx6238, nx6248, nx6258, nx6268, nx6278, nx6288, nx6300, nx6312, nx6324, 
      nx6336, nx6348, nx6360, nx6372, nx6384, nx6396, nx6408, nx6420, nx6432, 
      nx6444, nx6456, nx6468, nx6480, nx6490, nx6500, nx6510, nx6520, nx6530, 
      nx6540, nx6550, nx6560, nx6570, nx6580, nx6590, nx6600, nx6610, nx6620, 
      nx6630, nx6640, nx6652, nx6664, nx6676, nx6688, nx6700, nx6712, nx6724, 
      nx6736, nx6748, nx6760, nx6772, nx6784, nx6796, nx6808, nx6820, nx6832, 
      nx6842, nx6852, nx6862, nx6872, nx6882, nx6892, nx6902, nx6912, nx6922, 
      nx6932, nx6942, nx6952, nx6962, nx6972, nx6982, nx6992, nx7002, nx7018, 
      nx7028, nx7036, nx7060, nx7084, nx7108, nx7132, nx7156, nx7180, nx7204, 
      nx7228, nx7252, nx7276, nx7300, nx7324, nx7348, nx7372, nx7392, nx7414, 
      nx7436, nx7458, nx7480, nx7502, nx7524, nx7546, nx7568, nx7590, nx7612, 
      nx7634, nx7656, nx7678, nx7700, nx7722, nx7744, nx7768, nx7792, nx7816, 
      nx7840, nx7864, nx7888, nx7912, nx7936, nx7960, nx7984, nx8008, nx8032, 
      nx8056, nx8080, nx8104, nx8124, nx8146, nx8168, nx8190, nx8212, nx8234, 
      nx8256, nx8278, nx8300, nx8322, nx8344, nx8366, nx8388, nx8410, nx8432, 
      nx8454, nx8476, nx7201, nx7205, nx7209, nx7215, nx7221, nx7227, nx7233, 
      nx7239, nx7245, nx7251, nx7257, nx7263, nx7269, nx7275, nx7281, nx7287, 
      nx7293, nx7295, nx7301, nx7305, nx7311, nx7317, nx7323, nx7329, nx7335, 
      nx7341, nx7347, nx7353, nx7359, nx7365, nx7371, nx7377, nx7383, nx7389, 
      nx7395, nx7401, nx7407, nx7413, nx7419, nx7425, nx7431, nx7437, nx7441, 
      nx7447, nx7453, nx7459, nx7463, nx7469, nx7475, nx7481, nx7483, nx7489, 
      nx7495, nx7501, nx7507, nx7513, nx7519, nx7525, nx7529, nx7535, nx7541, 
      nx7547, nx7551, nx7557, nx7563, nx7569, nx7573, nx7579, nx7585, nx7591, 
      nx7595, nx7601, nx7607, nx7613, nx7617, nx7623, nx7629, nx7635, nx7639, 
      nx7645, nx7651, nx7657, nx7661, nx7663, nx7669, nx7675, nx7681, nx7687, 
      nx7693, nx7699, nx7705, nx7711, nx7717, nx7723, nx7727, nx7733, nx7739, 
      nx7745, nx7749, nx7755, nx7761, nx7767, nx7773, nx7779, nx7785, nx7791, 
      nx7797, nx7803, nx7809, nx7815, nx7821, nx7827, nx7833, nx7839, nx7845, 
      nx7851, nx7853, nx7859, nx7865, nx7869, nx7875, nx7881, nx7887, nx7893, 
      nx7899, nx7905, nx7911, nx7917, nx7923, nx7929, nx7935, nx7941, nx7947, 
      nx8423, nx8429, nx8435, nx8441, nx8447, nx8453, nx8459, nx8465, nx8471, 
      nx8477, nx8481, nx8485, nx8489, nx8493, nx8497, nx8501, nx8505, nx8509, 
      nx8513, nx8517, nx8521, nx8525, nx8529, nx8533, nx8537, nx8541, nx8545, 
      nx8549, nx8553, nx8557, nx8561, nx8565, nx8569, nx8573, nx8577, nx8581, 
      nx8585, nx8589, nx8593, nx8597, nx8601, nx8605, nx8609, nx8613, nx8617, 
      nx8621, nx8625, nx8629, nx8633, nx8637, nx8641, nx8645, nx8649, nx8653, 
      nx8657, nx8661, nx8665, nx8669, nx8673, nx8677, nx8681, nx8685, nx8689, 
      nx8693, nx8697, nx8701, nx8705, nx8709, nx8713, nx8717, nx8721, nx8725, 
      nx8729, nx8733, nx8737, nx8741, nx8745, nx8749, nx8753, nx8757, nx8761, 
      nx8765, nx8769, nx8773, nx8777, nx8781, nx8785, nx8789, nx8793, nx8797, 
      nx8801, nx8805, nx8809, nx8813, nx8817, nx8821, nx8825, nx8829, nx8833, 
      nx8837, nx8841, nx8845, nx8849, nx8853, nx8857, nx8861, nx8865, nx8869, 
      nx8873, nx8877, nx8881, nx8885, nx8889, nx8893, nx8897, nx8901, nx8905, 
      nx8909, nx8913, nx8917, nx8921, nx8925, nx8929, nx8933, nx8937, nx8941, 
      nx8945, nx8949, nx8953, nx8957, nx8961, nx8965, nx8969, nx8973, nx8977, 
      nx8981, nx8985, nx8989, nx8993, nx8997, nx9001, nx9005, nx9009, nx9013, 
      nx9017, nx9021, nx9025, nx9029, nx9033, nx9037, nx9041, nx9045, nx9049, 
      nx9053, nx9057, nx9061, nx9065, nx9069, nx9073, nx9077, nx9341, nx9345, 
      nx9349, nx9353, nx9357, nx9361, nx9365, nx9369, nx9373, nx9377, nx9381, 
      nx9385, nx9389, nx9393, nx9397, nx9401, nx9403, nx9407, nx9411, nx9415, 
      nx9419, nx9423, nx9427, nx9431, nx9435, nx9439, nx9443, nx9447, nx9451, 
      nx9455, nx9459, nx9463, nx9467, nx9471, nx9475, nx9479, nx9483, nx9487, 
      nx9491, nx9495, nx9499, nx9503, nx9507, nx9511, nx9515, nx9519, nx9523, 
      nx9527, nx9531, nx9533, nx9537, nx9541, nx9545, nx9549, nx9553, nx9557, 
      nx9561, nx9565, nx9569, nx9573, nx9577, nx9581, nx9585, nx9589, nx9593, 
      nx9597, nx9601, nx9605, nx9609, nx9613, nx9617, nx9621, nx9625, nx9629, 
      nx9633, nx9637, nx9641, nx9645, nx9649, nx9653, nx9657, nx9661, nx9663, 
      nx9667, nx9671, nx9675, nx9679, nx9683, nx9687, nx9691, nx9695, nx9699, 
      nx9703, nx9707, nx9711, nx9715, nx9719, nx9723, nx9727, nx9731, nx9734, 
      nx9737, nx9739, nx9742, nx9746, nx9748, nx9752, nx9754, nx9758, nx9760, 
      nx9764, nx9766, nx9770, nx9772, nx9776, nx9778, nx9782, nx9784, nx9788, 
      nx9790, nx9794, nx9796, nx9800, nx9802, nx9806, nx9808, nx9812, nx9814, 
      nx9818, nx9820, nx9824, nx9826, nx9830, nx9832, nx9834, nx9838, nx9840, 
      nx9844, nx9846, nx9850, nx9852, nx9856, nx9858, nx9862, nx9864, nx9868, 
      nx9870, nx9874, nx9876, nx9880, nx9882, nx9886, nx9888, nx9892, nx9894, 
      nx9898, nx9900, nx9904, nx9906, nx9910, nx9912, nx9916, nx9918, nx9922, 
      nx9924, nx9928, nx9930, nx9934, nx9936, nx9940, nx9942, nx9946, nx9948, 
      nx9952, nx9954, nx9958, nx9960, nx9964, nx9966, nx9970, nx9972, nx9976, 
      nx9978, nx9982, nx9984, nx9988, nx9990, nx9994, nx9996, nx10000, 
      nx10002, nx10006, nx10008, nx10012, nx10014, nx10018, nx10020, nx10024, 
      nx10026, nx10028, nx10032, nx10034, nx10038, nx10040, nx10044, nx10046, 
      nx10050, nx10052, nx10056, nx10058, nx10062, nx10064, nx10068, nx10070, 
      nx10074, nx10076, nx10080, nx10082, nx10086, nx10088, nx10092, nx10094, 
      nx10098, nx10100, nx10104, nx10106, nx10110, nx10112, nx10116, nx10118, 
      nx10122, nx10124, nx10133, nx10135, nx10137, nx10139, nx10141, nx10143, 
      nx10145, nx10147, nx10149, nx10151, nx10153, nx10155, nx10157, nx10159, 
      nx10161, nx10163, nx10165, nx10167, nx10169, nx10171, nx10173, nx10175, 
      nx10177, nx10179, nx10181, nx10183, nx10185, nx10187, nx10189, nx10191, 
      nx10193, nx10195, nx10197, nx10199, nx10201, nx10203, nx10205, nx10207, 
      nx10209, nx10211, nx10213, nx10215, nx10217, nx10219, nx10221, nx10223, 
      nx10225, nx10227, nx10229, nx10231, nx10233, nx10235, nx10237, nx10239, 
      nx10241, nx10243, nx10245, nx10247, nx10249, nx10251, nx10253, nx10255, 
      nx10257, nx10259, nx10261, nx10263, nx10265, nx10267, nx10269, nx10271, 
      nx10273, nx10275, nx10277, nx10279, nx10281, nx10283, nx10285, nx10287, 
      nx10289, nx10291, nx10293, nx10295, nx10297, nx10299, nx10301, nx10303, 
      nx10305, nx10307, nx10309, nx10311, nx10313, nx10315, nx10317, nx10319, 
      nx10321, nx10323, nx10325, nx10327, nx10329, nx10331, nx10333, nx10335, 
      nx10337, nx10339, nx10341, nx10343, nx10345, nx10347, nx10349, nx10351, 
      nx10353, nx10355, nx10357, nx10359, nx10361, nx10365, nx10367, nx10369, 
      nx10373, nx10375, nx10377, nx10383, nx10385, nx10387, nx10391, nx10393, 
      nx10395, nx10397, nx10399, nx10401, nx10403, nx10405, nx10407, nx10409, 
      nx10411, nx10413, nx10415, nx10417, nx10419, nx10421, nx10423, nx10425, 
      nx10427, nx10429, nx10431, nx10433, nx10435, nx10437, nx10439, nx10441, 
      nx10443, nx10445, nx10447, nx10449, nx10451, nx10453, nx10455, nx10457, 
      nx10459, nx10461, nx10463, nx10465, nx10467, nx10469, nx10471, nx10473, 
      nx10475, nx10477, nx10479, nx10481, nx10483, nx10485, nx10487, nx10489, 
      nx10491, nx10493, nx10495, nx10497, nx10499, nx10501, nx10503, nx10505, 
      nx10507, nx10509, nx10511, nx10513, nx10515, nx10519, nx10521, nx10523, 
      nx10529, nx10531, nx10533, nx10537, nx10539, nx10541, nx10547, nx10549, 
      nx10551, nx10553, nx10555, nx10557, nx10559, nx10561, nx10563, nx10565, 
      nx10567, nx10569, nx10571, nx10573, nx10575, nx10577, nx10579, nx10581, 
      nx10583, nx10585, nx10587, nx10589, nx10591, nx10593, nx10595, nx10603, 
      nx10611, nx10621, nx10623, nx10625, nx10627, nx10629, nx10631, nx10633, 
      nx10635, nx10637, nx10639, nx10641, nx10643, nx10645, nx10647, nx10649, 
      nx10651, nx10653, nx10655, nx10657, nx10659, nx10661, nx10663, nx10665, 
      nx10667, nx10669, nx10671, nx10673, nx10675, nx10677, nx10679, nx10681, 
      nx10683, nx10685, nx10687, nx10689, nx10691, nx10693, nx10695, nx10697, 
      nx10699, nx10701, nx10703, nx10705, nx10707, nx10709, nx10711, nx10713, 
      nx10715, nx10717, nx10719, nx10721, nx10723, nx10725, nx10727, nx10729, 
      nx10731, nx10733, nx10735, nx10737, nx10739, nx10741, nx10743, nx10745, 
      nx10747, nx10749, nx10757, nx10765, nx10773, nx10781, nx10783, nx10785, 
      nx10787, nx10789, nx10791, nx10793, nx10795, nx10797, nx10799, nx10801, 
      nx10803, nx10805, nx10807, nx10809, nx10811, nx10813, nx10815, nx10817, 
      nx10819, nx10821, nx10823, nx10825, nx10827, nx10829, nx10831, nx10833, 
      nx10835, nx10837, nx10839, nx10841, nx10843, nx10845, nx10847, nx10849, 
      nx10851, nx10853, nx10855, nx10857, nx10859, nx10861, nx10863, nx10865, 
      nx10867, nx10869, nx10871, nx10873, nx10875, nx10877, nx10879, nx10881, 
      nx10883, nx10885, nx10887, nx10889, nx10891, nx10893, nx10895, nx10897, 
      nx10899, nx10901, nx10903, nx10905, nx10907, nx10909, nx10911, nx10913, 
      nx10915, nx10917, nx10919, nx10921, nx10923, nx10925, nx10927, nx10929, 
      nx10931, nx10933, nx10935, nx10937, nx10939, nx10941, nx10943, nx10945, 
      nx10947, nx10949, nx10951, nx10953, nx10955, nx10957, nx10959, nx10961, 
      nx10963, nx10965, nx10967, nx10969, nx10971, nx10973, nx10979, nx10981, 
      nx10983, nx10985, nx10987, nx10989, nx10991, nx10993, nx10995, nx10997, 
      nx10999, nx11005, nx11007, nx11009, nx11011, nx11013, nx11015, nx11017, 
      nx11019, nx11021, nx11023, nx11025, nx11027, nx11029, nx11031, nx11033, 
      nx11035, nx11037, nx11039, nx11041, nx11043, nx11045, nx11047, nx11049, 
      nx11051, nx11053, nx11055, nx11057, nx11059, nx11061, nx11063, nx11065, 
      nx11067, nx11069, nx11071, nx11073, nx11075, nx11077, nx11079, nx11081, 
      nx11083, nx11085, nx11087, nx11089, nx11091, nx11093, nx11095, nx11097, 
      nx11099, nx11101, nx11103, nx11105, nx11107, nx11109, nx11111, nx11113, 
      nx11115, nx11117, nx11119, nx11121, nx11123, nx11125, nx11127, nx11129, 
      nx11131, nx11133, nx11135, nx11137, nx11139, nx11141, nx11143, nx11145, 
      nx11147, nx11149, nx11151, nx11153, nx11155, nx11157, nx11159, nx11161, 
      nx11163, nx11165, nx11167, nx11169, nx11171, nx11173, nx11175, nx11177, 
      nx11179, nx11181, nx11183, nx11185, nx11187, nx11189, nx11191, nx11193, 
      nx11195, nx11197, nx11199, nx11201, nx11203, nx11205, nx11207, nx11209, 
      nx11211, nx11213, nx11215, nx11217, nx11219, nx11221, nx11223, nx11225, 
      nx11227, nx11229, nx11231, nx11233, nx11235, nx11237, nx11239, nx11241, 
      nx11245, nx11247, nx11249, nx11251, nx11253, nx11255, nx11257, nx11259, 
      nx11261, nx11263, nx11265, nx11267, nx11269, nx11271, nx11273, nx11275, 
      nx11277, nx11279, nx11281, nx11283, nx11285, nx11287, nx11289, nx11291, 
      nx11293, nx11295, nx11297, nx11299, nx11301, nx11303, nx11305, nx11307, 
      nx11309, nx11311, nx11313, nx11315, nx11317, nx11319, nx11321, nx11323, 
      nx11325, nx11327, nx11329, nx11331, nx11333, nx11335, nx11337, nx11339, 
      nx11341, nx11343, nx11345, nx11347, nx11349, nx11351, nx11353, nx11355, 
      nx11357, nx11359, nx11361, nx11363, nx11365, nx11367, nx11369, nx11371, 
      nx11373, nx11375, nx11377, nx11379, nx11381, nx11383, nx11385, nx11387, 
      nx11389, nx11391, nx11393, nx11395, nx11397, nx11399, nx11401, nx11403, 
      nx11405, nx11407, nx11409, nx11411, nx11413, nx11415, nx11417, nx11419, 
      nx11421, nx11423, nx11425, nx11427, nx11429, nx11431, nx11433, nx11435, 
      nx11437, nx11439, nx11441, nx11443, nx11445, nx11447, nx11449, nx11451, 
      nx11453, nx11455, nx11457, nx11459, nx11461, nx11463, nx11465, nx11467, 
      nx11469, nx11471, nx11473, nx11475, nx11477, nx11479, nx11481, nx11483, 
      nx11485, nx11487, nx11489, nx11491, nx11493, nx11495, nx11497, nx11499, 
      nx11501, nx11503, nx11505, nx11511, nx11517, nx11519, nx11524, nx11525
   : std_logic ;

begin
   lat_d_arr_24_0 : latch port map ( Q=>d_arr_24_0, D=>nx18, CLK=>nx10133);
   ix19 : ao22 port map ( Y=>nx18, A0=>d_arr_mux_24_0, A1=>nx11245, B0=>
      d_arr_mul_24_0, B1=>nx10365);
   ix13 : nor02ii port map ( Y=>nx12, A0=>nx11245, A1=>sel_mul);
   ix9 : or03 port map ( Y=>nx8, A0=>sel_merge2, A1=>sel_relu, A2=>nx4);
   lat_d_arr_24_1 : latch port map ( Q=>d_arr_24_1, D=>nx28, CLK=>nx10133);
   ix29 : ao22 port map ( Y=>nx28, A0=>d_arr_mux_24_1, A1=>nx11245, B0=>
      d_arr_mul_24_1, B1=>nx10365);
   lat_d_arr_24_2 : latch port map ( Q=>d_arr_24_2, D=>nx36, CLK=>nx10133);
   ix37 : ao22 port map ( Y=>nx36, A0=>d_arr_mux_24_2, A1=>nx11245, B0=>
      d_arr_mul_24_2, B1=>nx10365);
   lat_d_arr_24_3 : latch port map ( Q=>d_arr_24_3, D=>nx44, CLK=>nx10133);
   ix45 : ao22 port map ( Y=>nx44, A0=>d_arr_mux_24_3, A1=>nx11245, B0=>
      d_arr_mul_24_3, B1=>nx10365);
   lat_d_arr_24_4 : latch port map ( Q=>d_arr_24_4, D=>nx52, CLK=>nx10133);
   ix53 : ao22 port map ( Y=>nx52, A0=>d_arr_mux_24_4, A1=>nx11245, B0=>
      d_arr_mul_24_4, B1=>nx10365);
   lat_d_arr_24_5 : latch port map ( Q=>d_arr_24_5, D=>nx60, CLK=>nx10133);
   ix61 : ao22 port map ( Y=>nx60, A0=>d_arr_mux_24_5, A1=>nx11245, B0=>
      d_arr_mul_24_5, B1=>nx10365);
   lat_d_arr_24_6 : latch port map ( Q=>d_arr_24_6, D=>nx68, CLK=>nx10133);
   ix69 : ao22 port map ( Y=>nx68, A0=>d_arr_mux_24_6, A1=>nx11247, B0=>
      d_arr_mul_24_6, B1=>nx10365);
   lat_d_arr_24_7 : latch port map ( Q=>d_arr_24_7, D=>nx76, CLK=>nx10135);
   ix77 : ao22 port map ( Y=>nx76, A0=>d_arr_mux_24_7, A1=>nx11247, B0=>
      d_arr_mul_24_7, B1=>nx10367);
   lat_d_arr_24_8 : latch port map ( Q=>d_arr_24_8, D=>nx84, CLK=>nx10135);
   ix85 : ao22 port map ( Y=>nx84, A0=>d_arr_mux_24_8, A1=>nx11247, B0=>
      d_arr_mul_24_8, B1=>nx10367);
   lat_d_arr_24_9 : latch port map ( Q=>d_arr_24_9, D=>nx92, CLK=>nx10135);
   ix93 : ao22 port map ( Y=>nx92, A0=>d_arr_mux_24_9, A1=>nx11247, B0=>
      d_arr_mul_24_9, B1=>nx10367);
   lat_d_arr_24_10 : latch port map ( Q=>d_arr_24_10, D=>nx100, CLK=>nx10135
   );
   ix101 : ao22 port map ( Y=>nx100, A0=>d_arr_mux_24_10, A1=>nx11247, B0=>
      d_arr_mul_24_10, B1=>nx10367);
   lat_d_arr_24_11 : latch port map ( Q=>d_arr_24_11, D=>nx108, CLK=>nx10135
   );
   ix109 : ao22 port map ( Y=>nx108, A0=>d_arr_mux_24_11, A1=>nx11247, B0=>
      d_arr_mul_24_11, B1=>nx10367);
   lat_d_arr_24_12 : latch port map ( Q=>d_arr_24_12, D=>nx116, CLK=>nx10135
   );
   ix117 : ao22 port map ( Y=>nx116, A0=>d_arr_mux_24_12, A1=>nx11247, B0=>
      d_arr_mul_24_12, B1=>nx10367);
   lat_d_arr_24_13 : latch port map ( Q=>d_arr_24_13, D=>nx124, CLK=>nx10135
   );
   ix125 : ao22 port map ( Y=>nx124, A0=>d_arr_mux_24_13, A1=>nx11249, B0=>
      d_arr_mul_24_13, B1=>nx10367);
   lat_d_arr_24_14 : latch port map ( Q=>d_arr_24_14, D=>nx132, CLK=>nx10137
   );
   ix133 : ao22 port map ( Y=>nx132, A0=>d_arr_mux_24_14, A1=>nx11249, B0=>
      d_arr_mul_24_14, B1=>nx10369);
   lat_d_arr_24_15 : latch port map ( Q=>d_arr_24_15, D=>nx140, CLK=>nx10137
   );
   lat_d_arr_24_16 : latch port map ( Q=>d_arr_24_16, D=>nx146, CLK=>nx10137
   );
   lat_d_arr_24_17 : latch port map ( Q=>d_arr_24_17, D=>nx152, CLK=>nx10137
   );
   lat_d_arr_24_18 : latch port map ( Q=>d_arr_24_18, D=>nx158, CLK=>nx10137
   );
   lat_d_arr_24_19 : latch port map ( Q=>d_arr_24_19, D=>nx164, CLK=>nx10137
   );
   lat_d_arr_24_20 : latch port map ( Q=>d_arr_24_20, D=>nx170, CLK=>nx10137
   );
   lat_d_arr_24_21 : latch port map ( Q=>d_arr_24_21, D=>nx176, CLK=>nx10139
   );
   lat_d_arr_24_22 : latch port map ( Q=>d_arr_24_22, D=>nx182, CLK=>nx10139
   );
   lat_d_arr_24_23 : latch port map ( Q=>d_arr_24_23, D=>nx188, CLK=>nx10139
   );
   lat_d_arr_24_24 : latch port map ( Q=>d_arr_24_24, D=>nx194, CLK=>nx10139
   );
   lat_d_arr_24_25 : latch port map ( Q=>d_arr_24_25, D=>nx200, CLK=>nx10139
   );
   lat_d_arr_24_26 : latch port map ( Q=>d_arr_24_26, D=>nx206, CLK=>nx10139
   );
   lat_d_arr_24_27 : latch port map ( Q=>d_arr_24_27, D=>nx212, CLK=>nx10139
   );
   lat_d_arr_24_28 : latch port map ( Q=>d_arr_24_28, D=>nx218, CLK=>nx10141
   );
   lat_d_arr_24_29 : latch port map ( Q=>d_arr_24_29, D=>nx224, CLK=>nx10141
   );
   lat_d_arr_24_30 : latch port map ( Q=>d_arr_24_30, D=>nx230, CLK=>nx10141
   );
   lat_d_arr_24_31 : latch port map ( Q=>d_arr_24_31, D=>nx236, CLK=>nx10141
   );
   lat_d_arr_23_0 : latch port map ( Q=>d_arr_23_0, D=>nx244, CLK=>nx10141);
   ix245 : ao22 port map ( Y=>nx244, A0=>d_arr_mux_23_0, A1=>nx11249, B0=>
      d_arr_mul_23_0, B1=>nx10373);
   lat_d_arr_23_1 : latch port map ( Q=>d_arr_23_1, D=>nx252, CLK=>nx10141);
   ix253 : ao22 port map ( Y=>nx252, A0=>d_arr_mux_23_1, A1=>nx11249, B0=>
      d_arr_mul_23_1, B1=>nx10373);
   lat_d_arr_23_2 : latch port map ( Q=>d_arr_23_2, D=>nx260, CLK=>nx10141);
   ix261 : ao22 port map ( Y=>nx260, A0=>d_arr_mux_23_2, A1=>nx11249, B0=>
      d_arr_mul_23_2, B1=>nx10373);
   lat_d_arr_23_3 : latch port map ( Q=>d_arr_23_3, D=>nx268, CLK=>nx10143);
   ix269 : ao22 port map ( Y=>nx268, A0=>d_arr_mux_23_3, A1=>nx11249, B0=>
      d_arr_mul_23_3, B1=>nx10375);
   lat_d_arr_23_4 : latch port map ( Q=>d_arr_23_4, D=>nx276, CLK=>nx10143);
   ix277 : ao22 port map ( Y=>nx276, A0=>d_arr_mux_23_4, A1=>nx11249, B0=>
      d_arr_mul_23_4, B1=>nx10375);
   lat_d_arr_23_5 : latch port map ( Q=>d_arr_23_5, D=>nx284, CLK=>nx10143);
   ix285 : ao22 port map ( Y=>nx284, A0=>d_arr_mux_23_5, A1=>nx11251, B0=>
      d_arr_mul_23_5, B1=>nx10375);
   lat_d_arr_23_6 : latch port map ( Q=>d_arr_23_6, D=>nx292, CLK=>nx10143);
   ix293 : ao22 port map ( Y=>nx292, A0=>d_arr_mux_23_6, A1=>nx11251, B0=>
      d_arr_mul_23_6, B1=>nx10375);
   lat_d_arr_23_7 : latch port map ( Q=>d_arr_23_7, D=>nx300, CLK=>nx10143);
   ix301 : ao22 port map ( Y=>nx300, A0=>d_arr_mux_23_7, A1=>nx11251, B0=>
      d_arr_mul_23_7, B1=>nx10375);
   lat_d_arr_23_8 : latch port map ( Q=>d_arr_23_8, D=>nx308, CLK=>nx10143);
   ix309 : ao22 port map ( Y=>nx308, A0=>d_arr_mux_23_8, A1=>nx11251, B0=>
      d_arr_mul_23_8, B1=>nx10375);
   lat_d_arr_23_9 : latch port map ( Q=>d_arr_23_9, D=>nx316, CLK=>nx10143);
   ix317 : ao22 port map ( Y=>nx316, A0=>d_arr_mux_23_9, A1=>nx11251, B0=>
      d_arr_mul_23_9, B1=>nx10375);
   lat_d_arr_23_10 : latch port map ( Q=>d_arr_23_10, D=>nx324, CLK=>nx10145
   );
   ix325 : ao22 port map ( Y=>nx324, A0=>d_arr_mux_23_10, A1=>nx11251, B0=>
      d_arr_mul_23_10, B1=>nx10377);
   lat_d_arr_23_11 : latch port map ( Q=>d_arr_23_11, D=>nx332, CLK=>nx10145
   );
   ix333 : ao22 port map ( Y=>nx332, A0=>d_arr_mux_23_11, A1=>nx11251, B0=>
      d_arr_mul_23_11, B1=>nx10377);
   lat_d_arr_23_12 : latch port map ( Q=>d_arr_23_12, D=>nx340, CLK=>nx10145
   );
   ix341 : ao22 port map ( Y=>nx340, A0=>d_arr_mux_23_12, A1=>nx11253, B0=>
      d_arr_mul_23_12, B1=>nx10377);
   lat_d_arr_23_13 : latch port map ( Q=>d_arr_23_13, D=>nx348, CLK=>nx10145
   );
   ix349 : ao22 port map ( Y=>nx348, A0=>d_arr_mux_23_13, A1=>nx11253, B0=>
      d_arr_mul_23_13, B1=>nx10377);
   lat_d_arr_23_14 : latch port map ( Q=>d_arr_23_14, D=>nx356, CLK=>nx10145
   );
   ix357 : ao22 port map ( Y=>nx356, A0=>d_arr_mux_23_14, A1=>nx11253, B0=>
      d_arr_mul_23_14, B1=>nx10377);
   lat_d_arr_23_15 : latch port map ( Q=>d_arr_23_15, D=>nx364, CLK=>nx10145
   );
   lat_d_arr_23_16 : latch port map ( Q=>d_arr_23_16, D=>nx370, CLK=>nx10145
   );
   lat_d_arr_23_17 : latch port map ( Q=>d_arr_23_17, D=>nx376, CLK=>nx10147
   );
   lat_d_arr_23_18 : latch port map ( Q=>d_arr_23_18, D=>nx382, CLK=>nx10147
   );
   lat_d_arr_23_19 : latch port map ( Q=>d_arr_23_19, D=>nx388, CLK=>nx10147
   );
   lat_d_arr_23_20 : latch port map ( Q=>d_arr_23_20, D=>nx394, CLK=>nx10147
   );
   lat_d_arr_23_21 : latch port map ( Q=>d_arr_23_21, D=>nx400, CLK=>nx10147
   );
   lat_d_arr_23_22 : latch port map ( Q=>d_arr_23_22, D=>nx406, CLK=>nx10147
   );
   lat_d_arr_23_23 : latch port map ( Q=>d_arr_23_23, D=>nx412, CLK=>nx10147
   );
   lat_d_arr_23_24 : latch port map ( Q=>d_arr_23_24, D=>nx418, CLK=>nx10149
   );
   lat_d_arr_23_25 : latch port map ( Q=>d_arr_23_25, D=>nx424, CLK=>nx10149
   );
   lat_d_arr_23_26 : latch port map ( Q=>d_arr_23_26, D=>nx430, CLK=>nx10149
   );
   lat_d_arr_23_27 : latch port map ( Q=>d_arr_23_27, D=>nx436, CLK=>nx10149
   );
   lat_d_arr_23_28 : latch port map ( Q=>d_arr_23_28, D=>nx442, CLK=>nx10149
   );
   lat_d_arr_23_29 : latch port map ( Q=>d_arr_23_29, D=>nx448, CLK=>nx10149
   );
   lat_d_arr_23_30 : latch port map ( Q=>d_arr_23_30, D=>nx454, CLK=>nx10149
   );
   lat_d_arr_23_31 : latch port map ( Q=>d_arr_23_31, D=>nx460, CLK=>nx10151
   );
   lat_d_arr_22_0 : latch port map ( Q=>d_arr_22_0, D=>nx468, CLK=>nx10151);
   ix469 : ao22 port map ( Y=>nx468, A0=>d_arr_mux_22_0, A1=>nx11253, B0=>
      d_arr_mul_22_0, B1=>nx10383);
   lat_d_arr_22_1 : latch port map ( Q=>d_arr_22_1, D=>nx476, CLK=>nx10151);
   ix477 : ao22 port map ( Y=>nx476, A0=>d_arr_mux_22_1, A1=>nx11253, B0=>
      d_arr_mul_22_1, B1=>nx10383);
   lat_d_arr_22_2 : latch port map ( Q=>d_arr_22_2, D=>nx484, CLK=>nx10151);
   ix485 : ao22 port map ( Y=>nx484, A0=>d_arr_mux_22_2, A1=>nx11253, B0=>
      d_arr_mul_22_2, B1=>nx10383);
   lat_d_arr_22_3 : latch port map ( Q=>d_arr_22_3, D=>nx492, CLK=>nx10151);
   ix493 : ao22 port map ( Y=>nx492, A0=>d_arr_mux_22_3, A1=>nx11253, B0=>
      d_arr_mul_22_3, B1=>nx10383);
   lat_d_arr_22_4 : latch port map ( Q=>d_arr_22_4, D=>nx500, CLK=>nx10151);
   ix501 : ao22 port map ( Y=>nx500, A0=>d_arr_mux_22_4, A1=>nx11255, B0=>
      d_arr_mul_22_4, B1=>nx10383);
   lat_d_arr_22_5 : latch port map ( Q=>d_arr_22_5, D=>nx508, CLK=>nx10151);
   ix509 : ao22 port map ( Y=>nx508, A0=>d_arr_mux_22_5, A1=>nx11255, B0=>
      d_arr_mul_22_5, B1=>nx10383);
   lat_d_arr_22_6 : latch port map ( Q=>d_arr_22_6, D=>nx516, CLK=>nx10153);
   ix517 : ao22 port map ( Y=>nx516, A0=>d_arr_mux_22_6, A1=>nx11255, B0=>
      d_arr_mul_22_6, B1=>nx10385);
   lat_d_arr_22_7 : latch port map ( Q=>d_arr_22_7, D=>nx524, CLK=>nx10153);
   ix525 : ao22 port map ( Y=>nx524, A0=>d_arr_mux_22_7, A1=>nx11255, B0=>
      d_arr_mul_22_7, B1=>nx10385);
   lat_d_arr_22_8 : latch port map ( Q=>d_arr_22_8, D=>nx532, CLK=>nx10153);
   ix533 : ao22 port map ( Y=>nx532, A0=>d_arr_mux_22_8, A1=>nx11255, B0=>
      d_arr_mul_22_8, B1=>nx10385);
   lat_d_arr_22_9 : latch port map ( Q=>d_arr_22_9, D=>nx540, CLK=>nx10153);
   ix541 : ao22 port map ( Y=>nx540, A0=>d_arr_mux_22_9, A1=>nx11255, B0=>
      d_arr_mul_22_9, B1=>nx10385);
   lat_d_arr_22_10 : latch port map ( Q=>d_arr_22_10, D=>nx548, CLK=>nx10153
   );
   ix549 : ao22 port map ( Y=>nx548, A0=>d_arr_mux_22_10, A1=>nx11255, B0=>
      d_arr_mul_22_10, B1=>nx10385);
   lat_d_arr_22_11 : latch port map ( Q=>d_arr_22_11, D=>nx556, CLK=>nx10153
   );
   ix557 : ao22 port map ( Y=>nx556, A0=>d_arr_mux_22_11, A1=>nx11257, B0=>
      d_arr_mul_22_11, B1=>nx10385);
   lat_d_arr_22_12 : latch port map ( Q=>d_arr_22_12, D=>nx564, CLK=>nx10153
   );
   ix565 : ao22 port map ( Y=>nx564, A0=>d_arr_mux_22_12, A1=>nx11257, B0=>
      d_arr_mul_22_12, B1=>nx10385);
   lat_d_arr_22_13 : latch port map ( Q=>d_arr_22_13, D=>nx572, CLK=>nx10155
   );
   ix573 : ao22 port map ( Y=>nx572, A0=>d_arr_mux_22_13, A1=>nx11257, B0=>
      d_arr_mul_22_13, B1=>nx10387);
   lat_d_arr_22_14 : latch port map ( Q=>d_arr_22_14, D=>nx580, CLK=>nx10155
   );
   ix581 : ao22 port map ( Y=>nx580, A0=>d_arr_mux_22_14, A1=>nx11257, B0=>
      d_arr_mul_22_14, B1=>nx10387);
   lat_d_arr_22_15 : latch port map ( Q=>d_arr_22_15, D=>nx588, CLK=>nx10155
   );
   lat_d_arr_22_16 : latch port map ( Q=>d_arr_22_16, D=>nx594, CLK=>nx10155
   );
   lat_d_arr_22_17 : latch port map ( Q=>d_arr_22_17, D=>nx600, CLK=>nx10155
   );
   lat_d_arr_22_18 : latch port map ( Q=>d_arr_22_18, D=>nx606, CLK=>nx10155
   );
   lat_d_arr_22_19 : latch port map ( Q=>d_arr_22_19, D=>nx612, CLK=>nx10155
   );
   lat_d_arr_22_20 : latch port map ( Q=>d_arr_22_20, D=>nx618, CLK=>nx10157
   );
   lat_d_arr_22_21 : latch port map ( Q=>d_arr_22_21, D=>nx624, CLK=>nx10157
   );
   lat_d_arr_22_22 : latch port map ( Q=>d_arr_22_22, D=>nx630, CLK=>nx10157
   );
   lat_d_arr_22_23 : latch port map ( Q=>d_arr_22_23, D=>nx636, CLK=>nx10157
   );
   lat_d_arr_22_24 : latch port map ( Q=>d_arr_22_24, D=>nx642, CLK=>nx10157
   );
   lat_d_arr_22_25 : latch port map ( Q=>d_arr_22_25, D=>nx648, CLK=>nx10157
   );
   lat_d_arr_22_26 : latch port map ( Q=>d_arr_22_26, D=>nx654, CLK=>nx10157
   );
   lat_d_arr_22_27 : latch port map ( Q=>d_arr_22_27, D=>nx660, CLK=>nx10159
   );
   lat_d_arr_22_28 : latch port map ( Q=>d_arr_22_28, D=>nx666, CLK=>nx10159
   );
   lat_d_arr_22_29 : latch port map ( Q=>d_arr_22_29, D=>nx672, CLK=>nx10159
   );
   lat_d_arr_22_30 : latch port map ( Q=>d_arr_22_30, D=>nx678, CLK=>nx10159
   );
   lat_d_arr_22_31 : latch port map ( Q=>d_arr_22_31, D=>nx684, CLK=>nx10159
   );
   lat_d_arr_21_0 : latch port map ( Q=>d_arr_21_0, D=>nx700, CLK=>nx10159);
   ix701 : inv01 port map ( Y=>nx700, A=>nx7201);
   ix7202 : aoi222 port map ( Y=>nx7201, A0=>d_arr_mux_21_0, A1=>nx11257, B0
      =>d_arr_mul_21_0, B1=>nx10391, C0=>d_arr_add_21_0, C1=>nx10621);
   ix695 : nor03_2x port map ( Y=>nx694, A0=>nx7205, A1=>nx11257, A2=>
      sel_mul);
   ix7206 : inv01 port map ( Y=>nx7205, A=>sel_add);
   lat_d_arr_21_1 : latch port map ( Q=>d_arr_21_1, D=>nx712, CLK=>nx10159);
   ix713 : inv01 port map ( Y=>nx712, A=>nx7209);
   ix7210 : aoi222 port map ( Y=>nx7209, A0=>d_arr_mux_21_1, A1=>nx11257, B0
      =>d_arr_mul_21_1, B1=>nx10391, C0=>d_arr_add_21_1, C1=>nx10621);
   lat_d_arr_21_2 : latch port map ( Q=>d_arr_21_2, D=>nx724, CLK=>nx10161);
   ix725 : inv01 port map ( Y=>nx724, A=>nx7215);
   ix7216 : aoi222 port map ( Y=>nx7215, A0=>d_arr_mux_21_2, A1=>nx11259, B0
      =>d_arr_mul_21_2, B1=>nx10393, C0=>d_arr_add_21_2, C1=>nx10621);
   lat_d_arr_21_3 : latch port map ( Q=>d_arr_21_3, D=>nx736, CLK=>nx10161);
   ix737 : inv01 port map ( Y=>nx736, A=>nx7221);
   ix7222 : aoi222 port map ( Y=>nx7221, A0=>d_arr_mux_21_3, A1=>nx11259, B0
      =>d_arr_mul_21_3, B1=>nx10393, C0=>d_arr_add_21_3, C1=>nx10621);
   lat_d_arr_21_4 : latch port map ( Q=>d_arr_21_4, D=>nx748, CLK=>nx10161);
   ix749 : inv01 port map ( Y=>nx748, A=>nx7227);
   ix7228 : aoi222 port map ( Y=>nx7227, A0=>d_arr_mux_21_4, A1=>nx11259, B0
      =>d_arr_mul_21_4, B1=>nx10393, C0=>d_arr_add_21_4, C1=>nx10621);
   lat_d_arr_21_5 : latch port map ( Q=>d_arr_21_5, D=>nx760, CLK=>nx10161);
   ix761 : inv01 port map ( Y=>nx760, A=>nx7233);
   ix7234 : aoi222 port map ( Y=>nx7233, A0=>d_arr_mux_21_5, A1=>nx11259, B0
      =>d_arr_mul_21_5, B1=>nx10393, C0=>d_arr_add_21_5, C1=>nx10621);
   lat_d_arr_21_6 : latch port map ( Q=>d_arr_21_6, D=>nx772, CLK=>nx10161);
   ix773 : inv01 port map ( Y=>nx772, A=>nx7239);
   ix7240 : aoi222 port map ( Y=>nx7239, A0=>d_arr_mux_21_6, A1=>nx11259, B0
      =>d_arr_mul_21_6, B1=>nx10393, C0=>d_arr_add_21_6, C1=>nx10621);
   lat_d_arr_21_7 : latch port map ( Q=>d_arr_21_7, D=>nx784, CLK=>nx10161);
   ix785 : inv01 port map ( Y=>nx784, A=>nx7245);
   ix7246 : aoi222 port map ( Y=>nx7245, A0=>d_arr_mux_21_7, A1=>nx11259, B0
      =>d_arr_mul_21_7, B1=>nx10393, C0=>d_arr_add_21_7, C1=>nx10623);
   lat_d_arr_21_8 : latch port map ( Q=>d_arr_21_8, D=>nx796, CLK=>nx10161);
   ix797 : inv01 port map ( Y=>nx796, A=>nx7251);
   ix7252 : aoi222 port map ( Y=>nx7251, A0=>d_arr_mux_21_8, A1=>nx11259, B0
      =>d_arr_mul_21_8, B1=>nx10393, C0=>d_arr_add_21_8, C1=>nx10623);
   lat_d_arr_21_9 : latch port map ( Q=>d_arr_21_9, D=>nx808, CLK=>nx10163);
   ix809 : inv01 port map ( Y=>nx808, A=>nx7257);
   ix7258 : aoi222 port map ( Y=>nx7257, A0=>d_arr_mux_21_9, A1=>nx11261, B0
      =>d_arr_mul_21_9, B1=>nx10395, C0=>d_arr_add_21_9, C1=>nx10623);
   lat_d_arr_21_10 : latch port map ( Q=>d_arr_21_10, D=>nx820, CLK=>nx10163
   );
   ix821 : inv01 port map ( Y=>nx820, A=>nx7263);
   ix7264 : aoi222 port map ( Y=>nx7263, A0=>d_arr_mux_21_10, A1=>nx11261, 
      B0=>d_arr_mul_21_10, B1=>nx10395, C0=>d_arr_add_21_10, C1=>nx10623);
   lat_d_arr_21_11 : latch port map ( Q=>d_arr_21_11, D=>nx832, CLK=>nx10163
   );
   ix833 : inv01 port map ( Y=>nx832, A=>nx7269);
   ix7270 : aoi222 port map ( Y=>nx7269, A0=>d_arr_mux_21_11, A1=>nx11261, 
      B0=>d_arr_mul_21_11, B1=>nx10395, C0=>d_arr_add_21_11, C1=>nx10623);
   lat_d_arr_21_12 : latch port map ( Q=>d_arr_21_12, D=>nx844, CLK=>nx10163
   );
   ix845 : inv01 port map ( Y=>nx844, A=>nx7275);
   ix7276 : aoi222 port map ( Y=>nx7275, A0=>d_arr_mux_21_12, A1=>nx11261, 
      B0=>d_arr_mul_21_12, B1=>nx10395, C0=>d_arr_add_21_12, C1=>nx10623);
   lat_d_arr_21_13 : latch port map ( Q=>d_arr_21_13, D=>nx856, CLK=>nx10163
   );
   ix857 : inv01 port map ( Y=>nx856, A=>nx7281);
   ix7282 : aoi222 port map ( Y=>nx7281, A0=>d_arr_mux_21_13, A1=>nx11261, 
      B0=>d_arr_mul_21_13, B1=>nx10395, C0=>d_arr_add_21_13, C1=>nx10623);
   lat_d_arr_21_14 : latch port map ( Q=>d_arr_21_14, D=>nx868, CLK=>nx10163
   );
   ix869 : inv01 port map ( Y=>nx868, A=>nx7287);
   ix7288 : aoi222 port map ( Y=>nx7287, A0=>d_arr_mux_21_14, A1=>nx11261, 
      B0=>d_arr_mul_21_14, B1=>nx10395, C0=>d_arr_add_21_14, C1=>nx10625);
   lat_d_arr_21_15 : latch port map ( Q=>d_arr_21_15, D=>nx880, CLK=>nx10163
   );
   ix881 : nand02 port map ( Y=>nx880, A0=>nx7293, A1=>nx10845);
   ix7294 : aoi22 port map ( Y=>nx7293, A0=>d_arr_mul_21_15, A1=>nx10395, B0
      =>d_arr_add_21_15, B1=>nx10625);
   ix7296 : nand02 port map ( Y=>nx7295, A0=>d_arr_mux_21_31, A1=>nx11261);
   lat_d_arr_21_16 : latch port map ( Q=>d_arr_21_16, D=>nx890, CLK=>nx10165
   );
   ix891 : nand02 port map ( Y=>nx890, A0=>nx7301, A1=>nx10845);
   ix7302 : aoi22 port map ( Y=>nx7301, A0=>d_arr_mul_21_16, A1=>nx10397, B0
      =>d_arr_add_21_16, B1=>nx10625);
   lat_d_arr_21_17 : latch port map ( Q=>d_arr_21_17, D=>nx900, CLK=>nx10165
   );
   ix901 : nand02 port map ( Y=>nx900, A0=>nx7305, A1=>nx10845);
   ix7306 : aoi22 port map ( Y=>nx7305, A0=>d_arr_mul_21_17, A1=>nx10397, B0
      =>d_arr_add_21_17, B1=>nx10625);
   lat_d_arr_21_18 : latch port map ( Q=>d_arr_21_18, D=>nx910, CLK=>nx10165
   );
   ix911 : nand02 port map ( Y=>nx910, A0=>nx7311, A1=>nx10845);
   ix7312 : aoi22 port map ( Y=>nx7311, A0=>d_arr_mul_21_18, A1=>nx10397, B0
      =>d_arr_add_21_18, B1=>nx10625);
   lat_d_arr_21_19 : latch port map ( Q=>d_arr_21_19, D=>nx920, CLK=>nx10165
   );
   ix921 : nand02 port map ( Y=>nx920, A0=>nx7317, A1=>nx10845);
   ix7318 : aoi22 port map ( Y=>nx7317, A0=>d_arr_mul_21_19, A1=>nx10397, B0
      =>d_arr_add_21_19, B1=>nx10625);
   lat_d_arr_21_20 : latch port map ( Q=>d_arr_21_20, D=>nx930, CLK=>nx10165
   );
   ix931 : nand02 port map ( Y=>nx930, A0=>nx7323, A1=>nx10845);
   ix7324 : aoi22 port map ( Y=>nx7323, A0=>d_arr_mul_21_20, A1=>nx10397, B0
      =>d_arr_add_21_20, B1=>nx10625);
   lat_d_arr_21_21 : latch port map ( Q=>d_arr_21_21, D=>nx940, CLK=>nx10165
   );
   ix941 : nand02 port map ( Y=>nx940, A0=>nx7329, A1=>nx10845);
   ix7330 : aoi22 port map ( Y=>nx7329, A0=>d_arr_mul_21_21, A1=>nx10397, B0
      =>d_arr_add_21_21, B1=>nx10627);
   lat_d_arr_21_22 : latch port map ( Q=>d_arr_21_22, D=>nx950, CLK=>nx10165
   );
   ix951 : nand02 port map ( Y=>nx950, A0=>nx7335, A1=>nx10847);
   ix7336 : aoi22 port map ( Y=>nx7335, A0=>d_arr_mul_21_22, A1=>nx10397, B0
      =>d_arr_add_21_22, B1=>nx10627);
   lat_d_arr_21_23 : latch port map ( Q=>d_arr_21_23, D=>nx960, CLK=>nx10167
   );
   ix961 : nand02 port map ( Y=>nx960, A0=>nx7341, A1=>nx10847);
   ix7342 : aoi22 port map ( Y=>nx7341, A0=>d_arr_mul_21_23, A1=>nx10399, B0
      =>d_arr_add_21_23, B1=>nx10627);
   lat_d_arr_21_24 : latch port map ( Q=>d_arr_21_24, D=>nx970, CLK=>nx10167
   );
   ix971 : nand02 port map ( Y=>nx970, A0=>nx7347, A1=>nx10847);
   ix7348 : aoi22 port map ( Y=>nx7347, A0=>d_arr_mul_21_24, A1=>nx10399, B0
      =>d_arr_add_21_24, B1=>nx10627);
   lat_d_arr_21_25 : latch port map ( Q=>d_arr_21_25, D=>nx980, CLK=>nx10167
   );
   ix981 : nand02 port map ( Y=>nx980, A0=>nx7353, A1=>nx10847);
   ix7354 : aoi22 port map ( Y=>nx7353, A0=>d_arr_mul_21_25, A1=>nx10399, B0
      =>d_arr_add_21_25, B1=>nx10627);
   lat_d_arr_21_26 : latch port map ( Q=>d_arr_21_26, D=>nx990, CLK=>nx10167
   );
   ix991 : nand02 port map ( Y=>nx990, A0=>nx7359, A1=>nx10847);
   ix7360 : aoi22 port map ( Y=>nx7359, A0=>d_arr_mul_21_26, A1=>nx10399, B0
      =>d_arr_add_21_26, B1=>nx10627);
   lat_d_arr_21_27 : latch port map ( Q=>d_arr_21_27, D=>nx1000, CLK=>
      nx10167);
   ix1001 : nand02 port map ( Y=>nx1000, A0=>nx7365, A1=>nx10847);
   ix7366 : aoi22 port map ( Y=>nx7365, A0=>d_arr_mul_21_27, A1=>nx10399, B0
      =>d_arr_add_21_27, B1=>nx10627);
   lat_d_arr_21_28 : latch port map ( Q=>d_arr_21_28, D=>nx1010, CLK=>
      nx10167);
   ix1011 : nand02 port map ( Y=>nx1010, A0=>nx7371, A1=>nx10847);
   ix7372 : aoi22 port map ( Y=>nx7371, A0=>d_arr_mul_21_28, A1=>nx10399, B0
      =>d_arr_add_21_28, B1=>nx10629);
   lat_d_arr_21_29 : latch port map ( Q=>d_arr_21_29, D=>nx1020, CLK=>
      nx10167);
   ix1021 : nand02 port map ( Y=>nx1020, A0=>nx7377, A1=>nx7295);
   ix7378 : aoi22 port map ( Y=>nx7377, A0=>d_arr_mul_21_29, A1=>nx10399, B0
      =>d_arr_add_21_29, B1=>nx10629);
   lat_d_arr_21_30 : latch port map ( Q=>d_arr_21_30, D=>nx1030, CLK=>
      nx10169);
   ix1031 : nand02 port map ( Y=>nx1030, A0=>nx7383, A1=>nx7295);
   ix7384 : aoi22 port map ( Y=>nx7383, A0=>d_arr_mul_21_30, A1=>nx10401, B0
      =>d_arr_add_21_30, B1=>nx10629);
   lat_d_arr_21_31 : latch port map ( Q=>d_arr_21_31, D=>nx1040, CLK=>
      nx10169);
   ix1041 : nand02 port map ( Y=>nx1040, A0=>nx7389, A1=>nx7295);
   ix7390 : aoi22 port map ( Y=>nx7389, A0=>d_arr_mul_21_31, A1=>nx10401, B0
      =>d_arr_add_21_31, B1=>nx10629);
   lat_d_arr_20_0 : latch port map ( Q=>d_arr_20_0, D=>nx1052, CLK=>nx10169
   );
   ix1053 : inv01 port map ( Y=>nx1052, A=>nx7395);
   ix7396 : aoi222 port map ( Y=>nx7395, A0=>d_arr_mux_20_0, A1=>nx11263, B0
      =>d_arr_mul_20_0, B1=>nx10401, C0=>d_arr_add_20_0, C1=>nx10629);
   lat_d_arr_20_1 : latch port map ( Q=>d_arr_20_1, D=>nx1064, CLK=>nx10169
   );
   ix1065 : inv01 port map ( Y=>nx1064, A=>nx7401);
   ix7402 : aoi222 port map ( Y=>nx7401, A0=>d_arr_mux_20_1, A1=>nx11263, B0
      =>d_arr_mul_20_1, B1=>nx10401, C0=>d_arr_add_20_1, C1=>nx10629);
   lat_d_arr_20_2 : latch port map ( Q=>d_arr_20_2, D=>nx1076, CLK=>nx10169
   );
   ix1077 : inv01 port map ( Y=>nx1076, A=>nx7407);
   ix7408 : aoi222 port map ( Y=>nx7407, A0=>d_arr_mux_20_2, A1=>nx11263, B0
      =>d_arr_mul_20_2, B1=>nx10401, C0=>d_arr_add_20_2, C1=>nx10629);
   lat_d_arr_20_3 : latch port map ( Q=>d_arr_20_3, D=>nx1088, CLK=>nx10169
   );
   ix1089 : inv01 port map ( Y=>nx1088, A=>nx7413);
   ix7414 : aoi222 port map ( Y=>nx7413, A0=>d_arr_mux_20_3, A1=>nx11263, B0
      =>d_arr_mul_20_3, B1=>nx10401, C0=>d_arr_add_20_3, C1=>nx10631);
   lat_d_arr_20_4 : latch port map ( Q=>d_arr_20_4, D=>nx1100, CLK=>nx10169
   );
   ix1101 : inv01 port map ( Y=>nx1100, A=>nx7419);
   ix7420 : aoi222 port map ( Y=>nx7419, A0=>d_arr_mux_20_4, A1=>nx11263, B0
      =>d_arr_mul_20_4, B1=>nx10401, C0=>d_arr_add_20_4, C1=>nx10631);
   lat_d_arr_20_5 : latch port map ( Q=>d_arr_20_5, D=>nx1112, CLK=>nx10171
   );
   ix1113 : inv01 port map ( Y=>nx1112, A=>nx7425);
   ix7426 : aoi222 port map ( Y=>nx7425, A0=>d_arr_mux_20_5, A1=>nx11263, B0
      =>d_arr_mul_20_5, B1=>nx10403, C0=>d_arr_add_20_5, C1=>nx10631);
   lat_d_arr_20_6 : latch port map ( Q=>d_arr_20_6, D=>nx1124, CLK=>nx10171
   );
   ix1125 : inv01 port map ( Y=>nx1124, A=>nx7431);
   ix7432 : aoi222 port map ( Y=>nx7431, A0=>d_arr_mux_20_6, A1=>nx11263, B0
      =>d_arr_mul_20_6, B1=>nx10403, C0=>d_arr_add_20_6, C1=>nx10631);
   lat_d_arr_20_7 : latch port map ( Q=>d_arr_20_7, D=>nx1136, CLK=>nx10171
   );
   ix1137 : inv01 port map ( Y=>nx1136, A=>nx7437);
   ix7438 : aoi222 port map ( Y=>nx7437, A0=>d_arr_mux_20_7, A1=>nx11265, B0
      =>d_arr_mul_20_7, B1=>nx10403, C0=>d_arr_add_20_7, C1=>nx10631);
   lat_d_arr_20_8 : latch port map ( Q=>d_arr_20_8, D=>nx1148, CLK=>nx10171
   );
   ix1149 : inv01 port map ( Y=>nx1148, A=>nx7441);
   ix7442 : aoi222 port map ( Y=>nx7441, A0=>d_arr_mux_20_8, A1=>nx11265, B0
      =>d_arr_mul_20_8, B1=>nx10403, C0=>d_arr_add_20_8, C1=>nx10631);
   lat_d_arr_20_9 : latch port map ( Q=>d_arr_20_9, D=>nx1160, CLK=>nx10171
   );
   ix1161 : inv01 port map ( Y=>nx1160, A=>nx7447);
   ix7448 : aoi222 port map ( Y=>nx7447, A0=>d_arr_mux_20_9, A1=>nx11265, B0
      =>d_arr_mul_20_9, B1=>nx10403, C0=>d_arr_add_20_9, C1=>nx10631);
   lat_d_arr_20_10 : latch port map ( Q=>d_arr_20_10, D=>nx1172, CLK=>
      nx10171);
   ix1173 : inv01 port map ( Y=>nx1172, A=>nx7453);
   ix7454 : aoi222 port map ( Y=>nx7453, A0=>d_arr_mux_20_10, A1=>nx11265, 
      B0=>d_arr_mul_20_10, B1=>nx10403, C0=>d_arr_add_20_10, C1=>nx10633);
   lat_d_arr_20_11 : latch port map ( Q=>d_arr_20_11, D=>nx1184, CLK=>
      nx10171);
   ix1185 : inv01 port map ( Y=>nx1184, A=>nx7459);
   ix7460 : aoi222 port map ( Y=>nx7459, A0=>d_arr_mux_20_11, A1=>nx11265, 
      B0=>d_arr_mul_20_11, B1=>nx10403, C0=>d_arr_add_20_11, C1=>nx10633);
   lat_d_arr_20_12 : latch port map ( Q=>d_arr_20_12, D=>nx1196, CLK=>
      nx10173);
   ix1197 : inv01 port map ( Y=>nx1196, A=>nx7463);
   ix7464 : aoi222 port map ( Y=>nx7463, A0=>d_arr_mux_20_12, A1=>nx11265, 
      B0=>d_arr_mul_20_12, B1=>nx10405, C0=>d_arr_add_20_12, C1=>nx10633);
   lat_d_arr_20_13 : latch port map ( Q=>d_arr_20_13, D=>nx1208, CLK=>
      nx10173);
   ix1209 : inv01 port map ( Y=>nx1208, A=>nx7469);
   ix7470 : aoi222 port map ( Y=>nx7469, A0=>d_arr_mux_20_13, A1=>nx11265, 
      B0=>d_arr_mul_20_13, B1=>nx10405, C0=>d_arr_add_20_13, C1=>nx10633);
   lat_d_arr_20_14 : latch port map ( Q=>d_arr_20_14, D=>nx1220, CLK=>
      nx10173);
   ix1221 : inv01 port map ( Y=>nx1220, A=>nx7475);
   ix7476 : aoi222 port map ( Y=>nx7475, A0=>d_arr_mux_20_14, A1=>nx11267, 
      B0=>d_arr_mul_20_14, B1=>nx10405, C0=>d_arr_add_20_14, C1=>nx10633);
   lat_d_arr_20_15 : latch port map ( Q=>d_arr_20_15, D=>nx1232, CLK=>
      nx10173);
   ix1233 : nand02 port map ( Y=>nx1232, A0=>nx7481, A1=>nx10849);
   ix7482 : aoi22 port map ( Y=>nx7481, A0=>d_arr_mul_20_15, A1=>nx10405, B0
      =>d_arr_add_20_15, B1=>nx10633);
   ix7484 : nand02 port map ( Y=>nx7483, A0=>d_arr_mux_20_31, A1=>nx11267);
   lat_d_arr_20_16 : latch port map ( Q=>d_arr_20_16, D=>nx1242, CLK=>
      nx10173);
   ix1243 : nand02 port map ( Y=>nx1242, A0=>nx7489, A1=>nx10849);
   ix7490 : aoi22 port map ( Y=>nx7489, A0=>d_arr_mul_20_16, A1=>nx10405, B0
      =>d_arr_add_20_16, B1=>nx10633);
   lat_d_arr_20_17 : latch port map ( Q=>d_arr_20_17, D=>nx1252, CLK=>
      nx10173);
   ix1253 : nand02 port map ( Y=>nx1252, A0=>nx7495, A1=>nx10849);
   ix7496 : aoi22 port map ( Y=>nx7495, A0=>d_arr_mul_20_17, A1=>nx10405, B0
      =>d_arr_add_20_17, B1=>nx10635);
   lat_d_arr_20_18 : latch port map ( Q=>d_arr_20_18, D=>nx1262, CLK=>
      nx10173);
   ix1263 : nand02 port map ( Y=>nx1262, A0=>nx7501, A1=>nx10849);
   ix7502 : aoi22 port map ( Y=>nx7501, A0=>d_arr_mul_20_18, A1=>nx10405, B0
      =>d_arr_add_20_18, B1=>nx10635);
   lat_d_arr_20_19 : latch port map ( Q=>d_arr_20_19, D=>nx1272, CLK=>
      nx10175);
   ix1273 : nand02 port map ( Y=>nx1272, A0=>nx7507, A1=>nx10849);
   ix7508 : aoi22 port map ( Y=>nx7507, A0=>d_arr_mul_20_19, A1=>nx10407, B0
      =>d_arr_add_20_19, B1=>nx10635);
   lat_d_arr_20_20 : latch port map ( Q=>d_arr_20_20, D=>nx1282, CLK=>
      nx10175);
   ix1283 : nand02 port map ( Y=>nx1282, A0=>nx7513, A1=>nx10849);
   ix7514 : aoi22 port map ( Y=>nx7513, A0=>d_arr_mul_20_20, A1=>nx10407, B0
      =>d_arr_add_20_20, B1=>nx10635);
   lat_d_arr_20_21 : latch port map ( Q=>d_arr_20_21, D=>nx1292, CLK=>
      nx10175);
   ix1293 : nand02 port map ( Y=>nx1292, A0=>nx7519, A1=>nx10849);
   ix7520 : aoi22 port map ( Y=>nx7519, A0=>d_arr_mul_20_21, A1=>nx10407, B0
      =>d_arr_add_20_21, B1=>nx10635);
   lat_d_arr_20_22 : latch port map ( Q=>d_arr_20_22, D=>nx1302, CLK=>
      nx10175);
   ix1303 : nand02 port map ( Y=>nx1302, A0=>nx7525, A1=>nx10851);
   ix7526 : aoi22 port map ( Y=>nx7525, A0=>d_arr_mul_20_22, A1=>nx10407, B0
      =>d_arr_add_20_22, B1=>nx10635);
   lat_d_arr_20_23 : latch port map ( Q=>d_arr_20_23, D=>nx1312, CLK=>
      nx10175);
   ix1313 : nand02 port map ( Y=>nx1312, A0=>nx7529, A1=>nx10851);
   ix7530 : aoi22 port map ( Y=>nx7529, A0=>d_arr_mul_20_23, A1=>nx10407, B0
      =>d_arr_add_20_23, B1=>nx10635);
   lat_d_arr_20_24 : latch port map ( Q=>d_arr_20_24, D=>nx1322, CLK=>
      nx10175);
   ix1323 : nand02 port map ( Y=>nx1322, A0=>nx7535, A1=>nx10851);
   ix7536 : aoi22 port map ( Y=>nx7535, A0=>d_arr_mul_20_24, A1=>nx10407, B0
      =>d_arr_add_20_24, B1=>nx10637);
   lat_d_arr_20_25 : latch port map ( Q=>d_arr_20_25, D=>nx1332, CLK=>
      nx10175);
   ix1333 : nand02 port map ( Y=>nx1332, A0=>nx7541, A1=>nx10851);
   ix7542 : aoi22 port map ( Y=>nx7541, A0=>d_arr_mul_20_25, A1=>nx10407, B0
      =>d_arr_add_20_25, B1=>nx10637);
   lat_d_arr_20_26 : latch port map ( Q=>d_arr_20_26, D=>nx1342, CLK=>
      nx10177);
   ix1343 : nand02 port map ( Y=>nx1342, A0=>nx7547, A1=>nx10851);
   ix7548 : aoi22 port map ( Y=>nx7547, A0=>d_arr_mul_20_26, A1=>nx10409, B0
      =>d_arr_add_20_26, B1=>nx10637);
   lat_d_arr_20_27 : latch port map ( Q=>d_arr_20_27, D=>nx1352, CLK=>
      nx10177);
   ix1353 : nand02 port map ( Y=>nx1352, A0=>nx7551, A1=>nx10851);
   ix7552 : aoi22 port map ( Y=>nx7551, A0=>d_arr_mul_20_27, A1=>nx10409, B0
      =>d_arr_add_20_27, B1=>nx10637);
   lat_d_arr_20_28 : latch port map ( Q=>d_arr_20_28, D=>nx1362, CLK=>
      nx10177);
   ix1363 : nand02 port map ( Y=>nx1362, A0=>nx7557, A1=>nx10851);
   ix7558 : aoi22 port map ( Y=>nx7557, A0=>d_arr_mul_20_28, A1=>nx10409, B0
      =>d_arr_add_20_28, B1=>nx10637);
   lat_d_arr_20_29 : latch port map ( Q=>d_arr_20_29, D=>nx1372, CLK=>
      nx10177);
   ix1373 : nand02 port map ( Y=>nx1372, A0=>nx7563, A1=>nx7483);
   ix7564 : aoi22 port map ( Y=>nx7563, A0=>d_arr_mul_20_29, A1=>nx10409, B0
      =>d_arr_add_20_29, B1=>nx10637);
   lat_d_arr_20_30 : latch port map ( Q=>d_arr_20_30, D=>nx1382, CLK=>
      nx10177);
   ix1383 : nand02 port map ( Y=>nx1382, A0=>nx7569, A1=>nx7483);
   ix7570 : aoi22 port map ( Y=>nx7569, A0=>d_arr_mul_20_30, A1=>nx10409, B0
      =>d_arr_add_20_30, B1=>nx10637);
   lat_d_arr_20_31 : latch port map ( Q=>d_arr_20_31, D=>nx1392, CLK=>
      nx10177);
   ix1393 : nand02 port map ( Y=>nx1392, A0=>nx7573, A1=>nx7483);
   ix7574 : aoi22 port map ( Y=>nx7573, A0=>d_arr_mul_20_31, A1=>nx10409, B0
      =>d_arr_add_20_31, B1=>nx10639);
   lat_d_arr_19_0 : latch port map ( Q=>d_arr_19_0, D=>nx1404, CLK=>nx10177
   );
   ix1405 : inv01 port map ( Y=>nx1404, A=>nx7579);
   ix7580 : aoi222 port map ( Y=>nx7579, A0=>d_arr_mux_19_0, A1=>nx11267, B0
      =>d_arr_mul_19_0, B1=>nx10409, C0=>d_arr_add_19_0, C1=>nx10639);
   lat_d_arr_19_1 : latch port map ( Q=>d_arr_19_1, D=>nx1416, CLK=>nx10179
   );
   ix1417 : inv01 port map ( Y=>nx1416, A=>nx7585);
   ix7586 : aoi222 port map ( Y=>nx7585, A0=>d_arr_mux_19_1, A1=>nx11267, B0
      =>d_arr_mul_19_1, B1=>nx10411, C0=>d_arr_add_19_1, C1=>nx10639);
   lat_d_arr_19_2 : latch port map ( Q=>d_arr_19_2, D=>nx1428, CLK=>nx10179
   );
   ix1429 : inv01 port map ( Y=>nx1428, A=>nx7591);
   ix7592 : aoi222 port map ( Y=>nx7591, A0=>d_arr_mux_19_2, A1=>nx11267, B0
      =>d_arr_mul_19_2, B1=>nx10411, C0=>d_arr_add_19_2, C1=>nx10639);
   lat_d_arr_19_3 : latch port map ( Q=>d_arr_19_3, D=>nx1440, CLK=>nx10179
   );
   ix1441 : inv01 port map ( Y=>nx1440, A=>nx7595);
   ix7596 : aoi222 port map ( Y=>nx7595, A0=>d_arr_mux_19_3, A1=>nx11267, B0
      =>d_arr_mul_19_3, B1=>nx10411, C0=>d_arr_add_19_3, C1=>nx10639);
   lat_d_arr_19_4 : latch port map ( Q=>d_arr_19_4, D=>nx1452, CLK=>nx10179
   );
   ix1453 : inv01 port map ( Y=>nx1452, A=>nx7601);
   ix7602 : aoi222 port map ( Y=>nx7601, A0=>d_arr_mux_19_4, A1=>nx11267, B0
      =>d_arr_mul_19_4, B1=>nx10411, C0=>d_arr_add_19_4, C1=>nx10639);
   lat_d_arr_19_5 : latch port map ( Q=>d_arr_19_5, D=>nx1464, CLK=>nx10179
   );
   ix1465 : inv01 port map ( Y=>nx1464, A=>nx7607);
   ix7608 : aoi222 port map ( Y=>nx7607, A0=>d_arr_mux_19_5, A1=>nx11269, B0
      =>d_arr_mul_19_5, B1=>nx10411, C0=>d_arr_add_19_5, C1=>nx10639);
   lat_d_arr_19_6 : latch port map ( Q=>d_arr_19_6, D=>nx1476, CLK=>nx10179
   );
   ix1477 : inv01 port map ( Y=>nx1476, A=>nx7613);
   ix7614 : aoi222 port map ( Y=>nx7613, A0=>d_arr_mux_19_6, A1=>nx11269, B0
      =>d_arr_mul_19_6, B1=>nx10411, C0=>d_arr_add_19_6, C1=>nx10641);
   lat_d_arr_19_7 : latch port map ( Q=>d_arr_19_7, D=>nx1488, CLK=>nx10179
   );
   ix1489 : inv01 port map ( Y=>nx1488, A=>nx7617);
   ix7618 : aoi222 port map ( Y=>nx7617, A0=>d_arr_mux_19_7, A1=>nx11269, B0
      =>d_arr_mul_19_7, B1=>nx10411, C0=>d_arr_add_19_7, C1=>nx10641);
   lat_d_arr_19_8 : latch port map ( Q=>d_arr_19_8, D=>nx1500, CLK=>nx10181
   );
   ix1501 : inv01 port map ( Y=>nx1500, A=>nx7623);
   ix7624 : aoi222 port map ( Y=>nx7623, A0=>d_arr_mux_19_8, A1=>nx11269, B0
      =>d_arr_mul_19_8, B1=>nx10413, C0=>d_arr_add_19_8, C1=>nx10641);
   lat_d_arr_19_9 : latch port map ( Q=>d_arr_19_9, D=>nx1512, CLK=>nx10181
   );
   ix1513 : inv01 port map ( Y=>nx1512, A=>nx7629);
   ix7630 : aoi222 port map ( Y=>nx7629, A0=>d_arr_mux_19_9, A1=>nx11269, B0
      =>d_arr_mul_19_9, B1=>nx10413, C0=>d_arr_add_19_9, C1=>nx10641);
   lat_d_arr_19_10 : latch port map ( Q=>d_arr_19_10, D=>nx1524, CLK=>
      nx10181);
   ix1525 : inv01 port map ( Y=>nx1524, A=>nx7635);
   ix7636 : aoi222 port map ( Y=>nx7635, A0=>d_arr_mux_19_10, A1=>nx11269, 
      B0=>d_arr_mul_19_10, B1=>nx10413, C0=>d_arr_add_19_10, C1=>nx10641);
   lat_d_arr_19_11 : latch port map ( Q=>d_arr_19_11, D=>nx1536, CLK=>
      nx10181);
   ix1537 : inv01 port map ( Y=>nx1536, A=>nx7639);
   ix7640 : aoi222 port map ( Y=>nx7639, A0=>d_arr_mux_19_11, A1=>nx11269, 
      B0=>d_arr_mul_19_11, B1=>nx10413, C0=>d_arr_add_19_11, C1=>nx10641);
   lat_d_arr_19_12 : latch port map ( Q=>d_arr_19_12, D=>nx1548, CLK=>
      nx10181);
   ix1549 : inv01 port map ( Y=>nx1548, A=>nx7645);
   ix7646 : aoi222 port map ( Y=>nx7645, A0=>d_arr_mux_19_12, A1=>nx11271, 
      B0=>d_arr_mul_19_12, B1=>nx10413, C0=>d_arr_add_19_12, C1=>nx10641);
   lat_d_arr_19_13 : latch port map ( Q=>d_arr_19_13, D=>nx1560, CLK=>
      nx10181);
   ix1561 : inv01 port map ( Y=>nx1560, A=>nx7651);
   ix7652 : aoi222 port map ( Y=>nx7651, A0=>d_arr_mux_19_13, A1=>nx11271, 
      B0=>d_arr_mul_19_13, B1=>nx10413, C0=>d_arr_add_19_13, C1=>nx10643);
   lat_d_arr_19_14 : latch port map ( Q=>d_arr_19_14, D=>nx1572, CLK=>
      nx10181);
   ix1573 : inv01 port map ( Y=>nx1572, A=>nx7657);
   ix7658 : aoi222 port map ( Y=>nx7657, A0=>d_arr_mux_19_14, A1=>nx11271, 
      B0=>d_arr_mul_19_14, B1=>nx10413, C0=>d_arr_add_19_14, C1=>nx10643);
   lat_d_arr_19_15 : latch port map ( Q=>d_arr_19_15, D=>nx1584, CLK=>
      nx10183);
   ix1585 : nand02 port map ( Y=>nx1584, A0=>nx7661, A1=>nx10853);
   ix7662 : aoi22 port map ( Y=>nx7661, A0=>d_arr_mul_19_15, A1=>nx10415, B0
      =>d_arr_add_19_15, B1=>nx10643);
   ix7664 : nand02 port map ( Y=>nx7663, A0=>d_arr_mux_19_31, A1=>nx11271);
   lat_d_arr_19_16 : latch port map ( Q=>d_arr_19_16, D=>nx1594, CLK=>
      nx10183);
   ix1595 : nand02 port map ( Y=>nx1594, A0=>nx7669, A1=>nx10853);
   ix7670 : aoi22 port map ( Y=>nx7669, A0=>d_arr_mul_19_16, A1=>nx10415, B0
      =>d_arr_add_19_16, B1=>nx10643);
   lat_d_arr_19_17 : latch port map ( Q=>d_arr_19_17, D=>nx1604, CLK=>
      nx10183);
   ix1605 : nand02 port map ( Y=>nx1604, A0=>nx7675, A1=>nx10853);
   ix7676 : aoi22 port map ( Y=>nx7675, A0=>d_arr_mul_19_17, A1=>nx10415, B0
      =>d_arr_add_19_17, B1=>nx10643);
   lat_d_arr_19_18 : latch port map ( Q=>d_arr_19_18, D=>nx1614, CLK=>
      nx10183);
   ix1615 : nand02 port map ( Y=>nx1614, A0=>nx7681, A1=>nx10853);
   ix7682 : aoi22 port map ( Y=>nx7681, A0=>d_arr_mul_19_18, A1=>nx10415, B0
      =>d_arr_add_19_18, B1=>nx10643);
   lat_d_arr_19_19 : latch port map ( Q=>d_arr_19_19, D=>nx1624, CLK=>
      nx10183);
   ix1625 : nand02 port map ( Y=>nx1624, A0=>nx7687, A1=>nx10853);
   ix7688 : aoi22 port map ( Y=>nx7687, A0=>d_arr_mul_19_19, A1=>nx10415, B0
      =>d_arr_add_19_19, B1=>nx10643);
   lat_d_arr_19_20 : latch port map ( Q=>d_arr_19_20, D=>nx1634, CLK=>
      nx10183);
   ix1635 : nand02 port map ( Y=>nx1634, A0=>nx7693, A1=>nx10853);
   ix7694 : aoi22 port map ( Y=>nx7693, A0=>d_arr_mul_19_20, A1=>nx10415, B0
      =>d_arr_add_19_20, B1=>nx10645);
   lat_d_arr_19_21 : latch port map ( Q=>d_arr_19_21, D=>nx1644, CLK=>
      nx10183);
   ix1645 : nand02 port map ( Y=>nx1644, A0=>nx7699, A1=>nx10853);
   ix7700 : aoi22 port map ( Y=>nx7699, A0=>d_arr_mul_19_21, A1=>nx10415, B0
      =>d_arr_add_19_21, B1=>nx10645);
   lat_d_arr_19_22 : latch port map ( Q=>d_arr_19_22, D=>nx1654, CLK=>
      nx10185);
   ix1655 : nand02 port map ( Y=>nx1654, A0=>nx7705, A1=>nx10855);
   ix7706 : aoi22 port map ( Y=>nx7705, A0=>d_arr_mul_19_22, A1=>nx10417, B0
      =>d_arr_add_19_22, B1=>nx10645);
   lat_d_arr_19_23 : latch port map ( Q=>d_arr_19_23, D=>nx1664, CLK=>
      nx10185);
   ix1665 : nand02 port map ( Y=>nx1664, A0=>nx7711, A1=>nx10855);
   ix7712 : aoi22 port map ( Y=>nx7711, A0=>d_arr_mul_19_23, A1=>nx10417, B0
      =>d_arr_add_19_23, B1=>nx10645);
   lat_d_arr_19_24 : latch port map ( Q=>d_arr_19_24, D=>nx1674, CLK=>
      nx10185);
   ix1675 : nand02 port map ( Y=>nx1674, A0=>nx7717, A1=>nx10855);
   ix7718 : aoi22 port map ( Y=>nx7717, A0=>d_arr_mul_19_24, A1=>nx10417, B0
      =>d_arr_add_19_24, B1=>nx10645);
   lat_d_arr_19_25 : latch port map ( Q=>d_arr_19_25, D=>nx1684, CLK=>
      nx10185);
   ix1685 : nand02 port map ( Y=>nx1684, A0=>nx7723, A1=>nx10855);
   ix7724 : aoi22 port map ( Y=>nx7723, A0=>d_arr_mul_19_25, A1=>nx10417, B0
      =>d_arr_add_19_25, B1=>nx10645);
   lat_d_arr_19_26 : latch port map ( Q=>d_arr_19_26, D=>nx1694, CLK=>
      nx10185);
   ix1695 : nand02 port map ( Y=>nx1694, A0=>nx7727, A1=>nx10855);
   ix7728 : aoi22 port map ( Y=>nx7727, A0=>d_arr_mul_19_26, A1=>nx10417, B0
      =>d_arr_add_19_26, B1=>nx10645);
   lat_d_arr_19_27 : latch port map ( Q=>d_arr_19_27, D=>nx1704, CLK=>
      nx10185);
   ix1705 : nand02 port map ( Y=>nx1704, A0=>nx7733, A1=>nx10855);
   ix7734 : aoi22 port map ( Y=>nx7733, A0=>d_arr_mul_19_27, A1=>nx10417, B0
      =>d_arr_add_19_27, B1=>nx10647);
   lat_d_arr_19_28 : latch port map ( Q=>d_arr_19_28, D=>nx1714, CLK=>
      nx10185);
   ix1715 : nand02 port map ( Y=>nx1714, A0=>nx7739, A1=>nx10855);
   ix7740 : aoi22 port map ( Y=>nx7739, A0=>d_arr_mul_19_28, A1=>nx10417, B0
      =>d_arr_add_19_28, B1=>nx10647);
   lat_d_arr_19_29 : latch port map ( Q=>d_arr_19_29, D=>nx1724, CLK=>
      nx10187);
   ix1725 : nand02 port map ( Y=>nx1724, A0=>nx7745, A1=>nx7663);
   ix7746 : aoi22 port map ( Y=>nx7745, A0=>d_arr_mul_19_29, A1=>nx10419, B0
      =>d_arr_add_19_29, B1=>nx10647);
   lat_d_arr_19_30 : latch port map ( Q=>d_arr_19_30, D=>nx1734, CLK=>
      nx10187);
   ix1735 : nand02 port map ( Y=>nx1734, A0=>nx7749, A1=>nx7663);
   ix7750 : aoi22 port map ( Y=>nx7749, A0=>d_arr_mul_19_30, A1=>nx10419, B0
      =>d_arr_add_19_30, B1=>nx10647);
   lat_d_arr_19_31 : latch port map ( Q=>d_arr_19_31, D=>nx1744, CLK=>
      nx10187);
   ix1745 : nand02 port map ( Y=>nx1744, A0=>nx7755, A1=>nx7663);
   ix7756 : aoi22 port map ( Y=>nx7755, A0=>d_arr_mul_19_31, A1=>nx10419, B0
      =>d_arr_add_19_31, B1=>nx10647);
   lat_d_arr_18_0 : latch port map ( Q=>d_arr_18_0, D=>nx1756, CLK=>nx10187
   );
   ix1757 : inv01 port map ( Y=>nx1756, A=>nx7761);
   ix7762 : aoi222 port map ( Y=>nx7761, A0=>d_arr_mux_18_0, A1=>nx11271, B0
      =>d_arr_mul_18_0, B1=>nx10419, C0=>d_arr_add_18_0, C1=>nx10647);
   lat_d_arr_18_1 : latch port map ( Q=>d_arr_18_1, D=>nx1768, CLK=>nx10187
   );
   ix1769 : inv01 port map ( Y=>nx1768, A=>nx7767);
   ix7768 : aoi222 port map ( Y=>nx7767, A0=>d_arr_mux_18_1, A1=>nx11271, B0
      =>d_arr_mul_18_1, B1=>nx10419, C0=>d_arr_add_18_1, C1=>nx10647);
   lat_d_arr_18_2 : latch port map ( Q=>d_arr_18_2, D=>nx1780, CLK=>nx10187
   );
   ix1781 : inv01 port map ( Y=>nx1780, A=>nx7773);
   ix7774 : aoi222 port map ( Y=>nx7773, A0=>d_arr_mux_18_2, A1=>nx11271, B0
      =>d_arr_mul_18_2, B1=>nx10419, C0=>d_arr_add_18_2, C1=>nx10649);
   lat_d_arr_18_3 : latch port map ( Q=>d_arr_18_3, D=>nx1792, CLK=>nx10187
   );
   ix1793 : inv01 port map ( Y=>nx1792, A=>nx7779);
   ix7780 : aoi222 port map ( Y=>nx7779, A0=>d_arr_mux_18_3, A1=>nx11273, B0
      =>d_arr_mul_18_3, B1=>nx10419, C0=>d_arr_add_18_3, C1=>nx10649);
   lat_d_arr_18_4 : latch port map ( Q=>d_arr_18_4, D=>nx1804, CLK=>nx10189
   );
   ix1805 : inv01 port map ( Y=>nx1804, A=>nx7785);
   ix7786 : aoi222 port map ( Y=>nx7785, A0=>d_arr_mux_18_4, A1=>nx11273, B0
      =>d_arr_mul_18_4, B1=>nx10421, C0=>d_arr_add_18_4, C1=>nx10649);
   lat_d_arr_18_5 : latch port map ( Q=>d_arr_18_5, D=>nx1816, CLK=>nx10189
   );
   ix1817 : inv01 port map ( Y=>nx1816, A=>nx7791);
   ix7792 : aoi222 port map ( Y=>nx7791, A0=>d_arr_mux_18_5, A1=>nx11273, B0
      =>d_arr_mul_18_5, B1=>nx10421, C0=>d_arr_add_18_5, C1=>nx10649);
   lat_d_arr_18_6 : latch port map ( Q=>d_arr_18_6, D=>nx1828, CLK=>nx10189
   );
   ix1829 : inv01 port map ( Y=>nx1828, A=>nx7797);
   ix7798 : aoi222 port map ( Y=>nx7797, A0=>d_arr_mux_18_6, A1=>nx11273, B0
      =>d_arr_mul_18_6, B1=>nx10421, C0=>d_arr_add_18_6, C1=>nx10649);
   lat_d_arr_18_7 : latch port map ( Q=>d_arr_18_7, D=>nx1840, CLK=>nx10189
   );
   ix1841 : inv01 port map ( Y=>nx1840, A=>nx7803);
   ix7804 : aoi222 port map ( Y=>nx7803, A0=>d_arr_mux_18_7, A1=>nx11273, B0
      =>d_arr_mul_18_7, B1=>nx10421, C0=>d_arr_add_18_7, C1=>nx10649);
   lat_d_arr_18_8 : latch port map ( Q=>d_arr_18_8, D=>nx1852, CLK=>nx10189
   );
   ix1853 : inv01 port map ( Y=>nx1852, A=>nx7809);
   ix7810 : aoi222 port map ( Y=>nx7809, A0=>d_arr_mux_18_8, A1=>nx11273, B0
      =>d_arr_mul_18_8, B1=>nx10421, C0=>d_arr_add_18_8, C1=>nx10649);
   lat_d_arr_18_9 : latch port map ( Q=>d_arr_18_9, D=>nx1864, CLK=>nx10189
   );
   ix1865 : inv01 port map ( Y=>nx1864, A=>nx7815);
   ix7816 : aoi222 port map ( Y=>nx7815, A0=>d_arr_mux_18_9, A1=>nx11273, B0
      =>d_arr_mul_18_9, B1=>nx10421, C0=>d_arr_add_18_9, C1=>nx10651);
   lat_d_arr_18_10 : latch port map ( Q=>d_arr_18_10, D=>nx1876, CLK=>
      nx10189);
   ix1877 : inv01 port map ( Y=>nx1876, A=>nx7821);
   ix7822 : aoi222 port map ( Y=>nx7821, A0=>d_arr_mux_18_10, A1=>nx11275, 
      B0=>d_arr_mul_18_10, B1=>nx10421, C0=>d_arr_add_18_10, C1=>nx10651);
   lat_d_arr_18_11 : latch port map ( Q=>d_arr_18_11, D=>nx1888, CLK=>
      nx10191);
   ix1889 : inv01 port map ( Y=>nx1888, A=>nx7827);
   ix7828 : aoi222 port map ( Y=>nx7827, A0=>d_arr_mux_18_11, A1=>nx11275, 
      B0=>d_arr_mul_18_11, B1=>nx10423, C0=>d_arr_add_18_11, C1=>nx10651);
   lat_d_arr_18_12 : latch port map ( Q=>d_arr_18_12, D=>nx1900, CLK=>
      nx10191);
   ix1901 : inv01 port map ( Y=>nx1900, A=>nx7833);
   ix7834 : aoi222 port map ( Y=>nx7833, A0=>d_arr_mux_18_12, A1=>nx11275, 
      B0=>d_arr_mul_18_12, B1=>nx10423, C0=>d_arr_add_18_12, C1=>nx10651);
   lat_d_arr_18_13 : latch port map ( Q=>d_arr_18_13, D=>nx1912, CLK=>
      nx10191);
   ix1913 : inv01 port map ( Y=>nx1912, A=>nx7839);
   ix7840 : aoi222 port map ( Y=>nx7839, A0=>d_arr_mux_18_13, A1=>nx11275, 
      B0=>d_arr_mul_18_13, B1=>nx10423, C0=>d_arr_add_18_13, C1=>nx10651);
   lat_d_arr_18_14 : latch port map ( Q=>d_arr_18_14, D=>nx1924, CLK=>
      nx10191);
   ix1925 : inv01 port map ( Y=>nx1924, A=>nx7845);
   ix7846 : aoi222 port map ( Y=>nx7845, A0=>d_arr_mux_18_14, A1=>nx11275, 
      B0=>d_arr_mul_18_14, B1=>nx10423, C0=>d_arr_add_18_14, C1=>nx10651);
   lat_d_arr_18_15 : latch port map ( Q=>d_arr_18_15, D=>nx1936, CLK=>
      nx10191);
   ix1937 : nand02 port map ( Y=>nx1936, A0=>nx7851, A1=>nx10857);
   ix7852 : aoi22 port map ( Y=>nx7851, A0=>d_arr_mul_18_15, A1=>nx10423, B0
      =>d_arr_add_18_15, B1=>nx10651);
   ix7854 : nand02 port map ( Y=>nx7853, A0=>d_arr_mux_18_31, A1=>nx11275);
   lat_d_arr_18_16 : latch port map ( Q=>d_arr_18_16, D=>nx1946, CLK=>
      nx10191);
   ix1947 : nand02 port map ( Y=>nx1946, A0=>nx7859, A1=>nx10857);
   ix7860 : aoi22 port map ( Y=>nx7859, A0=>d_arr_mul_18_16, A1=>nx10423, B0
      =>d_arr_add_18_16, B1=>nx10653);
   lat_d_arr_18_17 : latch port map ( Q=>d_arr_18_17, D=>nx1956, CLK=>
      nx10191);
   ix1957 : nand02 port map ( Y=>nx1956, A0=>nx7865, A1=>nx10857);
   ix7866 : aoi22 port map ( Y=>nx7865, A0=>d_arr_mul_18_17, A1=>nx10423, B0
      =>d_arr_add_18_17, B1=>nx10653);
   lat_d_arr_18_18 : latch port map ( Q=>d_arr_18_18, D=>nx1966, CLK=>
      nx10193);
   ix1967 : nand02 port map ( Y=>nx1966, A0=>nx7869, A1=>nx10857);
   ix7870 : aoi22 port map ( Y=>nx7869, A0=>d_arr_mul_18_18, A1=>nx10425, B0
      =>d_arr_add_18_18, B1=>nx10653);
   lat_d_arr_18_19 : latch port map ( Q=>d_arr_18_19, D=>nx1976, CLK=>
      nx10193);
   ix1977 : nand02 port map ( Y=>nx1976, A0=>nx7875, A1=>nx10857);
   ix7876 : aoi22 port map ( Y=>nx7875, A0=>d_arr_mul_18_19, A1=>nx10425, B0
      =>d_arr_add_18_19, B1=>nx10653);
   lat_d_arr_18_20 : latch port map ( Q=>d_arr_18_20, D=>nx1986, CLK=>
      nx10193);
   ix1987 : nand02 port map ( Y=>nx1986, A0=>nx7881, A1=>nx10857);
   ix7882 : aoi22 port map ( Y=>nx7881, A0=>d_arr_mul_18_20, A1=>nx10425, B0
      =>d_arr_add_18_20, B1=>nx10653);
   lat_d_arr_18_21 : latch port map ( Q=>d_arr_18_21, D=>nx1996, CLK=>
      nx10193);
   ix1997 : nand02 port map ( Y=>nx1996, A0=>nx7887, A1=>nx10857);
   ix7888 : aoi22 port map ( Y=>nx7887, A0=>d_arr_mul_18_21, A1=>nx10425, B0
      =>d_arr_add_18_21, B1=>nx10653);
   lat_d_arr_18_22 : latch port map ( Q=>d_arr_18_22, D=>nx2006, CLK=>
      nx10193);
   ix2007 : nand02 port map ( Y=>nx2006, A0=>nx7893, A1=>nx10859);
   ix7894 : aoi22 port map ( Y=>nx7893, A0=>d_arr_mul_18_22, A1=>nx10425, B0
      =>d_arr_add_18_22, B1=>nx10653);
   lat_d_arr_18_23 : latch port map ( Q=>d_arr_18_23, D=>nx2016, CLK=>
      nx10193);
   ix2017 : nand02 port map ( Y=>nx2016, A0=>nx7899, A1=>nx10859);
   ix7900 : aoi22 port map ( Y=>nx7899, A0=>d_arr_mul_18_23, A1=>nx10425, B0
      =>d_arr_add_18_23, B1=>nx10655);
   lat_d_arr_18_24 : latch port map ( Q=>d_arr_18_24, D=>nx2026, CLK=>
      nx10193);
   ix2027 : nand02 port map ( Y=>nx2026, A0=>nx7905, A1=>nx10859);
   ix7906 : aoi22 port map ( Y=>nx7905, A0=>d_arr_mul_18_24, A1=>nx10425, B0
      =>d_arr_add_18_24, B1=>nx10655);
   lat_d_arr_18_25 : latch port map ( Q=>d_arr_18_25, D=>nx2036, CLK=>
      nx10195);
   ix2037 : nand02 port map ( Y=>nx2036, A0=>nx7911, A1=>nx10859);
   ix7912 : aoi22 port map ( Y=>nx7911, A0=>d_arr_mul_18_25, A1=>nx10427, B0
      =>d_arr_add_18_25, B1=>nx10655);
   lat_d_arr_18_26 : latch port map ( Q=>d_arr_18_26, D=>nx2046, CLK=>
      nx10195);
   ix2047 : nand02 port map ( Y=>nx2046, A0=>nx7917, A1=>nx10859);
   ix7918 : aoi22 port map ( Y=>nx7917, A0=>d_arr_mul_18_26, A1=>nx10427, B0
      =>d_arr_add_18_26, B1=>nx10655);
   lat_d_arr_18_27 : latch port map ( Q=>d_arr_18_27, D=>nx2056, CLK=>
      nx10195);
   ix2057 : nand02 port map ( Y=>nx2056, A0=>nx7923, A1=>nx10859);
   ix7924 : aoi22 port map ( Y=>nx7923, A0=>d_arr_mul_18_27, A1=>nx10427, B0
      =>d_arr_add_18_27, B1=>nx10655);
   lat_d_arr_18_28 : latch port map ( Q=>d_arr_18_28, D=>nx2066, CLK=>
      nx10195);
   ix2067 : nand02 port map ( Y=>nx2066, A0=>nx7929, A1=>nx10859);
   ix7930 : aoi22 port map ( Y=>nx7929, A0=>d_arr_mul_18_28, A1=>nx10427, B0
      =>d_arr_add_18_28, B1=>nx10655);
   lat_d_arr_18_29 : latch port map ( Q=>d_arr_18_29, D=>nx2076, CLK=>
      nx10195);
   ix2077 : nand02 port map ( Y=>nx2076, A0=>nx7935, A1=>nx7853);
   ix7936 : aoi22 port map ( Y=>nx7935, A0=>d_arr_mul_18_29, A1=>nx10427, B0
      =>d_arr_add_18_29, B1=>nx10655);
   lat_d_arr_18_30 : latch port map ( Q=>d_arr_18_30, D=>nx2086, CLK=>
      nx10195);
   ix2087 : nand02 port map ( Y=>nx2086, A0=>nx7941, A1=>nx7853);
   ix7942 : aoi22 port map ( Y=>nx7941, A0=>d_arr_mul_18_30, A1=>nx10427, B0
      =>d_arr_add_18_30, B1=>nx10657);
   lat_d_arr_18_31 : latch port map ( Q=>d_arr_18_31, D=>nx2096, CLK=>
      nx10195);
   ix2097 : nand02 port map ( Y=>nx2096, A0=>nx7947, A1=>nx7853);
   ix7948 : aoi22 port map ( Y=>nx7947, A0=>d_arr_mul_18_31, A1=>nx10427, B0
      =>d_arr_add_18_31, B1=>nx10657);
   lat_d_arr_17_0 : latch port map ( Q=>d_arr_17_0, D=>nx2104, CLK=>nx10197
   );
   ix2105 : ao22 port map ( Y=>nx2104, A0=>d_arr_mux_17_0, A1=>nx11275, B0=>
      d_arr_mul_17_0, B1=>nx10429);
   lat_d_arr_17_1 : latch port map ( Q=>d_arr_17_1, D=>nx2112, CLK=>nx10197
   );
   ix2113 : ao22 port map ( Y=>nx2112, A0=>d_arr_mux_17_1, A1=>nx11277, B0=>
      d_arr_mul_17_1, B1=>nx10429);
   lat_d_arr_17_2 : latch port map ( Q=>d_arr_17_2, D=>nx2120, CLK=>nx10197
   );
   ix2121 : ao22 port map ( Y=>nx2120, A0=>d_arr_mux_17_2, A1=>nx11277, B0=>
      d_arr_mul_17_2, B1=>nx10429);
   lat_d_arr_17_3 : latch port map ( Q=>d_arr_17_3, D=>nx2128, CLK=>nx10197
   );
   ix2129 : ao22 port map ( Y=>nx2128, A0=>d_arr_mux_17_3, A1=>nx11277, B0=>
      d_arr_mul_17_3, B1=>nx10429);
   lat_d_arr_17_4 : latch port map ( Q=>d_arr_17_4, D=>nx2136, CLK=>nx10197
   );
   ix2137 : ao22 port map ( Y=>nx2136, A0=>d_arr_mux_17_4, A1=>nx11277, B0=>
      d_arr_mul_17_4, B1=>nx10429);
   lat_d_arr_17_5 : latch port map ( Q=>d_arr_17_5, D=>nx2144, CLK=>nx10197
   );
   ix2145 : ao22 port map ( Y=>nx2144, A0=>d_arr_mux_17_5, A1=>nx11277, B0=>
      d_arr_mul_17_5, B1=>nx10429);
   lat_d_arr_17_6 : latch port map ( Q=>d_arr_17_6, D=>nx2152, CLK=>nx10197
   );
   ix2153 : ao22 port map ( Y=>nx2152, A0=>d_arr_mux_17_6, A1=>nx11277, B0=>
      d_arr_mul_17_6, B1=>nx10429);
   lat_d_arr_17_7 : latch port map ( Q=>d_arr_17_7, D=>nx2160, CLK=>nx10199
   );
   ix2161 : ao22 port map ( Y=>nx2160, A0=>d_arr_mux_17_7, A1=>nx11277, B0=>
      d_arr_mul_17_7, B1=>nx10431);
   lat_d_arr_17_8 : latch port map ( Q=>d_arr_17_8, D=>nx2168, CLK=>nx10199
   );
   ix2169 : ao22 port map ( Y=>nx2168, A0=>d_arr_mux_17_8, A1=>nx11279, B0=>
      d_arr_mul_17_8, B1=>nx10431);
   lat_d_arr_17_9 : latch port map ( Q=>d_arr_17_9, D=>nx2176, CLK=>nx10199
   );
   ix2177 : ao22 port map ( Y=>nx2176, A0=>d_arr_mux_17_9, A1=>nx11279, B0=>
      d_arr_mul_17_9, B1=>nx10431);
   lat_d_arr_17_10 : latch port map ( Q=>d_arr_17_10, D=>nx2184, CLK=>
      nx10199);
   ix2185 : ao22 port map ( Y=>nx2184, A0=>d_arr_mux_17_10, A1=>nx11279, B0
      =>d_arr_mul_17_10, B1=>nx10431);
   lat_d_arr_17_11 : latch port map ( Q=>d_arr_17_11, D=>nx2192, CLK=>
      nx10199);
   ix2193 : ao22 port map ( Y=>nx2192, A0=>d_arr_mux_17_11, A1=>nx11279, B0
      =>d_arr_mul_17_11, B1=>nx10431);
   lat_d_arr_17_12 : latch port map ( Q=>d_arr_17_12, D=>nx2200, CLK=>
      nx10199);
   ix2201 : ao22 port map ( Y=>nx2200, A0=>d_arr_mux_17_12, A1=>nx11279, B0
      =>d_arr_mul_17_12, B1=>nx10431);
   lat_d_arr_17_13 : latch port map ( Q=>d_arr_17_13, D=>nx2208, CLK=>
      nx10199);
   ix2209 : ao22 port map ( Y=>nx2208, A0=>d_arr_mux_17_13, A1=>nx11279, B0
      =>d_arr_mul_17_13, B1=>nx10431);
   lat_d_arr_17_14 : latch port map ( Q=>d_arr_17_14, D=>nx2216, CLK=>
      nx10201);
   ix2217 : ao22 port map ( Y=>nx2216, A0=>d_arr_mux_17_14, A1=>nx11279, B0
      =>d_arr_mul_17_14, B1=>nx10433);
   lat_d_arr_17_15 : latch port map ( Q=>d_arr_17_15, D=>nx2224, CLK=>
      nx10201);
   ix2225 : ao22 port map ( Y=>nx2224, A0=>d_arr_mux_17_15, A1=>nx11281, B0
      =>d_arr_mul_17_15, B1=>nx10433);
   lat_d_arr_17_16 : latch port map ( Q=>d_arr_17_16, D=>nx2232, CLK=>
      nx10201);
   ix2233 : ao22 port map ( Y=>nx2232, A0=>d_arr_mux_17_16, A1=>nx11281, B0
      =>d_arr_mul_17_16, B1=>nx10433);
   lat_d_arr_17_17 : latch port map ( Q=>d_arr_17_17, D=>nx2240, CLK=>
      nx10201);
   ix2241 : ao22 port map ( Y=>nx2240, A0=>d_arr_mux_17_17, A1=>nx11281, B0
      =>d_arr_mul_17_17, B1=>nx10433);
   lat_d_arr_17_18 : latch port map ( Q=>d_arr_17_18, D=>nx2248, CLK=>
      nx10201);
   ix2249 : ao22 port map ( Y=>nx2248, A0=>d_arr_mux_17_18, A1=>nx11281, B0
      =>d_arr_mul_17_18, B1=>nx10433);
   lat_d_arr_17_19 : latch port map ( Q=>d_arr_17_19, D=>nx2256, CLK=>
      nx10201);
   ix2257 : ao22 port map ( Y=>nx2256, A0=>d_arr_mux_17_19, A1=>nx11281, B0
      =>d_arr_mul_17_19, B1=>nx10433);
   lat_d_arr_17_20 : latch port map ( Q=>d_arr_17_20, D=>nx2264, CLK=>
      nx10201);
   ix2265 : ao22 port map ( Y=>nx2264, A0=>d_arr_mux_17_20, A1=>nx11281, B0
      =>d_arr_mul_17_20, B1=>nx10433);
   lat_d_arr_17_21 : latch port map ( Q=>d_arr_17_21, D=>nx2272, CLK=>
      nx10203);
   ix2273 : ao22 port map ( Y=>nx2272, A0=>d_arr_mux_17_21, A1=>nx11281, B0
      =>d_arr_mul_17_21, B1=>nx10435);
   lat_d_arr_17_22 : latch port map ( Q=>d_arr_17_22, D=>nx2280, CLK=>
      nx10203);
   ix2281 : ao22 port map ( Y=>nx2280, A0=>d_arr_mux_17_22, A1=>nx11283, B0
      =>d_arr_mul_17_22, B1=>nx10435);
   lat_d_arr_17_23 : latch port map ( Q=>d_arr_17_23, D=>nx2288, CLK=>
      nx10203);
   ix2289 : ao22 port map ( Y=>nx2288, A0=>d_arr_mux_17_23, A1=>nx11283, B0
      =>d_arr_mul_17_23, B1=>nx10435);
   lat_d_arr_17_24 : latch port map ( Q=>d_arr_17_24, D=>nx2296, CLK=>
      nx10203);
   ix2297 : ao22 port map ( Y=>nx2296, A0=>d_arr_mux_17_24, A1=>nx11283, B0
      =>d_arr_mul_17_24, B1=>nx10435);
   lat_d_arr_17_25 : latch port map ( Q=>d_arr_17_25, D=>nx2304, CLK=>
      nx10203);
   ix2305 : ao22 port map ( Y=>nx2304, A0=>d_arr_mux_17_25, A1=>nx11283, B0
      =>d_arr_mul_17_25, B1=>nx10435);
   lat_d_arr_17_26 : latch port map ( Q=>d_arr_17_26, D=>nx2312, CLK=>
      nx10203);
   ix2313 : ao22 port map ( Y=>nx2312, A0=>d_arr_mux_17_26, A1=>nx11283, B0
      =>d_arr_mul_17_26, B1=>nx10435);
   lat_d_arr_17_27 : latch port map ( Q=>d_arr_17_27, D=>nx2320, CLK=>
      nx10203);
   ix2321 : ao22 port map ( Y=>nx2320, A0=>d_arr_mux_17_27, A1=>nx11283, B0
      =>d_arr_mul_17_27, B1=>nx10435);
   lat_d_arr_17_28 : latch port map ( Q=>d_arr_17_28, D=>nx2328, CLK=>
      nx10205);
   ix2329 : ao22 port map ( Y=>nx2328, A0=>d_arr_mux_17_28, A1=>nx11283, B0
      =>d_arr_mul_17_28, B1=>nx10437);
   lat_d_arr_17_29 : latch port map ( Q=>d_arr_17_29, D=>nx2336, CLK=>
      nx10205);
   ix2337 : ao22 port map ( Y=>nx2336, A0=>d_arr_mux_17_29, A1=>nx11285, B0
      =>d_arr_mul_17_29, B1=>nx10437);
   lat_d_arr_17_30 : latch port map ( Q=>d_arr_17_30, D=>nx2344, CLK=>
      nx10205);
   ix2345 : ao22 port map ( Y=>nx2344, A0=>d_arr_mux_17_30, A1=>nx11285, B0
      =>d_arr_mul_17_30, B1=>nx10437);
   lat_d_arr_17_31 : latch port map ( Q=>d_arr_17_31, D=>nx2352, CLK=>
      nx10205);
   ix2353 : ao22 port map ( Y=>nx2352, A0=>d_arr_mux_17_31, A1=>nx11285, B0
      =>d_arr_mul_17_31, B1=>nx10437);
   lat_d_arr_16_0 : latch port map ( Q=>d_arr_16_0, D=>nx2360, CLK=>nx10205
   );
   ix2361 : ao22 port map ( Y=>nx2360, A0=>d_arr_mux_16_0, A1=>nx11285, B0=>
      d_arr_mul_16_0, B1=>nx10437);
   lat_d_arr_16_1 : latch port map ( Q=>d_arr_16_1, D=>nx2368, CLK=>nx10205
   );
   ix2369 : ao22 port map ( Y=>nx2368, A0=>d_arr_mux_16_1, A1=>nx11285, B0=>
      d_arr_mul_16_1, B1=>nx10437);
   lat_d_arr_16_2 : latch port map ( Q=>d_arr_16_2, D=>nx2376, CLK=>nx10205
   );
   ix2377 : ao22 port map ( Y=>nx2376, A0=>d_arr_mux_16_2, A1=>nx11285, B0=>
      d_arr_mul_16_2, B1=>nx10437);
   lat_d_arr_16_3 : latch port map ( Q=>d_arr_16_3, D=>nx2384, CLK=>nx10207
   );
   ix2385 : ao22 port map ( Y=>nx2384, A0=>d_arr_mux_16_3, A1=>nx11285, B0=>
      d_arr_mul_16_3, B1=>nx10439);
   lat_d_arr_16_4 : latch port map ( Q=>d_arr_16_4, D=>nx2392, CLK=>nx10207
   );
   ix2393 : ao22 port map ( Y=>nx2392, A0=>d_arr_mux_16_4, A1=>nx11287, B0=>
      d_arr_mul_16_4, B1=>nx10439);
   lat_d_arr_16_5 : latch port map ( Q=>d_arr_16_5, D=>nx2400, CLK=>nx10207
   );
   ix2401 : ao22 port map ( Y=>nx2400, A0=>d_arr_mux_16_5, A1=>nx11287, B0=>
      d_arr_mul_16_5, B1=>nx10439);
   lat_d_arr_16_6 : latch port map ( Q=>d_arr_16_6, D=>nx2408, CLK=>nx10207
   );
   ix2409 : ao22 port map ( Y=>nx2408, A0=>d_arr_mux_16_6, A1=>nx11287, B0=>
      d_arr_mul_16_6, B1=>nx10439);
   lat_d_arr_16_7 : latch port map ( Q=>d_arr_16_7, D=>nx2416, CLK=>nx10207
   );
   ix2417 : ao22 port map ( Y=>nx2416, A0=>d_arr_mux_16_7, A1=>nx11287, B0=>
      d_arr_mul_16_7, B1=>nx10439);
   lat_d_arr_16_8 : latch port map ( Q=>d_arr_16_8, D=>nx2424, CLK=>nx10207
   );
   ix2425 : ao22 port map ( Y=>nx2424, A0=>d_arr_mux_16_8, A1=>nx11287, B0=>
      d_arr_mul_16_8, B1=>nx10439);
   lat_d_arr_16_9 : latch port map ( Q=>d_arr_16_9, D=>nx2432, CLK=>nx10207
   );
   ix2433 : ao22 port map ( Y=>nx2432, A0=>d_arr_mux_16_9, A1=>nx11287, B0=>
      d_arr_mul_16_9, B1=>nx10439);
   lat_d_arr_16_10 : latch port map ( Q=>d_arr_16_10, D=>nx2440, CLK=>
      nx10209);
   ix2441 : ao22 port map ( Y=>nx2440, A0=>d_arr_mux_16_10, A1=>nx11287, B0
      =>d_arr_mul_16_10, B1=>nx10441);
   lat_d_arr_16_11 : latch port map ( Q=>d_arr_16_11, D=>nx2448, CLK=>
      nx10209);
   ix2449 : ao22 port map ( Y=>nx2448, A0=>d_arr_mux_16_11, A1=>nx11289, B0
      =>d_arr_mul_16_11, B1=>nx10441);
   lat_d_arr_16_12 : latch port map ( Q=>d_arr_16_12, D=>nx2456, CLK=>
      nx10209);
   ix2457 : ao22 port map ( Y=>nx2456, A0=>d_arr_mux_16_12, A1=>nx11289, B0
      =>d_arr_mul_16_12, B1=>nx10441);
   lat_d_arr_16_13 : latch port map ( Q=>d_arr_16_13, D=>nx2464, CLK=>
      nx10209);
   ix2465 : ao22 port map ( Y=>nx2464, A0=>d_arr_mux_16_13, A1=>nx11289, B0
      =>d_arr_mul_16_13, B1=>nx10441);
   lat_d_arr_16_14 : latch port map ( Q=>d_arr_16_14, D=>nx2472, CLK=>
      nx10209);
   ix2473 : ao22 port map ( Y=>nx2472, A0=>d_arr_mux_16_14, A1=>nx11289, B0
      =>d_arr_mul_16_14, B1=>nx10441);
   lat_d_arr_16_15 : latch port map ( Q=>d_arr_16_15, D=>nx2480, CLK=>
      nx10209);
   ix2481 : ao22 port map ( Y=>nx2480, A0=>d_arr_mux_16_15, A1=>nx11289, B0
      =>d_arr_mul_16_15, B1=>nx10441);
   lat_d_arr_16_16 : latch port map ( Q=>d_arr_16_16, D=>nx2488, CLK=>
      nx10209);
   ix2489 : ao22 port map ( Y=>nx2488, A0=>d_arr_mux_16_16, A1=>nx11289, B0
      =>d_arr_mul_16_16, B1=>nx10441);
   lat_d_arr_16_17 : latch port map ( Q=>d_arr_16_17, D=>nx2496, CLK=>
      nx10211);
   ix2497 : ao22 port map ( Y=>nx2496, A0=>d_arr_mux_16_17, A1=>nx11289, B0
      =>d_arr_mul_16_17, B1=>nx10443);
   lat_d_arr_16_18 : latch port map ( Q=>d_arr_16_18, D=>nx2504, CLK=>
      nx10211);
   ix2505 : ao22 port map ( Y=>nx2504, A0=>d_arr_mux_16_18, A1=>nx11291, B0
      =>d_arr_mul_16_18, B1=>nx10443);
   lat_d_arr_16_19 : latch port map ( Q=>d_arr_16_19, D=>nx2512, CLK=>
      nx10211);
   ix2513 : ao22 port map ( Y=>nx2512, A0=>d_arr_mux_16_19, A1=>nx11291, B0
      =>d_arr_mul_16_19, B1=>nx10443);
   lat_d_arr_16_20 : latch port map ( Q=>d_arr_16_20, D=>nx2520, CLK=>
      nx10211);
   ix2521 : ao22 port map ( Y=>nx2520, A0=>d_arr_mux_16_20, A1=>nx11291, B0
      =>d_arr_mul_16_20, B1=>nx10443);
   lat_d_arr_16_21 : latch port map ( Q=>d_arr_16_21, D=>nx2528, CLK=>
      nx10211);
   ix2529 : ao22 port map ( Y=>nx2528, A0=>d_arr_mux_16_21, A1=>nx11291, B0
      =>d_arr_mul_16_21, B1=>nx10443);
   lat_d_arr_16_22 : latch port map ( Q=>d_arr_16_22, D=>nx2536, CLK=>
      nx10211);
   ix2537 : ao22 port map ( Y=>nx2536, A0=>d_arr_mux_16_22, A1=>nx11291, B0
      =>d_arr_mul_16_22, B1=>nx10443);
   lat_d_arr_16_23 : latch port map ( Q=>d_arr_16_23, D=>nx2544, CLK=>
      nx10211);
   ix2545 : ao22 port map ( Y=>nx2544, A0=>d_arr_mux_16_23, A1=>nx11291, B0
      =>d_arr_mul_16_23, B1=>nx10443);
   lat_d_arr_16_24 : latch port map ( Q=>d_arr_16_24, D=>nx2552, CLK=>
      nx10213);
   ix2553 : ao22 port map ( Y=>nx2552, A0=>d_arr_mux_16_24, A1=>nx11291, B0
      =>d_arr_mul_16_24, B1=>nx10445);
   lat_d_arr_16_25 : latch port map ( Q=>d_arr_16_25, D=>nx2560, CLK=>
      nx10213);
   ix2561 : ao22 port map ( Y=>nx2560, A0=>d_arr_mux_16_25, A1=>nx11293, B0
      =>d_arr_mul_16_25, B1=>nx10445);
   lat_d_arr_16_26 : latch port map ( Q=>d_arr_16_26, D=>nx2568, CLK=>
      nx10213);
   ix2569 : ao22 port map ( Y=>nx2568, A0=>d_arr_mux_16_26, A1=>nx11293, B0
      =>d_arr_mul_16_26, B1=>nx10445);
   lat_d_arr_16_27 : latch port map ( Q=>d_arr_16_27, D=>nx2576, CLK=>
      nx10213);
   ix2577 : ao22 port map ( Y=>nx2576, A0=>d_arr_mux_16_27, A1=>nx11293, B0
      =>d_arr_mul_16_27, B1=>nx10445);
   lat_d_arr_16_28 : latch port map ( Q=>d_arr_16_28, D=>nx2584, CLK=>
      nx10213);
   ix2585 : ao22 port map ( Y=>nx2584, A0=>d_arr_mux_16_28, A1=>nx11293, B0
      =>d_arr_mul_16_28, B1=>nx10445);
   lat_d_arr_16_29 : latch port map ( Q=>d_arr_16_29, D=>nx2592, CLK=>
      nx10213);
   ix2593 : ao22 port map ( Y=>nx2592, A0=>d_arr_mux_16_29, A1=>nx11293, B0
      =>d_arr_mul_16_29, B1=>nx10445);
   lat_d_arr_16_30 : latch port map ( Q=>d_arr_16_30, D=>nx2600, CLK=>
      nx10213);
   ix2601 : ao22 port map ( Y=>nx2600, A0=>d_arr_mux_16_30, A1=>nx11293, B0
      =>d_arr_mul_16_30, B1=>nx10445);
   lat_d_arr_16_31 : latch port map ( Q=>d_arr_16_31, D=>nx2608, CLK=>
      nx10215);
   ix2609 : ao22 port map ( Y=>nx2608, A0=>d_arr_mux_16_31, A1=>nx11293, B0
      =>d_arr_mul_16_31, B1=>nx10447);
   lat_d_arr_15_0 : latch port map ( Q=>d_arr_15_0, D=>nx2616, CLK=>nx10215
   );
   ix2617 : ao22 port map ( Y=>nx2616, A0=>d_arr_mux_15_0, A1=>nx11295, B0=>
      d_arr_mul_15_0, B1=>nx10447);
   lat_d_arr_15_1 : latch port map ( Q=>d_arr_15_1, D=>nx2624, CLK=>nx10215
   );
   ix2625 : ao22 port map ( Y=>nx2624, A0=>d_arr_mux_15_1, A1=>nx11295, B0=>
      d_arr_mul_15_1, B1=>nx10447);
   lat_d_arr_15_2 : latch port map ( Q=>d_arr_15_2, D=>nx2632, CLK=>nx10215
   );
   ix2633 : ao22 port map ( Y=>nx2632, A0=>d_arr_mux_15_2, A1=>nx11295, B0=>
      d_arr_mul_15_2, B1=>nx10447);
   lat_d_arr_15_3 : latch port map ( Q=>d_arr_15_3, D=>nx2640, CLK=>nx10215
   );
   ix2641 : ao22 port map ( Y=>nx2640, A0=>d_arr_mux_15_3, A1=>nx11295, B0=>
      d_arr_mul_15_3, B1=>nx10447);
   lat_d_arr_15_4 : latch port map ( Q=>d_arr_15_4, D=>nx2648, CLK=>nx10215
   );
   ix2649 : ao22 port map ( Y=>nx2648, A0=>d_arr_mux_15_4, A1=>nx11295, B0=>
      d_arr_mul_15_4, B1=>nx10447);
   lat_d_arr_15_5 : latch port map ( Q=>d_arr_15_5, D=>nx2656, CLK=>nx10215
   );
   ix2657 : ao22 port map ( Y=>nx2656, A0=>d_arr_mux_15_5, A1=>nx11295, B0=>
      d_arr_mul_15_5, B1=>nx10447);
   lat_d_arr_15_6 : latch port map ( Q=>d_arr_15_6, D=>nx2664, CLK=>nx10217
   );
   ix2665 : ao22 port map ( Y=>nx2664, A0=>d_arr_mux_15_6, A1=>nx11295, B0=>
      d_arr_mul_15_6, B1=>nx10449);
   lat_d_arr_15_7 : latch port map ( Q=>d_arr_15_7, D=>nx2672, CLK=>nx10217
   );
   ix2673 : ao22 port map ( Y=>nx2672, A0=>d_arr_mux_15_7, A1=>nx11297, B0=>
      d_arr_mul_15_7, B1=>nx10449);
   lat_d_arr_15_8 : latch port map ( Q=>d_arr_15_8, D=>nx2680, CLK=>nx10217
   );
   ix2681 : ao22 port map ( Y=>nx2680, A0=>d_arr_mux_15_8, A1=>nx11297, B0=>
      d_arr_mul_15_8, B1=>nx10449);
   lat_d_arr_15_9 : latch port map ( Q=>d_arr_15_9, D=>nx2688, CLK=>nx10217
   );
   ix2689 : ao22 port map ( Y=>nx2688, A0=>d_arr_mux_15_9, A1=>nx11297, B0=>
      d_arr_mul_15_9, B1=>nx10449);
   lat_d_arr_15_10 : latch port map ( Q=>d_arr_15_10, D=>nx2696, CLK=>
      nx10217);
   ix2697 : ao22 port map ( Y=>nx2696, A0=>d_arr_mux_15_10, A1=>nx11297, B0
      =>d_arr_mul_15_10, B1=>nx10449);
   lat_d_arr_15_11 : latch port map ( Q=>d_arr_15_11, D=>nx2704, CLK=>
      nx10217);
   ix2705 : ao22 port map ( Y=>nx2704, A0=>d_arr_mux_15_11, A1=>nx11297, B0
      =>d_arr_mul_15_11, B1=>nx10449);
   lat_d_arr_15_12 : latch port map ( Q=>d_arr_15_12, D=>nx2712, CLK=>
      nx10217);
   ix2713 : ao22 port map ( Y=>nx2712, A0=>d_arr_mux_15_12, A1=>nx11297, B0
      =>d_arr_mul_15_12, B1=>nx10449);
   lat_d_arr_15_13 : latch port map ( Q=>d_arr_15_13, D=>nx2720, CLK=>
      nx10219);
   ix2721 : ao22 port map ( Y=>nx2720, A0=>d_arr_mux_15_13, A1=>nx11297, B0
      =>d_arr_mul_15_13, B1=>nx10451);
   lat_d_arr_15_14 : latch port map ( Q=>d_arr_15_14, D=>nx2728, CLK=>
      nx10219);
   ix2729 : ao22 port map ( Y=>nx2728, A0=>d_arr_mux_15_14, A1=>nx11299, B0
      =>d_arr_mul_15_14, B1=>nx10451);
   lat_d_arr_15_15 : latch port map ( Q=>d_arr_15_15, D=>nx2736, CLK=>
      nx10219);
   ix2737 : ao22 port map ( Y=>nx2736, A0=>d_arr_mux_15_15, A1=>nx11299, B0
      =>d_arr_mul_15_15, B1=>nx10451);
   lat_d_arr_15_16 : latch port map ( Q=>d_arr_15_16, D=>nx2744, CLK=>
      nx10219);
   ix2745 : ao22 port map ( Y=>nx2744, A0=>d_arr_mux_15_16, A1=>nx11299, B0
      =>d_arr_mul_15_16, B1=>nx10451);
   lat_d_arr_15_17 : latch port map ( Q=>d_arr_15_17, D=>nx2752, CLK=>
      nx10219);
   ix2753 : ao22 port map ( Y=>nx2752, A0=>d_arr_mux_15_17, A1=>nx11299, B0
      =>d_arr_mul_15_17, B1=>nx10451);
   lat_d_arr_15_18 : latch port map ( Q=>d_arr_15_18, D=>nx2760, CLK=>
      nx10219);
   ix2761 : ao22 port map ( Y=>nx2760, A0=>d_arr_mux_15_18, A1=>nx11299, B0
      =>d_arr_mul_15_18, B1=>nx10451);
   lat_d_arr_15_19 : latch port map ( Q=>d_arr_15_19, D=>nx2768, CLK=>
      nx10219);
   ix2769 : ao22 port map ( Y=>nx2768, A0=>d_arr_mux_15_19, A1=>nx11299, B0
      =>d_arr_mul_15_19, B1=>nx10451);
   lat_d_arr_15_20 : latch port map ( Q=>d_arr_15_20, D=>nx2776, CLK=>
      nx10221);
   ix2777 : ao22 port map ( Y=>nx2776, A0=>d_arr_mux_15_20, A1=>nx11299, B0
      =>d_arr_mul_15_20, B1=>nx10453);
   lat_d_arr_15_21 : latch port map ( Q=>d_arr_15_21, D=>nx2784, CLK=>
      nx10221);
   ix2785 : ao22 port map ( Y=>nx2784, A0=>d_arr_mux_15_21, A1=>nx11301, B0
      =>d_arr_mul_15_21, B1=>nx10453);
   lat_d_arr_15_22 : latch port map ( Q=>d_arr_15_22, D=>nx2792, CLK=>
      nx10221);
   ix2793 : ao22 port map ( Y=>nx2792, A0=>d_arr_mux_15_22, A1=>nx11301, B0
      =>d_arr_mul_15_22, B1=>nx10453);
   lat_d_arr_15_23 : latch port map ( Q=>d_arr_15_23, D=>nx2800, CLK=>
      nx10221);
   ix2801 : ao22 port map ( Y=>nx2800, A0=>d_arr_mux_15_23, A1=>nx11301, B0
      =>d_arr_mul_15_23, B1=>nx10453);
   lat_d_arr_15_24 : latch port map ( Q=>d_arr_15_24, D=>nx2808, CLK=>
      nx10221);
   ix2809 : ao22 port map ( Y=>nx2808, A0=>d_arr_mux_15_24, A1=>nx11301, B0
      =>d_arr_mul_15_24, B1=>nx10453);
   lat_d_arr_15_25 : latch port map ( Q=>d_arr_15_25, D=>nx2816, CLK=>
      nx10221);
   ix2817 : ao22 port map ( Y=>nx2816, A0=>d_arr_mux_15_25, A1=>nx11301, B0
      =>d_arr_mul_15_25, B1=>nx10453);
   lat_d_arr_15_26 : latch port map ( Q=>d_arr_15_26, D=>nx2824, CLK=>
      nx10221);
   ix2825 : ao22 port map ( Y=>nx2824, A0=>d_arr_mux_15_26, A1=>nx11301, B0
      =>d_arr_mul_15_26, B1=>nx10453);
   lat_d_arr_15_27 : latch port map ( Q=>d_arr_15_27, D=>nx2832, CLK=>
      nx10223);
   ix2833 : ao22 port map ( Y=>nx2832, A0=>d_arr_mux_15_27, A1=>nx11301, B0
      =>d_arr_mul_15_27, B1=>nx10455);
   lat_d_arr_15_28 : latch port map ( Q=>d_arr_15_28, D=>nx2840, CLK=>
      nx10223);
   ix2841 : ao22 port map ( Y=>nx2840, A0=>d_arr_mux_15_28, A1=>nx11303, B0
      =>d_arr_mul_15_28, B1=>nx10455);
   lat_d_arr_15_29 : latch port map ( Q=>d_arr_15_29, D=>nx2848, CLK=>
      nx10223);
   ix2849 : ao22 port map ( Y=>nx2848, A0=>d_arr_mux_15_29, A1=>nx11303, B0
      =>d_arr_mul_15_29, B1=>nx10455);
   lat_d_arr_15_30 : latch port map ( Q=>d_arr_15_30, D=>nx2856, CLK=>
      nx10223);
   ix2857 : ao22 port map ( Y=>nx2856, A0=>d_arr_mux_15_30, A1=>nx11303, B0
      =>d_arr_mul_15_30, B1=>nx10455);
   lat_d_arr_15_31 : latch port map ( Q=>d_arr_15_31, D=>nx2864, CLK=>
      nx10223);
   ix2865 : ao22 port map ( Y=>nx2864, A0=>d_arr_mux_15_31, A1=>nx11303, B0
      =>d_arr_mul_15_31, B1=>nx10455);
   lat_d_arr_14_0 : latch port map ( Q=>d_arr_14_0, D=>nx2872, CLK=>nx10223
   );
   ix2873 : ao22 port map ( Y=>nx2872, A0=>d_arr_mux_14_0, A1=>nx11303, B0=>
      d_arr_mul_14_0, B1=>nx10455);
   lat_d_arr_14_1 : latch port map ( Q=>d_arr_14_1, D=>nx2880, CLK=>nx10223
   );
   ix2881 : ao22 port map ( Y=>nx2880, A0=>d_arr_mux_14_1, A1=>nx11303, B0=>
      d_arr_mul_14_1, B1=>nx10455);
   lat_d_arr_14_2 : latch port map ( Q=>d_arr_14_2, D=>nx2888, CLK=>nx10225
   );
   ix2889 : ao22 port map ( Y=>nx2888, A0=>d_arr_mux_14_2, A1=>nx11303, B0=>
      d_arr_mul_14_2, B1=>nx10457);
   lat_d_arr_14_3 : latch port map ( Q=>d_arr_14_3, D=>nx2896, CLK=>nx10225
   );
   ix2897 : ao22 port map ( Y=>nx2896, A0=>d_arr_mux_14_3, A1=>nx11305, B0=>
      d_arr_mul_14_3, B1=>nx10457);
   lat_d_arr_14_4 : latch port map ( Q=>d_arr_14_4, D=>nx2904, CLK=>nx10225
   );
   ix2905 : ao22 port map ( Y=>nx2904, A0=>d_arr_mux_14_4, A1=>nx11305, B0=>
      d_arr_mul_14_4, B1=>nx10457);
   lat_d_arr_14_5 : latch port map ( Q=>d_arr_14_5, D=>nx2912, CLK=>nx10225
   );
   ix2913 : ao22 port map ( Y=>nx2912, A0=>d_arr_mux_14_5, A1=>nx11305, B0=>
      d_arr_mul_14_5, B1=>nx10457);
   lat_d_arr_14_6 : latch port map ( Q=>d_arr_14_6, D=>nx2920, CLK=>nx10225
   );
   ix2921 : ao22 port map ( Y=>nx2920, A0=>d_arr_mux_14_6, A1=>nx11305, B0=>
      d_arr_mul_14_6, B1=>nx10457);
   lat_d_arr_14_7 : latch port map ( Q=>d_arr_14_7, D=>nx2928, CLK=>nx10225
   );
   ix2929 : ao22 port map ( Y=>nx2928, A0=>d_arr_mux_14_7, A1=>nx11305, B0=>
      d_arr_mul_14_7, B1=>nx10457);
   lat_d_arr_14_8 : latch port map ( Q=>d_arr_14_8, D=>nx2936, CLK=>nx10225
   );
   ix2937 : ao22 port map ( Y=>nx2936, A0=>d_arr_mux_14_8, A1=>nx11305, B0=>
      d_arr_mul_14_8, B1=>nx10457);
   lat_d_arr_14_9 : latch port map ( Q=>d_arr_14_9, D=>nx2944, CLK=>nx10227
   );
   ix2945 : ao22 port map ( Y=>nx2944, A0=>d_arr_mux_14_9, A1=>nx11305, B0=>
      d_arr_mul_14_9, B1=>nx10459);
   lat_d_arr_14_10 : latch port map ( Q=>d_arr_14_10, D=>nx2952, CLK=>
      nx10227);
   ix2953 : ao22 port map ( Y=>nx2952, A0=>d_arr_mux_14_10, A1=>nx11307, B0
      =>d_arr_mul_14_10, B1=>nx10459);
   lat_d_arr_14_11 : latch port map ( Q=>d_arr_14_11, D=>nx2960, CLK=>
      nx10227);
   ix2961 : ao22 port map ( Y=>nx2960, A0=>d_arr_mux_14_11, A1=>nx11307, B0
      =>d_arr_mul_14_11, B1=>nx10459);
   lat_d_arr_14_12 : latch port map ( Q=>d_arr_14_12, D=>nx2968, CLK=>
      nx10227);
   ix2969 : ao22 port map ( Y=>nx2968, A0=>d_arr_mux_14_12, A1=>nx11307, B0
      =>d_arr_mul_14_12, B1=>nx10459);
   lat_d_arr_14_13 : latch port map ( Q=>d_arr_14_13, D=>nx2976, CLK=>
      nx10227);
   ix2977 : ao22 port map ( Y=>nx2976, A0=>d_arr_mux_14_13, A1=>nx11307, B0
      =>d_arr_mul_14_13, B1=>nx10459);
   lat_d_arr_14_14 : latch port map ( Q=>d_arr_14_14, D=>nx2984, CLK=>
      nx10227);
   ix2985 : ao22 port map ( Y=>nx2984, A0=>d_arr_mux_14_14, A1=>nx11307, B0
      =>d_arr_mul_14_14, B1=>nx10459);
   lat_d_arr_14_15 : latch port map ( Q=>d_arr_14_15, D=>nx2992, CLK=>
      nx10227);
   ix2993 : ao22 port map ( Y=>nx2992, A0=>d_arr_mux_14_15, A1=>nx11307, B0
      =>d_arr_mul_14_15, B1=>nx10459);
   lat_d_arr_14_16 : latch port map ( Q=>d_arr_14_16, D=>nx3000, CLK=>
      nx10229);
   ix3001 : ao22 port map ( Y=>nx3000, A0=>d_arr_mux_14_16, A1=>nx11307, B0
      =>d_arr_mul_14_16, B1=>nx10461);
   lat_d_arr_14_17 : latch port map ( Q=>d_arr_14_17, D=>nx3008, CLK=>
      nx10229);
   ix3009 : ao22 port map ( Y=>nx3008, A0=>d_arr_mux_14_17, A1=>nx11309, B0
      =>d_arr_mul_14_17, B1=>nx10461);
   lat_d_arr_14_18 : latch port map ( Q=>d_arr_14_18, D=>nx3016, CLK=>
      nx10229);
   ix3017 : ao22 port map ( Y=>nx3016, A0=>d_arr_mux_14_18, A1=>nx11309, B0
      =>d_arr_mul_14_18, B1=>nx10461);
   lat_d_arr_14_19 : latch port map ( Q=>d_arr_14_19, D=>nx3024, CLK=>
      nx10229);
   ix3025 : ao22 port map ( Y=>nx3024, A0=>d_arr_mux_14_19, A1=>nx11309, B0
      =>d_arr_mul_14_19, B1=>nx10461);
   lat_d_arr_14_20 : latch port map ( Q=>d_arr_14_20, D=>nx3032, CLK=>
      nx10229);
   ix3033 : ao22 port map ( Y=>nx3032, A0=>d_arr_mux_14_20, A1=>nx11309, B0
      =>d_arr_mul_14_20, B1=>nx10461);
   lat_d_arr_14_21 : latch port map ( Q=>d_arr_14_21, D=>nx3040, CLK=>
      nx10229);
   ix3041 : ao22 port map ( Y=>nx3040, A0=>d_arr_mux_14_21, A1=>nx11309, B0
      =>d_arr_mul_14_21, B1=>nx10461);
   lat_d_arr_14_22 : latch port map ( Q=>d_arr_14_22, D=>nx3048, CLK=>
      nx10229);
   ix3049 : ao22 port map ( Y=>nx3048, A0=>d_arr_mux_14_22, A1=>nx11309, B0
      =>d_arr_mul_14_22, B1=>nx10461);
   lat_d_arr_14_23 : latch port map ( Q=>d_arr_14_23, D=>nx3056, CLK=>
      nx10231);
   ix3057 : ao22 port map ( Y=>nx3056, A0=>d_arr_mux_14_23, A1=>nx11309, B0
      =>d_arr_mul_14_23, B1=>nx10463);
   lat_d_arr_14_24 : latch port map ( Q=>d_arr_14_24, D=>nx3064, CLK=>
      nx10231);
   ix3065 : ao22 port map ( Y=>nx3064, A0=>d_arr_mux_14_24, A1=>nx11311, B0
      =>d_arr_mul_14_24, B1=>nx10463);
   lat_d_arr_14_25 : latch port map ( Q=>d_arr_14_25, D=>nx3072, CLK=>
      nx10231);
   ix3073 : ao22 port map ( Y=>nx3072, A0=>d_arr_mux_14_25, A1=>nx11311, B0
      =>d_arr_mul_14_25, B1=>nx10463);
   lat_d_arr_14_26 : latch port map ( Q=>d_arr_14_26, D=>nx3080, CLK=>
      nx10231);
   ix3081 : ao22 port map ( Y=>nx3080, A0=>d_arr_mux_14_26, A1=>nx11311, B0
      =>d_arr_mul_14_26, B1=>nx10463);
   lat_d_arr_14_27 : latch port map ( Q=>d_arr_14_27, D=>nx3088, CLK=>
      nx10231);
   ix3089 : ao22 port map ( Y=>nx3088, A0=>d_arr_mux_14_27, A1=>nx11311, B0
      =>d_arr_mul_14_27, B1=>nx10463);
   lat_d_arr_14_28 : latch port map ( Q=>d_arr_14_28, D=>nx3096, CLK=>
      nx10231);
   ix3097 : ao22 port map ( Y=>nx3096, A0=>d_arr_mux_14_28, A1=>nx11311, B0
      =>d_arr_mul_14_28, B1=>nx10463);
   lat_d_arr_14_29 : latch port map ( Q=>d_arr_14_29, D=>nx3104, CLK=>
      nx10231);
   ix3105 : ao22 port map ( Y=>nx3104, A0=>d_arr_mux_14_29, A1=>nx11311, B0
      =>d_arr_mul_14_29, B1=>nx10463);
   lat_d_arr_14_30 : latch port map ( Q=>d_arr_14_30, D=>nx3112, CLK=>
      nx10233);
   ix3113 : ao22 port map ( Y=>nx3112, A0=>d_arr_mux_14_30, A1=>nx11311, B0
      =>d_arr_mul_14_30, B1=>nx10465);
   lat_d_arr_14_31 : latch port map ( Q=>d_arr_14_31, D=>nx3120, CLK=>
      nx10233);
   ix3121 : ao22 port map ( Y=>nx3120, A0=>d_arr_mux_14_31, A1=>nx11313, B0
      =>d_arr_mul_14_31, B1=>nx10465);
   lat_d_arr_13_0 : latch port map ( Q=>d_arr_13_0, D=>nx3132, CLK=>nx10233
   );
   ix3133 : inv01 port map ( Y=>nx3132, A=>nx8423);
   ix8424 : aoi222 port map ( Y=>nx8423, A0=>d_arr_mux_13_0, A1=>nx11313, B0
      =>d_arr_mul_13_0, B1=>nx10465, C0=>d_arr_add_13_0, C1=>nx10657);
   lat_d_arr_13_1 : latch port map ( Q=>d_arr_13_1, D=>nx3144, CLK=>nx10233
   );
   ix3145 : inv01 port map ( Y=>nx3144, A=>nx8429);
   ix8430 : aoi222 port map ( Y=>nx8429, A0=>d_arr_mux_13_1, A1=>nx11313, B0
      =>d_arr_mul_13_1, B1=>nx10465, C0=>d_arr_add_13_1, C1=>nx10657);
   lat_d_arr_13_2 : latch port map ( Q=>d_arr_13_2, D=>nx3156, CLK=>nx10233
   );
   ix3157 : inv01 port map ( Y=>nx3156, A=>nx8435);
   ix8436 : aoi222 port map ( Y=>nx8435, A0=>d_arr_mux_13_2, A1=>nx11313, B0
      =>d_arr_mul_13_2, B1=>nx10465, C0=>d_arr_add_13_2, C1=>nx10657);
   lat_d_arr_13_3 : latch port map ( Q=>d_arr_13_3, D=>nx3168, CLK=>nx10233
   );
   ix3169 : inv01 port map ( Y=>nx3168, A=>nx8441);
   ix8442 : aoi222 port map ( Y=>nx8441, A0=>d_arr_mux_13_3, A1=>nx11313, B0
      =>d_arr_mul_13_3, B1=>nx10465, C0=>d_arr_add_13_3, C1=>nx10657);
   lat_d_arr_13_4 : latch port map ( Q=>d_arr_13_4, D=>nx3180, CLK=>nx10233
   );
   ix3181 : inv01 port map ( Y=>nx3180, A=>nx8447);
   ix8448 : aoi222 port map ( Y=>nx8447, A0=>d_arr_mux_13_4, A1=>nx11313, B0
      =>d_arr_mul_13_4, B1=>nx10465, C0=>d_arr_add_13_4, C1=>nx10657);
   lat_d_arr_13_5 : latch port map ( Q=>d_arr_13_5, D=>nx3192, CLK=>nx10235
   );
   ix3193 : inv01 port map ( Y=>nx3192, A=>nx8453);
   ix8454 : aoi222 port map ( Y=>nx8453, A0=>d_arr_mux_13_5, A1=>nx11313, B0
      =>d_arr_mul_13_5, B1=>nx10467, C0=>d_arr_add_13_5, C1=>nx10659);
   lat_d_arr_13_6 : latch port map ( Q=>d_arr_13_6, D=>nx3204, CLK=>nx10235
   );
   ix3205 : inv01 port map ( Y=>nx3204, A=>nx8459);
   ix8460 : aoi222 port map ( Y=>nx8459, A0=>d_arr_mux_13_6, A1=>nx11315, B0
      =>d_arr_mul_13_6, B1=>nx10467, C0=>d_arr_add_13_6, C1=>nx10659);
   lat_d_arr_13_7 : latch port map ( Q=>d_arr_13_7, D=>nx3216, CLK=>nx10235
   );
   ix3217 : inv01 port map ( Y=>nx3216, A=>nx8465);
   ix8466 : aoi222 port map ( Y=>nx8465, A0=>d_arr_mux_13_7, A1=>nx11315, B0
      =>d_arr_mul_13_7, B1=>nx10467, C0=>d_arr_add_13_7, C1=>nx10659);
   lat_d_arr_13_8 : latch port map ( Q=>d_arr_13_8, D=>nx3228, CLK=>nx10235
   );
   ix3229 : inv01 port map ( Y=>nx3228, A=>nx8471);
   ix8472 : aoi222 port map ( Y=>nx8471, A0=>d_arr_mux_13_8, A1=>nx11315, B0
      =>d_arr_mul_13_8, B1=>nx10467, C0=>d_arr_add_13_8, C1=>nx10659);
   lat_d_arr_13_9 : latch port map ( Q=>d_arr_13_9, D=>nx3240, CLK=>nx10235
   );
   ix3241 : inv01 port map ( Y=>nx3240, A=>nx8477);
   ix8478 : aoi222 port map ( Y=>nx8477, A0=>d_arr_mux_13_9, A1=>nx11315, B0
      =>d_arr_mul_13_9, B1=>nx10467, C0=>d_arr_add_13_9, C1=>nx10659);
   lat_d_arr_13_10 : latch port map ( Q=>d_arr_13_10, D=>nx3252, CLK=>
      nx10235);
   ix3253 : inv01 port map ( Y=>nx3252, A=>nx8481);
   ix8482 : aoi222 port map ( Y=>nx8481, A0=>d_arr_mux_13_10, A1=>nx11315, 
      B0=>d_arr_mul_13_10, B1=>nx10467, C0=>d_arr_add_13_10, C1=>nx10659);
   lat_d_arr_13_11 : latch port map ( Q=>d_arr_13_11, D=>nx3264, CLK=>
      nx10235);
   ix3265 : inv01 port map ( Y=>nx3264, A=>nx8485);
   ix8486 : aoi222 port map ( Y=>nx8485, A0=>d_arr_mux_13_11, A1=>nx11315, 
      B0=>d_arr_mul_13_11, B1=>nx10467, C0=>d_arr_add_13_11, C1=>nx10659);
   lat_d_arr_13_12 : latch port map ( Q=>d_arr_13_12, D=>nx3276, CLK=>
      nx10237);
   ix3277 : inv01 port map ( Y=>nx3276, A=>nx8489);
   ix8490 : aoi222 port map ( Y=>nx8489, A0=>d_arr_mux_13_12, A1=>nx11315, 
      B0=>d_arr_mul_13_12, B1=>nx10469, C0=>d_arr_add_13_12, C1=>nx10661);
   lat_d_arr_13_13 : latch port map ( Q=>d_arr_13_13, D=>nx3288, CLK=>
      nx10237);
   ix3289 : inv01 port map ( Y=>nx3288, A=>nx8493);
   ix8494 : aoi222 port map ( Y=>nx8493, A0=>d_arr_mux_13_13, A1=>nx11317, 
      B0=>d_arr_mul_13_13, B1=>nx10469, C0=>d_arr_add_13_13, C1=>nx10661);
   lat_d_arr_13_14 : latch port map ( Q=>d_arr_13_14, D=>nx3300, CLK=>
      nx10237);
   ix3301 : inv01 port map ( Y=>nx3300, A=>nx8497);
   ix8498 : aoi222 port map ( Y=>nx8497, A0=>d_arr_mux_13_14, A1=>nx11317, 
      B0=>d_arr_mul_13_14, B1=>nx10469, C0=>d_arr_add_13_14, C1=>nx10661);
   lat_d_arr_13_15 : latch port map ( Q=>d_arr_13_15, D=>nx3312, CLK=>
      nx10237);
   ix3313 : inv01 port map ( Y=>nx3312, A=>nx8501);
   ix8502 : aoi222 port map ( Y=>nx8501, A0=>d_arr_mux_13_15, A1=>nx11317, 
      B0=>d_arr_mul_13_15, B1=>nx10469, C0=>d_arr_add_13_15, C1=>nx10661);
   lat_d_arr_13_16 : latch port map ( Q=>d_arr_13_16, D=>nx3324, CLK=>
      nx10237);
   ix3325 : inv01 port map ( Y=>nx3324, A=>nx8505);
   ix8506 : aoi222 port map ( Y=>nx8505, A0=>d_arr_mux_13_16, A1=>nx11317, 
      B0=>d_arr_mul_13_16, B1=>nx10469, C0=>d_arr_add_13_16, C1=>nx10661);
   lat_d_arr_13_17 : latch port map ( Q=>d_arr_13_17, D=>nx3336, CLK=>
      nx10237);
   ix3337 : inv01 port map ( Y=>nx3336, A=>nx8509);
   ix8510 : aoi222 port map ( Y=>nx8509, A0=>d_arr_mux_13_17, A1=>nx11317, 
      B0=>d_arr_mul_13_17, B1=>nx10469, C0=>d_arr_add_13_17, C1=>nx10661);
   lat_d_arr_13_18 : latch port map ( Q=>d_arr_13_18, D=>nx3348, CLK=>
      nx10237);
   ix3349 : inv01 port map ( Y=>nx3348, A=>nx8513);
   ix8514 : aoi222 port map ( Y=>nx8513, A0=>d_arr_mux_13_18, A1=>nx11317, 
      B0=>d_arr_mul_13_18, B1=>nx10469, C0=>d_arr_add_13_18, C1=>nx10661);
   lat_d_arr_13_19 : latch port map ( Q=>d_arr_13_19, D=>nx3360, CLK=>
      nx10239);
   ix3361 : inv01 port map ( Y=>nx3360, A=>nx8517);
   ix8518 : aoi222 port map ( Y=>nx8517, A0=>d_arr_mux_13_19, A1=>nx11317, 
      B0=>d_arr_mul_13_19, B1=>nx10471, C0=>d_arr_add_13_19, C1=>nx10663);
   lat_d_arr_13_20 : latch port map ( Q=>d_arr_13_20, D=>nx3372, CLK=>
      nx10239);
   ix3373 : inv01 port map ( Y=>nx3372, A=>nx8521);
   ix8522 : aoi222 port map ( Y=>nx8521, A0=>d_arr_mux_13_20, A1=>nx11319, 
      B0=>d_arr_mul_13_20, B1=>nx10471, C0=>d_arr_add_13_20, C1=>nx10663);
   lat_d_arr_13_21 : latch port map ( Q=>d_arr_13_21, D=>nx3384, CLK=>
      nx10239);
   ix3385 : inv01 port map ( Y=>nx3384, A=>nx8525);
   ix8526 : aoi222 port map ( Y=>nx8525, A0=>d_arr_mux_13_21, A1=>nx11319, 
      B0=>d_arr_mul_13_21, B1=>nx10471, C0=>d_arr_add_13_21, C1=>nx10663);
   lat_d_arr_13_22 : latch port map ( Q=>d_arr_13_22, D=>nx3396, CLK=>
      nx10239);
   ix3397 : inv01 port map ( Y=>nx3396, A=>nx8529);
   ix8530 : aoi222 port map ( Y=>nx8529, A0=>d_arr_mux_13_22, A1=>nx11319, 
      B0=>d_arr_mul_13_22, B1=>nx10471, C0=>d_arr_add_13_22, C1=>nx10663);
   lat_d_arr_13_23 : latch port map ( Q=>d_arr_13_23, D=>nx3408, CLK=>
      nx10239);
   ix3409 : inv01 port map ( Y=>nx3408, A=>nx8533);
   ix8534 : aoi222 port map ( Y=>nx8533, A0=>d_arr_mux_13_23, A1=>nx11319, 
      B0=>d_arr_mul_13_23, B1=>nx10471, C0=>d_arr_add_13_23, C1=>nx10663);
   lat_d_arr_13_24 : latch port map ( Q=>d_arr_13_24, D=>nx3420, CLK=>
      nx10239);
   ix3421 : inv01 port map ( Y=>nx3420, A=>nx8537);
   ix8538 : aoi222 port map ( Y=>nx8537, A0=>d_arr_mux_13_24, A1=>nx11319, 
      B0=>d_arr_mul_13_24, B1=>nx10471, C0=>d_arr_add_13_24, C1=>nx10663);
   lat_d_arr_13_25 : latch port map ( Q=>d_arr_13_25, D=>nx3432, CLK=>
      nx10239);
   ix3433 : inv01 port map ( Y=>nx3432, A=>nx8541);
   ix8542 : aoi222 port map ( Y=>nx8541, A0=>d_arr_mux_13_25, A1=>nx11319, 
      B0=>d_arr_mul_13_25, B1=>nx10471, C0=>d_arr_add_13_25, C1=>nx10663);
   lat_d_arr_13_26 : latch port map ( Q=>d_arr_13_26, D=>nx3444, CLK=>
      nx10241);
   ix3445 : inv01 port map ( Y=>nx3444, A=>nx8545);
   ix8546 : aoi222 port map ( Y=>nx8545, A0=>d_arr_mux_13_26, A1=>nx11319, 
      B0=>d_arr_mul_13_26, B1=>nx10473, C0=>d_arr_add_13_26, C1=>nx10665);
   lat_d_arr_13_27 : latch port map ( Q=>d_arr_13_27, D=>nx3456, CLK=>
      nx10241);
   ix3457 : inv01 port map ( Y=>nx3456, A=>nx8549);
   ix8550 : aoi222 port map ( Y=>nx8549, A0=>d_arr_mux_13_27, A1=>nx11321, 
      B0=>d_arr_mul_13_27, B1=>nx10473, C0=>d_arr_add_13_27, C1=>nx10665);
   lat_d_arr_13_28 : latch port map ( Q=>d_arr_13_28, D=>nx3468, CLK=>
      nx10241);
   ix3469 : inv01 port map ( Y=>nx3468, A=>nx8553);
   ix8554 : aoi222 port map ( Y=>nx8553, A0=>d_arr_mux_13_28, A1=>nx11321, 
      B0=>d_arr_mul_13_28, B1=>nx10473, C0=>d_arr_add_13_28, C1=>nx10665);
   lat_d_arr_13_29 : latch port map ( Q=>d_arr_13_29, D=>nx3480, CLK=>
      nx10241);
   ix3481 : inv01 port map ( Y=>nx3480, A=>nx8557);
   ix8558 : aoi222 port map ( Y=>nx8557, A0=>d_arr_mux_13_29, A1=>nx11321, 
      B0=>d_arr_mul_13_29, B1=>nx10473, C0=>d_arr_add_13_29, C1=>nx10665);
   lat_d_arr_13_30 : latch port map ( Q=>d_arr_13_30, D=>nx3492, CLK=>
      nx10241);
   ix3493 : inv01 port map ( Y=>nx3492, A=>nx8561);
   ix8562 : aoi222 port map ( Y=>nx8561, A0=>d_arr_mux_13_30, A1=>nx11321, 
      B0=>d_arr_mul_13_30, B1=>nx10473, C0=>d_arr_add_13_30, C1=>nx10665);
   lat_d_arr_13_31 : latch port map ( Q=>d_arr_13_31, D=>nx3504, CLK=>
      nx10241);
   ix3505 : inv01 port map ( Y=>nx3504, A=>nx8565);
   ix8566 : aoi222 port map ( Y=>nx8565, A0=>d_arr_mux_13_31, A1=>nx11321, 
      B0=>d_arr_mul_13_31, B1=>nx10473, C0=>d_arr_add_13_31, C1=>nx10665);
   lat_d_arr_12_0 : latch port map ( Q=>d_arr_12_0, D=>nx3516, CLK=>nx10241
   );
   ix3517 : inv01 port map ( Y=>nx3516, A=>nx8569);
   ix8570 : aoi222 port map ( Y=>nx8569, A0=>d_arr_mux_12_0, A1=>nx11321, B0
      =>d_arr_mul_12_0, B1=>nx10473, C0=>d_arr_add_12_0, C1=>nx10665);
   lat_d_arr_12_1 : latch port map ( Q=>d_arr_12_1, D=>nx3528, CLK=>nx10243
   );
   ix3529 : inv01 port map ( Y=>nx3528, A=>nx8573);
   ix8574 : aoi222 port map ( Y=>nx8573, A0=>d_arr_mux_12_1, A1=>nx11321, B0
      =>d_arr_mul_12_1, B1=>nx10475, C0=>d_arr_add_12_1, C1=>nx10667);
   lat_d_arr_12_2 : latch port map ( Q=>d_arr_12_2, D=>nx3540, CLK=>nx10243
   );
   ix3541 : inv01 port map ( Y=>nx3540, A=>nx8577);
   ix8578 : aoi222 port map ( Y=>nx8577, A0=>d_arr_mux_12_2, A1=>nx11323, B0
      =>d_arr_mul_12_2, B1=>nx10475, C0=>d_arr_add_12_2, C1=>nx10667);
   lat_d_arr_12_3 : latch port map ( Q=>d_arr_12_3, D=>nx3552, CLK=>nx10243
   );
   ix3553 : inv01 port map ( Y=>nx3552, A=>nx8581);
   ix8582 : aoi222 port map ( Y=>nx8581, A0=>d_arr_mux_12_3, A1=>nx11323, B0
      =>d_arr_mul_12_3, B1=>nx10475, C0=>d_arr_add_12_3, C1=>nx10667);
   lat_d_arr_12_4 : latch port map ( Q=>d_arr_12_4, D=>nx3564, CLK=>nx10243
   );
   ix3565 : inv01 port map ( Y=>nx3564, A=>nx8585);
   ix8586 : aoi222 port map ( Y=>nx8585, A0=>d_arr_mux_12_4, A1=>nx11323, B0
      =>d_arr_mul_12_4, B1=>nx10475, C0=>d_arr_add_12_4, C1=>nx10667);
   lat_d_arr_12_5 : latch port map ( Q=>d_arr_12_5, D=>nx3576, CLK=>nx10243
   );
   ix3577 : inv01 port map ( Y=>nx3576, A=>nx8589);
   ix8590 : aoi222 port map ( Y=>nx8589, A0=>d_arr_mux_12_5, A1=>nx11323, B0
      =>d_arr_mul_12_5, B1=>nx10475, C0=>d_arr_add_12_5, C1=>nx10667);
   lat_d_arr_12_6 : latch port map ( Q=>d_arr_12_6, D=>nx3588, CLK=>nx10243
   );
   ix3589 : inv01 port map ( Y=>nx3588, A=>nx8593);
   ix8594 : aoi222 port map ( Y=>nx8593, A0=>d_arr_mux_12_6, A1=>nx11323, B0
      =>d_arr_mul_12_6, B1=>nx10475, C0=>d_arr_add_12_6, C1=>nx10667);
   lat_d_arr_12_7 : latch port map ( Q=>d_arr_12_7, D=>nx3600, CLK=>nx10243
   );
   ix3601 : inv01 port map ( Y=>nx3600, A=>nx8597);
   ix8598 : aoi222 port map ( Y=>nx8597, A0=>d_arr_mux_12_7, A1=>nx11323, B0
      =>d_arr_mul_12_7, B1=>nx10475, C0=>d_arr_add_12_7, C1=>nx10667);
   lat_d_arr_12_8 : latch port map ( Q=>d_arr_12_8, D=>nx3612, CLK=>nx10245
   );
   ix3613 : inv01 port map ( Y=>nx3612, A=>nx8601);
   ix8602 : aoi222 port map ( Y=>nx8601, A0=>d_arr_mux_12_8, A1=>nx11323, B0
      =>d_arr_mul_12_8, B1=>nx10477, C0=>d_arr_add_12_8, C1=>nx10669);
   lat_d_arr_12_9 : latch port map ( Q=>d_arr_12_9, D=>nx3624, CLK=>nx10245
   );
   ix3625 : inv01 port map ( Y=>nx3624, A=>nx8605);
   ix8606 : aoi222 port map ( Y=>nx8605, A0=>d_arr_mux_12_9, A1=>nx11325, B0
      =>d_arr_mul_12_9, B1=>nx10477, C0=>d_arr_add_12_9, C1=>nx10669);
   lat_d_arr_12_10 : latch port map ( Q=>d_arr_12_10, D=>nx3636, CLK=>
      nx10245);
   ix3637 : inv01 port map ( Y=>nx3636, A=>nx8609);
   ix8610 : aoi222 port map ( Y=>nx8609, A0=>d_arr_mux_12_10, A1=>nx11325, 
      B0=>d_arr_mul_12_10, B1=>nx10477, C0=>d_arr_add_12_10, C1=>nx10669);
   lat_d_arr_12_11 : latch port map ( Q=>d_arr_12_11, D=>nx3648, CLK=>
      nx10245);
   ix3649 : inv01 port map ( Y=>nx3648, A=>nx8613);
   ix8614 : aoi222 port map ( Y=>nx8613, A0=>d_arr_mux_12_11, A1=>nx11325, 
      B0=>d_arr_mul_12_11, B1=>nx10477, C0=>d_arr_add_12_11, C1=>nx10669);
   lat_d_arr_12_12 : latch port map ( Q=>d_arr_12_12, D=>nx3660, CLK=>
      nx10245);
   ix3661 : inv01 port map ( Y=>nx3660, A=>nx8617);
   ix8618 : aoi222 port map ( Y=>nx8617, A0=>d_arr_mux_12_12, A1=>nx11325, 
      B0=>d_arr_mul_12_12, B1=>nx10477, C0=>d_arr_add_12_12, C1=>nx10669);
   lat_d_arr_12_13 : latch port map ( Q=>d_arr_12_13, D=>nx3672, CLK=>
      nx10245);
   ix3673 : inv01 port map ( Y=>nx3672, A=>nx8621);
   ix8622 : aoi222 port map ( Y=>nx8621, A0=>d_arr_mux_12_13, A1=>nx11325, 
      B0=>d_arr_mul_12_13, B1=>nx10477, C0=>d_arr_add_12_13, C1=>nx10669);
   lat_d_arr_12_14 : latch port map ( Q=>d_arr_12_14, D=>nx3684, CLK=>
      nx10245);
   ix3685 : inv01 port map ( Y=>nx3684, A=>nx8625);
   ix8626 : aoi222 port map ( Y=>nx8625, A0=>d_arr_mux_12_14, A1=>nx11325, 
      B0=>d_arr_mul_12_14, B1=>nx10477, C0=>d_arr_add_12_14, C1=>nx10669);
   lat_d_arr_12_15 : latch port map ( Q=>d_arr_12_15, D=>nx3696, CLK=>
      nx10247);
   ix3697 : inv01 port map ( Y=>nx3696, A=>nx8629);
   ix8630 : aoi222 port map ( Y=>nx8629, A0=>d_arr_mux_12_15, A1=>nx11325, 
      B0=>d_arr_mul_12_15, B1=>nx10479, C0=>d_arr_add_12_15, C1=>nx10671);
   lat_d_arr_12_16 : latch port map ( Q=>d_arr_12_16, D=>nx3708, CLK=>
      nx10247);
   ix3709 : inv01 port map ( Y=>nx3708, A=>nx8633);
   ix8634 : aoi222 port map ( Y=>nx8633, A0=>d_arr_mux_12_16, A1=>nx11327, 
      B0=>d_arr_mul_12_16, B1=>nx10479, C0=>d_arr_add_12_16, C1=>nx10671);
   lat_d_arr_12_17 : latch port map ( Q=>d_arr_12_17, D=>nx3720, CLK=>
      nx10247);
   ix3721 : inv01 port map ( Y=>nx3720, A=>nx8637);
   ix8638 : aoi222 port map ( Y=>nx8637, A0=>d_arr_mux_12_17, A1=>nx11327, 
      B0=>d_arr_mul_12_17, B1=>nx10479, C0=>d_arr_add_12_17, C1=>nx10671);
   lat_d_arr_12_18 : latch port map ( Q=>d_arr_12_18, D=>nx3732, CLK=>
      nx10247);
   ix3733 : inv01 port map ( Y=>nx3732, A=>nx8641);
   ix8642 : aoi222 port map ( Y=>nx8641, A0=>d_arr_mux_12_18, A1=>nx11327, 
      B0=>d_arr_mul_12_18, B1=>nx10479, C0=>d_arr_add_12_18, C1=>nx10671);
   lat_d_arr_12_19 : latch port map ( Q=>d_arr_12_19, D=>nx3744, CLK=>
      nx10247);
   ix3745 : inv01 port map ( Y=>nx3744, A=>nx8645);
   ix8646 : aoi222 port map ( Y=>nx8645, A0=>d_arr_mux_12_19, A1=>nx11327, 
      B0=>d_arr_mul_12_19, B1=>nx10479, C0=>d_arr_add_12_19, C1=>nx10671);
   lat_d_arr_12_20 : latch port map ( Q=>d_arr_12_20, D=>nx3756, CLK=>
      nx10247);
   ix3757 : inv01 port map ( Y=>nx3756, A=>nx8649);
   ix8650 : aoi222 port map ( Y=>nx8649, A0=>d_arr_mux_12_20, A1=>nx11327, 
      B0=>d_arr_mul_12_20, B1=>nx10479, C0=>d_arr_add_12_20, C1=>nx10671);
   lat_d_arr_12_21 : latch port map ( Q=>d_arr_12_21, D=>nx3768, CLK=>
      nx10247);
   ix3769 : inv01 port map ( Y=>nx3768, A=>nx8653);
   ix8654 : aoi222 port map ( Y=>nx8653, A0=>d_arr_mux_12_21, A1=>nx11327, 
      B0=>d_arr_mul_12_21, B1=>nx10479, C0=>d_arr_add_12_21, C1=>nx10671);
   lat_d_arr_12_22 : latch port map ( Q=>d_arr_12_22, D=>nx3780, CLK=>
      nx10249);
   ix3781 : inv01 port map ( Y=>nx3780, A=>nx8657);
   ix8658 : aoi222 port map ( Y=>nx8657, A0=>d_arr_mux_12_22, A1=>nx11327, 
      B0=>d_arr_mul_12_22, B1=>nx10481, C0=>d_arr_add_12_22, C1=>nx10673);
   lat_d_arr_12_23 : latch port map ( Q=>d_arr_12_23, D=>nx3792, CLK=>
      nx10249);
   ix3793 : inv01 port map ( Y=>nx3792, A=>nx8661);
   ix8662 : aoi222 port map ( Y=>nx8661, A0=>d_arr_mux_12_23, A1=>nx11329, 
      B0=>d_arr_mul_12_23, B1=>nx10481, C0=>d_arr_add_12_23, C1=>nx10673);
   lat_d_arr_12_24 : latch port map ( Q=>d_arr_12_24, D=>nx3804, CLK=>
      nx10249);
   ix3805 : inv01 port map ( Y=>nx3804, A=>nx8665);
   ix8666 : aoi222 port map ( Y=>nx8665, A0=>d_arr_mux_12_24, A1=>nx11329, 
      B0=>d_arr_mul_12_24, B1=>nx10481, C0=>d_arr_add_12_24, C1=>nx10673);
   lat_d_arr_12_25 : latch port map ( Q=>d_arr_12_25, D=>nx3816, CLK=>
      nx10249);
   ix3817 : inv01 port map ( Y=>nx3816, A=>nx8669);
   ix8670 : aoi222 port map ( Y=>nx8669, A0=>d_arr_mux_12_25, A1=>nx11329, 
      B0=>d_arr_mul_12_25, B1=>nx10481, C0=>d_arr_add_12_25, C1=>nx10673);
   lat_d_arr_12_26 : latch port map ( Q=>d_arr_12_26, D=>nx3828, CLK=>
      nx10249);
   ix3829 : inv01 port map ( Y=>nx3828, A=>nx8673);
   ix8674 : aoi222 port map ( Y=>nx8673, A0=>d_arr_mux_12_26, A1=>nx11329, 
      B0=>d_arr_mul_12_26, B1=>nx10481, C0=>d_arr_add_12_26, C1=>nx10673);
   lat_d_arr_12_27 : latch port map ( Q=>d_arr_12_27, D=>nx3840, CLK=>
      nx10249);
   ix3841 : inv01 port map ( Y=>nx3840, A=>nx8677);
   ix8678 : aoi222 port map ( Y=>nx8677, A0=>d_arr_mux_12_27, A1=>nx11329, 
      B0=>d_arr_mul_12_27, B1=>nx10481, C0=>d_arr_add_12_27, C1=>nx10673);
   lat_d_arr_12_28 : latch port map ( Q=>d_arr_12_28, D=>nx3852, CLK=>
      nx10249);
   ix3853 : inv01 port map ( Y=>nx3852, A=>nx8681);
   ix8682 : aoi222 port map ( Y=>nx8681, A0=>d_arr_mux_12_28, A1=>nx11329, 
      B0=>d_arr_mul_12_28, B1=>nx10481, C0=>d_arr_add_12_28, C1=>nx10673);
   lat_d_arr_12_29 : latch port map ( Q=>d_arr_12_29, D=>nx3864, CLK=>
      nx10251);
   ix3865 : inv01 port map ( Y=>nx3864, A=>nx8685);
   ix8686 : aoi222 port map ( Y=>nx8685, A0=>d_arr_mux_12_29, A1=>nx11329, 
      B0=>d_arr_mul_12_29, B1=>nx10483, C0=>d_arr_add_12_29, C1=>nx10675);
   lat_d_arr_12_30 : latch port map ( Q=>d_arr_12_30, D=>nx3876, CLK=>
      nx10251);
   ix3877 : inv01 port map ( Y=>nx3876, A=>nx8689);
   ix8690 : aoi222 port map ( Y=>nx8689, A0=>d_arr_mux_12_30, A1=>nx11331, 
      B0=>d_arr_mul_12_30, B1=>nx10483, C0=>d_arr_add_12_30, C1=>nx10675);
   lat_d_arr_12_31 : latch port map ( Q=>d_arr_12_31, D=>nx3888, CLK=>
      nx10251);
   ix3889 : inv01 port map ( Y=>nx3888, A=>nx8693);
   ix8694 : aoi222 port map ( Y=>nx8693, A0=>d_arr_mux_12_31, A1=>nx11331, 
      B0=>d_arr_mul_12_31, B1=>nx10483, C0=>d_arr_add_12_31, C1=>nx10675);
   lat_d_arr_11_0 : latch port map ( Q=>d_arr_11_0, D=>nx3900, CLK=>nx10251
   );
   ix3901 : inv01 port map ( Y=>nx3900, A=>nx8697);
   ix8698 : aoi222 port map ( Y=>nx8697, A0=>d_arr_mux_11_0, A1=>nx11331, B0
      =>d_arr_mul_11_0, B1=>nx10483, C0=>d_arr_add_11_0, C1=>nx10675);
   lat_d_arr_11_1 : latch port map ( Q=>d_arr_11_1, D=>nx3912, CLK=>nx10251
   );
   ix3913 : inv01 port map ( Y=>nx3912, A=>nx8701);
   ix8702 : aoi222 port map ( Y=>nx8701, A0=>d_arr_mux_11_1, A1=>nx11331, B0
      =>d_arr_mul_11_1, B1=>nx10483, C0=>d_arr_add_11_1, C1=>nx10675);
   lat_d_arr_11_2 : latch port map ( Q=>d_arr_11_2, D=>nx3924, CLK=>nx10251
   );
   ix3925 : inv01 port map ( Y=>nx3924, A=>nx8705);
   ix8706 : aoi222 port map ( Y=>nx8705, A0=>d_arr_mux_11_2, A1=>nx11331, B0
      =>d_arr_mul_11_2, B1=>nx10483, C0=>d_arr_add_11_2, C1=>nx10675);
   lat_d_arr_11_3 : latch port map ( Q=>d_arr_11_3, D=>nx3936, CLK=>nx10251
   );
   ix3937 : inv01 port map ( Y=>nx3936, A=>nx8709);
   ix8710 : aoi222 port map ( Y=>nx8709, A0=>d_arr_mux_11_3, A1=>nx11331, B0
      =>d_arr_mul_11_3, B1=>nx10483, C0=>d_arr_add_11_3, C1=>nx10675);
   lat_d_arr_11_4 : latch port map ( Q=>d_arr_11_4, D=>nx3948, CLK=>nx10253
   );
   ix3949 : inv01 port map ( Y=>nx3948, A=>nx8713);
   ix8714 : aoi222 port map ( Y=>nx8713, A0=>d_arr_mux_11_4, A1=>nx11331, B0
      =>d_arr_mul_11_4, B1=>nx10485, C0=>d_arr_add_11_4, C1=>nx10677);
   lat_d_arr_11_5 : latch port map ( Q=>d_arr_11_5, D=>nx3960, CLK=>nx10253
   );
   ix3961 : inv01 port map ( Y=>nx3960, A=>nx8717);
   ix8718 : aoi222 port map ( Y=>nx8717, A0=>d_arr_mux_11_5, A1=>nx11333, B0
      =>d_arr_mul_11_5, B1=>nx10485, C0=>d_arr_add_11_5, C1=>nx10677);
   lat_d_arr_11_6 : latch port map ( Q=>d_arr_11_6, D=>nx3972, CLK=>nx10253
   );
   ix3973 : inv01 port map ( Y=>nx3972, A=>nx8721);
   ix8722 : aoi222 port map ( Y=>nx8721, A0=>d_arr_mux_11_6, A1=>nx11333, B0
      =>d_arr_mul_11_6, B1=>nx10485, C0=>d_arr_add_11_6, C1=>nx10677);
   lat_d_arr_11_7 : latch port map ( Q=>d_arr_11_7, D=>nx3984, CLK=>nx10253
   );
   ix3985 : inv01 port map ( Y=>nx3984, A=>nx8725);
   ix8726 : aoi222 port map ( Y=>nx8725, A0=>d_arr_mux_11_7, A1=>nx11333, B0
      =>d_arr_mul_11_7, B1=>nx10485, C0=>d_arr_add_11_7, C1=>nx10677);
   lat_d_arr_11_8 : latch port map ( Q=>d_arr_11_8, D=>nx3996, CLK=>nx10253
   );
   ix3997 : inv01 port map ( Y=>nx3996, A=>nx8729);
   ix8730 : aoi222 port map ( Y=>nx8729, A0=>d_arr_mux_11_8, A1=>nx11333, B0
      =>d_arr_mul_11_8, B1=>nx10485, C0=>d_arr_add_11_8, C1=>nx10677);
   lat_d_arr_11_9 : latch port map ( Q=>d_arr_11_9, D=>nx4008, CLK=>nx10253
   );
   ix4009 : inv01 port map ( Y=>nx4008, A=>nx8733);
   ix8734 : aoi222 port map ( Y=>nx8733, A0=>d_arr_mux_11_9, A1=>nx11333, B0
      =>d_arr_mul_11_9, B1=>nx10485, C0=>d_arr_add_11_9, C1=>nx10677);
   lat_d_arr_11_10 : latch port map ( Q=>d_arr_11_10, D=>nx4020, CLK=>
      nx10253);
   ix4021 : inv01 port map ( Y=>nx4020, A=>nx8737);
   ix8738 : aoi222 port map ( Y=>nx8737, A0=>d_arr_mux_11_10, A1=>nx11333, 
      B0=>d_arr_mul_11_10, B1=>nx10485, C0=>d_arr_add_11_10, C1=>nx10677);
   lat_d_arr_11_11 : latch port map ( Q=>d_arr_11_11, D=>nx4032, CLK=>
      nx10255);
   ix4033 : inv01 port map ( Y=>nx4032, A=>nx8741);
   ix8742 : aoi222 port map ( Y=>nx8741, A0=>d_arr_mux_11_11, A1=>nx11333, 
      B0=>d_arr_mul_11_11, B1=>nx10487, C0=>d_arr_add_11_11, C1=>nx10679);
   lat_d_arr_11_12 : latch port map ( Q=>d_arr_11_12, D=>nx4044, CLK=>
      nx10255);
   ix4045 : inv01 port map ( Y=>nx4044, A=>nx8745);
   ix8746 : aoi222 port map ( Y=>nx8745, A0=>d_arr_mux_11_12, A1=>nx11335, 
      B0=>d_arr_mul_11_12, B1=>nx10487, C0=>d_arr_add_11_12, C1=>nx10679);
   lat_d_arr_11_13 : latch port map ( Q=>d_arr_11_13, D=>nx4056, CLK=>
      nx10255);
   ix4057 : inv01 port map ( Y=>nx4056, A=>nx8749);
   ix8750 : aoi222 port map ( Y=>nx8749, A0=>d_arr_mux_11_13, A1=>nx11335, 
      B0=>d_arr_mul_11_13, B1=>nx10487, C0=>d_arr_add_11_13, C1=>nx10679);
   lat_d_arr_11_14 : latch port map ( Q=>d_arr_11_14, D=>nx4068, CLK=>
      nx10255);
   ix4069 : inv01 port map ( Y=>nx4068, A=>nx8753);
   ix8754 : aoi222 port map ( Y=>nx8753, A0=>d_arr_mux_11_14, A1=>nx11335, 
      B0=>d_arr_mul_11_14, B1=>nx10487, C0=>d_arr_add_11_14, C1=>nx10679);
   lat_d_arr_11_15 : latch port map ( Q=>d_arr_11_15, D=>nx4080, CLK=>
      nx10255);
   ix4081 : inv01 port map ( Y=>nx4080, A=>nx8757);
   ix8758 : aoi222 port map ( Y=>nx8757, A0=>d_arr_mux_11_15, A1=>nx11335, 
      B0=>d_arr_mul_11_15, B1=>nx10487, C0=>d_arr_add_11_15, C1=>nx10679);
   lat_d_arr_11_16 : latch port map ( Q=>d_arr_11_16, D=>nx4092, CLK=>
      nx10255);
   ix4093 : inv01 port map ( Y=>nx4092, A=>nx8761);
   ix8762 : aoi222 port map ( Y=>nx8761, A0=>d_arr_mux_11_16, A1=>nx11335, 
      B0=>d_arr_mul_11_16, B1=>nx10487, C0=>d_arr_add_11_16, C1=>nx10679);
   lat_d_arr_11_17 : latch port map ( Q=>d_arr_11_17, D=>nx4104, CLK=>
      nx10255);
   ix4105 : inv01 port map ( Y=>nx4104, A=>nx8765);
   ix8766 : aoi222 port map ( Y=>nx8765, A0=>d_arr_mux_11_17, A1=>nx11335, 
      B0=>d_arr_mul_11_17, B1=>nx10487, C0=>d_arr_add_11_17, C1=>nx10679);
   lat_d_arr_11_18 : latch port map ( Q=>d_arr_11_18, D=>nx4116, CLK=>
      nx10257);
   ix4117 : inv01 port map ( Y=>nx4116, A=>nx8769);
   ix8770 : aoi222 port map ( Y=>nx8769, A0=>d_arr_mux_11_18, A1=>nx11335, 
      B0=>d_arr_mul_11_18, B1=>nx10489, C0=>d_arr_add_11_18, C1=>nx10681);
   lat_d_arr_11_19 : latch port map ( Q=>d_arr_11_19, D=>nx4128, CLK=>
      nx10257);
   ix4129 : inv01 port map ( Y=>nx4128, A=>nx8773);
   ix8774 : aoi222 port map ( Y=>nx8773, A0=>d_arr_mux_11_19, A1=>nx11337, 
      B0=>d_arr_mul_11_19, B1=>nx10489, C0=>d_arr_add_11_19, C1=>nx10681);
   lat_d_arr_11_20 : latch port map ( Q=>d_arr_11_20, D=>nx4140, CLK=>
      nx10257);
   ix4141 : inv01 port map ( Y=>nx4140, A=>nx8777);
   ix8778 : aoi222 port map ( Y=>nx8777, A0=>d_arr_mux_11_20, A1=>nx11337, 
      B0=>d_arr_mul_11_20, B1=>nx10489, C0=>d_arr_add_11_20, C1=>nx10681);
   lat_d_arr_11_21 : latch port map ( Q=>d_arr_11_21, D=>nx4152, CLK=>
      nx10257);
   ix4153 : inv01 port map ( Y=>nx4152, A=>nx8781);
   ix8782 : aoi222 port map ( Y=>nx8781, A0=>d_arr_mux_11_21, A1=>nx11337, 
      B0=>d_arr_mul_11_21, B1=>nx10489, C0=>d_arr_add_11_21, C1=>nx10681);
   lat_d_arr_11_22 : latch port map ( Q=>d_arr_11_22, D=>nx4164, CLK=>
      nx10257);
   ix4165 : inv01 port map ( Y=>nx4164, A=>nx8785);
   ix8786 : aoi222 port map ( Y=>nx8785, A0=>d_arr_mux_11_22, A1=>nx11337, 
      B0=>d_arr_mul_11_22, B1=>nx10489, C0=>d_arr_add_11_22, C1=>nx10681);
   lat_d_arr_11_23 : latch port map ( Q=>d_arr_11_23, D=>nx4176, CLK=>
      nx10257);
   ix4177 : inv01 port map ( Y=>nx4176, A=>nx8789);
   ix8790 : aoi222 port map ( Y=>nx8789, A0=>d_arr_mux_11_23, A1=>nx11337, 
      B0=>d_arr_mul_11_23, B1=>nx10489, C0=>d_arr_add_11_23, C1=>nx10681);
   lat_d_arr_11_24 : latch port map ( Q=>d_arr_11_24, D=>nx4188, CLK=>
      nx10257);
   ix4189 : inv01 port map ( Y=>nx4188, A=>nx8793);
   ix8794 : aoi222 port map ( Y=>nx8793, A0=>d_arr_mux_11_24, A1=>nx11337, 
      B0=>d_arr_mul_11_24, B1=>nx10489, C0=>d_arr_add_11_24, C1=>nx10681);
   lat_d_arr_11_25 : latch port map ( Q=>d_arr_11_25, D=>nx4200, CLK=>
      nx10259);
   ix4201 : inv01 port map ( Y=>nx4200, A=>nx8797);
   ix8798 : aoi222 port map ( Y=>nx8797, A0=>d_arr_mux_11_25, A1=>nx11337, 
      B0=>d_arr_mul_11_25, B1=>nx10491, C0=>d_arr_add_11_25, C1=>nx10683);
   lat_d_arr_11_26 : latch port map ( Q=>d_arr_11_26, D=>nx4212, CLK=>
      nx10259);
   ix4213 : inv01 port map ( Y=>nx4212, A=>nx8801);
   ix8802 : aoi222 port map ( Y=>nx8801, A0=>d_arr_mux_11_26, A1=>nx11339, 
      B0=>d_arr_mul_11_26, B1=>nx10491, C0=>d_arr_add_11_26, C1=>nx10683);
   lat_d_arr_11_27 : latch port map ( Q=>d_arr_11_27, D=>nx4224, CLK=>
      nx10259);
   ix4225 : inv01 port map ( Y=>nx4224, A=>nx8805);
   ix8806 : aoi222 port map ( Y=>nx8805, A0=>d_arr_mux_11_27, A1=>nx11339, 
      B0=>d_arr_mul_11_27, B1=>nx10491, C0=>d_arr_add_11_27, C1=>nx10683);
   lat_d_arr_11_28 : latch port map ( Q=>d_arr_11_28, D=>nx4236, CLK=>
      nx10259);
   ix4237 : inv01 port map ( Y=>nx4236, A=>nx8809);
   ix8810 : aoi222 port map ( Y=>nx8809, A0=>d_arr_mux_11_28, A1=>nx11339, 
      B0=>d_arr_mul_11_28, B1=>nx10491, C0=>d_arr_add_11_28, C1=>nx10683);
   lat_d_arr_11_29 : latch port map ( Q=>d_arr_11_29, D=>nx4248, CLK=>
      nx10259);
   ix4249 : inv01 port map ( Y=>nx4248, A=>nx8813);
   ix8814 : aoi222 port map ( Y=>nx8813, A0=>d_arr_mux_11_29, A1=>nx11339, 
      B0=>d_arr_mul_11_29, B1=>nx10491, C0=>d_arr_add_11_29, C1=>nx10683);
   lat_d_arr_11_30 : latch port map ( Q=>d_arr_11_30, D=>nx4260, CLK=>
      nx10259);
   ix4261 : inv01 port map ( Y=>nx4260, A=>nx8817);
   ix8818 : aoi222 port map ( Y=>nx8817, A0=>d_arr_mux_11_30, A1=>nx11339, 
      B0=>d_arr_mul_11_30, B1=>nx10491, C0=>d_arr_add_11_30, C1=>nx10683);
   lat_d_arr_11_31 : latch port map ( Q=>d_arr_11_31, D=>nx4272, CLK=>
      nx10259);
   ix4273 : inv01 port map ( Y=>nx4272, A=>nx8821);
   ix8822 : aoi222 port map ( Y=>nx8821, A0=>d_arr_mux_11_31, A1=>nx11339, 
      B0=>d_arr_mul_11_31, B1=>nx10491, C0=>d_arr_add_11_31, C1=>nx10683);
   lat_d_arr_10_0 : latch port map ( Q=>d_arr_10_0, D=>nx4284, CLK=>nx10261
   );
   ix4285 : inv01 port map ( Y=>nx4284, A=>nx8825);
   ix8826 : aoi222 port map ( Y=>nx8825, A0=>d_arr_mux_10_0, A1=>nx11339, B0
      =>d_arr_mul_10_0, B1=>nx10493, C0=>d_arr_add_10_0, C1=>nx10685);
   lat_d_arr_10_1 : latch port map ( Q=>d_arr_10_1, D=>nx4296, CLK=>nx10261
   );
   ix4297 : inv01 port map ( Y=>nx4296, A=>nx8829);
   ix8830 : aoi222 port map ( Y=>nx8829, A0=>d_arr_mux_10_1, A1=>nx11341, B0
      =>d_arr_mul_10_1, B1=>nx10493, C0=>d_arr_add_10_1, C1=>nx10685);
   lat_d_arr_10_2 : latch port map ( Q=>d_arr_10_2, D=>nx4308, CLK=>nx10261
   );
   ix4309 : inv01 port map ( Y=>nx4308, A=>nx8833);
   ix8834 : aoi222 port map ( Y=>nx8833, A0=>d_arr_mux_10_2, A1=>nx11341, B0
      =>d_arr_mul_10_2, B1=>nx10493, C0=>d_arr_add_10_2, C1=>nx10685);
   lat_d_arr_10_3 : latch port map ( Q=>d_arr_10_3, D=>nx4320, CLK=>nx10261
   );
   ix4321 : inv01 port map ( Y=>nx4320, A=>nx8837);
   ix8838 : aoi222 port map ( Y=>nx8837, A0=>d_arr_mux_10_3, A1=>nx11341, B0
      =>d_arr_mul_10_3, B1=>nx10493, C0=>d_arr_add_10_3, C1=>nx10685);
   lat_d_arr_10_4 : latch port map ( Q=>d_arr_10_4, D=>nx4332, CLK=>nx10261
   );
   ix4333 : inv01 port map ( Y=>nx4332, A=>nx8841);
   ix8842 : aoi222 port map ( Y=>nx8841, A0=>d_arr_mux_10_4, A1=>nx11341, B0
      =>d_arr_mul_10_4, B1=>nx10493, C0=>d_arr_add_10_4, C1=>nx10685);
   lat_d_arr_10_5 : latch port map ( Q=>d_arr_10_5, D=>nx4344, CLK=>nx10261
   );
   ix4345 : inv01 port map ( Y=>nx4344, A=>nx8845);
   ix8846 : aoi222 port map ( Y=>nx8845, A0=>d_arr_mux_10_5, A1=>nx11341, B0
      =>d_arr_mul_10_5, B1=>nx10493, C0=>d_arr_add_10_5, C1=>nx10685);
   lat_d_arr_10_6 : latch port map ( Q=>d_arr_10_6, D=>nx4356, CLK=>nx10261
   );
   ix4357 : inv01 port map ( Y=>nx4356, A=>nx8849);
   ix8850 : aoi222 port map ( Y=>nx8849, A0=>d_arr_mux_10_6, A1=>nx11341, B0
      =>d_arr_mul_10_6, B1=>nx10493, C0=>d_arr_add_10_6, C1=>nx10685);
   lat_d_arr_10_7 : latch port map ( Q=>d_arr_10_7, D=>nx4368, CLK=>nx10263
   );
   ix4369 : inv01 port map ( Y=>nx4368, A=>nx8853);
   ix8854 : aoi222 port map ( Y=>nx8853, A0=>d_arr_mux_10_7, A1=>nx11341, B0
      =>d_arr_mul_10_7, B1=>nx10495, C0=>d_arr_add_10_7, C1=>nx10687);
   lat_d_arr_10_8 : latch port map ( Q=>d_arr_10_8, D=>nx4380, CLK=>nx10263
   );
   ix4381 : inv01 port map ( Y=>nx4380, A=>nx8857);
   ix8858 : aoi222 port map ( Y=>nx8857, A0=>d_arr_mux_10_8, A1=>nx11343, B0
      =>d_arr_mul_10_8, B1=>nx10495, C0=>d_arr_add_10_8, C1=>nx10687);
   lat_d_arr_10_9 : latch port map ( Q=>d_arr_10_9, D=>nx4392, CLK=>nx10263
   );
   ix4393 : inv01 port map ( Y=>nx4392, A=>nx8861);
   ix8862 : aoi222 port map ( Y=>nx8861, A0=>d_arr_mux_10_9, A1=>nx11343, B0
      =>d_arr_mul_10_9, B1=>nx10495, C0=>d_arr_add_10_9, C1=>nx10687);
   lat_d_arr_10_10 : latch port map ( Q=>d_arr_10_10, D=>nx4404, CLK=>
      nx10263);
   ix4405 : inv01 port map ( Y=>nx4404, A=>nx8865);
   ix8866 : aoi222 port map ( Y=>nx8865, A0=>d_arr_mux_10_10, A1=>nx11343, 
      B0=>d_arr_mul_10_10, B1=>nx10495, C0=>d_arr_add_10_10, C1=>nx10687);
   lat_d_arr_10_11 : latch port map ( Q=>d_arr_10_11, D=>nx4416, CLK=>
      nx10263);
   ix4417 : inv01 port map ( Y=>nx4416, A=>nx8869);
   ix8870 : aoi222 port map ( Y=>nx8869, A0=>d_arr_mux_10_11, A1=>nx11343, 
      B0=>d_arr_mul_10_11, B1=>nx10495, C0=>d_arr_add_10_11, C1=>nx10687);
   lat_d_arr_10_12 : latch port map ( Q=>d_arr_10_12, D=>nx4428, CLK=>
      nx10263);
   ix4429 : inv01 port map ( Y=>nx4428, A=>nx8873);
   ix8874 : aoi222 port map ( Y=>nx8873, A0=>d_arr_mux_10_12, A1=>nx11343, 
      B0=>d_arr_mul_10_12, B1=>nx10495, C0=>d_arr_add_10_12, C1=>nx10687);
   lat_d_arr_10_13 : latch port map ( Q=>d_arr_10_13, D=>nx4440, CLK=>
      nx10263);
   ix4441 : inv01 port map ( Y=>nx4440, A=>nx8877);
   ix8878 : aoi222 port map ( Y=>nx8877, A0=>d_arr_mux_10_13, A1=>nx11343, 
      B0=>d_arr_mul_10_13, B1=>nx10495, C0=>d_arr_add_10_13, C1=>nx10687);
   lat_d_arr_10_14 : latch port map ( Q=>d_arr_10_14, D=>nx4452, CLK=>
      nx10265);
   ix4453 : inv01 port map ( Y=>nx4452, A=>nx8881);
   ix8882 : aoi222 port map ( Y=>nx8881, A0=>d_arr_mux_10_14, A1=>nx11343, 
      B0=>d_arr_mul_10_14, B1=>nx10497, C0=>d_arr_add_10_14, C1=>nx10689);
   lat_d_arr_10_15 : latch port map ( Q=>d_arr_10_15, D=>nx4464, CLK=>
      nx10265);
   ix4465 : inv01 port map ( Y=>nx4464, A=>nx8885);
   ix8886 : aoi222 port map ( Y=>nx8885, A0=>d_arr_mux_10_15, A1=>nx11345, 
      B0=>d_arr_mul_10_15, B1=>nx10497, C0=>d_arr_add_10_15, C1=>nx10689);
   lat_d_arr_10_16 : latch port map ( Q=>d_arr_10_16, D=>nx4476, CLK=>
      nx10265);
   ix4477 : inv01 port map ( Y=>nx4476, A=>nx8889);
   ix8890 : aoi222 port map ( Y=>nx8889, A0=>d_arr_mux_10_16, A1=>nx11345, 
      B0=>d_arr_mul_10_16, B1=>nx10497, C0=>d_arr_add_10_16, C1=>nx10689);
   lat_d_arr_10_17 : latch port map ( Q=>d_arr_10_17, D=>nx4488, CLK=>
      nx10265);
   ix4489 : inv01 port map ( Y=>nx4488, A=>nx8893);
   ix8894 : aoi222 port map ( Y=>nx8893, A0=>d_arr_mux_10_17, A1=>nx11345, 
      B0=>d_arr_mul_10_17, B1=>nx10497, C0=>d_arr_add_10_17, C1=>nx10689);
   lat_d_arr_10_18 : latch port map ( Q=>d_arr_10_18, D=>nx4500, CLK=>
      nx10265);
   ix4501 : inv01 port map ( Y=>nx4500, A=>nx8897);
   ix8898 : aoi222 port map ( Y=>nx8897, A0=>d_arr_mux_10_18, A1=>nx11345, 
      B0=>d_arr_mul_10_18, B1=>nx10497, C0=>d_arr_add_10_18, C1=>nx10689);
   lat_d_arr_10_19 : latch port map ( Q=>d_arr_10_19, D=>nx4512, CLK=>
      nx10265);
   ix4513 : inv01 port map ( Y=>nx4512, A=>nx8901);
   ix8902 : aoi222 port map ( Y=>nx8901, A0=>d_arr_mux_10_19, A1=>nx11345, 
      B0=>d_arr_mul_10_19, B1=>nx10497, C0=>d_arr_add_10_19, C1=>nx10689);
   lat_d_arr_10_20 : latch port map ( Q=>d_arr_10_20, D=>nx4524, CLK=>
      nx10265);
   ix4525 : inv01 port map ( Y=>nx4524, A=>nx8905);
   ix8906 : aoi222 port map ( Y=>nx8905, A0=>d_arr_mux_10_20, A1=>nx11345, 
      B0=>d_arr_mul_10_20, B1=>nx10497, C0=>d_arr_add_10_20, C1=>nx10689);
   lat_d_arr_10_21 : latch port map ( Q=>d_arr_10_21, D=>nx4536, CLK=>
      nx10267);
   ix4537 : inv01 port map ( Y=>nx4536, A=>nx8909);
   ix8910 : aoi222 port map ( Y=>nx8909, A0=>d_arr_mux_10_21, A1=>nx11345, 
      B0=>d_arr_mul_10_21, B1=>nx10499, C0=>d_arr_add_10_21, C1=>nx10691);
   lat_d_arr_10_22 : latch port map ( Q=>d_arr_10_22, D=>nx4548, CLK=>
      nx10267);
   ix4549 : inv01 port map ( Y=>nx4548, A=>nx8913);
   ix8914 : aoi222 port map ( Y=>nx8913, A0=>d_arr_mux_10_22, A1=>nx11347, 
      B0=>d_arr_mul_10_22, B1=>nx10499, C0=>d_arr_add_10_22, C1=>nx10691);
   lat_d_arr_10_23 : latch port map ( Q=>d_arr_10_23, D=>nx4560, CLK=>
      nx10267);
   ix4561 : inv01 port map ( Y=>nx4560, A=>nx8917);
   ix8918 : aoi222 port map ( Y=>nx8917, A0=>d_arr_mux_10_23, A1=>nx11347, 
      B0=>d_arr_mul_10_23, B1=>nx10499, C0=>d_arr_add_10_23, C1=>nx10691);
   lat_d_arr_10_24 : latch port map ( Q=>d_arr_10_24, D=>nx4572, CLK=>
      nx10267);
   ix4573 : inv01 port map ( Y=>nx4572, A=>nx8921);
   ix8922 : aoi222 port map ( Y=>nx8921, A0=>d_arr_mux_10_24, A1=>nx11347, 
      B0=>d_arr_mul_10_24, B1=>nx10499, C0=>d_arr_add_10_24, C1=>nx10691);
   lat_d_arr_10_25 : latch port map ( Q=>d_arr_10_25, D=>nx4584, CLK=>
      nx10267);
   ix4585 : inv01 port map ( Y=>nx4584, A=>nx8925);
   ix8926 : aoi222 port map ( Y=>nx8925, A0=>d_arr_mux_10_25, A1=>nx11347, 
      B0=>d_arr_mul_10_25, B1=>nx10499, C0=>d_arr_add_10_25, C1=>nx10691);
   lat_d_arr_10_26 : latch port map ( Q=>d_arr_10_26, D=>nx4596, CLK=>
      nx10267);
   ix4597 : inv01 port map ( Y=>nx4596, A=>nx8929);
   ix8930 : aoi222 port map ( Y=>nx8929, A0=>d_arr_mux_10_26, A1=>nx11347, 
      B0=>d_arr_mul_10_26, B1=>nx10499, C0=>d_arr_add_10_26, C1=>nx10691);
   lat_d_arr_10_27 : latch port map ( Q=>d_arr_10_27, D=>nx4608, CLK=>
      nx10267);
   ix4609 : inv01 port map ( Y=>nx4608, A=>nx8933);
   ix8934 : aoi222 port map ( Y=>nx8933, A0=>d_arr_mux_10_27, A1=>nx11347, 
      B0=>d_arr_mul_10_27, B1=>nx10499, C0=>d_arr_add_10_27, C1=>nx10691);
   lat_d_arr_10_28 : latch port map ( Q=>d_arr_10_28, D=>nx4620, CLK=>
      nx10269);
   ix4621 : inv01 port map ( Y=>nx4620, A=>nx8937);
   ix8938 : aoi222 port map ( Y=>nx8937, A0=>d_arr_mux_10_28, A1=>nx11347, 
      B0=>d_arr_mul_10_28, B1=>nx10501, C0=>d_arr_add_10_28, C1=>nx10693);
   lat_d_arr_10_29 : latch port map ( Q=>d_arr_10_29, D=>nx4632, CLK=>
      nx10269);
   ix4633 : inv01 port map ( Y=>nx4632, A=>nx8941);
   ix8942 : aoi222 port map ( Y=>nx8941, A0=>d_arr_mux_10_29, A1=>nx11349, 
      B0=>d_arr_mul_10_29, B1=>nx10501, C0=>d_arr_add_10_29, C1=>nx10693);
   lat_d_arr_10_30 : latch port map ( Q=>d_arr_10_30, D=>nx4644, CLK=>
      nx10269);
   ix4645 : inv01 port map ( Y=>nx4644, A=>nx8945);
   ix8946 : aoi222 port map ( Y=>nx8945, A0=>d_arr_mux_10_30, A1=>nx11349, 
      B0=>d_arr_mul_10_30, B1=>nx10501, C0=>d_arr_add_10_30, C1=>nx10693);
   lat_d_arr_10_31 : latch port map ( Q=>d_arr_10_31, D=>nx4656, CLK=>
      nx10269);
   ix4657 : inv01 port map ( Y=>nx4656, A=>nx8949);
   ix8950 : aoi222 port map ( Y=>nx8949, A0=>d_arr_mux_10_31, A1=>nx11349, 
      B0=>d_arr_mul_10_31, B1=>nx10501, C0=>d_arr_add_10_31, C1=>nx10693);
   lat_d_arr_9_0 : latch port map ( Q=>d_arr_9_0, D=>nx4668, CLK=>nx10269);
   ix4669 : inv01 port map ( Y=>nx4668, A=>nx8953);
   ix8954 : aoi222 port map ( Y=>nx8953, A0=>d_arr_mux_9_0, A1=>nx11349, B0
      =>d_arr_mul_9_0, B1=>nx10501, C0=>d_arr_add_9_0, C1=>nx10693);
   lat_d_arr_9_1 : latch port map ( Q=>d_arr_9_1, D=>nx4680, CLK=>nx10269);
   ix4681 : inv01 port map ( Y=>nx4680, A=>nx8957);
   ix8958 : aoi222 port map ( Y=>nx8957, A0=>d_arr_mux_9_1, A1=>nx11349, B0
      =>d_arr_mul_9_1, B1=>nx10501, C0=>d_arr_add_9_1, C1=>nx10693);
   lat_d_arr_9_2 : latch port map ( Q=>d_arr_9_2, D=>nx4692, CLK=>nx10269);
   ix4693 : inv01 port map ( Y=>nx4692, A=>nx8961);
   ix8962 : aoi222 port map ( Y=>nx8961, A0=>d_arr_mux_9_2, A1=>nx11349, B0
      =>d_arr_mul_9_2, B1=>nx10501, C0=>d_arr_add_9_2, C1=>nx10693);
   lat_d_arr_9_3 : latch port map ( Q=>d_arr_9_3, D=>nx4704, CLK=>nx10271);
   ix4705 : inv01 port map ( Y=>nx4704, A=>nx8965);
   ix8966 : aoi222 port map ( Y=>nx8965, A0=>d_arr_mux_9_3, A1=>nx11349, B0
      =>d_arr_mul_9_3, B1=>nx10503, C0=>d_arr_add_9_3, C1=>nx10695);
   lat_d_arr_9_4 : latch port map ( Q=>d_arr_9_4, D=>nx4716, CLK=>nx10271);
   ix4717 : inv01 port map ( Y=>nx4716, A=>nx8969);
   ix8970 : aoi222 port map ( Y=>nx8969, A0=>d_arr_mux_9_4, A1=>nx11351, B0
      =>d_arr_mul_9_4, B1=>nx10503, C0=>d_arr_add_9_4, C1=>nx10695);
   lat_d_arr_9_5 : latch port map ( Q=>d_arr_9_5, D=>nx4728, CLK=>nx10271);
   ix4729 : inv01 port map ( Y=>nx4728, A=>nx8973);
   ix8974 : aoi222 port map ( Y=>nx8973, A0=>d_arr_mux_9_5, A1=>nx11351, B0
      =>d_arr_mul_9_5, B1=>nx10503, C0=>d_arr_add_9_5, C1=>nx10695);
   lat_d_arr_9_6 : latch port map ( Q=>d_arr_9_6, D=>nx4740, CLK=>nx10271);
   ix4741 : inv01 port map ( Y=>nx4740, A=>nx8977);
   ix8978 : aoi222 port map ( Y=>nx8977, A0=>d_arr_mux_9_6, A1=>nx11351, B0
      =>d_arr_mul_9_6, B1=>nx10503, C0=>d_arr_add_9_6, C1=>nx10695);
   lat_d_arr_9_7 : latch port map ( Q=>d_arr_9_7, D=>nx4752, CLK=>nx10271);
   ix4753 : inv01 port map ( Y=>nx4752, A=>nx8981);
   ix8982 : aoi222 port map ( Y=>nx8981, A0=>d_arr_mux_9_7, A1=>nx11351, B0
      =>d_arr_mul_9_7, B1=>nx10503, C0=>d_arr_add_9_7, C1=>nx10695);
   lat_d_arr_9_8 : latch port map ( Q=>d_arr_9_8, D=>nx4764, CLK=>nx10271);
   ix4765 : inv01 port map ( Y=>nx4764, A=>nx8985);
   ix8986 : aoi222 port map ( Y=>nx8985, A0=>d_arr_mux_9_8, A1=>nx11351, B0
      =>d_arr_mul_9_8, B1=>nx10503, C0=>d_arr_add_9_8, C1=>nx10695);
   lat_d_arr_9_9 : latch port map ( Q=>d_arr_9_9, D=>nx4776, CLK=>nx10271);
   ix4777 : inv01 port map ( Y=>nx4776, A=>nx8989);
   ix8990 : aoi222 port map ( Y=>nx8989, A0=>d_arr_mux_9_9, A1=>nx11351, B0
      =>d_arr_mul_9_9, B1=>nx10503, C0=>d_arr_add_9_9, C1=>nx10695);
   lat_d_arr_9_10 : latch port map ( Q=>d_arr_9_10, D=>nx4788, CLK=>nx10273
   );
   ix4789 : inv01 port map ( Y=>nx4788, A=>nx8993);
   ix8994 : aoi222 port map ( Y=>nx8993, A0=>d_arr_mux_9_10, A1=>nx11351, B0
      =>d_arr_mul_9_10, B1=>nx10505, C0=>d_arr_add_9_10, C1=>nx10697);
   lat_d_arr_9_11 : latch port map ( Q=>d_arr_9_11, D=>nx4800, CLK=>nx10273
   );
   ix4801 : inv01 port map ( Y=>nx4800, A=>nx8997);
   ix8998 : aoi222 port map ( Y=>nx8997, A0=>d_arr_mux_9_11, A1=>nx11353, B0
      =>d_arr_mul_9_11, B1=>nx10505, C0=>d_arr_add_9_11, C1=>nx10697);
   lat_d_arr_9_12 : latch port map ( Q=>d_arr_9_12, D=>nx4812, CLK=>nx10273
   );
   ix4813 : inv01 port map ( Y=>nx4812, A=>nx9001);
   ix9002 : aoi222 port map ( Y=>nx9001, A0=>d_arr_mux_9_12, A1=>nx11353, B0
      =>d_arr_mul_9_12, B1=>nx10505, C0=>d_arr_add_9_12, C1=>nx10697);
   lat_d_arr_9_13 : latch port map ( Q=>d_arr_9_13, D=>nx4824, CLK=>nx10273
   );
   ix4825 : inv01 port map ( Y=>nx4824, A=>nx9005);
   ix9006 : aoi222 port map ( Y=>nx9005, A0=>d_arr_mux_9_13, A1=>nx11353, B0
      =>d_arr_mul_9_13, B1=>nx10505, C0=>d_arr_add_9_13, C1=>nx10697);
   lat_d_arr_9_14 : latch port map ( Q=>d_arr_9_14, D=>nx4836, CLK=>nx10273
   );
   ix4837 : inv01 port map ( Y=>nx4836, A=>nx9009);
   ix9010 : aoi222 port map ( Y=>nx9009, A0=>d_arr_mux_9_14, A1=>nx11353, B0
      =>d_arr_mul_9_14, B1=>nx10505, C0=>d_arr_add_9_14, C1=>nx10697);
   lat_d_arr_9_15 : latch port map ( Q=>d_arr_9_15, D=>nx4848, CLK=>nx10273
   );
   ix4849 : inv01 port map ( Y=>nx4848, A=>nx9013);
   ix9014 : aoi222 port map ( Y=>nx9013, A0=>d_arr_mux_9_15, A1=>nx11353, B0
      =>d_arr_mul_9_15, B1=>nx10505, C0=>d_arr_add_9_15, C1=>nx10697);
   lat_d_arr_9_16 : latch port map ( Q=>d_arr_9_16, D=>nx4860, CLK=>nx10273
   );
   ix4861 : inv01 port map ( Y=>nx4860, A=>nx9017);
   ix9018 : aoi222 port map ( Y=>nx9017, A0=>d_arr_mux_9_16, A1=>nx11353, B0
      =>d_arr_mul_9_16, B1=>nx10505, C0=>d_arr_add_9_16, C1=>nx10697);
   lat_d_arr_9_17 : latch port map ( Q=>d_arr_9_17, D=>nx4872, CLK=>nx10275
   );
   ix4873 : inv01 port map ( Y=>nx4872, A=>nx9021);
   ix9022 : aoi222 port map ( Y=>nx9021, A0=>d_arr_mux_9_17, A1=>nx11353, B0
      =>d_arr_mul_9_17, B1=>nx10507, C0=>d_arr_add_9_17, C1=>nx10699);
   lat_d_arr_9_18 : latch port map ( Q=>d_arr_9_18, D=>nx4884, CLK=>nx10275
   );
   ix4885 : inv01 port map ( Y=>nx4884, A=>nx9025);
   ix9026 : aoi222 port map ( Y=>nx9025, A0=>d_arr_mux_9_18, A1=>nx11355, B0
      =>d_arr_mul_9_18, B1=>nx10507, C0=>d_arr_add_9_18, C1=>nx10699);
   lat_d_arr_9_19 : latch port map ( Q=>d_arr_9_19, D=>nx4896, CLK=>nx10275
   );
   ix4897 : inv01 port map ( Y=>nx4896, A=>nx9029);
   ix9030 : aoi222 port map ( Y=>nx9029, A0=>d_arr_mux_9_19, A1=>nx11355, B0
      =>d_arr_mul_9_19, B1=>nx10507, C0=>d_arr_add_9_19, C1=>nx10699);
   lat_d_arr_9_20 : latch port map ( Q=>d_arr_9_20, D=>nx4908, CLK=>nx10275
   );
   ix4909 : inv01 port map ( Y=>nx4908, A=>nx9033);
   ix9034 : aoi222 port map ( Y=>nx9033, A0=>d_arr_mux_9_20, A1=>nx11355, B0
      =>d_arr_mul_9_20, B1=>nx10507, C0=>d_arr_add_9_20, C1=>nx10699);
   lat_d_arr_9_21 : latch port map ( Q=>d_arr_9_21, D=>nx4920, CLK=>nx10275
   );
   ix4921 : inv01 port map ( Y=>nx4920, A=>nx9037);
   ix9038 : aoi222 port map ( Y=>nx9037, A0=>d_arr_mux_9_21, A1=>nx11355, B0
      =>d_arr_mul_9_21, B1=>nx10507, C0=>d_arr_add_9_21, C1=>nx10699);
   lat_d_arr_9_22 : latch port map ( Q=>d_arr_9_22, D=>nx4932, CLK=>nx10275
   );
   ix4933 : inv01 port map ( Y=>nx4932, A=>nx9041);
   ix9042 : aoi222 port map ( Y=>nx9041, A0=>d_arr_mux_9_22, A1=>nx11355, B0
      =>d_arr_mul_9_22, B1=>nx10507, C0=>d_arr_add_9_22, C1=>nx10699);
   lat_d_arr_9_23 : latch port map ( Q=>d_arr_9_23, D=>nx4944, CLK=>nx10275
   );
   ix4945 : inv01 port map ( Y=>nx4944, A=>nx9045);
   ix9046 : aoi222 port map ( Y=>nx9045, A0=>d_arr_mux_9_23, A1=>nx11355, B0
      =>d_arr_mul_9_23, B1=>nx10507, C0=>d_arr_add_9_23, C1=>nx10699);
   lat_d_arr_9_24 : latch port map ( Q=>d_arr_9_24, D=>nx4956, CLK=>nx10277
   );
   ix4957 : inv01 port map ( Y=>nx4956, A=>nx9049);
   ix9050 : aoi222 port map ( Y=>nx9049, A0=>d_arr_mux_9_24, A1=>nx11355, B0
      =>d_arr_mul_9_24, B1=>nx10509, C0=>d_arr_add_9_24, C1=>nx10701);
   lat_d_arr_9_25 : latch port map ( Q=>d_arr_9_25, D=>nx4968, CLK=>nx10277
   );
   ix4969 : inv01 port map ( Y=>nx4968, A=>nx9053);
   ix9054 : aoi222 port map ( Y=>nx9053, A0=>d_arr_mux_9_25, A1=>nx11357, B0
      =>d_arr_mul_9_25, B1=>nx10509, C0=>d_arr_add_9_25, C1=>nx10701);
   lat_d_arr_9_26 : latch port map ( Q=>d_arr_9_26, D=>nx4980, CLK=>nx10277
   );
   ix4981 : inv01 port map ( Y=>nx4980, A=>nx9057);
   ix9058 : aoi222 port map ( Y=>nx9057, A0=>d_arr_mux_9_26, A1=>nx11357, B0
      =>d_arr_mul_9_26, B1=>nx10509, C0=>d_arr_add_9_26, C1=>nx10701);
   lat_d_arr_9_27 : latch port map ( Q=>d_arr_9_27, D=>nx4992, CLK=>nx10277
   );
   ix4993 : inv01 port map ( Y=>nx4992, A=>nx9061);
   ix9062 : aoi222 port map ( Y=>nx9061, A0=>d_arr_mux_9_27, A1=>nx11357, B0
      =>d_arr_mul_9_27, B1=>nx10509, C0=>d_arr_add_9_27, C1=>nx10701);
   lat_d_arr_9_28 : latch port map ( Q=>d_arr_9_28, D=>nx5004, CLK=>nx10277
   );
   ix5005 : inv01 port map ( Y=>nx5004, A=>nx9065);
   ix9066 : aoi222 port map ( Y=>nx9065, A0=>d_arr_mux_9_28, A1=>nx11357, B0
      =>d_arr_mul_9_28, B1=>nx10509, C0=>d_arr_add_9_28, C1=>nx10701);
   lat_d_arr_9_29 : latch port map ( Q=>d_arr_9_29, D=>nx5016, CLK=>nx10277
   );
   ix5017 : inv01 port map ( Y=>nx5016, A=>nx9069);
   ix9070 : aoi222 port map ( Y=>nx9069, A0=>d_arr_mux_9_29, A1=>nx11357, B0
      =>d_arr_mul_9_29, B1=>nx10509, C0=>d_arr_add_9_29, C1=>nx10701);
   lat_d_arr_9_30 : latch port map ( Q=>d_arr_9_30, D=>nx5028, CLK=>nx10277
   );
   ix5029 : inv01 port map ( Y=>nx5028, A=>nx9073);
   ix9074 : aoi222 port map ( Y=>nx9073, A0=>d_arr_mux_9_30, A1=>nx11357, B0
      =>d_arr_mul_9_30, B1=>nx10509, C0=>d_arr_add_9_30, C1=>nx10701);
   lat_d_arr_9_31 : latch port map ( Q=>d_arr_9_31, D=>nx5040, CLK=>nx10279
   );
   ix5041 : inv01 port map ( Y=>nx5040, A=>nx9077);
   ix9078 : aoi222 port map ( Y=>nx9077, A0=>d_arr_mux_9_31, A1=>nx11357, B0
      =>d_arr_mul_9_31, B1=>nx10511, C0=>d_arr_add_9_31, C1=>nx10703);
   lat_d_arr_8_0 : latch port map ( Q=>d_arr_8_0, D=>nx5048, CLK=>nx10279);
   ix5049 : ao22 port map ( Y=>nx5048, A0=>d_arr_mux_8_0, A1=>nx11359, B0=>
      d_arr_mul_8_0, B1=>nx10511);
   lat_d_arr_8_1 : latch port map ( Q=>d_arr_8_1, D=>nx5056, CLK=>nx10279);
   ix5057 : ao22 port map ( Y=>nx5056, A0=>d_arr_mux_8_1, A1=>nx11359, B0=>
      d_arr_mul_8_1, B1=>nx10511);
   lat_d_arr_8_2 : latch port map ( Q=>d_arr_8_2, D=>nx5064, CLK=>nx10279);
   ix5065 : ao22 port map ( Y=>nx5064, A0=>d_arr_mux_8_2, A1=>nx11359, B0=>
      d_arr_mul_8_2, B1=>nx10511);
   lat_d_arr_8_3 : latch port map ( Q=>d_arr_8_3, D=>nx5072, CLK=>nx10279);
   ix5073 : ao22 port map ( Y=>nx5072, A0=>d_arr_mux_8_3, A1=>nx11359, B0=>
      d_arr_mul_8_3, B1=>nx10511);
   lat_d_arr_8_4 : latch port map ( Q=>d_arr_8_4, D=>nx5080, CLK=>nx10279);
   ix5081 : ao22 port map ( Y=>nx5080, A0=>d_arr_mux_8_4, A1=>nx11359, B0=>
      d_arr_mul_8_4, B1=>nx10511);
   lat_d_arr_8_5 : latch port map ( Q=>d_arr_8_5, D=>nx5088, CLK=>nx10279);
   ix5089 : ao22 port map ( Y=>nx5088, A0=>d_arr_mux_8_5, A1=>nx11359, B0=>
      d_arr_mul_8_5, B1=>nx10511);
   lat_d_arr_8_6 : latch port map ( Q=>d_arr_8_6, D=>nx5096, CLK=>nx10281);
   ix5097 : ao22 port map ( Y=>nx5096, A0=>d_arr_mux_8_6, A1=>nx11359, B0=>
      d_arr_mul_8_6, B1=>nx10513);
   lat_d_arr_8_7 : latch port map ( Q=>d_arr_8_7, D=>nx5104, CLK=>nx10281);
   ix5105 : ao22 port map ( Y=>nx5104, A0=>d_arr_mux_8_7, A1=>nx11361, B0=>
      d_arr_mul_8_7, B1=>nx10513);
   lat_d_arr_8_8 : latch port map ( Q=>d_arr_8_8, D=>nx5112, CLK=>nx10281);
   ix5113 : ao22 port map ( Y=>nx5112, A0=>d_arr_mux_8_8, A1=>nx11361, B0=>
      d_arr_mul_8_8, B1=>nx10513);
   lat_d_arr_8_9 : latch port map ( Q=>d_arr_8_9, D=>nx5120, CLK=>nx10281);
   ix5121 : ao22 port map ( Y=>nx5120, A0=>d_arr_mux_8_9, A1=>nx11361, B0=>
      d_arr_mul_8_9, B1=>nx10513);
   lat_d_arr_8_10 : latch port map ( Q=>d_arr_8_10, D=>nx5128, CLK=>nx10281
   );
   ix5129 : ao22 port map ( Y=>nx5128, A0=>d_arr_mux_8_10, A1=>nx11361, B0=>
      d_arr_mul_8_10, B1=>nx10513);
   lat_d_arr_8_11 : latch port map ( Q=>d_arr_8_11, D=>nx5136, CLK=>nx10281
   );
   ix5137 : ao22 port map ( Y=>nx5136, A0=>d_arr_mux_8_11, A1=>nx11361, B0=>
      d_arr_mul_8_11, B1=>nx10513);
   lat_d_arr_8_12 : latch port map ( Q=>d_arr_8_12, D=>nx5144, CLK=>nx10281
   );
   ix5145 : ao22 port map ( Y=>nx5144, A0=>d_arr_mux_8_12, A1=>nx11361, B0=>
      d_arr_mul_8_12, B1=>nx10513);
   lat_d_arr_8_13 : latch port map ( Q=>d_arr_8_13, D=>nx5152, CLK=>nx10283
   );
   ix5153 : ao22 port map ( Y=>nx5152, A0=>d_arr_mux_8_13, A1=>nx11361, B0=>
      d_arr_mul_8_13, B1=>nx10515);
   lat_d_arr_8_14 : latch port map ( Q=>d_arr_8_14, D=>nx5160, CLK=>nx10283
   );
   ix5161 : ao22 port map ( Y=>nx5160, A0=>d_arr_mux_8_14, A1=>nx11363, B0=>
      d_arr_mul_8_14, B1=>nx10515);
   lat_d_arr_8_15 : latch port map ( Q=>d_arr_8_15, D=>nx5168, CLK=>nx10283
   );
   lat_d_arr_8_16 : latch port map ( Q=>d_arr_8_16, D=>nx5174, CLK=>nx10283
   );
   lat_d_arr_8_17 : latch port map ( Q=>d_arr_8_17, D=>nx5180, CLK=>nx10283
   );
   lat_d_arr_8_18 : latch port map ( Q=>d_arr_8_18, D=>nx5186, CLK=>nx10283
   );
   lat_d_arr_8_19 : latch port map ( Q=>d_arr_8_19, D=>nx5192, CLK=>nx10283
   );
   lat_d_arr_8_20 : latch port map ( Q=>d_arr_8_20, D=>nx5198, CLK=>nx10285
   );
   lat_d_arr_8_21 : latch port map ( Q=>d_arr_8_21, D=>nx5204, CLK=>nx10285
   );
   lat_d_arr_8_22 : latch port map ( Q=>d_arr_8_22, D=>nx5210, CLK=>nx10285
   );
   lat_d_arr_8_23 : latch port map ( Q=>d_arr_8_23, D=>nx5216, CLK=>nx10285
   );
   lat_d_arr_8_24 : latch port map ( Q=>d_arr_8_24, D=>nx5222, CLK=>nx10285
   );
   lat_d_arr_8_25 : latch port map ( Q=>d_arr_8_25, D=>nx5228, CLK=>nx10285
   );
   lat_d_arr_8_26 : latch port map ( Q=>d_arr_8_26, D=>nx5234, CLK=>nx10285
   );
   lat_d_arr_8_27 : latch port map ( Q=>d_arr_8_27, D=>nx5240, CLK=>nx10287
   );
   lat_d_arr_8_28 : latch port map ( Q=>d_arr_8_28, D=>nx5246, CLK=>nx10287
   );
   lat_d_arr_8_29 : latch port map ( Q=>d_arr_8_29, D=>nx5252, CLK=>nx10287
   );
   lat_d_arr_8_30 : latch port map ( Q=>d_arr_8_30, D=>nx5258, CLK=>nx10287
   );
   lat_d_arr_8_31 : latch port map ( Q=>d_arr_8_31, D=>nx5264, CLK=>nx10287
   );
   lat_d_arr_7_0 : latch port map ( Q=>d_arr_7_0, D=>nx5272, CLK=>nx10287);
   ix5273 : ao22 port map ( Y=>nx5272, A0=>d_arr_mux_7_0, A1=>nx11363, B0=>
      d_arr_mul_7_0, B1=>nx10519);
   lat_d_arr_7_1 : latch port map ( Q=>d_arr_7_1, D=>nx5280, CLK=>nx10287);
   ix5281 : ao22 port map ( Y=>nx5280, A0=>d_arr_mux_7_1, A1=>nx11363, B0=>
      d_arr_mul_7_1, B1=>nx10519);
   lat_d_arr_7_2 : latch port map ( Q=>d_arr_7_2, D=>nx5288, CLK=>nx10289);
   ix5289 : ao22 port map ( Y=>nx5288, A0=>d_arr_mux_7_2, A1=>nx11363, B0=>
      d_arr_mul_7_2, B1=>nx10521);
   lat_d_arr_7_3 : latch port map ( Q=>d_arr_7_3, D=>nx5296, CLK=>nx10289);
   ix5297 : ao22 port map ( Y=>nx5296, A0=>d_arr_mux_7_3, A1=>nx11363, B0=>
      d_arr_mul_7_3, B1=>nx10521);
   lat_d_arr_7_4 : latch port map ( Q=>d_arr_7_4, D=>nx5304, CLK=>nx10289);
   ix5305 : ao22 port map ( Y=>nx5304, A0=>d_arr_mux_7_4, A1=>nx11363, B0=>
      d_arr_mul_7_4, B1=>nx10521);
   lat_d_arr_7_5 : latch port map ( Q=>d_arr_7_5, D=>nx5312, CLK=>nx10289);
   ix5313 : ao22 port map ( Y=>nx5312, A0=>d_arr_mux_7_5, A1=>nx11363, B0=>
      d_arr_mul_7_5, B1=>nx10521);
   lat_d_arr_7_6 : latch port map ( Q=>d_arr_7_6, D=>nx5320, CLK=>nx10289);
   ix5321 : ao22 port map ( Y=>nx5320, A0=>d_arr_mux_7_6, A1=>nx11365, B0=>
      d_arr_mul_7_6, B1=>nx10521);
   lat_d_arr_7_7 : latch port map ( Q=>d_arr_7_7, D=>nx5328, CLK=>nx10289);
   ix5329 : ao22 port map ( Y=>nx5328, A0=>d_arr_mux_7_7, A1=>nx11365, B0=>
      d_arr_mul_7_7, B1=>nx10521);
   lat_d_arr_7_8 : latch port map ( Q=>d_arr_7_8, D=>nx5336, CLK=>nx10289);
   ix5337 : ao22 port map ( Y=>nx5336, A0=>d_arr_mux_7_8, A1=>nx11365, B0=>
      d_arr_mul_7_8, B1=>nx10521);
   lat_d_arr_7_9 : latch port map ( Q=>d_arr_7_9, D=>nx5344, CLK=>nx10291);
   ix5345 : ao22 port map ( Y=>nx5344, A0=>d_arr_mux_7_9, A1=>nx11365, B0=>
      d_arr_mul_7_9, B1=>nx10523);
   lat_d_arr_7_10 : latch port map ( Q=>d_arr_7_10, D=>nx5352, CLK=>nx10291
   );
   ix5353 : ao22 port map ( Y=>nx5352, A0=>d_arr_mux_7_10, A1=>nx11365, B0=>
      d_arr_mul_7_10, B1=>nx10523);
   lat_d_arr_7_11 : latch port map ( Q=>d_arr_7_11, D=>nx5360, CLK=>nx10291
   );
   ix5361 : ao22 port map ( Y=>nx5360, A0=>d_arr_mux_7_11, A1=>nx11365, B0=>
      d_arr_mul_7_11, B1=>nx10523);
   lat_d_arr_7_12 : latch port map ( Q=>d_arr_7_12, D=>nx5368, CLK=>nx10291
   );
   ix5369 : ao22 port map ( Y=>nx5368, A0=>d_arr_mux_7_12, A1=>nx11365, B0=>
      d_arr_mul_7_12, B1=>nx10523);
   lat_d_arr_7_13 : latch port map ( Q=>d_arr_7_13, D=>nx5376, CLK=>nx10291
   );
   ix5377 : ao22 port map ( Y=>nx5376, A0=>d_arr_mux_7_13, A1=>nx11367, B0=>
      d_arr_mul_7_13, B1=>nx10523);
   lat_d_arr_7_14 : latch port map ( Q=>d_arr_7_14, D=>nx5384, CLK=>nx10291
   );
   ix5385 : ao22 port map ( Y=>nx5384, A0=>d_arr_mux_7_14, A1=>nx11367, B0=>
      d_arr_mul_7_14, B1=>nx10523);
   lat_d_arr_7_15 : latch port map ( Q=>d_arr_7_15, D=>nx5392, CLK=>nx10291
   );
   lat_d_arr_7_16 : latch port map ( Q=>d_arr_7_16, D=>nx5398, CLK=>nx10293
   );
   lat_d_arr_7_17 : latch port map ( Q=>d_arr_7_17, D=>nx5404, CLK=>nx10293
   );
   lat_d_arr_7_18 : latch port map ( Q=>d_arr_7_18, D=>nx5410, CLK=>nx10293
   );
   lat_d_arr_7_19 : latch port map ( Q=>d_arr_7_19, D=>nx5416, CLK=>nx10293
   );
   lat_d_arr_7_20 : latch port map ( Q=>d_arr_7_20, D=>nx5422, CLK=>nx10293
   );
   lat_d_arr_7_21 : latch port map ( Q=>d_arr_7_21, D=>nx5428, CLK=>nx10293
   );
   lat_d_arr_7_22 : latch port map ( Q=>d_arr_7_22, D=>nx5434, CLK=>nx10293
   );
   lat_d_arr_7_23 : latch port map ( Q=>d_arr_7_23, D=>nx5440, CLK=>nx10295
   );
   lat_d_arr_7_24 : latch port map ( Q=>d_arr_7_24, D=>nx5446, CLK=>nx10295
   );
   lat_d_arr_7_25 : latch port map ( Q=>d_arr_7_25, D=>nx5452, CLK=>nx10295
   );
   lat_d_arr_7_26 : latch port map ( Q=>d_arr_7_26, D=>nx5458, CLK=>nx10295
   );
   lat_d_arr_7_27 : latch port map ( Q=>d_arr_7_27, D=>nx5464, CLK=>nx10295
   );
   lat_d_arr_7_28 : latch port map ( Q=>d_arr_7_28, D=>nx5470, CLK=>nx10295
   );
   lat_d_arr_7_29 : latch port map ( Q=>d_arr_7_29, D=>nx5476, CLK=>nx10295
   );
   lat_d_arr_7_30 : latch port map ( Q=>d_arr_7_30, D=>nx5482, CLK=>nx10297
   );
   lat_d_arr_7_31 : latch port map ( Q=>d_arr_7_31, D=>nx5488, CLK=>nx10297
   );
   lat_d_arr_6_0 : latch port map ( Q=>d_arr_6_0, D=>nx5496, CLK=>nx10297);
   ix5497 : ao22 port map ( Y=>nx5496, A0=>d_arr_mux_6_0, A1=>nx11367, B0=>
      d_arr_mul_6_0, B1=>nx10529);
   lat_d_arr_6_1 : latch port map ( Q=>d_arr_6_1, D=>nx5504, CLK=>nx10297);
   ix5505 : ao22 port map ( Y=>nx5504, A0=>d_arr_mux_6_1, A1=>nx11367, B0=>
      d_arr_mul_6_1, B1=>nx10529);
   lat_d_arr_6_2 : latch port map ( Q=>d_arr_6_2, D=>nx5512, CLK=>nx10297);
   ix5513 : ao22 port map ( Y=>nx5512, A0=>d_arr_mux_6_2, A1=>nx11367, B0=>
      d_arr_mul_6_2, B1=>nx10529);
   lat_d_arr_6_3 : latch port map ( Q=>d_arr_6_3, D=>nx5520, CLK=>nx10297);
   ix5521 : ao22 port map ( Y=>nx5520, A0=>d_arr_mux_6_3, A1=>nx11367, B0=>
      d_arr_mul_6_3, B1=>nx10529);
   lat_d_arr_6_4 : latch port map ( Q=>d_arr_6_4, D=>nx5528, CLK=>nx10297);
   ix5529 : ao22 port map ( Y=>nx5528, A0=>d_arr_mux_6_4, A1=>nx11367, B0=>
      d_arr_mul_6_4, B1=>nx10529);
   lat_d_arr_6_5 : latch port map ( Q=>d_arr_6_5, D=>nx5536, CLK=>nx10299);
   ix5537 : ao22 port map ( Y=>nx5536, A0=>d_arr_mux_6_5, A1=>nx11369, B0=>
      d_arr_mul_6_5, B1=>nx10531);
   lat_d_arr_6_6 : latch port map ( Q=>d_arr_6_6, D=>nx5544, CLK=>nx10299);
   ix5545 : ao22 port map ( Y=>nx5544, A0=>d_arr_mux_6_6, A1=>nx11369, B0=>
      d_arr_mul_6_6, B1=>nx10531);
   lat_d_arr_6_7 : latch port map ( Q=>d_arr_6_7, D=>nx5552, CLK=>nx10299);
   ix5553 : ao22 port map ( Y=>nx5552, A0=>d_arr_mux_6_7, A1=>nx11369, B0=>
      d_arr_mul_6_7, B1=>nx10531);
   lat_d_arr_6_8 : latch port map ( Q=>d_arr_6_8, D=>nx5560, CLK=>nx10299);
   ix5561 : ao22 port map ( Y=>nx5560, A0=>d_arr_mux_6_8, A1=>nx11369, B0=>
      d_arr_mul_6_8, B1=>nx10531);
   lat_d_arr_6_9 : latch port map ( Q=>d_arr_6_9, D=>nx5568, CLK=>nx10299);
   ix5569 : ao22 port map ( Y=>nx5568, A0=>d_arr_mux_6_9, A1=>nx11369, B0=>
      d_arr_mul_6_9, B1=>nx10531);
   lat_d_arr_6_10 : latch port map ( Q=>d_arr_6_10, D=>nx5576, CLK=>nx10299
   );
   ix5577 : ao22 port map ( Y=>nx5576, A0=>d_arr_mux_6_10, A1=>nx11369, B0=>
      d_arr_mul_6_10, B1=>nx10531);
   lat_d_arr_6_11 : latch port map ( Q=>d_arr_6_11, D=>nx5584, CLK=>nx10299
   );
   ix5585 : ao22 port map ( Y=>nx5584, A0=>d_arr_mux_6_11, A1=>nx11369, B0=>
      d_arr_mul_6_11, B1=>nx10531);
   lat_d_arr_6_12 : latch port map ( Q=>d_arr_6_12, D=>nx5592, CLK=>nx10301
   );
   ix5593 : ao22 port map ( Y=>nx5592, A0=>d_arr_mux_6_12, A1=>nx11371, B0=>
      d_arr_mul_6_12, B1=>nx10533);
   lat_d_arr_6_13 : latch port map ( Q=>d_arr_6_13, D=>nx5600, CLK=>nx10301
   );
   ix5601 : ao22 port map ( Y=>nx5600, A0=>d_arr_mux_6_13, A1=>nx11371, B0=>
      d_arr_mul_6_13, B1=>nx10533);
   lat_d_arr_6_14 : latch port map ( Q=>d_arr_6_14, D=>nx5608, CLK=>nx10301
   );
   ix5609 : ao22 port map ( Y=>nx5608, A0=>d_arr_mux_6_14, A1=>nx11371, B0=>
      d_arr_mul_6_14, B1=>nx10533);
   lat_d_arr_6_15 : latch port map ( Q=>d_arr_6_15, D=>nx5616, CLK=>nx10301
   );
   lat_d_arr_6_16 : latch port map ( Q=>d_arr_6_16, D=>nx5622, CLK=>nx10301
   );
   lat_d_arr_6_17 : latch port map ( Q=>d_arr_6_17, D=>nx5628, CLK=>nx10301
   );
   lat_d_arr_6_18 : latch port map ( Q=>d_arr_6_18, D=>nx5634, CLK=>nx10301
   );
   lat_d_arr_6_19 : latch port map ( Q=>d_arr_6_19, D=>nx5640, CLK=>nx10303
   );
   lat_d_arr_6_20 : latch port map ( Q=>d_arr_6_20, D=>nx5646, CLK=>nx10303
   );
   lat_d_arr_6_21 : latch port map ( Q=>d_arr_6_21, D=>nx5652, CLK=>nx10303
   );
   lat_d_arr_6_22 : latch port map ( Q=>d_arr_6_22, D=>nx5658, CLK=>nx10303
   );
   lat_d_arr_6_23 : latch port map ( Q=>d_arr_6_23, D=>nx5664, CLK=>nx10303
   );
   lat_d_arr_6_24 : latch port map ( Q=>d_arr_6_24, D=>nx5670, CLK=>nx10303
   );
   lat_d_arr_6_25 : latch port map ( Q=>d_arr_6_25, D=>nx5676, CLK=>nx10303
   );
   lat_d_arr_6_26 : latch port map ( Q=>d_arr_6_26, D=>nx5682, CLK=>nx10305
   );
   lat_d_arr_6_27 : latch port map ( Q=>d_arr_6_27, D=>nx5688, CLK=>nx10305
   );
   lat_d_arr_6_28 : latch port map ( Q=>d_arr_6_28, D=>nx5694, CLK=>nx10305
   );
   lat_d_arr_6_29 : latch port map ( Q=>d_arr_6_29, D=>nx5700, CLK=>nx10305
   );
   lat_d_arr_6_30 : latch port map ( Q=>d_arr_6_30, D=>nx5706, CLK=>nx10305
   );
   lat_d_arr_6_31 : latch port map ( Q=>d_arr_6_31, D=>nx5712, CLK=>nx10305
   );
   lat_d_arr_5_0 : latch port map ( Q=>d_arr_5_0, D=>nx5720, CLK=>nx10305);
   ix5721 : ao22 port map ( Y=>nx5720, A0=>d_arr_mux_5_0, A1=>nx11371, B0=>
      d_arr_mul_5_0, B1=>nx10537);
   lat_d_arr_5_1 : latch port map ( Q=>d_arr_5_1, D=>nx5728, CLK=>nx10307);
   ix5729 : ao22 port map ( Y=>nx5728, A0=>d_arr_mux_5_1, A1=>nx11371, B0=>
      d_arr_mul_5_1, B1=>nx10539);
   lat_d_arr_5_2 : latch port map ( Q=>d_arr_5_2, D=>nx5736, CLK=>nx10307);
   ix5737 : ao22 port map ( Y=>nx5736, A0=>d_arr_mux_5_2, A1=>nx11371, B0=>
      d_arr_mul_5_2, B1=>nx10539);
   lat_d_arr_5_3 : latch port map ( Q=>d_arr_5_3, D=>nx5744, CLK=>nx10307);
   ix5745 : ao22 port map ( Y=>nx5744, A0=>d_arr_mux_5_3, A1=>nx11371, B0=>
      d_arr_mul_5_3, B1=>nx10539);
   lat_d_arr_5_4 : latch port map ( Q=>d_arr_5_4, D=>nx5752, CLK=>nx10307);
   ix5753 : ao22 port map ( Y=>nx5752, A0=>d_arr_mux_5_4, A1=>nx11373, B0=>
      d_arr_mul_5_4, B1=>nx10539);
   lat_d_arr_5_5 : latch port map ( Q=>d_arr_5_5, D=>nx5760, CLK=>nx10307);
   ix5761 : ao22 port map ( Y=>nx5760, A0=>d_arr_mux_5_5, A1=>nx11373, B0=>
      d_arr_mul_5_5, B1=>nx10539);
   lat_d_arr_5_6 : latch port map ( Q=>d_arr_5_6, D=>nx5768, CLK=>nx10307);
   ix5769 : ao22 port map ( Y=>nx5768, A0=>d_arr_mux_5_6, A1=>nx11373, B0=>
      d_arr_mul_5_6, B1=>nx10539);
   lat_d_arr_5_7 : latch port map ( Q=>d_arr_5_7, D=>nx5776, CLK=>nx10307);
   ix5777 : ao22 port map ( Y=>nx5776, A0=>d_arr_mux_5_7, A1=>nx11373, B0=>
      d_arr_mul_5_7, B1=>nx10539);
   lat_d_arr_5_8 : latch port map ( Q=>d_arr_5_8, D=>nx5784, CLK=>nx10309);
   ix5785 : ao22 port map ( Y=>nx5784, A0=>d_arr_mux_5_8, A1=>nx11373, B0=>
      d_arr_mul_5_8, B1=>nx10541);
   lat_d_arr_5_9 : latch port map ( Q=>d_arr_5_9, D=>nx5792, CLK=>nx10309);
   ix5793 : ao22 port map ( Y=>nx5792, A0=>d_arr_mux_5_9, A1=>nx11373, B0=>
      d_arr_mul_5_9, B1=>nx10541);
   lat_d_arr_5_10 : latch port map ( Q=>d_arr_5_10, D=>nx5800, CLK=>nx10309
   );
   ix5801 : ao22 port map ( Y=>nx5800, A0=>d_arr_mux_5_10, A1=>nx11373, B0=>
      d_arr_mul_5_10, B1=>nx10541);
   lat_d_arr_5_11 : latch port map ( Q=>d_arr_5_11, D=>nx5808, CLK=>nx10309
   );
   ix5809 : ao22 port map ( Y=>nx5808, A0=>d_arr_mux_5_11, A1=>nx11375, B0=>
      d_arr_mul_5_11, B1=>nx10541);
   lat_d_arr_5_12 : latch port map ( Q=>d_arr_5_12, D=>nx5816, CLK=>nx10309
   );
   ix5817 : ao22 port map ( Y=>nx5816, A0=>d_arr_mux_5_12, A1=>nx11375, B0=>
      d_arr_mul_5_12, B1=>nx10541);
   lat_d_arr_5_13 : latch port map ( Q=>d_arr_5_13, D=>nx5824, CLK=>nx10309
   );
   ix5825 : ao22 port map ( Y=>nx5824, A0=>d_arr_mux_5_13, A1=>nx11375, B0=>
      d_arr_mul_5_13, B1=>nx10541);
   lat_d_arr_5_14 : latch port map ( Q=>d_arr_5_14, D=>nx5832, CLK=>nx10309
   );
   ix5833 : ao22 port map ( Y=>nx5832, A0=>d_arr_mux_5_14, A1=>nx11375, B0=>
      d_arr_mul_5_14, B1=>nx10541);
   lat_d_arr_5_15 : latch port map ( Q=>d_arr_5_15, D=>nx5840, CLK=>nx10311
   );
   lat_d_arr_5_16 : latch port map ( Q=>d_arr_5_16, D=>nx5846, CLK=>nx10311
   );
   lat_d_arr_5_17 : latch port map ( Q=>d_arr_5_17, D=>nx5852, CLK=>nx10311
   );
   lat_d_arr_5_18 : latch port map ( Q=>d_arr_5_18, D=>nx5858, CLK=>nx10311
   );
   lat_d_arr_5_19 : latch port map ( Q=>d_arr_5_19, D=>nx5864, CLK=>nx10311
   );
   lat_d_arr_5_20 : latch port map ( Q=>d_arr_5_20, D=>nx5870, CLK=>nx10311
   );
   lat_d_arr_5_21 : latch port map ( Q=>d_arr_5_21, D=>nx5876, CLK=>nx10311
   );
   lat_d_arr_5_22 : latch port map ( Q=>d_arr_5_22, D=>nx5882, CLK=>nx10313
   );
   lat_d_arr_5_23 : latch port map ( Q=>d_arr_5_23, D=>nx5888, CLK=>nx10313
   );
   lat_d_arr_5_24 : latch port map ( Q=>d_arr_5_24, D=>nx5894, CLK=>nx10313
   );
   lat_d_arr_5_25 : latch port map ( Q=>d_arr_5_25, D=>nx5900, CLK=>nx10313
   );
   lat_d_arr_5_26 : latch port map ( Q=>d_arr_5_26, D=>nx5906, CLK=>nx10313
   );
   lat_d_arr_5_27 : latch port map ( Q=>d_arr_5_27, D=>nx5912, CLK=>nx10313
   );
   lat_d_arr_5_28 : latch port map ( Q=>d_arr_5_28, D=>nx5918, CLK=>nx10313
   );
   lat_d_arr_5_29 : latch port map ( Q=>d_arr_5_29, D=>nx5924, CLK=>nx10315
   );
   lat_d_arr_5_30 : latch port map ( Q=>d_arr_5_30, D=>nx5930, CLK=>nx10315
   );
   lat_d_arr_5_31 : latch port map ( Q=>d_arr_5_31, D=>nx5936, CLK=>nx10315
   );
   lat_d_arr_4_0 : latch port map ( Q=>d_arr_4_0, D=>nx5948, CLK=>nx10315);
   ix5949 : inv01 port map ( Y=>nx5948, A=>nx9341);
   ix9342 : aoi222 port map ( Y=>nx9341, A0=>d_arr_mux_4_0, A1=>nx11375, B0
      =>d_arr_mul_4_0, B1=>nx10547, C0=>d_arr_add_4_0, C1=>nx10703);
   lat_d_arr_4_1 : latch port map ( Q=>d_arr_4_1, D=>nx5960, CLK=>nx10315);
   ix5961 : inv01 port map ( Y=>nx5960, A=>nx9345);
   ix9346 : aoi222 port map ( Y=>nx9345, A0=>d_arr_mux_4_1, A1=>nx11375, B0
      =>d_arr_mul_4_1, B1=>nx10547, C0=>d_arr_add_4_1, C1=>nx10703);
   lat_d_arr_4_2 : latch port map ( Q=>d_arr_4_2, D=>nx5972, CLK=>nx10315);
   ix5973 : inv01 port map ( Y=>nx5972, A=>nx9349);
   ix9350 : aoi222 port map ( Y=>nx9349, A0=>d_arr_mux_4_2, A1=>nx11375, B0
      =>d_arr_mul_4_2, B1=>nx10547, C0=>d_arr_add_4_2, C1=>nx10703);
   lat_d_arr_4_3 : latch port map ( Q=>d_arr_4_3, D=>nx5984, CLK=>nx10315);
   ix5985 : inv01 port map ( Y=>nx5984, A=>nx9353);
   ix9354 : aoi222 port map ( Y=>nx9353, A0=>d_arr_mux_4_3, A1=>nx11377, B0
      =>d_arr_mul_4_3, B1=>nx10547, C0=>d_arr_add_4_3, C1=>nx10703);
   lat_d_arr_4_4 : latch port map ( Q=>d_arr_4_4, D=>nx5996, CLK=>nx10317);
   ix5997 : inv01 port map ( Y=>nx5996, A=>nx9357);
   ix9358 : aoi222 port map ( Y=>nx9357, A0=>d_arr_mux_4_4, A1=>nx11377, B0
      =>d_arr_mul_4_4, B1=>nx10549, C0=>d_arr_add_4_4, C1=>nx10703);
   lat_d_arr_4_5 : latch port map ( Q=>d_arr_4_5, D=>nx6008, CLK=>nx10317);
   ix6009 : inv01 port map ( Y=>nx6008, A=>nx9361);
   ix9362 : aoi222 port map ( Y=>nx9361, A0=>d_arr_mux_4_5, A1=>nx11377, B0
      =>d_arr_mul_4_5, B1=>nx10549, C0=>d_arr_add_4_5, C1=>nx10703);
   lat_d_arr_4_6 : latch port map ( Q=>d_arr_4_6, D=>nx6020, CLK=>nx10317);
   ix6021 : inv01 port map ( Y=>nx6020, A=>nx9365);
   ix9366 : aoi222 port map ( Y=>nx9365, A0=>d_arr_mux_4_6, A1=>nx11377, B0
      =>d_arr_mul_4_6, B1=>nx10549, C0=>d_arr_add_4_6, C1=>nx10705);
   lat_d_arr_4_7 : latch port map ( Q=>d_arr_4_7, D=>nx6032, CLK=>nx10317);
   ix6033 : inv01 port map ( Y=>nx6032, A=>nx9369);
   ix9370 : aoi222 port map ( Y=>nx9369, A0=>d_arr_mux_4_7, A1=>nx11377, B0
      =>d_arr_mul_4_7, B1=>nx10549, C0=>d_arr_add_4_7, C1=>nx10705);
   lat_d_arr_4_8 : latch port map ( Q=>d_arr_4_8, D=>nx6044, CLK=>nx10317);
   ix6045 : inv01 port map ( Y=>nx6044, A=>nx9373);
   ix9374 : aoi222 port map ( Y=>nx9373, A0=>d_arr_mux_4_8, A1=>nx11377, B0
      =>d_arr_mul_4_8, B1=>nx10549, C0=>d_arr_add_4_8, C1=>nx10705);
   lat_d_arr_4_9 : latch port map ( Q=>d_arr_4_9, D=>nx6056, CLK=>nx10317);
   ix6057 : inv01 port map ( Y=>nx6056, A=>nx9377);
   ix9378 : aoi222 port map ( Y=>nx9377, A0=>d_arr_mux_4_9, A1=>nx11377, B0
      =>d_arr_mul_4_9, B1=>nx10549, C0=>d_arr_add_4_9, C1=>nx10705);
   lat_d_arr_4_10 : latch port map ( Q=>d_arr_4_10, D=>nx6068, CLK=>nx10317
   );
   ix6069 : inv01 port map ( Y=>nx6068, A=>nx9381);
   ix9382 : aoi222 port map ( Y=>nx9381, A0=>d_arr_mux_4_10, A1=>nx11379, B0
      =>d_arr_mul_4_10, B1=>nx10549, C0=>d_arr_add_4_10, C1=>nx10705);
   lat_d_arr_4_11 : latch port map ( Q=>d_arr_4_11, D=>nx6080, CLK=>nx10319
   );
   ix6081 : inv01 port map ( Y=>nx6080, A=>nx9385);
   ix9386 : aoi222 port map ( Y=>nx9385, A0=>d_arr_mux_4_11, A1=>nx11379, B0
      =>d_arr_mul_4_11, B1=>nx10551, C0=>d_arr_add_4_11, C1=>nx10705);
   lat_d_arr_4_12 : latch port map ( Q=>d_arr_4_12, D=>nx6092, CLK=>nx10319
   );
   ix6093 : inv01 port map ( Y=>nx6092, A=>nx9389);
   ix9390 : aoi222 port map ( Y=>nx9389, A0=>d_arr_mux_4_12, A1=>nx11379, B0
      =>d_arr_mul_4_12, B1=>nx10551, C0=>d_arr_add_4_12, C1=>nx10705);
   lat_d_arr_4_13 : latch port map ( Q=>d_arr_4_13, D=>nx6104, CLK=>nx10319
   );
   ix6105 : inv01 port map ( Y=>nx6104, A=>nx9393);
   ix9394 : aoi222 port map ( Y=>nx9393, A0=>d_arr_mux_4_13, A1=>nx11379, B0
      =>d_arr_mul_4_13, B1=>nx10551, C0=>d_arr_add_4_13, C1=>nx10707);
   lat_d_arr_4_14 : latch port map ( Q=>d_arr_4_14, D=>nx6116, CLK=>nx10319
   );
   ix6117 : inv01 port map ( Y=>nx6116, A=>nx9397);
   ix9398 : aoi222 port map ( Y=>nx9397, A0=>d_arr_mux_4_14, A1=>nx11379, B0
      =>d_arr_mul_4_14, B1=>nx10551, C0=>d_arr_add_4_14, C1=>nx10707);
   lat_d_arr_4_15 : latch port map ( Q=>d_arr_4_15, D=>nx6128, CLK=>nx10319
   );
   ix6129 : nand02 port map ( Y=>nx6128, A0=>nx9401, A1=>nx10861);
   ix9402 : aoi22 port map ( Y=>nx9401, A0=>d_arr_mul_4_15, A1=>nx10551, B0
      =>d_arr_add_4_15, B1=>nx10707);
   ix9404 : nand02 port map ( Y=>nx9403, A0=>d_arr_mux_4_31, A1=>nx11379);
   lat_d_arr_4_16 : latch port map ( Q=>d_arr_4_16, D=>nx6138, CLK=>nx10319
   );
   ix6139 : nand02 port map ( Y=>nx6138, A0=>nx9407, A1=>nx10861);
   ix9408 : aoi22 port map ( Y=>nx9407, A0=>d_arr_mul_4_16, A1=>nx10551, B0
      =>d_arr_add_4_16, B1=>nx10707);
   lat_d_arr_4_17 : latch port map ( Q=>d_arr_4_17, D=>nx6148, CLK=>nx10319
   );
   ix6149 : nand02 port map ( Y=>nx6148, A0=>nx9411, A1=>nx10861);
   ix9412 : aoi22 port map ( Y=>nx9411, A0=>d_arr_mul_4_17, A1=>nx10551, B0
      =>d_arr_add_4_17, B1=>nx10707);
   lat_d_arr_4_18 : latch port map ( Q=>d_arr_4_18, D=>nx6158, CLK=>nx10321
   );
   ix6159 : nand02 port map ( Y=>nx6158, A0=>nx9415, A1=>nx10861);
   ix9416 : aoi22 port map ( Y=>nx9415, A0=>d_arr_mul_4_18, A1=>nx10553, B0
      =>d_arr_add_4_18, B1=>nx10707);
   lat_d_arr_4_19 : latch port map ( Q=>d_arr_4_19, D=>nx6168, CLK=>nx10321
   );
   ix6169 : nand02 port map ( Y=>nx6168, A0=>nx9419, A1=>nx10861);
   ix9420 : aoi22 port map ( Y=>nx9419, A0=>d_arr_mul_4_19, A1=>nx10553, B0
      =>d_arr_add_4_19, B1=>nx10707);
   lat_d_arr_4_20 : latch port map ( Q=>d_arr_4_20, D=>nx6178, CLK=>nx10321
   );
   ix6179 : nand02 port map ( Y=>nx6178, A0=>nx9423, A1=>nx10861);
   ix9424 : aoi22 port map ( Y=>nx9423, A0=>d_arr_mul_4_20, A1=>nx10553, B0
      =>d_arr_add_4_20, B1=>nx10709);
   lat_d_arr_4_21 : latch port map ( Q=>d_arr_4_21, D=>nx6188, CLK=>nx10321
   );
   ix6189 : nand02 port map ( Y=>nx6188, A0=>nx9427, A1=>nx10861);
   ix9428 : aoi22 port map ( Y=>nx9427, A0=>d_arr_mul_4_21, A1=>nx10553, B0
      =>d_arr_add_4_21, B1=>nx10709);
   lat_d_arr_4_22 : latch port map ( Q=>d_arr_4_22, D=>nx6198, CLK=>nx10321
   );
   ix6199 : nand02 port map ( Y=>nx6198, A0=>nx9431, A1=>nx10863);
   ix9432 : aoi22 port map ( Y=>nx9431, A0=>d_arr_mul_4_22, A1=>nx10553, B0
      =>d_arr_add_4_22, B1=>nx10709);
   lat_d_arr_4_23 : latch port map ( Q=>d_arr_4_23, D=>nx6208, CLK=>nx10321
   );
   ix6209 : nand02 port map ( Y=>nx6208, A0=>nx9435, A1=>nx10863);
   ix9436 : aoi22 port map ( Y=>nx9435, A0=>d_arr_mul_4_23, A1=>nx10553, B0
      =>d_arr_add_4_23, B1=>nx10709);
   lat_d_arr_4_24 : latch port map ( Q=>d_arr_4_24, D=>nx6218, CLK=>nx10321
   );
   ix6219 : nand02 port map ( Y=>nx6218, A0=>nx9439, A1=>nx10863);
   ix9440 : aoi22 port map ( Y=>nx9439, A0=>d_arr_mul_4_24, A1=>nx10553, B0
      =>d_arr_add_4_24, B1=>nx10709);
   lat_d_arr_4_25 : latch port map ( Q=>d_arr_4_25, D=>nx6228, CLK=>nx10323
   );
   ix6229 : nand02 port map ( Y=>nx6228, A0=>nx9443, A1=>nx10863);
   ix9444 : aoi22 port map ( Y=>nx9443, A0=>d_arr_mul_4_25, A1=>nx10555, B0
      =>d_arr_add_4_25, B1=>nx10709);
   lat_d_arr_4_26 : latch port map ( Q=>d_arr_4_26, D=>nx6238, CLK=>nx10323
   );
   ix6239 : nand02 port map ( Y=>nx6238, A0=>nx9447, A1=>nx10863);
   ix9448 : aoi22 port map ( Y=>nx9447, A0=>d_arr_mul_4_26, A1=>nx10555, B0
      =>d_arr_add_4_26, B1=>nx10709);
   lat_d_arr_4_27 : latch port map ( Q=>d_arr_4_27, D=>nx6248, CLK=>nx10323
   );
   ix6249 : nand02 port map ( Y=>nx6248, A0=>nx9451, A1=>nx10863);
   ix9452 : aoi22 port map ( Y=>nx9451, A0=>d_arr_mul_4_27, A1=>nx10555, B0
      =>d_arr_add_4_27, B1=>nx10711);
   lat_d_arr_4_28 : latch port map ( Q=>d_arr_4_28, D=>nx6258, CLK=>nx10323
   );
   ix6259 : nand02 port map ( Y=>nx6258, A0=>nx9455, A1=>nx10863);
   ix9456 : aoi22 port map ( Y=>nx9455, A0=>d_arr_mul_4_28, A1=>nx10555, B0
      =>d_arr_add_4_28, B1=>nx10711);
   lat_d_arr_4_29 : latch port map ( Q=>d_arr_4_29, D=>nx6268, CLK=>nx10323
   );
   ix6269 : nand02 port map ( Y=>nx6268, A0=>nx9459, A1=>nx9403);
   ix9460 : aoi22 port map ( Y=>nx9459, A0=>d_arr_mul_4_29, A1=>nx10555, B0
      =>d_arr_add_4_29, B1=>nx10711);
   lat_d_arr_4_30 : latch port map ( Q=>d_arr_4_30, D=>nx6278, CLK=>nx10323
   );
   ix6279 : nand02 port map ( Y=>nx6278, A0=>nx9463, A1=>nx9403);
   ix9464 : aoi22 port map ( Y=>nx9463, A0=>d_arr_mul_4_30, A1=>nx10555, B0
      =>d_arr_add_4_30, B1=>nx10711);
   lat_d_arr_4_31 : latch port map ( Q=>d_arr_4_31, D=>nx6288, CLK=>nx10323
   );
   ix6289 : nand02 port map ( Y=>nx6288, A0=>nx9467, A1=>nx9403);
   ix9468 : aoi22 port map ( Y=>nx9467, A0=>d_arr_mul_4_31, A1=>nx10555, B0
      =>d_arr_add_4_31, B1=>nx10711);
   lat_d_arr_3_0 : latch port map ( Q=>d_arr_3_0, D=>nx6300, CLK=>nx10325);
   ix6301 : inv01 port map ( Y=>nx6300, A=>nx9471);
   ix9472 : aoi222 port map ( Y=>nx9471, A0=>d_arr_mux_3_0, A1=>nx11379, B0
      =>d_arr_mul_3_0, B1=>nx10557, C0=>d_arr_add_3_0, C1=>nx10711);
   lat_d_arr_3_1 : latch port map ( Q=>d_arr_3_1, D=>nx6312, CLK=>nx10325);
   ix6313 : inv01 port map ( Y=>nx6312, A=>nx9475);
   ix9476 : aoi222 port map ( Y=>nx9475, A0=>d_arr_mux_3_1, A1=>nx11381, B0
      =>d_arr_mul_3_1, B1=>nx10557, C0=>d_arr_add_3_1, C1=>nx10711);
   lat_d_arr_3_2 : latch port map ( Q=>d_arr_3_2, D=>nx6324, CLK=>nx10325);
   ix6325 : inv01 port map ( Y=>nx6324, A=>nx9479);
   ix9480 : aoi222 port map ( Y=>nx9479, A0=>d_arr_mux_3_2, A1=>nx11381, B0
      =>d_arr_mul_3_2, B1=>nx10557, C0=>d_arr_add_3_2, C1=>nx10713);
   lat_d_arr_3_3 : latch port map ( Q=>d_arr_3_3, D=>nx6336, CLK=>nx10325);
   ix6337 : inv01 port map ( Y=>nx6336, A=>nx9483);
   ix9484 : aoi222 port map ( Y=>nx9483, A0=>d_arr_mux_3_3, A1=>nx11381, B0
      =>d_arr_mul_3_3, B1=>nx10557, C0=>d_arr_add_3_3, C1=>nx10713);
   lat_d_arr_3_4 : latch port map ( Q=>d_arr_3_4, D=>nx6348, CLK=>nx10325);
   ix6349 : inv01 port map ( Y=>nx6348, A=>nx9487);
   ix9488 : aoi222 port map ( Y=>nx9487, A0=>d_arr_mux_3_4, A1=>nx11381, B0
      =>d_arr_mul_3_4, B1=>nx10557, C0=>d_arr_add_3_4, C1=>nx10713);
   lat_d_arr_3_5 : latch port map ( Q=>d_arr_3_5, D=>nx6360, CLK=>nx10325);
   ix6361 : inv01 port map ( Y=>nx6360, A=>nx9491);
   ix9492 : aoi222 port map ( Y=>nx9491, A0=>d_arr_mux_3_5, A1=>nx11381, B0
      =>d_arr_mul_3_5, B1=>nx10557, C0=>d_arr_add_3_5, C1=>nx10713);
   lat_d_arr_3_6 : latch port map ( Q=>d_arr_3_6, D=>nx6372, CLK=>nx10325);
   ix6373 : inv01 port map ( Y=>nx6372, A=>nx9495);
   ix9496 : aoi222 port map ( Y=>nx9495, A0=>d_arr_mux_3_6, A1=>nx11381, B0
      =>d_arr_mul_3_6, B1=>nx10557, C0=>d_arr_add_3_6, C1=>nx10713);
   lat_d_arr_3_7 : latch port map ( Q=>d_arr_3_7, D=>nx6384, CLK=>nx10327);
   ix6385 : inv01 port map ( Y=>nx6384, A=>nx9499);
   ix9500 : aoi222 port map ( Y=>nx9499, A0=>d_arr_mux_3_7, A1=>nx11381, B0
      =>d_arr_mul_3_7, B1=>nx10559, C0=>d_arr_add_3_7, C1=>nx10713);
   lat_d_arr_3_8 : latch port map ( Q=>d_arr_3_8, D=>nx6396, CLK=>nx10327);
   ix6397 : inv01 port map ( Y=>nx6396, A=>nx9503);
   ix9504 : aoi222 port map ( Y=>nx9503, A0=>d_arr_mux_3_8, A1=>nx11383, B0
      =>d_arr_mul_3_8, B1=>nx10559, C0=>d_arr_add_3_8, C1=>nx10713);
   lat_d_arr_3_9 : latch port map ( Q=>d_arr_3_9, D=>nx6408, CLK=>nx10327);
   ix6409 : inv01 port map ( Y=>nx6408, A=>nx9507);
   ix9508 : aoi222 port map ( Y=>nx9507, A0=>d_arr_mux_3_9, A1=>nx11383, B0
      =>d_arr_mul_3_9, B1=>nx10559, C0=>d_arr_add_3_9, C1=>nx10715);
   lat_d_arr_3_10 : latch port map ( Q=>d_arr_3_10, D=>nx6420, CLK=>nx10327
   );
   ix6421 : inv01 port map ( Y=>nx6420, A=>nx9511);
   ix9512 : aoi222 port map ( Y=>nx9511, A0=>d_arr_mux_3_10, A1=>nx11383, B0
      =>d_arr_mul_3_10, B1=>nx10559, C0=>d_arr_add_3_10, C1=>nx10715);
   lat_d_arr_3_11 : latch port map ( Q=>d_arr_3_11, D=>nx6432, CLK=>nx10327
   );
   ix6433 : inv01 port map ( Y=>nx6432, A=>nx9515);
   ix9516 : aoi222 port map ( Y=>nx9515, A0=>d_arr_mux_3_11, A1=>nx11383, B0
      =>d_arr_mul_3_11, B1=>nx10559, C0=>d_arr_add_3_11, C1=>nx10715);
   lat_d_arr_3_12 : latch port map ( Q=>d_arr_3_12, D=>nx6444, CLK=>nx10327
   );
   ix6445 : inv01 port map ( Y=>nx6444, A=>nx9519);
   ix9520 : aoi222 port map ( Y=>nx9519, A0=>d_arr_mux_3_12, A1=>nx11383, B0
      =>d_arr_mul_3_12, B1=>nx10559, C0=>d_arr_add_3_12, C1=>nx10715);
   lat_d_arr_3_13 : latch port map ( Q=>d_arr_3_13, D=>nx6456, CLK=>nx10327
   );
   ix6457 : inv01 port map ( Y=>nx6456, A=>nx9523);
   ix9524 : aoi222 port map ( Y=>nx9523, A0=>d_arr_mux_3_13, A1=>nx11383, B0
      =>d_arr_mul_3_13, B1=>nx10559, C0=>d_arr_add_3_13, C1=>nx10715);
   lat_d_arr_3_14 : latch port map ( Q=>d_arr_3_14, D=>nx6468, CLK=>nx10329
   );
   ix6469 : inv01 port map ( Y=>nx6468, A=>nx9527);
   ix9528 : aoi222 port map ( Y=>nx9527, A0=>d_arr_mux_3_14, A1=>nx11383, B0
      =>d_arr_mul_3_14, B1=>nx10561, C0=>d_arr_add_3_14, C1=>nx10715);
   lat_d_arr_3_15 : latch port map ( Q=>d_arr_3_15, D=>nx6480, CLK=>nx10329
   );
   ix6481 : nand02 port map ( Y=>nx6480, A0=>nx9531, A1=>nx10865);
   ix9532 : aoi22 port map ( Y=>nx9531, A0=>d_arr_mul_3_15, A1=>nx10561, B0
      =>d_arr_add_3_15, B1=>nx10715);
   ix9534 : nand02 port map ( Y=>nx9533, A0=>d_arr_mux_3_31, A1=>nx11385);
   lat_d_arr_3_16 : latch port map ( Q=>d_arr_3_16, D=>nx6490, CLK=>nx10329
   );
   ix6491 : nand02 port map ( Y=>nx6490, A0=>nx9537, A1=>nx10865);
   ix9538 : aoi22 port map ( Y=>nx9537, A0=>d_arr_mul_3_16, A1=>nx10561, B0
      =>d_arr_add_3_16, B1=>nx10717);
   lat_d_arr_3_17 : latch port map ( Q=>d_arr_3_17, D=>nx6500, CLK=>nx10329
   );
   ix6501 : nand02 port map ( Y=>nx6500, A0=>nx9541, A1=>nx10865);
   ix9542 : aoi22 port map ( Y=>nx9541, A0=>d_arr_mul_3_17, A1=>nx10561, B0
      =>d_arr_add_3_17, B1=>nx10717);
   lat_d_arr_3_18 : latch port map ( Q=>d_arr_3_18, D=>nx6510, CLK=>nx10329
   );
   ix6511 : nand02 port map ( Y=>nx6510, A0=>nx9545, A1=>nx10865);
   ix9546 : aoi22 port map ( Y=>nx9545, A0=>d_arr_mul_3_18, A1=>nx10561, B0
      =>d_arr_add_3_18, B1=>nx10717);
   lat_d_arr_3_19 : latch port map ( Q=>d_arr_3_19, D=>nx6520, CLK=>nx10329
   );
   ix6521 : nand02 port map ( Y=>nx6520, A0=>nx9549, A1=>nx10865);
   ix9550 : aoi22 port map ( Y=>nx9549, A0=>d_arr_mul_3_19, A1=>nx10561, B0
      =>d_arr_add_3_19, B1=>nx10717);
   lat_d_arr_3_20 : latch port map ( Q=>d_arr_3_20, D=>nx6530, CLK=>nx10329
   );
   ix6531 : nand02 port map ( Y=>nx6530, A0=>nx9553, A1=>nx10865);
   ix9554 : aoi22 port map ( Y=>nx9553, A0=>d_arr_mul_3_20, A1=>nx10561, B0
      =>d_arr_add_3_20, B1=>nx10717);
   lat_d_arr_3_21 : latch port map ( Q=>d_arr_3_21, D=>nx6540, CLK=>nx10331
   );
   ix6541 : nand02 port map ( Y=>nx6540, A0=>nx9557, A1=>nx10865);
   ix9558 : aoi22 port map ( Y=>nx9557, A0=>d_arr_mul_3_21, A1=>nx10563, B0
      =>d_arr_add_3_21, B1=>nx10717);
   lat_d_arr_3_22 : latch port map ( Q=>d_arr_3_22, D=>nx6550, CLK=>nx10331
   );
   ix6551 : nand02 port map ( Y=>nx6550, A0=>nx9561, A1=>nx10867);
   ix9562 : aoi22 port map ( Y=>nx9561, A0=>d_arr_mul_3_22, A1=>nx10563, B0
      =>d_arr_add_3_22, B1=>nx10717);
   lat_d_arr_3_23 : latch port map ( Q=>d_arr_3_23, D=>nx6560, CLK=>nx10331
   );
   ix6561 : nand02 port map ( Y=>nx6560, A0=>nx9565, A1=>nx10867);
   ix9566 : aoi22 port map ( Y=>nx9565, A0=>d_arr_mul_3_23, A1=>nx10563, B0
      =>d_arr_add_3_23, B1=>nx10719);
   lat_d_arr_3_24 : latch port map ( Q=>d_arr_3_24, D=>nx6570, CLK=>nx10331
   );
   ix6571 : nand02 port map ( Y=>nx6570, A0=>nx9569, A1=>nx10867);
   ix9570 : aoi22 port map ( Y=>nx9569, A0=>d_arr_mul_3_24, A1=>nx10563, B0
      =>d_arr_add_3_24, B1=>nx10719);
   lat_d_arr_3_25 : latch port map ( Q=>d_arr_3_25, D=>nx6580, CLK=>nx10331
   );
   ix6581 : nand02 port map ( Y=>nx6580, A0=>nx9573, A1=>nx10867);
   ix9574 : aoi22 port map ( Y=>nx9573, A0=>d_arr_mul_3_25, A1=>nx10563, B0
      =>d_arr_add_3_25, B1=>nx10719);
   lat_d_arr_3_26 : latch port map ( Q=>d_arr_3_26, D=>nx6590, CLK=>nx10331
   );
   ix6591 : nand02 port map ( Y=>nx6590, A0=>nx9577, A1=>nx10867);
   ix9578 : aoi22 port map ( Y=>nx9577, A0=>d_arr_mul_3_26, A1=>nx10563, B0
      =>d_arr_add_3_26, B1=>nx10719);
   lat_d_arr_3_27 : latch port map ( Q=>d_arr_3_27, D=>nx6600, CLK=>nx10331
   );
   ix6601 : nand02 port map ( Y=>nx6600, A0=>nx9581, A1=>nx10867);
   ix9582 : aoi22 port map ( Y=>nx9581, A0=>d_arr_mul_3_27, A1=>nx10563, B0
      =>d_arr_add_3_27, B1=>nx10719);
   lat_d_arr_3_28 : latch port map ( Q=>d_arr_3_28, D=>nx6610, CLK=>nx10333
   );
   ix6611 : nand02 port map ( Y=>nx6610, A0=>nx9585, A1=>nx10867);
   ix9586 : aoi22 port map ( Y=>nx9585, A0=>d_arr_mul_3_28, A1=>nx10565, B0
      =>d_arr_add_3_28, B1=>nx10719);
   lat_d_arr_3_29 : latch port map ( Q=>d_arr_3_29, D=>nx6620, CLK=>nx10333
   );
   ix6621 : nand02 port map ( Y=>nx6620, A0=>nx9589, A1=>nx9533);
   ix9590 : aoi22 port map ( Y=>nx9589, A0=>d_arr_mul_3_29, A1=>nx10565, B0
      =>d_arr_add_3_29, B1=>nx10719);
   lat_d_arr_3_30 : latch port map ( Q=>d_arr_3_30, D=>nx6630, CLK=>nx10333
   );
   ix6631 : nand02 port map ( Y=>nx6630, A0=>nx9593, A1=>nx9533);
   ix9594 : aoi22 port map ( Y=>nx9593, A0=>d_arr_mul_3_30, A1=>nx10565, B0
      =>d_arr_add_3_30, B1=>nx10721);
   lat_d_arr_3_31 : latch port map ( Q=>d_arr_3_31, D=>nx6640, CLK=>nx10333
   );
   ix6641 : nand02 port map ( Y=>nx6640, A0=>nx9597, A1=>nx9533);
   ix9598 : aoi22 port map ( Y=>nx9597, A0=>d_arr_mul_3_31, A1=>nx10565, B0
      =>d_arr_add_3_31, B1=>nx10721);
   lat_d_arr_2_0 : latch port map ( Q=>d_arr_2_0, D=>nx6652, CLK=>nx10333);
   ix6653 : inv01 port map ( Y=>nx6652, A=>nx9601);
   ix9602 : aoi222 port map ( Y=>nx9601, A0=>d_arr_mux_2_0, A1=>nx11385, B0
      =>d_arr_mul_2_0, B1=>nx10565, C0=>d_arr_add_2_0, C1=>nx10721);
   lat_d_arr_2_1 : latch port map ( Q=>d_arr_2_1, D=>nx6664, CLK=>nx10333);
   ix6665 : inv01 port map ( Y=>nx6664, A=>nx9605);
   ix9606 : aoi222 port map ( Y=>nx9605, A0=>d_arr_mux_2_1, A1=>nx11385, B0
      =>d_arr_mul_2_1, B1=>nx10565, C0=>d_arr_add_2_1, C1=>nx10721);
   lat_d_arr_2_2 : latch port map ( Q=>d_arr_2_2, D=>nx6676, CLK=>nx10333);
   ix6677 : inv01 port map ( Y=>nx6676, A=>nx9609);
   ix9610 : aoi222 port map ( Y=>nx9609, A0=>d_arr_mux_2_2, A1=>nx11385, B0
      =>d_arr_mul_2_2, B1=>nx10565, C0=>d_arr_add_2_2, C1=>nx10721);
   lat_d_arr_2_3 : latch port map ( Q=>d_arr_2_3, D=>nx6688, CLK=>nx10335);
   ix6689 : inv01 port map ( Y=>nx6688, A=>nx9613);
   ix9614 : aoi222 port map ( Y=>nx9613, A0=>d_arr_mux_2_3, A1=>nx11385, B0
      =>d_arr_mul_2_3, B1=>nx10567, C0=>d_arr_add_2_3, C1=>nx10721);
   lat_d_arr_2_4 : latch port map ( Q=>d_arr_2_4, D=>nx6700, CLK=>nx10335);
   ix6701 : inv01 port map ( Y=>nx6700, A=>nx9617);
   ix9618 : aoi222 port map ( Y=>nx9617, A0=>d_arr_mux_2_4, A1=>nx11385, B0
      =>d_arr_mul_2_4, B1=>nx10567, C0=>d_arr_add_2_4, C1=>nx10721);
   lat_d_arr_2_5 : latch port map ( Q=>d_arr_2_5, D=>nx6712, CLK=>nx10335);
   ix6713 : inv01 port map ( Y=>nx6712, A=>nx9621);
   ix9622 : aoi222 port map ( Y=>nx9621, A0=>d_arr_mux_2_5, A1=>nx11385, B0
      =>d_arr_mul_2_5, B1=>nx10567, C0=>d_arr_add_2_5, C1=>nx10723);
   lat_d_arr_2_6 : latch port map ( Q=>d_arr_2_6, D=>nx6724, CLK=>nx10335);
   ix6725 : inv01 port map ( Y=>nx6724, A=>nx9625);
   ix9626 : aoi222 port map ( Y=>nx9625, A0=>d_arr_mux_2_6, A1=>nx11387, B0
      =>d_arr_mul_2_6, B1=>nx10567, C0=>d_arr_add_2_6, C1=>nx10723);
   lat_d_arr_2_7 : latch port map ( Q=>d_arr_2_7, D=>nx6736, CLK=>nx10335);
   ix6737 : inv01 port map ( Y=>nx6736, A=>nx9629);
   ix9630 : aoi222 port map ( Y=>nx9629, A0=>d_arr_mux_2_7, A1=>nx11387, B0
      =>d_arr_mul_2_7, B1=>nx10567, C0=>d_arr_add_2_7, C1=>nx10723);
   lat_d_arr_2_8 : latch port map ( Q=>d_arr_2_8, D=>nx6748, CLK=>nx10335);
   ix6749 : inv01 port map ( Y=>nx6748, A=>nx9633);
   ix9634 : aoi222 port map ( Y=>nx9633, A0=>d_arr_mux_2_8, A1=>nx11387, B0
      =>d_arr_mul_2_8, B1=>nx10567, C0=>d_arr_add_2_8, C1=>nx10723);
   lat_d_arr_2_9 : latch port map ( Q=>d_arr_2_9, D=>nx6760, CLK=>nx10335);
   ix6761 : inv01 port map ( Y=>nx6760, A=>nx9637);
   ix9638 : aoi222 port map ( Y=>nx9637, A0=>d_arr_mux_2_9, A1=>nx11387, B0
      =>d_arr_mul_2_9, B1=>nx10567, C0=>d_arr_add_2_9, C1=>nx10723);
   lat_d_arr_2_10 : latch port map ( Q=>d_arr_2_10, D=>nx6772, CLK=>nx10337
   );
   ix6773 : inv01 port map ( Y=>nx6772, A=>nx9641);
   ix9642 : aoi222 port map ( Y=>nx9641, A0=>d_arr_mux_2_10, A1=>nx11387, B0
      =>d_arr_mul_2_10, B1=>nx10569, C0=>d_arr_add_2_10, C1=>nx10723);
   lat_d_arr_2_11 : latch port map ( Q=>d_arr_2_11, D=>nx6784, CLK=>nx10337
   );
   ix6785 : inv01 port map ( Y=>nx6784, A=>nx9645);
   ix9646 : aoi222 port map ( Y=>nx9645, A0=>d_arr_mux_2_11, A1=>nx11387, B0
      =>d_arr_mul_2_11, B1=>nx10569, C0=>d_arr_add_2_11, C1=>nx10723);
   lat_d_arr_2_12 : latch port map ( Q=>d_arr_2_12, D=>nx6796, CLK=>nx10337
   );
   ix6797 : inv01 port map ( Y=>nx6796, A=>nx9649);
   ix9650 : aoi222 port map ( Y=>nx9649, A0=>d_arr_mux_2_12, A1=>nx11387, B0
      =>d_arr_mul_2_12, B1=>nx10569, C0=>d_arr_add_2_12, C1=>nx10725);
   lat_d_arr_2_13 : latch port map ( Q=>d_arr_2_13, D=>nx6808, CLK=>nx10337
   );
   ix6809 : inv01 port map ( Y=>nx6808, A=>nx9653);
   ix9654 : aoi222 port map ( Y=>nx9653, A0=>d_arr_mux_2_13, A1=>nx11389, B0
      =>d_arr_mul_2_13, B1=>nx10569, C0=>d_arr_add_2_13, C1=>nx10725);
   lat_d_arr_2_14 : latch port map ( Q=>d_arr_2_14, D=>nx6820, CLK=>nx10337
   );
   ix6821 : inv01 port map ( Y=>nx6820, A=>nx9657);
   ix9658 : aoi222 port map ( Y=>nx9657, A0=>d_arr_mux_2_14, A1=>nx11389, B0
      =>d_arr_mul_2_14, B1=>nx10569, C0=>d_arr_add_2_14, C1=>nx10725);
   lat_d_arr_2_15 : latch port map ( Q=>d_arr_2_15, D=>nx6832, CLK=>nx10337
   );
   ix6833 : nand02 port map ( Y=>nx6832, A0=>nx9661, A1=>nx10869);
   ix9662 : aoi22 port map ( Y=>nx9661, A0=>d_arr_mul_2_15, A1=>nx10569, B0
      =>d_arr_add_2_15, B1=>nx10725);
   ix9664 : nand02 port map ( Y=>nx9663, A0=>d_arr_mux_2_31, A1=>nx11389);
   lat_d_arr_2_16 : latch port map ( Q=>d_arr_2_16, D=>nx6842, CLK=>nx10337
   );
   ix6843 : nand02 port map ( Y=>nx6842, A0=>nx9667, A1=>nx10869);
   ix9668 : aoi22 port map ( Y=>nx9667, A0=>d_arr_mul_2_16, A1=>nx10569, B0
      =>d_arr_add_2_16, B1=>nx10725);
   lat_d_arr_2_17 : latch port map ( Q=>d_arr_2_17, D=>nx6852, CLK=>nx10339
   );
   ix6853 : nand02 port map ( Y=>nx6852, A0=>nx9671, A1=>nx10869);
   ix9672 : aoi22 port map ( Y=>nx9671, A0=>d_arr_mul_2_17, A1=>nx10571, B0
      =>d_arr_add_2_17, B1=>nx10725);
   lat_d_arr_2_18 : latch port map ( Q=>d_arr_2_18, D=>nx6862, CLK=>nx10339
   );
   ix6863 : nand02 port map ( Y=>nx6862, A0=>nx9675, A1=>nx10869);
   ix9676 : aoi22 port map ( Y=>nx9675, A0=>d_arr_mul_2_18, A1=>nx10571, B0
      =>d_arr_add_2_18, B1=>nx10725);
   lat_d_arr_2_19 : latch port map ( Q=>d_arr_2_19, D=>nx6872, CLK=>nx10339
   );
   ix6873 : nand02 port map ( Y=>nx6872, A0=>nx9679, A1=>nx10869);
   ix9680 : aoi22 port map ( Y=>nx9679, A0=>d_arr_mul_2_19, A1=>nx10571, B0
      =>d_arr_add_2_19, B1=>nx10727);
   lat_d_arr_2_20 : latch port map ( Q=>d_arr_2_20, D=>nx6882, CLK=>nx10339
   );
   ix6883 : nand02 port map ( Y=>nx6882, A0=>nx9683, A1=>nx10869);
   ix9684 : aoi22 port map ( Y=>nx9683, A0=>d_arr_mul_2_20, A1=>nx10571, B0
      =>d_arr_add_2_20, B1=>nx10727);
   lat_d_arr_2_21 : latch port map ( Q=>d_arr_2_21, D=>nx6892, CLK=>nx10339
   );
   ix6893 : nand02 port map ( Y=>nx6892, A0=>nx9687, A1=>nx10869);
   ix9688 : aoi22 port map ( Y=>nx9687, A0=>d_arr_mul_2_21, A1=>nx10571, B0
      =>d_arr_add_2_21, B1=>nx10727);
   lat_d_arr_2_22 : latch port map ( Q=>d_arr_2_22, D=>nx6902, CLK=>nx10339
   );
   ix6903 : nand02 port map ( Y=>nx6902, A0=>nx9691, A1=>nx10871);
   ix9692 : aoi22 port map ( Y=>nx9691, A0=>d_arr_mul_2_22, A1=>nx10571, B0
      =>d_arr_add_2_22, B1=>nx10727);
   lat_d_arr_2_23 : latch port map ( Q=>d_arr_2_23, D=>nx6912, CLK=>nx10339
   );
   ix6913 : nand02 port map ( Y=>nx6912, A0=>nx9695, A1=>nx10871);
   ix9696 : aoi22 port map ( Y=>nx9695, A0=>d_arr_mul_2_23, A1=>nx10571, B0
      =>d_arr_add_2_23, B1=>nx10727);
   lat_d_arr_2_24 : latch port map ( Q=>d_arr_2_24, D=>nx6922, CLK=>nx10341
   );
   ix6923 : nand02 port map ( Y=>nx6922, A0=>nx9699, A1=>nx10871);
   ix9700 : aoi22 port map ( Y=>nx9699, A0=>d_arr_mul_2_24, A1=>nx10573, B0
      =>d_arr_add_2_24, B1=>nx10727);
   lat_d_arr_2_25 : latch port map ( Q=>d_arr_2_25, D=>nx6932, CLK=>nx10341
   );
   ix6933 : nand02 port map ( Y=>nx6932, A0=>nx9703, A1=>nx10871);
   ix9704 : aoi22 port map ( Y=>nx9703, A0=>d_arr_mul_2_25, A1=>nx10573, B0
      =>d_arr_add_2_25, B1=>nx10727);
   lat_d_arr_2_26 : latch port map ( Q=>d_arr_2_26, D=>nx6942, CLK=>nx10341
   );
   ix6943 : nand02 port map ( Y=>nx6942, A0=>nx9707, A1=>nx10871);
   ix9708 : aoi22 port map ( Y=>nx9707, A0=>d_arr_mul_2_26, A1=>nx10573, B0
      =>d_arr_add_2_26, B1=>nx10729);
   lat_d_arr_2_27 : latch port map ( Q=>d_arr_2_27, D=>nx6952, CLK=>nx10341
   );
   ix6953 : nand02 port map ( Y=>nx6952, A0=>nx9711, A1=>nx10871);
   ix9712 : aoi22 port map ( Y=>nx9711, A0=>d_arr_mul_2_27, A1=>nx10573, B0
      =>d_arr_add_2_27, B1=>nx10729);
   lat_d_arr_2_28 : latch port map ( Q=>d_arr_2_28, D=>nx6962, CLK=>nx10341
   );
   ix6963 : nand02 port map ( Y=>nx6962, A0=>nx9715, A1=>nx10871);
   ix9716 : aoi22 port map ( Y=>nx9715, A0=>d_arr_mul_2_28, A1=>nx10573, B0
      =>d_arr_add_2_28, B1=>nx10729);
   lat_d_arr_2_29 : latch port map ( Q=>d_arr_2_29, D=>nx6972, CLK=>nx10341
   );
   ix6973 : nand02 port map ( Y=>nx6972, A0=>nx9719, A1=>nx9663);
   ix9720 : aoi22 port map ( Y=>nx9719, A0=>d_arr_mul_2_29, A1=>nx10573, B0
      =>d_arr_add_2_29, B1=>nx10729);
   lat_d_arr_2_30 : latch port map ( Q=>d_arr_2_30, D=>nx6982, CLK=>nx10341
   );
   ix6983 : nand02 port map ( Y=>nx6982, A0=>nx9723, A1=>nx9663);
   ix9724 : aoi22 port map ( Y=>nx9723, A0=>d_arr_mul_2_30, A1=>nx10573, B0
      =>d_arr_add_2_30, B1=>nx10729);
   lat_d_arr_2_31 : latch port map ( Q=>d_arr_2_31, D=>nx6992, CLK=>nx10343
   );
   ix6993 : nand02 port map ( Y=>nx6992, A0=>nx9727, A1=>nx9663);
   ix9728 : aoi22 port map ( Y=>nx9727, A0=>d_arr_mul_2_31, A1=>nx10575, B0
      =>d_arr_add_2_31, B1=>nx10729);
   lat_d_arr_1_0 : latch port map ( Q=>d_arr_1_0, D=>nx7036, CLK=>nx10343);
   ix7037 : nand02 port map ( Y=>nx7036, A0=>nx9731, A1=>nx9739);
   ix9732 : aoi222 port map ( Y=>nx9731, A0=>d_arr_mux_1_0, A1=>nx11389, B0
      =>d_arr_merge2_1_0, B1=>nx10805, C0=>d_arr_relu_1_0, C1=>nx10827);
   ix7019 : and02 port map ( Y=>nx7018, A0=>sel_merge2, A1=>nx9734);
   ix9735 : nor04 port map ( Y=>nx9734, A0=>sel_add, A1=>sel_merge1, A2=>
      nx11389, A3=>sel_mul);
   ix7029 : and03 port map ( Y=>nx7028, A0=>nx9734, A1=>sel_relu, A2=>nx9737
   );
   ix9738 : inv01 port map ( Y=>nx9737, A=>sel_merge2);
   ix9740 : aoi222 port map ( Y=>nx9739, A0=>d_arr_mul_1_0, A1=>nx10575, B0
      =>d_arr_add_1_0, B1=>nx10729, C0=>d_arr_merge1_1_0, C1=>nx10783);
   ix7003 : nor04 port map ( Y=>nx7002, A0=>nx11389, A1=>sel_mul, A2=>nx9742, 
      A3=>sel_add);
   ix9743 : inv01 port map ( Y=>nx9742, A=>sel_merge1);
   lat_d_arr_1_1 : latch port map ( Q=>d_arr_1_1, D=>nx7060, CLK=>nx10343);
   ix7061 : nand02 port map ( Y=>nx7060, A0=>nx9746, A1=>nx9748);
   ix9747 : aoi222 port map ( Y=>nx9746, A0=>d_arr_mux_1_1, A1=>nx11389, B0
      =>d_arr_merge2_1_1, B1=>nx10805, C0=>d_arr_relu_1_1, C1=>nx10827);
   ix9749 : aoi222 port map ( Y=>nx9748, A0=>d_arr_mul_1_1, A1=>nx10575, B0
      =>d_arr_add_1_1, B1=>nx10731, C0=>d_arr_merge1_1_1, C1=>nx10783);
   lat_d_arr_1_2 : latch port map ( Q=>d_arr_1_2, D=>nx7084, CLK=>nx10343);
   ix7085 : nand02 port map ( Y=>nx7084, A0=>nx9752, A1=>nx9754);
   ix9753 : aoi222 port map ( Y=>nx9752, A0=>d_arr_mux_1_2, A1=>nx11391, B0
      =>d_arr_merge2_1_2, B1=>nx10805, C0=>d_arr_relu_1_2, C1=>nx10827);
   ix9755 : aoi222 port map ( Y=>nx9754, A0=>d_arr_mul_1_2, A1=>nx10575, B0
      =>d_arr_add_1_2, B1=>nx10731, C0=>d_arr_merge1_1_2, C1=>nx10783);
   lat_d_arr_1_3 : latch port map ( Q=>d_arr_1_3, D=>nx7108, CLK=>nx10343);
   ix7109 : nand02 port map ( Y=>nx7108, A0=>nx9758, A1=>nx9760);
   ix9759 : aoi222 port map ( Y=>nx9758, A0=>d_arr_mux_1_3, A1=>nx11391, B0
      =>d_arr_merge2_1_3, B1=>nx10805, C0=>d_arr_relu_1_3, C1=>nx10827);
   ix9761 : aoi222 port map ( Y=>nx9760, A0=>d_arr_mul_1_3, A1=>nx10575, B0
      =>d_arr_add_1_3, B1=>nx10731, C0=>d_arr_merge1_1_3, C1=>nx10783);
   lat_d_arr_1_4 : latch port map ( Q=>d_arr_1_4, D=>nx7132, CLK=>nx10343);
   ix7133 : nand02 port map ( Y=>nx7132, A0=>nx9764, A1=>nx9766);
   ix9765 : aoi222 port map ( Y=>nx9764, A0=>d_arr_mux_1_4, A1=>nx11391, B0
      =>d_arr_merge2_1_4, B1=>nx10805, C0=>d_arr_relu_1_4, C1=>nx10827);
   ix9767 : aoi222 port map ( Y=>nx9766, A0=>d_arr_mul_1_4, A1=>nx10575, B0
      =>d_arr_add_1_4, B1=>nx10731, C0=>d_arr_merge1_1_4, C1=>nx10783);
   lat_d_arr_1_5 : latch port map ( Q=>d_arr_1_5, D=>nx7156, CLK=>nx10343);
   ix7157 : nand02 port map ( Y=>nx7156, A0=>nx9770, A1=>nx9772);
   ix9771 : aoi222 port map ( Y=>nx9770, A0=>d_arr_mux_1_5, A1=>nx11391, B0
      =>d_arr_merge2_1_5, B1=>nx10805, C0=>d_arr_relu_1_5, C1=>nx10827);
   ix9773 : aoi222 port map ( Y=>nx9772, A0=>d_arr_mul_1_5, A1=>nx10575, B0
      =>d_arr_add_1_5, B1=>nx10731, C0=>d_arr_merge1_1_5, C1=>nx10783);
   lat_d_arr_1_6 : latch port map ( Q=>d_arr_1_6, D=>nx7180, CLK=>nx10345);
   ix7181 : nand02 port map ( Y=>nx7180, A0=>nx9776, A1=>nx9778);
   ix9777 : aoi222 port map ( Y=>nx9776, A0=>d_arr_mux_1_6, A1=>nx11391, B0
      =>d_arr_merge2_1_6, B1=>nx10805, C0=>d_arr_relu_1_6, C1=>nx10827);
   ix9779 : aoi222 port map ( Y=>nx9778, A0=>d_arr_mul_1_6, A1=>nx10577, B0
      =>d_arr_add_1_6, B1=>nx10731, C0=>d_arr_merge1_1_6, C1=>nx10783);
   lat_d_arr_1_7 : latch port map ( Q=>d_arr_1_7, D=>nx7204, CLK=>nx10345);
   ix7205 : nand02 port map ( Y=>nx7204, A0=>nx9782, A1=>nx9784);
   ix9783 : aoi222 port map ( Y=>nx9782, A0=>d_arr_mux_1_7, A1=>nx11391, B0
      =>d_arr_merge2_1_7, B1=>nx10807, C0=>d_arr_relu_1_7, C1=>nx10829);
   ix9785 : aoi222 port map ( Y=>nx9784, A0=>d_arr_mul_1_7, A1=>nx10577, B0
      =>d_arr_add_1_7, B1=>nx10731, C0=>d_arr_merge1_1_7, C1=>nx10785);
   lat_d_arr_1_8 : latch port map ( Q=>d_arr_1_8, D=>nx7228, CLK=>nx10345);
   ix7229 : nand02 port map ( Y=>nx7228, A0=>nx9788, A1=>nx9790);
   ix9789 : aoi222 port map ( Y=>nx9788, A0=>d_arr_mux_1_8, A1=>nx11391, B0
      =>d_arr_merge2_1_8, B1=>nx10807, C0=>d_arr_relu_1_8, C1=>nx10829);
   ix9791 : aoi222 port map ( Y=>nx9790, A0=>d_arr_mul_1_8, A1=>nx10577, B0
      =>d_arr_add_1_8, B1=>nx10733, C0=>d_arr_merge1_1_8, C1=>nx10785);
   lat_d_arr_1_9 : latch port map ( Q=>d_arr_1_9, D=>nx7252, CLK=>nx10345);
   ix7253 : nand02 port map ( Y=>nx7252, A0=>nx9794, A1=>nx9796);
   ix9795 : aoi222 port map ( Y=>nx9794, A0=>d_arr_mux_1_9, A1=>nx11393, B0
      =>d_arr_merge2_1_9, B1=>nx10807, C0=>d_arr_relu_1_9, C1=>nx10829);
   ix9797 : aoi222 port map ( Y=>nx9796, A0=>d_arr_mul_1_9, A1=>nx10577, B0
      =>d_arr_add_1_9, B1=>nx10733, C0=>d_arr_merge1_1_9, C1=>nx10785);
   lat_d_arr_1_10 : latch port map ( Q=>d_arr_1_10, D=>nx7276, CLK=>nx10345
   );
   ix7277 : nand02 port map ( Y=>nx7276, A0=>nx9800, A1=>nx9802);
   ix9801 : aoi222 port map ( Y=>nx9800, A0=>d_arr_mux_1_10, A1=>nx11393, B0
      =>d_arr_merge2_1_10, B1=>nx10807, C0=>d_arr_relu_1_10, C1=>nx10829);
   ix9803 : aoi222 port map ( Y=>nx9802, A0=>d_arr_mul_1_10, A1=>nx10577, B0
      =>d_arr_add_1_10, B1=>nx10733, C0=>d_arr_merge1_1_10, C1=>nx10785);
   lat_d_arr_1_11 : latch port map ( Q=>d_arr_1_11, D=>nx7300, CLK=>nx10345
   );
   ix7301 : nand02 port map ( Y=>nx7300, A0=>nx9806, A1=>nx9808);
   ix9807 : aoi222 port map ( Y=>nx9806, A0=>d_arr_mux_1_11, A1=>nx11393, B0
      =>d_arr_merge2_1_11, B1=>nx10807, C0=>d_arr_relu_1_11, C1=>nx10829);
   ix9809 : aoi222 port map ( Y=>nx9808, A0=>d_arr_mul_1_11, A1=>nx10577, B0
      =>d_arr_add_1_11, B1=>nx10733, C0=>d_arr_merge1_1_11, C1=>nx10785);
   lat_d_arr_1_12 : latch port map ( Q=>d_arr_1_12, D=>nx7324, CLK=>nx10345
   );
   ix7325 : nand02 port map ( Y=>nx7324, A0=>nx9812, A1=>nx9814);
   ix9813 : aoi222 port map ( Y=>nx9812, A0=>d_arr_mux_1_12, A1=>nx11393, B0
      =>d_arr_merge2_1_12, B1=>nx10807, C0=>d_arr_relu_1_12, C1=>nx10829);
   ix9815 : aoi222 port map ( Y=>nx9814, A0=>d_arr_mul_1_12, A1=>nx10577, B0
      =>d_arr_add_1_12, B1=>nx10733, C0=>d_arr_merge1_1_12, C1=>nx10785);
   lat_d_arr_1_13 : latch port map ( Q=>d_arr_1_13, D=>nx7348, CLK=>nx10347
   );
   ix7349 : nand02 port map ( Y=>nx7348, A0=>nx9818, A1=>nx9820);
   ix9819 : aoi222 port map ( Y=>nx9818, A0=>d_arr_mux_1_13, A1=>nx11393, B0
      =>d_arr_merge2_1_13, B1=>nx10807, C0=>d_arr_relu_1_13, C1=>nx10829);
   ix9821 : aoi222 port map ( Y=>nx9820, A0=>d_arr_mul_1_13, A1=>nx10579, B0
      =>d_arr_add_1_13, B1=>nx10733, C0=>d_arr_merge1_1_13, C1=>nx10785);
   lat_d_arr_1_14 : latch port map ( Q=>d_arr_1_14, D=>nx7372, CLK=>nx10347
   );
   ix7373 : nand02 port map ( Y=>nx7372, A0=>nx9824, A1=>nx9826);
   ix9825 : aoi222 port map ( Y=>nx9824, A0=>d_arr_mux_1_14, A1=>nx11393, B0
      =>d_arr_merge2_1_14, B1=>nx10809, C0=>d_arr_relu_1_14, C1=>nx10831);
   ix9827 : aoi222 port map ( Y=>nx9826, A0=>d_arr_mul_1_14, A1=>nx10579, B0
      =>d_arr_add_1_14, B1=>nx10733, C0=>d_arr_merge1_1_14, C1=>nx10787);
   lat_d_arr_1_15 : latch port map ( Q=>d_arr_1_15, D=>nx7392, CLK=>nx10347
   );
   ix7393 : nand03 port map ( Y=>nx7392, A0=>nx9830, A1=>nx10873, A2=>nx9834
   );
   ix9831 : nand02 port map ( Y=>nx9830, A0=>d_arr_merge2_1_15, A1=>nx10809
   );
   ix9833 : nand02 port map ( Y=>nx9832, A0=>d_arr_mux_1_31, A1=>nx11393);
   ix9835 : aoi222 port map ( Y=>nx9834, A0=>d_arr_mul_1_15, A1=>nx10579, B0
      =>d_arr_add_1_15, B1=>nx10735, C0=>d_arr_merge1_1_15, C1=>nx10787);
   lat_d_arr_1_16 : latch port map ( Q=>d_arr_1_16, D=>nx7414, CLK=>nx10347
   );
   ix7415 : nand03 port map ( Y=>nx7414, A0=>nx9838, A1=>nx10873, A2=>nx9840
   );
   ix9839 : aoi22 port map ( Y=>nx9838, A0=>d_arr_merge2_1_16, A1=>nx10809, 
      B0=>d_arr_relu_1_16, B1=>nx10831);
   ix9841 : aoi222 port map ( Y=>nx9840, A0=>d_arr_mul_1_16, A1=>nx10579, B0
      =>d_arr_add_1_16, B1=>nx10735, C0=>d_arr_merge1_1_16, C1=>nx10787);
   lat_d_arr_1_17 : latch port map ( Q=>d_arr_1_17, D=>nx7436, CLK=>nx10347
   );
   ix7437 : nand03 port map ( Y=>nx7436, A0=>nx9844, A1=>nx10873, A2=>nx9846
   );
   ix9845 : aoi22 port map ( Y=>nx9844, A0=>d_arr_merge2_1_17, A1=>nx10809, 
      B0=>d_arr_relu_1_17, B1=>nx10831);
   ix9847 : aoi222 port map ( Y=>nx9846, A0=>d_arr_mul_1_17, A1=>nx10579, B0
      =>d_arr_add_1_17, B1=>nx10735, C0=>d_arr_merge1_1_17, C1=>nx10787);
   lat_d_arr_1_18 : latch port map ( Q=>d_arr_1_18, D=>nx7458, CLK=>nx10347
   );
   ix7459 : nand03 port map ( Y=>nx7458, A0=>nx9850, A1=>nx10873, A2=>nx9852
   );
   ix9851 : aoi22 port map ( Y=>nx9850, A0=>d_arr_merge2_1_18, A1=>nx10809, 
      B0=>d_arr_relu_1_18, B1=>nx10831);
   ix9853 : aoi222 port map ( Y=>nx9852, A0=>d_arr_mul_1_18, A1=>nx10579, B0
      =>d_arr_add_1_18, B1=>nx10735, C0=>d_arr_merge1_1_18, C1=>nx10787);
   lat_d_arr_1_19 : latch port map ( Q=>d_arr_1_19, D=>nx7480, CLK=>nx10347
   );
   ix7481 : nand03 port map ( Y=>nx7480, A0=>nx9856, A1=>nx10873, A2=>nx9858
   );
   ix9857 : aoi22 port map ( Y=>nx9856, A0=>d_arr_merge2_1_19, A1=>nx10809, 
      B0=>d_arr_relu_1_19, B1=>nx10831);
   ix9859 : aoi222 port map ( Y=>nx9858, A0=>d_arr_mul_1_19, A1=>nx10579, B0
      =>d_arr_add_1_19, B1=>nx10735, C0=>d_arr_merge1_1_19, C1=>nx10787);
   lat_d_arr_1_20 : latch port map ( Q=>d_arr_1_20, D=>nx7502, CLK=>nx10349
   );
   ix7503 : nand03 port map ( Y=>nx7502, A0=>nx9862, A1=>nx10873, A2=>nx9864
   );
   ix9863 : aoi22 port map ( Y=>nx9862, A0=>d_arr_merge2_1_20, A1=>nx10809, 
      B0=>d_arr_relu_1_20, B1=>nx10831);
   ix9865 : aoi222 port map ( Y=>nx9864, A0=>d_arr_mul_1_20, A1=>nx10581, B0
      =>d_arr_add_1_20, B1=>nx10735, C0=>d_arr_merge1_1_20, C1=>nx10787);
   lat_d_arr_1_21 : latch port map ( Q=>d_arr_1_21, D=>nx7524, CLK=>nx10349
   );
   ix7525 : nand03 port map ( Y=>nx7524, A0=>nx9868, A1=>nx10873, A2=>nx9870
   );
   ix9869 : aoi22 port map ( Y=>nx9868, A0=>d_arr_merge2_1_21, A1=>nx10811, 
      B0=>d_arr_relu_1_21, B1=>nx10831);
   ix9871 : aoi222 port map ( Y=>nx9870, A0=>d_arr_mul_1_21, A1=>nx10581, B0
      =>d_arr_add_1_21, B1=>nx10735, C0=>d_arr_merge1_1_21, C1=>nx10789);
   lat_d_arr_1_22 : latch port map ( Q=>d_arr_1_22, D=>nx7546, CLK=>nx10349
   );
   ix7547 : nand03 port map ( Y=>nx7546, A0=>nx9874, A1=>nx10875, A2=>nx9876
   );
   ix9875 : aoi22 port map ( Y=>nx9874, A0=>d_arr_merge2_1_22, A1=>nx10811, 
      B0=>d_arr_relu_1_22, B1=>nx10833);
   ix9877 : aoi222 port map ( Y=>nx9876, A0=>d_arr_mul_1_22, A1=>nx10581, B0
      =>d_arr_add_1_22, B1=>nx10737, C0=>d_arr_merge1_1_22, C1=>nx10789);
   lat_d_arr_1_23 : latch port map ( Q=>d_arr_1_23, D=>nx7568, CLK=>nx10349
   );
   ix7569 : nand03 port map ( Y=>nx7568, A0=>nx9880, A1=>nx10875, A2=>nx9882
   );
   ix9881 : aoi22 port map ( Y=>nx9880, A0=>d_arr_merge2_1_23, A1=>nx10811, 
      B0=>d_arr_relu_1_23, B1=>nx10833);
   ix9883 : aoi222 port map ( Y=>nx9882, A0=>d_arr_mul_1_23, A1=>nx10581, B0
      =>d_arr_add_1_23, B1=>nx10737, C0=>d_arr_merge1_1_23, C1=>nx10789);
   lat_d_arr_1_24 : latch port map ( Q=>d_arr_1_24, D=>nx7590, CLK=>nx10349
   );
   ix7591 : nand03 port map ( Y=>nx7590, A0=>nx9886, A1=>nx10875, A2=>nx9888
   );
   ix9887 : aoi22 port map ( Y=>nx9886, A0=>d_arr_merge2_1_24, A1=>nx10811, 
      B0=>d_arr_relu_1_24, B1=>nx10833);
   ix9889 : aoi222 port map ( Y=>nx9888, A0=>d_arr_mul_1_24, A1=>nx10581, B0
      =>d_arr_add_1_24, B1=>nx10737, C0=>d_arr_merge1_1_24, C1=>nx10789);
   lat_d_arr_1_25 : latch port map ( Q=>d_arr_1_25, D=>nx7612, CLK=>nx10349
   );
   ix7613 : nand03 port map ( Y=>nx7612, A0=>nx9892, A1=>nx10875, A2=>nx9894
   );
   ix9893 : aoi22 port map ( Y=>nx9892, A0=>d_arr_merge2_1_25, A1=>nx10811, 
      B0=>d_arr_relu_1_25, B1=>nx10833);
   ix9895 : aoi222 port map ( Y=>nx9894, A0=>d_arr_mul_1_25, A1=>nx10581, B0
      =>d_arr_add_1_25, B1=>nx10737, C0=>d_arr_merge1_1_25, C1=>nx10789);
   lat_d_arr_1_26 : latch port map ( Q=>d_arr_1_26, D=>nx7634, CLK=>nx10349
   );
   ix7635 : nand03 port map ( Y=>nx7634, A0=>nx9898, A1=>nx10875, A2=>nx9900
   );
   ix9899 : aoi22 port map ( Y=>nx9898, A0=>d_arr_merge2_1_26, A1=>nx10811, 
      B0=>d_arr_relu_1_26, B1=>nx10833);
   ix9901 : aoi222 port map ( Y=>nx9900, A0=>d_arr_mul_1_26, A1=>nx10581, B0
      =>d_arr_add_1_26, B1=>nx10737, C0=>d_arr_merge1_1_26, C1=>nx10789);
   lat_d_arr_1_27 : latch port map ( Q=>d_arr_1_27, D=>nx7656, CLK=>nx10351
   );
   ix7657 : nand03 port map ( Y=>nx7656, A0=>nx9904, A1=>nx10875, A2=>nx9906
   );
   ix9905 : aoi22 port map ( Y=>nx9904, A0=>d_arr_merge2_1_27, A1=>nx10811, 
      B0=>d_arr_relu_1_27, B1=>nx10833);
   ix9907 : aoi222 port map ( Y=>nx9906, A0=>d_arr_mul_1_27, A1=>nx10583, B0
      =>d_arr_add_1_27, B1=>nx10737, C0=>d_arr_merge1_1_27, C1=>nx10789);
   lat_d_arr_1_28 : latch port map ( Q=>d_arr_1_28, D=>nx7678, CLK=>nx10351
   );
   ix7679 : nand03 port map ( Y=>nx7678, A0=>nx9910, A1=>nx10875, A2=>nx9912
   );
   ix9911 : aoi22 port map ( Y=>nx9910, A0=>d_arr_merge2_1_28, A1=>nx10813, 
      B0=>d_arr_relu_1_28, B1=>nx10833);
   ix9913 : aoi222 port map ( Y=>nx9912, A0=>d_arr_mul_1_28, A1=>nx10583, B0
      =>d_arr_add_1_28, B1=>nx10737, C0=>d_arr_merge1_1_28, C1=>nx10791);
   lat_d_arr_1_29 : latch port map ( Q=>d_arr_1_29, D=>nx7700, CLK=>nx10351
   );
   ix7701 : nand03 port map ( Y=>nx7700, A0=>nx9916, A1=>nx9832, A2=>nx9918
   );
   ix9917 : aoi22 port map ( Y=>nx9916, A0=>d_arr_merge2_1_29, A1=>nx10813, 
      B0=>d_arr_relu_1_29, B1=>nx10835);
   ix9919 : aoi222 port map ( Y=>nx9918, A0=>d_arr_mul_1_29, A1=>nx10583, B0
      =>d_arr_add_1_29, B1=>nx10739, C0=>d_arr_merge1_1_29, C1=>nx10791);
   lat_d_arr_1_30 : latch port map ( Q=>d_arr_1_30, D=>nx7722, CLK=>nx10351
   );
   ix7723 : nand03 port map ( Y=>nx7722, A0=>nx9922, A1=>nx9832, A2=>nx9924
   );
   ix9923 : aoi22 port map ( Y=>nx9922, A0=>d_arr_merge2_1_30, A1=>nx10813, 
      B0=>d_arr_relu_1_30, B1=>nx10835);
   ix9925 : aoi222 port map ( Y=>nx9924, A0=>d_arr_mul_1_30, A1=>nx10583, B0
      =>d_arr_add_1_30, B1=>nx10739, C0=>d_arr_merge1_1_30, C1=>nx10791);
   lat_d_arr_1_31 : latch port map ( Q=>d_arr_1_31, D=>nx7744, CLK=>nx10351
   );
   ix7745 : nand03 port map ( Y=>nx7744, A0=>nx9928, A1=>nx9832, A2=>nx9930
   );
   ix9929 : aoi22 port map ( Y=>nx9928, A0=>d_arr_merge2_1_31, A1=>nx10813, 
      B0=>d_arr_relu_1_31, B1=>nx10835);
   ix9931 : aoi222 port map ( Y=>nx9930, A0=>d_arr_mul_1_31, A1=>nx10583, B0
      =>d_arr_add_1_31, B1=>nx10739, C0=>d_arr_merge1_1_31, C1=>nx10791);
   lat_d_arr_0_0 : latch port map ( Q=>d_arr_0_0, D=>nx7768, CLK=>nx10351);
   ix7769 : nand02 port map ( Y=>nx7768, A0=>nx9934, A1=>nx9936);
   ix9935 : aoi222 port map ( Y=>nx9934, A0=>d_arr_mux_0_0, A1=>nx11395, B0
      =>d_arr_merge2_0_0, B1=>nx10813, C0=>d_arr_relu_0_0, C1=>nx10835);
   ix9937 : aoi222 port map ( Y=>nx9936, A0=>d_arr_mul_0_0, A1=>nx10583, B0
      =>d_arr_add_0_0, B1=>nx10739, C0=>d_arr_merge1_0_0, C1=>nx10791);
   lat_d_arr_0_1 : latch port map ( Q=>d_arr_0_1, D=>nx7792, CLK=>nx10351);
   ix7793 : nand02 port map ( Y=>nx7792, A0=>nx9940, A1=>nx9942);
   ix9941 : aoi222 port map ( Y=>nx9940, A0=>d_arr_mux_0_1, A1=>nx11395, B0
      =>d_arr_merge2_0_1, B1=>nx10813, C0=>d_arr_relu_0_1, C1=>nx10835);
   ix9943 : aoi222 port map ( Y=>nx9942, A0=>d_arr_mul_0_1, A1=>nx10583, B0
      =>d_arr_add_0_1, B1=>nx10739, C0=>d_arr_merge1_0_1, C1=>nx10791);
   lat_d_arr_0_2 : latch port map ( Q=>d_arr_0_2, D=>nx7816, CLK=>nx10353);
   ix7817 : nand02 port map ( Y=>nx7816, A0=>nx9946, A1=>nx9948);
   ix9947 : aoi222 port map ( Y=>nx9946, A0=>d_arr_mux_0_2, A1=>nx11395, B0
      =>d_arr_merge2_0_2, B1=>nx10813, C0=>d_arr_relu_0_2, C1=>nx10835);
   ix9949 : aoi222 port map ( Y=>nx9948, A0=>d_arr_mul_0_2, A1=>nx10585, B0
      =>d_arr_add_0_2, B1=>nx10739, C0=>d_arr_merge1_0_2, C1=>nx10791);
   lat_d_arr_0_3 : latch port map ( Q=>d_arr_0_3, D=>nx7840, CLK=>nx10353);
   ix7841 : nand02 port map ( Y=>nx7840, A0=>nx9952, A1=>nx9954);
   ix9953 : aoi222 port map ( Y=>nx9952, A0=>d_arr_mux_0_3, A1=>nx11395, B0
      =>d_arr_merge2_0_3, B1=>nx10815, C0=>d_arr_relu_0_3, C1=>nx10835);
   ix9955 : aoi222 port map ( Y=>nx9954, A0=>d_arr_mul_0_3, A1=>nx10585, B0
      =>d_arr_add_0_3, B1=>nx10739, C0=>d_arr_merge1_0_3, C1=>nx10793);
   lat_d_arr_0_4 : latch port map ( Q=>d_arr_0_4, D=>nx7864, CLK=>nx10353);
   ix7865 : nand02 port map ( Y=>nx7864, A0=>nx9958, A1=>nx9960);
   ix9959 : aoi222 port map ( Y=>nx9958, A0=>d_arr_mux_0_4, A1=>nx11395, B0
      =>d_arr_merge2_0_4, B1=>nx10815, C0=>d_arr_relu_0_4, C1=>nx10837);
   ix9961 : aoi222 port map ( Y=>nx9960, A0=>d_arr_mul_0_4, A1=>nx10585, B0
      =>d_arr_add_0_4, B1=>nx10741, C0=>d_arr_merge1_0_4, C1=>nx10793);
   lat_d_arr_0_5 : latch port map ( Q=>d_arr_0_5, D=>nx7888, CLK=>nx10353);
   ix7889 : nand02 port map ( Y=>nx7888, A0=>nx9964, A1=>nx9966);
   ix9965 : aoi222 port map ( Y=>nx9964, A0=>d_arr_mux_0_5, A1=>nx11395, B0
      =>d_arr_merge2_0_5, B1=>nx10815, C0=>d_arr_relu_0_5, C1=>nx10837);
   ix9967 : aoi222 port map ( Y=>nx9966, A0=>d_arr_mul_0_5, A1=>nx10585, B0
      =>d_arr_add_0_5, B1=>nx10741, C0=>d_arr_merge1_0_5, C1=>nx10793);
   lat_d_arr_0_6 : latch port map ( Q=>d_arr_0_6, D=>nx7912, CLK=>nx10353);
   ix7913 : nand02 port map ( Y=>nx7912, A0=>nx9970, A1=>nx9972);
   ix9971 : aoi222 port map ( Y=>nx9970, A0=>d_arr_mux_0_6, A1=>nx11395, B0
      =>d_arr_merge2_0_6, B1=>nx10815, C0=>d_arr_relu_0_6, C1=>nx10837);
   ix9973 : aoi222 port map ( Y=>nx9972, A0=>d_arr_mul_0_6, A1=>nx10585, B0
      =>d_arr_add_0_6, B1=>nx10741, C0=>d_arr_merge1_0_6, C1=>nx10793);
   lat_d_arr_0_7 : latch port map ( Q=>d_arr_0_7, D=>nx7936, CLK=>nx10353);
   ix7937 : nand02 port map ( Y=>nx7936, A0=>nx9976, A1=>nx9978);
   ix9977 : aoi222 port map ( Y=>nx9976, A0=>d_arr_mux_0_7, A1=>nx11397, B0
      =>d_arr_merge2_0_7, B1=>nx10815, C0=>d_arr_relu_0_7, C1=>nx10837);
   ix9979 : aoi222 port map ( Y=>nx9978, A0=>d_arr_mul_0_7, A1=>nx10585, B0
      =>d_arr_add_0_7, B1=>nx10741, C0=>d_arr_merge1_0_7, C1=>nx10793);
   lat_d_arr_0_8 : latch port map ( Q=>d_arr_0_8, D=>nx7960, CLK=>nx10353);
   ix7961 : nand02 port map ( Y=>nx7960, A0=>nx9982, A1=>nx9984);
   ix9983 : aoi222 port map ( Y=>nx9982, A0=>d_arr_mux_0_8, A1=>nx11397, B0
      =>d_arr_merge2_0_8, B1=>nx10815, C0=>d_arr_relu_0_8, C1=>nx10837);
   ix9985 : aoi222 port map ( Y=>nx9984, A0=>d_arr_mul_0_8, A1=>nx10585, B0
      =>d_arr_add_0_8, B1=>nx10741, C0=>d_arr_merge1_0_8, C1=>nx10793);
   lat_d_arr_0_9 : latch port map ( Q=>d_arr_0_9, D=>nx7984, CLK=>nx10355);
   ix7985 : nand02 port map ( Y=>nx7984, A0=>nx9988, A1=>nx9990);
   ix9989 : aoi222 port map ( Y=>nx9988, A0=>d_arr_mux_0_9, A1=>nx11397, B0
      =>d_arr_merge2_0_9, B1=>nx10815, C0=>d_arr_relu_0_9, C1=>nx10837);
   ix9991 : aoi222 port map ( Y=>nx9990, A0=>d_arr_mul_0_9, A1=>nx10587, B0
      =>d_arr_add_0_9, B1=>nx10741, C0=>d_arr_merge1_0_9, C1=>nx10793);
   lat_d_arr_0_10 : latch port map ( Q=>d_arr_0_10, D=>nx8008, CLK=>nx10355
   );
   ix8009 : nand02 port map ( Y=>nx8008, A0=>nx9994, A1=>nx9996);
   ix9995 : aoi222 port map ( Y=>nx9994, A0=>d_arr_mux_0_10, A1=>nx11397, B0
      =>d_arr_merge2_0_10, B1=>nx10817, C0=>d_arr_relu_0_10, C1=>nx10837);
   ix9997 : aoi222 port map ( Y=>nx9996, A0=>d_arr_mul_0_10, A1=>nx10587, B0
      =>d_arr_add_0_10, B1=>nx10741, C0=>d_arr_merge1_0_10, C1=>nx10795);
   lat_d_arr_0_11 : latch port map ( Q=>d_arr_0_11, D=>nx8032, CLK=>nx10355
   );
   ix8033 : nand02 port map ( Y=>nx8032, A0=>nx10000, A1=>nx10002);
   ix10001 : aoi222 port map ( Y=>nx10000, A0=>d_arr_mux_0_11, A1=>nx11397, 
      B0=>d_arr_merge2_0_11, B1=>nx10817, C0=>d_arr_relu_0_11, C1=>nx10839);
   ix10003 : aoi222 port map ( Y=>nx10002, A0=>d_arr_mul_0_11, A1=>nx10587, 
      B0=>d_arr_add_0_11, B1=>nx10743, C0=>d_arr_merge1_0_11, C1=>nx10795);
   lat_d_arr_0_12 : latch port map ( Q=>d_arr_0_12, D=>nx8056, CLK=>nx10355
   );
   ix8057 : nand02 port map ( Y=>nx8056, A0=>nx10006, A1=>nx10008);
   ix10007 : aoi222 port map ( Y=>nx10006, A0=>d_arr_mux_0_12, A1=>nx11397, 
      B0=>d_arr_merge2_0_12, B1=>nx10817, C0=>d_arr_relu_0_12, C1=>nx10839);
   ix10009 : aoi222 port map ( Y=>nx10008, A0=>d_arr_mul_0_12, A1=>nx10587, 
      B0=>d_arr_add_0_12, B1=>nx10743, C0=>d_arr_merge1_0_12, C1=>nx10795);
   lat_d_arr_0_13 : latch port map ( Q=>d_arr_0_13, D=>nx8080, CLK=>nx10355
   );
   ix8081 : nand02 port map ( Y=>nx8080, A0=>nx10012, A1=>nx10014);
   ix10013 : aoi222 port map ( Y=>nx10012, A0=>d_arr_mux_0_13, A1=>nx11397, 
      B0=>d_arr_merge2_0_13, B1=>nx10817, C0=>d_arr_relu_0_13, C1=>nx10839);
   ix10015 : aoi222 port map ( Y=>nx10014, A0=>d_arr_mul_0_13, A1=>nx10587, 
      B0=>d_arr_add_0_13, B1=>nx10743, C0=>d_arr_merge1_0_13, C1=>nx10795);
   lat_d_arr_0_14 : latch port map ( Q=>d_arr_0_14, D=>nx8104, CLK=>nx10355
   );
   ix8105 : nand02 port map ( Y=>nx8104, A0=>nx10018, A1=>nx10020);
   ix10019 : aoi222 port map ( Y=>nx10018, A0=>d_arr_mux_0_14, A1=>nx11399, 
      B0=>d_arr_merge2_0_14, B1=>nx10817, C0=>d_arr_relu_0_14, C1=>nx10839);
   ix10021 : aoi222 port map ( Y=>nx10020, A0=>d_arr_mul_0_14, A1=>nx10587, 
      B0=>d_arr_add_0_14, B1=>nx10743, C0=>d_arr_merge1_0_14, C1=>nx10795);
   lat_d_arr_0_15 : latch port map ( Q=>d_arr_0_15, D=>nx8124, CLK=>nx10355
   );
   ix8125 : nand03 port map ( Y=>nx8124, A0=>nx10024, A1=>nx10877, A2=>
      nx10028);
   ix10025 : nand02 port map ( Y=>nx10024, A0=>d_arr_merge2_0_15, A1=>
      nx10817);
   ix10027 : nand02 port map ( Y=>nx10026, A0=>d_arr_mux_0_31, A1=>nx11399);
   ix10029 : aoi222 port map ( Y=>nx10028, A0=>d_arr_mul_0_15, A1=>nx10587, 
      B0=>d_arr_add_0_15, B1=>nx10743, C0=>d_arr_merge1_0_15, C1=>nx10795);
   lat_d_arr_0_16 : latch port map ( Q=>d_arr_0_16, D=>nx8146, CLK=>nx10357
   );
   ix8147 : nand03 port map ( Y=>nx8146, A0=>nx10032, A1=>nx10877, A2=>
      nx10034);
   ix10033 : aoi22 port map ( Y=>nx10032, A0=>d_arr_merge2_0_16, A1=>nx10817, 
      B0=>d_arr_relu_0_16, B1=>nx10839);
   ix10035 : aoi222 port map ( Y=>nx10034, A0=>d_arr_mul_0_16, A1=>nx10589, 
      B0=>d_arr_add_0_16, B1=>nx10743, C0=>d_arr_merge1_0_16, C1=>nx10795);
   lat_d_arr_0_17 : latch port map ( Q=>d_arr_0_17, D=>nx8168, CLK=>nx10357
   );
   ix8169 : nand03 port map ( Y=>nx8168, A0=>nx10038, A1=>nx10877, A2=>
      nx10040);
   ix10039 : aoi22 port map ( Y=>nx10038, A0=>d_arr_merge2_0_17, A1=>nx10819, 
      B0=>d_arr_relu_0_17, B1=>nx10839);
   ix10041 : aoi222 port map ( Y=>nx10040, A0=>d_arr_mul_0_17, A1=>nx10589, 
      B0=>d_arr_add_0_17, B1=>nx10743, C0=>d_arr_merge1_0_17, C1=>nx10797);
   lat_d_arr_0_18 : latch port map ( Q=>d_arr_0_18, D=>nx8190, CLK=>nx10357
   );
   ix8191 : nand03 port map ( Y=>nx8190, A0=>nx10044, A1=>nx10877, A2=>
      nx10046);
   ix10045 : aoi22 port map ( Y=>nx10044, A0=>d_arr_merge2_0_18, A1=>nx10819, 
      B0=>d_arr_relu_0_18, B1=>nx10839);
   ix10047 : aoi222 port map ( Y=>nx10046, A0=>d_arr_mul_0_18, A1=>nx10589, 
      B0=>d_arr_add_0_18, B1=>nx10745, C0=>d_arr_merge1_0_18, C1=>nx10797);
   lat_d_arr_0_19 : latch port map ( Q=>d_arr_0_19, D=>nx8212, CLK=>nx10357
   );
   ix8213 : nand03 port map ( Y=>nx8212, A0=>nx10050, A1=>nx10877, A2=>
      nx10052);
   ix10051 : aoi22 port map ( Y=>nx10050, A0=>d_arr_merge2_0_19, A1=>nx10819, 
      B0=>d_arr_relu_0_19, B1=>nx10841);
   ix10053 : aoi222 port map ( Y=>nx10052, A0=>d_arr_mul_0_19, A1=>nx10589, 
      B0=>d_arr_add_0_19, B1=>nx10745, C0=>d_arr_merge1_0_19, C1=>nx10797);
   lat_d_arr_0_20 : latch port map ( Q=>d_arr_0_20, D=>nx8234, CLK=>nx10357
   );
   ix8235 : nand03 port map ( Y=>nx8234, A0=>nx10056, A1=>nx10877, A2=>
      nx10058);
   ix10057 : aoi22 port map ( Y=>nx10056, A0=>d_arr_merge2_0_20, A1=>nx10819, 
      B0=>d_arr_relu_0_20, B1=>nx10841);
   ix10059 : aoi222 port map ( Y=>nx10058, A0=>d_arr_mul_0_20, A1=>nx10589, 
      B0=>d_arr_add_0_20, B1=>nx10745, C0=>d_arr_merge1_0_20, C1=>nx10797);
   lat_d_arr_0_21 : latch port map ( Q=>d_arr_0_21, D=>nx8256, CLK=>nx10357
   );
   ix8257 : nand03 port map ( Y=>nx8256, A0=>nx10062, A1=>nx10877, A2=>
      nx10064);
   ix10063 : aoi22 port map ( Y=>nx10062, A0=>d_arr_merge2_0_21, A1=>nx10819, 
      B0=>d_arr_relu_0_21, B1=>nx10841);
   ix10065 : aoi222 port map ( Y=>nx10064, A0=>d_arr_mul_0_21, A1=>nx10589, 
      B0=>d_arr_add_0_21, B1=>nx10745, C0=>d_arr_merge1_0_21, C1=>nx10797);
   lat_d_arr_0_22 : latch port map ( Q=>d_arr_0_22, D=>nx8278, CLK=>nx10357
   );
   ix8279 : nand03 port map ( Y=>nx8278, A0=>nx10068, A1=>nx10879, A2=>
      nx10070);
   ix10069 : aoi22 port map ( Y=>nx10068, A0=>d_arr_merge2_0_22, A1=>nx10819, 
      B0=>d_arr_relu_0_22, B1=>nx10841);
   ix10071 : aoi222 port map ( Y=>nx10070, A0=>d_arr_mul_0_22, A1=>nx10589, 
      B0=>d_arr_add_0_22, B1=>nx10745, C0=>d_arr_merge1_0_22, C1=>nx10797);
   lat_d_arr_0_23 : latch port map ( Q=>d_arr_0_23, D=>nx8300, CLK=>nx10359
   );
   ix8301 : nand03 port map ( Y=>nx8300, A0=>nx10074, A1=>nx10879, A2=>
      nx10076);
   ix10075 : aoi22 port map ( Y=>nx10074, A0=>d_arr_merge2_0_23, A1=>nx10819, 
      B0=>d_arr_relu_0_23, B1=>nx10841);
   ix10077 : aoi222 port map ( Y=>nx10076, A0=>d_arr_mul_0_23, A1=>nx10591, 
      B0=>d_arr_add_0_23, B1=>nx10745, C0=>d_arr_merge1_0_23, C1=>nx10797);
   lat_d_arr_0_24 : latch port map ( Q=>d_arr_0_24, D=>nx8322, CLK=>nx10359
   );
   ix8323 : nand03 port map ( Y=>nx8322, A0=>nx10080, A1=>nx10879, A2=>
      nx10082);
   ix10081 : aoi22 port map ( Y=>nx10080, A0=>d_arr_merge2_0_24, A1=>nx10821, 
      B0=>d_arr_relu_0_24, B1=>nx10841);
   ix10083 : aoi222 port map ( Y=>nx10082, A0=>d_arr_mul_0_24, A1=>nx10591, 
      B0=>d_arr_add_0_24, B1=>nx10745, C0=>d_arr_merge1_0_24, C1=>nx10799);
   lat_d_arr_0_25 : latch port map ( Q=>d_arr_0_25, D=>nx8344, CLK=>nx10359
   );
   ix8345 : nand03 port map ( Y=>nx8344, A0=>nx10086, A1=>nx10879, A2=>
      nx10088);
   ix10087 : aoi22 port map ( Y=>nx10086, A0=>d_arr_merge2_0_25, A1=>nx10821, 
      B0=>d_arr_relu_0_25, B1=>nx10841);
   ix10089 : aoi222 port map ( Y=>nx10088, A0=>d_arr_mul_0_25, A1=>nx10591, 
      B0=>d_arr_add_0_25, B1=>nx10747, C0=>d_arr_merge1_0_25, C1=>nx10799);
   lat_d_arr_0_26 : latch port map ( Q=>d_arr_0_26, D=>nx8366, CLK=>nx10359
   );
   ix8367 : nand03 port map ( Y=>nx8366, A0=>nx10092, A1=>nx10879, A2=>
      nx10094);
   ix10093 : aoi22 port map ( Y=>nx10092, A0=>d_arr_merge2_0_26, A1=>nx10821, 
      B0=>d_arr_relu_0_26, B1=>nx10843);
   ix10095 : aoi222 port map ( Y=>nx10094, A0=>d_arr_mul_0_26, A1=>nx10591, 
      B0=>d_arr_add_0_26, B1=>nx10747, C0=>d_arr_merge1_0_26, C1=>nx10799);
   lat_d_arr_0_27 : latch port map ( Q=>d_arr_0_27, D=>nx8388, CLK=>nx10359
   );
   ix8389 : nand03 port map ( Y=>nx8388, A0=>nx10098, A1=>nx10879, A2=>
      nx10100);
   ix10099 : aoi22 port map ( Y=>nx10098, A0=>d_arr_merge2_0_27, A1=>nx10821, 
      B0=>d_arr_relu_0_27, B1=>nx10843);
   ix10101 : aoi222 port map ( Y=>nx10100, A0=>d_arr_mul_0_27, A1=>nx10591, 
      B0=>d_arr_add_0_27, B1=>nx10747, C0=>d_arr_merge1_0_27, C1=>nx10799);
   lat_d_arr_0_28 : latch port map ( Q=>d_arr_0_28, D=>nx8410, CLK=>nx10359
   );
   ix8411 : nand03 port map ( Y=>nx8410, A0=>nx10104, A1=>nx10879, A2=>
      nx10106);
   ix10105 : aoi22 port map ( Y=>nx10104, A0=>d_arr_merge2_0_28, A1=>nx10821, 
      B0=>d_arr_relu_0_28, B1=>nx10843);
   ix10107 : aoi222 port map ( Y=>nx10106, A0=>d_arr_mul_0_28, A1=>nx10591, 
      B0=>d_arr_add_0_28, B1=>nx10747, C0=>d_arr_merge1_0_28, C1=>nx10799);
   lat_d_arr_0_29 : latch port map ( Q=>d_arr_0_29, D=>nx8432, CLK=>nx10359
   );
   ix8433 : nand03 port map ( Y=>nx8432, A0=>nx10110, A1=>nx10026, A2=>
      nx10112);
   ix10111 : aoi22 port map ( Y=>nx10110, A0=>d_arr_merge2_0_29, A1=>nx10821, 
      B0=>d_arr_relu_0_29, B1=>nx10843);
   ix10113 : aoi222 port map ( Y=>nx10112, A0=>d_arr_mul_0_29, A1=>nx10591, 
      B0=>d_arr_add_0_29, B1=>nx10747, C0=>d_arr_merge1_0_29, C1=>nx10799);
   lat_d_arr_0_30 : latch port map ( Q=>d_arr_0_30, D=>nx8454, CLK=>nx10361
   );
   ix8455 : nand03 port map ( Y=>nx8454, A0=>nx10116, A1=>nx10026, A2=>
      nx10118);
   ix10117 : aoi22 port map ( Y=>nx10116, A0=>d_arr_merge2_0_30, A1=>nx10821, 
      B0=>d_arr_relu_0_30, B1=>nx10843);
   ix10119 : aoi222 port map ( Y=>nx10118, A0=>d_arr_mul_0_30, A1=>nx10593, 
      B0=>d_arr_add_0_30, B1=>nx10747, C0=>d_arr_merge1_0_30, C1=>nx10799);
   lat_d_arr_0_31 : latch port map ( Q=>d_arr_0_31, D=>nx8476, CLK=>nx10361
   );
   ix8477 : nand03 port map ( Y=>nx8476, A0=>nx10122, A1=>nx10026, A2=>
      nx10124);
   ix10123 : aoi22 port map ( Y=>nx10122, A0=>d_arr_merge2_0_31, A1=>nx10823, 
      B0=>d_arr_relu_0_31, B1=>nx10843);
   ix10125 : aoi222 port map ( Y=>nx10124, A0=>d_arr_mul_0_31, A1=>nx10593, 
      B0=>d_arr_add_0_31, B1=>nx10747, C0=>d_arr_merge1_0_31, C1=>nx10801);
   ix5 : inv01 port map ( Y=>nx4, A=>nx9734);
   ix10132 : inv02 port map ( Y=>nx10133, A=>nx10995);
   ix10134 : inv02 port map ( Y=>nx10135, A=>nx10995);
   ix10136 : inv02 port map ( Y=>nx10137, A=>nx10995);
   ix10138 : inv02 port map ( Y=>nx10139, A=>nx10995);
   ix10140 : inv02 port map ( Y=>nx10141, A=>nx10995);
   ix10142 : inv02 port map ( Y=>nx10143, A=>nx10995);
   ix10144 : inv02 port map ( Y=>nx10145, A=>nx10995);
   ix10146 : inv02 port map ( Y=>nx10147, A=>nx10883);
   ix10148 : inv02 port map ( Y=>nx10149, A=>nx10883);
   ix10150 : inv02 port map ( Y=>nx10151, A=>nx10883);
   ix10152 : inv02 port map ( Y=>nx10153, A=>nx10883);
   ix10154 : inv02 port map ( Y=>nx10155, A=>nx10883);
   ix10156 : inv02 port map ( Y=>nx10157, A=>nx10883);
   ix10158 : inv02 port map ( Y=>nx10159, A=>nx10883);
   ix10160 : inv02 port map ( Y=>nx10161, A=>nx10885);
   ix10162 : inv02 port map ( Y=>nx10163, A=>nx10885);
   ix10164 : inv02 port map ( Y=>nx10165, A=>nx10885);
   ix10166 : inv02 port map ( Y=>nx10167, A=>nx10885);
   ix10168 : inv02 port map ( Y=>nx10169, A=>nx10885);
   ix10170 : inv02 port map ( Y=>nx10171, A=>nx10885);
   ix10172 : inv02 port map ( Y=>nx10173, A=>nx10885);
   ix10174 : inv02 port map ( Y=>nx10175, A=>nx10887);
   ix10176 : inv02 port map ( Y=>nx10177, A=>nx10887);
   ix10178 : inv02 port map ( Y=>nx10179, A=>nx10887);
   ix10180 : inv02 port map ( Y=>nx10181, A=>nx10887);
   ix10182 : inv02 port map ( Y=>nx10183, A=>nx10887);
   ix10184 : inv02 port map ( Y=>nx10185, A=>nx10887);
   ix10186 : inv02 port map ( Y=>nx10187, A=>nx10887);
   ix10188 : inv02 port map ( Y=>nx10189, A=>nx10889);
   ix10190 : inv02 port map ( Y=>nx10191, A=>nx10889);
   ix10192 : inv02 port map ( Y=>nx10193, A=>nx10889);
   ix10194 : inv02 port map ( Y=>nx10195, A=>nx10889);
   ix10196 : inv02 port map ( Y=>nx10197, A=>nx10889);
   ix10198 : inv02 port map ( Y=>nx10199, A=>nx10889);
   ix10200 : inv02 port map ( Y=>nx10201, A=>nx10889);
   ix10202 : inv02 port map ( Y=>nx10203, A=>nx10891);
   ix10204 : inv02 port map ( Y=>nx10205, A=>nx10891);
   ix10206 : inv02 port map ( Y=>nx10207, A=>nx10891);
   ix10208 : inv02 port map ( Y=>nx10209, A=>nx10891);
   ix10210 : inv02 port map ( Y=>nx10211, A=>nx10891);
   ix10212 : inv02 port map ( Y=>nx10213, A=>nx10891);
   ix10214 : inv02 port map ( Y=>nx10215, A=>nx10891);
   ix10216 : inv02 port map ( Y=>nx10217, A=>nx10893);
   ix10218 : inv02 port map ( Y=>nx10219, A=>nx10893);
   ix10220 : inv02 port map ( Y=>nx10221, A=>nx10893);
   ix10222 : inv02 port map ( Y=>nx10223, A=>nx10893);
   ix10224 : inv02 port map ( Y=>nx10225, A=>nx10893);
   ix10226 : inv02 port map ( Y=>nx10227, A=>nx10893);
   ix10228 : inv02 port map ( Y=>nx10229, A=>nx10893);
   ix10230 : inv02 port map ( Y=>nx10231, A=>nx10895);
   ix10232 : inv02 port map ( Y=>nx10233, A=>nx10895);
   ix10234 : inv02 port map ( Y=>nx10235, A=>nx10895);
   ix10236 : inv02 port map ( Y=>nx10237, A=>nx10895);
   ix10238 : inv02 port map ( Y=>nx10239, A=>nx10895);
   ix10240 : inv02 port map ( Y=>nx10241, A=>nx10895);
   ix10242 : inv02 port map ( Y=>nx10243, A=>nx10895);
   ix10244 : inv02 port map ( Y=>nx10245, A=>nx10897);
   ix10246 : inv02 port map ( Y=>nx10247, A=>nx10897);
   ix10248 : inv02 port map ( Y=>nx10249, A=>nx10897);
   ix10250 : inv02 port map ( Y=>nx10251, A=>nx10897);
   ix10252 : inv02 port map ( Y=>nx10253, A=>nx10897);
   ix10254 : inv02 port map ( Y=>nx10255, A=>nx10897);
   ix10256 : inv02 port map ( Y=>nx10257, A=>nx10897);
   ix10258 : inv02 port map ( Y=>nx10259, A=>nx10899);
   ix10260 : inv02 port map ( Y=>nx10261, A=>nx10899);
   ix10262 : inv02 port map ( Y=>nx10263, A=>nx10899);
   ix10264 : inv02 port map ( Y=>nx10265, A=>nx10899);
   ix10266 : inv02 port map ( Y=>nx10267, A=>nx10899);
   ix10268 : inv02 port map ( Y=>nx10269, A=>nx10899);
   ix10270 : inv02 port map ( Y=>nx10271, A=>nx10899);
   ix10272 : inv02 port map ( Y=>nx10273, A=>nx10901);
   ix10274 : inv02 port map ( Y=>nx10275, A=>nx10901);
   ix10276 : inv02 port map ( Y=>nx10277, A=>nx10901);
   ix10278 : inv02 port map ( Y=>nx10279, A=>nx10901);
   ix10280 : inv02 port map ( Y=>nx10281, A=>nx10901);
   ix10282 : inv02 port map ( Y=>nx10283, A=>nx10901);
   ix10284 : inv02 port map ( Y=>nx10285, A=>nx10901);
   ix10286 : inv02 port map ( Y=>nx10287, A=>nx10903);
   ix10288 : inv02 port map ( Y=>nx10289, A=>nx10903);
   ix10290 : inv02 port map ( Y=>nx10291, A=>nx10903);
   ix10292 : inv02 port map ( Y=>nx10293, A=>nx10903);
   ix10294 : inv02 port map ( Y=>nx10295, A=>nx10903);
   ix10296 : inv02 port map ( Y=>nx10297, A=>nx10903);
   ix10298 : inv02 port map ( Y=>nx10299, A=>nx10903);
   ix10300 : inv02 port map ( Y=>nx10301, A=>nx10905);
   ix10302 : inv02 port map ( Y=>nx10303, A=>nx10905);
   ix10304 : inv02 port map ( Y=>nx10305, A=>nx10905);
   ix10306 : inv02 port map ( Y=>nx10307, A=>nx10905);
   ix10308 : inv02 port map ( Y=>nx10309, A=>nx10905);
   ix10310 : inv02 port map ( Y=>nx10311, A=>nx10905);
   ix10312 : inv02 port map ( Y=>nx10313, A=>nx10905);
   ix10314 : inv02 port map ( Y=>nx10315, A=>nx10907);
   ix10316 : inv02 port map ( Y=>nx10317, A=>nx10907);
   ix10318 : inv02 port map ( Y=>nx10319, A=>nx10907);
   ix10320 : inv02 port map ( Y=>nx10321, A=>nx10907);
   ix10322 : inv02 port map ( Y=>nx10323, A=>nx10907);
   ix10324 : inv02 port map ( Y=>nx10325, A=>nx10907);
   ix10326 : inv02 port map ( Y=>nx10327, A=>nx10907);
   ix10328 : inv02 port map ( Y=>nx10329, A=>nx10909);
   ix10330 : inv02 port map ( Y=>nx10331, A=>nx10909);
   ix10332 : inv02 port map ( Y=>nx10333, A=>nx10909);
   ix10334 : inv02 port map ( Y=>nx10335, A=>nx10909);
   ix10336 : inv02 port map ( Y=>nx10337, A=>nx10909);
   ix10338 : inv02 port map ( Y=>nx10339, A=>nx10909);
   ix10340 : inv02 port map ( Y=>nx10341, A=>nx10909);
   ix10342 : inv02 port map ( Y=>nx10343, A=>nx10911);
   ix10344 : inv02 port map ( Y=>nx10345, A=>nx10911);
   ix10346 : inv02 port map ( Y=>nx10347, A=>nx10911);
   ix10348 : inv02 port map ( Y=>nx10349, A=>nx10911);
   ix10350 : inv02 port map ( Y=>nx10351, A=>nx10911);
   ix10352 : inv02 port map ( Y=>nx10353, A=>nx10911);
   ix10354 : inv02 port map ( Y=>nx10355, A=>nx10911);
   ix10356 : inv02 port map ( Y=>nx10357, A=>nx10913);
   ix10358 : inv02 port map ( Y=>nx10359, A=>nx10913);
   ix10360 : inv02 port map ( Y=>nx10361, A=>nx10913);
   ix10364 : inv02 port map ( Y=>nx10365, A=>nx11471);
   ix10366 : inv02 port map ( Y=>nx10367, A=>nx11471);
   ix10368 : inv02 port map ( Y=>nx10369, A=>nx11471);
   ix10372 : inv02 port map ( Y=>nx10373, A=>nx11471);
   ix10374 : inv02 port map ( Y=>nx10375, A=>nx11471);
   ix10376 : inv02 port map ( Y=>nx10377, A=>nx11471);
   ix10382 : inv02 port map ( Y=>nx10383, A=>nx11435);
   ix10384 : inv02 port map ( Y=>nx10385, A=>nx11435);
   ix10386 : inv02 port map ( Y=>nx10387, A=>nx11435);
   ix10390 : inv02 port map ( Y=>nx10391, A=>nx11435);
   ix10392 : inv02 port map ( Y=>nx10393, A=>nx10919);
   ix10394 : inv02 port map ( Y=>nx10395, A=>nx10919);
   ix10396 : inv02 port map ( Y=>nx10397, A=>nx10919);
   ix10398 : inv02 port map ( Y=>nx10399, A=>nx10919);
   ix10400 : inv02 port map ( Y=>nx10401, A=>nx10919);
   ix10402 : inv02 port map ( Y=>nx10403, A=>nx10919);
   ix10404 : inv02 port map ( Y=>nx10405, A=>nx10919);
   ix10406 : inv02 port map ( Y=>nx10407, A=>nx10921);
   ix10408 : inv02 port map ( Y=>nx10409, A=>nx10921);
   ix10410 : inv02 port map ( Y=>nx10411, A=>nx10921);
   ix10412 : inv02 port map ( Y=>nx10413, A=>nx10921);
   ix10414 : inv02 port map ( Y=>nx10415, A=>nx10921);
   ix10416 : inv02 port map ( Y=>nx10417, A=>nx10921);
   ix10418 : inv02 port map ( Y=>nx10419, A=>nx10921);
   ix10420 : inv02 port map ( Y=>nx10421, A=>nx10923);
   ix10422 : inv02 port map ( Y=>nx10423, A=>nx10923);
   ix10424 : inv02 port map ( Y=>nx10425, A=>nx10923);
   ix10426 : inv02 port map ( Y=>nx10427, A=>nx10923);
   ix10428 : inv02 port map ( Y=>nx10429, A=>nx10923);
   ix10430 : inv02 port map ( Y=>nx10431, A=>nx10923);
   ix10432 : inv02 port map ( Y=>nx10433, A=>nx10923);
   ix10434 : inv02 port map ( Y=>nx10435, A=>nx10925);
   ix10436 : inv02 port map ( Y=>nx10437, A=>nx10925);
   ix10438 : inv02 port map ( Y=>nx10439, A=>nx10925);
   ix10440 : inv02 port map ( Y=>nx10441, A=>nx10925);
   ix10442 : inv02 port map ( Y=>nx10443, A=>nx10925);
   ix10444 : inv02 port map ( Y=>nx10445, A=>nx10925);
   ix10446 : inv02 port map ( Y=>nx10447, A=>nx10925);
   ix10448 : inv02 port map ( Y=>nx10449, A=>nx10927);
   ix10450 : inv02 port map ( Y=>nx10451, A=>nx10927);
   ix10452 : inv02 port map ( Y=>nx10453, A=>nx10927);
   ix10454 : inv02 port map ( Y=>nx10455, A=>nx10927);
   ix10456 : inv02 port map ( Y=>nx10457, A=>nx10927);
   ix10458 : inv02 port map ( Y=>nx10459, A=>nx10927);
   ix10460 : inv02 port map ( Y=>nx10461, A=>nx10927);
   ix10462 : inv02 port map ( Y=>nx10463, A=>nx10929);
   ix10464 : inv02 port map ( Y=>nx10465, A=>nx10929);
   ix10466 : inv02 port map ( Y=>nx10467, A=>nx10929);
   ix10468 : inv02 port map ( Y=>nx10469, A=>nx10929);
   ix10470 : inv02 port map ( Y=>nx10471, A=>nx10929);
   ix10472 : inv02 port map ( Y=>nx10473, A=>nx10929);
   ix10474 : inv02 port map ( Y=>nx10475, A=>nx10929);
   ix10476 : inv02 port map ( Y=>nx10477, A=>nx10931);
   ix10478 : inv02 port map ( Y=>nx10479, A=>nx10931);
   ix10480 : inv02 port map ( Y=>nx10481, A=>nx10931);
   ix10482 : inv02 port map ( Y=>nx10483, A=>nx10931);
   ix10484 : inv02 port map ( Y=>nx10485, A=>nx10931);
   ix10486 : inv02 port map ( Y=>nx10487, A=>nx10931);
   ix10488 : inv02 port map ( Y=>nx10489, A=>nx10931);
   ix10490 : inv02 port map ( Y=>nx10491, A=>nx10933);
   ix10492 : inv02 port map ( Y=>nx10493, A=>nx10933);
   ix10494 : inv02 port map ( Y=>nx10495, A=>nx10933);
   ix10496 : inv02 port map ( Y=>nx10497, A=>nx10933);
   ix10498 : inv02 port map ( Y=>nx10499, A=>nx10933);
   ix10500 : inv02 port map ( Y=>nx10501, A=>nx10933);
   ix10502 : inv02 port map ( Y=>nx10503, A=>nx10933);
   ix10504 : inv02 port map ( Y=>nx10505, A=>nx11445);
   ix10506 : inv02 port map ( Y=>nx10507, A=>nx11445);
   ix10508 : inv02 port map ( Y=>nx10509, A=>nx11445);
   ix10510 : inv02 port map ( Y=>nx10511, A=>nx11445);
   ix10512 : inv02 port map ( Y=>nx10513, A=>nx11445);
   ix10514 : inv02 port map ( Y=>nx10515, A=>nx11445);
   ix10518 : inv02 port map ( Y=>nx10519, A=>nx11449);
   ix10520 : inv02 port map ( Y=>nx10521, A=>nx11449);
   ix10522 : inv02 port map ( Y=>nx10523, A=>nx11449);
   ix10528 : inv02 port map ( Y=>nx10529, A=>nx11449);
   ix10530 : inv02 port map ( Y=>nx10531, A=>nx11449);
   ix10532 : inv02 port map ( Y=>nx10533, A=>nx11455);
   ix10536 : inv02 port map ( Y=>nx10537, A=>nx11455);
   ix10538 : inv02 port map ( Y=>nx10539, A=>nx11455);
   ix10540 : inv02 port map ( Y=>nx10541, A=>nx11455);
   ix10546 : inv02 port map ( Y=>nx10547, A=>nx11463);
   ix10548 : inv02 port map ( Y=>nx10549, A=>nx11463);
   ix10550 : inv02 port map ( Y=>nx10551, A=>nx11463);
   ix10552 : inv02 port map ( Y=>nx10553, A=>nx11463);
   ix10554 : inv02 port map ( Y=>nx10555, A=>nx11463);
   ix10556 : inv02 port map ( Y=>nx10557, A=>nx11463);
   ix10558 : inv02 port map ( Y=>nx10559, A=>nx11463);
   ix10560 : inv02 port map ( Y=>nx10561, A=>nx10943);
   ix10562 : inv02 port map ( Y=>nx10563, A=>nx10943);
   ix10564 : inv02 port map ( Y=>nx10565, A=>nx10943);
   ix10566 : inv02 port map ( Y=>nx10567, A=>nx10943);
   ix10568 : inv02 port map ( Y=>nx10569, A=>nx10943);
   ix10570 : inv02 port map ( Y=>nx10571, A=>nx10943);
   ix10572 : inv02 port map ( Y=>nx10573, A=>nx10943);
   ix10574 : inv02 port map ( Y=>nx10575, A=>nx10945);
   ix10576 : inv02 port map ( Y=>nx10577, A=>nx10945);
   ix10578 : inv02 port map ( Y=>nx10579, A=>nx10945);
   ix10580 : inv02 port map ( Y=>nx10581, A=>nx10945);
   ix10582 : inv02 port map ( Y=>nx10583, A=>nx10945);
   ix10584 : inv02 port map ( Y=>nx10585, A=>nx10945);
   ix10586 : inv02 port map ( Y=>nx10587, A=>nx10945);
   ix10588 : inv02 port map ( Y=>nx10589, A=>nx10947);
   ix10590 : inv02 port map ( Y=>nx10591, A=>nx10947);
   ix10592 : inv02 port map ( Y=>nx10593, A=>nx10947);
   ix10620 : inv02 port map ( Y=>nx10621, A=>nx10999);
   ix10622 : inv02 port map ( Y=>nx10623, A=>nx10999);
   ix10624 : inv02 port map ( Y=>nx10625, A=>nx10999);
   ix10626 : inv02 port map ( Y=>nx10627, A=>nx10999);
   ix10628 : inv02 port map ( Y=>nx10629, A=>nx10999);
   ix10630 : inv02 port map ( Y=>nx10631, A=>nx10999);
   ix10632 : inv02 port map ( Y=>nx10633, A=>nx10949);
   ix10634 : inv02 port map ( Y=>nx10635, A=>nx10951);
   ix10636 : inv02 port map ( Y=>nx10637, A=>nx10951);
   ix10638 : inv02 port map ( Y=>nx10639, A=>nx10951);
   ix10640 : inv02 port map ( Y=>nx10641, A=>nx10951);
   ix10642 : inv02 port map ( Y=>nx10643, A=>nx10951);
   ix10644 : inv02 port map ( Y=>nx10645, A=>nx10951);
   ix10646 : inv02 port map ( Y=>nx10647, A=>nx10951);
   ix10648 : inv02 port map ( Y=>nx10649, A=>nx10953);
   ix10650 : inv02 port map ( Y=>nx10651, A=>nx10953);
   ix10652 : inv02 port map ( Y=>nx10653, A=>nx10953);
   ix10654 : inv02 port map ( Y=>nx10655, A=>nx10953);
   ix10656 : inv02 port map ( Y=>nx10657, A=>nx10953);
   ix10658 : inv02 port map ( Y=>nx10659, A=>nx10953);
   ix10660 : inv02 port map ( Y=>nx10661, A=>nx10953);
   ix10662 : inv02 port map ( Y=>nx10663, A=>nx10955);
   ix10664 : inv02 port map ( Y=>nx10665, A=>nx10955);
   ix10666 : inv02 port map ( Y=>nx10667, A=>nx10955);
   ix10668 : inv02 port map ( Y=>nx10669, A=>nx10955);
   ix10670 : inv02 port map ( Y=>nx10671, A=>nx10955);
   ix10672 : inv02 port map ( Y=>nx10673, A=>nx10955);
   ix10674 : inv02 port map ( Y=>nx10675, A=>nx10955);
   ix10676 : inv02 port map ( Y=>nx10677, A=>nx10957);
   ix10678 : inv02 port map ( Y=>nx10679, A=>nx10957);
   ix10680 : inv02 port map ( Y=>nx10681, A=>nx10957);
   ix10682 : inv02 port map ( Y=>nx10683, A=>nx10957);
   ix10684 : inv02 port map ( Y=>nx10685, A=>nx10957);
   ix10686 : inv02 port map ( Y=>nx10687, A=>nx10957);
   ix10688 : inv02 port map ( Y=>nx10689, A=>nx10957);
   ix10690 : inv02 port map ( Y=>nx10691, A=>nx10959);
   ix10692 : inv02 port map ( Y=>nx10693, A=>nx10959);
   ix10694 : inv02 port map ( Y=>nx10695, A=>nx10959);
   ix10696 : inv02 port map ( Y=>nx10697, A=>nx10959);
   ix10698 : inv02 port map ( Y=>nx10699, A=>nx10959);
   ix10700 : inv02 port map ( Y=>nx10701, A=>nx10959);
   ix10702 : inv02 port map ( Y=>nx10703, A=>nx10959);
   ix10704 : inv02 port map ( Y=>nx10705, A=>nx10961);
   ix10706 : inv02 port map ( Y=>nx10707, A=>nx10961);
   ix10708 : inv02 port map ( Y=>nx10709, A=>nx10961);
   ix10710 : inv02 port map ( Y=>nx10711, A=>nx10961);
   ix10712 : inv02 port map ( Y=>nx10713, A=>nx10961);
   ix10714 : inv02 port map ( Y=>nx10715, A=>nx10961);
   ix10716 : inv02 port map ( Y=>nx10717, A=>nx10961);
   ix10718 : inv02 port map ( Y=>nx10719, A=>nx10963);
   ix10720 : inv02 port map ( Y=>nx10721, A=>nx10963);
   ix10722 : inv02 port map ( Y=>nx10723, A=>nx10963);
   ix10724 : inv02 port map ( Y=>nx10725, A=>nx10963);
   ix10726 : inv02 port map ( Y=>nx10727, A=>nx10963);
   ix10728 : inv02 port map ( Y=>nx10729, A=>nx10963);
   ix10730 : inv02 port map ( Y=>nx10731, A=>nx10963);
   ix10732 : inv02 port map ( Y=>nx10733, A=>nx10965);
   ix10734 : inv02 port map ( Y=>nx10735, A=>nx10965);
   ix10736 : inv02 port map ( Y=>nx10737, A=>nx10965);
   ix10738 : inv02 port map ( Y=>nx10739, A=>nx10965);
   ix10740 : inv02 port map ( Y=>nx10741, A=>nx10965);
   ix10742 : inv02 port map ( Y=>nx10743, A=>nx10965);
   ix10744 : inv02 port map ( Y=>nx10745, A=>nx10965);
   ix10746 : inv02 port map ( Y=>nx10747, A=>nx10967);
   ix10780 : inv01 port map ( Y=>nx10781, A=>nx7002);
   ix10782 : inv02 port map ( Y=>nx10783, A=>nx10969);
   ix10784 : inv02 port map ( Y=>nx10785, A=>nx10969);
   ix10786 : inv02 port map ( Y=>nx10787, A=>nx10969);
   ix10788 : inv02 port map ( Y=>nx10789, A=>nx10969);
   ix10790 : inv02 port map ( Y=>nx10791, A=>nx10969);
   ix10792 : inv02 port map ( Y=>nx10793, A=>nx10781);
   ix10794 : inv02 port map ( Y=>nx10795, A=>nx10781);
   ix10796 : inv02 port map ( Y=>nx10797, A=>nx10781);
   ix10798 : inv02 port map ( Y=>nx10799, A=>nx10781);
   ix10800 : inv02 port map ( Y=>nx10801, A=>nx10781);
   ix10802 : inv01 port map ( Y=>nx10803, A=>nx7018);
   ix10804 : inv02 port map ( Y=>nx10805, A=>nx10971);
   ix10806 : inv02 port map ( Y=>nx10807, A=>nx10971);
   ix10808 : inv02 port map ( Y=>nx10809, A=>nx10971);
   ix10810 : inv02 port map ( Y=>nx10811, A=>nx10971);
   ix10812 : inv02 port map ( Y=>nx10813, A=>nx10971);
   ix10814 : inv02 port map ( Y=>nx10815, A=>nx10803);
   ix10816 : inv02 port map ( Y=>nx10817, A=>nx10803);
   ix10818 : inv02 port map ( Y=>nx10819, A=>nx10803);
   ix10820 : inv02 port map ( Y=>nx10821, A=>nx10803);
   ix10822 : inv02 port map ( Y=>nx10823, A=>nx10803);
   ix10824 : inv01 port map ( Y=>nx10825, A=>nx7028);
   ix10826 : inv02 port map ( Y=>nx10827, A=>nx10973);
   ix10828 : inv02 port map ( Y=>nx10829, A=>nx10973);
   ix10830 : inv02 port map ( Y=>nx10831, A=>nx10973);
   ix10832 : inv02 port map ( Y=>nx10833, A=>nx10973);
   ix10834 : inv02 port map ( Y=>nx10835, A=>nx10973);
   ix10836 : inv02 port map ( Y=>nx10837, A=>nx10825);
   ix10838 : inv02 port map ( Y=>nx10839, A=>nx10825);
   ix10840 : inv02 port map ( Y=>nx10841, A=>nx10825);
   ix10842 : inv02 port map ( Y=>nx10843, A=>nx10825);
   ix10844 : nand02 port map ( Y=>nx10845, A0=>d_arr_mux_21_31, A1=>nx11399
   );
   ix10846 : nand02 port map ( Y=>nx10847, A0=>d_arr_mux_21_31, A1=>nx11399
   );
   ix10848 : nand02 port map ( Y=>nx10849, A0=>d_arr_mux_20_31, A1=>nx11399
   );
   ix10850 : nand02 port map ( Y=>nx10851, A0=>d_arr_mux_20_31, A1=>nx11399
   );
   ix10852 : nand02 port map ( Y=>nx10853, A0=>d_arr_mux_19_31, A1=>nx11399
   );
   ix10854 : nand02 port map ( Y=>nx10855, A0=>d_arr_mux_19_31, A1=>nx11401
   );
   ix10856 : nand02 port map ( Y=>nx10857, A0=>d_arr_mux_18_31, A1=>nx11401
   );
   ix10858 : nand02 port map ( Y=>nx10859, A0=>d_arr_mux_18_31, A1=>nx11401
   );
   ix10860 : nand02 port map ( Y=>nx10861, A0=>d_arr_mux_4_31, A1=>nx11401);
   ix10862 : nand02 port map ( Y=>nx10863, A0=>d_arr_mux_4_31, A1=>nx11401);
   ix10864 : nand02 port map ( Y=>nx10865, A0=>d_arr_mux_3_31, A1=>nx11401);
   ix10866 : nand02 port map ( Y=>nx10867, A0=>d_arr_mux_3_31, A1=>nx11401);
   ix10868 : nand02 port map ( Y=>nx10869, A0=>d_arr_mux_2_31, A1=>nx11501);
   ix10870 : nand02 port map ( Y=>nx10871, A0=>d_arr_mux_2_31, A1=>nx11501);
   ix10872 : nand02 port map ( Y=>nx10873, A0=>d_arr_mux_1_31, A1=>nx11501);
   ix10874 : nand02 port map ( Y=>nx10875, A0=>d_arr_mux_1_31, A1=>nx11501);
   ix10876 : nand02 port map ( Y=>nx10877, A0=>d_arr_mux_0_31, A1=>nx11501);
   ix10878 : nand02 port map ( Y=>nx10879, A0=>d_arr_mux_0_31, A1=>nx11501);
   ix10880 : inv02 port map ( Y=>nx10881, A=>nx8);
   ix10882 : inv02 port map ( Y=>nx10883, A=>nx10979);
   ix10884 : inv02 port map ( Y=>nx10885, A=>nx10979);
   ix10886 : inv02 port map ( Y=>nx10887, A=>nx10979);
   ix10888 : inv02 port map ( Y=>nx10889, A=>nx10979);
   ix10890 : inv02 port map ( Y=>nx10891, A=>nx10979);
   ix10892 : inv02 port map ( Y=>nx10893, A=>nx10979);
   ix10894 : inv02 port map ( Y=>nx10895, A=>nx10979);
   ix10896 : inv02 port map ( Y=>nx10897, A=>nx10981);
   ix10898 : inv02 port map ( Y=>nx10899, A=>nx10981);
   ix10900 : inv02 port map ( Y=>nx10901, A=>nx10981);
   ix10902 : inv02 port map ( Y=>nx10903, A=>nx10981);
   ix10904 : inv02 port map ( Y=>nx10905, A=>nx10981);
   ix10906 : inv02 port map ( Y=>nx10907, A=>nx10981);
   ix10908 : inv02 port map ( Y=>nx10909, A=>nx10981);
   ix10910 : inv02 port map ( Y=>nx10911, A=>nx10983);
   ix10912 : inv02 port map ( Y=>nx10913, A=>nx10983);
   ix10914 : inv02 port map ( Y=>nx10915, A=>nx12);
   ix10916 : inv02 port map ( Y=>nx10917, A=>nx11465);
   ix10918 : inv02 port map ( Y=>nx10919, A=>nx11465);
   ix10920 : inv02 port map ( Y=>nx10921, A=>nx11465);
   ix10922 : inv02 port map ( Y=>nx10923, A=>nx11465);
   ix10924 : inv02 port map ( Y=>nx10925, A=>nx11465);
   ix10926 : inv02 port map ( Y=>nx10927, A=>nx11465);
   ix10928 : inv02 port map ( Y=>nx10929, A=>nx11465);
   ix10930 : inv02 port map ( Y=>nx10931, A=>nx11467);
   ix10932 : inv02 port map ( Y=>nx10933, A=>nx11467);
   ix10934 : inv02 port map ( Y=>nx10935, A=>nx11467);
   ix10936 : inv02 port map ( Y=>nx10937, A=>nx11467);
   ix10938 : inv02 port map ( Y=>nx10939, A=>nx11467);
   ix10940 : inv02 port map ( Y=>nx10941, A=>nx11467);
   ix10942 : inv02 port map ( Y=>nx10943, A=>nx11467);
   ix10944 : inv02 port map ( Y=>nx10945, A=>nx10989);
   ix10946 : inv02 port map ( Y=>nx10947, A=>nx10989);
   ix10948 : inv02 port map ( Y=>nx10949, A=>nx694);
   ix10950 : inv02 port map ( Y=>nx10951, A=>nx10991);
   ix10952 : inv02 port map ( Y=>nx10953, A=>nx10991);
   ix10954 : inv02 port map ( Y=>nx10955, A=>nx10991);
   ix10956 : inv02 port map ( Y=>nx10957, A=>nx10991);
   ix10958 : inv02 port map ( Y=>nx10959, A=>nx10991);
   ix10960 : inv02 port map ( Y=>nx10961, A=>nx10993);
   ix10962 : inv02 port map ( Y=>nx10963, A=>nx10993);
   ix10964 : inv02 port map ( Y=>nx10965, A=>nx10993);
   ix10966 : inv02 port map ( Y=>nx10967, A=>nx10993);
   ix10968 : inv01 port map ( Y=>nx10969, A=>nx7002);
   ix10970 : inv01 port map ( Y=>nx10971, A=>nx7018);
   ix10972 : inv01 port map ( Y=>nx10973, A=>nx7028);
   ix10978 : inv02 port map ( Y=>nx10979, A=>nx10881);
   ix10980 : inv02 port map ( Y=>nx10981, A=>nx10881);
   ix10982 : inv02 port map ( Y=>nx10983, A=>nx10881);
   ix10984 : inv02 port map ( Y=>nx10985, A=>nx10915);
   ix10986 : inv02 port map ( Y=>nx10987, A=>nx10915);
   ix10988 : inv02 port map ( Y=>nx10989, A=>nx10915);
   ix10990 : inv01 port map ( Y=>nx10991, A=>nx10999);
   ix10992 : inv01 port map ( Y=>nx10993, A=>nx10949);
   ix10994 : inv02 port map ( Y=>nx10995, A=>nx8);
   ix10996 : inv02 port map ( Y=>nx10997, A=>nx11511);
   ix10998 : inv02 port map ( Y=>nx10999, A=>nx694);
   ix141 : oai21 port map ( Y=>nx140, A0=>nx11005, A1=>nx11471, B0=>nx11407
   );
   ix11004 : inv01 port map ( Y=>nx11005, A=>d_arr_mul_24_15);
   ix137 : nand02 port map ( Y=>nx10595, A0=>nx11501, A1=>d_arr_mux_24_31);
   ix147 : oai21 port map ( Y=>nx146, A0=>nx11007, A1=>nx11473, B0=>nx11407
   );
   ix11006 : inv01 port map ( Y=>nx11007, A=>d_arr_mul_24_16);
   ix153 : oai21 port map ( Y=>nx152, A0=>nx11009, A1=>nx11473, B0=>nx11407
   );
   ix11008 : inv01 port map ( Y=>nx11009, A=>d_arr_mul_24_17);
   ix159 : oai21 port map ( Y=>nx158, A0=>nx11011, A1=>nx11473, B0=>nx11407
   );
   ix11010 : inv01 port map ( Y=>nx11011, A=>d_arr_mul_24_18);
   ix165 : oai21 port map ( Y=>nx164, A0=>nx11013, A1=>nx11473, B0=>nx11407
   );
   ix11012 : inv01 port map ( Y=>nx11013, A=>d_arr_mul_24_19);
   ix171 : oai21 port map ( Y=>nx170, A0=>nx11015, A1=>nx11473, B0=>nx11407
   );
   ix11014 : inv01 port map ( Y=>nx11015, A=>d_arr_mul_24_20);
   ix177 : oai21 port map ( Y=>nx176, A0=>nx11017, A1=>nx11473, B0=>nx11407
   );
   ix11016 : inv01 port map ( Y=>nx11017, A=>d_arr_mul_24_21);
   ix183 : oai21 port map ( Y=>nx182, A0=>nx11019, A1=>nx11473, B0=>nx11409
   );
   ix11018 : inv01 port map ( Y=>nx11019, A=>d_arr_mul_24_22);
   ix189 : oai21 port map ( Y=>nx188, A0=>nx11021, A1=>nx11475, B0=>nx11409
   );
   ix11020 : inv01 port map ( Y=>nx11021, A=>d_arr_mul_24_23);
   ix195 : oai21 port map ( Y=>nx194, A0=>nx11023, A1=>nx11475, B0=>nx11409
   );
   ix11022 : inv01 port map ( Y=>nx11023, A=>d_arr_mul_24_24);
   ix201 : oai21 port map ( Y=>nx200, A0=>nx11025, A1=>nx11475, B0=>nx11409
   );
   ix11024 : inv01 port map ( Y=>nx11025, A=>d_arr_mul_24_25);
   ix207 : oai21 port map ( Y=>nx206, A0=>nx11027, A1=>nx11475, B0=>nx11409
   );
   ix11026 : inv01 port map ( Y=>nx11027, A=>d_arr_mul_24_26);
   ix213 : oai21 port map ( Y=>nx212, A0=>nx11029, A1=>nx11475, B0=>nx11409
   );
   ix11028 : inv01 port map ( Y=>nx11029, A=>d_arr_mul_24_27);
   ix219 : oai21 port map ( Y=>nx218, A0=>nx11031, A1=>nx11475, B0=>nx11409
   );
   ix11030 : inv01 port map ( Y=>nx11031, A=>d_arr_mul_24_28);
   ix225 : oai21 port map ( Y=>nx224, A0=>nx11033, A1=>nx11475, B0=>nx10595
   );
   ix11032 : inv01 port map ( Y=>nx11033, A=>d_arr_mul_24_29);
   ix231 : oai21 port map ( Y=>nx230, A0=>nx11035, A1=>nx10997, B0=>nx10595
   );
   ix11034 : inv01 port map ( Y=>nx11035, A=>d_arr_mul_24_30);
   ix237 : oai21 port map ( Y=>nx236, A0=>nx11037, A1=>nx10997, B0=>nx10595
   );
   ix11036 : inv01 port map ( Y=>nx11037, A=>d_arr_mul_24_31);
   ix365 : oai21 port map ( Y=>nx364, A0=>nx11039, A1=>nx10997, B0=>nx11411
   );
   ix11038 : inv01 port map ( Y=>nx11039, A=>d_arr_mul_23_15);
   ix361 : nand02 port map ( Y=>nx10603, A0=>nx11503, A1=>d_arr_mux_23_31);
   ix371 : oai21 port map ( Y=>nx370, A0=>nx11041, A1=>nx10997, B0=>nx11411
   );
   ix11040 : inv01 port map ( Y=>nx11041, A=>d_arr_mul_23_16);
   ix377 : oai21 port map ( Y=>nx376, A0=>nx11043, A1=>nx11435, B0=>nx11411
   );
   ix11042 : inv01 port map ( Y=>nx11043, A=>d_arr_mul_23_17);
   ix383 : oai21 port map ( Y=>nx382, A0=>nx11045, A1=>nx11435, B0=>nx11411
   );
   ix11044 : inv01 port map ( Y=>nx11045, A=>d_arr_mul_23_18);
   ix389 : oai21 port map ( Y=>nx388, A0=>nx11047, A1=>nx11435, B0=>nx11411
   );
   ix11046 : inv01 port map ( Y=>nx11047, A=>d_arr_mul_23_19);
   ix395 : oai21 port map ( Y=>nx394, A0=>nx11049, A1=>nx11437, B0=>nx11411
   );
   ix11048 : inv01 port map ( Y=>nx11049, A=>d_arr_mul_23_20);
   ix401 : oai21 port map ( Y=>nx400, A0=>nx11051, A1=>nx11437, B0=>nx11411
   );
   ix11050 : inv01 port map ( Y=>nx11051, A=>d_arr_mul_23_21);
   ix407 : oai21 port map ( Y=>nx406, A0=>nx11053, A1=>nx11437, B0=>nx11413
   );
   ix11052 : inv01 port map ( Y=>nx11053, A=>d_arr_mul_23_22);
   ix413 : oai21 port map ( Y=>nx412, A0=>nx11055, A1=>nx11437, B0=>nx11413
   );
   ix11054 : inv01 port map ( Y=>nx11055, A=>d_arr_mul_23_23);
   ix419 : oai21 port map ( Y=>nx418, A0=>nx11057, A1=>nx11437, B0=>nx11413
   );
   ix11056 : inv01 port map ( Y=>nx11057, A=>d_arr_mul_23_24);
   ix425 : oai21 port map ( Y=>nx424, A0=>nx11059, A1=>nx11437, B0=>nx11413
   );
   ix11058 : inv01 port map ( Y=>nx11059, A=>d_arr_mul_23_25);
   ix431 : oai21 port map ( Y=>nx430, A0=>nx11061, A1=>nx11437, B0=>nx11413
   );
   ix11060 : inv01 port map ( Y=>nx11061, A=>d_arr_mul_23_26);
   ix437 : oai21 port map ( Y=>nx436, A0=>nx11063, A1=>nx11439, B0=>nx11413
   );
   ix11062 : inv01 port map ( Y=>nx11063, A=>d_arr_mul_23_27);
   ix443 : oai21 port map ( Y=>nx442, A0=>nx11065, A1=>nx11439, B0=>nx11413
   );
   ix11064 : inv01 port map ( Y=>nx11065, A=>d_arr_mul_23_28);
   ix449 : oai21 port map ( Y=>nx448, A0=>nx11067, A1=>nx11439, B0=>nx10603
   );
   ix11066 : inv01 port map ( Y=>nx11067, A=>d_arr_mul_23_29);
   ix455 : oai21 port map ( Y=>nx454, A0=>nx11069, A1=>nx11439, B0=>nx10603
   );
   ix11068 : inv01 port map ( Y=>nx11069, A=>d_arr_mul_23_30);
   ix461 : oai21 port map ( Y=>nx460, A0=>nx11071, A1=>nx11439, B0=>nx10603
   );
   ix11070 : inv01 port map ( Y=>nx11071, A=>d_arr_mul_23_31);
   ix589 : oai21 port map ( Y=>nx588, A0=>nx11073, A1=>nx11439, B0=>nx11415
   );
   ix11072 : inv01 port map ( Y=>nx11073, A=>d_arr_mul_22_15);
   ix585 : nand02 port map ( Y=>nx10611, A0=>nx11503, A1=>d_arr_mux_22_31);
   ix595 : oai21 port map ( Y=>nx594, A0=>nx11075, A1=>nx11439, B0=>nx11415
   );
   ix11074 : inv01 port map ( Y=>nx11075, A=>d_arr_mul_22_16);
   ix601 : oai21 port map ( Y=>nx600, A0=>nx11077, A1=>nx11441, B0=>nx11415
   );
   ix11076 : inv01 port map ( Y=>nx11077, A=>d_arr_mul_22_17);
   ix607 : oai21 port map ( Y=>nx606, A0=>nx11079, A1=>nx11441, B0=>nx11415
   );
   ix11078 : inv01 port map ( Y=>nx11079, A=>d_arr_mul_22_18);
   ix613 : oai21 port map ( Y=>nx612, A0=>nx11081, A1=>nx11441, B0=>nx11415
   );
   ix11080 : inv01 port map ( Y=>nx11081, A=>d_arr_mul_22_19);
   ix619 : oai21 port map ( Y=>nx618, A0=>nx11083, A1=>nx11441, B0=>nx11415
   );
   ix11082 : inv01 port map ( Y=>nx11083, A=>d_arr_mul_22_20);
   ix625 : oai21 port map ( Y=>nx624, A0=>nx11085, A1=>nx11441, B0=>nx11415
   );
   ix11084 : inv01 port map ( Y=>nx11085, A=>d_arr_mul_22_21);
   ix631 : oai21 port map ( Y=>nx630, A0=>nx11087, A1=>nx11441, B0=>nx11417
   );
   ix11086 : inv01 port map ( Y=>nx11087, A=>d_arr_mul_22_22);
   ix637 : oai21 port map ( Y=>nx636, A0=>nx11089, A1=>nx11441, B0=>nx11417
   );
   ix11088 : inv01 port map ( Y=>nx11089, A=>d_arr_mul_22_23);
   ix643 : oai21 port map ( Y=>nx642, A0=>nx11091, A1=>nx11443, B0=>nx11417
   );
   ix11090 : inv01 port map ( Y=>nx11091, A=>d_arr_mul_22_24);
   ix649 : oai21 port map ( Y=>nx648, A0=>nx11093, A1=>nx11443, B0=>nx11417
   );
   ix11092 : inv01 port map ( Y=>nx11093, A=>d_arr_mul_22_25);
   ix655 : oai21 port map ( Y=>nx654, A0=>nx11095, A1=>nx11443, B0=>nx11417
   );
   ix11094 : inv01 port map ( Y=>nx11095, A=>d_arr_mul_22_26);
   ix661 : oai21 port map ( Y=>nx660, A0=>nx11097, A1=>nx11443, B0=>nx11417
   );
   ix11096 : inv01 port map ( Y=>nx11097, A=>d_arr_mul_22_27);
   ix667 : oai21 port map ( Y=>nx666, A0=>nx11099, A1=>nx11443, B0=>nx11417
   );
   ix11098 : inv01 port map ( Y=>nx11099, A=>d_arr_mul_22_28);
   ix673 : oai21 port map ( Y=>nx672, A0=>nx11101, A1=>nx11443, B0=>nx10611
   );
   ix11100 : inv01 port map ( Y=>nx11101, A=>d_arr_mul_22_29);
   ix679 : oai21 port map ( Y=>nx678, A0=>nx11103, A1=>nx11443, B0=>nx10611
   );
   ix11102 : inv01 port map ( Y=>nx11103, A=>d_arr_mul_22_30);
   ix685 : oai21 port map ( Y=>nx684, A0=>nx11105, A1=>nx10917, B0=>nx10611
   );
   ix11104 : inv01 port map ( Y=>nx11105, A=>d_arr_mul_22_31);
   ix5169 : oai21 port map ( Y=>nx5168, A0=>nx11107, A1=>nx11445, B0=>
      nx11419);
   ix11106 : inv01 port map ( Y=>nx11107, A=>d_arr_mul_8_15);
   ix5165 : nand02 port map ( Y=>nx10749, A0=>nx11503, A1=>d_arr_mux_8_31);
   ix5175 : oai21 port map ( Y=>nx5174, A0=>nx11109, A1=>nx11447, B0=>
      nx11419);
   ix11108 : inv01 port map ( Y=>nx11109, A=>d_arr_mul_8_16);
   ix5181 : oai21 port map ( Y=>nx5180, A0=>nx11111, A1=>nx11447, B0=>
      nx11419);
   ix11110 : inv01 port map ( Y=>nx11111, A=>d_arr_mul_8_17);
   ix5187 : oai21 port map ( Y=>nx5186, A0=>nx11113, A1=>nx11447, B0=>
      nx11419);
   ix11112 : inv01 port map ( Y=>nx11113, A=>d_arr_mul_8_18);
   ix5193 : oai21 port map ( Y=>nx5192, A0=>nx11115, A1=>nx11447, B0=>
      nx11419);
   ix11114 : inv01 port map ( Y=>nx11115, A=>d_arr_mul_8_19);
   ix5199 : oai21 port map ( Y=>nx5198, A0=>nx11117, A1=>nx11447, B0=>
      nx11419);
   ix11116 : inv01 port map ( Y=>nx11117, A=>d_arr_mul_8_20);
   ix5205 : oai21 port map ( Y=>nx5204, A0=>nx11119, A1=>nx11447, B0=>
      nx11419);
   ix11118 : inv01 port map ( Y=>nx11119, A=>d_arr_mul_8_21);
   ix5211 : oai21 port map ( Y=>nx5210, A0=>nx11121, A1=>nx11447, B0=>
      nx11421);
   ix11120 : inv01 port map ( Y=>nx11121, A=>d_arr_mul_8_22);
   ix5217 : oai21 port map ( Y=>nx5216, A0=>nx11123, A1=>nx10935, B0=>
      nx11421);
   ix11122 : inv01 port map ( Y=>nx11123, A=>d_arr_mul_8_23);
   ix5223 : oai21 port map ( Y=>nx5222, A0=>nx11125, A1=>nx10935, B0=>
      nx11421);
   ix11124 : inv01 port map ( Y=>nx11125, A=>d_arr_mul_8_24);
   ix5229 : oai21 port map ( Y=>nx5228, A0=>nx11127, A1=>nx10935, B0=>
      nx11421);
   ix11126 : inv01 port map ( Y=>nx11127, A=>d_arr_mul_8_25);
   ix5235 : oai21 port map ( Y=>nx5234, A0=>nx11129, A1=>nx10935, B0=>
      nx11421);
   ix11128 : inv01 port map ( Y=>nx11129, A=>d_arr_mul_8_26);
   ix5241 : oai21 port map ( Y=>nx5240, A0=>nx11131, A1=>nx11449, B0=>
      nx11421);
   ix11130 : inv01 port map ( Y=>nx11131, A=>d_arr_mul_8_27);
   ix5247 : oai21 port map ( Y=>nx5246, A0=>nx11133, A1=>nx11449, B0=>
      nx11421);
   ix11132 : inv01 port map ( Y=>nx11133, A=>d_arr_mul_8_28);
   ix5253 : oai21 port map ( Y=>nx5252, A0=>nx11135, A1=>nx11451, B0=>
      nx10749);
   ix11134 : inv01 port map ( Y=>nx11135, A=>d_arr_mul_8_29);
   ix5259 : oai21 port map ( Y=>nx5258, A0=>nx11137, A1=>nx11451, B0=>
      nx10749);
   ix11136 : inv01 port map ( Y=>nx11137, A=>d_arr_mul_8_30);
   ix5265 : oai21 port map ( Y=>nx5264, A0=>nx11139, A1=>nx11451, B0=>
      nx10749);
   ix11138 : inv01 port map ( Y=>nx11139, A=>d_arr_mul_8_31);
   ix5393 : oai21 port map ( Y=>nx5392, A0=>nx11141, A1=>nx11451, B0=>
      nx11423);
   ix11140 : inv01 port map ( Y=>nx11141, A=>d_arr_mul_7_15);
   ix5389 : nand02 port map ( Y=>nx10757, A0=>nx11503, A1=>d_arr_mux_7_31);
   ix5399 : oai21 port map ( Y=>nx5398, A0=>nx11143, A1=>nx11451, B0=>
      nx11423);
   ix11142 : inv01 port map ( Y=>nx11143, A=>d_arr_mul_7_16);
   ix5405 : oai21 port map ( Y=>nx5404, A0=>nx11145, A1=>nx11451, B0=>
      nx11423);
   ix11144 : inv01 port map ( Y=>nx11145, A=>d_arr_mul_7_17);
   ix5411 : oai21 port map ( Y=>nx5410, A0=>nx11147, A1=>nx11451, B0=>
      nx11423);
   ix11146 : inv01 port map ( Y=>nx11147, A=>d_arr_mul_7_18);
   ix5417 : oai21 port map ( Y=>nx5416, A0=>nx11149, A1=>nx11453, B0=>
      nx11423);
   ix11148 : inv01 port map ( Y=>nx11149, A=>d_arr_mul_7_19);
   ix5423 : oai21 port map ( Y=>nx5422, A0=>nx11151, A1=>nx11453, B0=>
      nx11423);
   ix11150 : inv01 port map ( Y=>nx11151, A=>d_arr_mul_7_20);
   ix5429 : oai21 port map ( Y=>nx5428, A0=>nx11153, A1=>nx11453, B0=>
      nx11423);
   ix11152 : inv01 port map ( Y=>nx11153, A=>d_arr_mul_7_21);
   ix5435 : oai21 port map ( Y=>nx5434, A0=>nx11155, A1=>nx11453, B0=>
      nx11425);
   ix11154 : inv01 port map ( Y=>nx11155, A=>d_arr_mul_7_22);
   ix5441 : oai21 port map ( Y=>nx5440, A0=>nx11157, A1=>nx11453, B0=>
      nx11425);
   ix11156 : inv01 port map ( Y=>nx11157, A=>d_arr_mul_7_23);
   ix5447 : oai21 port map ( Y=>nx5446, A0=>nx11159, A1=>nx11453, B0=>
      nx11425);
   ix11158 : inv01 port map ( Y=>nx11159, A=>d_arr_mul_7_24);
   ix5453 : oai21 port map ( Y=>nx5452, A0=>nx11161, A1=>nx11453, B0=>
      nx11425);
   ix11160 : inv01 port map ( Y=>nx11161, A=>d_arr_mul_7_25);
   ix5459 : oai21 port map ( Y=>nx5458, A0=>nx11163, A1=>nx10937, B0=>
      nx11425);
   ix11162 : inv01 port map ( Y=>nx11163, A=>d_arr_mul_7_26);
   ix5465 : oai21 port map ( Y=>nx5464, A0=>nx11165, A1=>nx10937, B0=>
      nx11425);
   ix11164 : inv01 port map ( Y=>nx11165, A=>d_arr_mul_7_27);
   ix5471 : oai21 port map ( Y=>nx5470, A0=>nx11167, A1=>nx10937, B0=>
      nx11425);
   ix11166 : inv01 port map ( Y=>nx11167, A=>d_arr_mul_7_28);
   ix5477 : oai21 port map ( Y=>nx5476, A0=>nx11169, A1=>nx10937, B0=>
      nx10757);
   ix11168 : inv01 port map ( Y=>nx11169, A=>d_arr_mul_7_29);
   ix5483 : oai21 port map ( Y=>nx5482, A0=>nx11171, A1=>nx10937, B0=>
      nx10757);
   ix11170 : inv01 port map ( Y=>nx11171, A=>d_arr_mul_7_30);
   ix5489 : oai21 port map ( Y=>nx5488, A0=>nx11173, A1=>nx10937, B0=>
      nx10757);
   ix11172 : inv01 port map ( Y=>nx11173, A=>d_arr_mul_7_31);
   ix5617 : oai21 port map ( Y=>nx5616, A0=>nx11175, A1=>nx11455, B0=>
      nx11427);
   ix11174 : inv01 port map ( Y=>nx11175, A=>d_arr_mul_6_15);
   ix5613 : nand02 port map ( Y=>nx10765, A0=>nx11503, A1=>d_arr_mux_6_31);
   ix5623 : oai21 port map ( Y=>nx5622, A0=>nx11177, A1=>nx11455, B0=>
      nx11427);
   ix11176 : inv01 port map ( Y=>nx11177, A=>d_arr_mul_6_16);
   ix5629 : oai21 port map ( Y=>nx5628, A0=>nx11179, A1=>nx11455, B0=>
      nx11427);
   ix11178 : inv01 port map ( Y=>nx11179, A=>d_arr_mul_6_17);
   ix5635 : oai21 port map ( Y=>nx5634, A0=>nx11181, A1=>nx11457, B0=>
      nx11427);
   ix11180 : inv01 port map ( Y=>nx11181, A=>d_arr_mul_6_18);
   ix5641 : oai21 port map ( Y=>nx5640, A0=>nx11183, A1=>nx11457, B0=>
      nx11427);
   ix11182 : inv01 port map ( Y=>nx11183, A=>d_arr_mul_6_19);
   ix5647 : oai21 port map ( Y=>nx5646, A0=>nx11185, A1=>nx11457, B0=>
      nx11427);
   ix11184 : inv01 port map ( Y=>nx11185, A=>d_arr_mul_6_20);
   ix5653 : oai21 port map ( Y=>nx5652, A0=>nx11187, A1=>nx11457, B0=>
      nx11427);
   ix11186 : inv01 port map ( Y=>nx11187, A=>d_arr_mul_6_21);
   ix5659 : oai21 port map ( Y=>nx5658, A0=>nx11189, A1=>nx11457, B0=>
      nx11429);
   ix11188 : inv01 port map ( Y=>nx11189, A=>d_arr_mul_6_22);
   ix5665 : oai21 port map ( Y=>nx5664, A0=>nx11191, A1=>nx11457, B0=>
      nx11429);
   ix11190 : inv01 port map ( Y=>nx11191, A=>d_arr_mul_6_23);
   ix5671 : oai21 port map ( Y=>nx5670, A0=>nx11193, A1=>nx11457, B0=>
      nx11429);
   ix11192 : inv01 port map ( Y=>nx11193, A=>d_arr_mul_6_24);
   ix5677 : oai21 port map ( Y=>nx5676, A0=>nx11195, A1=>nx11459, B0=>
      nx11429);
   ix11194 : inv01 port map ( Y=>nx11195, A=>d_arr_mul_6_25);
   ix5683 : oai21 port map ( Y=>nx5682, A0=>nx11197, A1=>nx11459, B0=>
      nx11429);
   ix11196 : inv01 port map ( Y=>nx11197, A=>d_arr_mul_6_26);
   ix5689 : oai21 port map ( Y=>nx5688, A0=>nx11199, A1=>nx11459, B0=>
      nx11429);
   ix11198 : inv01 port map ( Y=>nx11199, A=>d_arr_mul_6_27);
   ix5695 : oai21 port map ( Y=>nx5694, A0=>nx11201, A1=>nx11459, B0=>
      nx11429);
   ix11200 : inv01 port map ( Y=>nx11201, A=>d_arr_mul_6_28);
   ix5701 : oai21 port map ( Y=>nx5700, A0=>nx11203, A1=>nx11459, B0=>
      nx10765);
   ix11202 : inv01 port map ( Y=>nx11203, A=>d_arr_mul_6_29);
   ix5707 : oai21 port map ( Y=>nx5706, A0=>nx11205, A1=>nx11459, B0=>
      nx10765);
   ix11204 : inv01 port map ( Y=>nx11205, A=>d_arr_mul_6_30);
   ix5713 : oai21 port map ( Y=>nx5712, A0=>nx11207, A1=>nx11459, B0=>
      nx10765);
   ix11206 : inv01 port map ( Y=>nx11207, A=>d_arr_mul_6_31);
   ix5841 : oai21 port map ( Y=>nx5840, A0=>nx11209, A1=>nx11461, B0=>
      nx11431);
   ix11208 : inv01 port map ( Y=>nx11209, A=>d_arr_mul_5_15);
   ix5837 : nand02 port map ( Y=>nx10773, A0=>nx11503, A1=>d_arr_mux_5_31);
   ix5847 : oai21 port map ( Y=>nx5846, A0=>nx11211, A1=>nx11461, B0=>
      nx11431);
   ix11210 : inv01 port map ( Y=>nx11211, A=>d_arr_mul_5_16);
   ix5853 : oai21 port map ( Y=>nx5852, A0=>nx11213, A1=>nx11461, B0=>
      nx11431);
   ix11212 : inv01 port map ( Y=>nx11213, A=>d_arr_mul_5_17);
   ix5859 : oai21 port map ( Y=>nx5858, A0=>nx11215, A1=>nx11461, B0=>
      nx11431);
   ix11214 : inv01 port map ( Y=>nx11215, A=>d_arr_mul_5_18);
   ix5865 : oai21 port map ( Y=>nx5864, A0=>nx11217, A1=>nx11461, B0=>
      nx11431);
   ix11216 : inv01 port map ( Y=>nx11217, A=>d_arr_mul_5_19);
   ix5871 : oai21 port map ( Y=>nx5870, A0=>nx11219, A1=>nx11461, B0=>
      nx11431);
   ix11218 : inv01 port map ( Y=>nx11219, A=>d_arr_mul_5_20);
   ix5877 : oai21 port map ( Y=>nx5876, A0=>nx11221, A1=>nx11461, B0=>
      nx11431);
   ix11220 : inv01 port map ( Y=>nx11221, A=>d_arr_mul_5_21);
   ix5883 : oai21 port map ( Y=>nx5882, A0=>nx11223, A1=>nx10939, B0=>
      nx11433);
   ix11222 : inv01 port map ( Y=>nx11223, A=>d_arr_mul_5_22);
   ix5889 : oai21 port map ( Y=>nx5888, A0=>nx11225, A1=>nx10939, B0=>
      nx11433);
   ix11224 : inv01 port map ( Y=>nx11225, A=>d_arr_mul_5_23);
   ix5895 : oai21 port map ( Y=>nx5894, A0=>nx11227, A1=>nx10939, B0=>
      nx11433);
   ix11226 : inv01 port map ( Y=>nx11227, A=>d_arr_mul_5_24);
   ix5901 : oai21 port map ( Y=>nx5900, A0=>nx11229, A1=>nx10939, B0=>
      nx11433);
   ix11228 : inv01 port map ( Y=>nx11229, A=>d_arr_mul_5_25);
   ix5907 : oai21 port map ( Y=>nx5906, A0=>nx11231, A1=>nx10939, B0=>
      nx11433);
   ix11230 : inv01 port map ( Y=>nx11231, A=>d_arr_mul_5_26);
   ix5913 : oai21 port map ( Y=>nx5912, A0=>nx11233, A1=>nx10939, B0=>
      nx11433);
   ix11232 : inv01 port map ( Y=>nx11233, A=>d_arr_mul_5_27);
   ix5919 : oai21 port map ( Y=>nx5918, A0=>nx11235, A1=>nx10939, B0=>
      nx11433);
   ix11234 : inv01 port map ( Y=>nx11235, A=>d_arr_mul_5_28);
   ix5925 : oai21 port map ( Y=>nx5924, A0=>nx11237, A1=>nx10941, B0=>
      nx10773);
   ix11236 : inv01 port map ( Y=>nx11237, A=>d_arr_mul_5_29);
   ix5931 : oai21 port map ( Y=>nx5930, A0=>nx11239, A1=>nx10941, B0=>
      nx10773);
   ix11238 : inv01 port map ( Y=>nx11239, A=>d_arr_mul_5_30);
   ix5937 : oai21 port map ( Y=>nx5936, A0=>nx11241, A1=>nx10941, B0=>
      nx10773);
   ix11240 : inv01 port map ( Y=>nx11241, A=>d_arr_mul_5_31);
   ix11244 : inv02 port map ( Y=>nx11245, A=>nx11524);
   ix11246 : inv02 port map ( Y=>nx11247, A=>nx11524);
   ix11248 : inv02 port map ( Y=>nx11249, A=>nx11524);
   ix11250 : inv02 port map ( Y=>nx11251, A=>nx11524);
   ix11252 : inv02 port map ( Y=>nx11253, A=>nx11525);
   ix11254 : inv02 port map ( Y=>nx11255, A=>nx11525);
   ix11256 : inv02 port map ( Y=>nx11257, A=>nx11525);
   ix11258 : inv02 port map ( Y=>nx11259, A=>nx11479);
   ix11260 : inv02 port map ( Y=>nx11261, A=>nx11479);
   ix11262 : inv02 port map ( Y=>nx11263, A=>nx11479);
   ix11264 : inv02 port map ( Y=>nx11265, A=>nx11479);
   ix11266 : inv02 port map ( Y=>nx11267, A=>nx11479);
   ix11268 : inv02 port map ( Y=>nx11269, A=>nx11479);
   ix11270 : inv02 port map ( Y=>nx11271, A=>nx11479);
   ix11272 : inv02 port map ( Y=>nx11273, A=>nx11481);
   ix11274 : inv02 port map ( Y=>nx11275, A=>nx11481);
   ix11276 : inv02 port map ( Y=>nx11277, A=>nx11481);
   ix11278 : inv02 port map ( Y=>nx11279, A=>nx11481);
   ix11280 : inv02 port map ( Y=>nx11281, A=>nx11481);
   ix11282 : inv02 port map ( Y=>nx11283, A=>nx11481);
   ix11284 : inv02 port map ( Y=>nx11285, A=>nx11481);
   ix11286 : inv02 port map ( Y=>nx11287, A=>nx11483);
   ix11288 : inv02 port map ( Y=>nx11289, A=>nx11483);
   ix11290 : inv02 port map ( Y=>nx11291, A=>nx11483);
   ix11292 : inv02 port map ( Y=>nx11293, A=>nx11483);
   ix11294 : inv02 port map ( Y=>nx11295, A=>nx11483);
   ix11296 : inv02 port map ( Y=>nx11297, A=>nx11483);
   ix11298 : inv02 port map ( Y=>nx11299, A=>nx11483);
   ix11300 : inv02 port map ( Y=>nx11301, A=>nx11485);
   ix11302 : inv02 port map ( Y=>nx11303, A=>nx11485);
   ix11304 : inv02 port map ( Y=>nx11305, A=>nx11485);
   ix11306 : inv02 port map ( Y=>nx11307, A=>nx11485);
   ix11308 : inv02 port map ( Y=>nx11309, A=>nx11485);
   ix11310 : inv02 port map ( Y=>nx11311, A=>nx11485);
   ix11312 : inv02 port map ( Y=>nx11313, A=>nx11485);
   ix11314 : inv02 port map ( Y=>nx11315, A=>nx11487);
   ix11316 : inv02 port map ( Y=>nx11317, A=>nx11487);
   ix11318 : inv02 port map ( Y=>nx11319, A=>nx11487);
   ix11320 : inv02 port map ( Y=>nx11321, A=>nx11487);
   ix11322 : inv02 port map ( Y=>nx11323, A=>nx11487);
   ix11324 : inv02 port map ( Y=>nx11325, A=>nx11487);
   ix11326 : inv02 port map ( Y=>nx11327, A=>nx11487);
   ix11328 : inv02 port map ( Y=>nx11329, A=>nx11489);
   ix11330 : inv02 port map ( Y=>nx11331, A=>nx11489);
   ix11332 : inv02 port map ( Y=>nx11333, A=>nx11489);
   ix11334 : inv02 port map ( Y=>nx11335, A=>nx11489);
   ix11336 : inv02 port map ( Y=>nx11337, A=>nx11489);
   ix11338 : inv02 port map ( Y=>nx11339, A=>nx11489);
   ix11340 : inv02 port map ( Y=>nx11341, A=>nx11489);
   ix11342 : inv02 port map ( Y=>nx11343, A=>nx11491);
   ix11344 : inv02 port map ( Y=>nx11345, A=>nx11491);
   ix11346 : inv02 port map ( Y=>nx11347, A=>nx11491);
   ix11348 : inv02 port map ( Y=>nx11349, A=>nx11491);
   ix11350 : inv02 port map ( Y=>nx11351, A=>nx11491);
   ix11352 : inv02 port map ( Y=>nx11353, A=>nx11491);
   ix11354 : inv02 port map ( Y=>nx11355, A=>nx11491);
   ix11356 : inv02 port map ( Y=>nx11357, A=>nx11493);
   ix11358 : inv02 port map ( Y=>nx11359, A=>nx11493);
   ix11360 : inv02 port map ( Y=>nx11361, A=>nx11493);
   ix11362 : inv02 port map ( Y=>nx11363, A=>nx11493);
   ix11364 : inv02 port map ( Y=>nx11365, A=>nx11493);
   ix11366 : inv02 port map ( Y=>nx11367, A=>nx11493);
   ix11368 : inv02 port map ( Y=>nx11369, A=>nx11493);
   ix11370 : inv02 port map ( Y=>nx11371, A=>nx11495);
   ix11372 : inv02 port map ( Y=>nx11373, A=>nx11495);
   ix11374 : inv02 port map ( Y=>nx11375, A=>nx11495);
   ix11376 : inv02 port map ( Y=>nx11377, A=>nx11495);
   ix11378 : inv02 port map ( Y=>nx11379, A=>nx11495);
   ix11380 : inv02 port map ( Y=>nx11381, A=>nx11495);
   ix11382 : inv02 port map ( Y=>nx11383, A=>nx11495);
   ix11384 : inv02 port map ( Y=>nx11385, A=>nx11497);
   ix11386 : inv02 port map ( Y=>nx11387, A=>nx11497);
   ix11388 : inv02 port map ( Y=>nx11389, A=>nx11497);
   ix11390 : inv02 port map ( Y=>nx11391, A=>nx11497);
   ix11392 : inv02 port map ( Y=>nx11393, A=>nx11497);
   ix11394 : inv02 port map ( Y=>nx11395, A=>nx11497);
   ix11396 : inv02 port map ( Y=>nx11397, A=>nx11497);
   ix11398 : inv02 port map ( Y=>nx11399, A=>nx11499);
   ix11400 : inv02 port map ( Y=>nx11401, A=>nx11499);
   ix11402 : inv02 port map ( Y=>nx11403, A=>nx11499);
   ix11404 : inv02 port map ( Y=>nx11405, A=>nx11499);
   ix11406 : nand02 port map ( Y=>nx11407, A0=>nx11403, A1=>d_arr_mux_24_31
   );
   ix11408 : nand02 port map ( Y=>nx11409, A0=>nx11403, A1=>d_arr_mux_24_31
   );
   ix11410 : nand02 port map ( Y=>nx11411, A0=>nx11503, A1=>d_arr_mux_23_31
   );
   ix11412 : nand02 port map ( Y=>nx11413, A0=>nx11505, A1=>d_arr_mux_23_31
   );
   ix11414 : nand02 port map ( Y=>nx11415, A0=>nx11505, A1=>d_arr_mux_22_31
   );
   ix11416 : nand02 port map ( Y=>nx11417, A0=>nx11505, A1=>d_arr_mux_22_31
   );
   ix11418 : nand02 port map ( Y=>nx11419, A0=>nx11505, A1=>d_arr_mux_8_31);
   ix11420 : nand02 port map ( Y=>nx11421, A0=>nx11505, A1=>d_arr_mux_8_31);
   ix11422 : nand02 port map ( Y=>nx11423, A0=>nx11505, A1=>d_arr_mux_7_31);
   ix11424 : nand02 port map ( Y=>nx11425, A0=>nx11505, A1=>d_arr_mux_7_31);
   ix11426 : nand02 port map ( Y=>nx11427, A0=>nx11405, A1=>d_arr_mux_6_31);
   ix11428 : nand02 port map ( Y=>nx11429, A0=>nx11405, A1=>d_arr_mux_6_31);
   ix11430 : nand02 port map ( Y=>nx11431, A0=>nx11405, A1=>d_arr_mux_5_31);
   ix11432 : nand02 port map ( Y=>nx11433, A0=>nx11405, A1=>d_arr_mux_5_31);
   ix11434 : inv02 port map ( Y=>nx11435, A=>nx10985);
   ix11436 : inv02 port map ( Y=>nx11437, A=>nx10985);
   ix11438 : inv02 port map ( Y=>nx11439, A=>nx10985);
   ix11440 : inv02 port map ( Y=>nx11441, A=>nx10985);
   ix11442 : inv02 port map ( Y=>nx11443, A=>nx10985);
   ix11444 : inv02 port map ( Y=>nx11445, A=>nx11469);
   ix11446 : inv02 port map ( Y=>nx11447, A=>nx11469);
   ix11448 : inv02 port map ( Y=>nx11449, A=>nx11469);
   ix11450 : inv02 port map ( Y=>nx11451, A=>nx11469);
   ix11452 : inv02 port map ( Y=>nx11453, A=>nx11469);
   ix11454 : inv02 port map ( Y=>nx11455, A=>nx11469);
   ix11456 : inv02 port map ( Y=>nx11457, A=>nx11469);
   ix11458 : inv02 port map ( Y=>nx11459, A=>nx10987);
   ix11460 : inv02 port map ( Y=>nx11461, A=>nx10987);
   ix11462 : inv02 port map ( Y=>nx11463, A=>nx10987);
   ix11464 : inv02 port map ( Y=>nx11465, A=>nx10915);
   ix11466 : inv02 port map ( Y=>nx11467, A=>nx10915);
   ix11468 : inv02 port map ( Y=>nx11469, A=>nx10915);
   ix11470 : inv02 port map ( Y=>nx11471, A=>nx11511);
   ix11472 : inv02 port map ( Y=>nx11473, A=>nx11511);
   ix11474 : inv02 port map ( Y=>nx11475, A=>nx11511);
   ix11476 : inv02 port map ( Y=>nx11477, A=>sel_mux);
   ix11478 : inv02 port map ( Y=>nx11479, A=>nx11517);
   ix11480 : inv02 port map ( Y=>nx11481, A=>nx11517);
   ix11482 : inv02 port map ( Y=>nx11483, A=>nx11517);
   ix11484 : inv02 port map ( Y=>nx11485, A=>nx11517);
   ix11486 : inv02 port map ( Y=>nx11487, A=>nx11517);
   ix11488 : inv02 port map ( Y=>nx11489, A=>nx11517);
   ix11490 : inv02 port map ( Y=>nx11491, A=>nx11517);
   ix11492 : inv02 port map ( Y=>nx11493, A=>nx11519);
   ix11494 : inv02 port map ( Y=>nx11495, A=>nx11519);
   ix11496 : inv02 port map ( Y=>nx11497, A=>nx11519);
   ix11498 : inv02 port map ( Y=>nx11499, A=>nx11519);
   ix11500 : inv02 port map ( Y=>nx11501, A=>nx11499);
   ix11502 : inv02 port map ( Y=>nx11503, A=>nx11499);
   ix11504 : inv02 port map ( Y=>nx11505, A=>nx11499);
   ix11510 : inv01 port map ( Y=>nx11511, A=>nx10915);
   ix11516 : inv02 port map ( Y=>nx11517, A=>nx11525);
   ix11518 : inv02 port map ( Y=>nx11519, A=>nx11525);
   ix11526 : buf16 port map ( Y=>nx11524, A=>nx11477);
   ix11527 : buf16 port map ( Y=>nx11525, A=>nx11477);
end Behavioral_unfold_3297_0 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity MuxLayer is
   port (
      img_data_0_31 : IN std_logic ;
      img_data_0_30 : IN std_logic ;
      img_data_0_29 : IN std_logic ;
      img_data_0_28 : IN std_logic ;
      img_data_0_27 : IN std_logic ;
      img_data_0_26 : IN std_logic ;
      img_data_0_25 : IN std_logic ;
      img_data_0_24 : IN std_logic ;
      img_data_0_23 : IN std_logic ;
      img_data_0_22 : IN std_logic ;
      img_data_0_21 : IN std_logic ;
      img_data_0_20 : IN std_logic ;
      img_data_0_19 : IN std_logic ;
      img_data_0_18 : IN std_logic ;
      img_data_0_17 : IN std_logic ;
      img_data_0_16 : IN std_logic ;
      img_data_0_15 : IN std_logic ;
      img_data_0_14 : IN std_logic ;
      img_data_0_13 : IN std_logic ;
      img_data_0_12 : IN std_logic ;
      img_data_0_11 : IN std_logic ;
      img_data_0_10 : IN std_logic ;
      img_data_0_9 : IN std_logic ;
      img_data_0_8 : IN std_logic ;
      img_data_0_7 : IN std_logic ;
      img_data_0_6 : IN std_logic ;
      img_data_0_5 : IN std_logic ;
      img_data_0_4 : IN std_logic ;
      img_data_0_3 : IN std_logic ;
      img_data_0_2 : IN std_logic ;
      img_data_0_1 : IN std_logic ;
      img_data_0_0 : IN std_logic ;
      img_data_1_31 : IN std_logic ;
      img_data_1_30 : IN std_logic ;
      img_data_1_29 : IN std_logic ;
      img_data_1_28 : IN std_logic ;
      img_data_1_27 : IN std_logic ;
      img_data_1_26 : IN std_logic ;
      img_data_1_25 : IN std_logic ;
      img_data_1_24 : IN std_logic ;
      img_data_1_23 : IN std_logic ;
      img_data_1_22 : IN std_logic ;
      img_data_1_21 : IN std_logic ;
      img_data_1_20 : IN std_logic ;
      img_data_1_19 : IN std_logic ;
      img_data_1_18 : IN std_logic ;
      img_data_1_17 : IN std_logic ;
      img_data_1_16 : IN std_logic ;
      img_data_1_15 : IN std_logic ;
      img_data_1_14 : IN std_logic ;
      img_data_1_13 : IN std_logic ;
      img_data_1_12 : IN std_logic ;
      img_data_1_11 : IN std_logic ;
      img_data_1_10 : IN std_logic ;
      img_data_1_9 : IN std_logic ;
      img_data_1_8 : IN std_logic ;
      img_data_1_7 : IN std_logic ;
      img_data_1_6 : IN std_logic ;
      img_data_1_5 : IN std_logic ;
      img_data_1_4 : IN std_logic ;
      img_data_1_3 : IN std_logic ;
      img_data_1_2 : IN std_logic ;
      img_data_1_1 : IN std_logic ;
      img_data_1_0 : IN std_logic ;
      img_data_2_31 : IN std_logic ;
      img_data_2_30 : IN std_logic ;
      img_data_2_29 : IN std_logic ;
      img_data_2_28 : IN std_logic ;
      img_data_2_27 : IN std_logic ;
      img_data_2_26 : IN std_logic ;
      img_data_2_25 : IN std_logic ;
      img_data_2_24 : IN std_logic ;
      img_data_2_23 : IN std_logic ;
      img_data_2_22 : IN std_logic ;
      img_data_2_21 : IN std_logic ;
      img_data_2_20 : IN std_logic ;
      img_data_2_19 : IN std_logic ;
      img_data_2_18 : IN std_logic ;
      img_data_2_17 : IN std_logic ;
      img_data_2_16 : IN std_logic ;
      img_data_2_15 : IN std_logic ;
      img_data_2_14 : IN std_logic ;
      img_data_2_13 : IN std_logic ;
      img_data_2_12 : IN std_logic ;
      img_data_2_11 : IN std_logic ;
      img_data_2_10 : IN std_logic ;
      img_data_2_9 : IN std_logic ;
      img_data_2_8 : IN std_logic ;
      img_data_2_7 : IN std_logic ;
      img_data_2_6 : IN std_logic ;
      img_data_2_5 : IN std_logic ;
      img_data_2_4 : IN std_logic ;
      img_data_2_3 : IN std_logic ;
      img_data_2_2 : IN std_logic ;
      img_data_2_1 : IN std_logic ;
      img_data_2_0 : IN std_logic ;
      img_data_3_31 : IN std_logic ;
      img_data_3_30 : IN std_logic ;
      img_data_3_29 : IN std_logic ;
      img_data_3_28 : IN std_logic ;
      img_data_3_27 : IN std_logic ;
      img_data_3_26 : IN std_logic ;
      img_data_3_25 : IN std_logic ;
      img_data_3_24 : IN std_logic ;
      img_data_3_23 : IN std_logic ;
      img_data_3_22 : IN std_logic ;
      img_data_3_21 : IN std_logic ;
      img_data_3_20 : IN std_logic ;
      img_data_3_19 : IN std_logic ;
      img_data_3_18 : IN std_logic ;
      img_data_3_17 : IN std_logic ;
      img_data_3_16 : IN std_logic ;
      img_data_3_15 : IN std_logic ;
      img_data_3_14 : IN std_logic ;
      img_data_3_13 : IN std_logic ;
      img_data_3_12 : IN std_logic ;
      img_data_3_11 : IN std_logic ;
      img_data_3_10 : IN std_logic ;
      img_data_3_9 : IN std_logic ;
      img_data_3_8 : IN std_logic ;
      img_data_3_7 : IN std_logic ;
      img_data_3_6 : IN std_logic ;
      img_data_3_5 : IN std_logic ;
      img_data_3_4 : IN std_logic ;
      img_data_3_3 : IN std_logic ;
      img_data_3_2 : IN std_logic ;
      img_data_3_1 : IN std_logic ;
      img_data_3_0 : IN std_logic ;
      img_data_4_31 : IN std_logic ;
      img_data_4_30 : IN std_logic ;
      img_data_4_29 : IN std_logic ;
      img_data_4_28 : IN std_logic ;
      img_data_4_27 : IN std_logic ;
      img_data_4_26 : IN std_logic ;
      img_data_4_25 : IN std_logic ;
      img_data_4_24 : IN std_logic ;
      img_data_4_23 : IN std_logic ;
      img_data_4_22 : IN std_logic ;
      img_data_4_21 : IN std_logic ;
      img_data_4_20 : IN std_logic ;
      img_data_4_19 : IN std_logic ;
      img_data_4_18 : IN std_logic ;
      img_data_4_17 : IN std_logic ;
      img_data_4_16 : IN std_logic ;
      img_data_4_15 : IN std_logic ;
      img_data_4_14 : IN std_logic ;
      img_data_4_13 : IN std_logic ;
      img_data_4_12 : IN std_logic ;
      img_data_4_11 : IN std_logic ;
      img_data_4_10 : IN std_logic ;
      img_data_4_9 : IN std_logic ;
      img_data_4_8 : IN std_logic ;
      img_data_4_7 : IN std_logic ;
      img_data_4_6 : IN std_logic ;
      img_data_4_5 : IN std_logic ;
      img_data_4_4 : IN std_logic ;
      img_data_4_3 : IN std_logic ;
      img_data_4_2 : IN std_logic ;
      img_data_4_1 : IN std_logic ;
      img_data_4_0 : IN std_logic ;
      img_data_5_31 : IN std_logic ;
      img_data_5_30 : IN std_logic ;
      img_data_5_29 : IN std_logic ;
      img_data_5_28 : IN std_logic ;
      img_data_5_27 : IN std_logic ;
      img_data_5_26 : IN std_logic ;
      img_data_5_25 : IN std_logic ;
      img_data_5_24 : IN std_logic ;
      img_data_5_23 : IN std_logic ;
      img_data_5_22 : IN std_logic ;
      img_data_5_21 : IN std_logic ;
      img_data_5_20 : IN std_logic ;
      img_data_5_19 : IN std_logic ;
      img_data_5_18 : IN std_logic ;
      img_data_5_17 : IN std_logic ;
      img_data_5_16 : IN std_logic ;
      img_data_5_15 : IN std_logic ;
      img_data_5_14 : IN std_logic ;
      img_data_5_13 : IN std_logic ;
      img_data_5_12 : IN std_logic ;
      img_data_5_11 : IN std_logic ;
      img_data_5_10 : IN std_logic ;
      img_data_5_9 : IN std_logic ;
      img_data_5_8 : IN std_logic ;
      img_data_5_7 : IN std_logic ;
      img_data_5_6 : IN std_logic ;
      img_data_5_5 : IN std_logic ;
      img_data_5_4 : IN std_logic ;
      img_data_5_3 : IN std_logic ;
      img_data_5_2 : IN std_logic ;
      img_data_5_1 : IN std_logic ;
      img_data_5_0 : IN std_logic ;
      img_data_6_31 : IN std_logic ;
      img_data_6_30 : IN std_logic ;
      img_data_6_29 : IN std_logic ;
      img_data_6_28 : IN std_logic ;
      img_data_6_27 : IN std_logic ;
      img_data_6_26 : IN std_logic ;
      img_data_6_25 : IN std_logic ;
      img_data_6_24 : IN std_logic ;
      img_data_6_23 : IN std_logic ;
      img_data_6_22 : IN std_logic ;
      img_data_6_21 : IN std_logic ;
      img_data_6_20 : IN std_logic ;
      img_data_6_19 : IN std_logic ;
      img_data_6_18 : IN std_logic ;
      img_data_6_17 : IN std_logic ;
      img_data_6_16 : IN std_logic ;
      img_data_6_15 : IN std_logic ;
      img_data_6_14 : IN std_logic ;
      img_data_6_13 : IN std_logic ;
      img_data_6_12 : IN std_logic ;
      img_data_6_11 : IN std_logic ;
      img_data_6_10 : IN std_logic ;
      img_data_6_9 : IN std_logic ;
      img_data_6_8 : IN std_logic ;
      img_data_6_7 : IN std_logic ;
      img_data_6_6 : IN std_logic ;
      img_data_6_5 : IN std_logic ;
      img_data_6_4 : IN std_logic ;
      img_data_6_3 : IN std_logic ;
      img_data_6_2 : IN std_logic ;
      img_data_6_1 : IN std_logic ;
      img_data_6_0 : IN std_logic ;
      img_data_7_31 : IN std_logic ;
      img_data_7_30 : IN std_logic ;
      img_data_7_29 : IN std_logic ;
      img_data_7_28 : IN std_logic ;
      img_data_7_27 : IN std_logic ;
      img_data_7_26 : IN std_logic ;
      img_data_7_25 : IN std_logic ;
      img_data_7_24 : IN std_logic ;
      img_data_7_23 : IN std_logic ;
      img_data_7_22 : IN std_logic ;
      img_data_7_21 : IN std_logic ;
      img_data_7_20 : IN std_logic ;
      img_data_7_19 : IN std_logic ;
      img_data_7_18 : IN std_logic ;
      img_data_7_17 : IN std_logic ;
      img_data_7_16 : IN std_logic ;
      img_data_7_15 : IN std_logic ;
      img_data_7_14 : IN std_logic ;
      img_data_7_13 : IN std_logic ;
      img_data_7_12 : IN std_logic ;
      img_data_7_11 : IN std_logic ;
      img_data_7_10 : IN std_logic ;
      img_data_7_9 : IN std_logic ;
      img_data_7_8 : IN std_logic ;
      img_data_7_7 : IN std_logic ;
      img_data_7_6 : IN std_logic ;
      img_data_7_5 : IN std_logic ;
      img_data_7_4 : IN std_logic ;
      img_data_7_3 : IN std_logic ;
      img_data_7_2 : IN std_logic ;
      img_data_7_1 : IN std_logic ;
      img_data_7_0 : IN std_logic ;
      img_data_8_31 : IN std_logic ;
      img_data_8_30 : IN std_logic ;
      img_data_8_29 : IN std_logic ;
      img_data_8_28 : IN std_logic ;
      img_data_8_27 : IN std_logic ;
      img_data_8_26 : IN std_logic ;
      img_data_8_25 : IN std_logic ;
      img_data_8_24 : IN std_logic ;
      img_data_8_23 : IN std_logic ;
      img_data_8_22 : IN std_logic ;
      img_data_8_21 : IN std_logic ;
      img_data_8_20 : IN std_logic ;
      img_data_8_19 : IN std_logic ;
      img_data_8_18 : IN std_logic ;
      img_data_8_17 : IN std_logic ;
      img_data_8_16 : IN std_logic ;
      img_data_8_15 : IN std_logic ;
      img_data_8_14 : IN std_logic ;
      img_data_8_13 : IN std_logic ;
      img_data_8_12 : IN std_logic ;
      img_data_8_11 : IN std_logic ;
      img_data_8_10 : IN std_logic ;
      img_data_8_9 : IN std_logic ;
      img_data_8_8 : IN std_logic ;
      img_data_8_7 : IN std_logic ;
      img_data_8_6 : IN std_logic ;
      img_data_8_5 : IN std_logic ;
      img_data_8_4 : IN std_logic ;
      img_data_8_3 : IN std_logic ;
      img_data_8_2 : IN std_logic ;
      img_data_8_1 : IN std_logic ;
      img_data_8_0 : IN std_logic ;
      img_data_9_31 : IN std_logic ;
      img_data_9_30 : IN std_logic ;
      img_data_9_29 : IN std_logic ;
      img_data_9_28 : IN std_logic ;
      img_data_9_27 : IN std_logic ;
      img_data_9_26 : IN std_logic ;
      img_data_9_25 : IN std_logic ;
      img_data_9_24 : IN std_logic ;
      img_data_9_23 : IN std_logic ;
      img_data_9_22 : IN std_logic ;
      img_data_9_21 : IN std_logic ;
      img_data_9_20 : IN std_logic ;
      img_data_9_19 : IN std_logic ;
      img_data_9_18 : IN std_logic ;
      img_data_9_17 : IN std_logic ;
      img_data_9_16 : IN std_logic ;
      img_data_9_15 : IN std_logic ;
      img_data_9_14 : IN std_logic ;
      img_data_9_13 : IN std_logic ;
      img_data_9_12 : IN std_logic ;
      img_data_9_11 : IN std_logic ;
      img_data_9_10 : IN std_logic ;
      img_data_9_9 : IN std_logic ;
      img_data_9_8 : IN std_logic ;
      img_data_9_7 : IN std_logic ;
      img_data_9_6 : IN std_logic ;
      img_data_9_5 : IN std_logic ;
      img_data_9_4 : IN std_logic ;
      img_data_9_3 : IN std_logic ;
      img_data_9_2 : IN std_logic ;
      img_data_9_1 : IN std_logic ;
      img_data_9_0 : IN std_logic ;
      img_data_10_31 : IN std_logic ;
      img_data_10_30 : IN std_logic ;
      img_data_10_29 : IN std_logic ;
      img_data_10_28 : IN std_logic ;
      img_data_10_27 : IN std_logic ;
      img_data_10_26 : IN std_logic ;
      img_data_10_25 : IN std_logic ;
      img_data_10_24 : IN std_logic ;
      img_data_10_23 : IN std_logic ;
      img_data_10_22 : IN std_logic ;
      img_data_10_21 : IN std_logic ;
      img_data_10_20 : IN std_logic ;
      img_data_10_19 : IN std_logic ;
      img_data_10_18 : IN std_logic ;
      img_data_10_17 : IN std_logic ;
      img_data_10_16 : IN std_logic ;
      img_data_10_15 : IN std_logic ;
      img_data_10_14 : IN std_logic ;
      img_data_10_13 : IN std_logic ;
      img_data_10_12 : IN std_logic ;
      img_data_10_11 : IN std_logic ;
      img_data_10_10 : IN std_logic ;
      img_data_10_9 : IN std_logic ;
      img_data_10_8 : IN std_logic ;
      img_data_10_7 : IN std_logic ;
      img_data_10_6 : IN std_logic ;
      img_data_10_5 : IN std_logic ;
      img_data_10_4 : IN std_logic ;
      img_data_10_3 : IN std_logic ;
      img_data_10_2 : IN std_logic ;
      img_data_10_1 : IN std_logic ;
      img_data_10_0 : IN std_logic ;
      img_data_11_31 : IN std_logic ;
      img_data_11_30 : IN std_logic ;
      img_data_11_29 : IN std_logic ;
      img_data_11_28 : IN std_logic ;
      img_data_11_27 : IN std_logic ;
      img_data_11_26 : IN std_logic ;
      img_data_11_25 : IN std_logic ;
      img_data_11_24 : IN std_logic ;
      img_data_11_23 : IN std_logic ;
      img_data_11_22 : IN std_logic ;
      img_data_11_21 : IN std_logic ;
      img_data_11_20 : IN std_logic ;
      img_data_11_19 : IN std_logic ;
      img_data_11_18 : IN std_logic ;
      img_data_11_17 : IN std_logic ;
      img_data_11_16 : IN std_logic ;
      img_data_11_15 : IN std_logic ;
      img_data_11_14 : IN std_logic ;
      img_data_11_13 : IN std_logic ;
      img_data_11_12 : IN std_logic ;
      img_data_11_11 : IN std_logic ;
      img_data_11_10 : IN std_logic ;
      img_data_11_9 : IN std_logic ;
      img_data_11_8 : IN std_logic ;
      img_data_11_7 : IN std_logic ;
      img_data_11_6 : IN std_logic ;
      img_data_11_5 : IN std_logic ;
      img_data_11_4 : IN std_logic ;
      img_data_11_3 : IN std_logic ;
      img_data_11_2 : IN std_logic ;
      img_data_11_1 : IN std_logic ;
      img_data_11_0 : IN std_logic ;
      img_data_12_31 : IN std_logic ;
      img_data_12_30 : IN std_logic ;
      img_data_12_29 : IN std_logic ;
      img_data_12_28 : IN std_logic ;
      img_data_12_27 : IN std_logic ;
      img_data_12_26 : IN std_logic ;
      img_data_12_25 : IN std_logic ;
      img_data_12_24 : IN std_logic ;
      img_data_12_23 : IN std_logic ;
      img_data_12_22 : IN std_logic ;
      img_data_12_21 : IN std_logic ;
      img_data_12_20 : IN std_logic ;
      img_data_12_19 : IN std_logic ;
      img_data_12_18 : IN std_logic ;
      img_data_12_17 : IN std_logic ;
      img_data_12_16 : IN std_logic ;
      img_data_12_15 : IN std_logic ;
      img_data_12_14 : IN std_logic ;
      img_data_12_13 : IN std_logic ;
      img_data_12_12 : IN std_logic ;
      img_data_12_11 : IN std_logic ;
      img_data_12_10 : IN std_logic ;
      img_data_12_9 : IN std_logic ;
      img_data_12_8 : IN std_logic ;
      img_data_12_7 : IN std_logic ;
      img_data_12_6 : IN std_logic ;
      img_data_12_5 : IN std_logic ;
      img_data_12_4 : IN std_logic ;
      img_data_12_3 : IN std_logic ;
      img_data_12_2 : IN std_logic ;
      img_data_12_1 : IN std_logic ;
      img_data_12_0 : IN std_logic ;
      img_data_13_31 : IN std_logic ;
      img_data_13_30 : IN std_logic ;
      img_data_13_29 : IN std_logic ;
      img_data_13_28 : IN std_logic ;
      img_data_13_27 : IN std_logic ;
      img_data_13_26 : IN std_logic ;
      img_data_13_25 : IN std_logic ;
      img_data_13_24 : IN std_logic ;
      img_data_13_23 : IN std_logic ;
      img_data_13_22 : IN std_logic ;
      img_data_13_21 : IN std_logic ;
      img_data_13_20 : IN std_logic ;
      img_data_13_19 : IN std_logic ;
      img_data_13_18 : IN std_logic ;
      img_data_13_17 : IN std_logic ;
      img_data_13_16 : IN std_logic ;
      img_data_13_15 : IN std_logic ;
      img_data_13_14 : IN std_logic ;
      img_data_13_13 : IN std_logic ;
      img_data_13_12 : IN std_logic ;
      img_data_13_11 : IN std_logic ;
      img_data_13_10 : IN std_logic ;
      img_data_13_9 : IN std_logic ;
      img_data_13_8 : IN std_logic ;
      img_data_13_7 : IN std_logic ;
      img_data_13_6 : IN std_logic ;
      img_data_13_5 : IN std_logic ;
      img_data_13_4 : IN std_logic ;
      img_data_13_3 : IN std_logic ;
      img_data_13_2 : IN std_logic ;
      img_data_13_1 : IN std_logic ;
      img_data_13_0 : IN std_logic ;
      img_data_14_31 : IN std_logic ;
      img_data_14_30 : IN std_logic ;
      img_data_14_29 : IN std_logic ;
      img_data_14_28 : IN std_logic ;
      img_data_14_27 : IN std_logic ;
      img_data_14_26 : IN std_logic ;
      img_data_14_25 : IN std_logic ;
      img_data_14_24 : IN std_logic ;
      img_data_14_23 : IN std_logic ;
      img_data_14_22 : IN std_logic ;
      img_data_14_21 : IN std_logic ;
      img_data_14_20 : IN std_logic ;
      img_data_14_19 : IN std_logic ;
      img_data_14_18 : IN std_logic ;
      img_data_14_17 : IN std_logic ;
      img_data_14_16 : IN std_logic ;
      img_data_14_15 : IN std_logic ;
      img_data_14_14 : IN std_logic ;
      img_data_14_13 : IN std_logic ;
      img_data_14_12 : IN std_logic ;
      img_data_14_11 : IN std_logic ;
      img_data_14_10 : IN std_logic ;
      img_data_14_9 : IN std_logic ;
      img_data_14_8 : IN std_logic ;
      img_data_14_7 : IN std_logic ;
      img_data_14_6 : IN std_logic ;
      img_data_14_5 : IN std_logic ;
      img_data_14_4 : IN std_logic ;
      img_data_14_3 : IN std_logic ;
      img_data_14_2 : IN std_logic ;
      img_data_14_1 : IN std_logic ;
      img_data_14_0 : IN std_logic ;
      img_data_15_31 : IN std_logic ;
      img_data_15_30 : IN std_logic ;
      img_data_15_29 : IN std_logic ;
      img_data_15_28 : IN std_logic ;
      img_data_15_27 : IN std_logic ;
      img_data_15_26 : IN std_logic ;
      img_data_15_25 : IN std_logic ;
      img_data_15_24 : IN std_logic ;
      img_data_15_23 : IN std_logic ;
      img_data_15_22 : IN std_logic ;
      img_data_15_21 : IN std_logic ;
      img_data_15_20 : IN std_logic ;
      img_data_15_19 : IN std_logic ;
      img_data_15_18 : IN std_logic ;
      img_data_15_17 : IN std_logic ;
      img_data_15_16 : IN std_logic ;
      img_data_15_15 : IN std_logic ;
      img_data_15_14 : IN std_logic ;
      img_data_15_13 : IN std_logic ;
      img_data_15_12 : IN std_logic ;
      img_data_15_11 : IN std_logic ;
      img_data_15_10 : IN std_logic ;
      img_data_15_9 : IN std_logic ;
      img_data_15_8 : IN std_logic ;
      img_data_15_7 : IN std_logic ;
      img_data_15_6 : IN std_logic ;
      img_data_15_5 : IN std_logic ;
      img_data_15_4 : IN std_logic ;
      img_data_15_3 : IN std_logic ;
      img_data_15_2 : IN std_logic ;
      img_data_15_1 : IN std_logic ;
      img_data_15_0 : IN std_logic ;
      img_data_16_31 : IN std_logic ;
      img_data_16_30 : IN std_logic ;
      img_data_16_29 : IN std_logic ;
      img_data_16_28 : IN std_logic ;
      img_data_16_27 : IN std_logic ;
      img_data_16_26 : IN std_logic ;
      img_data_16_25 : IN std_logic ;
      img_data_16_24 : IN std_logic ;
      img_data_16_23 : IN std_logic ;
      img_data_16_22 : IN std_logic ;
      img_data_16_21 : IN std_logic ;
      img_data_16_20 : IN std_logic ;
      img_data_16_19 : IN std_logic ;
      img_data_16_18 : IN std_logic ;
      img_data_16_17 : IN std_logic ;
      img_data_16_16 : IN std_logic ;
      img_data_16_15 : IN std_logic ;
      img_data_16_14 : IN std_logic ;
      img_data_16_13 : IN std_logic ;
      img_data_16_12 : IN std_logic ;
      img_data_16_11 : IN std_logic ;
      img_data_16_10 : IN std_logic ;
      img_data_16_9 : IN std_logic ;
      img_data_16_8 : IN std_logic ;
      img_data_16_7 : IN std_logic ;
      img_data_16_6 : IN std_logic ;
      img_data_16_5 : IN std_logic ;
      img_data_16_4 : IN std_logic ;
      img_data_16_3 : IN std_logic ;
      img_data_16_2 : IN std_logic ;
      img_data_16_1 : IN std_logic ;
      img_data_16_0 : IN std_logic ;
      img_data_17_31 : IN std_logic ;
      img_data_17_30 : IN std_logic ;
      img_data_17_29 : IN std_logic ;
      img_data_17_28 : IN std_logic ;
      img_data_17_27 : IN std_logic ;
      img_data_17_26 : IN std_logic ;
      img_data_17_25 : IN std_logic ;
      img_data_17_24 : IN std_logic ;
      img_data_17_23 : IN std_logic ;
      img_data_17_22 : IN std_logic ;
      img_data_17_21 : IN std_logic ;
      img_data_17_20 : IN std_logic ;
      img_data_17_19 : IN std_logic ;
      img_data_17_18 : IN std_logic ;
      img_data_17_17 : IN std_logic ;
      img_data_17_16 : IN std_logic ;
      img_data_17_15 : IN std_logic ;
      img_data_17_14 : IN std_logic ;
      img_data_17_13 : IN std_logic ;
      img_data_17_12 : IN std_logic ;
      img_data_17_11 : IN std_logic ;
      img_data_17_10 : IN std_logic ;
      img_data_17_9 : IN std_logic ;
      img_data_17_8 : IN std_logic ;
      img_data_17_7 : IN std_logic ;
      img_data_17_6 : IN std_logic ;
      img_data_17_5 : IN std_logic ;
      img_data_17_4 : IN std_logic ;
      img_data_17_3 : IN std_logic ;
      img_data_17_2 : IN std_logic ;
      img_data_17_1 : IN std_logic ;
      img_data_17_0 : IN std_logic ;
      img_data_18_31 : IN std_logic ;
      img_data_18_30 : IN std_logic ;
      img_data_18_29 : IN std_logic ;
      img_data_18_28 : IN std_logic ;
      img_data_18_27 : IN std_logic ;
      img_data_18_26 : IN std_logic ;
      img_data_18_25 : IN std_logic ;
      img_data_18_24 : IN std_logic ;
      img_data_18_23 : IN std_logic ;
      img_data_18_22 : IN std_logic ;
      img_data_18_21 : IN std_logic ;
      img_data_18_20 : IN std_logic ;
      img_data_18_19 : IN std_logic ;
      img_data_18_18 : IN std_logic ;
      img_data_18_17 : IN std_logic ;
      img_data_18_16 : IN std_logic ;
      img_data_18_15 : IN std_logic ;
      img_data_18_14 : IN std_logic ;
      img_data_18_13 : IN std_logic ;
      img_data_18_12 : IN std_logic ;
      img_data_18_11 : IN std_logic ;
      img_data_18_10 : IN std_logic ;
      img_data_18_9 : IN std_logic ;
      img_data_18_8 : IN std_logic ;
      img_data_18_7 : IN std_logic ;
      img_data_18_6 : IN std_logic ;
      img_data_18_5 : IN std_logic ;
      img_data_18_4 : IN std_logic ;
      img_data_18_3 : IN std_logic ;
      img_data_18_2 : IN std_logic ;
      img_data_18_1 : IN std_logic ;
      img_data_18_0 : IN std_logic ;
      img_data_19_31 : IN std_logic ;
      img_data_19_30 : IN std_logic ;
      img_data_19_29 : IN std_logic ;
      img_data_19_28 : IN std_logic ;
      img_data_19_27 : IN std_logic ;
      img_data_19_26 : IN std_logic ;
      img_data_19_25 : IN std_logic ;
      img_data_19_24 : IN std_logic ;
      img_data_19_23 : IN std_logic ;
      img_data_19_22 : IN std_logic ;
      img_data_19_21 : IN std_logic ;
      img_data_19_20 : IN std_logic ;
      img_data_19_19 : IN std_logic ;
      img_data_19_18 : IN std_logic ;
      img_data_19_17 : IN std_logic ;
      img_data_19_16 : IN std_logic ;
      img_data_19_15 : IN std_logic ;
      img_data_19_14 : IN std_logic ;
      img_data_19_13 : IN std_logic ;
      img_data_19_12 : IN std_logic ;
      img_data_19_11 : IN std_logic ;
      img_data_19_10 : IN std_logic ;
      img_data_19_9 : IN std_logic ;
      img_data_19_8 : IN std_logic ;
      img_data_19_7 : IN std_logic ;
      img_data_19_6 : IN std_logic ;
      img_data_19_5 : IN std_logic ;
      img_data_19_4 : IN std_logic ;
      img_data_19_3 : IN std_logic ;
      img_data_19_2 : IN std_logic ;
      img_data_19_1 : IN std_logic ;
      img_data_19_0 : IN std_logic ;
      img_data_20_31 : IN std_logic ;
      img_data_20_30 : IN std_logic ;
      img_data_20_29 : IN std_logic ;
      img_data_20_28 : IN std_logic ;
      img_data_20_27 : IN std_logic ;
      img_data_20_26 : IN std_logic ;
      img_data_20_25 : IN std_logic ;
      img_data_20_24 : IN std_logic ;
      img_data_20_23 : IN std_logic ;
      img_data_20_22 : IN std_logic ;
      img_data_20_21 : IN std_logic ;
      img_data_20_20 : IN std_logic ;
      img_data_20_19 : IN std_logic ;
      img_data_20_18 : IN std_logic ;
      img_data_20_17 : IN std_logic ;
      img_data_20_16 : IN std_logic ;
      img_data_20_15 : IN std_logic ;
      img_data_20_14 : IN std_logic ;
      img_data_20_13 : IN std_logic ;
      img_data_20_12 : IN std_logic ;
      img_data_20_11 : IN std_logic ;
      img_data_20_10 : IN std_logic ;
      img_data_20_9 : IN std_logic ;
      img_data_20_8 : IN std_logic ;
      img_data_20_7 : IN std_logic ;
      img_data_20_6 : IN std_logic ;
      img_data_20_5 : IN std_logic ;
      img_data_20_4 : IN std_logic ;
      img_data_20_3 : IN std_logic ;
      img_data_20_2 : IN std_logic ;
      img_data_20_1 : IN std_logic ;
      img_data_20_0 : IN std_logic ;
      img_data_21_31 : IN std_logic ;
      img_data_21_30 : IN std_logic ;
      img_data_21_29 : IN std_logic ;
      img_data_21_28 : IN std_logic ;
      img_data_21_27 : IN std_logic ;
      img_data_21_26 : IN std_logic ;
      img_data_21_25 : IN std_logic ;
      img_data_21_24 : IN std_logic ;
      img_data_21_23 : IN std_logic ;
      img_data_21_22 : IN std_logic ;
      img_data_21_21 : IN std_logic ;
      img_data_21_20 : IN std_logic ;
      img_data_21_19 : IN std_logic ;
      img_data_21_18 : IN std_logic ;
      img_data_21_17 : IN std_logic ;
      img_data_21_16 : IN std_logic ;
      img_data_21_15 : IN std_logic ;
      img_data_21_14 : IN std_logic ;
      img_data_21_13 : IN std_logic ;
      img_data_21_12 : IN std_logic ;
      img_data_21_11 : IN std_logic ;
      img_data_21_10 : IN std_logic ;
      img_data_21_9 : IN std_logic ;
      img_data_21_8 : IN std_logic ;
      img_data_21_7 : IN std_logic ;
      img_data_21_6 : IN std_logic ;
      img_data_21_5 : IN std_logic ;
      img_data_21_4 : IN std_logic ;
      img_data_21_3 : IN std_logic ;
      img_data_21_2 : IN std_logic ;
      img_data_21_1 : IN std_logic ;
      img_data_21_0 : IN std_logic ;
      img_data_22_31 : IN std_logic ;
      img_data_22_30 : IN std_logic ;
      img_data_22_29 : IN std_logic ;
      img_data_22_28 : IN std_logic ;
      img_data_22_27 : IN std_logic ;
      img_data_22_26 : IN std_logic ;
      img_data_22_25 : IN std_logic ;
      img_data_22_24 : IN std_logic ;
      img_data_22_23 : IN std_logic ;
      img_data_22_22 : IN std_logic ;
      img_data_22_21 : IN std_logic ;
      img_data_22_20 : IN std_logic ;
      img_data_22_19 : IN std_logic ;
      img_data_22_18 : IN std_logic ;
      img_data_22_17 : IN std_logic ;
      img_data_22_16 : IN std_logic ;
      img_data_22_15 : IN std_logic ;
      img_data_22_14 : IN std_logic ;
      img_data_22_13 : IN std_logic ;
      img_data_22_12 : IN std_logic ;
      img_data_22_11 : IN std_logic ;
      img_data_22_10 : IN std_logic ;
      img_data_22_9 : IN std_logic ;
      img_data_22_8 : IN std_logic ;
      img_data_22_7 : IN std_logic ;
      img_data_22_6 : IN std_logic ;
      img_data_22_5 : IN std_logic ;
      img_data_22_4 : IN std_logic ;
      img_data_22_3 : IN std_logic ;
      img_data_22_2 : IN std_logic ;
      img_data_22_1 : IN std_logic ;
      img_data_22_0 : IN std_logic ;
      img_data_23_31 : IN std_logic ;
      img_data_23_30 : IN std_logic ;
      img_data_23_29 : IN std_logic ;
      img_data_23_28 : IN std_logic ;
      img_data_23_27 : IN std_logic ;
      img_data_23_26 : IN std_logic ;
      img_data_23_25 : IN std_logic ;
      img_data_23_24 : IN std_logic ;
      img_data_23_23 : IN std_logic ;
      img_data_23_22 : IN std_logic ;
      img_data_23_21 : IN std_logic ;
      img_data_23_20 : IN std_logic ;
      img_data_23_19 : IN std_logic ;
      img_data_23_18 : IN std_logic ;
      img_data_23_17 : IN std_logic ;
      img_data_23_16 : IN std_logic ;
      img_data_23_15 : IN std_logic ;
      img_data_23_14 : IN std_logic ;
      img_data_23_13 : IN std_logic ;
      img_data_23_12 : IN std_logic ;
      img_data_23_11 : IN std_logic ;
      img_data_23_10 : IN std_logic ;
      img_data_23_9 : IN std_logic ;
      img_data_23_8 : IN std_logic ;
      img_data_23_7 : IN std_logic ;
      img_data_23_6 : IN std_logic ;
      img_data_23_5 : IN std_logic ;
      img_data_23_4 : IN std_logic ;
      img_data_23_3 : IN std_logic ;
      img_data_23_2 : IN std_logic ;
      img_data_23_1 : IN std_logic ;
      img_data_23_0 : IN std_logic ;
      img_data_24_31 : IN std_logic ;
      img_data_24_30 : IN std_logic ;
      img_data_24_29 : IN std_logic ;
      img_data_24_28 : IN std_logic ;
      img_data_24_27 : IN std_logic ;
      img_data_24_26 : IN std_logic ;
      img_data_24_25 : IN std_logic ;
      img_data_24_24 : IN std_logic ;
      img_data_24_23 : IN std_logic ;
      img_data_24_22 : IN std_logic ;
      img_data_24_21 : IN std_logic ;
      img_data_24_20 : IN std_logic ;
      img_data_24_19 : IN std_logic ;
      img_data_24_18 : IN std_logic ;
      img_data_24_17 : IN std_logic ;
      img_data_24_16 : IN std_logic ;
      img_data_24_15 : IN std_logic ;
      img_data_24_14 : IN std_logic ;
      img_data_24_13 : IN std_logic ;
      img_data_24_12 : IN std_logic ;
      img_data_24_11 : IN std_logic ;
      img_data_24_10 : IN std_logic ;
      img_data_24_9 : IN std_logic ;
      img_data_24_8 : IN std_logic ;
      img_data_24_7 : IN std_logic ;
      img_data_24_6 : IN std_logic ;
      img_data_24_5 : IN std_logic ;
      img_data_24_4 : IN std_logic ;
      img_data_24_3 : IN std_logic ;
      img_data_24_2 : IN std_logic ;
      img_data_24_1 : IN std_logic ;
      img_data_24_0 : IN std_logic ;
      filter_data_0_31 : IN std_logic ;
      filter_data_0_30 : IN std_logic ;
      filter_data_0_29 : IN std_logic ;
      filter_data_0_28 : IN std_logic ;
      filter_data_0_27 : IN std_logic ;
      filter_data_0_26 : IN std_logic ;
      filter_data_0_25 : IN std_logic ;
      filter_data_0_24 : IN std_logic ;
      filter_data_0_23 : IN std_logic ;
      filter_data_0_22 : IN std_logic ;
      filter_data_0_21 : IN std_logic ;
      filter_data_0_20 : IN std_logic ;
      filter_data_0_19 : IN std_logic ;
      filter_data_0_18 : IN std_logic ;
      filter_data_0_17 : IN std_logic ;
      filter_data_0_16 : IN std_logic ;
      filter_data_0_15 : IN std_logic ;
      filter_data_0_14 : IN std_logic ;
      filter_data_0_13 : IN std_logic ;
      filter_data_0_12 : IN std_logic ;
      filter_data_0_11 : IN std_logic ;
      filter_data_0_10 : IN std_logic ;
      filter_data_0_9 : IN std_logic ;
      filter_data_0_8 : IN std_logic ;
      filter_data_0_7 : IN std_logic ;
      filter_data_0_6 : IN std_logic ;
      filter_data_0_5 : IN std_logic ;
      filter_data_0_4 : IN std_logic ;
      filter_data_0_3 : IN std_logic ;
      filter_data_0_2 : IN std_logic ;
      filter_data_0_1 : IN std_logic ;
      filter_data_0_0 : IN std_logic ;
      filter_data_1_31 : IN std_logic ;
      filter_data_1_30 : IN std_logic ;
      filter_data_1_29 : IN std_logic ;
      filter_data_1_28 : IN std_logic ;
      filter_data_1_27 : IN std_logic ;
      filter_data_1_26 : IN std_logic ;
      filter_data_1_25 : IN std_logic ;
      filter_data_1_24 : IN std_logic ;
      filter_data_1_23 : IN std_logic ;
      filter_data_1_22 : IN std_logic ;
      filter_data_1_21 : IN std_logic ;
      filter_data_1_20 : IN std_logic ;
      filter_data_1_19 : IN std_logic ;
      filter_data_1_18 : IN std_logic ;
      filter_data_1_17 : IN std_logic ;
      filter_data_1_16 : IN std_logic ;
      filter_data_1_15 : IN std_logic ;
      filter_data_1_14 : IN std_logic ;
      filter_data_1_13 : IN std_logic ;
      filter_data_1_12 : IN std_logic ;
      filter_data_1_11 : IN std_logic ;
      filter_data_1_10 : IN std_logic ;
      filter_data_1_9 : IN std_logic ;
      filter_data_1_8 : IN std_logic ;
      filter_data_1_7 : IN std_logic ;
      filter_data_1_6 : IN std_logic ;
      filter_data_1_5 : IN std_logic ;
      filter_data_1_4 : IN std_logic ;
      filter_data_1_3 : IN std_logic ;
      filter_data_1_2 : IN std_logic ;
      filter_data_1_1 : IN std_logic ;
      filter_data_1_0 : IN std_logic ;
      filter_data_2_31 : IN std_logic ;
      filter_data_2_30 : IN std_logic ;
      filter_data_2_29 : IN std_logic ;
      filter_data_2_28 : IN std_logic ;
      filter_data_2_27 : IN std_logic ;
      filter_data_2_26 : IN std_logic ;
      filter_data_2_25 : IN std_logic ;
      filter_data_2_24 : IN std_logic ;
      filter_data_2_23 : IN std_logic ;
      filter_data_2_22 : IN std_logic ;
      filter_data_2_21 : IN std_logic ;
      filter_data_2_20 : IN std_logic ;
      filter_data_2_19 : IN std_logic ;
      filter_data_2_18 : IN std_logic ;
      filter_data_2_17 : IN std_logic ;
      filter_data_2_16 : IN std_logic ;
      filter_data_2_15 : IN std_logic ;
      filter_data_2_14 : IN std_logic ;
      filter_data_2_13 : IN std_logic ;
      filter_data_2_12 : IN std_logic ;
      filter_data_2_11 : IN std_logic ;
      filter_data_2_10 : IN std_logic ;
      filter_data_2_9 : IN std_logic ;
      filter_data_2_8 : IN std_logic ;
      filter_data_2_7 : IN std_logic ;
      filter_data_2_6 : IN std_logic ;
      filter_data_2_5 : IN std_logic ;
      filter_data_2_4 : IN std_logic ;
      filter_data_2_3 : IN std_logic ;
      filter_data_2_2 : IN std_logic ;
      filter_data_2_1 : IN std_logic ;
      filter_data_2_0 : IN std_logic ;
      filter_data_3_31 : IN std_logic ;
      filter_data_3_30 : IN std_logic ;
      filter_data_3_29 : IN std_logic ;
      filter_data_3_28 : IN std_logic ;
      filter_data_3_27 : IN std_logic ;
      filter_data_3_26 : IN std_logic ;
      filter_data_3_25 : IN std_logic ;
      filter_data_3_24 : IN std_logic ;
      filter_data_3_23 : IN std_logic ;
      filter_data_3_22 : IN std_logic ;
      filter_data_3_21 : IN std_logic ;
      filter_data_3_20 : IN std_logic ;
      filter_data_3_19 : IN std_logic ;
      filter_data_3_18 : IN std_logic ;
      filter_data_3_17 : IN std_logic ;
      filter_data_3_16 : IN std_logic ;
      filter_data_3_15 : IN std_logic ;
      filter_data_3_14 : IN std_logic ;
      filter_data_3_13 : IN std_logic ;
      filter_data_3_12 : IN std_logic ;
      filter_data_3_11 : IN std_logic ;
      filter_data_3_10 : IN std_logic ;
      filter_data_3_9 : IN std_logic ;
      filter_data_3_8 : IN std_logic ;
      filter_data_3_7 : IN std_logic ;
      filter_data_3_6 : IN std_logic ;
      filter_data_3_5 : IN std_logic ;
      filter_data_3_4 : IN std_logic ;
      filter_data_3_3 : IN std_logic ;
      filter_data_3_2 : IN std_logic ;
      filter_data_3_1 : IN std_logic ;
      filter_data_3_0 : IN std_logic ;
      filter_data_4_31 : IN std_logic ;
      filter_data_4_30 : IN std_logic ;
      filter_data_4_29 : IN std_logic ;
      filter_data_4_28 : IN std_logic ;
      filter_data_4_27 : IN std_logic ;
      filter_data_4_26 : IN std_logic ;
      filter_data_4_25 : IN std_logic ;
      filter_data_4_24 : IN std_logic ;
      filter_data_4_23 : IN std_logic ;
      filter_data_4_22 : IN std_logic ;
      filter_data_4_21 : IN std_logic ;
      filter_data_4_20 : IN std_logic ;
      filter_data_4_19 : IN std_logic ;
      filter_data_4_18 : IN std_logic ;
      filter_data_4_17 : IN std_logic ;
      filter_data_4_16 : IN std_logic ;
      filter_data_4_15 : IN std_logic ;
      filter_data_4_14 : IN std_logic ;
      filter_data_4_13 : IN std_logic ;
      filter_data_4_12 : IN std_logic ;
      filter_data_4_11 : IN std_logic ;
      filter_data_4_10 : IN std_logic ;
      filter_data_4_9 : IN std_logic ;
      filter_data_4_8 : IN std_logic ;
      filter_data_4_7 : IN std_logic ;
      filter_data_4_6 : IN std_logic ;
      filter_data_4_5 : IN std_logic ;
      filter_data_4_4 : IN std_logic ;
      filter_data_4_3 : IN std_logic ;
      filter_data_4_2 : IN std_logic ;
      filter_data_4_1 : IN std_logic ;
      filter_data_4_0 : IN std_logic ;
      filter_data_5_31 : IN std_logic ;
      filter_data_5_30 : IN std_logic ;
      filter_data_5_29 : IN std_logic ;
      filter_data_5_28 : IN std_logic ;
      filter_data_5_27 : IN std_logic ;
      filter_data_5_26 : IN std_logic ;
      filter_data_5_25 : IN std_logic ;
      filter_data_5_24 : IN std_logic ;
      filter_data_5_23 : IN std_logic ;
      filter_data_5_22 : IN std_logic ;
      filter_data_5_21 : IN std_logic ;
      filter_data_5_20 : IN std_logic ;
      filter_data_5_19 : IN std_logic ;
      filter_data_5_18 : IN std_logic ;
      filter_data_5_17 : IN std_logic ;
      filter_data_5_16 : IN std_logic ;
      filter_data_5_15 : IN std_logic ;
      filter_data_5_14 : IN std_logic ;
      filter_data_5_13 : IN std_logic ;
      filter_data_5_12 : IN std_logic ;
      filter_data_5_11 : IN std_logic ;
      filter_data_5_10 : IN std_logic ;
      filter_data_5_9 : IN std_logic ;
      filter_data_5_8 : IN std_logic ;
      filter_data_5_7 : IN std_logic ;
      filter_data_5_6 : IN std_logic ;
      filter_data_5_5 : IN std_logic ;
      filter_data_5_4 : IN std_logic ;
      filter_data_5_3 : IN std_logic ;
      filter_data_5_2 : IN std_logic ;
      filter_data_5_1 : IN std_logic ;
      filter_data_5_0 : IN std_logic ;
      filter_data_6_31 : IN std_logic ;
      filter_data_6_30 : IN std_logic ;
      filter_data_6_29 : IN std_logic ;
      filter_data_6_28 : IN std_logic ;
      filter_data_6_27 : IN std_logic ;
      filter_data_6_26 : IN std_logic ;
      filter_data_6_25 : IN std_logic ;
      filter_data_6_24 : IN std_logic ;
      filter_data_6_23 : IN std_logic ;
      filter_data_6_22 : IN std_logic ;
      filter_data_6_21 : IN std_logic ;
      filter_data_6_20 : IN std_logic ;
      filter_data_6_19 : IN std_logic ;
      filter_data_6_18 : IN std_logic ;
      filter_data_6_17 : IN std_logic ;
      filter_data_6_16 : IN std_logic ;
      filter_data_6_15 : IN std_logic ;
      filter_data_6_14 : IN std_logic ;
      filter_data_6_13 : IN std_logic ;
      filter_data_6_12 : IN std_logic ;
      filter_data_6_11 : IN std_logic ;
      filter_data_6_10 : IN std_logic ;
      filter_data_6_9 : IN std_logic ;
      filter_data_6_8 : IN std_logic ;
      filter_data_6_7 : IN std_logic ;
      filter_data_6_6 : IN std_logic ;
      filter_data_6_5 : IN std_logic ;
      filter_data_6_4 : IN std_logic ;
      filter_data_6_3 : IN std_logic ;
      filter_data_6_2 : IN std_logic ;
      filter_data_6_1 : IN std_logic ;
      filter_data_6_0 : IN std_logic ;
      filter_data_7_31 : IN std_logic ;
      filter_data_7_30 : IN std_logic ;
      filter_data_7_29 : IN std_logic ;
      filter_data_7_28 : IN std_logic ;
      filter_data_7_27 : IN std_logic ;
      filter_data_7_26 : IN std_logic ;
      filter_data_7_25 : IN std_logic ;
      filter_data_7_24 : IN std_logic ;
      filter_data_7_23 : IN std_logic ;
      filter_data_7_22 : IN std_logic ;
      filter_data_7_21 : IN std_logic ;
      filter_data_7_20 : IN std_logic ;
      filter_data_7_19 : IN std_logic ;
      filter_data_7_18 : IN std_logic ;
      filter_data_7_17 : IN std_logic ;
      filter_data_7_16 : IN std_logic ;
      filter_data_7_15 : IN std_logic ;
      filter_data_7_14 : IN std_logic ;
      filter_data_7_13 : IN std_logic ;
      filter_data_7_12 : IN std_logic ;
      filter_data_7_11 : IN std_logic ;
      filter_data_7_10 : IN std_logic ;
      filter_data_7_9 : IN std_logic ;
      filter_data_7_8 : IN std_logic ;
      filter_data_7_7 : IN std_logic ;
      filter_data_7_6 : IN std_logic ;
      filter_data_7_5 : IN std_logic ;
      filter_data_7_4 : IN std_logic ;
      filter_data_7_3 : IN std_logic ;
      filter_data_7_2 : IN std_logic ;
      filter_data_7_1 : IN std_logic ;
      filter_data_7_0 : IN std_logic ;
      filter_data_8_31 : IN std_logic ;
      filter_data_8_30 : IN std_logic ;
      filter_data_8_29 : IN std_logic ;
      filter_data_8_28 : IN std_logic ;
      filter_data_8_27 : IN std_logic ;
      filter_data_8_26 : IN std_logic ;
      filter_data_8_25 : IN std_logic ;
      filter_data_8_24 : IN std_logic ;
      filter_data_8_23 : IN std_logic ;
      filter_data_8_22 : IN std_logic ;
      filter_data_8_21 : IN std_logic ;
      filter_data_8_20 : IN std_logic ;
      filter_data_8_19 : IN std_logic ;
      filter_data_8_18 : IN std_logic ;
      filter_data_8_17 : IN std_logic ;
      filter_data_8_16 : IN std_logic ;
      filter_data_8_15 : IN std_logic ;
      filter_data_8_14 : IN std_logic ;
      filter_data_8_13 : IN std_logic ;
      filter_data_8_12 : IN std_logic ;
      filter_data_8_11 : IN std_logic ;
      filter_data_8_10 : IN std_logic ;
      filter_data_8_9 : IN std_logic ;
      filter_data_8_8 : IN std_logic ;
      filter_data_8_7 : IN std_logic ;
      filter_data_8_6 : IN std_logic ;
      filter_data_8_5 : IN std_logic ;
      filter_data_8_4 : IN std_logic ;
      filter_data_8_3 : IN std_logic ;
      filter_data_8_2 : IN std_logic ;
      filter_data_8_1 : IN std_logic ;
      filter_data_8_0 : IN std_logic ;
      filter_data_9_31 : IN std_logic ;
      filter_data_9_30 : IN std_logic ;
      filter_data_9_29 : IN std_logic ;
      filter_data_9_28 : IN std_logic ;
      filter_data_9_27 : IN std_logic ;
      filter_data_9_26 : IN std_logic ;
      filter_data_9_25 : IN std_logic ;
      filter_data_9_24 : IN std_logic ;
      filter_data_9_23 : IN std_logic ;
      filter_data_9_22 : IN std_logic ;
      filter_data_9_21 : IN std_logic ;
      filter_data_9_20 : IN std_logic ;
      filter_data_9_19 : IN std_logic ;
      filter_data_9_18 : IN std_logic ;
      filter_data_9_17 : IN std_logic ;
      filter_data_9_16 : IN std_logic ;
      filter_data_9_15 : IN std_logic ;
      filter_data_9_14 : IN std_logic ;
      filter_data_9_13 : IN std_logic ;
      filter_data_9_12 : IN std_logic ;
      filter_data_9_11 : IN std_logic ;
      filter_data_9_10 : IN std_logic ;
      filter_data_9_9 : IN std_logic ;
      filter_data_9_8 : IN std_logic ;
      filter_data_9_7 : IN std_logic ;
      filter_data_9_6 : IN std_logic ;
      filter_data_9_5 : IN std_logic ;
      filter_data_9_4 : IN std_logic ;
      filter_data_9_3 : IN std_logic ;
      filter_data_9_2 : IN std_logic ;
      filter_data_9_1 : IN std_logic ;
      filter_data_9_0 : IN std_logic ;
      filter_data_10_31 : IN std_logic ;
      filter_data_10_30 : IN std_logic ;
      filter_data_10_29 : IN std_logic ;
      filter_data_10_28 : IN std_logic ;
      filter_data_10_27 : IN std_logic ;
      filter_data_10_26 : IN std_logic ;
      filter_data_10_25 : IN std_logic ;
      filter_data_10_24 : IN std_logic ;
      filter_data_10_23 : IN std_logic ;
      filter_data_10_22 : IN std_logic ;
      filter_data_10_21 : IN std_logic ;
      filter_data_10_20 : IN std_logic ;
      filter_data_10_19 : IN std_logic ;
      filter_data_10_18 : IN std_logic ;
      filter_data_10_17 : IN std_logic ;
      filter_data_10_16 : IN std_logic ;
      filter_data_10_15 : IN std_logic ;
      filter_data_10_14 : IN std_logic ;
      filter_data_10_13 : IN std_logic ;
      filter_data_10_12 : IN std_logic ;
      filter_data_10_11 : IN std_logic ;
      filter_data_10_10 : IN std_logic ;
      filter_data_10_9 : IN std_logic ;
      filter_data_10_8 : IN std_logic ;
      filter_data_10_7 : IN std_logic ;
      filter_data_10_6 : IN std_logic ;
      filter_data_10_5 : IN std_logic ;
      filter_data_10_4 : IN std_logic ;
      filter_data_10_3 : IN std_logic ;
      filter_data_10_2 : IN std_logic ;
      filter_data_10_1 : IN std_logic ;
      filter_data_10_0 : IN std_logic ;
      filter_data_11_31 : IN std_logic ;
      filter_data_11_30 : IN std_logic ;
      filter_data_11_29 : IN std_logic ;
      filter_data_11_28 : IN std_logic ;
      filter_data_11_27 : IN std_logic ;
      filter_data_11_26 : IN std_logic ;
      filter_data_11_25 : IN std_logic ;
      filter_data_11_24 : IN std_logic ;
      filter_data_11_23 : IN std_logic ;
      filter_data_11_22 : IN std_logic ;
      filter_data_11_21 : IN std_logic ;
      filter_data_11_20 : IN std_logic ;
      filter_data_11_19 : IN std_logic ;
      filter_data_11_18 : IN std_logic ;
      filter_data_11_17 : IN std_logic ;
      filter_data_11_16 : IN std_logic ;
      filter_data_11_15 : IN std_logic ;
      filter_data_11_14 : IN std_logic ;
      filter_data_11_13 : IN std_logic ;
      filter_data_11_12 : IN std_logic ;
      filter_data_11_11 : IN std_logic ;
      filter_data_11_10 : IN std_logic ;
      filter_data_11_9 : IN std_logic ;
      filter_data_11_8 : IN std_logic ;
      filter_data_11_7 : IN std_logic ;
      filter_data_11_6 : IN std_logic ;
      filter_data_11_5 : IN std_logic ;
      filter_data_11_4 : IN std_logic ;
      filter_data_11_3 : IN std_logic ;
      filter_data_11_2 : IN std_logic ;
      filter_data_11_1 : IN std_logic ;
      filter_data_11_0 : IN std_logic ;
      filter_data_12_31 : IN std_logic ;
      filter_data_12_30 : IN std_logic ;
      filter_data_12_29 : IN std_logic ;
      filter_data_12_28 : IN std_logic ;
      filter_data_12_27 : IN std_logic ;
      filter_data_12_26 : IN std_logic ;
      filter_data_12_25 : IN std_logic ;
      filter_data_12_24 : IN std_logic ;
      filter_data_12_23 : IN std_logic ;
      filter_data_12_22 : IN std_logic ;
      filter_data_12_21 : IN std_logic ;
      filter_data_12_20 : IN std_logic ;
      filter_data_12_19 : IN std_logic ;
      filter_data_12_18 : IN std_logic ;
      filter_data_12_17 : IN std_logic ;
      filter_data_12_16 : IN std_logic ;
      filter_data_12_15 : IN std_logic ;
      filter_data_12_14 : IN std_logic ;
      filter_data_12_13 : IN std_logic ;
      filter_data_12_12 : IN std_logic ;
      filter_data_12_11 : IN std_logic ;
      filter_data_12_10 : IN std_logic ;
      filter_data_12_9 : IN std_logic ;
      filter_data_12_8 : IN std_logic ;
      filter_data_12_7 : IN std_logic ;
      filter_data_12_6 : IN std_logic ;
      filter_data_12_5 : IN std_logic ;
      filter_data_12_4 : IN std_logic ;
      filter_data_12_3 : IN std_logic ;
      filter_data_12_2 : IN std_logic ;
      filter_data_12_1 : IN std_logic ;
      filter_data_12_0 : IN std_logic ;
      filter_data_13_31 : IN std_logic ;
      filter_data_13_30 : IN std_logic ;
      filter_data_13_29 : IN std_logic ;
      filter_data_13_28 : IN std_logic ;
      filter_data_13_27 : IN std_logic ;
      filter_data_13_26 : IN std_logic ;
      filter_data_13_25 : IN std_logic ;
      filter_data_13_24 : IN std_logic ;
      filter_data_13_23 : IN std_logic ;
      filter_data_13_22 : IN std_logic ;
      filter_data_13_21 : IN std_logic ;
      filter_data_13_20 : IN std_logic ;
      filter_data_13_19 : IN std_logic ;
      filter_data_13_18 : IN std_logic ;
      filter_data_13_17 : IN std_logic ;
      filter_data_13_16 : IN std_logic ;
      filter_data_13_15 : IN std_logic ;
      filter_data_13_14 : IN std_logic ;
      filter_data_13_13 : IN std_logic ;
      filter_data_13_12 : IN std_logic ;
      filter_data_13_11 : IN std_logic ;
      filter_data_13_10 : IN std_logic ;
      filter_data_13_9 : IN std_logic ;
      filter_data_13_8 : IN std_logic ;
      filter_data_13_7 : IN std_logic ;
      filter_data_13_6 : IN std_logic ;
      filter_data_13_5 : IN std_logic ;
      filter_data_13_4 : IN std_logic ;
      filter_data_13_3 : IN std_logic ;
      filter_data_13_2 : IN std_logic ;
      filter_data_13_1 : IN std_logic ;
      filter_data_13_0 : IN std_logic ;
      filter_data_14_31 : IN std_logic ;
      filter_data_14_30 : IN std_logic ;
      filter_data_14_29 : IN std_logic ;
      filter_data_14_28 : IN std_logic ;
      filter_data_14_27 : IN std_logic ;
      filter_data_14_26 : IN std_logic ;
      filter_data_14_25 : IN std_logic ;
      filter_data_14_24 : IN std_logic ;
      filter_data_14_23 : IN std_logic ;
      filter_data_14_22 : IN std_logic ;
      filter_data_14_21 : IN std_logic ;
      filter_data_14_20 : IN std_logic ;
      filter_data_14_19 : IN std_logic ;
      filter_data_14_18 : IN std_logic ;
      filter_data_14_17 : IN std_logic ;
      filter_data_14_16 : IN std_logic ;
      filter_data_14_15 : IN std_logic ;
      filter_data_14_14 : IN std_logic ;
      filter_data_14_13 : IN std_logic ;
      filter_data_14_12 : IN std_logic ;
      filter_data_14_11 : IN std_logic ;
      filter_data_14_10 : IN std_logic ;
      filter_data_14_9 : IN std_logic ;
      filter_data_14_8 : IN std_logic ;
      filter_data_14_7 : IN std_logic ;
      filter_data_14_6 : IN std_logic ;
      filter_data_14_5 : IN std_logic ;
      filter_data_14_4 : IN std_logic ;
      filter_data_14_3 : IN std_logic ;
      filter_data_14_2 : IN std_logic ;
      filter_data_14_1 : IN std_logic ;
      filter_data_14_0 : IN std_logic ;
      filter_data_15_31 : IN std_logic ;
      filter_data_15_30 : IN std_logic ;
      filter_data_15_29 : IN std_logic ;
      filter_data_15_28 : IN std_logic ;
      filter_data_15_27 : IN std_logic ;
      filter_data_15_26 : IN std_logic ;
      filter_data_15_25 : IN std_logic ;
      filter_data_15_24 : IN std_logic ;
      filter_data_15_23 : IN std_logic ;
      filter_data_15_22 : IN std_logic ;
      filter_data_15_21 : IN std_logic ;
      filter_data_15_20 : IN std_logic ;
      filter_data_15_19 : IN std_logic ;
      filter_data_15_18 : IN std_logic ;
      filter_data_15_17 : IN std_logic ;
      filter_data_15_16 : IN std_logic ;
      filter_data_15_15 : IN std_logic ;
      filter_data_15_14 : IN std_logic ;
      filter_data_15_13 : IN std_logic ;
      filter_data_15_12 : IN std_logic ;
      filter_data_15_11 : IN std_logic ;
      filter_data_15_10 : IN std_logic ;
      filter_data_15_9 : IN std_logic ;
      filter_data_15_8 : IN std_logic ;
      filter_data_15_7 : IN std_logic ;
      filter_data_15_6 : IN std_logic ;
      filter_data_15_5 : IN std_logic ;
      filter_data_15_4 : IN std_logic ;
      filter_data_15_3 : IN std_logic ;
      filter_data_15_2 : IN std_logic ;
      filter_data_15_1 : IN std_logic ;
      filter_data_15_0 : IN std_logic ;
      filter_data_16_31 : IN std_logic ;
      filter_data_16_30 : IN std_logic ;
      filter_data_16_29 : IN std_logic ;
      filter_data_16_28 : IN std_logic ;
      filter_data_16_27 : IN std_logic ;
      filter_data_16_26 : IN std_logic ;
      filter_data_16_25 : IN std_logic ;
      filter_data_16_24 : IN std_logic ;
      filter_data_16_23 : IN std_logic ;
      filter_data_16_22 : IN std_logic ;
      filter_data_16_21 : IN std_logic ;
      filter_data_16_20 : IN std_logic ;
      filter_data_16_19 : IN std_logic ;
      filter_data_16_18 : IN std_logic ;
      filter_data_16_17 : IN std_logic ;
      filter_data_16_16 : IN std_logic ;
      filter_data_16_15 : IN std_logic ;
      filter_data_16_14 : IN std_logic ;
      filter_data_16_13 : IN std_logic ;
      filter_data_16_12 : IN std_logic ;
      filter_data_16_11 : IN std_logic ;
      filter_data_16_10 : IN std_logic ;
      filter_data_16_9 : IN std_logic ;
      filter_data_16_8 : IN std_logic ;
      filter_data_16_7 : IN std_logic ;
      filter_data_16_6 : IN std_logic ;
      filter_data_16_5 : IN std_logic ;
      filter_data_16_4 : IN std_logic ;
      filter_data_16_3 : IN std_logic ;
      filter_data_16_2 : IN std_logic ;
      filter_data_16_1 : IN std_logic ;
      filter_data_16_0 : IN std_logic ;
      filter_data_17_31 : IN std_logic ;
      filter_data_17_30 : IN std_logic ;
      filter_data_17_29 : IN std_logic ;
      filter_data_17_28 : IN std_logic ;
      filter_data_17_27 : IN std_logic ;
      filter_data_17_26 : IN std_logic ;
      filter_data_17_25 : IN std_logic ;
      filter_data_17_24 : IN std_logic ;
      filter_data_17_23 : IN std_logic ;
      filter_data_17_22 : IN std_logic ;
      filter_data_17_21 : IN std_logic ;
      filter_data_17_20 : IN std_logic ;
      filter_data_17_19 : IN std_logic ;
      filter_data_17_18 : IN std_logic ;
      filter_data_17_17 : IN std_logic ;
      filter_data_17_16 : IN std_logic ;
      filter_data_17_15 : IN std_logic ;
      filter_data_17_14 : IN std_logic ;
      filter_data_17_13 : IN std_logic ;
      filter_data_17_12 : IN std_logic ;
      filter_data_17_11 : IN std_logic ;
      filter_data_17_10 : IN std_logic ;
      filter_data_17_9 : IN std_logic ;
      filter_data_17_8 : IN std_logic ;
      filter_data_17_7 : IN std_logic ;
      filter_data_17_6 : IN std_logic ;
      filter_data_17_5 : IN std_logic ;
      filter_data_17_4 : IN std_logic ;
      filter_data_17_3 : IN std_logic ;
      filter_data_17_2 : IN std_logic ;
      filter_data_17_1 : IN std_logic ;
      filter_data_17_0 : IN std_logic ;
      filter_data_18_31 : IN std_logic ;
      filter_data_18_30 : IN std_logic ;
      filter_data_18_29 : IN std_logic ;
      filter_data_18_28 : IN std_logic ;
      filter_data_18_27 : IN std_logic ;
      filter_data_18_26 : IN std_logic ;
      filter_data_18_25 : IN std_logic ;
      filter_data_18_24 : IN std_logic ;
      filter_data_18_23 : IN std_logic ;
      filter_data_18_22 : IN std_logic ;
      filter_data_18_21 : IN std_logic ;
      filter_data_18_20 : IN std_logic ;
      filter_data_18_19 : IN std_logic ;
      filter_data_18_18 : IN std_logic ;
      filter_data_18_17 : IN std_logic ;
      filter_data_18_16 : IN std_logic ;
      filter_data_18_15 : IN std_logic ;
      filter_data_18_14 : IN std_logic ;
      filter_data_18_13 : IN std_logic ;
      filter_data_18_12 : IN std_logic ;
      filter_data_18_11 : IN std_logic ;
      filter_data_18_10 : IN std_logic ;
      filter_data_18_9 : IN std_logic ;
      filter_data_18_8 : IN std_logic ;
      filter_data_18_7 : IN std_logic ;
      filter_data_18_6 : IN std_logic ;
      filter_data_18_5 : IN std_logic ;
      filter_data_18_4 : IN std_logic ;
      filter_data_18_3 : IN std_logic ;
      filter_data_18_2 : IN std_logic ;
      filter_data_18_1 : IN std_logic ;
      filter_data_18_0 : IN std_logic ;
      filter_data_19_31 : IN std_logic ;
      filter_data_19_30 : IN std_logic ;
      filter_data_19_29 : IN std_logic ;
      filter_data_19_28 : IN std_logic ;
      filter_data_19_27 : IN std_logic ;
      filter_data_19_26 : IN std_logic ;
      filter_data_19_25 : IN std_logic ;
      filter_data_19_24 : IN std_logic ;
      filter_data_19_23 : IN std_logic ;
      filter_data_19_22 : IN std_logic ;
      filter_data_19_21 : IN std_logic ;
      filter_data_19_20 : IN std_logic ;
      filter_data_19_19 : IN std_logic ;
      filter_data_19_18 : IN std_logic ;
      filter_data_19_17 : IN std_logic ;
      filter_data_19_16 : IN std_logic ;
      filter_data_19_15 : IN std_logic ;
      filter_data_19_14 : IN std_logic ;
      filter_data_19_13 : IN std_logic ;
      filter_data_19_12 : IN std_logic ;
      filter_data_19_11 : IN std_logic ;
      filter_data_19_10 : IN std_logic ;
      filter_data_19_9 : IN std_logic ;
      filter_data_19_8 : IN std_logic ;
      filter_data_19_7 : IN std_logic ;
      filter_data_19_6 : IN std_logic ;
      filter_data_19_5 : IN std_logic ;
      filter_data_19_4 : IN std_logic ;
      filter_data_19_3 : IN std_logic ;
      filter_data_19_2 : IN std_logic ;
      filter_data_19_1 : IN std_logic ;
      filter_data_19_0 : IN std_logic ;
      filter_data_20_31 : IN std_logic ;
      filter_data_20_30 : IN std_logic ;
      filter_data_20_29 : IN std_logic ;
      filter_data_20_28 : IN std_logic ;
      filter_data_20_27 : IN std_logic ;
      filter_data_20_26 : IN std_logic ;
      filter_data_20_25 : IN std_logic ;
      filter_data_20_24 : IN std_logic ;
      filter_data_20_23 : IN std_logic ;
      filter_data_20_22 : IN std_logic ;
      filter_data_20_21 : IN std_logic ;
      filter_data_20_20 : IN std_logic ;
      filter_data_20_19 : IN std_logic ;
      filter_data_20_18 : IN std_logic ;
      filter_data_20_17 : IN std_logic ;
      filter_data_20_16 : IN std_logic ;
      filter_data_20_15 : IN std_logic ;
      filter_data_20_14 : IN std_logic ;
      filter_data_20_13 : IN std_logic ;
      filter_data_20_12 : IN std_logic ;
      filter_data_20_11 : IN std_logic ;
      filter_data_20_10 : IN std_logic ;
      filter_data_20_9 : IN std_logic ;
      filter_data_20_8 : IN std_logic ;
      filter_data_20_7 : IN std_logic ;
      filter_data_20_6 : IN std_logic ;
      filter_data_20_5 : IN std_logic ;
      filter_data_20_4 : IN std_logic ;
      filter_data_20_3 : IN std_logic ;
      filter_data_20_2 : IN std_logic ;
      filter_data_20_1 : IN std_logic ;
      filter_data_20_0 : IN std_logic ;
      filter_data_21_31 : IN std_logic ;
      filter_data_21_30 : IN std_logic ;
      filter_data_21_29 : IN std_logic ;
      filter_data_21_28 : IN std_logic ;
      filter_data_21_27 : IN std_logic ;
      filter_data_21_26 : IN std_logic ;
      filter_data_21_25 : IN std_logic ;
      filter_data_21_24 : IN std_logic ;
      filter_data_21_23 : IN std_logic ;
      filter_data_21_22 : IN std_logic ;
      filter_data_21_21 : IN std_logic ;
      filter_data_21_20 : IN std_logic ;
      filter_data_21_19 : IN std_logic ;
      filter_data_21_18 : IN std_logic ;
      filter_data_21_17 : IN std_logic ;
      filter_data_21_16 : IN std_logic ;
      filter_data_21_15 : IN std_logic ;
      filter_data_21_14 : IN std_logic ;
      filter_data_21_13 : IN std_logic ;
      filter_data_21_12 : IN std_logic ;
      filter_data_21_11 : IN std_logic ;
      filter_data_21_10 : IN std_logic ;
      filter_data_21_9 : IN std_logic ;
      filter_data_21_8 : IN std_logic ;
      filter_data_21_7 : IN std_logic ;
      filter_data_21_6 : IN std_logic ;
      filter_data_21_5 : IN std_logic ;
      filter_data_21_4 : IN std_logic ;
      filter_data_21_3 : IN std_logic ;
      filter_data_21_2 : IN std_logic ;
      filter_data_21_1 : IN std_logic ;
      filter_data_21_0 : IN std_logic ;
      filter_data_22_31 : IN std_logic ;
      filter_data_22_30 : IN std_logic ;
      filter_data_22_29 : IN std_logic ;
      filter_data_22_28 : IN std_logic ;
      filter_data_22_27 : IN std_logic ;
      filter_data_22_26 : IN std_logic ;
      filter_data_22_25 : IN std_logic ;
      filter_data_22_24 : IN std_logic ;
      filter_data_22_23 : IN std_logic ;
      filter_data_22_22 : IN std_logic ;
      filter_data_22_21 : IN std_logic ;
      filter_data_22_20 : IN std_logic ;
      filter_data_22_19 : IN std_logic ;
      filter_data_22_18 : IN std_logic ;
      filter_data_22_17 : IN std_logic ;
      filter_data_22_16 : IN std_logic ;
      filter_data_22_15 : IN std_logic ;
      filter_data_22_14 : IN std_logic ;
      filter_data_22_13 : IN std_logic ;
      filter_data_22_12 : IN std_logic ;
      filter_data_22_11 : IN std_logic ;
      filter_data_22_10 : IN std_logic ;
      filter_data_22_9 : IN std_logic ;
      filter_data_22_8 : IN std_logic ;
      filter_data_22_7 : IN std_logic ;
      filter_data_22_6 : IN std_logic ;
      filter_data_22_5 : IN std_logic ;
      filter_data_22_4 : IN std_logic ;
      filter_data_22_3 : IN std_logic ;
      filter_data_22_2 : IN std_logic ;
      filter_data_22_1 : IN std_logic ;
      filter_data_22_0 : IN std_logic ;
      filter_data_23_31 : IN std_logic ;
      filter_data_23_30 : IN std_logic ;
      filter_data_23_29 : IN std_logic ;
      filter_data_23_28 : IN std_logic ;
      filter_data_23_27 : IN std_logic ;
      filter_data_23_26 : IN std_logic ;
      filter_data_23_25 : IN std_logic ;
      filter_data_23_24 : IN std_logic ;
      filter_data_23_23 : IN std_logic ;
      filter_data_23_22 : IN std_logic ;
      filter_data_23_21 : IN std_logic ;
      filter_data_23_20 : IN std_logic ;
      filter_data_23_19 : IN std_logic ;
      filter_data_23_18 : IN std_logic ;
      filter_data_23_17 : IN std_logic ;
      filter_data_23_16 : IN std_logic ;
      filter_data_23_15 : IN std_logic ;
      filter_data_23_14 : IN std_logic ;
      filter_data_23_13 : IN std_logic ;
      filter_data_23_12 : IN std_logic ;
      filter_data_23_11 : IN std_logic ;
      filter_data_23_10 : IN std_logic ;
      filter_data_23_9 : IN std_logic ;
      filter_data_23_8 : IN std_logic ;
      filter_data_23_7 : IN std_logic ;
      filter_data_23_6 : IN std_logic ;
      filter_data_23_5 : IN std_logic ;
      filter_data_23_4 : IN std_logic ;
      filter_data_23_3 : IN std_logic ;
      filter_data_23_2 : IN std_logic ;
      filter_data_23_1 : IN std_logic ;
      filter_data_23_0 : IN std_logic ;
      filter_data_24_31 : IN std_logic ;
      filter_data_24_30 : IN std_logic ;
      filter_data_24_29 : IN std_logic ;
      filter_data_24_28 : IN std_logic ;
      filter_data_24_27 : IN std_logic ;
      filter_data_24_26 : IN std_logic ;
      filter_data_24_25 : IN std_logic ;
      filter_data_24_24 : IN std_logic ;
      filter_data_24_23 : IN std_logic ;
      filter_data_24_22 : IN std_logic ;
      filter_data_24_21 : IN std_logic ;
      filter_data_24_20 : IN std_logic ;
      filter_data_24_19 : IN std_logic ;
      filter_data_24_18 : IN std_logic ;
      filter_data_24_17 : IN std_logic ;
      filter_data_24_16 : IN std_logic ;
      filter_data_24_15 : IN std_logic ;
      filter_data_24_14 : IN std_logic ;
      filter_data_24_13 : IN std_logic ;
      filter_data_24_12 : IN std_logic ;
      filter_data_24_11 : IN std_logic ;
      filter_data_24_10 : IN std_logic ;
      filter_data_24_9 : IN std_logic ;
      filter_data_24_8 : IN std_logic ;
      filter_data_24_7 : IN std_logic ;
      filter_data_24_6 : IN std_logic ;
      filter_data_24_5 : IN std_logic ;
      filter_data_24_4 : IN std_logic ;
      filter_data_24_3 : IN std_logic ;
      filter_data_24_2 : IN std_logic ;
      filter_data_24_1 : IN std_logic ;
      filter_data_24_0 : IN std_logic ;
      filter_size : IN std_logic ;
      ordered_img_data_0_31 : OUT std_logic ;
      ordered_img_data_0_30 : OUT std_logic ;
      ordered_img_data_0_29 : OUT std_logic ;
      ordered_img_data_0_28 : OUT std_logic ;
      ordered_img_data_0_27 : OUT std_logic ;
      ordered_img_data_0_26 : OUT std_logic ;
      ordered_img_data_0_25 : OUT std_logic ;
      ordered_img_data_0_24 : OUT std_logic ;
      ordered_img_data_0_23 : OUT std_logic ;
      ordered_img_data_0_22 : OUT std_logic ;
      ordered_img_data_0_21 : OUT std_logic ;
      ordered_img_data_0_20 : OUT std_logic ;
      ordered_img_data_0_19 : OUT std_logic ;
      ordered_img_data_0_18 : OUT std_logic ;
      ordered_img_data_0_17 : OUT std_logic ;
      ordered_img_data_0_16 : OUT std_logic ;
      ordered_img_data_0_15 : OUT std_logic ;
      ordered_img_data_0_14 : OUT std_logic ;
      ordered_img_data_0_13 : OUT std_logic ;
      ordered_img_data_0_12 : OUT std_logic ;
      ordered_img_data_0_11 : OUT std_logic ;
      ordered_img_data_0_10 : OUT std_logic ;
      ordered_img_data_0_9 : OUT std_logic ;
      ordered_img_data_0_8 : OUT std_logic ;
      ordered_img_data_0_7 : OUT std_logic ;
      ordered_img_data_0_6 : OUT std_logic ;
      ordered_img_data_0_5 : OUT std_logic ;
      ordered_img_data_0_4 : OUT std_logic ;
      ordered_img_data_0_3 : OUT std_logic ;
      ordered_img_data_0_2 : OUT std_logic ;
      ordered_img_data_0_1 : OUT std_logic ;
      ordered_img_data_0_0 : OUT std_logic ;
      ordered_img_data_1_31 : OUT std_logic ;
      ordered_img_data_1_30 : OUT std_logic ;
      ordered_img_data_1_29 : OUT std_logic ;
      ordered_img_data_1_28 : OUT std_logic ;
      ordered_img_data_1_27 : OUT std_logic ;
      ordered_img_data_1_26 : OUT std_logic ;
      ordered_img_data_1_25 : OUT std_logic ;
      ordered_img_data_1_24 : OUT std_logic ;
      ordered_img_data_1_23 : OUT std_logic ;
      ordered_img_data_1_22 : OUT std_logic ;
      ordered_img_data_1_21 : OUT std_logic ;
      ordered_img_data_1_20 : OUT std_logic ;
      ordered_img_data_1_19 : OUT std_logic ;
      ordered_img_data_1_18 : OUT std_logic ;
      ordered_img_data_1_17 : OUT std_logic ;
      ordered_img_data_1_16 : OUT std_logic ;
      ordered_img_data_1_15 : OUT std_logic ;
      ordered_img_data_1_14 : OUT std_logic ;
      ordered_img_data_1_13 : OUT std_logic ;
      ordered_img_data_1_12 : OUT std_logic ;
      ordered_img_data_1_11 : OUT std_logic ;
      ordered_img_data_1_10 : OUT std_logic ;
      ordered_img_data_1_9 : OUT std_logic ;
      ordered_img_data_1_8 : OUT std_logic ;
      ordered_img_data_1_7 : OUT std_logic ;
      ordered_img_data_1_6 : OUT std_logic ;
      ordered_img_data_1_5 : OUT std_logic ;
      ordered_img_data_1_4 : OUT std_logic ;
      ordered_img_data_1_3 : OUT std_logic ;
      ordered_img_data_1_2 : OUT std_logic ;
      ordered_img_data_1_1 : OUT std_logic ;
      ordered_img_data_1_0 : OUT std_logic ;
      ordered_img_data_2_31 : OUT std_logic ;
      ordered_img_data_2_30 : OUT std_logic ;
      ordered_img_data_2_29 : OUT std_logic ;
      ordered_img_data_2_28 : OUT std_logic ;
      ordered_img_data_2_27 : OUT std_logic ;
      ordered_img_data_2_26 : OUT std_logic ;
      ordered_img_data_2_25 : OUT std_logic ;
      ordered_img_data_2_24 : OUT std_logic ;
      ordered_img_data_2_23 : OUT std_logic ;
      ordered_img_data_2_22 : OUT std_logic ;
      ordered_img_data_2_21 : OUT std_logic ;
      ordered_img_data_2_20 : OUT std_logic ;
      ordered_img_data_2_19 : OUT std_logic ;
      ordered_img_data_2_18 : OUT std_logic ;
      ordered_img_data_2_17 : OUT std_logic ;
      ordered_img_data_2_16 : OUT std_logic ;
      ordered_img_data_2_15 : OUT std_logic ;
      ordered_img_data_2_14 : OUT std_logic ;
      ordered_img_data_2_13 : OUT std_logic ;
      ordered_img_data_2_12 : OUT std_logic ;
      ordered_img_data_2_11 : OUT std_logic ;
      ordered_img_data_2_10 : OUT std_logic ;
      ordered_img_data_2_9 : OUT std_logic ;
      ordered_img_data_2_8 : OUT std_logic ;
      ordered_img_data_2_7 : OUT std_logic ;
      ordered_img_data_2_6 : OUT std_logic ;
      ordered_img_data_2_5 : OUT std_logic ;
      ordered_img_data_2_4 : OUT std_logic ;
      ordered_img_data_2_3 : OUT std_logic ;
      ordered_img_data_2_2 : OUT std_logic ;
      ordered_img_data_2_1 : OUT std_logic ;
      ordered_img_data_2_0 : OUT std_logic ;
      ordered_img_data_3_31 : OUT std_logic ;
      ordered_img_data_3_30 : OUT std_logic ;
      ordered_img_data_3_29 : OUT std_logic ;
      ordered_img_data_3_28 : OUT std_logic ;
      ordered_img_data_3_27 : OUT std_logic ;
      ordered_img_data_3_26 : OUT std_logic ;
      ordered_img_data_3_25 : OUT std_logic ;
      ordered_img_data_3_24 : OUT std_logic ;
      ordered_img_data_3_23 : OUT std_logic ;
      ordered_img_data_3_22 : OUT std_logic ;
      ordered_img_data_3_21 : OUT std_logic ;
      ordered_img_data_3_20 : OUT std_logic ;
      ordered_img_data_3_19 : OUT std_logic ;
      ordered_img_data_3_18 : OUT std_logic ;
      ordered_img_data_3_17 : OUT std_logic ;
      ordered_img_data_3_16 : OUT std_logic ;
      ordered_img_data_3_15 : OUT std_logic ;
      ordered_img_data_3_14 : OUT std_logic ;
      ordered_img_data_3_13 : OUT std_logic ;
      ordered_img_data_3_12 : OUT std_logic ;
      ordered_img_data_3_11 : OUT std_logic ;
      ordered_img_data_3_10 : OUT std_logic ;
      ordered_img_data_3_9 : OUT std_logic ;
      ordered_img_data_3_8 : OUT std_logic ;
      ordered_img_data_3_7 : OUT std_logic ;
      ordered_img_data_3_6 : OUT std_logic ;
      ordered_img_data_3_5 : OUT std_logic ;
      ordered_img_data_3_4 : OUT std_logic ;
      ordered_img_data_3_3 : OUT std_logic ;
      ordered_img_data_3_2 : OUT std_logic ;
      ordered_img_data_3_1 : OUT std_logic ;
      ordered_img_data_3_0 : OUT std_logic ;
      ordered_img_data_4_31 : OUT std_logic ;
      ordered_img_data_4_30 : OUT std_logic ;
      ordered_img_data_4_29 : OUT std_logic ;
      ordered_img_data_4_28 : OUT std_logic ;
      ordered_img_data_4_27 : OUT std_logic ;
      ordered_img_data_4_26 : OUT std_logic ;
      ordered_img_data_4_25 : OUT std_logic ;
      ordered_img_data_4_24 : OUT std_logic ;
      ordered_img_data_4_23 : OUT std_logic ;
      ordered_img_data_4_22 : OUT std_logic ;
      ordered_img_data_4_21 : OUT std_logic ;
      ordered_img_data_4_20 : OUT std_logic ;
      ordered_img_data_4_19 : OUT std_logic ;
      ordered_img_data_4_18 : OUT std_logic ;
      ordered_img_data_4_17 : OUT std_logic ;
      ordered_img_data_4_16 : OUT std_logic ;
      ordered_img_data_4_15 : OUT std_logic ;
      ordered_img_data_4_14 : OUT std_logic ;
      ordered_img_data_4_13 : OUT std_logic ;
      ordered_img_data_4_12 : OUT std_logic ;
      ordered_img_data_4_11 : OUT std_logic ;
      ordered_img_data_4_10 : OUT std_logic ;
      ordered_img_data_4_9 : OUT std_logic ;
      ordered_img_data_4_8 : OUT std_logic ;
      ordered_img_data_4_7 : OUT std_logic ;
      ordered_img_data_4_6 : OUT std_logic ;
      ordered_img_data_4_5 : OUT std_logic ;
      ordered_img_data_4_4 : OUT std_logic ;
      ordered_img_data_4_3 : OUT std_logic ;
      ordered_img_data_4_2 : OUT std_logic ;
      ordered_img_data_4_1 : OUT std_logic ;
      ordered_img_data_4_0 : OUT std_logic ;
      ordered_img_data_5_31 : OUT std_logic ;
      ordered_img_data_5_30 : OUT std_logic ;
      ordered_img_data_5_29 : OUT std_logic ;
      ordered_img_data_5_28 : OUT std_logic ;
      ordered_img_data_5_27 : OUT std_logic ;
      ordered_img_data_5_26 : OUT std_logic ;
      ordered_img_data_5_25 : OUT std_logic ;
      ordered_img_data_5_24 : OUT std_logic ;
      ordered_img_data_5_23 : OUT std_logic ;
      ordered_img_data_5_22 : OUT std_logic ;
      ordered_img_data_5_21 : OUT std_logic ;
      ordered_img_data_5_20 : OUT std_logic ;
      ordered_img_data_5_19 : OUT std_logic ;
      ordered_img_data_5_18 : OUT std_logic ;
      ordered_img_data_5_17 : OUT std_logic ;
      ordered_img_data_5_16 : OUT std_logic ;
      ordered_img_data_5_15 : OUT std_logic ;
      ordered_img_data_5_14 : OUT std_logic ;
      ordered_img_data_5_13 : OUT std_logic ;
      ordered_img_data_5_12 : OUT std_logic ;
      ordered_img_data_5_11 : OUT std_logic ;
      ordered_img_data_5_10 : OUT std_logic ;
      ordered_img_data_5_9 : OUT std_logic ;
      ordered_img_data_5_8 : OUT std_logic ;
      ordered_img_data_5_7 : OUT std_logic ;
      ordered_img_data_5_6 : OUT std_logic ;
      ordered_img_data_5_5 : OUT std_logic ;
      ordered_img_data_5_4 : OUT std_logic ;
      ordered_img_data_5_3 : OUT std_logic ;
      ordered_img_data_5_2 : OUT std_logic ;
      ordered_img_data_5_1 : OUT std_logic ;
      ordered_img_data_5_0 : OUT std_logic ;
      ordered_img_data_6_31 : OUT std_logic ;
      ordered_img_data_6_30 : OUT std_logic ;
      ordered_img_data_6_29 : OUT std_logic ;
      ordered_img_data_6_28 : OUT std_logic ;
      ordered_img_data_6_27 : OUT std_logic ;
      ordered_img_data_6_26 : OUT std_logic ;
      ordered_img_data_6_25 : OUT std_logic ;
      ordered_img_data_6_24 : OUT std_logic ;
      ordered_img_data_6_23 : OUT std_logic ;
      ordered_img_data_6_22 : OUT std_logic ;
      ordered_img_data_6_21 : OUT std_logic ;
      ordered_img_data_6_20 : OUT std_logic ;
      ordered_img_data_6_19 : OUT std_logic ;
      ordered_img_data_6_18 : OUT std_logic ;
      ordered_img_data_6_17 : OUT std_logic ;
      ordered_img_data_6_16 : OUT std_logic ;
      ordered_img_data_6_15 : OUT std_logic ;
      ordered_img_data_6_14 : OUT std_logic ;
      ordered_img_data_6_13 : OUT std_logic ;
      ordered_img_data_6_12 : OUT std_logic ;
      ordered_img_data_6_11 : OUT std_logic ;
      ordered_img_data_6_10 : OUT std_logic ;
      ordered_img_data_6_9 : OUT std_logic ;
      ordered_img_data_6_8 : OUT std_logic ;
      ordered_img_data_6_7 : OUT std_logic ;
      ordered_img_data_6_6 : OUT std_logic ;
      ordered_img_data_6_5 : OUT std_logic ;
      ordered_img_data_6_4 : OUT std_logic ;
      ordered_img_data_6_3 : OUT std_logic ;
      ordered_img_data_6_2 : OUT std_logic ;
      ordered_img_data_6_1 : OUT std_logic ;
      ordered_img_data_6_0 : OUT std_logic ;
      ordered_img_data_7_31 : OUT std_logic ;
      ordered_img_data_7_30 : OUT std_logic ;
      ordered_img_data_7_29 : OUT std_logic ;
      ordered_img_data_7_28 : OUT std_logic ;
      ordered_img_data_7_27 : OUT std_logic ;
      ordered_img_data_7_26 : OUT std_logic ;
      ordered_img_data_7_25 : OUT std_logic ;
      ordered_img_data_7_24 : OUT std_logic ;
      ordered_img_data_7_23 : OUT std_logic ;
      ordered_img_data_7_22 : OUT std_logic ;
      ordered_img_data_7_21 : OUT std_logic ;
      ordered_img_data_7_20 : OUT std_logic ;
      ordered_img_data_7_19 : OUT std_logic ;
      ordered_img_data_7_18 : OUT std_logic ;
      ordered_img_data_7_17 : OUT std_logic ;
      ordered_img_data_7_16 : OUT std_logic ;
      ordered_img_data_7_15 : OUT std_logic ;
      ordered_img_data_7_14 : OUT std_logic ;
      ordered_img_data_7_13 : OUT std_logic ;
      ordered_img_data_7_12 : OUT std_logic ;
      ordered_img_data_7_11 : OUT std_logic ;
      ordered_img_data_7_10 : OUT std_logic ;
      ordered_img_data_7_9 : OUT std_logic ;
      ordered_img_data_7_8 : OUT std_logic ;
      ordered_img_data_7_7 : OUT std_logic ;
      ordered_img_data_7_6 : OUT std_logic ;
      ordered_img_data_7_5 : OUT std_logic ;
      ordered_img_data_7_4 : OUT std_logic ;
      ordered_img_data_7_3 : OUT std_logic ;
      ordered_img_data_7_2 : OUT std_logic ;
      ordered_img_data_7_1 : OUT std_logic ;
      ordered_img_data_7_0 : OUT std_logic ;
      ordered_img_data_8_31 : OUT std_logic ;
      ordered_img_data_8_30 : OUT std_logic ;
      ordered_img_data_8_29 : OUT std_logic ;
      ordered_img_data_8_28 : OUT std_logic ;
      ordered_img_data_8_27 : OUT std_logic ;
      ordered_img_data_8_26 : OUT std_logic ;
      ordered_img_data_8_25 : OUT std_logic ;
      ordered_img_data_8_24 : OUT std_logic ;
      ordered_img_data_8_23 : OUT std_logic ;
      ordered_img_data_8_22 : OUT std_logic ;
      ordered_img_data_8_21 : OUT std_logic ;
      ordered_img_data_8_20 : OUT std_logic ;
      ordered_img_data_8_19 : OUT std_logic ;
      ordered_img_data_8_18 : OUT std_logic ;
      ordered_img_data_8_17 : OUT std_logic ;
      ordered_img_data_8_16 : OUT std_logic ;
      ordered_img_data_8_15 : OUT std_logic ;
      ordered_img_data_8_14 : OUT std_logic ;
      ordered_img_data_8_13 : OUT std_logic ;
      ordered_img_data_8_12 : OUT std_logic ;
      ordered_img_data_8_11 : OUT std_logic ;
      ordered_img_data_8_10 : OUT std_logic ;
      ordered_img_data_8_9 : OUT std_logic ;
      ordered_img_data_8_8 : OUT std_logic ;
      ordered_img_data_8_7 : OUT std_logic ;
      ordered_img_data_8_6 : OUT std_logic ;
      ordered_img_data_8_5 : OUT std_logic ;
      ordered_img_data_8_4 : OUT std_logic ;
      ordered_img_data_8_3 : OUT std_logic ;
      ordered_img_data_8_2 : OUT std_logic ;
      ordered_img_data_8_1 : OUT std_logic ;
      ordered_img_data_8_0 : OUT std_logic ;
      ordered_img_data_9_31 : OUT std_logic ;
      ordered_img_data_9_30 : OUT std_logic ;
      ordered_img_data_9_29 : OUT std_logic ;
      ordered_img_data_9_28 : OUT std_logic ;
      ordered_img_data_9_27 : OUT std_logic ;
      ordered_img_data_9_26 : OUT std_logic ;
      ordered_img_data_9_25 : OUT std_logic ;
      ordered_img_data_9_24 : OUT std_logic ;
      ordered_img_data_9_23 : OUT std_logic ;
      ordered_img_data_9_22 : OUT std_logic ;
      ordered_img_data_9_21 : OUT std_logic ;
      ordered_img_data_9_20 : OUT std_logic ;
      ordered_img_data_9_19 : OUT std_logic ;
      ordered_img_data_9_18 : OUT std_logic ;
      ordered_img_data_9_17 : OUT std_logic ;
      ordered_img_data_9_16 : OUT std_logic ;
      ordered_img_data_9_15 : OUT std_logic ;
      ordered_img_data_9_14 : OUT std_logic ;
      ordered_img_data_9_13 : OUT std_logic ;
      ordered_img_data_9_12 : OUT std_logic ;
      ordered_img_data_9_11 : OUT std_logic ;
      ordered_img_data_9_10 : OUT std_logic ;
      ordered_img_data_9_9 : OUT std_logic ;
      ordered_img_data_9_8 : OUT std_logic ;
      ordered_img_data_9_7 : OUT std_logic ;
      ordered_img_data_9_6 : OUT std_logic ;
      ordered_img_data_9_5 : OUT std_logic ;
      ordered_img_data_9_4 : OUT std_logic ;
      ordered_img_data_9_3 : OUT std_logic ;
      ordered_img_data_9_2 : OUT std_logic ;
      ordered_img_data_9_1 : OUT std_logic ;
      ordered_img_data_9_0 : OUT std_logic ;
      ordered_img_data_10_31 : OUT std_logic ;
      ordered_img_data_10_30 : OUT std_logic ;
      ordered_img_data_10_29 : OUT std_logic ;
      ordered_img_data_10_28 : OUT std_logic ;
      ordered_img_data_10_27 : OUT std_logic ;
      ordered_img_data_10_26 : OUT std_logic ;
      ordered_img_data_10_25 : OUT std_logic ;
      ordered_img_data_10_24 : OUT std_logic ;
      ordered_img_data_10_23 : OUT std_logic ;
      ordered_img_data_10_22 : OUT std_logic ;
      ordered_img_data_10_21 : OUT std_logic ;
      ordered_img_data_10_20 : OUT std_logic ;
      ordered_img_data_10_19 : OUT std_logic ;
      ordered_img_data_10_18 : OUT std_logic ;
      ordered_img_data_10_17 : OUT std_logic ;
      ordered_img_data_10_16 : OUT std_logic ;
      ordered_img_data_10_15 : OUT std_logic ;
      ordered_img_data_10_14 : OUT std_logic ;
      ordered_img_data_10_13 : OUT std_logic ;
      ordered_img_data_10_12 : OUT std_logic ;
      ordered_img_data_10_11 : OUT std_logic ;
      ordered_img_data_10_10 : OUT std_logic ;
      ordered_img_data_10_9 : OUT std_logic ;
      ordered_img_data_10_8 : OUT std_logic ;
      ordered_img_data_10_7 : OUT std_logic ;
      ordered_img_data_10_6 : OUT std_logic ;
      ordered_img_data_10_5 : OUT std_logic ;
      ordered_img_data_10_4 : OUT std_logic ;
      ordered_img_data_10_3 : OUT std_logic ;
      ordered_img_data_10_2 : OUT std_logic ;
      ordered_img_data_10_1 : OUT std_logic ;
      ordered_img_data_10_0 : OUT std_logic ;
      ordered_img_data_11_31 : OUT std_logic ;
      ordered_img_data_11_30 : OUT std_logic ;
      ordered_img_data_11_29 : OUT std_logic ;
      ordered_img_data_11_28 : OUT std_logic ;
      ordered_img_data_11_27 : OUT std_logic ;
      ordered_img_data_11_26 : OUT std_logic ;
      ordered_img_data_11_25 : OUT std_logic ;
      ordered_img_data_11_24 : OUT std_logic ;
      ordered_img_data_11_23 : OUT std_logic ;
      ordered_img_data_11_22 : OUT std_logic ;
      ordered_img_data_11_21 : OUT std_logic ;
      ordered_img_data_11_20 : OUT std_logic ;
      ordered_img_data_11_19 : OUT std_logic ;
      ordered_img_data_11_18 : OUT std_logic ;
      ordered_img_data_11_17 : OUT std_logic ;
      ordered_img_data_11_16 : OUT std_logic ;
      ordered_img_data_11_15 : OUT std_logic ;
      ordered_img_data_11_14 : OUT std_logic ;
      ordered_img_data_11_13 : OUT std_logic ;
      ordered_img_data_11_12 : OUT std_logic ;
      ordered_img_data_11_11 : OUT std_logic ;
      ordered_img_data_11_10 : OUT std_logic ;
      ordered_img_data_11_9 : OUT std_logic ;
      ordered_img_data_11_8 : OUT std_logic ;
      ordered_img_data_11_7 : OUT std_logic ;
      ordered_img_data_11_6 : OUT std_logic ;
      ordered_img_data_11_5 : OUT std_logic ;
      ordered_img_data_11_4 : OUT std_logic ;
      ordered_img_data_11_3 : OUT std_logic ;
      ordered_img_data_11_2 : OUT std_logic ;
      ordered_img_data_11_1 : OUT std_logic ;
      ordered_img_data_11_0 : OUT std_logic ;
      ordered_img_data_12_31 : OUT std_logic ;
      ordered_img_data_12_30 : OUT std_logic ;
      ordered_img_data_12_29 : OUT std_logic ;
      ordered_img_data_12_28 : OUT std_logic ;
      ordered_img_data_12_27 : OUT std_logic ;
      ordered_img_data_12_26 : OUT std_logic ;
      ordered_img_data_12_25 : OUT std_logic ;
      ordered_img_data_12_24 : OUT std_logic ;
      ordered_img_data_12_23 : OUT std_logic ;
      ordered_img_data_12_22 : OUT std_logic ;
      ordered_img_data_12_21 : OUT std_logic ;
      ordered_img_data_12_20 : OUT std_logic ;
      ordered_img_data_12_19 : OUT std_logic ;
      ordered_img_data_12_18 : OUT std_logic ;
      ordered_img_data_12_17 : OUT std_logic ;
      ordered_img_data_12_16 : OUT std_logic ;
      ordered_img_data_12_15 : OUT std_logic ;
      ordered_img_data_12_14 : OUT std_logic ;
      ordered_img_data_12_13 : OUT std_logic ;
      ordered_img_data_12_12 : OUT std_logic ;
      ordered_img_data_12_11 : OUT std_logic ;
      ordered_img_data_12_10 : OUT std_logic ;
      ordered_img_data_12_9 : OUT std_logic ;
      ordered_img_data_12_8 : OUT std_logic ;
      ordered_img_data_12_7 : OUT std_logic ;
      ordered_img_data_12_6 : OUT std_logic ;
      ordered_img_data_12_5 : OUT std_logic ;
      ordered_img_data_12_4 : OUT std_logic ;
      ordered_img_data_12_3 : OUT std_logic ;
      ordered_img_data_12_2 : OUT std_logic ;
      ordered_img_data_12_1 : OUT std_logic ;
      ordered_img_data_12_0 : OUT std_logic ;
      ordered_img_data_13_31 : OUT std_logic ;
      ordered_img_data_13_30 : OUT std_logic ;
      ordered_img_data_13_29 : OUT std_logic ;
      ordered_img_data_13_28 : OUT std_logic ;
      ordered_img_data_13_27 : OUT std_logic ;
      ordered_img_data_13_26 : OUT std_logic ;
      ordered_img_data_13_25 : OUT std_logic ;
      ordered_img_data_13_24 : OUT std_logic ;
      ordered_img_data_13_23 : OUT std_logic ;
      ordered_img_data_13_22 : OUT std_logic ;
      ordered_img_data_13_21 : OUT std_logic ;
      ordered_img_data_13_20 : OUT std_logic ;
      ordered_img_data_13_19 : OUT std_logic ;
      ordered_img_data_13_18 : OUT std_logic ;
      ordered_img_data_13_17 : OUT std_logic ;
      ordered_img_data_13_16 : OUT std_logic ;
      ordered_img_data_13_15 : OUT std_logic ;
      ordered_img_data_13_14 : OUT std_logic ;
      ordered_img_data_13_13 : OUT std_logic ;
      ordered_img_data_13_12 : OUT std_logic ;
      ordered_img_data_13_11 : OUT std_logic ;
      ordered_img_data_13_10 : OUT std_logic ;
      ordered_img_data_13_9 : OUT std_logic ;
      ordered_img_data_13_8 : OUT std_logic ;
      ordered_img_data_13_7 : OUT std_logic ;
      ordered_img_data_13_6 : OUT std_logic ;
      ordered_img_data_13_5 : OUT std_logic ;
      ordered_img_data_13_4 : OUT std_logic ;
      ordered_img_data_13_3 : OUT std_logic ;
      ordered_img_data_13_2 : OUT std_logic ;
      ordered_img_data_13_1 : OUT std_logic ;
      ordered_img_data_13_0 : OUT std_logic ;
      ordered_img_data_14_31 : OUT std_logic ;
      ordered_img_data_14_30 : OUT std_logic ;
      ordered_img_data_14_29 : OUT std_logic ;
      ordered_img_data_14_28 : OUT std_logic ;
      ordered_img_data_14_27 : OUT std_logic ;
      ordered_img_data_14_26 : OUT std_logic ;
      ordered_img_data_14_25 : OUT std_logic ;
      ordered_img_data_14_24 : OUT std_logic ;
      ordered_img_data_14_23 : OUT std_logic ;
      ordered_img_data_14_22 : OUT std_logic ;
      ordered_img_data_14_21 : OUT std_logic ;
      ordered_img_data_14_20 : OUT std_logic ;
      ordered_img_data_14_19 : OUT std_logic ;
      ordered_img_data_14_18 : OUT std_logic ;
      ordered_img_data_14_17 : OUT std_logic ;
      ordered_img_data_14_16 : OUT std_logic ;
      ordered_img_data_14_15 : OUT std_logic ;
      ordered_img_data_14_14 : OUT std_logic ;
      ordered_img_data_14_13 : OUT std_logic ;
      ordered_img_data_14_12 : OUT std_logic ;
      ordered_img_data_14_11 : OUT std_logic ;
      ordered_img_data_14_10 : OUT std_logic ;
      ordered_img_data_14_9 : OUT std_logic ;
      ordered_img_data_14_8 : OUT std_logic ;
      ordered_img_data_14_7 : OUT std_logic ;
      ordered_img_data_14_6 : OUT std_logic ;
      ordered_img_data_14_5 : OUT std_logic ;
      ordered_img_data_14_4 : OUT std_logic ;
      ordered_img_data_14_3 : OUT std_logic ;
      ordered_img_data_14_2 : OUT std_logic ;
      ordered_img_data_14_1 : OUT std_logic ;
      ordered_img_data_14_0 : OUT std_logic ;
      ordered_img_data_15_31 : OUT std_logic ;
      ordered_img_data_15_30 : OUT std_logic ;
      ordered_img_data_15_29 : OUT std_logic ;
      ordered_img_data_15_28 : OUT std_logic ;
      ordered_img_data_15_27 : OUT std_logic ;
      ordered_img_data_15_26 : OUT std_logic ;
      ordered_img_data_15_25 : OUT std_logic ;
      ordered_img_data_15_24 : OUT std_logic ;
      ordered_img_data_15_23 : OUT std_logic ;
      ordered_img_data_15_22 : OUT std_logic ;
      ordered_img_data_15_21 : OUT std_logic ;
      ordered_img_data_15_20 : OUT std_logic ;
      ordered_img_data_15_19 : OUT std_logic ;
      ordered_img_data_15_18 : OUT std_logic ;
      ordered_img_data_15_17 : OUT std_logic ;
      ordered_img_data_15_16 : OUT std_logic ;
      ordered_img_data_15_15 : OUT std_logic ;
      ordered_img_data_15_14 : OUT std_logic ;
      ordered_img_data_15_13 : OUT std_logic ;
      ordered_img_data_15_12 : OUT std_logic ;
      ordered_img_data_15_11 : OUT std_logic ;
      ordered_img_data_15_10 : OUT std_logic ;
      ordered_img_data_15_9 : OUT std_logic ;
      ordered_img_data_15_8 : OUT std_logic ;
      ordered_img_data_15_7 : OUT std_logic ;
      ordered_img_data_15_6 : OUT std_logic ;
      ordered_img_data_15_5 : OUT std_logic ;
      ordered_img_data_15_4 : OUT std_logic ;
      ordered_img_data_15_3 : OUT std_logic ;
      ordered_img_data_15_2 : OUT std_logic ;
      ordered_img_data_15_1 : OUT std_logic ;
      ordered_img_data_15_0 : OUT std_logic ;
      ordered_img_data_16_31 : OUT std_logic ;
      ordered_img_data_16_30 : OUT std_logic ;
      ordered_img_data_16_29 : OUT std_logic ;
      ordered_img_data_16_28 : OUT std_logic ;
      ordered_img_data_16_27 : OUT std_logic ;
      ordered_img_data_16_26 : OUT std_logic ;
      ordered_img_data_16_25 : OUT std_logic ;
      ordered_img_data_16_24 : OUT std_logic ;
      ordered_img_data_16_23 : OUT std_logic ;
      ordered_img_data_16_22 : OUT std_logic ;
      ordered_img_data_16_21 : OUT std_logic ;
      ordered_img_data_16_20 : OUT std_logic ;
      ordered_img_data_16_19 : OUT std_logic ;
      ordered_img_data_16_18 : OUT std_logic ;
      ordered_img_data_16_17 : OUT std_logic ;
      ordered_img_data_16_16 : OUT std_logic ;
      ordered_img_data_16_15 : OUT std_logic ;
      ordered_img_data_16_14 : OUT std_logic ;
      ordered_img_data_16_13 : OUT std_logic ;
      ordered_img_data_16_12 : OUT std_logic ;
      ordered_img_data_16_11 : OUT std_logic ;
      ordered_img_data_16_10 : OUT std_logic ;
      ordered_img_data_16_9 : OUT std_logic ;
      ordered_img_data_16_8 : OUT std_logic ;
      ordered_img_data_16_7 : OUT std_logic ;
      ordered_img_data_16_6 : OUT std_logic ;
      ordered_img_data_16_5 : OUT std_logic ;
      ordered_img_data_16_4 : OUT std_logic ;
      ordered_img_data_16_3 : OUT std_logic ;
      ordered_img_data_16_2 : OUT std_logic ;
      ordered_img_data_16_1 : OUT std_logic ;
      ordered_img_data_16_0 : OUT std_logic ;
      ordered_img_data_17_31 : OUT std_logic ;
      ordered_img_data_17_30 : OUT std_logic ;
      ordered_img_data_17_29 : OUT std_logic ;
      ordered_img_data_17_28 : OUT std_logic ;
      ordered_img_data_17_27 : OUT std_logic ;
      ordered_img_data_17_26 : OUT std_logic ;
      ordered_img_data_17_25 : OUT std_logic ;
      ordered_img_data_17_24 : OUT std_logic ;
      ordered_img_data_17_23 : OUT std_logic ;
      ordered_img_data_17_22 : OUT std_logic ;
      ordered_img_data_17_21 : OUT std_logic ;
      ordered_img_data_17_20 : OUT std_logic ;
      ordered_img_data_17_19 : OUT std_logic ;
      ordered_img_data_17_18 : OUT std_logic ;
      ordered_img_data_17_17 : OUT std_logic ;
      ordered_img_data_17_16 : OUT std_logic ;
      ordered_img_data_17_15 : OUT std_logic ;
      ordered_img_data_17_14 : OUT std_logic ;
      ordered_img_data_17_13 : OUT std_logic ;
      ordered_img_data_17_12 : OUT std_logic ;
      ordered_img_data_17_11 : OUT std_logic ;
      ordered_img_data_17_10 : OUT std_logic ;
      ordered_img_data_17_9 : OUT std_logic ;
      ordered_img_data_17_8 : OUT std_logic ;
      ordered_img_data_17_7 : OUT std_logic ;
      ordered_img_data_17_6 : OUT std_logic ;
      ordered_img_data_17_5 : OUT std_logic ;
      ordered_img_data_17_4 : OUT std_logic ;
      ordered_img_data_17_3 : OUT std_logic ;
      ordered_img_data_17_2 : OUT std_logic ;
      ordered_img_data_17_1 : OUT std_logic ;
      ordered_img_data_17_0 : OUT std_logic ;
      ordered_img_data_18_31 : OUT std_logic ;
      ordered_img_data_18_30 : OUT std_logic ;
      ordered_img_data_18_29 : OUT std_logic ;
      ordered_img_data_18_28 : OUT std_logic ;
      ordered_img_data_18_27 : OUT std_logic ;
      ordered_img_data_18_26 : OUT std_logic ;
      ordered_img_data_18_25 : OUT std_logic ;
      ordered_img_data_18_24 : OUT std_logic ;
      ordered_img_data_18_23 : OUT std_logic ;
      ordered_img_data_18_22 : OUT std_logic ;
      ordered_img_data_18_21 : OUT std_logic ;
      ordered_img_data_18_20 : OUT std_logic ;
      ordered_img_data_18_19 : OUT std_logic ;
      ordered_img_data_18_18 : OUT std_logic ;
      ordered_img_data_18_17 : OUT std_logic ;
      ordered_img_data_18_16 : OUT std_logic ;
      ordered_img_data_18_15 : OUT std_logic ;
      ordered_img_data_18_14 : OUT std_logic ;
      ordered_img_data_18_13 : OUT std_logic ;
      ordered_img_data_18_12 : OUT std_logic ;
      ordered_img_data_18_11 : OUT std_logic ;
      ordered_img_data_18_10 : OUT std_logic ;
      ordered_img_data_18_9 : OUT std_logic ;
      ordered_img_data_18_8 : OUT std_logic ;
      ordered_img_data_18_7 : OUT std_logic ;
      ordered_img_data_18_6 : OUT std_logic ;
      ordered_img_data_18_5 : OUT std_logic ;
      ordered_img_data_18_4 : OUT std_logic ;
      ordered_img_data_18_3 : OUT std_logic ;
      ordered_img_data_18_2 : OUT std_logic ;
      ordered_img_data_18_1 : OUT std_logic ;
      ordered_img_data_18_0 : OUT std_logic ;
      ordered_img_data_19_31 : OUT std_logic ;
      ordered_img_data_19_30 : OUT std_logic ;
      ordered_img_data_19_29 : OUT std_logic ;
      ordered_img_data_19_28 : OUT std_logic ;
      ordered_img_data_19_27 : OUT std_logic ;
      ordered_img_data_19_26 : OUT std_logic ;
      ordered_img_data_19_25 : OUT std_logic ;
      ordered_img_data_19_24 : OUT std_logic ;
      ordered_img_data_19_23 : OUT std_logic ;
      ordered_img_data_19_22 : OUT std_logic ;
      ordered_img_data_19_21 : OUT std_logic ;
      ordered_img_data_19_20 : OUT std_logic ;
      ordered_img_data_19_19 : OUT std_logic ;
      ordered_img_data_19_18 : OUT std_logic ;
      ordered_img_data_19_17 : OUT std_logic ;
      ordered_img_data_19_16 : OUT std_logic ;
      ordered_img_data_19_15 : OUT std_logic ;
      ordered_img_data_19_14 : OUT std_logic ;
      ordered_img_data_19_13 : OUT std_logic ;
      ordered_img_data_19_12 : OUT std_logic ;
      ordered_img_data_19_11 : OUT std_logic ;
      ordered_img_data_19_10 : OUT std_logic ;
      ordered_img_data_19_9 : OUT std_logic ;
      ordered_img_data_19_8 : OUT std_logic ;
      ordered_img_data_19_7 : OUT std_logic ;
      ordered_img_data_19_6 : OUT std_logic ;
      ordered_img_data_19_5 : OUT std_logic ;
      ordered_img_data_19_4 : OUT std_logic ;
      ordered_img_data_19_3 : OUT std_logic ;
      ordered_img_data_19_2 : OUT std_logic ;
      ordered_img_data_19_1 : OUT std_logic ;
      ordered_img_data_19_0 : OUT std_logic ;
      ordered_img_data_20_31 : OUT std_logic ;
      ordered_img_data_20_30 : OUT std_logic ;
      ordered_img_data_20_29 : OUT std_logic ;
      ordered_img_data_20_28 : OUT std_logic ;
      ordered_img_data_20_27 : OUT std_logic ;
      ordered_img_data_20_26 : OUT std_logic ;
      ordered_img_data_20_25 : OUT std_logic ;
      ordered_img_data_20_24 : OUT std_logic ;
      ordered_img_data_20_23 : OUT std_logic ;
      ordered_img_data_20_22 : OUT std_logic ;
      ordered_img_data_20_21 : OUT std_logic ;
      ordered_img_data_20_20 : OUT std_logic ;
      ordered_img_data_20_19 : OUT std_logic ;
      ordered_img_data_20_18 : OUT std_logic ;
      ordered_img_data_20_17 : OUT std_logic ;
      ordered_img_data_20_16 : OUT std_logic ;
      ordered_img_data_20_15 : OUT std_logic ;
      ordered_img_data_20_14 : OUT std_logic ;
      ordered_img_data_20_13 : OUT std_logic ;
      ordered_img_data_20_12 : OUT std_logic ;
      ordered_img_data_20_11 : OUT std_logic ;
      ordered_img_data_20_10 : OUT std_logic ;
      ordered_img_data_20_9 : OUT std_logic ;
      ordered_img_data_20_8 : OUT std_logic ;
      ordered_img_data_20_7 : OUT std_logic ;
      ordered_img_data_20_6 : OUT std_logic ;
      ordered_img_data_20_5 : OUT std_logic ;
      ordered_img_data_20_4 : OUT std_logic ;
      ordered_img_data_20_3 : OUT std_logic ;
      ordered_img_data_20_2 : OUT std_logic ;
      ordered_img_data_20_1 : OUT std_logic ;
      ordered_img_data_20_0 : OUT std_logic ;
      ordered_img_data_21_31 : OUT std_logic ;
      ordered_img_data_21_30 : OUT std_logic ;
      ordered_img_data_21_29 : OUT std_logic ;
      ordered_img_data_21_28 : OUT std_logic ;
      ordered_img_data_21_27 : OUT std_logic ;
      ordered_img_data_21_26 : OUT std_logic ;
      ordered_img_data_21_25 : OUT std_logic ;
      ordered_img_data_21_24 : OUT std_logic ;
      ordered_img_data_21_23 : OUT std_logic ;
      ordered_img_data_21_22 : OUT std_logic ;
      ordered_img_data_21_21 : OUT std_logic ;
      ordered_img_data_21_20 : OUT std_logic ;
      ordered_img_data_21_19 : OUT std_logic ;
      ordered_img_data_21_18 : OUT std_logic ;
      ordered_img_data_21_17 : OUT std_logic ;
      ordered_img_data_21_16 : OUT std_logic ;
      ordered_img_data_21_15 : OUT std_logic ;
      ordered_img_data_21_14 : OUT std_logic ;
      ordered_img_data_21_13 : OUT std_logic ;
      ordered_img_data_21_12 : OUT std_logic ;
      ordered_img_data_21_11 : OUT std_logic ;
      ordered_img_data_21_10 : OUT std_logic ;
      ordered_img_data_21_9 : OUT std_logic ;
      ordered_img_data_21_8 : OUT std_logic ;
      ordered_img_data_21_7 : OUT std_logic ;
      ordered_img_data_21_6 : OUT std_logic ;
      ordered_img_data_21_5 : OUT std_logic ;
      ordered_img_data_21_4 : OUT std_logic ;
      ordered_img_data_21_3 : OUT std_logic ;
      ordered_img_data_21_2 : OUT std_logic ;
      ordered_img_data_21_1 : OUT std_logic ;
      ordered_img_data_21_0 : OUT std_logic ;
      ordered_img_data_22_31 : OUT std_logic ;
      ordered_img_data_22_30 : OUT std_logic ;
      ordered_img_data_22_29 : OUT std_logic ;
      ordered_img_data_22_28 : OUT std_logic ;
      ordered_img_data_22_27 : OUT std_logic ;
      ordered_img_data_22_26 : OUT std_logic ;
      ordered_img_data_22_25 : OUT std_logic ;
      ordered_img_data_22_24 : OUT std_logic ;
      ordered_img_data_22_23 : OUT std_logic ;
      ordered_img_data_22_22 : OUT std_logic ;
      ordered_img_data_22_21 : OUT std_logic ;
      ordered_img_data_22_20 : OUT std_logic ;
      ordered_img_data_22_19 : OUT std_logic ;
      ordered_img_data_22_18 : OUT std_logic ;
      ordered_img_data_22_17 : OUT std_logic ;
      ordered_img_data_22_16 : OUT std_logic ;
      ordered_img_data_22_15 : OUT std_logic ;
      ordered_img_data_22_14 : OUT std_logic ;
      ordered_img_data_22_13 : OUT std_logic ;
      ordered_img_data_22_12 : OUT std_logic ;
      ordered_img_data_22_11 : OUT std_logic ;
      ordered_img_data_22_10 : OUT std_logic ;
      ordered_img_data_22_9 : OUT std_logic ;
      ordered_img_data_22_8 : OUT std_logic ;
      ordered_img_data_22_7 : OUT std_logic ;
      ordered_img_data_22_6 : OUT std_logic ;
      ordered_img_data_22_5 : OUT std_logic ;
      ordered_img_data_22_4 : OUT std_logic ;
      ordered_img_data_22_3 : OUT std_logic ;
      ordered_img_data_22_2 : OUT std_logic ;
      ordered_img_data_22_1 : OUT std_logic ;
      ordered_img_data_22_0 : OUT std_logic ;
      ordered_img_data_23_31 : OUT std_logic ;
      ordered_img_data_23_30 : OUT std_logic ;
      ordered_img_data_23_29 : OUT std_logic ;
      ordered_img_data_23_28 : OUT std_logic ;
      ordered_img_data_23_27 : OUT std_logic ;
      ordered_img_data_23_26 : OUT std_logic ;
      ordered_img_data_23_25 : OUT std_logic ;
      ordered_img_data_23_24 : OUT std_logic ;
      ordered_img_data_23_23 : OUT std_logic ;
      ordered_img_data_23_22 : OUT std_logic ;
      ordered_img_data_23_21 : OUT std_logic ;
      ordered_img_data_23_20 : OUT std_logic ;
      ordered_img_data_23_19 : OUT std_logic ;
      ordered_img_data_23_18 : OUT std_logic ;
      ordered_img_data_23_17 : OUT std_logic ;
      ordered_img_data_23_16 : OUT std_logic ;
      ordered_img_data_23_15 : OUT std_logic ;
      ordered_img_data_23_14 : OUT std_logic ;
      ordered_img_data_23_13 : OUT std_logic ;
      ordered_img_data_23_12 : OUT std_logic ;
      ordered_img_data_23_11 : OUT std_logic ;
      ordered_img_data_23_10 : OUT std_logic ;
      ordered_img_data_23_9 : OUT std_logic ;
      ordered_img_data_23_8 : OUT std_logic ;
      ordered_img_data_23_7 : OUT std_logic ;
      ordered_img_data_23_6 : OUT std_logic ;
      ordered_img_data_23_5 : OUT std_logic ;
      ordered_img_data_23_4 : OUT std_logic ;
      ordered_img_data_23_3 : OUT std_logic ;
      ordered_img_data_23_2 : OUT std_logic ;
      ordered_img_data_23_1 : OUT std_logic ;
      ordered_img_data_23_0 : OUT std_logic ;
      ordered_img_data_24_31 : OUT std_logic ;
      ordered_img_data_24_30 : OUT std_logic ;
      ordered_img_data_24_29 : OUT std_logic ;
      ordered_img_data_24_28 : OUT std_logic ;
      ordered_img_data_24_27 : OUT std_logic ;
      ordered_img_data_24_26 : OUT std_logic ;
      ordered_img_data_24_25 : OUT std_logic ;
      ordered_img_data_24_24 : OUT std_logic ;
      ordered_img_data_24_23 : OUT std_logic ;
      ordered_img_data_24_22 : OUT std_logic ;
      ordered_img_data_24_21 : OUT std_logic ;
      ordered_img_data_24_20 : OUT std_logic ;
      ordered_img_data_24_19 : OUT std_logic ;
      ordered_img_data_24_18 : OUT std_logic ;
      ordered_img_data_24_17 : OUT std_logic ;
      ordered_img_data_24_16 : OUT std_logic ;
      ordered_img_data_24_15 : OUT std_logic ;
      ordered_img_data_24_14 : OUT std_logic ;
      ordered_img_data_24_13 : OUT std_logic ;
      ordered_img_data_24_12 : OUT std_logic ;
      ordered_img_data_24_11 : OUT std_logic ;
      ordered_img_data_24_10 : OUT std_logic ;
      ordered_img_data_24_9 : OUT std_logic ;
      ordered_img_data_24_8 : OUT std_logic ;
      ordered_img_data_24_7 : OUT std_logic ;
      ordered_img_data_24_6 : OUT std_logic ;
      ordered_img_data_24_5 : OUT std_logic ;
      ordered_img_data_24_4 : OUT std_logic ;
      ordered_img_data_24_3 : OUT std_logic ;
      ordered_img_data_24_2 : OUT std_logic ;
      ordered_img_data_24_1 : OUT std_logic ;
      ordered_img_data_24_0 : OUT std_logic ;
      ordered_filter_data_0_31 : OUT std_logic ;
      ordered_filter_data_0_30 : OUT std_logic ;
      ordered_filter_data_0_29 : OUT std_logic ;
      ordered_filter_data_0_28 : OUT std_logic ;
      ordered_filter_data_0_27 : OUT std_logic ;
      ordered_filter_data_0_26 : OUT std_logic ;
      ordered_filter_data_0_25 : OUT std_logic ;
      ordered_filter_data_0_24 : OUT std_logic ;
      ordered_filter_data_0_23 : OUT std_logic ;
      ordered_filter_data_0_22 : OUT std_logic ;
      ordered_filter_data_0_21 : OUT std_logic ;
      ordered_filter_data_0_20 : OUT std_logic ;
      ordered_filter_data_0_19 : OUT std_logic ;
      ordered_filter_data_0_18 : OUT std_logic ;
      ordered_filter_data_0_17 : OUT std_logic ;
      ordered_filter_data_0_16 : OUT std_logic ;
      ordered_filter_data_0_15 : OUT std_logic ;
      ordered_filter_data_0_14 : OUT std_logic ;
      ordered_filter_data_0_13 : OUT std_logic ;
      ordered_filter_data_0_12 : OUT std_logic ;
      ordered_filter_data_0_11 : OUT std_logic ;
      ordered_filter_data_0_10 : OUT std_logic ;
      ordered_filter_data_0_9 : OUT std_logic ;
      ordered_filter_data_0_8 : OUT std_logic ;
      ordered_filter_data_0_7 : OUT std_logic ;
      ordered_filter_data_0_6 : OUT std_logic ;
      ordered_filter_data_0_5 : OUT std_logic ;
      ordered_filter_data_0_4 : OUT std_logic ;
      ordered_filter_data_0_3 : OUT std_logic ;
      ordered_filter_data_0_2 : OUT std_logic ;
      ordered_filter_data_0_1 : OUT std_logic ;
      ordered_filter_data_0_0 : OUT std_logic ;
      ordered_filter_data_1_31 : OUT std_logic ;
      ordered_filter_data_1_30 : OUT std_logic ;
      ordered_filter_data_1_29 : OUT std_logic ;
      ordered_filter_data_1_28 : OUT std_logic ;
      ordered_filter_data_1_27 : OUT std_logic ;
      ordered_filter_data_1_26 : OUT std_logic ;
      ordered_filter_data_1_25 : OUT std_logic ;
      ordered_filter_data_1_24 : OUT std_logic ;
      ordered_filter_data_1_23 : OUT std_logic ;
      ordered_filter_data_1_22 : OUT std_logic ;
      ordered_filter_data_1_21 : OUT std_logic ;
      ordered_filter_data_1_20 : OUT std_logic ;
      ordered_filter_data_1_19 : OUT std_logic ;
      ordered_filter_data_1_18 : OUT std_logic ;
      ordered_filter_data_1_17 : OUT std_logic ;
      ordered_filter_data_1_16 : OUT std_logic ;
      ordered_filter_data_1_15 : OUT std_logic ;
      ordered_filter_data_1_14 : OUT std_logic ;
      ordered_filter_data_1_13 : OUT std_logic ;
      ordered_filter_data_1_12 : OUT std_logic ;
      ordered_filter_data_1_11 : OUT std_logic ;
      ordered_filter_data_1_10 : OUT std_logic ;
      ordered_filter_data_1_9 : OUT std_logic ;
      ordered_filter_data_1_8 : OUT std_logic ;
      ordered_filter_data_1_7 : OUT std_logic ;
      ordered_filter_data_1_6 : OUT std_logic ;
      ordered_filter_data_1_5 : OUT std_logic ;
      ordered_filter_data_1_4 : OUT std_logic ;
      ordered_filter_data_1_3 : OUT std_logic ;
      ordered_filter_data_1_2 : OUT std_logic ;
      ordered_filter_data_1_1 : OUT std_logic ;
      ordered_filter_data_1_0 : OUT std_logic ;
      ordered_filter_data_2_31 : OUT std_logic ;
      ordered_filter_data_2_30 : OUT std_logic ;
      ordered_filter_data_2_29 : OUT std_logic ;
      ordered_filter_data_2_28 : OUT std_logic ;
      ordered_filter_data_2_27 : OUT std_logic ;
      ordered_filter_data_2_26 : OUT std_logic ;
      ordered_filter_data_2_25 : OUT std_logic ;
      ordered_filter_data_2_24 : OUT std_logic ;
      ordered_filter_data_2_23 : OUT std_logic ;
      ordered_filter_data_2_22 : OUT std_logic ;
      ordered_filter_data_2_21 : OUT std_logic ;
      ordered_filter_data_2_20 : OUT std_logic ;
      ordered_filter_data_2_19 : OUT std_logic ;
      ordered_filter_data_2_18 : OUT std_logic ;
      ordered_filter_data_2_17 : OUT std_logic ;
      ordered_filter_data_2_16 : OUT std_logic ;
      ordered_filter_data_2_15 : OUT std_logic ;
      ordered_filter_data_2_14 : OUT std_logic ;
      ordered_filter_data_2_13 : OUT std_logic ;
      ordered_filter_data_2_12 : OUT std_logic ;
      ordered_filter_data_2_11 : OUT std_logic ;
      ordered_filter_data_2_10 : OUT std_logic ;
      ordered_filter_data_2_9 : OUT std_logic ;
      ordered_filter_data_2_8 : OUT std_logic ;
      ordered_filter_data_2_7 : OUT std_logic ;
      ordered_filter_data_2_6 : OUT std_logic ;
      ordered_filter_data_2_5 : OUT std_logic ;
      ordered_filter_data_2_4 : OUT std_logic ;
      ordered_filter_data_2_3 : OUT std_logic ;
      ordered_filter_data_2_2 : OUT std_logic ;
      ordered_filter_data_2_1 : OUT std_logic ;
      ordered_filter_data_2_0 : OUT std_logic ;
      ordered_filter_data_3_31 : OUT std_logic ;
      ordered_filter_data_3_30 : OUT std_logic ;
      ordered_filter_data_3_29 : OUT std_logic ;
      ordered_filter_data_3_28 : OUT std_logic ;
      ordered_filter_data_3_27 : OUT std_logic ;
      ordered_filter_data_3_26 : OUT std_logic ;
      ordered_filter_data_3_25 : OUT std_logic ;
      ordered_filter_data_3_24 : OUT std_logic ;
      ordered_filter_data_3_23 : OUT std_logic ;
      ordered_filter_data_3_22 : OUT std_logic ;
      ordered_filter_data_3_21 : OUT std_logic ;
      ordered_filter_data_3_20 : OUT std_logic ;
      ordered_filter_data_3_19 : OUT std_logic ;
      ordered_filter_data_3_18 : OUT std_logic ;
      ordered_filter_data_3_17 : OUT std_logic ;
      ordered_filter_data_3_16 : OUT std_logic ;
      ordered_filter_data_3_15 : OUT std_logic ;
      ordered_filter_data_3_14 : OUT std_logic ;
      ordered_filter_data_3_13 : OUT std_logic ;
      ordered_filter_data_3_12 : OUT std_logic ;
      ordered_filter_data_3_11 : OUT std_logic ;
      ordered_filter_data_3_10 : OUT std_logic ;
      ordered_filter_data_3_9 : OUT std_logic ;
      ordered_filter_data_3_8 : OUT std_logic ;
      ordered_filter_data_3_7 : OUT std_logic ;
      ordered_filter_data_3_6 : OUT std_logic ;
      ordered_filter_data_3_5 : OUT std_logic ;
      ordered_filter_data_3_4 : OUT std_logic ;
      ordered_filter_data_3_3 : OUT std_logic ;
      ordered_filter_data_3_2 : OUT std_logic ;
      ordered_filter_data_3_1 : OUT std_logic ;
      ordered_filter_data_3_0 : OUT std_logic ;
      ordered_filter_data_4_31 : OUT std_logic ;
      ordered_filter_data_4_30 : OUT std_logic ;
      ordered_filter_data_4_29 : OUT std_logic ;
      ordered_filter_data_4_28 : OUT std_logic ;
      ordered_filter_data_4_27 : OUT std_logic ;
      ordered_filter_data_4_26 : OUT std_logic ;
      ordered_filter_data_4_25 : OUT std_logic ;
      ordered_filter_data_4_24 : OUT std_logic ;
      ordered_filter_data_4_23 : OUT std_logic ;
      ordered_filter_data_4_22 : OUT std_logic ;
      ordered_filter_data_4_21 : OUT std_logic ;
      ordered_filter_data_4_20 : OUT std_logic ;
      ordered_filter_data_4_19 : OUT std_logic ;
      ordered_filter_data_4_18 : OUT std_logic ;
      ordered_filter_data_4_17 : OUT std_logic ;
      ordered_filter_data_4_16 : OUT std_logic ;
      ordered_filter_data_4_15 : OUT std_logic ;
      ordered_filter_data_4_14 : OUT std_logic ;
      ordered_filter_data_4_13 : OUT std_logic ;
      ordered_filter_data_4_12 : OUT std_logic ;
      ordered_filter_data_4_11 : OUT std_logic ;
      ordered_filter_data_4_10 : OUT std_logic ;
      ordered_filter_data_4_9 : OUT std_logic ;
      ordered_filter_data_4_8 : OUT std_logic ;
      ordered_filter_data_4_7 : OUT std_logic ;
      ordered_filter_data_4_6 : OUT std_logic ;
      ordered_filter_data_4_5 : OUT std_logic ;
      ordered_filter_data_4_4 : OUT std_logic ;
      ordered_filter_data_4_3 : OUT std_logic ;
      ordered_filter_data_4_2 : OUT std_logic ;
      ordered_filter_data_4_1 : OUT std_logic ;
      ordered_filter_data_4_0 : OUT std_logic ;
      ordered_filter_data_5_31 : OUT std_logic ;
      ordered_filter_data_5_30 : OUT std_logic ;
      ordered_filter_data_5_29 : OUT std_logic ;
      ordered_filter_data_5_28 : OUT std_logic ;
      ordered_filter_data_5_27 : OUT std_logic ;
      ordered_filter_data_5_26 : OUT std_logic ;
      ordered_filter_data_5_25 : OUT std_logic ;
      ordered_filter_data_5_24 : OUT std_logic ;
      ordered_filter_data_5_23 : OUT std_logic ;
      ordered_filter_data_5_22 : OUT std_logic ;
      ordered_filter_data_5_21 : OUT std_logic ;
      ordered_filter_data_5_20 : OUT std_logic ;
      ordered_filter_data_5_19 : OUT std_logic ;
      ordered_filter_data_5_18 : OUT std_logic ;
      ordered_filter_data_5_17 : OUT std_logic ;
      ordered_filter_data_5_16 : OUT std_logic ;
      ordered_filter_data_5_15 : OUT std_logic ;
      ordered_filter_data_5_14 : OUT std_logic ;
      ordered_filter_data_5_13 : OUT std_logic ;
      ordered_filter_data_5_12 : OUT std_logic ;
      ordered_filter_data_5_11 : OUT std_logic ;
      ordered_filter_data_5_10 : OUT std_logic ;
      ordered_filter_data_5_9 : OUT std_logic ;
      ordered_filter_data_5_8 : OUT std_logic ;
      ordered_filter_data_5_7 : OUT std_logic ;
      ordered_filter_data_5_6 : OUT std_logic ;
      ordered_filter_data_5_5 : OUT std_logic ;
      ordered_filter_data_5_4 : OUT std_logic ;
      ordered_filter_data_5_3 : OUT std_logic ;
      ordered_filter_data_5_2 : OUT std_logic ;
      ordered_filter_data_5_1 : OUT std_logic ;
      ordered_filter_data_5_0 : OUT std_logic ;
      ordered_filter_data_6_31 : OUT std_logic ;
      ordered_filter_data_6_30 : OUT std_logic ;
      ordered_filter_data_6_29 : OUT std_logic ;
      ordered_filter_data_6_28 : OUT std_logic ;
      ordered_filter_data_6_27 : OUT std_logic ;
      ordered_filter_data_6_26 : OUT std_logic ;
      ordered_filter_data_6_25 : OUT std_logic ;
      ordered_filter_data_6_24 : OUT std_logic ;
      ordered_filter_data_6_23 : OUT std_logic ;
      ordered_filter_data_6_22 : OUT std_logic ;
      ordered_filter_data_6_21 : OUT std_logic ;
      ordered_filter_data_6_20 : OUT std_logic ;
      ordered_filter_data_6_19 : OUT std_logic ;
      ordered_filter_data_6_18 : OUT std_logic ;
      ordered_filter_data_6_17 : OUT std_logic ;
      ordered_filter_data_6_16 : OUT std_logic ;
      ordered_filter_data_6_15 : OUT std_logic ;
      ordered_filter_data_6_14 : OUT std_logic ;
      ordered_filter_data_6_13 : OUT std_logic ;
      ordered_filter_data_6_12 : OUT std_logic ;
      ordered_filter_data_6_11 : OUT std_logic ;
      ordered_filter_data_6_10 : OUT std_logic ;
      ordered_filter_data_6_9 : OUT std_logic ;
      ordered_filter_data_6_8 : OUT std_logic ;
      ordered_filter_data_6_7 : OUT std_logic ;
      ordered_filter_data_6_6 : OUT std_logic ;
      ordered_filter_data_6_5 : OUT std_logic ;
      ordered_filter_data_6_4 : OUT std_logic ;
      ordered_filter_data_6_3 : OUT std_logic ;
      ordered_filter_data_6_2 : OUT std_logic ;
      ordered_filter_data_6_1 : OUT std_logic ;
      ordered_filter_data_6_0 : OUT std_logic ;
      ordered_filter_data_7_31 : OUT std_logic ;
      ordered_filter_data_7_30 : OUT std_logic ;
      ordered_filter_data_7_29 : OUT std_logic ;
      ordered_filter_data_7_28 : OUT std_logic ;
      ordered_filter_data_7_27 : OUT std_logic ;
      ordered_filter_data_7_26 : OUT std_logic ;
      ordered_filter_data_7_25 : OUT std_logic ;
      ordered_filter_data_7_24 : OUT std_logic ;
      ordered_filter_data_7_23 : OUT std_logic ;
      ordered_filter_data_7_22 : OUT std_logic ;
      ordered_filter_data_7_21 : OUT std_logic ;
      ordered_filter_data_7_20 : OUT std_logic ;
      ordered_filter_data_7_19 : OUT std_logic ;
      ordered_filter_data_7_18 : OUT std_logic ;
      ordered_filter_data_7_17 : OUT std_logic ;
      ordered_filter_data_7_16 : OUT std_logic ;
      ordered_filter_data_7_15 : OUT std_logic ;
      ordered_filter_data_7_14 : OUT std_logic ;
      ordered_filter_data_7_13 : OUT std_logic ;
      ordered_filter_data_7_12 : OUT std_logic ;
      ordered_filter_data_7_11 : OUT std_logic ;
      ordered_filter_data_7_10 : OUT std_logic ;
      ordered_filter_data_7_9 : OUT std_logic ;
      ordered_filter_data_7_8 : OUT std_logic ;
      ordered_filter_data_7_7 : OUT std_logic ;
      ordered_filter_data_7_6 : OUT std_logic ;
      ordered_filter_data_7_5 : OUT std_logic ;
      ordered_filter_data_7_4 : OUT std_logic ;
      ordered_filter_data_7_3 : OUT std_logic ;
      ordered_filter_data_7_2 : OUT std_logic ;
      ordered_filter_data_7_1 : OUT std_logic ;
      ordered_filter_data_7_0 : OUT std_logic ;
      ordered_filter_data_8_31 : OUT std_logic ;
      ordered_filter_data_8_30 : OUT std_logic ;
      ordered_filter_data_8_29 : OUT std_logic ;
      ordered_filter_data_8_28 : OUT std_logic ;
      ordered_filter_data_8_27 : OUT std_logic ;
      ordered_filter_data_8_26 : OUT std_logic ;
      ordered_filter_data_8_25 : OUT std_logic ;
      ordered_filter_data_8_24 : OUT std_logic ;
      ordered_filter_data_8_23 : OUT std_logic ;
      ordered_filter_data_8_22 : OUT std_logic ;
      ordered_filter_data_8_21 : OUT std_logic ;
      ordered_filter_data_8_20 : OUT std_logic ;
      ordered_filter_data_8_19 : OUT std_logic ;
      ordered_filter_data_8_18 : OUT std_logic ;
      ordered_filter_data_8_17 : OUT std_logic ;
      ordered_filter_data_8_16 : OUT std_logic ;
      ordered_filter_data_8_15 : OUT std_logic ;
      ordered_filter_data_8_14 : OUT std_logic ;
      ordered_filter_data_8_13 : OUT std_logic ;
      ordered_filter_data_8_12 : OUT std_logic ;
      ordered_filter_data_8_11 : OUT std_logic ;
      ordered_filter_data_8_10 : OUT std_logic ;
      ordered_filter_data_8_9 : OUT std_logic ;
      ordered_filter_data_8_8 : OUT std_logic ;
      ordered_filter_data_8_7 : OUT std_logic ;
      ordered_filter_data_8_6 : OUT std_logic ;
      ordered_filter_data_8_5 : OUT std_logic ;
      ordered_filter_data_8_4 : OUT std_logic ;
      ordered_filter_data_8_3 : OUT std_logic ;
      ordered_filter_data_8_2 : OUT std_logic ;
      ordered_filter_data_8_1 : OUT std_logic ;
      ordered_filter_data_8_0 : OUT std_logic ;
      ordered_filter_data_9_31 : OUT std_logic ;
      ordered_filter_data_9_30 : OUT std_logic ;
      ordered_filter_data_9_29 : OUT std_logic ;
      ordered_filter_data_9_28 : OUT std_logic ;
      ordered_filter_data_9_27 : OUT std_logic ;
      ordered_filter_data_9_26 : OUT std_logic ;
      ordered_filter_data_9_25 : OUT std_logic ;
      ordered_filter_data_9_24 : OUT std_logic ;
      ordered_filter_data_9_23 : OUT std_logic ;
      ordered_filter_data_9_22 : OUT std_logic ;
      ordered_filter_data_9_21 : OUT std_logic ;
      ordered_filter_data_9_20 : OUT std_logic ;
      ordered_filter_data_9_19 : OUT std_logic ;
      ordered_filter_data_9_18 : OUT std_logic ;
      ordered_filter_data_9_17 : OUT std_logic ;
      ordered_filter_data_9_16 : OUT std_logic ;
      ordered_filter_data_9_15 : OUT std_logic ;
      ordered_filter_data_9_14 : OUT std_logic ;
      ordered_filter_data_9_13 : OUT std_logic ;
      ordered_filter_data_9_12 : OUT std_logic ;
      ordered_filter_data_9_11 : OUT std_logic ;
      ordered_filter_data_9_10 : OUT std_logic ;
      ordered_filter_data_9_9 : OUT std_logic ;
      ordered_filter_data_9_8 : OUT std_logic ;
      ordered_filter_data_9_7 : OUT std_logic ;
      ordered_filter_data_9_6 : OUT std_logic ;
      ordered_filter_data_9_5 : OUT std_logic ;
      ordered_filter_data_9_4 : OUT std_logic ;
      ordered_filter_data_9_3 : OUT std_logic ;
      ordered_filter_data_9_2 : OUT std_logic ;
      ordered_filter_data_9_1 : OUT std_logic ;
      ordered_filter_data_9_0 : OUT std_logic ;
      ordered_filter_data_10_31 : OUT std_logic ;
      ordered_filter_data_10_30 : OUT std_logic ;
      ordered_filter_data_10_29 : OUT std_logic ;
      ordered_filter_data_10_28 : OUT std_logic ;
      ordered_filter_data_10_27 : OUT std_logic ;
      ordered_filter_data_10_26 : OUT std_logic ;
      ordered_filter_data_10_25 : OUT std_logic ;
      ordered_filter_data_10_24 : OUT std_logic ;
      ordered_filter_data_10_23 : OUT std_logic ;
      ordered_filter_data_10_22 : OUT std_logic ;
      ordered_filter_data_10_21 : OUT std_logic ;
      ordered_filter_data_10_20 : OUT std_logic ;
      ordered_filter_data_10_19 : OUT std_logic ;
      ordered_filter_data_10_18 : OUT std_logic ;
      ordered_filter_data_10_17 : OUT std_logic ;
      ordered_filter_data_10_16 : OUT std_logic ;
      ordered_filter_data_10_15 : OUT std_logic ;
      ordered_filter_data_10_14 : OUT std_logic ;
      ordered_filter_data_10_13 : OUT std_logic ;
      ordered_filter_data_10_12 : OUT std_logic ;
      ordered_filter_data_10_11 : OUT std_logic ;
      ordered_filter_data_10_10 : OUT std_logic ;
      ordered_filter_data_10_9 : OUT std_logic ;
      ordered_filter_data_10_8 : OUT std_logic ;
      ordered_filter_data_10_7 : OUT std_logic ;
      ordered_filter_data_10_6 : OUT std_logic ;
      ordered_filter_data_10_5 : OUT std_logic ;
      ordered_filter_data_10_4 : OUT std_logic ;
      ordered_filter_data_10_3 : OUT std_logic ;
      ordered_filter_data_10_2 : OUT std_logic ;
      ordered_filter_data_10_1 : OUT std_logic ;
      ordered_filter_data_10_0 : OUT std_logic ;
      ordered_filter_data_11_31 : OUT std_logic ;
      ordered_filter_data_11_30 : OUT std_logic ;
      ordered_filter_data_11_29 : OUT std_logic ;
      ordered_filter_data_11_28 : OUT std_logic ;
      ordered_filter_data_11_27 : OUT std_logic ;
      ordered_filter_data_11_26 : OUT std_logic ;
      ordered_filter_data_11_25 : OUT std_logic ;
      ordered_filter_data_11_24 : OUT std_logic ;
      ordered_filter_data_11_23 : OUT std_logic ;
      ordered_filter_data_11_22 : OUT std_logic ;
      ordered_filter_data_11_21 : OUT std_logic ;
      ordered_filter_data_11_20 : OUT std_logic ;
      ordered_filter_data_11_19 : OUT std_logic ;
      ordered_filter_data_11_18 : OUT std_logic ;
      ordered_filter_data_11_17 : OUT std_logic ;
      ordered_filter_data_11_16 : OUT std_logic ;
      ordered_filter_data_11_15 : OUT std_logic ;
      ordered_filter_data_11_14 : OUT std_logic ;
      ordered_filter_data_11_13 : OUT std_logic ;
      ordered_filter_data_11_12 : OUT std_logic ;
      ordered_filter_data_11_11 : OUT std_logic ;
      ordered_filter_data_11_10 : OUT std_logic ;
      ordered_filter_data_11_9 : OUT std_logic ;
      ordered_filter_data_11_8 : OUT std_logic ;
      ordered_filter_data_11_7 : OUT std_logic ;
      ordered_filter_data_11_6 : OUT std_logic ;
      ordered_filter_data_11_5 : OUT std_logic ;
      ordered_filter_data_11_4 : OUT std_logic ;
      ordered_filter_data_11_3 : OUT std_logic ;
      ordered_filter_data_11_2 : OUT std_logic ;
      ordered_filter_data_11_1 : OUT std_logic ;
      ordered_filter_data_11_0 : OUT std_logic ;
      ordered_filter_data_12_31 : OUT std_logic ;
      ordered_filter_data_12_30 : OUT std_logic ;
      ordered_filter_data_12_29 : OUT std_logic ;
      ordered_filter_data_12_28 : OUT std_logic ;
      ordered_filter_data_12_27 : OUT std_logic ;
      ordered_filter_data_12_26 : OUT std_logic ;
      ordered_filter_data_12_25 : OUT std_logic ;
      ordered_filter_data_12_24 : OUT std_logic ;
      ordered_filter_data_12_23 : OUT std_logic ;
      ordered_filter_data_12_22 : OUT std_logic ;
      ordered_filter_data_12_21 : OUT std_logic ;
      ordered_filter_data_12_20 : OUT std_logic ;
      ordered_filter_data_12_19 : OUT std_logic ;
      ordered_filter_data_12_18 : OUT std_logic ;
      ordered_filter_data_12_17 : OUT std_logic ;
      ordered_filter_data_12_16 : OUT std_logic ;
      ordered_filter_data_12_15 : OUT std_logic ;
      ordered_filter_data_12_14 : OUT std_logic ;
      ordered_filter_data_12_13 : OUT std_logic ;
      ordered_filter_data_12_12 : OUT std_logic ;
      ordered_filter_data_12_11 : OUT std_logic ;
      ordered_filter_data_12_10 : OUT std_logic ;
      ordered_filter_data_12_9 : OUT std_logic ;
      ordered_filter_data_12_8 : OUT std_logic ;
      ordered_filter_data_12_7 : OUT std_logic ;
      ordered_filter_data_12_6 : OUT std_logic ;
      ordered_filter_data_12_5 : OUT std_logic ;
      ordered_filter_data_12_4 : OUT std_logic ;
      ordered_filter_data_12_3 : OUT std_logic ;
      ordered_filter_data_12_2 : OUT std_logic ;
      ordered_filter_data_12_1 : OUT std_logic ;
      ordered_filter_data_12_0 : OUT std_logic ;
      ordered_filter_data_13_31 : OUT std_logic ;
      ordered_filter_data_13_30 : OUT std_logic ;
      ordered_filter_data_13_29 : OUT std_logic ;
      ordered_filter_data_13_28 : OUT std_logic ;
      ordered_filter_data_13_27 : OUT std_logic ;
      ordered_filter_data_13_26 : OUT std_logic ;
      ordered_filter_data_13_25 : OUT std_logic ;
      ordered_filter_data_13_24 : OUT std_logic ;
      ordered_filter_data_13_23 : OUT std_logic ;
      ordered_filter_data_13_22 : OUT std_logic ;
      ordered_filter_data_13_21 : OUT std_logic ;
      ordered_filter_data_13_20 : OUT std_logic ;
      ordered_filter_data_13_19 : OUT std_logic ;
      ordered_filter_data_13_18 : OUT std_logic ;
      ordered_filter_data_13_17 : OUT std_logic ;
      ordered_filter_data_13_16 : OUT std_logic ;
      ordered_filter_data_13_15 : OUT std_logic ;
      ordered_filter_data_13_14 : OUT std_logic ;
      ordered_filter_data_13_13 : OUT std_logic ;
      ordered_filter_data_13_12 : OUT std_logic ;
      ordered_filter_data_13_11 : OUT std_logic ;
      ordered_filter_data_13_10 : OUT std_logic ;
      ordered_filter_data_13_9 : OUT std_logic ;
      ordered_filter_data_13_8 : OUT std_logic ;
      ordered_filter_data_13_7 : OUT std_logic ;
      ordered_filter_data_13_6 : OUT std_logic ;
      ordered_filter_data_13_5 : OUT std_logic ;
      ordered_filter_data_13_4 : OUT std_logic ;
      ordered_filter_data_13_3 : OUT std_logic ;
      ordered_filter_data_13_2 : OUT std_logic ;
      ordered_filter_data_13_1 : OUT std_logic ;
      ordered_filter_data_13_0 : OUT std_logic ;
      ordered_filter_data_14_31 : OUT std_logic ;
      ordered_filter_data_14_30 : OUT std_logic ;
      ordered_filter_data_14_29 : OUT std_logic ;
      ordered_filter_data_14_28 : OUT std_logic ;
      ordered_filter_data_14_27 : OUT std_logic ;
      ordered_filter_data_14_26 : OUT std_logic ;
      ordered_filter_data_14_25 : OUT std_logic ;
      ordered_filter_data_14_24 : OUT std_logic ;
      ordered_filter_data_14_23 : OUT std_logic ;
      ordered_filter_data_14_22 : OUT std_logic ;
      ordered_filter_data_14_21 : OUT std_logic ;
      ordered_filter_data_14_20 : OUT std_logic ;
      ordered_filter_data_14_19 : OUT std_logic ;
      ordered_filter_data_14_18 : OUT std_logic ;
      ordered_filter_data_14_17 : OUT std_logic ;
      ordered_filter_data_14_16 : OUT std_logic ;
      ordered_filter_data_14_15 : OUT std_logic ;
      ordered_filter_data_14_14 : OUT std_logic ;
      ordered_filter_data_14_13 : OUT std_logic ;
      ordered_filter_data_14_12 : OUT std_logic ;
      ordered_filter_data_14_11 : OUT std_logic ;
      ordered_filter_data_14_10 : OUT std_logic ;
      ordered_filter_data_14_9 : OUT std_logic ;
      ordered_filter_data_14_8 : OUT std_logic ;
      ordered_filter_data_14_7 : OUT std_logic ;
      ordered_filter_data_14_6 : OUT std_logic ;
      ordered_filter_data_14_5 : OUT std_logic ;
      ordered_filter_data_14_4 : OUT std_logic ;
      ordered_filter_data_14_3 : OUT std_logic ;
      ordered_filter_data_14_2 : OUT std_logic ;
      ordered_filter_data_14_1 : OUT std_logic ;
      ordered_filter_data_14_0 : OUT std_logic ;
      ordered_filter_data_15_31 : OUT std_logic ;
      ordered_filter_data_15_30 : OUT std_logic ;
      ordered_filter_data_15_29 : OUT std_logic ;
      ordered_filter_data_15_28 : OUT std_logic ;
      ordered_filter_data_15_27 : OUT std_logic ;
      ordered_filter_data_15_26 : OUT std_logic ;
      ordered_filter_data_15_25 : OUT std_logic ;
      ordered_filter_data_15_24 : OUT std_logic ;
      ordered_filter_data_15_23 : OUT std_logic ;
      ordered_filter_data_15_22 : OUT std_logic ;
      ordered_filter_data_15_21 : OUT std_logic ;
      ordered_filter_data_15_20 : OUT std_logic ;
      ordered_filter_data_15_19 : OUT std_logic ;
      ordered_filter_data_15_18 : OUT std_logic ;
      ordered_filter_data_15_17 : OUT std_logic ;
      ordered_filter_data_15_16 : OUT std_logic ;
      ordered_filter_data_15_15 : OUT std_logic ;
      ordered_filter_data_15_14 : OUT std_logic ;
      ordered_filter_data_15_13 : OUT std_logic ;
      ordered_filter_data_15_12 : OUT std_logic ;
      ordered_filter_data_15_11 : OUT std_logic ;
      ordered_filter_data_15_10 : OUT std_logic ;
      ordered_filter_data_15_9 : OUT std_logic ;
      ordered_filter_data_15_8 : OUT std_logic ;
      ordered_filter_data_15_7 : OUT std_logic ;
      ordered_filter_data_15_6 : OUT std_logic ;
      ordered_filter_data_15_5 : OUT std_logic ;
      ordered_filter_data_15_4 : OUT std_logic ;
      ordered_filter_data_15_3 : OUT std_logic ;
      ordered_filter_data_15_2 : OUT std_logic ;
      ordered_filter_data_15_1 : OUT std_logic ;
      ordered_filter_data_15_0 : OUT std_logic ;
      ordered_filter_data_16_31 : OUT std_logic ;
      ordered_filter_data_16_30 : OUT std_logic ;
      ordered_filter_data_16_29 : OUT std_logic ;
      ordered_filter_data_16_28 : OUT std_logic ;
      ordered_filter_data_16_27 : OUT std_logic ;
      ordered_filter_data_16_26 : OUT std_logic ;
      ordered_filter_data_16_25 : OUT std_logic ;
      ordered_filter_data_16_24 : OUT std_logic ;
      ordered_filter_data_16_23 : OUT std_logic ;
      ordered_filter_data_16_22 : OUT std_logic ;
      ordered_filter_data_16_21 : OUT std_logic ;
      ordered_filter_data_16_20 : OUT std_logic ;
      ordered_filter_data_16_19 : OUT std_logic ;
      ordered_filter_data_16_18 : OUT std_logic ;
      ordered_filter_data_16_17 : OUT std_logic ;
      ordered_filter_data_16_16 : OUT std_logic ;
      ordered_filter_data_16_15 : OUT std_logic ;
      ordered_filter_data_16_14 : OUT std_logic ;
      ordered_filter_data_16_13 : OUT std_logic ;
      ordered_filter_data_16_12 : OUT std_logic ;
      ordered_filter_data_16_11 : OUT std_logic ;
      ordered_filter_data_16_10 : OUT std_logic ;
      ordered_filter_data_16_9 : OUT std_logic ;
      ordered_filter_data_16_8 : OUT std_logic ;
      ordered_filter_data_16_7 : OUT std_logic ;
      ordered_filter_data_16_6 : OUT std_logic ;
      ordered_filter_data_16_5 : OUT std_logic ;
      ordered_filter_data_16_4 : OUT std_logic ;
      ordered_filter_data_16_3 : OUT std_logic ;
      ordered_filter_data_16_2 : OUT std_logic ;
      ordered_filter_data_16_1 : OUT std_logic ;
      ordered_filter_data_16_0 : OUT std_logic ;
      ordered_filter_data_17_31 : OUT std_logic ;
      ordered_filter_data_17_30 : OUT std_logic ;
      ordered_filter_data_17_29 : OUT std_logic ;
      ordered_filter_data_17_28 : OUT std_logic ;
      ordered_filter_data_17_27 : OUT std_logic ;
      ordered_filter_data_17_26 : OUT std_logic ;
      ordered_filter_data_17_25 : OUT std_logic ;
      ordered_filter_data_17_24 : OUT std_logic ;
      ordered_filter_data_17_23 : OUT std_logic ;
      ordered_filter_data_17_22 : OUT std_logic ;
      ordered_filter_data_17_21 : OUT std_logic ;
      ordered_filter_data_17_20 : OUT std_logic ;
      ordered_filter_data_17_19 : OUT std_logic ;
      ordered_filter_data_17_18 : OUT std_logic ;
      ordered_filter_data_17_17 : OUT std_logic ;
      ordered_filter_data_17_16 : OUT std_logic ;
      ordered_filter_data_17_15 : OUT std_logic ;
      ordered_filter_data_17_14 : OUT std_logic ;
      ordered_filter_data_17_13 : OUT std_logic ;
      ordered_filter_data_17_12 : OUT std_logic ;
      ordered_filter_data_17_11 : OUT std_logic ;
      ordered_filter_data_17_10 : OUT std_logic ;
      ordered_filter_data_17_9 : OUT std_logic ;
      ordered_filter_data_17_8 : OUT std_logic ;
      ordered_filter_data_17_7 : OUT std_logic ;
      ordered_filter_data_17_6 : OUT std_logic ;
      ordered_filter_data_17_5 : OUT std_logic ;
      ordered_filter_data_17_4 : OUT std_logic ;
      ordered_filter_data_17_3 : OUT std_logic ;
      ordered_filter_data_17_2 : OUT std_logic ;
      ordered_filter_data_17_1 : OUT std_logic ;
      ordered_filter_data_17_0 : OUT std_logic ;
      ordered_filter_data_18_31 : OUT std_logic ;
      ordered_filter_data_18_30 : OUT std_logic ;
      ordered_filter_data_18_29 : OUT std_logic ;
      ordered_filter_data_18_28 : OUT std_logic ;
      ordered_filter_data_18_27 : OUT std_logic ;
      ordered_filter_data_18_26 : OUT std_logic ;
      ordered_filter_data_18_25 : OUT std_logic ;
      ordered_filter_data_18_24 : OUT std_logic ;
      ordered_filter_data_18_23 : OUT std_logic ;
      ordered_filter_data_18_22 : OUT std_logic ;
      ordered_filter_data_18_21 : OUT std_logic ;
      ordered_filter_data_18_20 : OUT std_logic ;
      ordered_filter_data_18_19 : OUT std_logic ;
      ordered_filter_data_18_18 : OUT std_logic ;
      ordered_filter_data_18_17 : OUT std_logic ;
      ordered_filter_data_18_16 : OUT std_logic ;
      ordered_filter_data_18_15 : OUT std_logic ;
      ordered_filter_data_18_14 : OUT std_logic ;
      ordered_filter_data_18_13 : OUT std_logic ;
      ordered_filter_data_18_12 : OUT std_logic ;
      ordered_filter_data_18_11 : OUT std_logic ;
      ordered_filter_data_18_10 : OUT std_logic ;
      ordered_filter_data_18_9 : OUT std_logic ;
      ordered_filter_data_18_8 : OUT std_logic ;
      ordered_filter_data_18_7 : OUT std_logic ;
      ordered_filter_data_18_6 : OUT std_logic ;
      ordered_filter_data_18_5 : OUT std_logic ;
      ordered_filter_data_18_4 : OUT std_logic ;
      ordered_filter_data_18_3 : OUT std_logic ;
      ordered_filter_data_18_2 : OUT std_logic ;
      ordered_filter_data_18_1 : OUT std_logic ;
      ordered_filter_data_18_0 : OUT std_logic ;
      ordered_filter_data_19_31 : OUT std_logic ;
      ordered_filter_data_19_30 : OUT std_logic ;
      ordered_filter_data_19_29 : OUT std_logic ;
      ordered_filter_data_19_28 : OUT std_logic ;
      ordered_filter_data_19_27 : OUT std_logic ;
      ordered_filter_data_19_26 : OUT std_logic ;
      ordered_filter_data_19_25 : OUT std_logic ;
      ordered_filter_data_19_24 : OUT std_logic ;
      ordered_filter_data_19_23 : OUT std_logic ;
      ordered_filter_data_19_22 : OUT std_logic ;
      ordered_filter_data_19_21 : OUT std_logic ;
      ordered_filter_data_19_20 : OUT std_logic ;
      ordered_filter_data_19_19 : OUT std_logic ;
      ordered_filter_data_19_18 : OUT std_logic ;
      ordered_filter_data_19_17 : OUT std_logic ;
      ordered_filter_data_19_16 : OUT std_logic ;
      ordered_filter_data_19_15 : OUT std_logic ;
      ordered_filter_data_19_14 : OUT std_logic ;
      ordered_filter_data_19_13 : OUT std_logic ;
      ordered_filter_data_19_12 : OUT std_logic ;
      ordered_filter_data_19_11 : OUT std_logic ;
      ordered_filter_data_19_10 : OUT std_logic ;
      ordered_filter_data_19_9 : OUT std_logic ;
      ordered_filter_data_19_8 : OUT std_logic ;
      ordered_filter_data_19_7 : OUT std_logic ;
      ordered_filter_data_19_6 : OUT std_logic ;
      ordered_filter_data_19_5 : OUT std_logic ;
      ordered_filter_data_19_4 : OUT std_logic ;
      ordered_filter_data_19_3 : OUT std_logic ;
      ordered_filter_data_19_2 : OUT std_logic ;
      ordered_filter_data_19_1 : OUT std_logic ;
      ordered_filter_data_19_0 : OUT std_logic ;
      ordered_filter_data_20_31 : OUT std_logic ;
      ordered_filter_data_20_30 : OUT std_logic ;
      ordered_filter_data_20_29 : OUT std_logic ;
      ordered_filter_data_20_28 : OUT std_logic ;
      ordered_filter_data_20_27 : OUT std_logic ;
      ordered_filter_data_20_26 : OUT std_logic ;
      ordered_filter_data_20_25 : OUT std_logic ;
      ordered_filter_data_20_24 : OUT std_logic ;
      ordered_filter_data_20_23 : OUT std_logic ;
      ordered_filter_data_20_22 : OUT std_logic ;
      ordered_filter_data_20_21 : OUT std_logic ;
      ordered_filter_data_20_20 : OUT std_logic ;
      ordered_filter_data_20_19 : OUT std_logic ;
      ordered_filter_data_20_18 : OUT std_logic ;
      ordered_filter_data_20_17 : OUT std_logic ;
      ordered_filter_data_20_16 : OUT std_logic ;
      ordered_filter_data_20_15 : OUT std_logic ;
      ordered_filter_data_20_14 : OUT std_logic ;
      ordered_filter_data_20_13 : OUT std_logic ;
      ordered_filter_data_20_12 : OUT std_logic ;
      ordered_filter_data_20_11 : OUT std_logic ;
      ordered_filter_data_20_10 : OUT std_logic ;
      ordered_filter_data_20_9 : OUT std_logic ;
      ordered_filter_data_20_8 : OUT std_logic ;
      ordered_filter_data_20_7 : OUT std_logic ;
      ordered_filter_data_20_6 : OUT std_logic ;
      ordered_filter_data_20_5 : OUT std_logic ;
      ordered_filter_data_20_4 : OUT std_logic ;
      ordered_filter_data_20_3 : OUT std_logic ;
      ordered_filter_data_20_2 : OUT std_logic ;
      ordered_filter_data_20_1 : OUT std_logic ;
      ordered_filter_data_20_0 : OUT std_logic ;
      ordered_filter_data_21_31 : OUT std_logic ;
      ordered_filter_data_21_30 : OUT std_logic ;
      ordered_filter_data_21_29 : OUT std_logic ;
      ordered_filter_data_21_28 : OUT std_logic ;
      ordered_filter_data_21_27 : OUT std_logic ;
      ordered_filter_data_21_26 : OUT std_logic ;
      ordered_filter_data_21_25 : OUT std_logic ;
      ordered_filter_data_21_24 : OUT std_logic ;
      ordered_filter_data_21_23 : OUT std_logic ;
      ordered_filter_data_21_22 : OUT std_logic ;
      ordered_filter_data_21_21 : OUT std_logic ;
      ordered_filter_data_21_20 : OUT std_logic ;
      ordered_filter_data_21_19 : OUT std_logic ;
      ordered_filter_data_21_18 : OUT std_logic ;
      ordered_filter_data_21_17 : OUT std_logic ;
      ordered_filter_data_21_16 : OUT std_logic ;
      ordered_filter_data_21_15 : OUT std_logic ;
      ordered_filter_data_21_14 : OUT std_logic ;
      ordered_filter_data_21_13 : OUT std_logic ;
      ordered_filter_data_21_12 : OUT std_logic ;
      ordered_filter_data_21_11 : OUT std_logic ;
      ordered_filter_data_21_10 : OUT std_logic ;
      ordered_filter_data_21_9 : OUT std_logic ;
      ordered_filter_data_21_8 : OUT std_logic ;
      ordered_filter_data_21_7 : OUT std_logic ;
      ordered_filter_data_21_6 : OUT std_logic ;
      ordered_filter_data_21_5 : OUT std_logic ;
      ordered_filter_data_21_4 : OUT std_logic ;
      ordered_filter_data_21_3 : OUT std_logic ;
      ordered_filter_data_21_2 : OUT std_logic ;
      ordered_filter_data_21_1 : OUT std_logic ;
      ordered_filter_data_21_0 : OUT std_logic ;
      ordered_filter_data_22_31 : OUT std_logic ;
      ordered_filter_data_22_30 : OUT std_logic ;
      ordered_filter_data_22_29 : OUT std_logic ;
      ordered_filter_data_22_28 : OUT std_logic ;
      ordered_filter_data_22_27 : OUT std_logic ;
      ordered_filter_data_22_26 : OUT std_logic ;
      ordered_filter_data_22_25 : OUT std_logic ;
      ordered_filter_data_22_24 : OUT std_logic ;
      ordered_filter_data_22_23 : OUT std_logic ;
      ordered_filter_data_22_22 : OUT std_logic ;
      ordered_filter_data_22_21 : OUT std_logic ;
      ordered_filter_data_22_20 : OUT std_logic ;
      ordered_filter_data_22_19 : OUT std_logic ;
      ordered_filter_data_22_18 : OUT std_logic ;
      ordered_filter_data_22_17 : OUT std_logic ;
      ordered_filter_data_22_16 : OUT std_logic ;
      ordered_filter_data_22_15 : OUT std_logic ;
      ordered_filter_data_22_14 : OUT std_logic ;
      ordered_filter_data_22_13 : OUT std_logic ;
      ordered_filter_data_22_12 : OUT std_logic ;
      ordered_filter_data_22_11 : OUT std_logic ;
      ordered_filter_data_22_10 : OUT std_logic ;
      ordered_filter_data_22_9 : OUT std_logic ;
      ordered_filter_data_22_8 : OUT std_logic ;
      ordered_filter_data_22_7 : OUT std_logic ;
      ordered_filter_data_22_6 : OUT std_logic ;
      ordered_filter_data_22_5 : OUT std_logic ;
      ordered_filter_data_22_4 : OUT std_logic ;
      ordered_filter_data_22_3 : OUT std_logic ;
      ordered_filter_data_22_2 : OUT std_logic ;
      ordered_filter_data_22_1 : OUT std_logic ;
      ordered_filter_data_22_0 : OUT std_logic ;
      ordered_filter_data_23_31 : OUT std_logic ;
      ordered_filter_data_23_30 : OUT std_logic ;
      ordered_filter_data_23_29 : OUT std_logic ;
      ordered_filter_data_23_28 : OUT std_logic ;
      ordered_filter_data_23_27 : OUT std_logic ;
      ordered_filter_data_23_26 : OUT std_logic ;
      ordered_filter_data_23_25 : OUT std_logic ;
      ordered_filter_data_23_24 : OUT std_logic ;
      ordered_filter_data_23_23 : OUT std_logic ;
      ordered_filter_data_23_22 : OUT std_logic ;
      ordered_filter_data_23_21 : OUT std_logic ;
      ordered_filter_data_23_20 : OUT std_logic ;
      ordered_filter_data_23_19 : OUT std_logic ;
      ordered_filter_data_23_18 : OUT std_logic ;
      ordered_filter_data_23_17 : OUT std_logic ;
      ordered_filter_data_23_16 : OUT std_logic ;
      ordered_filter_data_23_15 : OUT std_logic ;
      ordered_filter_data_23_14 : OUT std_logic ;
      ordered_filter_data_23_13 : OUT std_logic ;
      ordered_filter_data_23_12 : OUT std_logic ;
      ordered_filter_data_23_11 : OUT std_logic ;
      ordered_filter_data_23_10 : OUT std_logic ;
      ordered_filter_data_23_9 : OUT std_logic ;
      ordered_filter_data_23_8 : OUT std_logic ;
      ordered_filter_data_23_7 : OUT std_logic ;
      ordered_filter_data_23_6 : OUT std_logic ;
      ordered_filter_data_23_5 : OUT std_logic ;
      ordered_filter_data_23_4 : OUT std_logic ;
      ordered_filter_data_23_3 : OUT std_logic ;
      ordered_filter_data_23_2 : OUT std_logic ;
      ordered_filter_data_23_1 : OUT std_logic ;
      ordered_filter_data_23_0 : OUT std_logic ;
      ordered_filter_data_24_31 : OUT std_logic ;
      ordered_filter_data_24_30 : OUT std_logic ;
      ordered_filter_data_24_29 : OUT std_logic ;
      ordered_filter_data_24_28 : OUT std_logic ;
      ordered_filter_data_24_27 : OUT std_logic ;
      ordered_filter_data_24_26 : OUT std_logic ;
      ordered_filter_data_24_25 : OUT std_logic ;
      ordered_filter_data_24_24 : OUT std_logic ;
      ordered_filter_data_24_23 : OUT std_logic ;
      ordered_filter_data_24_22 : OUT std_logic ;
      ordered_filter_data_24_21 : OUT std_logic ;
      ordered_filter_data_24_20 : OUT std_logic ;
      ordered_filter_data_24_19 : OUT std_logic ;
      ordered_filter_data_24_18 : OUT std_logic ;
      ordered_filter_data_24_17 : OUT std_logic ;
      ordered_filter_data_24_16 : OUT std_logic ;
      ordered_filter_data_24_15 : OUT std_logic ;
      ordered_filter_data_24_14 : OUT std_logic ;
      ordered_filter_data_24_13 : OUT std_logic ;
      ordered_filter_data_24_12 : OUT std_logic ;
      ordered_filter_data_24_11 : OUT std_logic ;
      ordered_filter_data_24_10 : OUT std_logic ;
      ordered_filter_data_24_9 : OUT std_logic ;
      ordered_filter_data_24_8 : OUT std_logic ;
      ordered_filter_data_24_7 : OUT std_logic ;
      ordered_filter_data_24_6 : OUT std_logic ;
      ordered_filter_data_24_5 : OUT std_logic ;
      ordered_filter_data_24_4 : OUT std_logic ;
      ordered_filter_data_24_3 : OUT std_logic ;
      ordered_filter_data_24_2 : OUT std_logic ;
      ordered_filter_data_24_1 : OUT std_logic ;
      ordered_filter_data_24_0 : OUT std_logic) ;
end MuxLayer ;

architecture Structural_unfold_3247_0 of MuxLayer is
   signal ordered_img_data_9_15_EXMPLR, ordered_img_data_10_15_EXMPLR, 
      ordered_img_data_11_15_EXMPLR, ordered_img_data_12_15_EXMPLR, 
      ordered_img_data_13_15_EXMPLR, ordered_img_data_14_15_EXMPLR, 
      ordered_img_data_15_15_EXMPLR, ordered_img_data_16_15_EXMPLR, 
      ordered_img_data_17_15_EXMPLR, ordered_filter_data_24_0_EXMPLR, nx1206, 
      nx1209, nx1211, nx1213, nx1215, nx1217, nx1219, nx1221, nx1223, nx1225, 
      nx1227, nx1229, nx1231, nx1233, nx1235, nx1237, nx1239, nx1241, nx1243, 
      nx1245, nx1247, nx1249, nx1251, nx1253, nx1255, nx1257, nx1259, nx1261, 
      nx1263, nx1265, nx1267, nx1269, nx1271, nx1273, nx1287, nx1301, nx1315, 
      nx1319, nx1321, nx1323, nx1317, nx1317_XX0_XREP32, nx1325, nx1331, 
      nx1345, nx1346, nx1354, nx1356, nx1358, nx1361, nx1363, nx1365, nx1367, 
      nx1369, nx1371, nx1373, nx1375, nx1377, nx1379, nx1381, nx1383, nx1385, 
      nx1387, nx1389, nx1391: std_logic ;

begin
   ordered_img_data_0_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_0_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_1_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_2_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_3_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_4_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_5_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_6_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_7_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_8_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_9_31 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_30 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_29 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_28 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_27 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_26 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_25 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_24 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_23 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_22 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_21 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_20 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_19 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_18 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_17 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_16 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_9_15 <= ordered_img_data_9_15_EXMPLR ;
   ordered_img_data_10_31 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_30 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_29 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_28 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_27 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_26 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_25 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_24 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_23 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_22 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_21 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_20 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_19 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_18 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_17 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_16 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_10_15 <= ordered_img_data_10_15_EXMPLR ;
   ordered_img_data_11_31 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_30 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_29 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_28 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_27 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_26 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_25 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_24 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_23 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_22 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_21 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_20 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_19 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_18 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_17 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_16 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_11_15 <= ordered_img_data_11_15_EXMPLR ;
   ordered_img_data_12_31 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_30 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_29 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_28 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_27 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_26 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_25 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_24 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_23 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_22 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_21 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_20 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_19 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_18 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_17 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_16 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_12_15 <= ordered_img_data_12_15_EXMPLR ;
   ordered_img_data_13_31 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_30 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_29 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_28 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_27 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_26 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_25 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_24 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_23 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_22 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_21 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_20 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_19 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_18 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_17 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_16 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_13_15 <= ordered_img_data_13_15_EXMPLR ;
   ordered_img_data_14_31 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_30 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_29 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_28 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_27 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_26 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_25 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_24 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_23 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_22 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_21 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_20 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_19 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_18 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_17 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_16 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_14_15 <= ordered_img_data_14_15_EXMPLR ;
   ordered_img_data_15_31 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_30 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_29 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_28 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_27 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_26 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_25 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_24 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_23 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_22 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_21 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_20 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_19 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_18 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_17 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_16 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_15_15 <= ordered_img_data_15_15_EXMPLR ;
   ordered_img_data_16_31 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_30 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_29 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_28 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_27 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_26 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_25 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_24 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_23 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_22 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_21 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_20 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_19 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_18 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_17 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_16 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_16_15 <= ordered_img_data_16_15_EXMPLR ;
   ordered_img_data_17_31 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_30 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_29 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_28 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_27 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_26 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_25 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_24 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_23 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_22 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_21 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_20 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_19 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_18 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_17 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_16 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_17_15 <= ordered_img_data_17_15_EXMPLR ;
   ordered_img_data_18_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_18_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_19_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_20_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_21_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_22_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_23_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_img_data_24_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_0_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_1_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_2_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_3_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_4_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_5_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_6_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_7_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_8_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_9_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_10_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_11_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_12_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_13_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_14_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_15_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_16_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_17_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_18_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_19_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_20_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_21_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_22_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_23_0 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_31 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_30 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_29 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_28 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_27 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_26 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_25 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_24 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_23 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_22 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_21 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_20 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_19 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_18 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_17 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_16 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_15 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_14 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_13 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_12 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_11 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_10 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_9 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_8 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_7 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_6 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_5 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_4 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_3 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_2 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_1 <= ordered_filter_data_24_0_EXMPLR ;
   ordered_filter_data_24_0 <= ordered_filter_data_24_0_EXMPLR ;
   ix46 : fake_gnd port map ( Y=>ordered_filter_data_24_0_EXMPLR);
   ix7 : mux21_ni port map ( Y=>ordered_filter_data_17_0, A0=>
      filter_data_17_0, A1=>filter_data_8_0, S0=>nx1206);
   ix15 : mux21_ni port map ( Y=>ordered_filter_data_17_1, A0=>
      filter_data_17_1, A1=>filter_data_8_1, S0=>nx1206);
   ix23 : mux21_ni port map ( Y=>ordered_filter_data_17_2, A0=>
      filter_data_17_2, A1=>filter_data_8_2, S0=>nx1206);
   ix31 : mux21_ni port map ( Y=>ordered_filter_data_17_3, A0=>
      filter_data_17_3, A1=>filter_data_8_3, S0=>nx1206);
   ix39 : mux21_ni port map ( Y=>ordered_filter_data_17_4, A0=>
      filter_data_17_4, A1=>filter_data_8_4, S0=>nx1206);
   ix47 : mux21_ni port map ( Y=>ordered_filter_data_17_5, A0=>
      filter_data_17_5, A1=>filter_data_8_5, S0=>nx1206);
   ix55 : mux21_ni port map ( Y=>ordered_filter_data_17_6, A0=>
      filter_data_17_6, A1=>filter_data_8_6, S0=>nx1206);
   ix63 : mux21_ni port map ( Y=>ordered_filter_data_17_7, A0=>
      filter_data_17_7, A1=>filter_data_8_7, S0=>nx1209);
   ix71 : mux21_ni port map ( Y=>ordered_filter_data_17_8, A0=>
      filter_data_17_8, A1=>filter_data_8_8, S0=>nx1209);
   ix79 : mux21_ni port map ( Y=>ordered_filter_data_17_9, A0=>
      filter_data_17_9, A1=>filter_data_8_9, S0=>nx1209);
   ix87 : mux21_ni port map ( Y=>ordered_filter_data_17_10, A0=>
      filter_data_17_10, A1=>filter_data_8_10, S0=>nx1209);
   ix95 : mux21_ni port map ( Y=>ordered_filter_data_17_11, A0=>
      filter_data_17_11, A1=>filter_data_8_11, S0=>nx1209);
   ix103 : mux21_ni port map ( Y=>ordered_filter_data_17_12, A0=>
      filter_data_17_12, A1=>filter_data_8_12, S0=>nx1209);
   ix111 : mux21_ni port map ( Y=>ordered_filter_data_17_13, A0=>
      filter_data_17_13, A1=>filter_data_8_13, S0=>nx1209);
   ix119 : mux21_ni port map ( Y=>ordered_filter_data_17_14, A0=>
      filter_data_17_14, A1=>filter_data_8_14, S0=>nx1211);
   ix127 : mux21_ni port map ( Y=>ordered_filter_data_17_15, A0=>
      filter_data_17_31, A1=>filter_data_8_31, S0=>nx1211);
   ix391 : mux21_ni port map ( Y=>ordered_filter_data_16_0, A0=>
      filter_data_16_0, A1=>filter_data_7_0, S0=>nx1211);
   ix399 : mux21_ni port map ( Y=>ordered_filter_data_16_1, A0=>
      filter_data_16_1, A1=>filter_data_7_1, S0=>nx1211);
   ix407 : mux21_ni port map ( Y=>ordered_filter_data_16_2, A0=>
      filter_data_16_2, A1=>filter_data_7_2, S0=>nx1211);
   ix415 : mux21_ni port map ( Y=>ordered_filter_data_16_3, A0=>
      filter_data_16_3, A1=>filter_data_7_3, S0=>nx1211);
   ix423 : mux21_ni port map ( Y=>ordered_filter_data_16_4, A0=>
      filter_data_16_4, A1=>filter_data_7_4, S0=>nx1211);
   ix431 : mux21_ni port map ( Y=>ordered_filter_data_16_5, A0=>
      filter_data_16_5, A1=>filter_data_7_5, S0=>nx1213);
   ix439 : mux21_ni port map ( Y=>ordered_filter_data_16_6, A0=>
      filter_data_16_6, A1=>filter_data_7_6, S0=>nx1213);
   ix447 : mux21_ni port map ( Y=>ordered_filter_data_16_7, A0=>
      filter_data_16_7, A1=>filter_data_7_7, S0=>nx1213);
   ix455 : mux21_ni port map ( Y=>ordered_filter_data_16_8, A0=>
      filter_data_16_8, A1=>filter_data_7_8, S0=>nx1213);
   ix463 : mux21_ni port map ( Y=>ordered_filter_data_16_9, A0=>
      filter_data_16_9, A1=>filter_data_7_9, S0=>nx1213);
   ix471 : mux21_ni port map ( Y=>ordered_filter_data_16_10, A0=>
      filter_data_16_10, A1=>filter_data_7_10, S0=>nx1213);
   ix479 : mux21_ni port map ( Y=>ordered_filter_data_16_11, A0=>
      filter_data_16_11, A1=>filter_data_7_11, S0=>nx1213);
   ix487 : mux21_ni port map ( Y=>ordered_filter_data_16_12, A0=>
      filter_data_16_12, A1=>filter_data_7_12, S0=>nx1215);
   ix495 : mux21_ni port map ( Y=>ordered_filter_data_16_13, A0=>
      filter_data_16_13, A1=>filter_data_7_13, S0=>nx1215);
   ix503 : mux21_ni port map ( Y=>ordered_filter_data_16_14, A0=>
      filter_data_16_14, A1=>filter_data_7_14, S0=>nx1215);
   ix511 : mux21_ni port map ( Y=>ordered_filter_data_16_15, A0=>
      filter_data_16_31, A1=>filter_data_7_31, S0=>nx1215);
   ix775 : mux21_ni port map ( Y=>ordered_filter_data_15_0, A0=>
      filter_data_15_0, A1=>filter_data_6_0, S0=>nx1215);
   ix783 : mux21_ni port map ( Y=>ordered_filter_data_15_1, A0=>
      filter_data_15_1, A1=>filter_data_6_1, S0=>nx1215);
   ix791 : mux21_ni port map ( Y=>ordered_filter_data_15_2, A0=>
      filter_data_15_2, A1=>filter_data_6_2, S0=>nx1215);
   ix799 : mux21_ni port map ( Y=>ordered_filter_data_15_3, A0=>
      filter_data_15_3, A1=>filter_data_6_3, S0=>nx1217);
   ix807 : mux21_ni port map ( Y=>ordered_filter_data_15_4, A0=>
      filter_data_15_4, A1=>filter_data_6_4, S0=>nx1217);
   ix815 : mux21_ni port map ( Y=>ordered_filter_data_15_5, A0=>
      filter_data_15_5, A1=>filter_data_6_5, S0=>nx1217);
   ix823 : mux21_ni port map ( Y=>ordered_filter_data_15_6, A0=>
      filter_data_15_6, A1=>filter_data_6_6, S0=>nx1217);
   ix831 : mux21_ni port map ( Y=>ordered_filter_data_15_7, A0=>
      filter_data_15_7, A1=>filter_data_6_7, S0=>nx1217);
   ix839 : mux21_ni port map ( Y=>ordered_filter_data_15_8, A0=>
      filter_data_15_8, A1=>filter_data_6_8, S0=>nx1217);
   ix847 : mux21_ni port map ( Y=>ordered_filter_data_15_9, A0=>
      filter_data_15_9, A1=>filter_data_6_9, S0=>nx1217);
   ix855 : mux21_ni port map ( Y=>ordered_filter_data_15_10, A0=>
      filter_data_15_10, A1=>filter_data_6_10, S0=>nx1219);
   ix863 : mux21_ni port map ( Y=>ordered_filter_data_15_11, A0=>
      filter_data_15_11, A1=>filter_data_6_11, S0=>nx1219);
   ix871 : mux21_ni port map ( Y=>ordered_filter_data_15_12, A0=>
      filter_data_15_12, A1=>filter_data_6_12, S0=>nx1219);
   ix879 : mux21_ni port map ( Y=>ordered_filter_data_15_13, A0=>
      filter_data_15_13, A1=>filter_data_6_13, S0=>nx1219);
   ix887 : mux21_ni port map ( Y=>ordered_filter_data_15_14, A0=>
      filter_data_15_14, A1=>filter_data_6_14, S0=>nx1219);
   ix895 : mux21_ni port map ( Y=>ordered_filter_data_15_15, A0=>
      filter_data_15_31, A1=>filter_data_6_31, S0=>nx1219);
   ix1159 : mux21_ni port map ( Y=>ordered_filter_data_14_0, A0=>
      filter_data_14_0, A1=>filter_data_5_0, S0=>nx1219);
   ix1167 : mux21_ni port map ( Y=>ordered_filter_data_14_1, A0=>
      filter_data_14_1, A1=>filter_data_5_1, S0=>nx1221);
   ix1175 : mux21_ni port map ( Y=>ordered_filter_data_14_2, A0=>
      filter_data_14_2, A1=>filter_data_5_2, S0=>nx1221);
   ix1183 : mux21_ni port map ( Y=>ordered_filter_data_14_3, A0=>
      filter_data_14_3, A1=>filter_data_5_3, S0=>nx1221);
   ix1191 : mux21_ni port map ( Y=>ordered_filter_data_14_4, A0=>
      filter_data_14_4, A1=>filter_data_5_4, S0=>nx1221);
   ix1199 : mux21_ni port map ( Y=>ordered_filter_data_14_5, A0=>
      filter_data_14_5, A1=>filter_data_5_5, S0=>nx1221);
   ix1207 : mux21_ni port map ( Y=>ordered_filter_data_14_6, A0=>
      filter_data_14_6, A1=>filter_data_5_6, S0=>nx1221);
   ix1215 : mux21_ni port map ( Y=>ordered_filter_data_14_7, A0=>
      filter_data_14_7, A1=>filter_data_5_7, S0=>nx1221);
   ix1223 : mux21_ni port map ( Y=>ordered_filter_data_14_8, A0=>
      filter_data_14_8, A1=>filter_data_5_8, S0=>nx1223);
   ix1231 : mux21_ni port map ( Y=>ordered_filter_data_14_9, A0=>
      filter_data_14_9, A1=>filter_data_5_9, S0=>nx1223);
   ix1239 : mux21_ni port map ( Y=>ordered_filter_data_14_10, A0=>
      filter_data_14_10, A1=>filter_data_5_10, S0=>nx1223);
   ix1247 : mux21_ni port map ( Y=>ordered_filter_data_14_11, A0=>
      filter_data_14_11, A1=>filter_data_5_11, S0=>nx1223);
   ix1255 : mux21_ni port map ( Y=>ordered_filter_data_14_12, A0=>
      filter_data_14_12, A1=>filter_data_5_12, S0=>nx1223);
   ix1263 : mux21_ni port map ( Y=>ordered_filter_data_14_13, A0=>
      filter_data_14_13, A1=>filter_data_5_13, S0=>nx1223);
   ix1271 : mux21_ni port map ( Y=>ordered_filter_data_14_14, A0=>
      filter_data_14_14, A1=>filter_data_5_14, S0=>nx1223);
   ix1279 : mux21_ni port map ( Y=>ordered_filter_data_14_15, A0=>
      filter_data_14_31, A1=>filter_data_5_31, S0=>nx1225);
   ix1543 : mux21_ni port map ( Y=>ordered_filter_data_13_0, A0=>
      filter_data_9_0, A1=>filter_data_4_0, S0=>nx1225);
   ix1551 : mux21_ni port map ( Y=>ordered_filter_data_13_1, A0=>
      filter_data_9_1, A1=>filter_data_4_1, S0=>nx1225);
   ix1559 : mux21_ni port map ( Y=>ordered_filter_data_13_2, A0=>
      filter_data_9_2, A1=>filter_data_4_2, S0=>nx1225);
   ix1567 : mux21_ni port map ( Y=>ordered_filter_data_13_3, A0=>
      filter_data_9_3, A1=>filter_data_4_3, S0=>nx1225);
   ix1575 : mux21_ni port map ( Y=>ordered_filter_data_13_4, A0=>
      filter_data_9_4, A1=>filter_data_4_4, S0=>nx1225);
   ix1583 : mux21_ni port map ( Y=>ordered_filter_data_13_5, A0=>
      filter_data_9_5, A1=>filter_data_4_5, S0=>nx1225);
   ix1591 : mux21_ni port map ( Y=>ordered_filter_data_13_6, A0=>
      filter_data_9_6, A1=>filter_data_4_6, S0=>nx1227);
   ix1599 : mux21_ni port map ( Y=>ordered_filter_data_13_7, A0=>
      filter_data_9_7, A1=>filter_data_4_7, S0=>nx1227);
   ix1607 : mux21_ni port map ( Y=>ordered_filter_data_13_8, A0=>
      filter_data_9_8, A1=>filter_data_4_8, S0=>nx1227);
   ix1615 : mux21_ni port map ( Y=>ordered_filter_data_13_9, A0=>
      filter_data_9_9, A1=>filter_data_4_9, S0=>nx1227);
   ix1623 : mux21_ni port map ( Y=>ordered_filter_data_13_10, A0=>
      filter_data_9_10, A1=>filter_data_4_10, S0=>nx1227);
   ix1631 : mux21_ni port map ( Y=>ordered_filter_data_13_11, A0=>
      filter_data_9_11, A1=>filter_data_4_11, S0=>nx1227);
   ix1639 : mux21_ni port map ( Y=>ordered_filter_data_13_12, A0=>
      filter_data_9_12, A1=>filter_data_4_12, S0=>nx1227);
   ix1647 : mux21_ni port map ( Y=>ordered_filter_data_13_13, A0=>
      filter_data_9_13, A1=>filter_data_4_13, S0=>nx1229);
   ix1655 : mux21_ni port map ( Y=>ordered_filter_data_13_14, A0=>
      filter_data_9_14, A1=>filter_data_4_14, S0=>nx1229);
   ix1663 : mux21_ni port map ( Y=>ordered_filter_data_13_15, A0=>
      filter_data_9_31, A1=>filter_data_4_31, S0=>nx1229);
   ix1927 : mux21_ni port map ( Y=>ordered_filter_data_12_0, A0=>
      filter_data_4_0, A1=>filter_data_3_0, S0=>nx1229);
   ix1935 : mux21_ni port map ( Y=>ordered_filter_data_12_1, A0=>
      filter_data_4_1, A1=>filter_data_3_1, S0=>nx1229);
   ix1943 : mux21_ni port map ( Y=>ordered_filter_data_12_2, A0=>
      filter_data_4_2, A1=>filter_data_3_2, S0=>nx1229);
   ix1951 : mux21_ni port map ( Y=>ordered_filter_data_12_3, A0=>
      filter_data_4_3, A1=>filter_data_3_3, S0=>nx1229);
   ix1959 : mux21_ni port map ( Y=>ordered_filter_data_12_4, A0=>
      filter_data_4_4, A1=>filter_data_3_4, S0=>nx1231);
   ix1967 : mux21_ni port map ( Y=>ordered_filter_data_12_5, A0=>
      filter_data_4_5, A1=>filter_data_3_5, S0=>nx1231);
   ix1975 : mux21_ni port map ( Y=>ordered_filter_data_12_6, A0=>
      filter_data_4_6, A1=>filter_data_3_6, S0=>nx1231);
   ix1983 : mux21_ni port map ( Y=>ordered_filter_data_12_7, A0=>
      filter_data_4_7, A1=>filter_data_3_7, S0=>nx1231);
   ix1991 : mux21_ni port map ( Y=>ordered_filter_data_12_8, A0=>
      filter_data_4_8, A1=>filter_data_3_8, S0=>nx1231);
   ix1999 : mux21_ni port map ( Y=>ordered_filter_data_12_9, A0=>
      filter_data_4_9, A1=>filter_data_3_9, S0=>nx1231);
   ix2007 : mux21_ni port map ( Y=>ordered_filter_data_12_10, A0=>
      filter_data_4_10, A1=>filter_data_3_10, S0=>nx1231);
   ix2015 : mux21_ni port map ( Y=>ordered_filter_data_12_11, A0=>
      filter_data_4_11, A1=>filter_data_3_11, S0=>nx1233);
   ix2023 : mux21_ni port map ( Y=>ordered_filter_data_12_12, A0=>
      filter_data_4_12, A1=>filter_data_3_12, S0=>nx1233);
   ix2031 : mux21_ni port map ( Y=>ordered_filter_data_12_13, A0=>
      filter_data_4_13, A1=>filter_data_3_13, S0=>nx1233);
   ix2039 : mux21_ni port map ( Y=>ordered_filter_data_12_14, A0=>
      filter_data_4_14, A1=>filter_data_3_14, S0=>nx1233);
   ix2047 : mux21_ni port map ( Y=>ordered_filter_data_12_15, A0=>
      filter_data_4_31, A1=>filter_data_3_31, S0=>nx1233);
   ix2311 : mux21_ni port map ( Y=>ordered_filter_data_11_0, A0=>
      filter_data_13_0, A1=>filter_data_2_0, S0=>nx1233);
   ix2319 : mux21_ni port map ( Y=>ordered_filter_data_11_1, A0=>
      filter_data_13_1, A1=>filter_data_2_1, S0=>nx1233);
   ix2327 : mux21_ni port map ( Y=>ordered_filter_data_11_2, A0=>
      filter_data_13_2, A1=>filter_data_2_2, S0=>nx1235);
   ix2335 : mux21_ni port map ( Y=>ordered_filter_data_11_3, A0=>
      filter_data_13_3, A1=>filter_data_2_3, S0=>nx1235);
   ix2343 : mux21_ni port map ( Y=>ordered_filter_data_11_4, A0=>
      filter_data_13_4, A1=>filter_data_2_4, S0=>nx1235);
   ix2351 : mux21_ni port map ( Y=>ordered_filter_data_11_5, A0=>
      filter_data_13_5, A1=>filter_data_2_5, S0=>nx1235);
   ix2359 : mux21_ni port map ( Y=>ordered_filter_data_11_6, A0=>
      filter_data_13_6, A1=>filter_data_2_6, S0=>nx1235);
   ix2367 : mux21_ni port map ( Y=>ordered_filter_data_11_7, A0=>
      filter_data_13_7, A1=>filter_data_2_7, S0=>nx1235);
   ix2375 : mux21_ni port map ( Y=>ordered_filter_data_11_8, A0=>
      filter_data_13_8, A1=>filter_data_2_8, S0=>nx1235);
   ix2383 : mux21_ni port map ( Y=>ordered_filter_data_11_9, A0=>
      filter_data_13_9, A1=>filter_data_2_9, S0=>nx1237);
   ix2391 : mux21_ni port map ( Y=>ordered_filter_data_11_10, A0=>
      filter_data_13_10, A1=>filter_data_2_10, S0=>nx1237);
   ix2399 : mux21_ni port map ( Y=>ordered_filter_data_11_11, A0=>
      filter_data_13_11, A1=>filter_data_2_11, S0=>nx1237);
   ix2407 : mux21_ni port map ( Y=>ordered_filter_data_11_12, A0=>
      filter_data_13_12, A1=>filter_data_2_12, S0=>nx1237);
   ix2415 : mux21_ni port map ( Y=>ordered_filter_data_11_13, A0=>
      filter_data_13_13, A1=>filter_data_2_13, S0=>nx1237);
   ix2423 : mux21_ni port map ( Y=>ordered_filter_data_11_14, A0=>
      filter_data_13_14, A1=>filter_data_2_14, S0=>nx1237);
   ix2431 : mux21_ni port map ( Y=>ordered_filter_data_11_15, A0=>
      filter_data_13_31, A1=>filter_data_2_31, S0=>nx1237);
   ix2567 : mux21_ni port map ( Y=>ordered_filter_data_10_0, A0=>
      filter_data_8_0, A1=>filter_data_1_0, S0=>nx1239);
   ix2575 : mux21_ni port map ( Y=>ordered_filter_data_10_1, A0=>
      filter_data_8_1, A1=>filter_data_1_1, S0=>nx1239);
   ix2583 : mux21_ni port map ( Y=>ordered_filter_data_10_2, A0=>
      filter_data_8_2, A1=>filter_data_1_2, S0=>nx1239);
   ix2591 : mux21_ni port map ( Y=>ordered_filter_data_10_3, A0=>
      filter_data_8_3, A1=>filter_data_1_3, S0=>nx1239);
   ix2599 : mux21_ni port map ( Y=>ordered_filter_data_10_4, A0=>
      filter_data_8_4, A1=>filter_data_1_4, S0=>nx1239);
   ix2607 : mux21_ni port map ( Y=>ordered_filter_data_10_5, A0=>
      filter_data_8_5, A1=>filter_data_1_5, S0=>nx1239);
   ix2615 : mux21_ni port map ( Y=>ordered_filter_data_10_6, A0=>
      filter_data_8_6, A1=>filter_data_1_6, S0=>nx1239);
   ix2623 : mux21_ni port map ( Y=>ordered_filter_data_10_7, A0=>
      filter_data_8_7, A1=>filter_data_1_7, S0=>nx1241);
   ix2631 : mux21_ni port map ( Y=>ordered_filter_data_10_8, A0=>
      filter_data_8_8, A1=>filter_data_1_8, S0=>nx1241);
   ix2639 : mux21_ni port map ( Y=>ordered_filter_data_10_9, A0=>
      filter_data_8_9, A1=>filter_data_1_9, S0=>nx1241);
   ix2647 : mux21_ni port map ( Y=>ordered_filter_data_10_10, A0=>
      filter_data_8_10, A1=>filter_data_1_10, S0=>nx1241);
   ix2655 : mux21_ni port map ( Y=>ordered_filter_data_10_11, A0=>
      filter_data_8_11, A1=>filter_data_1_11, S0=>nx1241);
   ix2663 : mux21_ni port map ( Y=>ordered_filter_data_10_12, A0=>
      filter_data_8_12, A1=>filter_data_1_12, S0=>nx1241);
   ix2671 : mux21_ni port map ( Y=>ordered_filter_data_10_13, A0=>
      filter_data_8_13, A1=>filter_data_1_13, S0=>nx1241);
   ix2679 : mux21_ni port map ( Y=>ordered_filter_data_10_14, A0=>
      filter_data_8_14, A1=>filter_data_1_14, S0=>nx1243);
   ix2687 : mux21_ni port map ( Y=>ordered_filter_data_10_15, A0=>
      filter_data_8_31, A1=>filter_data_1_31, S0=>nx1243);
   ix2823 : mux21_ni port map ( Y=>ordered_filter_data_9_0, A0=>
      filter_data_3_0, A1=>filter_data_0_0, S0=>nx1243);
   ix2831 : mux21_ni port map ( Y=>ordered_filter_data_9_1, A0=>
      filter_data_3_1, A1=>filter_data_0_1, S0=>nx1243);
   ix2839 : mux21_ni port map ( Y=>ordered_filter_data_9_2, A0=>
      filter_data_3_2, A1=>filter_data_0_2, S0=>nx1243);
   ix2847 : mux21_ni port map ( Y=>ordered_filter_data_9_3, A0=>
      filter_data_3_3, A1=>filter_data_0_3, S0=>nx1243);
   ix2855 : mux21_ni port map ( Y=>ordered_filter_data_9_4, A0=>
      filter_data_3_4, A1=>filter_data_0_4, S0=>nx1243);
   ix2863 : mux21_ni port map ( Y=>ordered_filter_data_9_5, A0=>
      filter_data_3_5, A1=>filter_data_0_5, S0=>nx1245);
   ix2871 : mux21_ni port map ( Y=>ordered_filter_data_9_6, A0=>
      filter_data_3_6, A1=>filter_data_0_6, S0=>nx1245);
   ix2879 : mux21_ni port map ( Y=>ordered_filter_data_9_7, A0=>
      filter_data_3_7, A1=>filter_data_0_7, S0=>nx1245);
   ix2887 : mux21_ni port map ( Y=>ordered_filter_data_9_8, A0=>
      filter_data_3_8, A1=>filter_data_0_8, S0=>nx1245);
   ix2895 : mux21_ni port map ( Y=>ordered_filter_data_9_9, A0=>
      filter_data_3_9, A1=>filter_data_0_9, S0=>nx1245);
   ix2903 : mux21_ni port map ( Y=>ordered_filter_data_9_10, A0=>
      filter_data_3_10, A1=>filter_data_0_10, S0=>nx1245);
   ix2911 : mux21_ni port map ( Y=>ordered_filter_data_9_11, A0=>
      filter_data_3_11, A1=>filter_data_0_11, S0=>nx1245);
   ix2919 : mux21_ni port map ( Y=>ordered_filter_data_9_12, A0=>
      filter_data_3_12, A1=>filter_data_0_12, S0=>nx1247);
   ix2927 : mux21_ni port map ( Y=>ordered_filter_data_9_13, A0=>
      filter_data_3_13, A1=>filter_data_0_13, S0=>nx1247);
   ix2935 : mux21_ni port map ( Y=>ordered_filter_data_9_14, A0=>
      filter_data_3_14, A1=>filter_data_0_14, S0=>nx1247);
   ix2943 : mux21_ni port map ( Y=>ordered_filter_data_9_15, A0=>
      filter_data_3_31, A1=>filter_data_0_31, S0=>nx1247);
   ix263 : mux21_ni port map ( Y=>ordered_filter_data_8_0, A0=>
      filter_data_12_0, A1=>filter_data_8_0, S0=>nx1247);
   ix271 : mux21_ni port map ( Y=>ordered_filter_data_8_1, A0=>
      filter_data_12_1, A1=>filter_data_8_1, S0=>nx1247);
   ix279 : mux21_ni port map ( Y=>ordered_filter_data_8_2, A0=>
      filter_data_12_2, A1=>filter_data_8_2, S0=>nx1247);
   ix287 : mux21_ni port map ( Y=>ordered_filter_data_8_3, A0=>
      filter_data_12_3, A1=>filter_data_8_3, S0=>nx1249);
   ix295 : mux21_ni port map ( Y=>ordered_filter_data_8_4, A0=>
      filter_data_12_4, A1=>filter_data_8_4, S0=>nx1249);
   ix303 : mux21_ni port map ( Y=>ordered_filter_data_8_5, A0=>
      filter_data_12_5, A1=>filter_data_8_5, S0=>nx1249);
   ix311 : mux21_ni port map ( Y=>ordered_filter_data_8_6, A0=>
      filter_data_12_6, A1=>filter_data_8_6, S0=>nx1249);
   ix319 : mux21_ni port map ( Y=>ordered_filter_data_8_7, A0=>
      filter_data_12_7, A1=>filter_data_8_7, S0=>nx1249);
   ix327 : mux21_ni port map ( Y=>ordered_filter_data_8_8, A0=>
      filter_data_12_8, A1=>filter_data_8_8, S0=>nx1249);
   ix335 : mux21_ni port map ( Y=>ordered_filter_data_8_9, A0=>
      filter_data_12_9, A1=>filter_data_8_9, S0=>nx1249);
   ix343 : mux21_ni port map ( Y=>ordered_filter_data_8_10, A0=>
      filter_data_12_10, A1=>filter_data_8_10, S0=>nx1251);
   ix351 : mux21_ni port map ( Y=>ordered_filter_data_8_11, A0=>
      filter_data_12_11, A1=>filter_data_8_11, S0=>nx1251);
   ix359 : mux21_ni port map ( Y=>ordered_filter_data_8_12, A0=>
      filter_data_12_12, A1=>filter_data_8_12, S0=>nx1251);
   ix367 : mux21_ni port map ( Y=>ordered_filter_data_8_13, A0=>
      filter_data_12_13, A1=>filter_data_8_13, S0=>nx1251);
   ix375 : mux21_ni port map ( Y=>ordered_filter_data_8_14, A0=>
      filter_data_12_14, A1=>filter_data_8_14, S0=>nx1251);
   ix383 : mux21_ni port map ( Y=>ordered_filter_data_8_15, A0=>
      filter_data_12_31, A1=>filter_data_8_31, S0=>nx1251);
   ix647 : mux21_ni port map ( Y=>ordered_filter_data_7_0, A0=>
      filter_data_11_0, A1=>filter_data_7_0, S0=>nx1251);
   ix655 : mux21_ni port map ( Y=>ordered_filter_data_7_1, A0=>
      filter_data_11_1, A1=>filter_data_7_1, S0=>nx1253);
   ix663 : mux21_ni port map ( Y=>ordered_filter_data_7_2, A0=>
      filter_data_11_2, A1=>filter_data_7_2, S0=>nx1253);
   ix671 : mux21_ni port map ( Y=>ordered_filter_data_7_3, A0=>
      filter_data_11_3, A1=>filter_data_7_3, S0=>nx1253);
   ix679 : mux21_ni port map ( Y=>ordered_filter_data_7_4, A0=>
      filter_data_11_4, A1=>filter_data_7_4, S0=>nx1253);
   ix687 : mux21_ni port map ( Y=>ordered_filter_data_7_5, A0=>
      filter_data_11_5, A1=>filter_data_7_5, S0=>nx1253);
   ix695 : mux21_ni port map ( Y=>ordered_filter_data_7_6, A0=>
      filter_data_11_6, A1=>filter_data_7_6, S0=>nx1253);
   ix703 : mux21_ni port map ( Y=>ordered_filter_data_7_7, A0=>
      filter_data_11_7, A1=>filter_data_7_7, S0=>nx1253);
   ix711 : mux21_ni port map ( Y=>ordered_filter_data_7_8, A0=>
      filter_data_11_8, A1=>filter_data_7_8, S0=>nx1255);
   ix719 : mux21_ni port map ( Y=>ordered_filter_data_7_9, A0=>
      filter_data_11_9, A1=>filter_data_7_9, S0=>nx1255);
   ix727 : mux21_ni port map ( Y=>ordered_filter_data_7_10, A0=>
      filter_data_11_10, A1=>filter_data_7_10, S0=>nx1255);
   ix735 : mux21_ni port map ( Y=>ordered_filter_data_7_11, A0=>
      filter_data_11_11, A1=>filter_data_7_11, S0=>nx1255);
   ix743 : mux21_ni port map ( Y=>ordered_filter_data_7_12, A0=>
      filter_data_11_12, A1=>filter_data_7_12, S0=>nx1255);
   ix751 : mux21_ni port map ( Y=>ordered_filter_data_7_13, A0=>
      filter_data_11_13, A1=>filter_data_7_13, S0=>nx1255);
   ix759 : mux21_ni port map ( Y=>ordered_filter_data_7_14, A0=>
      filter_data_11_14, A1=>filter_data_7_14, S0=>nx1255);
   ix767 : mux21_ni port map ( Y=>ordered_filter_data_7_15, A0=>
      filter_data_11_31, A1=>filter_data_7_31, S0=>nx1257);
   ix1031 : mux21_ni port map ( Y=>ordered_filter_data_6_0, A0=>
      filter_data_10_0, A1=>filter_data_6_0, S0=>nx1257);
   ix1039 : mux21_ni port map ( Y=>ordered_filter_data_6_1, A0=>
      filter_data_10_1, A1=>filter_data_6_1, S0=>nx1257);
   ix1047 : mux21_ni port map ( Y=>ordered_filter_data_6_2, A0=>
      filter_data_10_2, A1=>filter_data_6_2, S0=>nx1257);
   ix1055 : mux21_ni port map ( Y=>ordered_filter_data_6_3, A0=>
      filter_data_10_3, A1=>filter_data_6_3, S0=>nx1257);
   ix1063 : mux21_ni port map ( Y=>ordered_filter_data_6_4, A0=>
      filter_data_10_4, A1=>filter_data_6_4, S0=>nx1257);
   ix1071 : mux21_ni port map ( Y=>ordered_filter_data_6_5, A0=>
      filter_data_10_5, A1=>filter_data_6_5, S0=>nx1257);
   ix1079 : mux21_ni port map ( Y=>ordered_filter_data_6_6, A0=>
      filter_data_10_6, A1=>filter_data_6_6, S0=>nx1259);
   ix1087 : mux21_ni port map ( Y=>ordered_filter_data_6_7, A0=>
      filter_data_10_7, A1=>filter_data_6_7, S0=>nx1259);
   ix1095 : mux21_ni port map ( Y=>ordered_filter_data_6_8, A0=>
      filter_data_10_8, A1=>filter_data_6_8, S0=>nx1259);
   ix1103 : mux21_ni port map ( Y=>ordered_filter_data_6_9, A0=>
      filter_data_10_9, A1=>filter_data_6_9, S0=>nx1259);
   ix1111 : mux21_ni port map ( Y=>ordered_filter_data_6_10, A0=>
      filter_data_10_10, A1=>filter_data_6_10, S0=>nx1259);
   ix1119 : mux21_ni port map ( Y=>ordered_filter_data_6_11, A0=>
      filter_data_10_11, A1=>filter_data_6_11, S0=>nx1259);
   ix1127 : mux21_ni port map ( Y=>ordered_filter_data_6_12, A0=>
      filter_data_10_12, A1=>filter_data_6_12, S0=>nx1259);
   ix1135 : mux21_ni port map ( Y=>ordered_filter_data_6_13, A0=>
      filter_data_10_13, A1=>filter_data_6_13, S0=>nx1261);
   ix1143 : mux21_ni port map ( Y=>ordered_filter_data_6_14, A0=>
      filter_data_10_14, A1=>filter_data_6_14, S0=>nx1261);
   ix1151 : mux21_ni port map ( Y=>ordered_filter_data_6_15, A0=>
      filter_data_10_31, A1=>filter_data_6_31, S0=>nx1261);
   ix1415 : mux21_ni port map ( Y=>ordered_filter_data_5_0, A0=>
      filter_data_7_0, A1=>filter_data_5_0, S0=>nx1261);
   ix1423 : mux21_ni port map ( Y=>ordered_filter_data_5_1, A0=>
      filter_data_7_1, A1=>filter_data_5_1, S0=>nx1261);
   ix1431 : mux21_ni port map ( Y=>ordered_filter_data_5_2, A0=>
      filter_data_7_2, A1=>filter_data_5_2, S0=>nx1261);
   ix1439 : mux21_ni port map ( Y=>ordered_filter_data_5_3, A0=>
      filter_data_7_3, A1=>filter_data_5_3, S0=>nx1261);
   ix1447 : mux21_ni port map ( Y=>ordered_filter_data_5_4, A0=>
      filter_data_7_4, A1=>filter_data_5_4, S0=>nx1263);
   ix1455 : mux21_ni port map ( Y=>ordered_filter_data_5_5, A0=>
      filter_data_7_5, A1=>filter_data_5_5, S0=>nx1263);
   ix1463 : mux21_ni port map ( Y=>ordered_filter_data_5_6, A0=>
      filter_data_7_6, A1=>filter_data_5_6, S0=>nx1263);
   ix1471 : mux21_ni port map ( Y=>ordered_filter_data_5_7, A0=>
      filter_data_7_7, A1=>filter_data_5_7, S0=>nx1263);
   ix1479 : mux21_ni port map ( Y=>ordered_filter_data_5_8, A0=>
      filter_data_7_8, A1=>filter_data_5_8, S0=>nx1263);
   ix1487 : mux21_ni port map ( Y=>ordered_filter_data_5_9, A0=>
      filter_data_7_9, A1=>filter_data_5_9, S0=>nx1263);
   ix1495 : mux21_ni port map ( Y=>ordered_filter_data_5_10, A0=>
      filter_data_7_10, A1=>filter_data_5_10, S0=>nx1263);
   ix1503 : mux21_ni port map ( Y=>ordered_filter_data_5_11, A0=>
      filter_data_7_11, A1=>filter_data_5_11, S0=>nx1265);
   ix1511 : mux21_ni port map ( Y=>ordered_filter_data_5_12, A0=>
      filter_data_7_12, A1=>filter_data_5_12, S0=>nx1265);
   ix1519 : mux21_ni port map ( Y=>ordered_filter_data_5_13, A0=>
      filter_data_7_13, A1=>filter_data_5_13, S0=>nx1265);
   ix1527 : mux21_ni port map ( Y=>ordered_filter_data_5_14, A0=>
      filter_data_7_14, A1=>filter_data_5_14, S0=>nx1265);
   ix1535 : mux21_ni port map ( Y=>ordered_filter_data_5_15, A0=>
      filter_data_7_31, A1=>filter_data_5_31, S0=>nx1265);
   ix1799 : mux21_ni port map ( Y=>ordered_filter_data_4_0, A0=>
      filter_data_6_0, A1=>filter_data_4_0, S0=>nx1265);
   ix1807 : mux21_ni port map ( Y=>ordered_filter_data_4_1, A0=>
      filter_data_6_1, A1=>filter_data_4_1, S0=>nx1265);
   ix1815 : mux21_ni port map ( Y=>ordered_filter_data_4_2, A0=>
      filter_data_6_2, A1=>filter_data_4_2, S0=>nx1267);
   ix1823 : mux21_ni port map ( Y=>ordered_filter_data_4_3, A0=>
      filter_data_6_3, A1=>filter_data_4_3, S0=>nx1267);
   ix1831 : mux21_ni port map ( Y=>ordered_filter_data_4_4, A0=>
      filter_data_6_4, A1=>filter_data_4_4, S0=>nx1267);
   ix1839 : mux21_ni port map ( Y=>ordered_filter_data_4_5, A0=>
      filter_data_6_5, A1=>filter_data_4_5, S0=>nx1267);
   ix1847 : mux21_ni port map ( Y=>ordered_filter_data_4_6, A0=>
      filter_data_6_6, A1=>filter_data_4_6, S0=>nx1267);
   ix1855 : mux21_ni port map ( Y=>ordered_filter_data_4_7, A0=>
      filter_data_6_7, A1=>filter_data_4_7, S0=>nx1267);
   ix1863 : mux21_ni port map ( Y=>ordered_filter_data_4_8, A0=>
      filter_data_6_8, A1=>filter_data_4_8, S0=>nx1267);
   ix1871 : mux21_ni port map ( Y=>ordered_filter_data_4_9, A0=>
      filter_data_6_9, A1=>filter_data_4_9, S0=>nx1269);
   ix1879 : mux21_ni port map ( Y=>ordered_filter_data_4_10, A0=>
      filter_data_6_10, A1=>filter_data_4_10, S0=>nx1269);
   ix1887 : mux21_ni port map ( Y=>ordered_filter_data_4_11, A0=>
      filter_data_6_11, A1=>filter_data_4_11, S0=>nx1269);
   ix1895 : mux21_ni port map ( Y=>ordered_filter_data_4_12, A0=>
      filter_data_6_12, A1=>filter_data_4_12, S0=>nx1269);
   ix1903 : mux21_ni port map ( Y=>ordered_filter_data_4_13, A0=>
      filter_data_6_13, A1=>filter_data_4_13, S0=>nx1269);
   ix1911 : mux21_ni port map ( Y=>ordered_filter_data_4_14, A0=>
      filter_data_6_14, A1=>filter_data_4_14, S0=>nx1269);
   ix1919 : mux21_ni port map ( Y=>ordered_filter_data_4_15, A0=>
      filter_data_6_31, A1=>filter_data_4_31, S0=>nx1269);
   ix2183 : mux21_ni port map ( Y=>ordered_filter_data_3_0, A0=>
      filter_data_5_0, A1=>filter_data_3_0, S0=>nx1271);
   ix2191 : mux21_ni port map ( Y=>ordered_filter_data_3_1, A0=>
      filter_data_5_1, A1=>filter_data_3_1, S0=>nx1271);
   ix2199 : mux21_ni port map ( Y=>ordered_filter_data_3_2, A0=>
      filter_data_5_2, A1=>filter_data_3_2, S0=>nx1271);
   ix2207 : mux21_ni port map ( Y=>ordered_filter_data_3_3, A0=>
      filter_data_5_3, A1=>filter_data_3_3, S0=>nx1271);
   ix2215 : mux21_ni port map ( Y=>ordered_filter_data_3_4, A0=>
      filter_data_5_4, A1=>filter_data_3_4, S0=>nx1271);
   ix2223 : mux21_ni port map ( Y=>ordered_filter_data_3_5, A0=>
      filter_data_5_5, A1=>filter_data_3_5, S0=>nx1271);
   ix2231 : mux21_ni port map ( Y=>ordered_filter_data_3_6, A0=>
      filter_data_5_6, A1=>filter_data_3_6, S0=>nx1271);
   ix2239 : mux21_ni port map ( Y=>ordered_filter_data_3_7, A0=>
      filter_data_5_7, A1=>filter_data_3_7, S0=>nx1273);
   ix2247 : mux21_ni port map ( Y=>ordered_filter_data_3_8, A0=>
      filter_data_5_8, A1=>filter_data_3_8, S0=>nx1273);
   ix2255 : mux21_ni port map ( Y=>ordered_filter_data_3_9, A0=>
      filter_data_5_9, A1=>filter_data_3_9, S0=>nx1273);
   ix2263 : mux21_ni port map ( Y=>ordered_filter_data_3_10, A0=>
      filter_data_5_10, A1=>filter_data_3_10, S0=>nx1273);
   ix2271 : mux21_ni port map ( Y=>ordered_filter_data_3_11, A0=>
      filter_data_5_11, A1=>filter_data_3_11, S0=>nx1273);
   ix2279 : mux21_ni port map ( Y=>ordered_filter_data_3_12, A0=>
      filter_data_5_12, A1=>filter_data_3_12, S0=>nx1273);
   ix2287 : mux21_ni port map ( Y=>ordered_filter_data_3_13, A0=>
      filter_data_5_13, A1=>filter_data_3_13, S0=>nx1273);
   ix2295 : mux21_ni port map ( Y=>ordered_filter_data_3_14, A0=>
      filter_data_5_14, A1=>filter_data_3_14, S0=>nx1354);
   ix2303 : mux21_ni port map ( Y=>ordered_filter_data_3_15, A0=>
      filter_data_5_31, A1=>filter_data_3_31, S0=>nx1354);
   ix143 : mux21_ni port map ( Y=>ordered_img_data_17_1, A0=>img_data_17_1, 
      A1=>img_data_13_1, S0=>nx1354);
   ix151 : mux21_ni port map ( Y=>ordered_img_data_17_2, A0=>img_data_17_2, 
      A1=>img_data_13_2, S0=>nx1354);
   ix159 : mux21_ni port map ( Y=>ordered_img_data_17_3, A0=>img_data_17_3, 
      A1=>img_data_13_3, S0=>nx1354);
   ix167 : mux21_ni port map ( Y=>ordered_img_data_17_4, A0=>img_data_17_4, 
      A1=>img_data_13_4, S0=>nx1354);
   ix183 : mux21_ni port map ( Y=>ordered_img_data_17_6, A0=>img_data_17_6, 
      A1=>img_data_13_6, S0=>nx1354);
   ix191 : mux21_ni port map ( Y=>ordered_img_data_17_7, A0=>img_data_17_7, 
      A1=>img_data_13_7, S0=>nx1356);
   ix199 : mux21_ni port map ( Y=>ordered_img_data_17_8, A0=>img_data_17_8, 
      A1=>img_data_13_8, S0=>nx1356);
   ix207 : mux21_ni port map ( Y=>ordered_img_data_17_9, A0=>img_data_17_9, 
      A1=>img_data_13_9, S0=>nx1356);
   ix215 : mux21_ni port map ( Y=>ordered_img_data_17_10, A0=>img_data_17_10, 
      A1=>img_data_13_10, S0=>nx1356);
   ix223 : mux21_ni port map ( Y=>ordered_img_data_17_11, A0=>img_data_17_11, 
      A1=>img_data_13_11, S0=>nx1356);
   ix231 : mux21_ni port map ( Y=>ordered_img_data_17_12, A0=>img_data_17_12, 
      A1=>img_data_13_12, S0=>nx1356);
   ix239 : mux21_ni port map ( Y=>ordered_img_data_17_13, A0=>img_data_17_13, 
      A1=>img_data_13_13, S0=>nx1356);
   ix247 : mux21_ni port map ( Y=>ordered_img_data_17_14, A0=>img_data_17_14, 
      A1=>img_data_13_14, S0=>nx1358);
   ix255 : mux21_ni port map ( Y=>ordered_img_data_17_15_EXMPLR, A0=>
      img_data_17_31, A1=>img_data_13_31, S0=>nx1358);
   ix519 : mux21_ni port map ( Y=>ordered_img_data_16_0, A0=>img_data_16_0, 
      A1=>img_data_12_0, S0=>nx1358);
   ix535 : mux21_ni port map ( Y=>ordered_img_data_16_2, A0=>img_data_16_2, 
      A1=>img_data_12_2, S0=>nx1358);
   ix543 : mux21_ni port map ( Y=>ordered_img_data_16_3, A0=>img_data_16_3, 
      A1=>img_data_12_3, S0=>nx1358);
   ix551 : mux21_ni port map ( Y=>ordered_img_data_16_4, A0=>img_data_16_4, 
      A1=>img_data_12_4, S0=>nx1358);
   ix559 : mux21_ni port map ( Y=>ordered_img_data_16_5, A0=>img_data_16_5, 
      A1=>img_data_12_5, S0=>nx1358);
   ix567 : mux21_ni port map ( Y=>ordered_img_data_16_6, A0=>img_data_16_6, 
      A1=>img_data_12_6, S0=>nx1361);
   ix583 : mux21_ni port map ( Y=>ordered_img_data_16_8, A0=>img_data_16_8, 
      A1=>img_data_12_8, S0=>nx1361);
   ix591 : mux21_ni port map ( Y=>ordered_img_data_16_9, A0=>img_data_16_9, 
      A1=>img_data_12_9, S0=>nx1361);
   ix599 : mux21_ni port map ( Y=>ordered_img_data_16_10, A0=>img_data_16_10, 
      A1=>img_data_12_10, S0=>nx1361);
   ix607 : mux21_ni port map ( Y=>ordered_img_data_16_11, A0=>img_data_16_11, 
      A1=>img_data_12_11, S0=>nx1361);
   ix615 : mux21_ni port map ( Y=>ordered_img_data_16_12, A0=>img_data_16_12, 
      A1=>img_data_12_12, S0=>nx1361);
   ix623 : mux21_ni port map ( Y=>ordered_img_data_16_13, A0=>img_data_16_13, 
      A1=>img_data_12_13, S0=>nx1361);
   ix631 : mux21_ni port map ( Y=>ordered_img_data_16_14, A0=>img_data_16_14, 
      A1=>img_data_12_14, S0=>nx1363);
   ix639 : mux21_ni port map ( Y=>ordered_img_data_16_15_EXMPLR, A0=>
      img_data_16_31, A1=>img_data_12_31, S0=>nx1363);
   ix911 : mux21_ni port map ( Y=>ordered_img_data_15_1, A0=>img_data_15_1, 
      A1=>img_data_11_1, S0=>nx1363);
   ix919 : mux21_ni port map ( Y=>ordered_img_data_15_2, A0=>img_data_15_2, 
      A1=>img_data_11_2, S0=>nx1363);
   ix927 : mux21_ni port map ( Y=>ordered_img_data_15_3, A0=>img_data_15_3, 
      A1=>img_data_11_3, S0=>nx1363);
   ix935 : mux21_ni port map ( Y=>ordered_img_data_15_4, A0=>img_data_15_4, 
      A1=>img_data_11_4, S0=>nx1363);
   ix943 : mux21_ni port map ( Y=>ordered_img_data_15_5, A0=>img_data_15_5, 
      A1=>img_data_11_5, S0=>nx1363);
   ix951 : mux21_ni port map ( Y=>ordered_img_data_15_6, A0=>img_data_15_6, 
      A1=>img_data_11_6, S0=>nx1365);
   ix967 : mux21_ni port map ( Y=>ordered_img_data_15_8, A0=>img_data_15_8, 
      A1=>img_data_11_8, S0=>nx1287);
   ix975 : mux21_ni port map ( Y=>ordered_img_data_15_9, A0=>img_data_15_9, 
      A1=>img_data_11_9, S0=>nx1287);
   ix983 : mux21_ni port map ( Y=>ordered_img_data_15_10, A0=>img_data_15_10, 
      A1=>img_data_11_10, S0=>nx1287);
   ix991 : mux21_ni port map ( Y=>ordered_img_data_15_11, A0=>img_data_15_11, 
      A1=>img_data_11_11, S0=>nx1287);
   ix999 : mux21_ni port map ( Y=>ordered_img_data_15_12, A0=>img_data_15_12, 
      A1=>img_data_11_12, S0=>nx1287);
   ix1007 : mux21_ni port map ( Y=>ordered_img_data_15_13, A0=>
      img_data_15_13, A1=>img_data_11_13, S0=>nx1287);
   ix1015 : mux21_ni port map ( Y=>ordered_img_data_15_14, A0=>
      img_data_15_14, A1=>img_data_11_14, S0=>nx1287);
   ix1023 : mux21_ni port map ( Y=>ordered_img_data_15_15_EXMPLR, A0=>
      img_data_15_31, A1=>img_data_11_31, S0=>nx1365);
   ix1287 : mux21_ni port map ( Y=>ordered_img_data_14_0, A0=>img_data_14_0, 
      A1=>img_data_8_0, S0=>nx1365);
   ix1295 : mux21_ni port map ( Y=>ordered_img_data_14_1, A0=>img_data_14_1, 
      A1=>img_data_8_1, S0=>nx1365);
   ix1303 : mux21_ni port map ( Y=>ordered_img_data_14_2, A0=>img_data_14_2, 
      A1=>img_data_8_2, S0=>nx1365);
   ix1319 : mux21_ni port map ( Y=>ordered_img_data_14_4, A0=>img_data_14_4, 
      A1=>img_data_8_4, S0=>nx1365);
   ix1327 : mux21_ni port map ( Y=>ordered_img_data_14_5, A0=>img_data_14_5, 
      A1=>img_data_8_5, S0=>nx1365);
   ix1335 : mux21_ni port map ( Y=>ordered_img_data_14_6, A0=>img_data_14_6, 
      A1=>img_data_8_6, S0=>nx1367);
   ix1351 : mux21_ni port map ( Y=>ordered_img_data_14_8, A0=>img_data_14_8, 
      A1=>img_data_8_8, S0=>nx1367);
   ix1359 : mux21_ni port map ( Y=>ordered_img_data_14_9, A0=>img_data_14_9, 
      A1=>img_data_8_9, S0=>nx1367);
   ix1367 : mux21_ni port map ( Y=>ordered_img_data_14_10, A0=>
      img_data_14_10, A1=>img_data_8_10, S0=>nx1367);
   ix1375 : mux21_ni port map ( Y=>ordered_img_data_14_11, A0=>
      img_data_14_11, A1=>img_data_8_11, S0=>nx1367);
   ix1383 : mux21_ni port map ( Y=>ordered_img_data_14_12, A0=>
      img_data_14_12, A1=>img_data_8_12, S0=>nx1367);
   ix1391 : mux21_ni port map ( Y=>ordered_img_data_14_13, A0=>
      img_data_14_13, A1=>img_data_8_13, S0=>nx1367);
   ix1399 : mux21_ni port map ( Y=>ordered_img_data_14_14, A0=>
      img_data_14_14, A1=>img_data_8_14, S0=>nx1369);
   ix1407 : mux21_ni port map ( Y=>ordered_img_data_14_15_EXMPLR, A0=>
      img_data_14_31, A1=>img_data_8_31, S0=>nx1369);
   ix1671 : mux21_ni port map ( Y=>ordered_img_data_13_0, A0=>img_data_9_0, 
      A1=>img_data_7_0, S0=>nx1369);
   ix1679 : mux21_ni port map ( Y=>ordered_img_data_13_1, A0=>img_data_9_1, 
      A1=>img_data_7_1, S0=>nx1369);
   ix1687 : mux21_ni port map ( Y=>ordered_img_data_13_2, A0=>img_data_9_2, 
      A1=>img_data_7_2, S0=>nx1369);
   ix1703 : mux21_ni port map ( Y=>ordered_img_data_13_4, A0=>img_data_9_4, 
      A1=>img_data_7_4, S0=>nx1369);
   ix1719 : mux21_ni port map ( Y=>ordered_img_data_13_6, A0=>img_data_9_6, 
      A1=>img_data_7_6, S0=>nx1369);
   ix1727 : mux21_ni port map ( Y=>ordered_img_data_13_7, A0=>img_data_9_7, 
      A1=>img_data_7_7, S0=>nx1371);
   ix1735 : mux21_ni port map ( Y=>ordered_img_data_13_8, A0=>img_data_9_8, 
      A1=>img_data_7_8, S0=>nx1371);
   ix1743 : mux21_ni port map ( Y=>ordered_img_data_13_9, A0=>img_data_9_9, 
      A1=>img_data_7_9, S0=>nx1371);
   ix1751 : mux21_ni port map ( Y=>ordered_img_data_13_10, A0=>img_data_9_10, 
      A1=>img_data_7_10, S0=>nx1371);
   ix1759 : mux21_ni port map ( Y=>ordered_img_data_13_11, A0=>img_data_9_11, 
      A1=>img_data_7_11, S0=>nx1371);
   ix1767 : mux21_ni port map ( Y=>ordered_img_data_13_12, A0=>img_data_9_12, 
      A1=>img_data_7_12, S0=>nx1371);
   ix1775 : mux21_ni port map ( Y=>ordered_img_data_13_13, A0=>img_data_9_13, 
      A1=>img_data_7_13, S0=>nx1371);
   ix1783 : mux21_ni port map ( Y=>ordered_img_data_13_14, A0=>img_data_9_14, 
      A1=>img_data_7_14, S0=>nx1373);
   ix1791 : mux21_ni port map ( Y=>ordered_img_data_13_15_EXMPLR, A0=>
      img_data_9_31, A1=>img_data_7_31, S0=>nx1373);
   ix2063 : mux21_ni port map ( Y=>ordered_img_data_12_1, A0=>img_data_4_1, 
      A1=>img_data_6_1, S0=>nx1373);
   ix2071 : mux21_ni port map ( Y=>ordered_img_data_12_2, A0=>img_data_4_2, 
      A1=>img_data_6_2, S0=>nx1373);
   ix2079 : mux21_ni port map ( Y=>ordered_img_data_12_3, A0=>img_data_4_3, 
      A1=>img_data_6_3, S0=>nx1373);
   ix2095 : mux21_ni port map ( Y=>ordered_img_data_12_5, A0=>img_data_4_5, 
      A1=>img_data_6_5, S0=>nx1373);
   ix2103 : mux21_ni port map ( Y=>ordered_img_data_12_6, A0=>img_data_4_6, 
      A1=>img_data_6_6, S0=>nx1373);
   ix2111 : mux21_ni port map ( Y=>ordered_img_data_12_7, A0=>img_data_4_7, 
      A1=>img_data_6_7, S0=>nx1375);
   ix2119 : mux21_ni port map ( Y=>ordered_img_data_12_8, A0=>img_data_4_8, 
      A1=>img_data_6_8, S0=>nx1375);
   ix2127 : mux21_ni port map ( Y=>ordered_img_data_12_9, A0=>img_data_4_9, 
      A1=>img_data_6_9, S0=>nx1301);
   ix2135 : mux21_ni port map ( Y=>ordered_img_data_12_10, A0=>img_data_4_10, 
      A1=>img_data_6_10, S0=>nx1301);
   ix2143 : mux21_ni port map ( Y=>ordered_img_data_12_11, A0=>img_data_4_11, 
      A1=>img_data_6_11, S0=>nx1301);
   ix2151 : mux21_ni port map ( Y=>ordered_img_data_12_12, A0=>img_data_4_12, 
      A1=>img_data_6_12, S0=>nx1301);
   ix2159 : mux21_ni port map ( Y=>ordered_img_data_12_13, A0=>img_data_4_13, 
      A1=>img_data_6_13, S0=>nx1301);
   ix2167 : mux21_ni port map ( Y=>ordered_img_data_12_14, A0=>img_data_4_14, 
      A1=>img_data_6_14, S0=>nx1301);
   ix2175 : mux21_ni port map ( Y=>ordered_img_data_12_15_EXMPLR, A0=>
      img_data_4_31, A1=>img_data_6_31, S0=>nx1301);
   ix2439 : mux21_ni port map ( Y=>ordered_img_data_11_0, A0=>img_data_13_0, 
      A1=>img_data_3_0, S0=>nx1375);
   ix2447 : mux21_ni port map ( Y=>ordered_img_data_11_1, A0=>img_data_13_1, 
      A1=>img_data_3_1, S0=>nx1375);
   ix2463 : mux21_ni port map ( Y=>ordered_img_data_11_3, A0=>img_data_13_3, 
      A1=>img_data_3_3, S0=>nx1375);
   ix2471 : mux21_ni port map ( Y=>ordered_img_data_11_4, A0=>img_data_13_4, 
      A1=>img_data_3_4, S0=>nx1375);
   ix2479 : mux21_ni port map ( Y=>ordered_img_data_11_5, A0=>img_data_13_5, 
      A1=>img_data_3_5, S0=>nx1375);
   ix2487 : mux21_ni port map ( Y=>ordered_img_data_11_6, A0=>img_data_13_6, 
      A1=>img_data_3_6, S0=>nx1377);
   ix2503 : mux21_ni port map ( Y=>ordered_img_data_11_8, A0=>img_data_13_8, 
      A1=>img_data_3_8, S0=>nx1377);
   ix2511 : mux21_ni port map ( Y=>ordered_img_data_11_9, A0=>img_data_13_9, 
      A1=>img_data_3_9, S0=>nx1377);
   ix2519 : mux21_ni port map ( Y=>ordered_img_data_11_10, A0=>
      img_data_13_10, A1=>img_data_3_10, S0=>nx1377);
   ix2527 : mux21_ni port map ( Y=>ordered_img_data_11_11, A0=>
      img_data_13_11, A1=>img_data_3_11, S0=>nx1377);
   ix2535 : mux21_ni port map ( Y=>ordered_img_data_11_12, A0=>
      img_data_13_12, A1=>img_data_3_12, S0=>nx1377);
   ix2543 : mux21_ni port map ( Y=>ordered_img_data_11_13, A0=>
      img_data_13_13, A1=>img_data_3_13, S0=>nx1377);
   ix2551 : mux21_ni port map ( Y=>ordered_img_data_11_14, A0=>
      img_data_13_14, A1=>img_data_3_14, S0=>nx1379);
   ix2559 : mux21_ni port map ( Y=>ordered_img_data_11_15_EXMPLR, A0=>
      img_data_13_31, A1=>img_data_3_31, S0=>nx1379);
   ix2695 : mux21_ni port map ( Y=>ordered_img_data_10_0, A0=>img_data_8_0, 
      A1=>img_data_2_0, S0=>nx1379);
   ix2711 : mux21_ni port map ( Y=>ordered_img_data_10_2, A0=>img_data_8_2, 
      A1=>img_data_2_2, S0=>nx1379);
   ix2719 : mux21_ni port map ( Y=>ordered_img_data_10_3, A0=>img_data_8_3, 
      A1=>img_data_2_3, S0=>nx1379);
   ix2727 : mux21_ni port map ( Y=>ordered_img_data_10_4, A0=>img_data_8_4, 
      A1=>img_data_2_4, S0=>nx1379);
   ix2735 : mux21_ni port map ( Y=>ordered_img_data_10_5, A0=>img_data_8_5, 
      A1=>img_data_2_5, S0=>nx1379);
   ix2743 : mux21_ni port map ( Y=>ordered_img_data_10_6, A0=>img_data_8_6, 
      A1=>img_data_2_6, S0=>nx1381);
   ix2759 : mux21_ni port map ( Y=>ordered_img_data_10_8, A0=>img_data_8_8, 
      A1=>img_data_2_8, S0=>nx1381);
   ix2767 : mux21_ni port map ( Y=>ordered_img_data_10_9, A0=>img_data_8_9, 
      A1=>img_data_2_9, S0=>nx1381);
   ix2775 : mux21_ni port map ( Y=>ordered_img_data_10_10, A0=>img_data_8_10, 
      A1=>img_data_2_10, S0=>nx1381);
   ix2783 : mux21_ni port map ( Y=>ordered_img_data_10_11, A0=>img_data_8_11, 
      A1=>img_data_2_11, S0=>nx1381);
   ix2791 : mux21_ni port map ( Y=>ordered_img_data_10_12, A0=>img_data_8_12, 
      A1=>img_data_2_12, S0=>nx1381);
   ix2799 : mux21_ni port map ( Y=>ordered_img_data_10_13, A0=>img_data_8_13, 
      A1=>img_data_2_13, S0=>nx1381);
   ix2807 : mux21_ni port map ( Y=>ordered_img_data_10_14, A0=>img_data_8_14, 
      A1=>img_data_2_14, S0=>nx1383);
   ix2815 : mux21_ni port map ( Y=>ordered_img_data_10_15_EXMPLR, A0=>
      img_data_8_31, A1=>img_data_2_31, S0=>nx1383);
   ix2959 : mux21_ni port map ( Y=>ordered_img_data_9_1, A0=>img_data_3_1, 
      A1=>img_data_1_1, S0=>nx1383);
   ix2967 : mux21_ni port map ( Y=>ordered_img_data_9_2, A0=>img_data_3_2, 
      A1=>img_data_1_2, S0=>nx1383);
   ix2975 : mux21_ni port map ( Y=>ordered_img_data_9_3, A0=>img_data_3_3, 
      A1=>img_data_1_3, S0=>nx1383);
   ix2983 : mux21_ni port map ( Y=>ordered_img_data_9_4, A0=>img_data_3_4, 
      A1=>img_data_1_4, S0=>nx1383);
   ix2991 : mux21_ni port map ( Y=>ordered_img_data_9_5, A0=>img_data_3_5, 
      A1=>img_data_1_5, S0=>nx1383);
   ix2999 : mux21_ni port map ( Y=>ordered_img_data_9_6, A0=>img_data_3_6, 
      A1=>img_data_1_6, S0=>nx1385);
   ix3015 : mux21_ni port map ( Y=>ordered_img_data_9_8, A0=>img_data_3_8, 
      A1=>img_data_1_8, S0=>nx1385);
   ix3023 : mux21_ni port map ( Y=>ordered_img_data_9_9, A0=>img_data_3_9, 
      A1=>img_data_1_9, S0=>nx1385);
   ix3031 : mux21_ni port map ( Y=>ordered_img_data_9_10, A0=>img_data_3_10, 
      A1=>img_data_1_10, S0=>nx1315);
   ix3039 : mux21_ni port map ( Y=>ordered_img_data_9_11, A0=>img_data_3_11, 
      A1=>img_data_1_11, S0=>nx1315);
   ix3047 : mux21_ni port map ( Y=>ordered_img_data_9_12, A0=>img_data_3_12, 
      A1=>img_data_1_12, S0=>nx1315);
   ix3055 : mux21_ni port map ( Y=>ordered_img_data_9_13, A0=>img_data_3_13, 
      A1=>img_data_1_13, S0=>nx1315);
   ix3063 : mux21_ni port map ( Y=>ordered_img_data_9_14, A0=>img_data_3_14, 
      A1=>img_data_1_14, S0=>nx1315);
   ix3071 : mux21_ni port map ( Y=>ordered_img_data_9_15_EXMPLR, A0=>
      img_data_3_31, A1=>img_data_1_31, S0=>nx1315);
   ix1205 : inv02 port map ( Y=>nx1206, A=>nx1317);
   ix1208 : inv02 port map ( Y=>nx1209, A=>nx1317);
   ix1210 : inv02 port map ( Y=>nx1211, A=>nx1317);
   ix1212 : inv02 port map ( Y=>nx1213, A=>nx1317);
   ix1214 : inv02 port map ( Y=>nx1215, A=>nx1317);
   ix1216 : inv02 port map ( Y=>nx1217, A=>nx1317);
   ix1218 : inv02 port map ( Y=>nx1219, A=>nx1317);
   ix1220 : inv02 port map ( Y=>nx1221, A=>nx1319);
   ix1222 : inv02 port map ( Y=>nx1223, A=>nx1319);
   ix1224 : inv02 port map ( Y=>nx1225, A=>nx1319);
   ix1226 : inv02 port map ( Y=>nx1227, A=>nx1319);
   ix1228 : inv02 port map ( Y=>nx1229, A=>nx1319);
   ix1230 : inv02 port map ( Y=>nx1231, A=>nx1319);
   ix1232 : inv02 port map ( Y=>nx1233, A=>nx1319);
   ix1234 : inv02 port map ( Y=>nx1235, A=>nx1321);
   ix1236 : inv02 port map ( Y=>nx1237, A=>nx1321);
   ix1238 : inv02 port map ( Y=>nx1239, A=>nx1321);
   ix1240 : inv02 port map ( Y=>nx1241, A=>nx1321);
   ix1242 : inv02 port map ( Y=>nx1243, A=>nx1321);
   ix1244 : inv02 port map ( Y=>nx1245, A=>nx1321);
   ix1246 : inv02 port map ( Y=>nx1247, A=>nx1321);
   ix1248 : inv02 port map ( Y=>nx1249, A=>nx1323);
   ix1250 : inv02 port map ( Y=>nx1251, A=>nx1323);
   ix1252 : inv02 port map ( Y=>nx1253, A=>nx1323);
   ix1254 : inv02 port map ( Y=>nx1255, A=>nx1323);
   ix1256 : inv02 port map ( Y=>nx1257, A=>nx1323);
   ix1258 : inv02 port map ( Y=>nx1259, A=>nx1323);
   ix1260 : inv02 port map ( Y=>nx1261, A=>nx1323);
   ix1262 : inv02 port map ( Y=>nx1263, A=>nx1325);
   ix1264 : inv02 port map ( Y=>nx1265, A=>nx1325);
   ix1266 : inv02 port map ( Y=>nx1267, A=>nx1325);
   ix1268 : inv02 port map ( Y=>nx1269, A=>nx1325);
   ix1270 : inv02 port map ( Y=>nx1271, A=>nx1325);
   ix1272 : inv02 port map ( Y=>nx1273, A=>nx1325);
   ix1286 : inv02 port map ( Y=>nx1287, A=>nx1345);
   ix1300 : inv02 port map ( Y=>nx1301, A=>nx1345);
   ix1314 : inv02 port map ( Y=>nx1315, A=>nx1331);
   ix1318 : inv02 port map ( Y=>nx1319, A=>filter_size);
   ix1320 : inv02 port map ( Y=>nx1321, A=>nx1385);
   ix1322 : inv02 port map ( Y=>nx1323, A=>nx1385);
   ix1316 : inv02 port map ( Y=>nx1317, A=>nx1385);
   reg_ordered_img_data_14_3 : ao22 port map ( Y=>ordered_img_data_14_3, A0
      =>img_data_14_3, A1=>nx1345, B0=>img_data_8_3, B1=>nx1385);
   reg_ordered_img_data_12_4 : ao22 port map ( Y=>ordered_img_data_12_4, A0
      =>img_data_4_4, A1=>nx1345, B0=>img_data_6_4, B1=>nx1387);
   reg_ordered_img_data_13_3 : ao22 port map ( Y=>ordered_img_data_13_3, A0
      =>img_data_9_3, A1=>nx1345, B0=>img_data_7_3, B1=>nx1387);
   reg_ordered_img_data_13_5 : ao22 port map ( Y=>ordered_img_data_13_5, A0
      =>img_data_9_5, A1=>nx1345, B0=>img_data_7_5, B1=>nx1387);
   reg_ordered_img_data_14_7 : ao22 port map ( Y=>ordered_img_data_14_7, A0
      =>img_data_14_7, A1=>nx1345, B0=>img_data_8_7, B1=>nx1387);
   reg_ordered_img_data_12_0 : ao22 port map ( Y=>ordered_img_data_12_0, A0
      =>img_data_4_0, A1=>nx1346, B0=>img_data_6_0, B1=>nx1387);
   reg_ordered_img_data_15_7 : ao22 port map ( Y=>ordered_img_data_15_7, A0
      =>img_data_15_7, A1=>nx1346, B0=>img_data_11_7, B1=>nx1387);
   reg_ordered_img_data_11_2 : ao22 port map ( Y=>ordered_img_data_11_2, A0
      =>img_data_13_2, A1=>nx1346, B0=>img_data_3_2, B1=>nx1387);
   reg_ordered_img_data_15_0 : ao22 port map ( Y=>ordered_img_data_15_0, A0
      =>img_data_15_0, A1=>nx1346, B0=>img_data_11_0, B1=>nx1389);
   reg_ordered_img_data_16_7 : ao22 port map ( Y=>ordered_img_data_16_7, A0
      =>img_data_16_7, A1=>nx1346, B0=>img_data_12_7, B1=>nx1389);
   reg_ordered_img_data_17_5 : ao22 port map ( Y=>ordered_img_data_17_5, A0
      =>img_data_17_5, A1=>nx1346, B0=>img_data_13_5, B1=>nx1389);
   reg_nx1317_XX0_XREP32 : inv01 port map ( Y=>nx1317_XX0_XREP32, A=>nx1389
   );
   reg_ordered_img_data_16_1 : ao22 port map ( Y=>ordered_img_data_16_1, A0
      =>img_data_16_1, A1=>nx1346, B0=>img_data_12_1, B1=>nx1389);
   reg_nx1325 : inv02 port map ( Y=>nx1325, A=>nx1391);
   reg_ordered_img_data_17_0 : ao22 port map ( Y=>ordered_img_data_17_0, A0
      =>img_data_17_0, A1=>nx1325, B0=>img_data_13_0, B1=>nx1389);
   reg_ordered_img_data_9_7 : ao22 port map ( Y=>ordered_img_data_9_7, A0=>
      img_data_3_7, A1=>nx1331, B0=>img_data_1_7, B1=>nx1389);
   reg_ordered_img_data_10_1 : ao22 port map ( Y=>ordered_img_data_10_1, A0
      =>img_data_8_1, A1=>nx1331, B0=>img_data_2_1, B1=>nx1391);
   reg_ordered_img_data_10_7 : ao22 port map ( Y=>ordered_img_data_10_7, A0
      =>img_data_8_7, A1=>nx1331, B0=>img_data_2_7, B1=>nx1391);
   reg_ordered_img_data_11_7 : ao22 port map ( Y=>ordered_img_data_11_7, A0
      =>img_data_13_7, A1=>nx1331, B0=>img_data_3_7, B1=>nx1391);
   reg_nx1331 : inv01 port map ( Y=>nx1331, A=>nx1391);
   reg_ordered_img_data_9_0 : ao22 port map ( Y=>ordered_img_data_9_0, A0=>
      img_data_3_0, A1=>nx1331, B0=>img_data_1_0, B1=>nx1391);
   ix1347 : buf16 port map ( Y=>nx1345, A=>nx1317_XX0_XREP32);
   ix1348 : buf16 port map ( Y=>nx1346, A=>nx1317_XX0_XREP32);
   ix1353 : inv02 port map ( Y=>nx1354, A=>nx1319);
   ix1355 : inv02 port map ( Y=>nx1356, A=>nx1319);
   ix1357 : inv02 port map ( Y=>nx1358, A=>nx1319);
   ix1360 : inv02 port map ( Y=>nx1361, A=>nx1319);
   ix1362 : inv02 port map ( Y=>nx1363, A=>nx1319);
   ix1364 : inv02 port map ( Y=>nx1365, A=>nx1319);
   ix1366 : inv02 port map ( Y=>nx1367, A=>nx1319);
   ix1368 : inv02 port map ( Y=>nx1369, A=>nx1319);
   ix1370 : inv02 port map ( Y=>nx1371, A=>nx1319);
   ix1372 : inv02 port map ( Y=>nx1373, A=>nx1319);
   ix1374 : inv02 port map ( Y=>nx1375, A=>nx1319);
   ix1376 : inv02 port map ( Y=>nx1377, A=>nx1319);
   ix1378 : inv02 port map ( Y=>nx1379, A=>nx1319);
   ix1380 : inv02 port map ( Y=>nx1381, A=>nx1319);
   ix1382 : inv02 port map ( Y=>nx1383, A=>nx1319);
   ix1384 : inv02 port map ( Y=>nx1385, A=>nx1319);
   ix1386 : inv02 port map ( Y=>nx1387, A=>nx1319);
   ix1388 : inv02 port map ( Y=>nx1389, A=>nx1319);
   ix1390 : inv02 port map ( Y=>nx1391, A=>nx1319);
end Structural_unfold_3247_0 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity NAdder_32 is
   port (
      a : IN std_logic_vector (31 DOWNTO 0) ;
      b : IN std_logic_vector (31 DOWNTO 0) ;
      cin : IN std_logic ;
      s : OUT std_logic_vector (31 DOWNTO 0) ;
      cout : OUT std_logic) ;
end NAdder_32 ;

architecture DataFlow_unfold_2448 of NAdder_32 is
   signal nx2, nx16, nx18, nx32, nx34, nx48, nx50, nx64, nx66, nx80, nx82, 
      nx96, nx98, nx112, nx114, nx128, nx130, nx144, nx146, nx160, nx162, 
      nx176, nx178, nx210, nx224, nx226, nx240, nx153, nx155, nx159, nx163, 
      nx169, nx171, nx175, nx179, nx185, nx187, nx191, nx195, nx201, nx203, 
      nx207, nx211, nx217, nx219, nx223, nx227, nx233, nx235, nx239, nx243, 
      nx249, nx251, nx255, nx259, nx265, nx267, nx271, nx275, nx281, nx283, 
      nx287, nx291, nx297, nx299, nx303, nx307, nx313, nx315, nx318, nx321, 
      nx325, nx327, nx339, nx345, nx349, nx354, nx357, nx361, nx363, nx366, 
      nx369, nx373, nx375, nx385, nx386, nx387, nx388, nx208, nx389, nx390, 
      nx391, nx392, nx393, nx394, nx395, nx351, nx342, nx192, nx330, nx396, 
      nx333: std_logic ;

begin
   ix73 : fake_gnd port map ( Y=>cout);
   ix311 : xor2 port map ( Y=>s(0), A0=>b(0), A1=>a(0));
   ix305 : xor2 port map ( Y=>s(1), A0=>nx153, A1=>nx155);
   ix154 : nand02 port map ( Y=>nx153, A0=>b(0), A1=>a(0));
   ix156 : xnor2 port map ( Y=>nx155, A0=>a(1), A1=>b(1));
   ix303 : xor2 port map ( Y=>s(2), A0=>nx159, A1=>nx163);
   ix160 : aoi32 port map ( Y=>nx159, A0=>b(0), A1=>a(0), A2=>nx2, B0=>b(1), 
      B1=>a(1));
   ix164 : xnor2 port map ( Y=>nx163, A0=>a(2), A1=>b(2));
   ix301 : xnor2 port map ( Y=>s(3), A0=>nx16, A1=>nx171);
   ix17 : oai21 port map ( Y=>nx16, A0=>nx159, A1=>nx163, B0=>nx169);
   ix170 : nand02 port map ( Y=>nx169, A0=>b(2), A1=>a(2));
   ix172 : xnor2 port map ( Y=>nx171, A0=>a(3), A1=>b(3));
   ix299 : xor2 port map ( Y=>s(4), A0=>nx175, A1=>nx179);
   ix176 : aoi22 port map ( Y=>nx175, A0=>b(3), A1=>a(3), B0=>nx16, B1=>nx18
   );
   ix180 : xnor2 port map ( Y=>nx179, A0=>a(4), A1=>b(4));
   ix297 : xnor2 port map ( Y=>s(5), A0=>nx32, A1=>nx187);
   ix33 : oai21 port map ( Y=>nx32, A0=>nx175, A1=>nx179, B0=>nx185);
   ix186 : nand02 port map ( Y=>nx185, A0=>b(4), A1=>a(4));
   ix188 : xnor2 port map ( Y=>nx187, A0=>a(5), A1=>b(5));
   ix295 : xor2 port map ( Y=>s(6), A0=>nx191, A1=>nx195);
   ix192 : aoi22 port map ( Y=>nx191, A0=>b(5), A1=>a(5), B0=>nx32, B1=>nx34
   );
   ix196 : xnor2 port map ( Y=>nx195, A0=>a(6), A1=>b(6));
   ix293 : xnor2 port map ( Y=>s(7), A0=>nx48, A1=>nx203);
   ix49 : oai21 port map ( Y=>nx48, A0=>nx191, A1=>nx195, B0=>nx201);
   ix202 : nand02 port map ( Y=>nx201, A0=>b(6), A1=>a(6));
   ix204 : xnor2 port map ( Y=>nx203, A0=>a(7), A1=>b(7));
   ix291 : xor2 port map ( Y=>s(8), A0=>nx207, A1=>nx211);
   ix208 : aoi22 port map ( Y=>nx207, A0=>b(7), A1=>a(7), B0=>nx48, B1=>nx50
   );
   ix212 : xnor2 port map ( Y=>nx211, A0=>a(8), A1=>b(8));
   ix289 : xnor2 port map ( Y=>s(9), A0=>nx64, A1=>nx219);
   ix65 : oai21 port map ( Y=>nx64, A0=>nx207, A1=>nx211, B0=>nx217);
   ix218 : nand02 port map ( Y=>nx217, A0=>b(8), A1=>a(8));
   ix220 : xnor2 port map ( Y=>nx219, A0=>a(9), A1=>b(9));
   ix287 : xor2 port map ( Y=>s(10), A0=>nx223, A1=>nx227);
   ix224 : aoi22 port map ( Y=>nx223, A0=>b(9), A1=>a(9), B0=>nx64, B1=>nx66
   );
   ix228 : xnor2 port map ( Y=>nx227, A0=>a(10), A1=>b(10));
   ix285 : xnor2 port map ( Y=>s(11), A0=>nx80, A1=>nx235);
   ix81 : oai21 port map ( Y=>nx80, A0=>nx223, A1=>nx227, B0=>nx233);
   ix234 : nand02 port map ( Y=>nx233, A0=>b(10), A1=>a(10));
   ix236 : xnor2 port map ( Y=>nx235, A0=>a(11), A1=>b(11));
   ix283 : xor2 port map ( Y=>s(12), A0=>nx239, A1=>nx243);
   ix240 : aoi22 port map ( Y=>nx239, A0=>b(11), A1=>a(11), B0=>nx80, B1=>
      nx82);
   ix244 : xnor2 port map ( Y=>nx243, A0=>a(12), A1=>b(12));
   ix281 : xnor2 port map ( Y=>s(13), A0=>nx96, A1=>nx251);
   ix97 : oai21 port map ( Y=>nx96, A0=>nx239, A1=>nx243, B0=>nx249);
   ix250 : nand02 port map ( Y=>nx249, A0=>b(12), A1=>a(12));
   ix252 : xnor2 port map ( Y=>nx251, A0=>a(13), A1=>b(13));
   ix279 : xor2 port map ( Y=>s(14), A0=>nx255, A1=>nx259);
   ix256 : aoi22 port map ( Y=>nx255, A0=>b(13), A1=>a(13), B0=>nx96, B1=>
      nx98);
   ix260 : xnor2 port map ( Y=>nx259, A0=>a(14), A1=>b(14));
   ix277 : xnor2 port map ( Y=>s(15), A0=>nx112, A1=>nx267);
   ix113 : oai21 port map ( Y=>nx112, A0=>nx255, A1=>nx259, B0=>nx265);
   ix266 : nand02 port map ( Y=>nx265, A0=>b(14), A1=>a(14));
   ix268 : xnor2 port map ( Y=>nx267, A0=>a(15), A1=>b(15));
   ix275 : xor2 port map ( Y=>s(16), A0=>nx271, A1=>nx275);
   ix272 : aoi22 port map ( Y=>nx271, A0=>b(15), A1=>a(15), B0=>nx112, B1=>
      nx114);
   ix276 : xnor2 port map ( Y=>nx275, A0=>a(16), A1=>b(16));
   ix273 : xnor2 port map ( Y=>s(17), A0=>nx128, A1=>nx283);
   ix129 : oai21 port map ( Y=>nx128, A0=>nx271, A1=>nx275, B0=>nx281);
   ix282 : nand02 port map ( Y=>nx281, A0=>b(16), A1=>a(16));
   ix284 : xnor2 port map ( Y=>nx283, A0=>a(17), A1=>b(17));
   ix271 : xor2 port map ( Y=>s(18), A0=>nx287, A1=>nx291);
   ix288 : aoi22 port map ( Y=>nx287, A0=>b(17), A1=>a(17), B0=>nx128, B1=>
      nx130);
   ix292 : xnor2 port map ( Y=>nx291, A0=>a(18), A1=>b(18));
   ix269 : xnor2 port map ( Y=>s(19), A0=>nx144, A1=>nx299);
   ix145 : oai21 port map ( Y=>nx144, A0=>nx287, A1=>nx291, B0=>nx297);
   ix298 : nand02 port map ( Y=>nx297, A0=>b(18), A1=>a(18));
   ix300 : xnor2 port map ( Y=>nx299, A0=>a(19), A1=>b(19));
   ix267 : xor2 port map ( Y=>s(20), A0=>nx303, A1=>nx307);
   ix304 : aoi22 port map ( Y=>nx303, A0=>b(19), A1=>a(19), B0=>nx144, B1=>
      nx146);
   ix308 : xnor2 port map ( Y=>nx307, A0=>a(20), A1=>b(20));
   ix265 : xnor2 port map ( Y=>s(21), A0=>nx160, A1=>nx315);
   ix161 : oai21 port map ( Y=>nx160, A0=>nx303, A1=>nx307, B0=>nx313);
   ix314 : nand02 port map ( Y=>nx313, A0=>b(20), A1=>a(20));
   ix316 : xnor2 port map ( Y=>nx315, A0=>a(21), A1=>b(21));
   ix263 : xor2 port map ( Y=>s(22), A0=>nx318, A1=>nx321);
   ix319 : aoi22 port map ( Y=>nx318, A0=>b(21), A1=>a(21), B0=>nx160, B1=>
      nx162);
   ix322 : xnor2 port map ( Y=>nx321, A0=>a(22), A1=>b(22));
   ix261 : xnor2 port map ( Y=>s(23), A0=>nx176, A1=>nx327);
   ix177 : oai21 port map ( Y=>nx176, A0=>nx318, A1=>nx321, B0=>nx325);
   ix326 : nand02 port map ( Y=>nx325, A0=>b(22), A1=>a(22));
   ix328 : xnor2 port map ( Y=>nx327, A0=>a(23), A1=>b(23));
   ix259 : xor2 port map ( Y=>s(24), A0=>nx330, A1=>nx333);
   ix257 : xnor2 port map ( Y=>s(25), A0=>nx192, A1=>nx339);
   ix340 : xnor2 port map ( Y=>nx339, A0=>a(25), A1=>b(25));
   ix255 : xor2 port map ( Y=>s(26), A0=>nx342, A1=>nx345);
   ix346 : xnor2 port map ( Y=>nx345, A0=>a(26), A1=>b(26));
   ix350 : nand02 port map ( Y=>nx349, A0=>b(26), A1=>a(26));
   ix251 : xor2 port map ( Y=>s(28), A0=>nx354, A1=>nx357);
   ix355 : aoi22 port map ( Y=>nx354, A0=>b(27), A1=>a(27), B0=>nx395, B1=>
      nx210);
   ix358 : xnor2 port map ( Y=>nx357, A0=>a(28), A1=>b(28));
   ix249 : xnor2 port map ( Y=>s(29), A0=>nx224, A1=>nx363);
   ix225 : oai21 port map ( Y=>nx224, A0=>nx354, A1=>nx357, B0=>nx361);
   ix362 : nand02 port map ( Y=>nx361, A0=>b(28), A1=>a(28));
   ix364 : xnor2 port map ( Y=>nx363, A0=>a(29), A1=>b(29));
   ix247 : xor2 port map ( Y=>s(30), A0=>nx366, A1=>nx369);
   ix367 : aoi22 port map ( Y=>nx366, A0=>b(29), A1=>a(29), B0=>nx224, B1=>
      nx226);
   ix370 : xnor2 port map ( Y=>nx369, A0=>a(30), A1=>b(30));
   ix245 : xnor2 port map ( Y=>s(31), A0=>nx240, A1=>nx375);
   ix241 : oai21 port map ( Y=>nx240, A0=>nx366, A1=>nx369, B0=>nx373);
   ix374 : nand02 port map ( Y=>nx373, A0=>b(30), A1=>a(30));
   ix376 : xnor2 port map ( Y=>nx375, A0=>a(31), A1=>b(31));
   ix227 : inv01 port map ( Y=>nx226, A=>nx363);
   ix211 : inv01 port map ( Y=>nx210, A=>nx351);
   ix179 : inv01 port map ( Y=>nx178, A=>nx327);
   ix163 : inv01 port map ( Y=>nx162, A=>nx315);
   ix147 : inv01 port map ( Y=>nx146, A=>nx299);
   ix131 : inv01 port map ( Y=>nx130, A=>nx283);
   ix115 : inv01 port map ( Y=>nx114, A=>nx267);
   ix99 : inv01 port map ( Y=>nx98, A=>nx251);
   ix83 : inv01 port map ( Y=>nx82, A=>nx235);
   ix67 : inv01 port map ( Y=>nx66, A=>nx219);
   ix51 : inv01 port map ( Y=>nx50, A=>nx203);
   ix35 : inv01 port map ( Y=>nx34, A=>nx187);
   ix19 : inv01 port map ( Y=>nx18, A=>nx171);
   ix3 : inv01 port map ( Y=>nx2, A=>nx155);
   ix397 : or02 port map ( Y=>nx385, A0=>a(24), A1=>b(24));
   ix398 : and02 port map ( Y=>nx386, A0=>b(23), A1=>a(23));
   ix399 : aoi322 port map ( Y=>nx387, A0=>nx176, A1=>nx178, A2=>nx385, B0=>
      nx385, B1=>nx386, C0=>a(24), C1=>b(24));
   ix400 : nand02_2x port map ( Y=>nx388, A0=>b(25), A1=>a(25));
   reg_nx208 : oai321 port map ( Y=>nx208, A0=>nx387, A1=>nx345, A2=>nx339, 
      B0=>nx345, B1=>nx388, C0=>nx349);
   ix401 : inv02 port map ( Y=>nx389, A=>nx208);
   ix402 : inv02 port map ( Y=>nx390, A=>a(27));
   ix403 : inv02 port map ( Y=>nx391, A=>b(27));
   ix404 : aoi22 port map ( Y=>nx392, A0=>a(27), A1=>b(27), B0=>nx390, B1=>
      nx391);
   ix405 : oai22 port map ( Y=>nx393, A0=>nx391, A1=>a(27), B0=>nx390, B1=>
      b(27));
   ix406 : nand02_2x port map ( Y=>nx394, A0=>nx393, A1=>nx389);
   reg_s_27 : oai21 port map ( Y=>s(27), A0=>nx389, A1=>nx392, B0=>nx394);
   ix407 : inv02 port map ( Y=>nx395, A=>nx389);
   reg_nx351 : oai22 port map ( Y=>nx351, A0=>nx390, A1=>nx391, B0=>a(27), 
      B1=>b(27));
   reg_nx342 : ao22 port map ( Y=>nx342, A0=>nx388, A1=>nx387, B0=>nx339, B1
      =>nx388);
   reg_nx192 : inv01 port map ( Y=>nx192, A=>nx387);
   reg_nx330 : oai22 port map ( Y=>nx330, A0=>nx386, A1=>nx176, B0=>nx386, 
      B1=>nx178);
   ix408 : nor02_2x port map ( Y=>nx396, A0=>a(24), A1=>b(24));
   reg_nx333 : ao21 port map ( Y=>nx333, A0=>a(24), A1=>b(24), B0=>nx396);

end DataFlow_unfold_2448 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity MergeLayer is
   port (
      d_arr_0_31 : OUT std_logic ;
      d_arr_0_30 : OUT std_logic ;
      d_arr_0_29 : OUT std_logic ;
      d_arr_0_28 : OUT std_logic ;
      d_arr_0_27 : OUT std_logic ;
      d_arr_0_26 : OUT std_logic ;
      d_arr_0_25 : OUT std_logic ;
      d_arr_0_24 : OUT std_logic ;
      d_arr_0_23 : OUT std_logic ;
      d_arr_0_22 : OUT std_logic ;
      d_arr_0_21 : OUT std_logic ;
      d_arr_0_20 : OUT std_logic ;
      d_arr_0_19 : OUT std_logic ;
      d_arr_0_18 : OUT std_logic ;
      d_arr_0_17 : OUT std_logic ;
      d_arr_0_16 : OUT std_logic ;
      d_arr_0_15 : OUT std_logic ;
      d_arr_0_14 : OUT std_logic ;
      d_arr_0_13 : OUT std_logic ;
      d_arr_0_12 : OUT std_logic ;
      d_arr_0_11 : OUT std_logic ;
      d_arr_0_10 : OUT std_logic ;
      d_arr_0_9 : OUT std_logic ;
      d_arr_0_8 : OUT std_logic ;
      d_arr_0_7 : OUT std_logic ;
      d_arr_0_6 : OUT std_logic ;
      d_arr_0_5 : OUT std_logic ;
      d_arr_0_4 : OUT std_logic ;
      d_arr_0_3 : OUT std_logic ;
      d_arr_0_2 : OUT std_logic ;
      d_arr_0_1 : OUT std_logic ;
      d_arr_0_0 : OUT std_logic ;
      d_arr_1_31 : OUT std_logic ;
      d_arr_1_30 : OUT std_logic ;
      d_arr_1_29 : OUT std_logic ;
      d_arr_1_28 : OUT std_logic ;
      d_arr_1_27 : OUT std_logic ;
      d_arr_1_26 : OUT std_logic ;
      d_arr_1_25 : OUT std_logic ;
      d_arr_1_24 : OUT std_logic ;
      d_arr_1_23 : OUT std_logic ;
      d_arr_1_22 : OUT std_logic ;
      d_arr_1_21 : OUT std_logic ;
      d_arr_1_20 : OUT std_logic ;
      d_arr_1_19 : OUT std_logic ;
      d_arr_1_18 : OUT std_logic ;
      d_arr_1_17 : OUT std_logic ;
      d_arr_1_16 : OUT std_logic ;
      d_arr_1_15 : OUT std_logic ;
      d_arr_1_14 : OUT std_logic ;
      d_arr_1_13 : OUT std_logic ;
      d_arr_1_12 : OUT std_logic ;
      d_arr_1_11 : OUT std_logic ;
      d_arr_1_10 : OUT std_logic ;
      d_arr_1_9 : OUT std_logic ;
      d_arr_1_8 : OUT std_logic ;
      d_arr_1_7 : OUT std_logic ;
      d_arr_1_6 : OUT std_logic ;
      d_arr_1_5 : OUT std_logic ;
      d_arr_1_4 : OUT std_logic ;
      d_arr_1_3 : OUT std_logic ;
      d_arr_1_2 : OUT std_logic ;
      d_arr_1_1 : OUT std_logic ;
      d_arr_1_0 : OUT std_logic ;
      d_arr_2_31 : OUT std_logic ;
      d_arr_2_30 : OUT std_logic ;
      d_arr_2_29 : OUT std_logic ;
      d_arr_2_28 : OUT std_logic ;
      d_arr_2_27 : OUT std_logic ;
      d_arr_2_26 : OUT std_logic ;
      d_arr_2_25 : OUT std_logic ;
      d_arr_2_24 : OUT std_logic ;
      d_arr_2_23 : OUT std_logic ;
      d_arr_2_22 : OUT std_logic ;
      d_arr_2_21 : OUT std_logic ;
      d_arr_2_20 : OUT std_logic ;
      d_arr_2_19 : OUT std_logic ;
      d_arr_2_18 : OUT std_logic ;
      d_arr_2_17 : OUT std_logic ;
      d_arr_2_16 : OUT std_logic ;
      d_arr_2_15 : OUT std_logic ;
      d_arr_2_14 : OUT std_logic ;
      d_arr_2_13 : OUT std_logic ;
      d_arr_2_12 : OUT std_logic ;
      d_arr_2_11 : OUT std_logic ;
      d_arr_2_10 : OUT std_logic ;
      d_arr_2_9 : OUT std_logic ;
      d_arr_2_8 : OUT std_logic ;
      d_arr_2_7 : OUT std_logic ;
      d_arr_2_6 : OUT std_logic ;
      d_arr_2_5 : OUT std_logic ;
      d_arr_2_4 : OUT std_logic ;
      d_arr_2_3 : OUT std_logic ;
      d_arr_2_2 : OUT std_logic ;
      d_arr_2_1 : OUT std_logic ;
      d_arr_2_0 : OUT std_logic ;
      d_arr_3_31 : OUT std_logic ;
      d_arr_3_30 : OUT std_logic ;
      d_arr_3_29 : OUT std_logic ;
      d_arr_3_28 : OUT std_logic ;
      d_arr_3_27 : OUT std_logic ;
      d_arr_3_26 : OUT std_logic ;
      d_arr_3_25 : OUT std_logic ;
      d_arr_3_24 : OUT std_logic ;
      d_arr_3_23 : OUT std_logic ;
      d_arr_3_22 : OUT std_logic ;
      d_arr_3_21 : OUT std_logic ;
      d_arr_3_20 : OUT std_logic ;
      d_arr_3_19 : OUT std_logic ;
      d_arr_3_18 : OUT std_logic ;
      d_arr_3_17 : OUT std_logic ;
      d_arr_3_16 : OUT std_logic ;
      d_arr_3_15 : OUT std_logic ;
      d_arr_3_14 : OUT std_logic ;
      d_arr_3_13 : OUT std_logic ;
      d_arr_3_12 : OUT std_logic ;
      d_arr_3_11 : OUT std_logic ;
      d_arr_3_10 : OUT std_logic ;
      d_arr_3_9 : OUT std_logic ;
      d_arr_3_8 : OUT std_logic ;
      d_arr_3_7 : OUT std_logic ;
      d_arr_3_6 : OUT std_logic ;
      d_arr_3_5 : OUT std_logic ;
      d_arr_3_4 : OUT std_logic ;
      d_arr_3_3 : OUT std_logic ;
      d_arr_3_2 : OUT std_logic ;
      d_arr_3_1 : OUT std_logic ;
      d_arr_3_0 : OUT std_logic ;
      d_arr_4_31 : OUT std_logic ;
      d_arr_4_30 : OUT std_logic ;
      d_arr_4_29 : OUT std_logic ;
      d_arr_4_28 : OUT std_logic ;
      d_arr_4_27 : OUT std_logic ;
      d_arr_4_26 : OUT std_logic ;
      d_arr_4_25 : OUT std_logic ;
      d_arr_4_24 : OUT std_logic ;
      d_arr_4_23 : OUT std_logic ;
      d_arr_4_22 : OUT std_logic ;
      d_arr_4_21 : OUT std_logic ;
      d_arr_4_20 : OUT std_logic ;
      d_arr_4_19 : OUT std_logic ;
      d_arr_4_18 : OUT std_logic ;
      d_arr_4_17 : OUT std_logic ;
      d_arr_4_16 : OUT std_logic ;
      d_arr_4_15 : OUT std_logic ;
      d_arr_4_14 : OUT std_logic ;
      d_arr_4_13 : OUT std_logic ;
      d_arr_4_12 : OUT std_logic ;
      d_arr_4_11 : OUT std_logic ;
      d_arr_4_10 : OUT std_logic ;
      d_arr_4_9 : OUT std_logic ;
      d_arr_4_8 : OUT std_logic ;
      d_arr_4_7 : OUT std_logic ;
      d_arr_4_6 : OUT std_logic ;
      d_arr_4_5 : OUT std_logic ;
      d_arr_4_4 : OUT std_logic ;
      d_arr_4_3 : OUT std_logic ;
      d_arr_4_2 : OUT std_logic ;
      d_arr_4_1 : OUT std_logic ;
      d_arr_4_0 : OUT std_logic ;
      d_arr_5_31 : OUT std_logic ;
      d_arr_5_30 : OUT std_logic ;
      d_arr_5_29 : OUT std_logic ;
      d_arr_5_28 : OUT std_logic ;
      d_arr_5_27 : OUT std_logic ;
      d_arr_5_26 : OUT std_logic ;
      d_arr_5_25 : OUT std_logic ;
      d_arr_5_24 : OUT std_logic ;
      d_arr_5_23 : OUT std_logic ;
      d_arr_5_22 : OUT std_logic ;
      d_arr_5_21 : OUT std_logic ;
      d_arr_5_20 : OUT std_logic ;
      d_arr_5_19 : OUT std_logic ;
      d_arr_5_18 : OUT std_logic ;
      d_arr_5_17 : OUT std_logic ;
      d_arr_5_16 : OUT std_logic ;
      d_arr_5_15 : OUT std_logic ;
      d_arr_5_14 : OUT std_logic ;
      d_arr_5_13 : OUT std_logic ;
      d_arr_5_12 : OUT std_logic ;
      d_arr_5_11 : OUT std_logic ;
      d_arr_5_10 : OUT std_logic ;
      d_arr_5_9 : OUT std_logic ;
      d_arr_5_8 : OUT std_logic ;
      d_arr_5_7 : OUT std_logic ;
      d_arr_5_6 : OUT std_logic ;
      d_arr_5_5 : OUT std_logic ;
      d_arr_5_4 : OUT std_logic ;
      d_arr_5_3 : OUT std_logic ;
      d_arr_5_2 : OUT std_logic ;
      d_arr_5_1 : OUT std_logic ;
      d_arr_5_0 : OUT std_logic ;
      d_arr_6_31 : OUT std_logic ;
      d_arr_6_30 : OUT std_logic ;
      d_arr_6_29 : OUT std_logic ;
      d_arr_6_28 : OUT std_logic ;
      d_arr_6_27 : OUT std_logic ;
      d_arr_6_26 : OUT std_logic ;
      d_arr_6_25 : OUT std_logic ;
      d_arr_6_24 : OUT std_logic ;
      d_arr_6_23 : OUT std_logic ;
      d_arr_6_22 : OUT std_logic ;
      d_arr_6_21 : OUT std_logic ;
      d_arr_6_20 : OUT std_logic ;
      d_arr_6_19 : OUT std_logic ;
      d_arr_6_18 : OUT std_logic ;
      d_arr_6_17 : OUT std_logic ;
      d_arr_6_16 : OUT std_logic ;
      d_arr_6_15 : OUT std_logic ;
      d_arr_6_14 : OUT std_logic ;
      d_arr_6_13 : OUT std_logic ;
      d_arr_6_12 : OUT std_logic ;
      d_arr_6_11 : OUT std_logic ;
      d_arr_6_10 : OUT std_logic ;
      d_arr_6_9 : OUT std_logic ;
      d_arr_6_8 : OUT std_logic ;
      d_arr_6_7 : OUT std_logic ;
      d_arr_6_6 : OUT std_logic ;
      d_arr_6_5 : OUT std_logic ;
      d_arr_6_4 : OUT std_logic ;
      d_arr_6_3 : OUT std_logic ;
      d_arr_6_2 : OUT std_logic ;
      d_arr_6_1 : OUT std_logic ;
      d_arr_6_0 : OUT std_logic ;
      d_arr_7_31 : OUT std_logic ;
      d_arr_7_30 : OUT std_logic ;
      d_arr_7_29 : OUT std_logic ;
      d_arr_7_28 : OUT std_logic ;
      d_arr_7_27 : OUT std_logic ;
      d_arr_7_26 : OUT std_logic ;
      d_arr_7_25 : OUT std_logic ;
      d_arr_7_24 : OUT std_logic ;
      d_arr_7_23 : OUT std_logic ;
      d_arr_7_22 : OUT std_logic ;
      d_arr_7_21 : OUT std_logic ;
      d_arr_7_20 : OUT std_logic ;
      d_arr_7_19 : OUT std_logic ;
      d_arr_7_18 : OUT std_logic ;
      d_arr_7_17 : OUT std_logic ;
      d_arr_7_16 : OUT std_logic ;
      d_arr_7_15 : OUT std_logic ;
      d_arr_7_14 : OUT std_logic ;
      d_arr_7_13 : OUT std_logic ;
      d_arr_7_12 : OUT std_logic ;
      d_arr_7_11 : OUT std_logic ;
      d_arr_7_10 : OUT std_logic ;
      d_arr_7_9 : OUT std_logic ;
      d_arr_7_8 : OUT std_logic ;
      d_arr_7_7 : OUT std_logic ;
      d_arr_7_6 : OUT std_logic ;
      d_arr_7_5 : OUT std_logic ;
      d_arr_7_4 : OUT std_logic ;
      d_arr_7_3 : OUT std_logic ;
      d_arr_7_2 : OUT std_logic ;
      d_arr_7_1 : OUT std_logic ;
      d_arr_7_0 : OUT std_logic ;
      d_arr_8_31 : OUT std_logic ;
      d_arr_8_30 : OUT std_logic ;
      d_arr_8_29 : OUT std_logic ;
      d_arr_8_28 : OUT std_logic ;
      d_arr_8_27 : OUT std_logic ;
      d_arr_8_26 : OUT std_logic ;
      d_arr_8_25 : OUT std_logic ;
      d_arr_8_24 : OUT std_logic ;
      d_arr_8_23 : OUT std_logic ;
      d_arr_8_22 : OUT std_logic ;
      d_arr_8_21 : OUT std_logic ;
      d_arr_8_20 : OUT std_logic ;
      d_arr_8_19 : OUT std_logic ;
      d_arr_8_18 : OUT std_logic ;
      d_arr_8_17 : OUT std_logic ;
      d_arr_8_16 : OUT std_logic ;
      d_arr_8_15 : OUT std_logic ;
      d_arr_8_14 : OUT std_logic ;
      d_arr_8_13 : OUT std_logic ;
      d_arr_8_12 : OUT std_logic ;
      d_arr_8_11 : OUT std_logic ;
      d_arr_8_10 : OUT std_logic ;
      d_arr_8_9 : OUT std_logic ;
      d_arr_8_8 : OUT std_logic ;
      d_arr_8_7 : OUT std_logic ;
      d_arr_8_6 : OUT std_logic ;
      d_arr_8_5 : OUT std_logic ;
      d_arr_8_4 : OUT std_logic ;
      d_arr_8_3 : OUT std_logic ;
      d_arr_8_2 : OUT std_logic ;
      d_arr_8_1 : OUT std_logic ;
      d_arr_8_0 : OUT std_logic ;
      d_arr_9_31 : OUT std_logic ;
      d_arr_9_30 : OUT std_logic ;
      d_arr_9_29 : OUT std_logic ;
      d_arr_9_28 : OUT std_logic ;
      d_arr_9_27 : OUT std_logic ;
      d_arr_9_26 : OUT std_logic ;
      d_arr_9_25 : OUT std_logic ;
      d_arr_9_24 : OUT std_logic ;
      d_arr_9_23 : OUT std_logic ;
      d_arr_9_22 : OUT std_logic ;
      d_arr_9_21 : OUT std_logic ;
      d_arr_9_20 : OUT std_logic ;
      d_arr_9_19 : OUT std_logic ;
      d_arr_9_18 : OUT std_logic ;
      d_arr_9_17 : OUT std_logic ;
      d_arr_9_16 : OUT std_logic ;
      d_arr_9_15 : OUT std_logic ;
      d_arr_9_14 : OUT std_logic ;
      d_arr_9_13 : OUT std_logic ;
      d_arr_9_12 : OUT std_logic ;
      d_arr_9_11 : OUT std_logic ;
      d_arr_9_10 : OUT std_logic ;
      d_arr_9_9 : OUT std_logic ;
      d_arr_9_8 : OUT std_logic ;
      d_arr_9_7 : OUT std_logic ;
      d_arr_9_6 : OUT std_logic ;
      d_arr_9_5 : OUT std_logic ;
      d_arr_9_4 : OUT std_logic ;
      d_arr_9_3 : OUT std_logic ;
      d_arr_9_2 : OUT std_logic ;
      d_arr_9_1 : OUT std_logic ;
      d_arr_9_0 : OUT std_logic ;
      d_arr_10_31 : OUT std_logic ;
      d_arr_10_30 : OUT std_logic ;
      d_arr_10_29 : OUT std_logic ;
      d_arr_10_28 : OUT std_logic ;
      d_arr_10_27 : OUT std_logic ;
      d_arr_10_26 : OUT std_logic ;
      d_arr_10_25 : OUT std_logic ;
      d_arr_10_24 : OUT std_logic ;
      d_arr_10_23 : OUT std_logic ;
      d_arr_10_22 : OUT std_logic ;
      d_arr_10_21 : OUT std_logic ;
      d_arr_10_20 : OUT std_logic ;
      d_arr_10_19 : OUT std_logic ;
      d_arr_10_18 : OUT std_logic ;
      d_arr_10_17 : OUT std_logic ;
      d_arr_10_16 : OUT std_logic ;
      d_arr_10_15 : OUT std_logic ;
      d_arr_10_14 : OUT std_logic ;
      d_arr_10_13 : OUT std_logic ;
      d_arr_10_12 : OUT std_logic ;
      d_arr_10_11 : OUT std_logic ;
      d_arr_10_10 : OUT std_logic ;
      d_arr_10_9 : OUT std_logic ;
      d_arr_10_8 : OUT std_logic ;
      d_arr_10_7 : OUT std_logic ;
      d_arr_10_6 : OUT std_logic ;
      d_arr_10_5 : OUT std_logic ;
      d_arr_10_4 : OUT std_logic ;
      d_arr_10_3 : OUT std_logic ;
      d_arr_10_2 : OUT std_logic ;
      d_arr_10_1 : OUT std_logic ;
      d_arr_10_0 : OUT std_logic ;
      d_arr_11_31 : OUT std_logic ;
      d_arr_11_30 : OUT std_logic ;
      d_arr_11_29 : OUT std_logic ;
      d_arr_11_28 : OUT std_logic ;
      d_arr_11_27 : OUT std_logic ;
      d_arr_11_26 : OUT std_logic ;
      d_arr_11_25 : OUT std_logic ;
      d_arr_11_24 : OUT std_logic ;
      d_arr_11_23 : OUT std_logic ;
      d_arr_11_22 : OUT std_logic ;
      d_arr_11_21 : OUT std_logic ;
      d_arr_11_20 : OUT std_logic ;
      d_arr_11_19 : OUT std_logic ;
      d_arr_11_18 : OUT std_logic ;
      d_arr_11_17 : OUT std_logic ;
      d_arr_11_16 : OUT std_logic ;
      d_arr_11_15 : OUT std_logic ;
      d_arr_11_14 : OUT std_logic ;
      d_arr_11_13 : OUT std_logic ;
      d_arr_11_12 : OUT std_logic ;
      d_arr_11_11 : OUT std_logic ;
      d_arr_11_10 : OUT std_logic ;
      d_arr_11_9 : OUT std_logic ;
      d_arr_11_8 : OUT std_logic ;
      d_arr_11_7 : OUT std_logic ;
      d_arr_11_6 : OUT std_logic ;
      d_arr_11_5 : OUT std_logic ;
      d_arr_11_4 : OUT std_logic ;
      d_arr_11_3 : OUT std_logic ;
      d_arr_11_2 : OUT std_logic ;
      d_arr_11_1 : OUT std_logic ;
      d_arr_11_0 : OUT std_logic ;
      d_arr_12_31 : OUT std_logic ;
      d_arr_12_30 : OUT std_logic ;
      d_arr_12_29 : OUT std_logic ;
      d_arr_12_28 : OUT std_logic ;
      d_arr_12_27 : OUT std_logic ;
      d_arr_12_26 : OUT std_logic ;
      d_arr_12_25 : OUT std_logic ;
      d_arr_12_24 : OUT std_logic ;
      d_arr_12_23 : OUT std_logic ;
      d_arr_12_22 : OUT std_logic ;
      d_arr_12_21 : OUT std_logic ;
      d_arr_12_20 : OUT std_logic ;
      d_arr_12_19 : OUT std_logic ;
      d_arr_12_18 : OUT std_logic ;
      d_arr_12_17 : OUT std_logic ;
      d_arr_12_16 : OUT std_logic ;
      d_arr_12_15 : OUT std_logic ;
      d_arr_12_14 : OUT std_logic ;
      d_arr_12_13 : OUT std_logic ;
      d_arr_12_12 : OUT std_logic ;
      d_arr_12_11 : OUT std_logic ;
      d_arr_12_10 : OUT std_logic ;
      d_arr_12_9 : OUT std_logic ;
      d_arr_12_8 : OUT std_logic ;
      d_arr_12_7 : OUT std_logic ;
      d_arr_12_6 : OUT std_logic ;
      d_arr_12_5 : OUT std_logic ;
      d_arr_12_4 : OUT std_logic ;
      d_arr_12_3 : OUT std_logic ;
      d_arr_12_2 : OUT std_logic ;
      d_arr_12_1 : OUT std_logic ;
      d_arr_12_0 : OUT std_logic ;
      d_arr_13_31 : OUT std_logic ;
      d_arr_13_30 : OUT std_logic ;
      d_arr_13_29 : OUT std_logic ;
      d_arr_13_28 : OUT std_logic ;
      d_arr_13_27 : OUT std_logic ;
      d_arr_13_26 : OUT std_logic ;
      d_arr_13_25 : OUT std_logic ;
      d_arr_13_24 : OUT std_logic ;
      d_arr_13_23 : OUT std_logic ;
      d_arr_13_22 : OUT std_logic ;
      d_arr_13_21 : OUT std_logic ;
      d_arr_13_20 : OUT std_logic ;
      d_arr_13_19 : OUT std_logic ;
      d_arr_13_18 : OUT std_logic ;
      d_arr_13_17 : OUT std_logic ;
      d_arr_13_16 : OUT std_logic ;
      d_arr_13_15 : OUT std_logic ;
      d_arr_13_14 : OUT std_logic ;
      d_arr_13_13 : OUT std_logic ;
      d_arr_13_12 : OUT std_logic ;
      d_arr_13_11 : OUT std_logic ;
      d_arr_13_10 : OUT std_logic ;
      d_arr_13_9 : OUT std_logic ;
      d_arr_13_8 : OUT std_logic ;
      d_arr_13_7 : OUT std_logic ;
      d_arr_13_6 : OUT std_logic ;
      d_arr_13_5 : OUT std_logic ;
      d_arr_13_4 : OUT std_logic ;
      d_arr_13_3 : OUT std_logic ;
      d_arr_13_2 : OUT std_logic ;
      d_arr_13_1 : OUT std_logic ;
      d_arr_13_0 : OUT std_logic ;
      d_arr_14_31 : OUT std_logic ;
      d_arr_14_30 : OUT std_logic ;
      d_arr_14_29 : OUT std_logic ;
      d_arr_14_28 : OUT std_logic ;
      d_arr_14_27 : OUT std_logic ;
      d_arr_14_26 : OUT std_logic ;
      d_arr_14_25 : OUT std_logic ;
      d_arr_14_24 : OUT std_logic ;
      d_arr_14_23 : OUT std_logic ;
      d_arr_14_22 : OUT std_logic ;
      d_arr_14_21 : OUT std_logic ;
      d_arr_14_20 : OUT std_logic ;
      d_arr_14_19 : OUT std_logic ;
      d_arr_14_18 : OUT std_logic ;
      d_arr_14_17 : OUT std_logic ;
      d_arr_14_16 : OUT std_logic ;
      d_arr_14_15 : OUT std_logic ;
      d_arr_14_14 : OUT std_logic ;
      d_arr_14_13 : OUT std_logic ;
      d_arr_14_12 : OUT std_logic ;
      d_arr_14_11 : OUT std_logic ;
      d_arr_14_10 : OUT std_logic ;
      d_arr_14_9 : OUT std_logic ;
      d_arr_14_8 : OUT std_logic ;
      d_arr_14_7 : OUT std_logic ;
      d_arr_14_6 : OUT std_logic ;
      d_arr_14_5 : OUT std_logic ;
      d_arr_14_4 : OUT std_logic ;
      d_arr_14_3 : OUT std_logic ;
      d_arr_14_2 : OUT std_logic ;
      d_arr_14_1 : OUT std_logic ;
      d_arr_14_0 : OUT std_logic ;
      d_arr_15_31 : OUT std_logic ;
      d_arr_15_30 : OUT std_logic ;
      d_arr_15_29 : OUT std_logic ;
      d_arr_15_28 : OUT std_logic ;
      d_arr_15_27 : OUT std_logic ;
      d_arr_15_26 : OUT std_logic ;
      d_arr_15_25 : OUT std_logic ;
      d_arr_15_24 : OUT std_logic ;
      d_arr_15_23 : OUT std_logic ;
      d_arr_15_22 : OUT std_logic ;
      d_arr_15_21 : OUT std_logic ;
      d_arr_15_20 : OUT std_logic ;
      d_arr_15_19 : OUT std_logic ;
      d_arr_15_18 : OUT std_logic ;
      d_arr_15_17 : OUT std_logic ;
      d_arr_15_16 : OUT std_logic ;
      d_arr_15_15 : OUT std_logic ;
      d_arr_15_14 : OUT std_logic ;
      d_arr_15_13 : OUT std_logic ;
      d_arr_15_12 : OUT std_logic ;
      d_arr_15_11 : OUT std_logic ;
      d_arr_15_10 : OUT std_logic ;
      d_arr_15_9 : OUT std_logic ;
      d_arr_15_8 : OUT std_logic ;
      d_arr_15_7 : OUT std_logic ;
      d_arr_15_6 : OUT std_logic ;
      d_arr_15_5 : OUT std_logic ;
      d_arr_15_4 : OUT std_logic ;
      d_arr_15_3 : OUT std_logic ;
      d_arr_15_2 : OUT std_logic ;
      d_arr_15_1 : OUT std_logic ;
      d_arr_15_0 : OUT std_logic ;
      d_arr_16_31 : OUT std_logic ;
      d_arr_16_30 : OUT std_logic ;
      d_arr_16_29 : OUT std_logic ;
      d_arr_16_28 : OUT std_logic ;
      d_arr_16_27 : OUT std_logic ;
      d_arr_16_26 : OUT std_logic ;
      d_arr_16_25 : OUT std_logic ;
      d_arr_16_24 : OUT std_logic ;
      d_arr_16_23 : OUT std_logic ;
      d_arr_16_22 : OUT std_logic ;
      d_arr_16_21 : OUT std_logic ;
      d_arr_16_20 : OUT std_logic ;
      d_arr_16_19 : OUT std_logic ;
      d_arr_16_18 : OUT std_logic ;
      d_arr_16_17 : OUT std_logic ;
      d_arr_16_16 : OUT std_logic ;
      d_arr_16_15 : OUT std_logic ;
      d_arr_16_14 : OUT std_logic ;
      d_arr_16_13 : OUT std_logic ;
      d_arr_16_12 : OUT std_logic ;
      d_arr_16_11 : OUT std_logic ;
      d_arr_16_10 : OUT std_logic ;
      d_arr_16_9 : OUT std_logic ;
      d_arr_16_8 : OUT std_logic ;
      d_arr_16_7 : OUT std_logic ;
      d_arr_16_6 : OUT std_logic ;
      d_arr_16_5 : OUT std_logic ;
      d_arr_16_4 : OUT std_logic ;
      d_arr_16_3 : OUT std_logic ;
      d_arr_16_2 : OUT std_logic ;
      d_arr_16_1 : OUT std_logic ;
      d_arr_16_0 : OUT std_logic ;
      d_arr_17_31 : OUT std_logic ;
      d_arr_17_30 : OUT std_logic ;
      d_arr_17_29 : OUT std_logic ;
      d_arr_17_28 : OUT std_logic ;
      d_arr_17_27 : OUT std_logic ;
      d_arr_17_26 : OUT std_logic ;
      d_arr_17_25 : OUT std_logic ;
      d_arr_17_24 : OUT std_logic ;
      d_arr_17_23 : OUT std_logic ;
      d_arr_17_22 : OUT std_logic ;
      d_arr_17_21 : OUT std_logic ;
      d_arr_17_20 : OUT std_logic ;
      d_arr_17_19 : OUT std_logic ;
      d_arr_17_18 : OUT std_logic ;
      d_arr_17_17 : OUT std_logic ;
      d_arr_17_16 : OUT std_logic ;
      d_arr_17_15 : OUT std_logic ;
      d_arr_17_14 : OUT std_logic ;
      d_arr_17_13 : OUT std_logic ;
      d_arr_17_12 : OUT std_logic ;
      d_arr_17_11 : OUT std_logic ;
      d_arr_17_10 : OUT std_logic ;
      d_arr_17_9 : OUT std_logic ;
      d_arr_17_8 : OUT std_logic ;
      d_arr_17_7 : OUT std_logic ;
      d_arr_17_6 : OUT std_logic ;
      d_arr_17_5 : OUT std_logic ;
      d_arr_17_4 : OUT std_logic ;
      d_arr_17_3 : OUT std_logic ;
      d_arr_17_2 : OUT std_logic ;
      d_arr_17_1 : OUT std_logic ;
      d_arr_17_0 : OUT std_logic ;
      d_arr_18_31 : OUT std_logic ;
      d_arr_18_30 : OUT std_logic ;
      d_arr_18_29 : OUT std_logic ;
      d_arr_18_28 : OUT std_logic ;
      d_arr_18_27 : OUT std_logic ;
      d_arr_18_26 : OUT std_logic ;
      d_arr_18_25 : OUT std_logic ;
      d_arr_18_24 : OUT std_logic ;
      d_arr_18_23 : OUT std_logic ;
      d_arr_18_22 : OUT std_logic ;
      d_arr_18_21 : OUT std_logic ;
      d_arr_18_20 : OUT std_logic ;
      d_arr_18_19 : OUT std_logic ;
      d_arr_18_18 : OUT std_logic ;
      d_arr_18_17 : OUT std_logic ;
      d_arr_18_16 : OUT std_logic ;
      d_arr_18_15 : OUT std_logic ;
      d_arr_18_14 : OUT std_logic ;
      d_arr_18_13 : OUT std_logic ;
      d_arr_18_12 : OUT std_logic ;
      d_arr_18_11 : OUT std_logic ;
      d_arr_18_10 : OUT std_logic ;
      d_arr_18_9 : OUT std_logic ;
      d_arr_18_8 : OUT std_logic ;
      d_arr_18_7 : OUT std_logic ;
      d_arr_18_6 : OUT std_logic ;
      d_arr_18_5 : OUT std_logic ;
      d_arr_18_4 : OUT std_logic ;
      d_arr_18_3 : OUT std_logic ;
      d_arr_18_2 : OUT std_logic ;
      d_arr_18_1 : OUT std_logic ;
      d_arr_18_0 : OUT std_logic ;
      d_arr_19_31 : OUT std_logic ;
      d_arr_19_30 : OUT std_logic ;
      d_arr_19_29 : OUT std_logic ;
      d_arr_19_28 : OUT std_logic ;
      d_arr_19_27 : OUT std_logic ;
      d_arr_19_26 : OUT std_logic ;
      d_arr_19_25 : OUT std_logic ;
      d_arr_19_24 : OUT std_logic ;
      d_arr_19_23 : OUT std_logic ;
      d_arr_19_22 : OUT std_logic ;
      d_arr_19_21 : OUT std_logic ;
      d_arr_19_20 : OUT std_logic ;
      d_arr_19_19 : OUT std_logic ;
      d_arr_19_18 : OUT std_logic ;
      d_arr_19_17 : OUT std_logic ;
      d_arr_19_16 : OUT std_logic ;
      d_arr_19_15 : OUT std_logic ;
      d_arr_19_14 : OUT std_logic ;
      d_arr_19_13 : OUT std_logic ;
      d_arr_19_12 : OUT std_logic ;
      d_arr_19_11 : OUT std_logic ;
      d_arr_19_10 : OUT std_logic ;
      d_arr_19_9 : OUT std_logic ;
      d_arr_19_8 : OUT std_logic ;
      d_arr_19_7 : OUT std_logic ;
      d_arr_19_6 : OUT std_logic ;
      d_arr_19_5 : OUT std_logic ;
      d_arr_19_4 : OUT std_logic ;
      d_arr_19_3 : OUT std_logic ;
      d_arr_19_2 : OUT std_logic ;
      d_arr_19_1 : OUT std_logic ;
      d_arr_19_0 : OUT std_logic ;
      d_arr_20_31 : OUT std_logic ;
      d_arr_20_30 : OUT std_logic ;
      d_arr_20_29 : OUT std_logic ;
      d_arr_20_28 : OUT std_logic ;
      d_arr_20_27 : OUT std_logic ;
      d_arr_20_26 : OUT std_logic ;
      d_arr_20_25 : OUT std_logic ;
      d_arr_20_24 : OUT std_logic ;
      d_arr_20_23 : OUT std_logic ;
      d_arr_20_22 : OUT std_logic ;
      d_arr_20_21 : OUT std_logic ;
      d_arr_20_20 : OUT std_logic ;
      d_arr_20_19 : OUT std_logic ;
      d_arr_20_18 : OUT std_logic ;
      d_arr_20_17 : OUT std_logic ;
      d_arr_20_16 : OUT std_logic ;
      d_arr_20_15 : OUT std_logic ;
      d_arr_20_14 : OUT std_logic ;
      d_arr_20_13 : OUT std_logic ;
      d_arr_20_12 : OUT std_logic ;
      d_arr_20_11 : OUT std_logic ;
      d_arr_20_10 : OUT std_logic ;
      d_arr_20_9 : OUT std_logic ;
      d_arr_20_8 : OUT std_logic ;
      d_arr_20_7 : OUT std_logic ;
      d_arr_20_6 : OUT std_logic ;
      d_arr_20_5 : OUT std_logic ;
      d_arr_20_4 : OUT std_logic ;
      d_arr_20_3 : OUT std_logic ;
      d_arr_20_2 : OUT std_logic ;
      d_arr_20_1 : OUT std_logic ;
      d_arr_20_0 : OUT std_logic ;
      d_arr_21_31 : OUT std_logic ;
      d_arr_21_30 : OUT std_logic ;
      d_arr_21_29 : OUT std_logic ;
      d_arr_21_28 : OUT std_logic ;
      d_arr_21_27 : OUT std_logic ;
      d_arr_21_26 : OUT std_logic ;
      d_arr_21_25 : OUT std_logic ;
      d_arr_21_24 : OUT std_logic ;
      d_arr_21_23 : OUT std_logic ;
      d_arr_21_22 : OUT std_logic ;
      d_arr_21_21 : OUT std_logic ;
      d_arr_21_20 : OUT std_logic ;
      d_arr_21_19 : OUT std_logic ;
      d_arr_21_18 : OUT std_logic ;
      d_arr_21_17 : OUT std_logic ;
      d_arr_21_16 : OUT std_logic ;
      d_arr_21_15 : OUT std_logic ;
      d_arr_21_14 : OUT std_logic ;
      d_arr_21_13 : OUT std_logic ;
      d_arr_21_12 : OUT std_logic ;
      d_arr_21_11 : OUT std_logic ;
      d_arr_21_10 : OUT std_logic ;
      d_arr_21_9 : OUT std_logic ;
      d_arr_21_8 : OUT std_logic ;
      d_arr_21_7 : OUT std_logic ;
      d_arr_21_6 : OUT std_logic ;
      d_arr_21_5 : OUT std_logic ;
      d_arr_21_4 : OUT std_logic ;
      d_arr_21_3 : OUT std_logic ;
      d_arr_21_2 : OUT std_logic ;
      d_arr_21_1 : OUT std_logic ;
      d_arr_21_0 : OUT std_logic ;
      d_arr_22_31 : OUT std_logic ;
      d_arr_22_30 : OUT std_logic ;
      d_arr_22_29 : OUT std_logic ;
      d_arr_22_28 : OUT std_logic ;
      d_arr_22_27 : OUT std_logic ;
      d_arr_22_26 : OUT std_logic ;
      d_arr_22_25 : OUT std_logic ;
      d_arr_22_24 : OUT std_logic ;
      d_arr_22_23 : OUT std_logic ;
      d_arr_22_22 : OUT std_logic ;
      d_arr_22_21 : OUT std_logic ;
      d_arr_22_20 : OUT std_logic ;
      d_arr_22_19 : OUT std_logic ;
      d_arr_22_18 : OUT std_logic ;
      d_arr_22_17 : OUT std_logic ;
      d_arr_22_16 : OUT std_logic ;
      d_arr_22_15 : OUT std_logic ;
      d_arr_22_14 : OUT std_logic ;
      d_arr_22_13 : OUT std_logic ;
      d_arr_22_12 : OUT std_logic ;
      d_arr_22_11 : OUT std_logic ;
      d_arr_22_10 : OUT std_logic ;
      d_arr_22_9 : OUT std_logic ;
      d_arr_22_8 : OUT std_logic ;
      d_arr_22_7 : OUT std_logic ;
      d_arr_22_6 : OUT std_logic ;
      d_arr_22_5 : OUT std_logic ;
      d_arr_22_4 : OUT std_logic ;
      d_arr_22_3 : OUT std_logic ;
      d_arr_22_2 : OUT std_logic ;
      d_arr_22_1 : OUT std_logic ;
      d_arr_22_0 : OUT std_logic ;
      d_arr_23_31 : OUT std_logic ;
      d_arr_23_30 : OUT std_logic ;
      d_arr_23_29 : OUT std_logic ;
      d_arr_23_28 : OUT std_logic ;
      d_arr_23_27 : OUT std_logic ;
      d_arr_23_26 : OUT std_logic ;
      d_arr_23_25 : OUT std_logic ;
      d_arr_23_24 : OUT std_logic ;
      d_arr_23_23 : OUT std_logic ;
      d_arr_23_22 : OUT std_logic ;
      d_arr_23_21 : OUT std_logic ;
      d_arr_23_20 : OUT std_logic ;
      d_arr_23_19 : OUT std_logic ;
      d_arr_23_18 : OUT std_logic ;
      d_arr_23_17 : OUT std_logic ;
      d_arr_23_16 : OUT std_logic ;
      d_arr_23_15 : OUT std_logic ;
      d_arr_23_14 : OUT std_logic ;
      d_arr_23_13 : OUT std_logic ;
      d_arr_23_12 : OUT std_logic ;
      d_arr_23_11 : OUT std_logic ;
      d_arr_23_10 : OUT std_logic ;
      d_arr_23_9 : OUT std_logic ;
      d_arr_23_8 : OUT std_logic ;
      d_arr_23_7 : OUT std_logic ;
      d_arr_23_6 : OUT std_logic ;
      d_arr_23_5 : OUT std_logic ;
      d_arr_23_4 : OUT std_logic ;
      d_arr_23_3 : OUT std_logic ;
      d_arr_23_2 : OUT std_logic ;
      d_arr_23_1 : OUT std_logic ;
      d_arr_23_0 : OUT std_logic ;
      d_arr_24_31 : OUT std_logic ;
      d_arr_24_30 : OUT std_logic ;
      d_arr_24_29 : OUT std_logic ;
      d_arr_24_28 : OUT std_logic ;
      d_arr_24_27 : OUT std_logic ;
      d_arr_24_26 : OUT std_logic ;
      d_arr_24_25 : OUT std_logic ;
      d_arr_24_24 : OUT std_logic ;
      d_arr_24_23 : OUT std_logic ;
      d_arr_24_22 : OUT std_logic ;
      d_arr_24_21 : OUT std_logic ;
      d_arr_24_20 : OUT std_logic ;
      d_arr_24_19 : OUT std_logic ;
      d_arr_24_18 : OUT std_logic ;
      d_arr_24_17 : OUT std_logic ;
      d_arr_24_16 : OUT std_logic ;
      d_arr_24_15 : OUT std_logic ;
      d_arr_24_14 : OUT std_logic ;
      d_arr_24_13 : OUT std_logic ;
      d_arr_24_12 : OUT std_logic ;
      d_arr_24_11 : OUT std_logic ;
      d_arr_24_10 : OUT std_logic ;
      d_arr_24_9 : OUT std_logic ;
      d_arr_24_8 : OUT std_logic ;
      d_arr_24_7 : OUT std_logic ;
      d_arr_24_6 : OUT std_logic ;
      d_arr_24_5 : OUT std_logic ;
      d_arr_24_4 : OUT std_logic ;
      d_arr_24_3 : OUT std_logic ;
      d_arr_24_2 : OUT std_logic ;
      d_arr_24_1 : OUT std_logic ;
      d_arr_24_0 : OUT std_logic ;
      q_arr_0_31 : IN std_logic ;
      q_arr_0_30 : IN std_logic ;
      q_arr_0_29 : IN std_logic ;
      q_arr_0_28 : IN std_logic ;
      q_arr_0_27 : IN std_logic ;
      q_arr_0_26 : IN std_logic ;
      q_arr_0_25 : IN std_logic ;
      q_arr_0_24 : IN std_logic ;
      q_arr_0_23 : IN std_logic ;
      q_arr_0_22 : IN std_logic ;
      q_arr_0_21 : IN std_logic ;
      q_arr_0_20 : IN std_logic ;
      q_arr_0_19 : IN std_logic ;
      q_arr_0_18 : IN std_logic ;
      q_arr_0_17 : IN std_logic ;
      q_arr_0_16 : IN std_logic ;
      q_arr_0_15 : IN std_logic ;
      q_arr_0_14 : IN std_logic ;
      q_arr_0_13 : IN std_logic ;
      q_arr_0_12 : IN std_logic ;
      q_arr_0_11 : IN std_logic ;
      q_arr_0_10 : IN std_logic ;
      q_arr_0_9 : IN std_logic ;
      q_arr_0_8 : IN std_logic ;
      q_arr_0_7 : IN std_logic ;
      q_arr_0_6 : IN std_logic ;
      q_arr_0_5 : IN std_logic ;
      q_arr_0_4 : IN std_logic ;
      q_arr_0_3 : IN std_logic ;
      q_arr_0_2 : IN std_logic ;
      q_arr_0_1 : IN std_logic ;
      q_arr_0_0 : IN std_logic ;
      q_arr_1_31 : IN std_logic ;
      q_arr_1_30 : IN std_logic ;
      q_arr_1_29 : IN std_logic ;
      q_arr_1_28 : IN std_logic ;
      q_arr_1_27 : IN std_logic ;
      q_arr_1_26 : IN std_logic ;
      q_arr_1_25 : IN std_logic ;
      q_arr_1_24 : IN std_logic ;
      q_arr_1_23 : IN std_logic ;
      q_arr_1_22 : IN std_logic ;
      q_arr_1_21 : IN std_logic ;
      q_arr_1_20 : IN std_logic ;
      q_arr_1_19 : IN std_logic ;
      q_arr_1_18 : IN std_logic ;
      q_arr_1_17 : IN std_logic ;
      q_arr_1_16 : IN std_logic ;
      q_arr_1_15 : IN std_logic ;
      q_arr_1_14 : IN std_logic ;
      q_arr_1_13 : IN std_logic ;
      q_arr_1_12 : IN std_logic ;
      q_arr_1_11 : IN std_logic ;
      q_arr_1_10 : IN std_logic ;
      q_arr_1_9 : IN std_logic ;
      q_arr_1_8 : IN std_logic ;
      q_arr_1_7 : IN std_logic ;
      q_arr_1_6 : IN std_logic ;
      q_arr_1_5 : IN std_logic ;
      q_arr_1_4 : IN std_logic ;
      q_arr_1_3 : IN std_logic ;
      q_arr_1_2 : IN std_logic ;
      q_arr_1_1 : IN std_logic ;
      q_arr_1_0 : IN std_logic ;
      q_arr_2_31 : IN std_logic ;
      q_arr_2_30 : IN std_logic ;
      q_arr_2_29 : IN std_logic ;
      q_arr_2_28 : IN std_logic ;
      q_arr_2_27 : IN std_logic ;
      q_arr_2_26 : IN std_logic ;
      q_arr_2_25 : IN std_logic ;
      q_arr_2_24 : IN std_logic ;
      q_arr_2_23 : IN std_logic ;
      q_arr_2_22 : IN std_logic ;
      q_arr_2_21 : IN std_logic ;
      q_arr_2_20 : IN std_logic ;
      q_arr_2_19 : IN std_logic ;
      q_arr_2_18 : IN std_logic ;
      q_arr_2_17 : IN std_logic ;
      q_arr_2_16 : IN std_logic ;
      q_arr_2_15 : IN std_logic ;
      q_arr_2_14 : IN std_logic ;
      q_arr_2_13 : IN std_logic ;
      q_arr_2_12 : IN std_logic ;
      q_arr_2_11 : IN std_logic ;
      q_arr_2_10 : IN std_logic ;
      q_arr_2_9 : IN std_logic ;
      q_arr_2_8 : IN std_logic ;
      q_arr_2_7 : IN std_logic ;
      q_arr_2_6 : IN std_logic ;
      q_arr_2_5 : IN std_logic ;
      q_arr_2_4 : IN std_logic ;
      q_arr_2_3 : IN std_logic ;
      q_arr_2_2 : IN std_logic ;
      q_arr_2_1 : IN std_logic ;
      q_arr_2_0 : IN std_logic ;
      q_arr_3_31 : IN std_logic ;
      q_arr_3_30 : IN std_logic ;
      q_arr_3_29 : IN std_logic ;
      q_arr_3_28 : IN std_logic ;
      q_arr_3_27 : IN std_logic ;
      q_arr_3_26 : IN std_logic ;
      q_arr_3_25 : IN std_logic ;
      q_arr_3_24 : IN std_logic ;
      q_arr_3_23 : IN std_logic ;
      q_arr_3_22 : IN std_logic ;
      q_arr_3_21 : IN std_logic ;
      q_arr_3_20 : IN std_logic ;
      q_arr_3_19 : IN std_logic ;
      q_arr_3_18 : IN std_logic ;
      q_arr_3_17 : IN std_logic ;
      q_arr_3_16 : IN std_logic ;
      q_arr_3_15 : IN std_logic ;
      q_arr_3_14 : IN std_logic ;
      q_arr_3_13 : IN std_logic ;
      q_arr_3_12 : IN std_logic ;
      q_arr_3_11 : IN std_logic ;
      q_arr_3_10 : IN std_logic ;
      q_arr_3_9 : IN std_logic ;
      q_arr_3_8 : IN std_logic ;
      q_arr_3_7 : IN std_logic ;
      q_arr_3_6 : IN std_logic ;
      q_arr_3_5 : IN std_logic ;
      q_arr_3_4 : IN std_logic ;
      q_arr_3_3 : IN std_logic ;
      q_arr_3_2 : IN std_logic ;
      q_arr_3_1 : IN std_logic ;
      q_arr_3_0 : IN std_logic ;
      q_arr_4_31 : IN std_logic ;
      q_arr_4_30 : IN std_logic ;
      q_arr_4_29 : IN std_logic ;
      q_arr_4_28 : IN std_logic ;
      q_arr_4_27 : IN std_logic ;
      q_arr_4_26 : IN std_logic ;
      q_arr_4_25 : IN std_logic ;
      q_arr_4_24 : IN std_logic ;
      q_arr_4_23 : IN std_logic ;
      q_arr_4_22 : IN std_logic ;
      q_arr_4_21 : IN std_logic ;
      q_arr_4_20 : IN std_logic ;
      q_arr_4_19 : IN std_logic ;
      q_arr_4_18 : IN std_logic ;
      q_arr_4_17 : IN std_logic ;
      q_arr_4_16 : IN std_logic ;
      q_arr_4_15 : IN std_logic ;
      q_arr_4_14 : IN std_logic ;
      q_arr_4_13 : IN std_logic ;
      q_arr_4_12 : IN std_logic ;
      q_arr_4_11 : IN std_logic ;
      q_arr_4_10 : IN std_logic ;
      q_arr_4_9 : IN std_logic ;
      q_arr_4_8 : IN std_logic ;
      q_arr_4_7 : IN std_logic ;
      q_arr_4_6 : IN std_logic ;
      q_arr_4_5 : IN std_logic ;
      q_arr_4_4 : IN std_logic ;
      q_arr_4_3 : IN std_logic ;
      q_arr_4_2 : IN std_logic ;
      q_arr_4_1 : IN std_logic ;
      q_arr_4_0 : IN std_logic ;
      q_arr_5_31 : IN std_logic ;
      q_arr_5_30 : IN std_logic ;
      q_arr_5_29 : IN std_logic ;
      q_arr_5_28 : IN std_logic ;
      q_arr_5_27 : IN std_logic ;
      q_arr_5_26 : IN std_logic ;
      q_arr_5_25 : IN std_logic ;
      q_arr_5_24 : IN std_logic ;
      q_arr_5_23 : IN std_logic ;
      q_arr_5_22 : IN std_logic ;
      q_arr_5_21 : IN std_logic ;
      q_arr_5_20 : IN std_logic ;
      q_arr_5_19 : IN std_logic ;
      q_arr_5_18 : IN std_logic ;
      q_arr_5_17 : IN std_logic ;
      q_arr_5_16 : IN std_logic ;
      q_arr_5_15 : IN std_logic ;
      q_arr_5_14 : IN std_logic ;
      q_arr_5_13 : IN std_logic ;
      q_arr_5_12 : IN std_logic ;
      q_arr_5_11 : IN std_logic ;
      q_arr_5_10 : IN std_logic ;
      q_arr_5_9 : IN std_logic ;
      q_arr_5_8 : IN std_logic ;
      q_arr_5_7 : IN std_logic ;
      q_arr_5_6 : IN std_logic ;
      q_arr_5_5 : IN std_logic ;
      q_arr_5_4 : IN std_logic ;
      q_arr_5_3 : IN std_logic ;
      q_arr_5_2 : IN std_logic ;
      q_arr_5_1 : IN std_logic ;
      q_arr_5_0 : IN std_logic ;
      q_arr_6_31 : IN std_logic ;
      q_arr_6_30 : IN std_logic ;
      q_arr_6_29 : IN std_logic ;
      q_arr_6_28 : IN std_logic ;
      q_arr_6_27 : IN std_logic ;
      q_arr_6_26 : IN std_logic ;
      q_arr_6_25 : IN std_logic ;
      q_arr_6_24 : IN std_logic ;
      q_arr_6_23 : IN std_logic ;
      q_arr_6_22 : IN std_logic ;
      q_arr_6_21 : IN std_logic ;
      q_arr_6_20 : IN std_logic ;
      q_arr_6_19 : IN std_logic ;
      q_arr_6_18 : IN std_logic ;
      q_arr_6_17 : IN std_logic ;
      q_arr_6_16 : IN std_logic ;
      q_arr_6_15 : IN std_logic ;
      q_arr_6_14 : IN std_logic ;
      q_arr_6_13 : IN std_logic ;
      q_arr_6_12 : IN std_logic ;
      q_arr_6_11 : IN std_logic ;
      q_arr_6_10 : IN std_logic ;
      q_arr_6_9 : IN std_logic ;
      q_arr_6_8 : IN std_logic ;
      q_arr_6_7 : IN std_logic ;
      q_arr_6_6 : IN std_logic ;
      q_arr_6_5 : IN std_logic ;
      q_arr_6_4 : IN std_logic ;
      q_arr_6_3 : IN std_logic ;
      q_arr_6_2 : IN std_logic ;
      q_arr_6_1 : IN std_logic ;
      q_arr_6_0 : IN std_logic ;
      q_arr_7_31 : IN std_logic ;
      q_arr_7_30 : IN std_logic ;
      q_arr_7_29 : IN std_logic ;
      q_arr_7_28 : IN std_logic ;
      q_arr_7_27 : IN std_logic ;
      q_arr_7_26 : IN std_logic ;
      q_arr_7_25 : IN std_logic ;
      q_arr_7_24 : IN std_logic ;
      q_arr_7_23 : IN std_logic ;
      q_arr_7_22 : IN std_logic ;
      q_arr_7_21 : IN std_logic ;
      q_arr_7_20 : IN std_logic ;
      q_arr_7_19 : IN std_logic ;
      q_arr_7_18 : IN std_logic ;
      q_arr_7_17 : IN std_logic ;
      q_arr_7_16 : IN std_logic ;
      q_arr_7_15 : IN std_logic ;
      q_arr_7_14 : IN std_logic ;
      q_arr_7_13 : IN std_logic ;
      q_arr_7_12 : IN std_logic ;
      q_arr_7_11 : IN std_logic ;
      q_arr_7_10 : IN std_logic ;
      q_arr_7_9 : IN std_logic ;
      q_arr_7_8 : IN std_logic ;
      q_arr_7_7 : IN std_logic ;
      q_arr_7_6 : IN std_logic ;
      q_arr_7_5 : IN std_logic ;
      q_arr_7_4 : IN std_logic ;
      q_arr_7_3 : IN std_logic ;
      q_arr_7_2 : IN std_logic ;
      q_arr_7_1 : IN std_logic ;
      q_arr_7_0 : IN std_logic ;
      q_arr_8_31 : IN std_logic ;
      q_arr_8_30 : IN std_logic ;
      q_arr_8_29 : IN std_logic ;
      q_arr_8_28 : IN std_logic ;
      q_arr_8_27 : IN std_logic ;
      q_arr_8_26 : IN std_logic ;
      q_arr_8_25 : IN std_logic ;
      q_arr_8_24 : IN std_logic ;
      q_arr_8_23 : IN std_logic ;
      q_arr_8_22 : IN std_logic ;
      q_arr_8_21 : IN std_logic ;
      q_arr_8_20 : IN std_logic ;
      q_arr_8_19 : IN std_logic ;
      q_arr_8_18 : IN std_logic ;
      q_arr_8_17 : IN std_logic ;
      q_arr_8_16 : IN std_logic ;
      q_arr_8_15 : IN std_logic ;
      q_arr_8_14 : IN std_logic ;
      q_arr_8_13 : IN std_logic ;
      q_arr_8_12 : IN std_logic ;
      q_arr_8_11 : IN std_logic ;
      q_arr_8_10 : IN std_logic ;
      q_arr_8_9 : IN std_logic ;
      q_arr_8_8 : IN std_logic ;
      q_arr_8_7 : IN std_logic ;
      q_arr_8_6 : IN std_logic ;
      q_arr_8_5 : IN std_logic ;
      q_arr_8_4 : IN std_logic ;
      q_arr_8_3 : IN std_logic ;
      q_arr_8_2 : IN std_logic ;
      q_arr_8_1 : IN std_logic ;
      q_arr_8_0 : IN std_logic ;
      q_arr_9_31 : IN std_logic ;
      q_arr_9_30 : IN std_logic ;
      q_arr_9_29 : IN std_logic ;
      q_arr_9_28 : IN std_logic ;
      q_arr_9_27 : IN std_logic ;
      q_arr_9_26 : IN std_logic ;
      q_arr_9_25 : IN std_logic ;
      q_arr_9_24 : IN std_logic ;
      q_arr_9_23 : IN std_logic ;
      q_arr_9_22 : IN std_logic ;
      q_arr_9_21 : IN std_logic ;
      q_arr_9_20 : IN std_logic ;
      q_arr_9_19 : IN std_logic ;
      q_arr_9_18 : IN std_logic ;
      q_arr_9_17 : IN std_logic ;
      q_arr_9_16 : IN std_logic ;
      q_arr_9_15 : IN std_logic ;
      q_arr_9_14 : IN std_logic ;
      q_arr_9_13 : IN std_logic ;
      q_arr_9_12 : IN std_logic ;
      q_arr_9_11 : IN std_logic ;
      q_arr_9_10 : IN std_logic ;
      q_arr_9_9 : IN std_logic ;
      q_arr_9_8 : IN std_logic ;
      q_arr_9_7 : IN std_logic ;
      q_arr_9_6 : IN std_logic ;
      q_arr_9_5 : IN std_logic ;
      q_arr_9_4 : IN std_logic ;
      q_arr_9_3 : IN std_logic ;
      q_arr_9_2 : IN std_logic ;
      q_arr_9_1 : IN std_logic ;
      q_arr_9_0 : IN std_logic ;
      q_arr_10_31 : IN std_logic ;
      q_arr_10_30 : IN std_logic ;
      q_arr_10_29 : IN std_logic ;
      q_arr_10_28 : IN std_logic ;
      q_arr_10_27 : IN std_logic ;
      q_arr_10_26 : IN std_logic ;
      q_arr_10_25 : IN std_logic ;
      q_arr_10_24 : IN std_logic ;
      q_arr_10_23 : IN std_logic ;
      q_arr_10_22 : IN std_logic ;
      q_arr_10_21 : IN std_logic ;
      q_arr_10_20 : IN std_logic ;
      q_arr_10_19 : IN std_logic ;
      q_arr_10_18 : IN std_logic ;
      q_arr_10_17 : IN std_logic ;
      q_arr_10_16 : IN std_logic ;
      q_arr_10_15 : IN std_logic ;
      q_arr_10_14 : IN std_logic ;
      q_arr_10_13 : IN std_logic ;
      q_arr_10_12 : IN std_logic ;
      q_arr_10_11 : IN std_logic ;
      q_arr_10_10 : IN std_logic ;
      q_arr_10_9 : IN std_logic ;
      q_arr_10_8 : IN std_logic ;
      q_arr_10_7 : IN std_logic ;
      q_arr_10_6 : IN std_logic ;
      q_arr_10_5 : IN std_logic ;
      q_arr_10_4 : IN std_logic ;
      q_arr_10_3 : IN std_logic ;
      q_arr_10_2 : IN std_logic ;
      q_arr_10_1 : IN std_logic ;
      q_arr_10_0 : IN std_logic ;
      q_arr_11_31 : IN std_logic ;
      q_arr_11_30 : IN std_logic ;
      q_arr_11_29 : IN std_logic ;
      q_arr_11_28 : IN std_logic ;
      q_arr_11_27 : IN std_logic ;
      q_arr_11_26 : IN std_logic ;
      q_arr_11_25 : IN std_logic ;
      q_arr_11_24 : IN std_logic ;
      q_arr_11_23 : IN std_logic ;
      q_arr_11_22 : IN std_logic ;
      q_arr_11_21 : IN std_logic ;
      q_arr_11_20 : IN std_logic ;
      q_arr_11_19 : IN std_logic ;
      q_arr_11_18 : IN std_logic ;
      q_arr_11_17 : IN std_logic ;
      q_arr_11_16 : IN std_logic ;
      q_arr_11_15 : IN std_logic ;
      q_arr_11_14 : IN std_logic ;
      q_arr_11_13 : IN std_logic ;
      q_arr_11_12 : IN std_logic ;
      q_arr_11_11 : IN std_logic ;
      q_arr_11_10 : IN std_logic ;
      q_arr_11_9 : IN std_logic ;
      q_arr_11_8 : IN std_logic ;
      q_arr_11_7 : IN std_logic ;
      q_arr_11_6 : IN std_logic ;
      q_arr_11_5 : IN std_logic ;
      q_arr_11_4 : IN std_logic ;
      q_arr_11_3 : IN std_logic ;
      q_arr_11_2 : IN std_logic ;
      q_arr_11_1 : IN std_logic ;
      q_arr_11_0 : IN std_logic ;
      q_arr_12_31 : IN std_logic ;
      q_arr_12_30 : IN std_logic ;
      q_arr_12_29 : IN std_logic ;
      q_arr_12_28 : IN std_logic ;
      q_arr_12_27 : IN std_logic ;
      q_arr_12_26 : IN std_logic ;
      q_arr_12_25 : IN std_logic ;
      q_arr_12_24 : IN std_logic ;
      q_arr_12_23 : IN std_logic ;
      q_arr_12_22 : IN std_logic ;
      q_arr_12_21 : IN std_logic ;
      q_arr_12_20 : IN std_logic ;
      q_arr_12_19 : IN std_logic ;
      q_arr_12_18 : IN std_logic ;
      q_arr_12_17 : IN std_logic ;
      q_arr_12_16 : IN std_logic ;
      q_arr_12_15 : IN std_logic ;
      q_arr_12_14 : IN std_logic ;
      q_arr_12_13 : IN std_logic ;
      q_arr_12_12 : IN std_logic ;
      q_arr_12_11 : IN std_logic ;
      q_arr_12_10 : IN std_logic ;
      q_arr_12_9 : IN std_logic ;
      q_arr_12_8 : IN std_logic ;
      q_arr_12_7 : IN std_logic ;
      q_arr_12_6 : IN std_logic ;
      q_arr_12_5 : IN std_logic ;
      q_arr_12_4 : IN std_logic ;
      q_arr_12_3 : IN std_logic ;
      q_arr_12_2 : IN std_logic ;
      q_arr_12_1 : IN std_logic ;
      q_arr_12_0 : IN std_logic ;
      q_arr_13_31 : IN std_logic ;
      q_arr_13_30 : IN std_logic ;
      q_arr_13_29 : IN std_logic ;
      q_arr_13_28 : IN std_logic ;
      q_arr_13_27 : IN std_logic ;
      q_arr_13_26 : IN std_logic ;
      q_arr_13_25 : IN std_logic ;
      q_arr_13_24 : IN std_logic ;
      q_arr_13_23 : IN std_logic ;
      q_arr_13_22 : IN std_logic ;
      q_arr_13_21 : IN std_logic ;
      q_arr_13_20 : IN std_logic ;
      q_arr_13_19 : IN std_logic ;
      q_arr_13_18 : IN std_logic ;
      q_arr_13_17 : IN std_logic ;
      q_arr_13_16 : IN std_logic ;
      q_arr_13_15 : IN std_logic ;
      q_arr_13_14 : IN std_logic ;
      q_arr_13_13 : IN std_logic ;
      q_arr_13_12 : IN std_logic ;
      q_arr_13_11 : IN std_logic ;
      q_arr_13_10 : IN std_logic ;
      q_arr_13_9 : IN std_logic ;
      q_arr_13_8 : IN std_logic ;
      q_arr_13_7 : IN std_logic ;
      q_arr_13_6 : IN std_logic ;
      q_arr_13_5 : IN std_logic ;
      q_arr_13_4 : IN std_logic ;
      q_arr_13_3 : IN std_logic ;
      q_arr_13_2 : IN std_logic ;
      q_arr_13_1 : IN std_logic ;
      q_arr_13_0 : IN std_logic ;
      q_arr_14_31 : IN std_logic ;
      q_arr_14_30 : IN std_logic ;
      q_arr_14_29 : IN std_logic ;
      q_arr_14_28 : IN std_logic ;
      q_arr_14_27 : IN std_logic ;
      q_arr_14_26 : IN std_logic ;
      q_arr_14_25 : IN std_logic ;
      q_arr_14_24 : IN std_logic ;
      q_arr_14_23 : IN std_logic ;
      q_arr_14_22 : IN std_logic ;
      q_arr_14_21 : IN std_logic ;
      q_arr_14_20 : IN std_logic ;
      q_arr_14_19 : IN std_logic ;
      q_arr_14_18 : IN std_logic ;
      q_arr_14_17 : IN std_logic ;
      q_arr_14_16 : IN std_logic ;
      q_arr_14_15 : IN std_logic ;
      q_arr_14_14 : IN std_logic ;
      q_arr_14_13 : IN std_logic ;
      q_arr_14_12 : IN std_logic ;
      q_arr_14_11 : IN std_logic ;
      q_arr_14_10 : IN std_logic ;
      q_arr_14_9 : IN std_logic ;
      q_arr_14_8 : IN std_logic ;
      q_arr_14_7 : IN std_logic ;
      q_arr_14_6 : IN std_logic ;
      q_arr_14_5 : IN std_logic ;
      q_arr_14_4 : IN std_logic ;
      q_arr_14_3 : IN std_logic ;
      q_arr_14_2 : IN std_logic ;
      q_arr_14_1 : IN std_logic ;
      q_arr_14_0 : IN std_logic ;
      q_arr_15_31 : IN std_logic ;
      q_arr_15_30 : IN std_logic ;
      q_arr_15_29 : IN std_logic ;
      q_arr_15_28 : IN std_logic ;
      q_arr_15_27 : IN std_logic ;
      q_arr_15_26 : IN std_logic ;
      q_arr_15_25 : IN std_logic ;
      q_arr_15_24 : IN std_logic ;
      q_arr_15_23 : IN std_logic ;
      q_arr_15_22 : IN std_logic ;
      q_arr_15_21 : IN std_logic ;
      q_arr_15_20 : IN std_logic ;
      q_arr_15_19 : IN std_logic ;
      q_arr_15_18 : IN std_logic ;
      q_arr_15_17 : IN std_logic ;
      q_arr_15_16 : IN std_logic ;
      q_arr_15_15 : IN std_logic ;
      q_arr_15_14 : IN std_logic ;
      q_arr_15_13 : IN std_logic ;
      q_arr_15_12 : IN std_logic ;
      q_arr_15_11 : IN std_logic ;
      q_arr_15_10 : IN std_logic ;
      q_arr_15_9 : IN std_logic ;
      q_arr_15_8 : IN std_logic ;
      q_arr_15_7 : IN std_logic ;
      q_arr_15_6 : IN std_logic ;
      q_arr_15_5 : IN std_logic ;
      q_arr_15_4 : IN std_logic ;
      q_arr_15_3 : IN std_logic ;
      q_arr_15_2 : IN std_logic ;
      q_arr_15_1 : IN std_logic ;
      q_arr_15_0 : IN std_logic ;
      q_arr_16_31 : IN std_logic ;
      q_arr_16_30 : IN std_logic ;
      q_arr_16_29 : IN std_logic ;
      q_arr_16_28 : IN std_logic ;
      q_arr_16_27 : IN std_logic ;
      q_arr_16_26 : IN std_logic ;
      q_arr_16_25 : IN std_logic ;
      q_arr_16_24 : IN std_logic ;
      q_arr_16_23 : IN std_logic ;
      q_arr_16_22 : IN std_logic ;
      q_arr_16_21 : IN std_logic ;
      q_arr_16_20 : IN std_logic ;
      q_arr_16_19 : IN std_logic ;
      q_arr_16_18 : IN std_logic ;
      q_arr_16_17 : IN std_logic ;
      q_arr_16_16 : IN std_logic ;
      q_arr_16_15 : IN std_logic ;
      q_arr_16_14 : IN std_logic ;
      q_arr_16_13 : IN std_logic ;
      q_arr_16_12 : IN std_logic ;
      q_arr_16_11 : IN std_logic ;
      q_arr_16_10 : IN std_logic ;
      q_arr_16_9 : IN std_logic ;
      q_arr_16_8 : IN std_logic ;
      q_arr_16_7 : IN std_logic ;
      q_arr_16_6 : IN std_logic ;
      q_arr_16_5 : IN std_logic ;
      q_arr_16_4 : IN std_logic ;
      q_arr_16_3 : IN std_logic ;
      q_arr_16_2 : IN std_logic ;
      q_arr_16_1 : IN std_logic ;
      q_arr_16_0 : IN std_logic ;
      q_arr_17_31 : IN std_logic ;
      q_arr_17_30 : IN std_logic ;
      q_arr_17_29 : IN std_logic ;
      q_arr_17_28 : IN std_logic ;
      q_arr_17_27 : IN std_logic ;
      q_arr_17_26 : IN std_logic ;
      q_arr_17_25 : IN std_logic ;
      q_arr_17_24 : IN std_logic ;
      q_arr_17_23 : IN std_logic ;
      q_arr_17_22 : IN std_logic ;
      q_arr_17_21 : IN std_logic ;
      q_arr_17_20 : IN std_logic ;
      q_arr_17_19 : IN std_logic ;
      q_arr_17_18 : IN std_logic ;
      q_arr_17_17 : IN std_logic ;
      q_arr_17_16 : IN std_logic ;
      q_arr_17_15 : IN std_logic ;
      q_arr_17_14 : IN std_logic ;
      q_arr_17_13 : IN std_logic ;
      q_arr_17_12 : IN std_logic ;
      q_arr_17_11 : IN std_logic ;
      q_arr_17_10 : IN std_logic ;
      q_arr_17_9 : IN std_logic ;
      q_arr_17_8 : IN std_logic ;
      q_arr_17_7 : IN std_logic ;
      q_arr_17_6 : IN std_logic ;
      q_arr_17_5 : IN std_logic ;
      q_arr_17_4 : IN std_logic ;
      q_arr_17_3 : IN std_logic ;
      q_arr_17_2 : IN std_logic ;
      q_arr_17_1 : IN std_logic ;
      q_arr_17_0 : IN std_logic ;
      q_arr_18_31 : IN std_logic ;
      q_arr_18_30 : IN std_logic ;
      q_arr_18_29 : IN std_logic ;
      q_arr_18_28 : IN std_logic ;
      q_arr_18_27 : IN std_logic ;
      q_arr_18_26 : IN std_logic ;
      q_arr_18_25 : IN std_logic ;
      q_arr_18_24 : IN std_logic ;
      q_arr_18_23 : IN std_logic ;
      q_arr_18_22 : IN std_logic ;
      q_arr_18_21 : IN std_logic ;
      q_arr_18_20 : IN std_logic ;
      q_arr_18_19 : IN std_logic ;
      q_arr_18_18 : IN std_logic ;
      q_arr_18_17 : IN std_logic ;
      q_arr_18_16 : IN std_logic ;
      q_arr_18_15 : IN std_logic ;
      q_arr_18_14 : IN std_logic ;
      q_arr_18_13 : IN std_logic ;
      q_arr_18_12 : IN std_logic ;
      q_arr_18_11 : IN std_logic ;
      q_arr_18_10 : IN std_logic ;
      q_arr_18_9 : IN std_logic ;
      q_arr_18_8 : IN std_logic ;
      q_arr_18_7 : IN std_logic ;
      q_arr_18_6 : IN std_logic ;
      q_arr_18_5 : IN std_logic ;
      q_arr_18_4 : IN std_logic ;
      q_arr_18_3 : IN std_logic ;
      q_arr_18_2 : IN std_logic ;
      q_arr_18_1 : IN std_logic ;
      q_arr_18_0 : IN std_logic ;
      q_arr_19_31 : IN std_logic ;
      q_arr_19_30 : IN std_logic ;
      q_arr_19_29 : IN std_logic ;
      q_arr_19_28 : IN std_logic ;
      q_arr_19_27 : IN std_logic ;
      q_arr_19_26 : IN std_logic ;
      q_arr_19_25 : IN std_logic ;
      q_arr_19_24 : IN std_logic ;
      q_arr_19_23 : IN std_logic ;
      q_arr_19_22 : IN std_logic ;
      q_arr_19_21 : IN std_logic ;
      q_arr_19_20 : IN std_logic ;
      q_arr_19_19 : IN std_logic ;
      q_arr_19_18 : IN std_logic ;
      q_arr_19_17 : IN std_logic ;
      q_arr_19_16 : IN std_logic ;
      q_arr_19_15 : IN std_logic ;
      q_arr_19_14 : IN std_logic ;
      q_arr_19_13 : IN std_logic ;
      q_arr_19_12 : IN std_logic ;
      q_arr_19_11 : IN std_logic ;
      q_arr_19_10 : IN std_logic ;
      q_arr_19_9 : IN std_logic ;
      q_arr_19_8 : IN std_logic ;
      q_arr_19_7 : IN std_logic ;
      q_arr_19_6 : IN std_logic ;
      q_arr_19_5 : IN std_logic ;
      q_arr_19_4 : IN std_logic ;
      q_arr_19_3 : IN std_logic ;
      q_arr_19_2 : IN std_logic ;
      q_arr_19_1 : IN std_logic ;
      q_arr_19_0 : IN std_logic ;
      q_arr_20_31 : IN std_logic ;
      q_arr_20_30 : IN std_logic ;
      q_arr_20_29 : IN std_logic ;
      q_arr_20_28 : IN std_logic ;
      q_arr_20_27 : IN std_logic ;
      q_arr_20_26 : IN std_logic ;
      q_arr_20_25 : IN std_logic ;
      q_arr_20_24 : IN std_logic ;
      q_arr_20_23 : IN std_logic ;
      q_arr_20_22 : IN std_logic ;
      q_arr_20_21 : IN std_logic ;
      q_arr_20_20 : IN std_logic ;
      q_arr_20_19 : IN std_logic ;
      q_arr_20_18 : IN std_logic ;
      q_arr_20_17 : IN std_logic ;
      q_arr_20_16 : IN std_logic ;
      q_arr_20_15 : IN std_logic ;
      q_arr_20_14 : IN std_logic ;
      q_arr_20_13 : IN std_logic ;
      q_arr_20_12 : IN std_logic ;
      q_arr_20_11 : IN std_logic ;
      q_arr_20_10 : IN std_logic ;
      q_arr_20_9 : IN std_logic ;
      q_arr_20_8 : IN std_logic ;
      q_arr_20_7 : IN std_logic ;
      q_arr_20_6 : IN std_logic ;
      q_arr_20_5 : IN std_logic ;
      q_arr_20_4 : IN std_logic ;
      q_arr_20_3 : IN std_logic ;
      q_arr_20_2 : IN std_logic ;
      q_arr_20_1 : IN std_logic ;
      q_arr_20_0 : IN std_logic ;
      q_arr_21_31 : IN std_logic ;
      q_arr_21_30 : IN std_logic ;
      q_arr_21_29 : IN std_logic ;
      q_arr_21_28 : IN std_logic ;
      q_arr_21_27 : IN std_logic ;
      q_arr_21_26 : IN std_logic ;
      q_arr_21_25 : IN std_logic ;
      q_arr_21_24 : IN std_logic ;
      q_arr_21_23 : IN std_logic ;
      q_arr_21_22 : IN std_logic ;
      q_arr_21_21 : IN std_logic ;
      q_arr_21_20 : IN std_logic ;
      q_arr_21_19 : IN std_logic ;
      q_arr_21_18 : IN std_logic ;
      q_arr_21_17 : IN std_logic ;
      q_arr_21_16 : IN std_logic ;
      q_arr_21_15 : IN std_logic ;
      q_arr_21_14 : IN std_logic ;
      q_arr_21_13 : IN std_logic ;
      q_arr_21_12 : IN std_logic ;
      q_arr_21_11 : IN std_logic ;
      q_arr_21_10 : IN std_logic ;
      q_arr_21_9 : IN std_logic ;
      q_arr_21_8 : IN std_logic ;
      q_arr_21_7 : IN std_logic ;
      q_arr_21_6 : IN std_logic ;
      q_arr_21_5 : IN std_logic ;
      q_arr_21_4 : IN std_logic ;
      q_arr_21_3 : IN std_logic ;
      q_arr_21_2 : IN std_logic ;
      q_arr_21_1 : IN std_logic ;
      q_arr_21_0 : IN std_logic ;
      q_arr_22_31 : IN std_logic ;
      q_arr_22_30 : IN std_logic ;
      q_arr_22_29 : IN std_logic ;
      q_arr_22_28 : IN std_logic ;
      q_arr_22_27 : IN std_logic ;
      q_arr_22_26 : IN std_logic ;
      q_arr_22_25 : IN std_logic ;
      q_arr_22_24 : IN std_logic ;
      q_arr_22_23 : IN std_logic ;
      q_arr_22_22 : IN std_logic ;
      q_arr_22_21 : IN std_logic ;
      q_arr_22_20 : IN std_logic ;
      q_arr_22_19 : IN std_logic ;
      q_arr_22_18 : IN std_logic ;
      q_arr_22_17 : IN std_logic ;
      q_arr_22_16 : IN std_logic ;
      q_arr_22_15 : IN std_logic ;
      q_arr_22_14 : IN std_logic ;
      q_arr_22_13 : IN std_logic ;
      q_arr_22_12 : IN std_logic ;
      q_arr_22_11 : IN std_logic ;
      q_arr_22_10 : IN std_logic ;
      q_arr_22_9 : IN std_logic ;
      q_arr_22_8 : IN std_logic ;
      q_arr_22_7 : IN std_logic ;
      q_arr_22_6 : IN std_logic ;
      q_arr_22_5 : IN std_logic ;
      q_arr_22_4 : IN std_logic ;
      q_arr_22_3 : IN std_logic ;
      q_arr_22_2 : IN std_logic ;
      q_arr_22_1 : IN std_logic ;
      q_arr_22_0 : IN std_logic ;
      q_arr_23_31 : IN std_logic ;
      q_arr_23_30 : IN std_logic ;
      q_arr_23_29 : IN std_logic ;
      q_arr_23_28 : IN std_logic ;
      q_arr_23_27 : IN std_logic ;
      q_arr_23_26 : IN std_logic ;
      q_arr_23_25 : IN std_logic ;
      q_arr_23_24 : IN std_logic ;
      q_arr_23_23 : IN std_logic ;
      q_arr_23_22 : IN std_logic ;
      q_arr_23_21 : IN std_logic ;
      q_arr_23_20 : IN std_logic ;
      q_arr_23_19 : IN std_logic ;
      q_arr_23_18 : IN std_logic ;
      q_arr_23_17 : IN std_logic ;
      q_arr_23_16 : IN std_logic ;
      q_arr_23_15 : IN std_logic ;
      q_arr_23_14 : IN std_logic ;
      q_arr_23_13 : IN std_logic ;
      q_arr_23_12 : IN std_logic ;
      q_arr_23_11 : IN std_logic ;
      q_arr_23_10 : IN std_logic ;
      q_arr_23_9 : IN std_logic ;
      q_arr_23_8 : IN std_logic ;
      q_arr_23_7 : IN std_logic ;
      q_arr_23_6 : IN std_logic ;
      q_arr_23_5 : IN std_logic ;
      q_arr_23_4 : IN std_logic ;
      q_arr_23_3 : IN std_logic ;
      q_arr_23_2 : IN std_logic ;
      q_arr_23_1 : IN std_logic ;
      q_arr_23_0 : IN std_logic ;
      q_arr_24_31 : IN std_logic ;
      q_arr_24_30 : IN std_logic ;
      q_arr_24_29 : IN std_logic ;
      q_arr_24_28 : IN std_logic ;
      q_arr_24_27 : IN std_logic ;
      q_arr_24_26 : IN std_logic ;
      q_arr_24_25 : IN std_logic ;
      q_arr_24_24 : IN std_logic ;
      q_arr_24_23 : IN std_logic ;
      q_arr_24_22 : IN std_logic ;
      q_arr_24_21 : IN std_logic ;
      q_arr_24_20 : IN std_logic ;
      q_arr_24_19 : IN std_logic ;
      q_arr_24_18 : IN std_logic ;
      q_arr_24_17 : IN std_logic ;
      q_arr_24_16 : IN std_logic ;
      q_arr_24_15 : IN std_logic ;
      q_arr_24_14 : IN std_logic ;
      q_arr_24_13 : IN std_logic ;
      q_arr_24_12 : IN std_logic ;
      q_arr_24_11 : IN std_logic ;
      q_arr_24_10 : IN std_logic ;
      q_arr_24_9 : IN std_logic ;
      q_arr_24_8 : IN std_logic ;
      q_arr_24_7 : IN std_logic ;
      q_arr_24_6 : IN std_logic ;
      q_arr_24_5 : IN std_logic ;
      q_arr_24_4 : IN std_logic ;
      q_arr_24_3 : IN std_logic ;
      q_arr_24_2 : IN std_logic ;
      q_arr_24_1 : IN std_logic ;
      q_arr_24_0 : IN std_logic ;
      operation : IN std_logic ;
      filter_size : IN std_logic) ;
end MergeLayer ;

architecture Structural_unfold_3382_0 of MergeLayer is
   component NAdder_32
      port (
         a : IN std_logic_vector (31 DOWNTO 0) ;
         b : IN std_logic_vector (31 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (31 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal s1_31, s1_30, s1_29, s1_28, s1_27, s1_26, s1_25, s1_24, s1_23, 
      s1_22, s1_21, s1_20, s1_19, s1_18, s1_17, s1_16, s1_15, s1_14, s1_13, 
      s1_12, s1_11, s1_10, s1_9, s1_8, s1_7, s1_6, s1_5, s1_4, s1_3, s1_2, 
      s1_1, s1_0, s2_31, s2_30, s2_29, s2_28, s2_27, s2_26, s2_25, s2_24, 
      s2_23, s2_22, s2_21, s2_20, s2_19, s2_18, s2_17, s2_16, s2_15, s2_14, 
      s2_13, s2_12, s2_11, s2_10, s2_9, s2_8, s2_7, s2_6, s2_5, s2_4, s2_3, 
      s2_2, s2_1, s2_0, d_arr_24_0_EXMPLR, nx6, nx10, nx350, nx153, nx165, 
      nx169, nx173, nx177, nx181, nx185, nx189, nx193, nx197, nx201, nx205, 
      nx209, nx213, nx217, nx221, nx225, nx229, nx233, nx237, nx241, nx245, 
      nx249, nx253, nx257, nx261, nx265, nx277, nx279, nx285, nx287, nx291, 
      nx293, nx297, nx299, nx303, nx305, nx309, nx311, nx315, nx317, nx321, 
      nx323, nx327, nx329, nx333, nx335, nx339, nx341, nx345, nx347, nx351, 
      nx353, nx357, nx359, nx363, nx365, nx369, nx371, nx375, nx377, nx381, 
      nx383, nx387, nx389, nx393, nx395, nx399, nx401, nx405, nx407, nx411, 
      nx413, nx417, nx419, nx423, nx425, nx429, nx431, nx435, nx437, nx441, 
      nx445, nx458, nx460, nx462, nx464, nx466, nx469, nx471, nx473, nx475, 
      nx477, nx479, nx481, nx483, nx485, nx487, nx489, nx491, nx493, nx495, 
      nx497, nx499, nx501, nx503, nx505, nx507, nx509, nx511, nx513, nx515, 
      nx517, nx519, nx521, nx523, nx525, nx527, nx529, nx531, nx533, nx540, 
      nx542, nx550, nx553, nx555: std_logic ;
   
   signal DANGLING : std_logic_vector (1 downto 0 );

begin
   d_arr_2_31 <= d_arr_24_0_EXMPLR ;
   d_arr_2_30 <= d_arr_24_0_EXMPLR ;
   d_arr_2_29 <= d_arr_24_0_EXMPLR ;
   d_arr_2_28 <= d_arr_24_0_EXMPLR ;
   d_arr_2_27 <= d_arr_24_0_EXMPLR ;
   d_arr_2_26 <= d_arr_24_0_EXMPLR ;
   d_arr_2_25 <= d_arr_24_0_EXMPLR ;
   d_arr_2_24 <= d_arr_24_0_EXMPLR ;
   d_arr_2_23 <= d_arr_24_0_EXMPLR ;
   d_arr_2_22 <= d_arr_24_0_EXMPLR ;
   d_arr_2_21 <= d_arr_24_0_EXMPLR ;
   d_arr_2_20 <= d_arr_24_0_EXMPLR ;
   d_arr_2_19 <= d_arr_24_0_EXMPLR ;
   d_arr_2_18 <= d_arr_24_0_EXMPLR ;
   d_arr_2_17 <= d_arr_24_0_EXMPLR ;
   d_arr_2_16 <= d_arr_24_0_EXMPLR ;
   d_arr_2_15 <= d_arr_24_0_EXMPLR ;
   d_arr_2_14 <= d_arr_24_0_EXMPLR ;
   d_arr_2_13 <= d_arr_24_0_EXMPLR ;
   d_arr_2_12 <= d_arr_24_0_EXMPLR ;
   d_arr_2_11 <= d_arr_24_0_EXMPLR ;
   d_arr_2_10 <= d_arr_24_0_EXMPLR ;
   d_arr_2_9 <= d_arr_24_0_EXMPLR ;
   d_arr_2_8 <= d_arr_24_0_EXMPLR ;
   d_arr_2_7 <= d_arr_24_0_EXMPLR ;
   d_arr_2_6 <= d_arr_24_0_EXMPLR ;
   d_arr_2_5 <= d_arr_24_0_EXMPLR ;
   d_arr_2_4 <= d_arr_24_0_EXMPLR ;
   d_arr_2_3 <= d_arr_24_0_EXMPLR ;
   d_arr_2_2 <= d_arr_24_0_EXMPLR ;
   d_arr_2_1 <= d_arr_24_0_EXMPLR ;
   d_arr_2_0 <= d_arr_24_0_EXMPLR ;
   d_arr_3_31 <= d_arr_24_0_EXMPLR ;
   d_arr_3_30 <= d_arr_24_0_EXMPLR ;
   d_arr_3_29 <= d_arr_24_0_EXMPLR ;
   d_arr_3_28 <= d_arr_24_0_EXMPLR ;
   d_arr_3_27 <= d_arr_24_0_EXMPLR ;
   d_arr_3_26 <= d_arr_24_0_EXMPLR ;
   d_arr_3_25 <= d_arr_24_0_EXMPLR ;
   d_arr_3_24 <= d_arr_24_0_EXMPLR ;
   d_arr_3_23 <= d_arr_24_0_EXMPLR ;
   d_arr_3_22 <= d_arr_24_0_EXMPLR ;
   d_arr_3_21 <= d_arr_24_0_EXMPLR ;
   d_arr_3_20 <= d_arr_24_0_EXMPLR ;
   d_arr_3_19 <= d_arr_24_0_EXMPLR ;
   d_arr_3_18 <= d_arr_24_0_EXMPLR ;
   d_arr_3_17 <= d_arr_24_0_EXMPLR ;
   d_arr_3_16 <= d_arr_24_0_EXMPLR ;
   d_arr_3_15 <= d_arr_24_0_EXMPLR ;
   d_arr_3_14 <= d_arr_24_0_EXMPLR ;
   d_arr_3_13 <= d_arr_24_0_EXMPLR ;
   d_arr_3_12 <= d_arr_24_0_EXMPLR ;
   d_arr_3_11 <= d_arr_24_0_EXMPLR ;
   d_arr_3_10 <= d_arr_24_0_EXMPLR ;
   d_arr_3_9 <= d_arr_24_0_EXMPLR ;
   d_arr_3_8 <= d_arr_24_0_EXMPLR ;
   d_arr_3_7 <= d_arr_24_0_EXMPLR ;
   d_arr_3_6 <= d_arr_24_0_EXMPLR ;
   d_arr_3_5 <= d_arr_24_0_EXMPLR ;
   d_arr_3_4 <= d_arr_24_0_EXMPLR ;
   d_arr_3_3 <= d_arr_24_0_EXMPLR ;
   d_arr_3_2 <= d_arr_24_0_EXMPLR ;
   d_arr_3_1 <= d_arr_24_0_EXMPLR ;
   d_arr_3_0 <= d_arr_24_0_EXMPLR ;
   d_arr_4_31 <= d_arr_24_0_EXMPLR ;
   d_arr_4_30 <= d_arr_24_0_EXMPLR ;
   d_arr_4_29 <= d_arr_24_0_EXMPLR ;
   d_arr_4_28 <= d_arr_24_0_EXMPLR ;
   d_arr_4_27 <= d_arr_24_0_EXMPLR ;
   d_arr_4_26 <= d_arr_24_0_EXMPLR ;
   d_arr_4_25 <= d_arr_24_0_EXMPLR ;
   d_arr_4_24 <= d_arr_24_0_EXMPLR ;
   d_arr_4_23 <= d_arr_24_0_EXMPLR ;
   d_arr_4_22 <= d_arr_24_0_EXMPLR ;
   d_arr_4_21 <= d_arr_24_0_EXMPLR ;
   d_arr_4_20 <= d_arr_24_0_EXMPLR ;
   d_arr_4_19 <= d_arr_24_0_EXMPLR ;
   d_arr_4_18 <= d_arr_24_0_EXMPLR ;
   d_arr_4_17 <= d_arr_24_0_EXMPLR ;
   d_arr_4_16 <= d_arr_24_0_EXMPLR ;
   d_arr_4_15 <= d_arr_24_0_EXMPLR ;
   d_arr_4_14 <= d_arr_24_0_EXMPLR ;
   d_arr_4_13 <= d_arr_24_0_EXMPLR ;
   d_arr_4_12 <= d_arr_24_0_EXMPLR ;
   d_arr_4_11 <= d_arr_24_0_EXMPLR ;
   d_arr_4_10 <= d_arr_24_0_EXMPLR ;
   d_arr_4_9 <= d_arr_24_0_EXMPLR ;
   d_arr_4_8 <= d_arr_24_0_EXMPLR ;
   d_arr_4_7 <= d_arr_24_0_EXMPLR ;
   d_arr_4_6 <= d_arr_24_0_EXMPLR ;
   d_arr_4_5 <= d_arr_24_0_EXMPLR ;
   d_arr_4_4 <= d_arr_24_0_EXMPLR ;
   d_arr_4_3 <= d_arr_24_0_EXMPLR ;
   d_arr_4_2 <= d_arr_24_0_EXMPLR ;
   d_arr_4_1 <= d_arr_24_0_EXMPLR ;
   d_arr_4_0 <= d_arr_24_0_EXMPLR ;
   d_arr_5_31 <= d_arr_24_0_EXMPLR ;
   d_arr_5_30 <= d_arr_24_0_EXMPLR ;
   d_arr_5_29 <= d_arr_24_0_EXMPLR ;
   d_arr_5_28 <= d_arr_24_0_EXMPLR ;
   d_arr_5_27 <= d_arr_24_0_EXMPLR ;
   d_arr_5_26 <= d_arr_24_0_EXMPLR ;
   d_arr_5_25 <= d_arr_24_0_EXMPLR ;
   d_arr_5_24 <= d_arr_24_0_EXMPLR ;
   d_arr_5_23 <= d_arr_24_0_EXMPLR ;
   d_arr_5_22 <= d_arr_24_0_EXMPLR ;
   d_arr_5_21 <= d_arr_24_0_EXMPLR ;
   d_arr_5_20 <= d_arr_24_0_EXMPLR ;
   d_arr_5_19 <= d_arr_24_0_EXMPLR ;
   d_arr_5_18 <= d_arr_24_0_EXMPLR ;
   d_arr_5_17 <= d_arr_24_0_EXMPLR ;
   d_arr_5_16 <= d_arr_24_0_EXMPLR ;
   d_arr_5_15 <= d_arr_24_0_EXMPLR ;
   d_arr_5_14 <= d_arr_24_0_EXMPLR ;
   d_arr_5_13 <= d_arr_24_0_EXMPLR ;
   d_arr_5_12 <= d_arr_24_0_EXMPLR ;
   d_arr_5_11 <= d_arr_24_0_EXMPLR ;
   d_arr_5_10 <= d_arr_24_0_EXMPLR ;
   d_arr_5_9 <= d_arr_24_0_EXMPLR ;
   d_arr_5_8 <= d_arr_24_0_EXMPLR ;
   d_arr_5_7 <= d_arr_24_0_EXMPLR ;
   d_arr_5_6 <= d_arr_24_0_EXMPLR ;
   d_arr_5_5 <= d_arr_24_0_EXMPLR ;
   d_arr_5_4 <= d_arr_24_0_EXMPLR ;
   d_arr_5_3 <= d_arr_24_0_EXMPLR ;
   d_arr_5_2 <= d_arr_24_0_EXMPLR ;
   d_arr_5_1 <= d_arr_24_0_EXMPLR ;
   d_arr_5_0 <= d_arr_24_0_EXMPLR ;
   d_arr_6_31 <= d_arr_24_0_EXMPLR ;
   d_arr_6_30 <= d_arr_24_0_EXMPLR ;
   d_arr_6_29 <= d_arr_24_0_EXMPLR ;
   d_arr_6_28 <= d_arr_24_0_EXMPLR ;
   d_arr_6_27 <= d_arr_24_0_EXMPLR ;
   d_arr_6_26 <= d_arr_24_0_EXMPLR ;
   d_arr_6_25 <= d_arr_24_0_EXMPLR ;
   d_arr_6_24 <= d_arr_24_0_EXMPLR ;
   d_arr_6_23 <= d_arr_24_0_EXMPLR ;
   d_arr_6_22 <= d_arr_24_0_EXMPLR ;
   d_arr_6_21 <= d_arr_24_0_EXMPLR ;
   d_arr_6_20 <= d_arr_24_0_EXMPLR ;
   d_arr_6_19 <= d_arr_24_0_EXMPLR ;
   d_arr_6_18 <= d_arr_24_0_EXMPLR ;
   d_arr_6_17 <= d_arr_24_0_EXMPLR ;
   d_arr_6_16 <= d_arr_24_0_EXMPLR ;
   d_arr_6_15 <= d_arr_24_0_EXMPLR ;
   d_arr_6_14 <= d_arr_24_0_EXMPLR ;
   d_arr_6_13 <= d_arr_24_0_EXMPLR ;
   d_arr_6_12 <= d_arr_24_0_EXMPLR ;
   d_arr_6_11 <= d_arr_24_0_EXMPLR ;
   d_arr_6_10 <= d_arr_24_0_EXMPLR ;
   d_arr_6_9 <= d_arr_24_0_EXMPLR ;
   d_arr_6_8 <= d_arr_24_0_EXMPLR ;
   d_arr_6_7 <= d_arr_24_0_EXMPLR ;
   d_arr_6_6 <= d_arr_24_0_EXMPLR ;
   d_arr_6_5 <= d_arr_24_0_EXMPLR ;
   d_arr_6_4 <= d_arr_24_0_EXMPLR ;
   d_arr_6_3 <= d_arr_24_0_EXMPLR ;
   d_arr_6_2 <= d_arr_24_0_EXMPLR ;
   d_arr_6_1 <= d_arr_24_0_EXMPLR ;
   d_arr_6_0 <= d_arr_24_0_EXMPLR ;
   d_arr_7_31 <= d_arr_24_0_EXMPLR ;
   d_arr_7_30 <= d_arr_24_0_EXMPLR ;
   d_arr_7_29 <= d_arr_24_0_EXMPLR ;
   d_arr_7_28 <= d_arr_24_0_EXMPLR ;
   d_arr_7_27 <= d_arr_24_0_EXMPLR ;
   d_arr_7_26 <= d_arr_24_0_EXMPLR ;
   d_arr_7_25 <= d_arr_24_0_EXMPLR ;
   d_arr_7_24 <= d_arr_24_0_EXMPLR ;
   d_arr_7_23 <= d_arr_24_0_EXMPLR ;
   d_arr_7_22 <= d_arr_24_0_EXMPLR ;
   d_arr_7_21 <= d_arr_24_0_EXMPLR ;
   d_arr_7_20 <= d_arr_24_0_EXMPLR ;
   d_arr_7_19 <= d_arr_24_0_EXMPLR ;
   d_arr_7_18 <= d_arr_24_0_EXMPLR ;
   d_arr_7_17 <= d_arr_24_0_EXMPLR ;
   d_arr_7_16 <= d_arr_24_0_EXMPLR ;
   d_arr_7_15 <= d_arr_24_0_EXMPLR ;
   d_arr_7_14 <= d_arr_24_0_EXMPLR ;
   d_arr_7_13 <= d_arr_24_0_EXMPLR ;
   d_arr_7_12 <= d_arr_24_0_EXMPLR ;
   d_arr_7_11 <= d_arr_24_0_EXMPLR ;
   d_arr_7_10 <= d_arr_24_0_EXMPLR ;
   d_arr_7_9 <= d_arr_24_0_EXMPLR ;
   d_arr_7_8 <= d_arr_24_0_EXMPLR ;
   d_arr_7_7 <= d_arr_24_0_EXMPLR ;
   d_arr_7_6 <= d_arr_24_0_EXMPLR ;
   d_arr_7_5 <= d_arr_24_0_EXMPLR ;
   d_arr_7_4 <= d_arr_24_0_EXMPLR ;
   d_arr_7_3 <= d_arr_24_0_EXMPLR ;
   d_arr_7_2 <= d_arr_24_0_EXMPLR ;
   d_arr_7_1 <= d_arr_24_0_EXMPLR ;
   d_arr_7_0 <= d_arr_24_0_EXMPLR ;
   d_arr_8_31 <= d_arr_24_0_EXMPLR ;
   d_arr_8_30 <= d_arr_24_0_EXMPLR ;
   d_arr_8_29 <= d_arr_24_0_EXMPLR ;
   d_arr_8_28 <= d_arr_24_0_EXMPLR ;
   d_arr_8_27 <= d_arr_24_0_EXMPLR ;
   d_arr_8_26 <= d_arr_24_0_EXMPLR ;
   d_arr_8_25 <= d_arr_24_0_EXMPLR ;
   d_arr_8_24 <= d_arr_24_0_EXMPLR ;
   d_arr_8_23 <= d_arr_24_0_EXMPLR ;
   d_arr_8_22 <= d_arr_24_0_EXMPLR ;
   d_arr_8_21 <= d_arr_24_0_EXMPLR ;
   d_arr_8_20 <= d_arr_24_0_EXMPLR ;
   d_arr_8_19 <= d_arr_24_0_EXMPLR ;
   d_arr_8_18 <= d_arr_24_0_EXMPLR ;
   d_arr_8_17 <= d_arr_24_0_EXMPLR ;
   d_arr_8_16 <= d_arr_24_0_EXMPLR ;
   d_arr_8_15 <= d_arr_24_0_EXMPLR ;
   d_arr_8_14 <= d_arr_24_0_EXMPLR ;
   d_arr_8_13 <= d_arr_24_0_EXMPLR ;
   d_arr_8_12 <= d_arr_24_0_EXMPLR ;
   d_arr_8_11 <= d_arr_24_0_EXMPLR ;
   d_arr_8_10 <= d_arr_24_0_EXMPLR ;
   d_arr_8_9 <= d_arr_24_0_EXMPLR ;
   d_arr_8_8 <= d_arr_24_0_EXMPLR ;
   d_arr_8_7 <= d_arr_24_0_EXMPLR ;
   d_arr_8_6 <= d_arr_24_0_EXMPLR ;
   d_arr_8_5 <= d_arr_24_0_EXMPLR ;
   d_arr_8_4 <= d_arr_24_0_EXMPLR ;
   d_arr_8_3 <= d_arr_24_0_EXMPLR ;
   d_arr_8_2 <= d_arr_24_0_EXMPLR ;
   d_arr_8_1 <= d_arr_24_0_EXMPLR ;
   d_arr_8_0 <= d_arr_24_0_EXMPLR ;
   d_arr_9_31 <= d_arr_24_0_EXMPLR ;
   d_arr_9_30 <= d_arr_24_0_EXMPLR ;
   d_arr_9_29 <= d_arr_24_0_EXMPLR ;
   d_arr_9_28 <= d_arr_24_0_EXMPLR ;
   d_arr_9_27 <= d_arr_24_0_EXMPLR ;
   d_arr_9_26 <= d_arr_24_0_EXMPLR ;
   d_arr_9_25 <= d_arr_24_0_EXMPLR ;
   d_arr_9_24 <= d_arr_24_0_EXMPLR ;
   d_arr_9_23 <= d_arr_24_0_EXMPLR ;
   d_arr_9_22 <= d_arr_24_0_EXMPLR ;
   d_arr_9_21 <= d_arr_24_0_EXMPLR ;
   d_arr_9_20 <= d_arr_24_0_EXMPLR ;
   d_arr_9_19 <= d_arr_24_0_EXMPLR ;
   d_arr_9_18 <= d_arr_24_0_EXMPLR ;
   d_arr_9_17 <= d_arr_24_0_EXMPLR ;
   d_arr_9_16 <= d_arr_24_0_EXMPLR ;
   d_arr_9_15 <= d_arr_24_0_EXMPLR ;
   d_arr_9_14 <= d_arr_24_0_EXMPLR ;
   d_arr_9_13 <= d_arr_24_0_EXMPLR ;
   d_arr_9_12 <= d_arr_24_0_EXMPLR ;
   d_arr_9_11 <= d_arr_24_0_EXMPLR ;
   d_arr_9_10 <= d_arr_24_0_EXMPLR ;
   d_arr_9_9 <= d_arr_24_0_EXMPLR ;
   d_arr_9_8 <= d_arr_24_0_EXMPLR ;
   d_arr_9_7 <= d_arr_24_0_EXMPLR ;
   d_arr_9_6 <= d_arr_24_0_EXMPLR ;
   d_arr_9_5 <= d_arr_24_0_EXMPLR ;
   d_arr_9_4 <= d_arr_24_0_EXMPLR ;
   d_arr_9_3 <= d_arr_24_0_EXMPLR ;
   d_arr_9_2 <= d_arr_24_0_EXMPLR ;
   d_arr_9_1 <= d_arr_24_0_EXMPLR ;
   d_arr_9_0 <= d_arr_24_0_EXMPLR ;
   d_arr_10_31 <= d_arr_24_0_EXMPLR ;
   d_arr_10_30 <= d_arr_24_0_EXMPLR ;
   d_arr_10_29 <= d_arr_24_0_EXMPLR ;
   d_arr_10_28 <= d_arr_24_0_EXMPLR ;
   d_arr_10_27 <= d_arr_24_0_EXMPLR ;
   d_arr_10_26 <= d_arr_24_0_EXMPLR ;
   d_arr_10_25 <= d_arr_24_0_EXMPLR ;
   d_arr_10_24 <= d_arr_24_0_EXMPLR ;
   d_arr_10_23 <= d_arr_24_0_EXMPLR ;
   d_arr_10_22 <= d_arr_24_0_EXMPLR ;
   d_arr_10_21 <= d_arr_24_0_EXMPLR ;
   d_arr_10_20 <= d_arr_24_0_EXMPLR ;
   d_arr_10_19 <= d_arr_24_0_EXMPLR ;
   d_arr_10_18 <= d_arr_24_0_EXMPLR ;
   d_arr_10_17 <= d_arr_24_0_EXMPLR ;
   d_arr_10_16 <= d_arr_24_0_EXMPLR ;
   d_arr_10_15 <= d_arr_24_0_EXMPLR ;
   d_arr_10_14 <= d_arr_24_0_EXMPLR ;
   d_arr_10_13 <= d_arr_24_0_EXMPLR ;
   d_arr_10_12 <= d_arr_24_0_EXMPLR ;
   d_arr_10_11 <= d_arr_24_0_EXMPLR ;
   d_arr_10_10 <= d_arr_24_0_EXMPLR ;
   d_arr_10_9 <= d_arr_24_0_EXMPLR ;
   d_arr_10_8 <= d_arr_24_0_EXMPLR ;
   d_arr_10_7 <= d_arr_24_0_EXMPLR ;
   d_arr_10_6 <= d_arr_24_0_EXMPLR ;
   d_arr_10_5 <= d_arr_24_0_EXMPLR ;
   d_arr_10_4 <= d_arr_24_0_EXMPLR ;
   d_arr_10_3 <= d_arr_24_0_EXMPLR ;
   d_arr_10_2 <= d_arr_24_0_EXMPLR ;
   d_arr_10_1 <= d_arr_24_0_EXMPLR ;
   d_arr_10_0 <= d_arr_24_0_EXMPLR ;
   d_arr_11_31 <= d_arr_24_0_EXMPLR ;
   d_arr_11_30 <= d_arr_24_0_EXMPLR ;
   d_arr_11_29 <= d_arr_24_0_EXMPLR ;
   d_arr_11_28 <= d_arr_24_0_EXMPLR ;
   d_arr_11_27 <= d_arr_24_0_EXMPLR ;
   d_arr_11_26 <= d_arr_24_0_EXMPLR ;
   d_arr_11_25 <= d_arr_24_0_EXMPLR ;
   d_arr_11_24 <= d_arr_24_0_EXMPLR ;
   d_arr_11_23 <= d_arr_24_0_EXMPLR ;
   d_arr_11_22 <= d_arr_24_0_EXMPLR ;
   d_arr_11_21 <= d_arr_24_0_EXMPLR ;
   d_arr_11_20 <= d_arr_24_0_EXMPLR ;
   d_arr_11_19 <= d_arr_24_0_EXMPLR ;
   d_arr_11_18 <= d_arr_24_0_EXMPLR ;
   d_arr_11_17 <= d_arr_24_0_EXMPLR ;
   d_arr_11_16 <= d_arr_24_0_EXMPLR ;
   d_arr_11_15 <= d_arr_24_0_EXMPLR ;
   d_arr_11_14 <= d_arr_24_0_EXMPLR ;
   d_arr_11_13 <= d_arr_24_0_EXMPLR ;
   d_arr_11_12 <= d_arr_24_0_EXMPLR ;
   d_arr_11_11 <= d_arr_24_0_EXMPLR ;
   d_arr_11_10 <= d_arr_24_0_EXMPLR ;
   d_arr_11_9 <= d_arr_24_0_EXMPLR ;
   d_arr_11_8 <= d_arr_24_0_EXMPLR ;
   d_arr_11_7 <= d_arr_24_0_EXMPLR ;
   d_arr_11_6 <= d_arr_24_0_EXMPLR ;
   d_arr_11_5 <= d_arr_24_0_EXMPLR ;
   d_arr_11_4 <= d_arr_24_0_EXMPLR ;
   d_arr_11_3 <= d_arr_24_0_EXMPLR ;
   d_arr_11_2 <= d_arr_24_0_EXMPLR ;
   d_arr_11_1 <= d_arr_24_0_EXMPLR ;
   d_arr_11_0 <= d_arr_24_0_EXMPLR ;
   d_arr_12_31 <= d_arr_24_0_EXMPLR ;
   d_arr_12_30 <= d_arr_24_0_EXMPLR ;
   d_arr_12_29 <= d_arr_24_0_EXMPLR ;
   d_arr_12_28 <= d_arr_24_0_EXMPLR ;
   d_arr_12_27 <= d_arr_24_0_EXMPLR ;
   d_arr_12_26 <= d_arr_24_0_EXMPLR ;
   d_arr_12_25 <= d_arr_24_0_EXMPLR ;
   d_arr_12_24 <= d_arr_24_0_EXMPLR ;
   d_arr_12_23 <= d_arr_24_0_EXMPLR ;
   d_arr_12_22 <= d_arr_24_0_EXMPLR ;
   d_arr_12_21 <= d_arr_24_0_EXMPLR ;
   d_arr_12_20 <= d_arr_24_0_EXMPLR ;
   d_arr_12_19 <= d_arr_24_0_EXMPLR ;
   d_arr_12_18 <= d_arr_24_0_EXMPLR ;
   d_arr_12_17 <= d_arr_24_0_EXMPLR ;
   d_arr_12_16 <= d_arr_24_0_EXMPLR ;
   d_arr_12_15 <= d_arr_24_0_EXMPLR ;
   d_arr_12_14 <= d_arr_24_0_EXMPLR ;
   d_arr_12_13 <= d_arr_24_0_EXMPLR ;
   d_arr_12_12 <= d_arr_24_0_EXMPLR ;
   d_arr_12_11 <= d_arr_24_0_EXMPLR ;
   d_arr_12_10 <= d_arr_24_0_EXMPLR ;
   d_arr_12_9 <= d_arr_24_0_EXMPLR ;
   d_arr_12_8 <= d_arr_24_0_EXMPLR ;
   d_arr_12_7 <= d_arr_24_0_EXMPLR ;
   d_arr_12_6 <= d_arr_24_0_EXMPLR ;
   d_arr_12_5 <= d_arr_24_0_EXMPLR ;
   d_arr_12_4 <= d_arr_24_0_EXMPLR ;
   d_arr_12_3 <= d_arr_24_0_EXMPLR ;
   d_arr_12_2 <= d_arr_24_0_EXMPLR ;
   d_arr_12_1 <= d_arr_24_0_EXMPLR ;
   d_arr_12_0 <= d_arr_24_0_EXMPLR ;
   d_arr_13_31 <= d_arr_24_0_EXMPLR ;
   d_arr_13_30 <= d_arr_24_0_EXMPLR ;
   d_arr_13_29 <= d_arr_24_0_EXMPLR ;
   d_arr_13_28 <= d_arr_24_0_EXMPLR ;
   d_arr_13_27 <= d_arr_24_0_EXMPLR ;
   d_arr_13_26 <= d_arr_24_0_EXMPLR ;
   d_arr_13_25 <= d_arr_24_0_EXMPLR ;
   d_arr_13_24 <= d_arr_24_0_EXMPLR ;
   d_arr_13_23 <= d_arr_24_0_EXMPLR ;
   d_arr_13_22 <= d_arr_24_0_EXMPLR ;
   d_arr_13_21 <= d_arr_24_0_EXMPLR ;
   d_arr_13_20 <= d_arr_24_0_EXMPLR ;
   d_arr_13_19 <= d_arr_24_0_EXMPLR ;
   d_arr_13_18 <= d_arr_24_0_EXMPLR ;
   d_arr_13_17 <= d_arr_24_0_EXMPLR ;
   d_arr_13_16 <= d_arr_24_0_EXMPLR ;
   d_arr_13_15 <= d_arr_24_0_EXMPLR ;
   d_arr_13_14 <= d_arr_24_0_EXMPLR ;
   d_arr_13_13 <= d_arr_24_0_EXMPLR ;
   d_arr_13_12 <= d_arr_24_0_EXMPLR ;
   d_arr_13_11 <= d_arr_24_0_EXMPLR ;
   d_arr_13_10 <= d_arr_24_0_EXMPLR ;
   d_arr_13_9 <= d_arr_24_0_EXMPLR ;
   d_arr_13_8 <= d_arr_24_0_EXMPLR ;
   d_arr_13_7 <= d_arr_24_0_EXMPLR ;
   d_arr_13_6 <= d_arr_24_0_EXMPLR ;
   d_arr_13_5 <= d_arr_24_0_EXMPLR ;
   d_arr_13_4 <= d_arr_24_0_EXMPLR ;
   d_arr_13_3 <= d_arr_24_0_EXMPLR ;
   d_arr_13_2 <= d_arr_24_0_EXMPLR ;
   d_arr_13_1 <= d_arr_24_0_EXMPLR ;
   d_arr_13_0 <= d_arr_24_0_EXMPLR ;
   d_arr_14_31 <= d_arr_24_0_EXMPLR ;
   d_arr_14_30 <= d_arr_24_0_EXMPLR ;
   d_arr_14_29 <= d_arr_24_0_EXMPLR ;
   d_arr_14_28 <= d_arr_24_0_EXMPLR ;
   d_arr_14_27 <= d_arr_24_0_EXMPLR ;
   d_arr_14_26 <= d_arr_24_0_EXMPLR ;
   d_arr_14_25 <= d_arr_24_0_EXMPLR ;
   d_arr_14_24 <= d_arr_24_0_EXMPLR ;
   d_arr_14_23 <= d_arr_24_0_EXMPLR ;
   d_arr_14_22 <= d_arr_24_0_EXMPLR ;
   d_arr_14_21 <= d_arr_24_0_EXMPLR ;
   d_arr_14_20 <= d_arr_24_0_EXMPLR ;
   d_arr_14_19 <= d_arr_24_0_EXMPLR ;
   d_arr_14_18 <= d_arr_24_0_EXMPLR ;
   d_arr_14_17 <= d_arr_24_0_EXMPLR ;
   d_arr_14_16 <= d_arr_24_0_EXMPLR ;
   d_arr_14_15 <= d_arr_24_0_EXMPLR ;
   d_arr_14_14 <= d_arr_24_0_EXMPLR ;
   d_arr_14_13 <= d_arr_24_0_EXMPLR ;
   d_arr_14_12 <= d_arr_24_0_EXMPLR ;
   d_arr_14_11 <= d_arr_24_0_EXMPLR ;
   d_arr_14_10 <= d_arr_24_0_EXMPLR ;
   d_arr_14_9 <= d_arr_24_0_EXMPLR ;
   d_arr_14_8 <= d_arr_24_0_EXMPLR ;
   d_arr_14_7 <= d_arr_24_0_EXMPLR ;
   d_arr_14_6 <= d_arr_24_0_EXMPLR ;
   d_arr_14_5 <= d_arr_24_0_EXMPLR ;
   d_arr_14_4 <= d_arr_24_0_EXMPLR ;
   d_arr_14_3 <= d_arr_24_0_EXMPLR ;
   d_arr_14_2 <= d_arr_24_0_EXMPLR ;
   d_arr_14_1 <= d_arr_24_0_EXMPLR ;
   d_arr_14_0 <= d_arr_24_0_EXMPLR ;
   d_arr_15_31 <= d_arr_24_0_EXMPLR ;
   d_arr_15_30 <= d_arr_24_0_EXMPLR ;
   d_arr_15_29 <= d_arr_24_0_EXMPLR ;
   d_arr_15_28 <= d_arr_24_0_EXMPLR ;
   d_arr_15_27 <= d_arr_24_0_EXMPLR ;
   d_arr_15_26 <= d_arr_24_0_EXMPLR ;
   d_arr_15_25 <= d_arr_24_0_EXMPLR ;
   d_arr_15_24 <= d_arr_24_0_EXMPLR ;
   d_arr_15_23 <= d_arr_24_0_EXMPLR ;
   d_arr_15_22 <= d_arr_24_0_EXMPLR ;
   d_arr_15_21 <= d_arr_24_0_EXMPLR ;
   d_arr_15_20 <= d_arr_24_0_EXMPLR ;
   d_arr_15_19 <= d_arr_24_0_EXMPLR ;
   d_arr_15_18 <= d_arr_24_0_EXMPLR ;
   d_arr_15_17 <= d_arr_24_0_EXMPLR ;
   d_arr_15_16 <= d_arr_24_0_EXMPLR ;
   d_arr_15_15 <= d_arr_24_0_EXMPLR ;
   d_arr_15_14 <= d_arr_24_0_EXMPLR ;
   d_arr_15_13 <= d_arr_24_0_EXMPLR ;
   d_arr_15_12 <= d_arr_24_0_EXMPLR ;
   d_arr_15_11 <= d_arr_24_0_EXMPLR ;
   d_arr_15_10 <= d_arr_24_0_EXMPLR ;
   d_arr_15_9 <= d_arr_24_0_EXMPLR ;
   d_arr_15_8 <= d_arr_24_0_EXMPLR ;
   d_arr_15_7 <= d_arr_24_0_EXMPLR ;
   d_arr_15_6 <= d_arr_24_0_EXMPLR ;
   d_arr_15_5 <= d_arr_24_0_EXMPLR ;
   d_arr_15_4 <= d_arr_24_0_EXMPLR ;
   d_arr_15_3 <= d_arr_24_0_EXMPLR ;
   d_arr_15_2 <= d_arr_24_0_EXMPLR ;
   d_arr_15_1 <= d_arr_24_0_EXMPLR ;
   d_arr_15_0 <= d_arr_24_0_EXMPLR ;
   d_arr_16_31 <= d_arr_24_0_EXMPLR ;
   d_arr_16_30 <= d_arr_24_0_EXMPLR ;
   d_arr_16_29 <= d_arr_24_0_EXMPLR ;
   d_arr_16_28 <= d_arr_24_0_EXMPLR ;
   d_arr_16_27 <= d_arr_24_0_EXMPLR ;
   d_arr_16_26 <= d_arr_24_0_EXMPLR ;
   d_arr_16_25 <= d_arr_24_0_EXMPLR ;
   d_arr_16_24 <= d_arr_24_0_EXMPLR ;
   d_arr_16_23 <= d_arr_24_0_EXMPLR ;
   d_arr_16_22 <= d_arr_24_0_EXMPLR ;
   d_arr_16_21 <= d_arr_24_0_EXMPLR ;
   d_arr_16_20 <= d_arr_24_0_EXMPLR ;
   d_arr_16_19 <= d_arr_24_0_EXMPLR ;
   d_arr_16_18 <= d_arr_24_0_EXMPLR ;
   d_arr_16_17 <= d_arr_24_0_EXMPLR ;
   d_arr_16_16 <= d_arr_24_0_EXMPLR ;
   d_arr_16_15 <= d_arr_24_0_EXMPLR ;
   d_arr_16_14 <= d_arr_24_0_EXMPLR ;
   d_arr_16_13 <= d_arr_24_0_EXMPLR ;
   d_arr_16_12 <= d_arr_24_0_EXMPLR ;
   d_arr_16_11 <= d_arr_24_0_EXMPLR ;
   d_arr_16_10 <= d_arr_24_0_EXMPLR ;
   d_arr_16_9 <= d_arr_24_0_EXMPLR ;
   d_arr_16_8 <= d_arr_24_0_EXMPLR ;
   d_arr_16_7 <= d_arr_24_0_EXMPLR ;
   d_arr_16_6 <= d_arr_24_0_EXMPLR ;
   d_arr_16_5 <= d_arr_24_0_EXMPLR ;
   d_arr_16_4 <= d_arr_24_0_EXMPLR ;
   d_arr_16_3 <= d_arr_24_0_EXMPLR ;
   d_arr_16_2 <= d_arr_24_0_EXMPLR ;
   d_arr_16_1 <= d_arr_24_0_EXMPLR ;
   d_arr_16_0 <= d_arr_24_0_EXMPLR ;
   d_arr_17_31 <= d_arr_24_0_EXMPLR ;
   d_arr_17_30 <= d_arr_24_0_EXMPLR ;
   d_arr_17_29 <= d_arr_24_0_EXMPLR ;
   d_arr_17_28 <= d_arr_24_0_EXMPLR ;
   d_arr_17_27 <= d_arr_24_0_EXMPLR ;
   d_arr_17_26 <= d_arr_24_0_EXMPLR ;
   d_arr_17_25 <= d_arr_24_0_EXMPLR ;
   d_arr_17_24 <= d_arr_24_0_EXMPLR ;
   d_arr_17_23 <= d_arr_24_0_EXMPLR ;
   d_arr_17_22 <= d_arr_24_0_EXMPLR ;
   d_arr_17_21 <= d_arr_24_0_EXMPLR ;
   d_arr_17_20 <= d_arr_24_0_EXMPLR ;
   d_arr_17_19 <= d_arr_24_0_EXMPLR ;
   d_arr_17_18 <= d_arr_24_0_EXMPLR ;
   d_arr_17_17 <= d_arr_24_0_EXMPLR ;
   d_arr_17_16 <= d_arr_24_0_EXMPLR ;
   d_arr_17_15 <= d_arr_24_0_EXMPLR ;
   d_arr_17_14 <= d_arr_24_0_EXMPLR ;
   d_arr_17_13 <= d_arr_24_0_EXMPLR ;
   d_arr_17_12 <= d_arr_24_0_EXMPLR ;
   d_arr_17_11 <= d_arr_24_0_EXMPLR ;
   d_arr_17_10 <= d_arr_24_0_EXMPLR ;
   d_arr_17_9 <= d_arr_24_0_EXMPLR ;
   d_arr_17_8 <= d_arr_24_0_EXMPLR ;
   d_arr_17_7 <= d_arr_24_0_EXMPLR ;
   d_arr_17_6 <= d_arr_24_0_EXMPLR ;
   d_arr_17_5 <= d_arr_24_0_EXMPLR ;
   d_arr_17_4 <= d_arr_24_0_EXMPLR ;
   d_arr_17_3 <= d_arr_24_0_EXMPLR ;
   d_arr_17_2 <= d_arr_24_0_EXMPLR ;
   d_arr_17_1 <= d_arr_24_0_EXMPLR ;
   d_arr_17_0 <= d_arr_24_0_EXMPLR ;
   d_arr_18_31 <= d_arr_24_0_EXMPLR ;
   d_arr_18_30 <= d_arr_24_0_EXMPLR ;
   d_arr_18_29 <= d_arr_24_0_EXMPLR ;
   d_arr_18_28 <= d_arr_24_0_EXMPLR ;
   d_arr_18_27 <= d_arr_24_0_EXMPLR ;
   d_arr_18_26 <= d_arr_24_0_EXMPLR ;
   d_arr_18_25 <= d_arr_24_0_EXMPLR ;
   d_arr_18_24 <= d_arr_24_0_EXMPLR ;
   d_arr_18_23 <= d_arr_24_0_EXMPLR ;
   d_arr_18_22 <= d_arr_24_0_EXMPLR ;
   d_arr_18_21 <= d_arr_24_0_EXMPLR ;
   d_arr_18_20 <= d_arr_24_0_EXMPLR ;
   d_arr_18_19 <= d_arr_24_0_EXMPLR ;
   d_arr_18_18 <= d_arr_24_0_EXMPLR ;
   d_arr_18_17 <= d_arr_24_0_EXMPLR ;
   d_arr_18_16 <= d_arr_24_0_EXMPLR ;
   d_arr_18_15 <= d_arr_24_0_EXMPLR ;
   d_arr_18_14 <= d_arr_24_0_EXMPLR ;
   d_arr_18_13 <= d_arr_24_0_EXMPLR ;
   d_arr_18_12 <= d_arr_24_0_EXMPLR ;
   d_arr_18_11 <= d_arr_24_0_EXMPLR ;
   d_arr_18_10 <= d_arr_24_0_EXMPLR ;
   d_arr_18_9 <= d_arr_24_0_EXMPLR ;
   d_arr_18_8 <= d_arr_24_0_EXMPLR ;
   d_arr_18_7 <= d_arr_24_0_EXMPLR ;
   d_arr_18_6 <= d_arr_24_0_EXMPLR ;
   d_arr_18_5 <= d_arr_24_0_EXMPLR ;
   d_arr_18_4 <= d_arr_24_0_EXMPLR ;
   d_arr_18_3 <= d_arr_24_0_EXMPLR ;
   d_arr_18_2 <= d_arr_24_0_EXMPLR ;
   d_arr_18_1 <= d_arr_24_0_EXMPLR ;
   d_arr_18_0 <= d_arr_24_0_EXMPLR ;
   d_arr_19_31 <= d_arr_24_0_EXMPLR ;
   d_arr_19_30 <= d_arr_24_0_EXMPLR ;
   d_arr_19_29 <= d_arr_24_0_EXMPLR ;
   d_arr_19_28 <= d_arr_24_0_EXMPLR ;
   d_arr_19_27 <= d_arr_24_0_EXMPLR ;
   d_arr_19_26 <= d_arr_24_0_EXMPLR ;
   d_arr_19_25 <= d_arr_24_0_EXMPLR ;
   d_arr_19_24 <= d_arr_24_0_EXMPLR ;
   d_arr_19_23 <= d_arr_24_0_EXMPLR ;
   d_arr_19_22 <= d_arr_24_0_EXMPLR ;
   d_arr_19_21 <= d_arr_24_0_EXMPLR ;
   d_arr_19_20 <= d_arr_24_0_EXMPLR ;
   d_arr_19_19 <= d_arr_24_0_EXMPLR ;
   d_arr_19_18 <= d_arr_24_0_EXMPLR ;
   d_arr_19_17 <= d_arr_24_0_EXMPLR ;
   d_arr_19_16 <= d_arr_24_0_EXMPLR ;
   d_arr_19_15 <= d_arr_24_0_EXMPLR ;
   d_arr_19_14 <= d_arr_24_0_EXMPLR ;
   d_arr_19_13 <= d_arr_24_0_EXMPLR ;
   d_arr_19_12 <= d_arr_24_0_EXMPLR ;
   d_arr_19_11 <= d_arr_24_0_EXMPLR ;
   d_arr_19_10 <= d_arr_24_0_EXMPLR ;
   d_arr_19_9 <= d_arr_24_0_EXMPLR ;
   d_arr_19_8 <= d_arr_24_0_EXMPLR ;
   d_arr_19_7 <= d_arr_24_0_EXMPLR ;
   d_arr_19_6 <= d_arr_24_0_EXMPLR ;
   d_arr_19_5 <= d_arr_24_0_EXMPLR ;
   d_arr_19_4 <= d_arr_24_0_EXMPLR ;
   d_arr_19_3 <= d_arr_24_0_EXMPLR ;
   d_arr_19_2 <= d_arr_24_0_EXMPLR ;
   d_arr_19_1 <= d_arr_24_0_EXMPLR ;
   d_arr_19_0 <= d_arr_24_0_EXMPLR ;
   d_arr_20_31 <= d_arr_24_0_EXMPLR ;
   d_arr_20_30 <= d_arr_24_0_EXMPLR ;
   d_arr_20_29 <= d_arr_24_0_EXMPLR ;
   d_arr_20_28 <= d_arr_24_0_EXMPLR ;
   d_arr_20_27 <= d_arr_24_0_EXMPLR ;
   d_arr_20_26 <= d_arr_24_0_EXMPLR ;
   d_arr_20_25 <= d_arr_24_0_EXMPLR ;
   d_arr_20_24 <= d_arr_24_0_EXMPLR ;
   d_arr_20_23 <= d_arr_24_0_EXMPLR ;
   d_arr_20_22 <= d_arr_24_0_EXMPLR ;
   d_arr_20_21 <= d_arr_24_0_EXMPLR ;
   d_arr_20_20 <= d_arr_24_0_EXMPLR ;
   d_arr_20_19 <= d_arr_24_0_EXMPLR ;
   d_arr_20_18 <= d_arr_24_0_EXMPLR ;
   d_arr_20_17 <= d_arr_24_0_EXMPLR ;
   d_arr_20_16 <= d_arr_24_0_EXMPLR ;
   d_arr_20_15 <= d_arr_24_0_EXMPLR ;
   d_arr_20_14 <= d_arr_24_0_EXMPLR ;
   d_arr_20_13 <= d_arr_24_0_EXMPLR ;
   d_arr_20_12 <= d_arr_24_0_EXMPLR ;
   d_arr_20_11 <= d_arr_24_0_EXMPLR ;
   d_arr_20_10 <= d_arr_24_0_EXMPLR ;
   d_arr_20_9 <= d_arr_24_0_EXMPLR ;
   d_arr_20_8 <= d_arr_24_0_EXMPLR ;
   d_arr_20_7 <= d_arr_24_0_EXMPLR ;
   d_arr_20_6 <= d_arr_24_0_EXMPLR ;
   d_arr_20_5 <= d_arr_24_0_EXMPLR ;
   d_arr_20_4 <= d_arr_24_0_EXMPLR ;
   d_arr_20_3 <= d_arr_24_0_EXMPLR ;
   d_arr_20_2 <= d_arr_24_0_EXMPLR ;
   d_arr_20_1 <= d_arr_24_0_EXMPLR ;
   d_arr_20_0 <= d_arr_24_0_EXMPLR ;
   d_arr_21_31 <= d_arr_24_0_EXMPLR ;
   d_arr_21_30 <= d_arr_24_0_EXMPLR ;
   d_arr_21_29 <= d_arr_24_0_EXMPLR ;
   d_arr_21_28 <= d_arr_24_0_EXMPLR ;
   d_arr_21_27 <= d_arr_24_0_EXMPLR ;
   d_arr_21_26 <= d_arr_24_0_EXMPLR ;
   d_arr_21_25 <= d_arr_24_0_EXMPLR ;
   d_arr_21_24 <= d_arr_24_0_EXMPLR ;
   d_arr_21_23 <= d_arr_24_0_EXMPLR ;
   d_arr_21_22 <= d_arr_24_0_EXMPLR ;
   d_arr_21_21 <= d_arr_24_0_EXMPLR ;
   d_arr_21_20 <= d_arr_24_0_EXMPLR ;
   d_arr_21_19 <= d_arr_24_0_EXMPLR ;
   d_arr_21_18 <= d_arr_24_0_EXMPLR ;
   d_arr_21_17 <= d_arr_24_0_EXMPLR ;
   d_arr_21_16 <= d_arr_24_0_EXMPLR ;
   d_arr_21_15 <= d_arr_24_0_EXMPLR ;
   d_arr_21_14 <= d_arr_24_0_EXMPLR ;
   d_arr_21_13 <= d_arr_24_0_EXMPLR ;
   d_arr_21_12 <= d_arr_24_0_EXMPLR ;
   d_arr_21_11 <= d_arr_24_0_EXMPLR ;
   d_arr_21_10 <= d_arr_24_0_EXMPLR ;
   d_arr_21_9 <= d_arr_24_0_EXMPLR ;
   d_arr_21_8 <= d_arr_24_0_EXMPLR ;
   d_arr_21_7 <= d_arr_24_0_EXMPLR ;
   d_arr_21_6 <= d_arr_24_0_EXMPLR ;
   d_arr_21_5 <= d_arr_24_0_EXMPLR ;
   d_arr_21_4 <= d_arr_24_0_EXMPLR ;
   d_arr_21_3 <= d_arr_24_0_EXMPLR ;
   d_arr_21_2 <= d_arr_24_0_EXMPLR ;
   d_arr_21_1 <= d_arr_24_0_EXMPLR ;
   d_arr_21_0 <= d_arr_24_0_EXMPLR ;
   d_arr_22_31 <= d_arr_24_0_EXMPLR ;
   d_arr_22_30 <= d_arr_24_0_EXMPLR ;
   d_arr_22_29 <= d_arr_24_0_EXMPLR ;
   d_arr_22_28 <= d_arr_24_0_EXMPLR ;
   d_arr_22_27 <= d_arr_24_0_EXMPLR ;
   d_arr_22_26 <= d_arr_24_0_EXMPLR ;
   d_arr_22_25 <= d_arr_24_0_EXMPLR ;
   d_arr_22_24 <= d_arr_24_0_EXMPLR ;
   d_arr_22_23 <= d_arr_24_0_EXMPLR ;
   d_arr_22_22 <= d_arr_24_0_EXMPLR ;
   d_arr_22_21 <= d_arr_24_0_EXMPLR ;
   d_arr_22_20 <= d_arr_24_0_EXMPLR ;
   d_arr_22_19 <= d_arr_24_0_EXMPLR ;
   d_arr_22_18 <= d_arr_24_0_EXMPLR ;
   d_arr_22_17 <= d_arr_24_0_EXMPLR ;
   d_arr_22_16 <= d_arr_24_0_EXMPLR ;
   d_arr_22_15 <= d_arr_24_0_EXMPLR ;
   d_arr_22_14 <= d_arr_24_0_EXMPLR ;
   d_arr_22_13 <= d_arr_24_0_EXMPLR ;
   d_arr_22_12 <= d_arr_24_0_EXMPLR ;
   d_arr_22_11 <= d_arr_24_0_EXMPLR ;
   d_arr_22_10 <= d_arr_24_0_EXMPLR ;
   d_arr_22_9 <= d_arr_24_0_EXMPLR ;
   d_arr_22_8 <= d_arr_24_0_EXMPLR ;
   d_arr_22_7 <= d_arr_24_0_EXMPLR ;
   d_arr_22_6 <= d_arr_24_0_EXMPLR ;
   d_arr_22_5 <= d_arr_24_0_EXMPLR ;
   d_arr_22_4 <= d_arr_24_0_EXMPLR ;
   d_arr_22_3 <= d_arr_24_0_EXMPLR ;
   d_arr_22_2 <= d_arr_24_0_EXMPLR ;
   d_arr_22_1 <= d_arr_24_0_EXMPLR ;
   d_arr_22_0 <= d_arr_24_0_EXMPLR ;
   d_arr_23_31 <= d_arr_24_0_EXMPLR ;
   d_arr_23_30 <= d_arr_24_0_EXMPLR ;
   d_arr_23_29 <= d_arr_24_0_EXMPLR ;
   d_arr_23_28 <= d_arr_24_0_EXMPLR ;
   d_arr_23_27 <= d_arr_24_0_EXMPLR ;
   d_arr_23_26 <= d_arr_24_0_EXMPLR ;
   d_arr_23_25 <= d_arr_24_0_EXMPLR ;
   d_arr_23_24 <= d_arr_24_0_EXMPLR ;
   d_arr_23_23 <= d_arr_24_0_EXMPLR ;
   d_arr_23_22 <= d_arr_24_0_EXMPLR ;
   d_arr_23_21 <= d_arr_24_0_EXMPLR ;
   d_arr_23_20 <= d_arr_24_0_EXMPLR ;
   d_arr_23_19 <= d_arr_24_0_EXMPLR ;
   d_arr_23_18 <= d_arr_24_0_EXMPLR ;
   d_arr_23_17 <= d_arr_24_0_EXMPLR ;
   d_arr_23_16 <= d_arr_24_0_EXMPLR ;
   d_arr_23_15 <= d_arr_24_0_EXMPLR ;
   d_arr_23_14 <= d_arr_24_0_EXMPLR ;
   d_arr_23_13 <= d_arr_24_0_EXMPLR ;
   d_arr_23_12 <= d_arr_24_0_EXMPLR ;
   d_arr_23_11 <= d_arr_24_0_EXMPLR ;
   d_arr_23_10 <= d_arr_24_0_EXMPLR ;
   d_arr_23_9 <= d_arr_24_0_EXMPLR ;
   d_arr_23_8 <= d_arr_24_0_EXMPLR ;
   d_arr_23_7 <= d_arr_24_0_EXMPLR ;
   d_arr_23_6 <= d_arr_24_0_EXMPLR ;
   d_arr_23_5 <= d_arr_24_0_EXMPLR ;
   d_arr_23_4 <= d_arr_24_0_EXMPLR ;
   d_arr_23_3 <= d_arr_24_0_EXMPLR ;
   d_arr_23_2 <= d_arr_24_0_EXMPLR ;
   d_arr_23_1 <= d_arr_24_0_EXMPLR ;
   d_arr_23_0 <= d_arr_24_0_EXMPLR ;
   d_arr_24_31 <= d_arr_24_0_EXMPLR ;
   d_arr_24_30 <= d_arr_24_0_EXMPLR ;
   d_arr_24_29 <= d_arr_24_0_EXMPLR ;
   d_arr_24_28 <= d_arr_24_0_EXMPLR ;
   d_arr_24_27 <= d_arr_24_0_EXMPLR ;
   d_arr_24_26 <= d_arr_24_0_EXMPLR ;
   d_arr_24_25 <= d_arr_24_0_EXMPLR ;
   d_arr_24_24 <= d_arr_24_0_EXMPLR ;
   d_arr_24_23 <= d_arr_24_0_EXMPLR ;
   d_arr_24_22 <= d_arr_24_0_EXMPLR ;
   d_arr_24_21 <= d_arr_24_0_EXMPLR ;
   d_arr_24_20 <= d_arr_24_0_EXMPLR ;
   d_arr_24_19 <= d_arr_24_0_EXMPLR ;
   d_arr_24_18 <= d_arr_24_0_EXMPLR ;
   d_arr_24_17 <= d_arr_24_0_EXMPLR ;
   d_arr_24_16 <= d_arr_24_0_EXMPLR ;
   d_arr_24_15 <= d_arr_24_0_EXMPLR ;
   d_arr_24_14 <= d_arr_24_0_EXMPLR ;
   d_arr_24_13 <= d_arr_24_0_EXMPLR ;
   d_arr_24_12 <= d_arr_24_0_EXMPLR ;
   d_arr_24_11 <= d_arr_24_0_EXMPLR ;
   d_arr_24_10 <= d_arr_24_0_EXMPLR ;
   d_arr_24_9 <= d_arr_24_0_EXMPLR ;
   d_arr_24_8 <= d_arr_24_0_EXMPLR ;
   d_arr_24_7 <= d_arr_24_0_EXMPLR ;
   d_arr_24_6 <= d_arr_24_0_EXMPLR ;
   d_arr_24_5 <= d_arr_24_0_EXMPLR ;
   d_arr_24_4 <= d_arr_24_0_EXMPLR ;
   d_arr_24_3 <= d_arr_24_0_EXMPLR ;
   d_arr_24_2 <= d_arr_24_0_EXMPLR ;
   d_arr_24_1 <= d_arr_24_0_EXMPLR ;
   d_arr_24_0 <= d_arr_24_0_EXMPLR ;
   adder1_gen : NAdder_32 port map ( a(31)=>q_arr_9_31, a(30)=>q_arr_9_30, 
      a(29)=>q_arr_9_29, a(28)=>q_arr_9_28, a(27)=>nx550, a(26)=>q_arr_9_26, 
      a(25)=>q_arr_9_25, a(24)=>nx555, a(23)=>q_arr_9_23, a(22)=>q_arr_9_22, 
      a(21)=>q_arr_9_21, a(20)=>q_arr_9_20, a(19)=>q_arr_9_19, a(18)=>
      q_arr_9_18, a(17)=>q_arr_9_17, a(16)=>q_arr_9_16, a(15)=>q_arr_9_15, 
      a(14)=>q_arr_9_14, a(13)=>q_arr_9_13, a(12)=>q_arr_9_12, a(11)=>
      q_arr_9_11, a(10)=>q_arr_9_10, a(9)=>q_arr_9_9, a(8)=>q_arr_9_8, a(7)
      =>q_arr_9_7, a(6)=>q_arr_9_6, a(5)=>q_arr_9_5, a(4)=>q_arr_9_4, a(3)=>
      q_arr_9_3, a(2)=>q_arr_9_2, a(1)=>q_arr_9_1, a(0)=>q_arr_9_0, b(31)=>
      q_arr_18_31, b(30)=>q_arr_18_30, b(29)=>q_arr_18_29, b(28)=>
      q_arr_18_28, b(27)=>q_arr_18_27, b(26)=>q_arr_18_26, b(25)=>
      q_arr_18_25, b(24)=>q_arr_18_24, b(23)=>q_arr_18_23, b(22)=>
      q_arr_18_22, b(21)=>q_arr_18_21, b(20)=>q_arr_18_20, b(19)=>
      q_arr_18_19, b(18)=>q_arr_18_18, b(17)=>q_arr_18_17, b(16)=>
      q_arr_18_16, b(15)=>q_arr_18_15, b(14)=>q_arr_18_14, b(13)=>
      q_arr_18_13, b(12)=>q_arr_18_12, b(11)=>q_arr_18_11, b(10)=>
      q_arr_18_10, b(9)=>q_arr_18_9, b(8)=>q_arr_18_8, b(7)=>q_arr_18_7, 
      b(6)=>q_arr_18_6, b(5)=>q_arr_18_5, b(4)=>q_arr_18_4, b(3)=>q_arr_18_3, 
      b(2)=>q_arr_18_2, b(1)=>q_arr_18_1, b(0)=>q_arr_18_0, cin=>
      d_arr_24_0_EXMPLR, s(31)=>s1_31, s(30)=>s1_30, s(29)=>s1_29, s(28)=>
      s1_28, s(27)=>s1_27, s(26)=>s1_26, s(25)=>s1_25, s(24)=>s1_24, s(23)=>
      s1_23, s(22)=>s1_22, s(21)=>s1_21, s(20)=>s1_20, s(19)=>s1_19, s(18)=>
      s1_18, s(17)=>s1_17, s(16)=>s1_16, s(15)=>s1_15, s(14)=>s1_14, s(13)=>
      s1_13, s(12)=>s1_12, s(11)=>s1_11, s(10)=>s1_10, s(9)=>s1_9, s(8)=>
      s1_8, s(7)=>s1_7, s(6)=>s1_6, s(5)=>s1_5, s(4)=>s1_4, s(3)=>s1_3, s(2)
      =>s1_2, s(1)=>s1_1, s(0)=>s1_0, cout=>DANGLING(0));
   adder2_gen : NAdder_32 port map ( a(31)=>q_arr_0_31, a(30)=>q_arr_0_30, 
      a(29)=>q_arr_0_29, a(28)=>q_arr_0_28, a(27)=>q_arr_0_27, a(26)=>
      q_arr_0_26, a(25)=>q_arr_0_25, a(24)=>q_arr_0_24, a(23)=>q_arr_0_23, 
      a(22)=>q_arr_0_22, a(21)=>q_arr_0_21, a(20)=>q_arr_0_20, a(19)=>
      q_arr_0_19, a(18)=>q_arr_0_18, a(17)=>q_arr_0_17, a(16)=>q_arr_0_16, 
      a(15)=>q_arr_0_15, a(14)=>q_arr_0_14, a(13)=>q_arr_0_13, a(12)=>
      q_arr_0_12, a(11)=>q_arr_0_11, a(10)=>q_arr_0_10, a(9)=>q_arr_0_9, 
      a(8)=>q_arr_0_8, a(7)=>q_arr_0_7, a(6)=>q_arr_0_6, a(5)=>q_arr_0_5, 
      a(4)=>q_arr_0_4, a(3)=>q_arr_0_3, a(2)=>q_arr_0_2, a(1)=>q_arr_0_1, 
      a(0)=>q_arr_0_0, b(31)=>s1_31, b(30)=>s1_30, b(29)=>s1_29, b(28)=>
      s1_28, b(27)=>s1_27, b(26)=>s1_26, b(25)=>s1_25, b(24)=>s1_24, b(23)=>
      s1_23, b(22)=>s1_22, b(21)=>s1_21, b(20)=>s1_20, b(19)=>s1_19, b(18)=>
      s1_18, b(17)=>s1_17, b(16)=>s1_16, b(15)=>s1_15, b(14)=>s1_14, b(13)=>
      s1_13, b(12)=>s1_12, b(11)=>s1_11, b(10)=>s1_10, b(9)=>s1_9, b(8)=>
      s1_8, b(7)=>s1_7, b(6)=>s1_6, b(5)=>s1_5, b(4)=>s1_4, b(3)=>s1_3, b(2)
      =>s1_2, b(1)=>s1_1, b(0)=>s1_0, cin=>d_arr_24_0_EXMPLR, s(31)=>s2_31, 
      s(30)=>s2_30, s(29)=>s2_29, s(28)=>s2_28, s(27)=>s2_27, s(26)=>s2_26, 
      s(25)=>s2_25, s(24)=>s2_24, s(23)=>s2_23, s(22)=>s2_22, s(21)=>s2_21, 
      s(20)=>s2_20, s(19)=>s2_19, s(18)=>s2_18, s(17)=>s2_17, s(16)=>s2_16, 
      s(15)=>s2_15, s(14)=>s2_14, s(13)=>s2_13, s(12)=>s2_12, s(11)=>s2_11, 
      s(10)=>s2_10, s(9)=>s2_9, s(8)=>s2_8, s(7)=>s2_7, s(6)=>s2_6, s(5)=>
      s2_5, s(4)=>s2_4, s(3)=>s2_3, s(2)=>s2_2, s(1)=>s2_1, s(0)=>s2_0, cout
      =>DANGLING(1));
   ix41 : fake_gnd port map ( Y=>d_arr_24_0_EXMPLR);
   ix17 : inv01 port map ( Y=>d_arr_1_0, A=>nx153);
   ix154 : aoi222 port map ( Y=>nx153, A0=>q_arr_9_0, A1=>nx521, B0=>
      q_arr_9_5, B1=>nx460, C0=>q_arr_9_3, C1=>nx479);
   ix29 : inv01 port map ( Y=>d_arr_1_1, A=>nx165);
   ix166 : aoi222 port map ( Y=>nx165, A0=>q_arr_9_1, A1=>nx521, B0=>
      q_arr_9_6, B1=>nx460, C0=>q_arr_9_4, C1=>nx479);
   ix43 : inv01 port map ( Y=>d_arr_1_2, A=>nx169);
   ix170 : aoi222 port map ( Y=>nx169, A0=>q_arr_9_2, A1=>nx521, B0=>
      q_arr_9_7, B1=>nx460, C0=>q_arr_9_5, C1=>nx479);
   ix53 : inv01 port map ( Y=>d_arr_1_3, A=>nx173);
   ix174 : aoi222 port map ( Y=>nx173, A0=>q_arr_9_3, A1=>nx521, B0=>
      q_arr_9_8, B1=>nx460, C0=>q_arr_9_6, C1=>nx479);
   ix65 : inv01 port map ( Y=>d_arr_1_4, A=>nx177);
   ix178 : aoi222 port map ( Y=>nx177, A0=>q_arr_9_4, A1=>nx521, B0=>
      q_arr_9_9, B1=>nx460, C0=>q_arr_9_7, C1=>nx479);
   ix77 : inv01 port map ( Y=>d_arr_1_5, A=>nx181);
   ix182 : aoi222 port map ( Y=>nx181, A0=>q_arr_9_5, A1=>nx523, B0=>
      q_arr_9_10, B1=>nx460, C0=>q_arr_9_8, C1=>nx479);
   ix89 : inv01 port map ( Y=>d_arr_1_6, A=>nx185);
   ix186 : aoi222 port map ( Y=>nx185, A0=>q_arr_9_6, A1=>nx523, B0=>
      q_arr_9_11, B1=>nx460, C0=>q_arr_9_9, C1=>nx479);
   ix101 : inv01 port map ( Y=>d_arr_1_7, A=>nx189);
   ix190 : aoi222 port map ( Y=>nx189, A0=>q_arr_9_7, A1=>nx523, B0=>
      q_arr_9_12, B1=>nx462, C0=>q_arr_9_10, C1=>nx481);
   ix113 : inv01 port map ( Y=>d_arr_1_8, A=>nx193);
   ix194 : aoi222 port map ( Y=>nx193, A0=>q_arr_9_8, A1=>nx523, B0=>
      q_arr_9_13, B1=>nx462, C0=>q_arr_9_11, C1=>nx481);
   ix125 : inv01 port map ( Y=>d_arr_1_9, A=>nx197);
   ix198 : aoi222 port map ( Y=>nx197, A0=>q_arr_9_9, A1=>nx523, B0=>
      q_arr_9_14, B1=>nx462, C0=>q_arr_9_12, C1=>nx481);
   ix137 : inv01 port map ( Y=>d_arr_1_10, A=>nx201);
   ix202 : aoi222 port map ( Y=>nx201, A0=>q_arr_9_10, A1=>nx523, B0=>
      q_arr_9_15, B1=>nx462, C0=>q_arr_9_13, C1=>nx481);
   ix149 : inv01 port map ( Y=>d_arr_1_11, A=>nx205);
   ix206 : aoi222 port map ( Y=>nx205, A0=>q_arr_9_11, A1=>nx523, B0=>
      q_arr_9_16, B1=>nx462, C0=>q_arr_9_14, C1=>nx481);
   ix161 : inv01 port map ( Y=>d_arr_1_12, A=>nx209);
   ix210 : aoi222 port map ( Y=>nx209, A0=>q_arr_9_12, A1=>nx525, B0=>
      q_arr_9_17, B1=>nx462, C0=>q_arr_9_15, C1=>nx481);
   ix173 : inv01 port map ( Y=>d_arr_1_13, A=>nx213);
   ix214 : aoi222 port map ( Y=>nx213, A0=>q_arr_9_13, A1=>nx525, B0=>
      q_arr_9_18, B1=>nx462, C0=>q_arr_9_16, C1=>nx481);
   ix185 : inv01 port map ( Y=>d_arr_1_14, A=>nx217);
   ix218 : aoi222 port map ( Y=>nx217, A0=>q_arr_9_14, A1=>nx525, B0=>
      q_arr_9_19, B1=>nx464, C0=>q_arr_9_17, C1=>nx483);
   ix197 : inv01 port map ( Y=>d_arr_1_15, A=>nx221);
   ix222 : aoi222 port map ( Y=>nx221, A0=>q_arr_9_15, A1=>nx525, B0=>
      q_arr_9_20, B1=>nx464, C0=>q_arr_9_18, C1=>nx483);
   ix209 : inv01 port map ( Y=>d_arr_1_16, A=>nx225);
   ix226 : aoi222 port map ( Y=>nx225, A0=>q_arr_9_16, A1=>nx525, B0=>
      q_arr_9_21, B1=>nx464, C0=>q_arr_9_19, C1=>nx483);
   ix221 : inv01 port map ( Y=>d_arr_1_17, A=>nx229);
   ix230 : aoi222 port map ( Y=>nx229, A0=>q_arr_9_17, A1=>nx525, B0=>
      q_arr_9_22, B1=>nx464, C0=>q_arr_9_20, C1=>nx483);
   ix233 : inv01 port map ( Y=>d_arr_1_18, A=>nx233);
   ix234 : aoi222 port map ( Y=>nx233, A0=>q_arr_9_18, A1=>nx525, B0=>
      q_arr_9_23, B1=>nx464, C0=>q_arr_9_21, C1=>nx483);
   ix245 : inv01 port map ( Y=>d_arr_1_19, A=>nx237);
   ix238 : aoi222 port map ( Y=>nx237, A0=>q_arr_9_19, A1=>nx527, B0=>nx555, 
      B1=>nx464, C0=>q_arr_9_22, C1=>nx483);
   ix257 : inv01 port map ( Y=>d_arr_1_20, A=>nx241);
   ix242 : aoi222 port map ( Y=>nx241, A0=>q_arr_9_20, A1=>nx527, B0=>
      q_arr_9_25, B1=>nx464, C0=>q_arr_9_23, C1=>nx483);
   ix269 : inv01 port map ( Y=>d_arr_1_21, A=>nx245);
   ix246 : aoi222 port map ( Y=>nx245, A0=>q_arr_9_21, A1=>nx527, B0=>
      q_arr_9_26, B1=>nx466, C0=>nx555, C1=>nx485);
   ix281 : inv01 port map ( Y=>d_arr_1_22, A=>nx249);
   ix250 : aoi222 port map ( Y=>nx249, A0=>q_arr_9_22, A1=>nx527, B0=>nx550, 
      B1=>nx466, C0=>q_arr_9_25, C1=>nx485);
   ix293 : inv01 port map ( Y=>d_arr_1_23, A=>nx253);
   ix254 : aoi222 port map ( Y=>nx253, A0=>q_arr_9_23, A1=>nx527, B0=>
      q_arr_9_28, B1=>nx466, C0=>q_arr_9_26, C1=>nx485);
   ix305 : inv01 port map ( Y=>d_arr_1_24, A=>nx257);
   ix258 : aoi222 port map ( Y=>nx257, A0=>nx555, A1=>nx527, B0=>q_arr_9_29, 
      B1=>nx466, C0=>nx550, C1=>nx485);
   ix317 : inv01 port map ( Y=>d_arr_1_25, A=>nx261);
   ix262 : aoi222 port map ( Y=>nx261, A0=>q_arr_9_25, A1=>nx527, B0=>
      q_arr_9_30, B1=>nx466, C0=>q_arr_9_28, C1=>nx485);
   ix329 : inv01 port map ( Y=>d_arr_1_26, A=>nx265);
   ix266 : aoi222 port map ( Y=>nx265, A0=>q_arr_9_26, A1=>nx529, B0=>
      q_arr_9_31, B1=>nx466, C0=>q_arr_9_29, C1=>nx485);
   ix337 : ao22 port map ( Y=>d_arr_1_27, A0=>nx553, A1=>nx529, B0=>
      q_arr_9_30, B1=>nx485);
   ix345 : ao22 port map ( Y=>d_arr_1_28, A0=>q_arr_9_28, A1=>nx529, B0=>
      q_arr_9_31, B1=>nx487);
   ix757 : nor02ii port map ( Y=>d_arr_1_29, A0=>nx540, A1=>q_arr_9_29);
   ix761 : nor02ii port map ( Y=>d_arr_1_30, A0=>nx540, A1=>q_arr_9_30);
   ix765 : nor02ii port map ( Y=>d_arr_1_31, A0=>nx540, A1=>q_arr_9_31);
   ix369 : nand02 port map ( Y=>d_arr_0_0, A0=>nx277, A1=>nx279);
   ix278 : aoi22 port map ( Y=>nx277, A0=>s2_5, A1=>nx466, B0=>q_arr_0_3, B1
      =>nx487);
   ix280 : aoi22 port map ( Y=>nx279, A0=>s2_0, A1=>nx499, B0=>q_arr_0_0, B1
      =>nx511);
   ix351 : nor02_2x port map ( Y=>nx350, A0=>filter_size, A1=>nx540);
   ix383 : nand02 port map ( Y=>d_arr_0_1, A0=>nx285, A1=>nx287);
   ix286 : aoi22 port map ( Y=>nx285, A0=>s2_6, A1=>nx469, B0=>q_arr_0_4, B1
      =>nx487);
   ix288 : aoi22 port map ( Y=>nx287, A0=>s2_1, A1=>nx499, B0=>q_arr_0_1, B1
      =>nx511);
   ix397 : nand02 port map ( Y=>d_arr_0_2, A0=>nx291, A1=>nx293);
   ix292 : aoi22 port map ( Y=>nx291, A0=>s2_7, A1=>nx469, B0=>q_arr_0_5, B1
      =>nx487);
   ix294 : aoi22 port map ( Y=>nx293, A0=>s2_2, A1=>nx499, B0=>q_arr_0_2, B1
      =>nx511);
   ix411 : nand02 port map ( Y=>d_arr_0_3, A0=>nx297, A1=>nx299);
   ix298 : aoi22 port map ( Y=>nx297, A0=>s2_8, A1=>nx469, B0=>q_arr_0_6, B1
      =>nx487);
   ix300 : aoi22 port map ( Y=>nx299, A0=>s2_3, A1=>nx499, B0=>q_arr_0_3, B1
      =>nx511);
   ix425 : nand02 port map ( Y=>d_arr_0_4, A0=>nx303, A1=>nx305);
   ix304 : aoi22 port map ( Y=>nx303, A0=>s2_9, A1=>nx469, B0=>q_arr_0_7, B1
      =>nx487);
   ix306 : aoi22 port map ( Y=>nx305, A0=>s2_4, A1=>nx499, B0=>q_arr_0_4, B1
      =>nx511);
   ix439 : nand02 port map ( Y=>d_arr_0_5, A0=>nx309, A1=>nx311);
   ix310 : aoi22 port map ( Y=>nx309, A0=>s2_10, A1=>nx469, B0=>q_arr_0_8, 
      B1=>nx487);
   ix312 : aoi22 port map ( Y=>nx311, A0=>s2_5, A1=>nx499, B0=>q_arr_0_5, B1
      =>nx511);
   ix453 : nand02 port map ( Y=>d_arr_0_6, A0=>nx315, A1=>nx317);
   ix316 : aoi22 port map ( Y=>nx315, A0=>s2_11, A1=>nx469, B0=>q_arr_0_9, 
      B1=>nx489);
   ix318 : aoi22 port map ( Y=>nx317, A0=>s2_6, A1=>nx499, B0=>q_arr_0_6, B1
      =>nx511);
   ix467 : nand02 port map ( Y=>d_arr_0_7, A0=>nx321, A1=>nx323);
   ix322 : aoi22 port map ( Y=>nx321, A0=>s2_12, A1=>nx469, B0=>q_arr_0_10, 
      B1=>nx489);
   ix324 : aoi22 port map ( Y=>nx323, A0=>s2_7, A1=>nx501, B0=>q_arr_0_7, B1
      =>nx513);
   ix481 : nand02 port map ( Y=>d_arr_0_8, A0=>nx327, A1=>nx329);
   ix328 : aoi22 port map ( Y=>nx327, A0=>s2_13, A1=>nx471, B0=>q_arr_0_11, 
      B1=>nx489);
   ix330 : aoi22 port map ( Y=>nx329, A0=>s2_8, A1=>nx501, B0=>q_arr_0_8, B1
      =>nx513);
   ix495 : nand02 port map ( Y=>d_arr_0_9, A0=>nx333, A1=>nx335);
   ix334 : aoi22 port map ( Y=>nx333, A0=>s2_14, A1=>nx471, B0=>q_arr_0_12, 
      B1=>nx489);
   ix336 : aoi22 port map ( Y=>nx335, A0=>s2_9, A1=>nx501, B0=>q_arr_0_9, B1
      =>nx513);
   ix509 : nand02 port map ( Y=>d_arr_0_10, A0=>nx339, A1=>nx341);
   ix340 : aoi22 port map ( Y=>nx339, A0=>s2_15, A1=>nx471, B0=>q_arr_0_13, 
      B1=>nx489);
   ix342 : aoi22 port map ( Y=>nx341, A0=>s2_10, A1=>nx501, B0=>q_arr_0_10, 
      B1=>nx513);
   ix523 : nand02 port map ( Y=>d_arr_0_11, A0=>nx345, A1=>nx347);
   ix346 : aoi22 port map ( Y=>nx345, A0=>s2_16, A1=>nx471, B0=>q_arr_0_14, 
      B1=>nx489);
   ix348 : aoi22 port map ( Y=>nx347, A0=>s2_11, A1=>nx501, B0=>q_arr_0_11, 
      B1=>nx513);
   ix537 : nand02 port map ( Y=>d_arr_0_12, A0=>nx351, A1=>nx353);
   ix352 : aoi22 port map ( Y=>nx351, A0=>s2_17, A1=>nx471, B0=>q_arr_0_15, 
      B1=>nx489);
   ix354 : aoi22 port map ( Y=>nx353, A0=>s2_12, A1=>nx501, B0=>q_arr_0_12, 
      B1=>nx513);
   ix551 : nand02 port map ( Y=>d_arr_0_13, A0=>nx357, A1=>nx359);
   ix358 : aoi22 port map ( Y=>nx357, A0=>s2_18, A1=>nx471, B0=>q_arr_0_16, 
      B1=>nx491);
   ix360 : aoi22 port map ( Y=>nx359, A0=>s2_13, A1=>nx501, B0=>q_arr_0_13, 
      B1=>nx513);
   ix565 : nand02 port map ( Y=>d_arr_0_14, A0=>nx363, A1=>nx365);
   ix364 : aoi22 port map ( Y=>nx363, A0=>s2_19, A1=>nx471, B0=>q_arr_0_17, 
      B1=>nx491);
   ix366 : aoi22 port map ( Y=>nx365, A0=>s2_14, A1=>nx503, B0=>q_arr_0_14, 
      B1=>nx515);
   ix579 : nand02 port map ( Y=>d_arr_0_15, A0=>nx369, A1=>nx371);
   ix370 : aoi22 port map ( Y=>nx369, A0=>s2_20, A1=>nx473, B0=>q_arr_0_18, 
      B1=>nx491);
   ix372 : aoi22 port map ( Y=>nx371, A0=>s2_15, A1=>nx503, B0=>q_arr_0_15, 
      B1=>nx515);
   ix593 : nand02 port map ( Y=>d_arr_0_16, A0=>nx375, A1=>nx377);
   ix376 : aoi22 port map ( Y=>nx375, A0=>s2_21, A1=>nx473, B0=>q_arr_0_19, 
      B1=>nx491);
   ix378 : aoi22 port map ( Y=>nx377, A0=>s2_16, A1=>nx503, B0=>q_arr_0_16, 
      B1=>nx515);
   ix607 : nand02 port map ( Y=>d_arr_0_17, A0=>nx381, A1=>nx383);
   ix382 : aoi22 port map ( Y=>nx381, A0=>s2_22, A1=>nx473, B0=>q_arr_0_20, 
      B1=>nx491);
   ix384 : aoi22 port map ( Y=>nx383, A0=>s2_17, A1=>nx503, B0=>q_arr_0_17, 
      B1=>nx515);
   ix621 : nand02 port map ( Y=>d_arr_0_18, A0=>nx387, A1=>nx389);
   ix388 : aoi22 port map ( Y=>nx387, A0=>s2_23, A1=>nx473, B0=>q_arr_0_21, 
      B1=>nx491);
   ix390 : aoi22 port map ( Y=>nx389, A0=>s2_18, A1=>nx503, B0=>q_arr_0_18, 
      B1=>nx515);
   ix635 : nand02 port map ( Y=>d_arr_0_19, A0=>nx393, A1=>nx395);
   ix394 : aoi22 port map ( Y=>nx393, A0=>s2_24, A1=>nx473, B0=>q_arr_0_22, 
      B1=>nx491);
   ix396 : aoi22 port map ( Y=>nx395, A0=>s2_19, A1=>nx503, B0=>q_arr_0_19, 
      B1=>nx515);
   ix649 : nand02 port map ( Y=>d_arr_0_20, A0=>nx399, A1=>nx401);
   ix400 : aoi22 port map ( Y=>nx399, A0=>s2_25, A1=>nx473, B0=>q_arr_0_23, 
      B1=>nx493);
   ix402 : aoi22 port map ( Y=>nx401, A0=>s2_20, A1=>nx503, B0=>q_arr_0_20, 
      B1=>nx515);
   ix663 : nand02 port map ( Y=>d_arr_0_21, A0=>nx405, A1=>nx407);
   ix406 : aoi22 port map ( Y=>nx405, A0=>s2_26, A1=>nx473, B0=>q_arr_0_24, 
      B1=>nx493);
   ix408 : aoi22 port map ( Y=>nx407, A0=>s2_21, A1=>nx505, B0=>q_arr_0_21, 
      B1=>nx517);
   ix677 : nand02 port map ( Y=>d_arr_0_22, A0=>nx411, A1=>nx413);
   ix412 : aoi22 port map ( Y=>nx411, A0=>s2_27, A1=>nx475, B0=>q_arr_0_25, 
      B1=>nx493);
   ix414 : aoi22 port map ( Y=>nx413, A0=>s2_22, A1=>nx505, B0=>q_arr_0_22, 
      B1=>nx517);
   ix691 : nand02 port map ( Y=>d_arr_0_23, A0=>nx417, A1=>nx419);
   ix418 : aoi22 port map ( Y=>nx417, A0=>s2_28, A1=>nx475, B0=>q_arr_0_26, 
      B1=>nx493);
   ix420 : aoi22 port map ( Y=>nx419, A0=>s2_23, A1=>nx505, B0=>q_arr_0_23, 
      B1=>nx517);
   ix705 : nand02 port map ( Y=>d_arr_0_24, A0=>nx423, A1=>nx425);
   ix424 : aoi22 port map ( Y=>nx423, A0=>s2_29, A1=>nx475, B0=>q_arr_0_27, 
      B1=>nx493);
   ix426 : aoi22 port map ( Y=>nx425, A0=>s2_24, A1=>nx505, B0=>q_arr_0_24, 
      B1=>nx517);
   ix719 : nand02 port map ( Y=>d_arr_0_25, A0=>nx429, A1=>nx431);
   ix430 : aoi22 port map ( Y=>nx429, A0=>s2_30, A1=>nx475, B0=>q_arr_0_28, 
      B1=>nx493);
   ix432 : aoi22 port map ( Y=>nx431, A0=>s2_25, A1=>nx505, B0=>q_arr_0_25, 
      B1=>nx517);
   ix733 : nand02 port map ( Y=>d_arr_0_26, A0=>nx435, A1=>nx437);
   ix436 : aoi22 port map ( Y=>nx435, A0=>s2_31, A1=>nx475, B0=>q_arr_0_29, 
      B1=>nx493);
   ix438 : aoi22 port map ( Y=>nx437, A0=>s2_26, A1=>nx505, B0=>q_arr_0_26, 
      B1=>nx517);
   ix743 : inv01 port map ( Y=>d_arr_0_27, A=>nx441);
   ix442 : aoi222 port map ( Y=>nx441, A0=>s2_27, A1=>nx505, B0=>q_arr_0_27, 
      B1=>nx517, C0=>q_arr_0_30, C1=>nx495);
   ix753 : inv01 port map ( Y=>d_arr_0_28, A=>nx445);
   ix446 : aoi222 port map ( Y=>nx445, A0=>s2_28, A1=>nx507, B0=>q_arr_0_28, 
      B1=>nx519, C0=>q_arr_0_31, C1=>nx495);
   ix771 : ao32 port map ( Y=>d_arr_0_29, A0=>q_arr_0_29, A1=>filter_size, 
      A2=>nx529, B0=>s2_29, B1=>nx507);
   ix777 : ao32 port map ( Y=>d_arr_0_30, A0=>q_arr_0_30, A1=>filter_size, 
      A2=>nx529, B0=>s2_30, B1=>nx507);
   ix783 : ao32 port map ( Y=>d_arr_0_31, A0=>q_arr_0_31, A1=>filter_size, 
      A2=>nx529, B0=>s2_31, B1=>nx507);
   ix457 : inv01 port map ( Y=>nx458, A=>nx6);
   ix459 : inv02 port map ( Y=>nx460, A=>nx531);
   ix461 : inv02 port map ( Y=>nx462, A=>nx531);
   ix463 : inv02 port map ( Y=>nx464, A=>nx531);
   ix465 : inv02 port map ( Y=>nx466, A=>nx531);
   ix468 : inv02 port map ( Y=>nx469, A=>nx531);
   ix470 : inv02 port map ( Y=>nx471, A=>nx458);
   ix472 : inv02 port map ( Y=>nx473, A=>nx458);
   ix474 : inv02 port map ( Y=>nx475, A=>nx458);
   ix476 : inv01 port map ( Y=>nx477, A=>nx10);
   ix478 : inv02 port map ( Y=>nx479, A=>nx533);
   ix480 : inv02 port map ( Y=>nx481, A=>nx533);
   ix482 : inv02 port map ( Y=>nx483, A=>nx533);
   ix484 : inv02 port map ( Y=>nx485, A=>nx533);
   ix486 : inv02 port map ( Y=>nx487, A=>nx533);
   ix488 : inv02 port map ( Y=>nx489, A=>nx477);
   ix490 : inv02 port map ( Y=>nx491, A=>nx477);
   ix492 : inv02 port map ( Y=>nx493, A=>nx477);
   ix494 : inv02 port map ( Y=>nx495, A=>nx477);
   ix496 : inv01 port map ( Y=>nx497, A=>nx350);
   ix498 : inv02 port map ( Y=>nx499, A=>nx497);
   ix500 : inv02 port map ( Y=>nx501, A=>nx497);
   ix502 : inv02 port map ( Y=>nx503, A=>nx497);
   ix504 : inv02 port map ( Y=>nx505, A=>nx497);
   ix506 : inv02 port map ( Y=>nx507, A=>nx497);
   ix510 : inv02 port map ( Y=>nx511, A=>nx509);
   ix512 : inv02 port map ( Y=>nx513, A=>nx509);
   ix514 : inv02 port map ( Y=>nx515, A=>nx509);
   ix516 : inv02 port map ( Y=>nx517, A=>nx509);
   ix518 : inv02 port map ( Y=>nx519, A=>nx509);
   ix520 : inv02 port map ( Y=>nx521, A=>operation);
   ix522 : inv02 port map ( Y=>nx523, A=>nx540);
   ix524 : inv02 port map ( Y=>nx525, A=>nx540);
   ix526 : inv02 port map ( Y=>nx527, A=>nx540);
   ix528 : inv02 port map ( Y=>nx529, A=>nx542);
   ix530 : inv01 port map ( Y=>nx531, A=>nx6);
   ix532 : inv01 port map ( Y=>nx533, A=>nx10);
   ix7 : nor02ii port map ( Y=>nx6, A0=>filter_size, A1=>nx542);
   ix11 : and02 port map ( Y=>nx10, A0=>filter_size, A1=>nx542);
   ix357 : nand02 port map ( Y=>nx509, A0=>filter_size, A1=>nx521);
   ix539 : inv02 port map ( Y=>nx540, A=>nx521);
   ix541 : inv02 port map ( Y=>nx542, A=>nx521);
   ix549 : buf02 port map ( Y=>nx550, A=>q_arr_9_27);
   ix552 : buf02 port map ( Y=>nx553, A=>q_arr_9_27);
   ix554 : buf02 port map ( Y=>nx555, A=>q_arr_9_24);
end Structural_unfold_3382_0 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity ReluLayer is
   port (
      d_arr_0_31 : OUT std_logic ;
      d_arr_0_30 : OUT std_logic ;
      d_arr_0_29 : OUT std_logic ;
      d_arr_0_28 : OUT std_logic ;
      d_arr_0_27 : OUT std_logic ;
      d_arr_0_26 : OUT std_logic ;
      d_arr_0_25 : OUT std_logic ;
      d_arr_0_24 : OUT std_logic ;
      d_arr_0_23 : OUT std_logic ;
      d_arr_0_22 : OUT std_logic ;
      d_arr_0_21 : OUT std_logic ;
      d_arr_0_20 : OUT std_logic ;
      d_arr_0_19 : OUT std_logic ;
      d_arr_0_18 : OUT std_logic ;
      d_arr_0_17 : OUT std_logic ;
      d_arr_0_16 : OUT std_logic ;
      d_arr_0_15 : OUT std_logic ;
      d_arr_0_14 : OUT std_logic ;
      d_arr_0_13 : OUT std_logic ;
      d_arr_0_12 : OUT std_logic ;
      d_arr_0_11 : OUT std_logic ;
      d_arr_0_10 : OUT std_logic ;
      d_arr_0_9 : OUT std_logic ;
      d_arr_0_8 : OUT std_logic ;
      d_arr_0_7 : OUT std_logic ;
      d_arr_0_6 : OUT std_logic ;
      d_arr_0_5 : OUT std_logic ;
      d_arr_0_4 : OUT std_logic ;
      d_arr_0_3 : OUT std_logic ;
      d_arr_0_2 : OUT std_logic ;
      d_arr_0_1 : OUT std_logic ;
      d_arr_0_0 : OUT std_logic ;
      d_arr_1_31 : OUT std_logic ;
      d_arr_1_30 : OUT std_logic ;
      d_arr_1_29 : OUT std_logic ;
      d_arr_1_28 : OUT std_logic ;
      d_arr_1_27 : OUT std_logic ;
      d_arr_1_26 : OUT std_logic ;
      d_arr_1_25 : OUT std_logic ;
      d_arr_1_24 : OUT std_logic ;
      d_arr_1_23 : OUT std_logic ;
      d_arr_1_22 : OUT std_logic ;
      d_arr_1_21 : OUT std_logic ;
      d_arr_1_20 : OUT std_logic ;
      d_arr_1_19 : OUT std_logic ;
      d_arr_1_18 : OUT std_logic ;
      d_arr_1_17 : OUT std_logic ;
      d_arr_1_16 : OUT std_logic ;
      d_arr_1_15 : OUT std_logic ;
      d_arr_1_14 : OUT std_logic ;
      d_arr_1_13 : OUT std_logic ;
      d_arr_1_12 : OUT std_logic ;
      d_arr_1_11 : OUT std_logic ;
      d_arr_1_10 : OUT std_logic ;
      d_arr_1_9 : OUT std_logic ;
      d_arr_1_8 : OUT std_logic ;
      d_arr_1_7 : OUT std_logic ;
      d_arr_1_6 : OUT std_logic ;
      d_arr_1_5 : OUT std_logic ;
      d_arr_1_4 : OUT std_logic ;
      d_arr_1_3 : OUT std_logic ;
      d_arr_1_2 : OUT std_logic ;
      d_arr_1_1 : OUT std_logic ;
      d_arr_1_0 : OUT std_logic ;
      d_arr_2_31 : OUT std_logic ;
      d_arr_2_30 : OUT std_logic ;
      d_arr_2_29 : OUT std_logic ;
      d_arr_2_28 : OUT std_logic ;
      d_arr_2_27 : OUT std_logic ;
      d_arr_2_26 : OUT std_logic ;
      d_arr_2_25 : OUT std_logic ;
      d_arr_2_24 : OUT std_logic ;
      d_arr_2_23 : OUT std_logic ;
      d_arr_2_22 : OUT std_logic ;
      d_arr_2_21 : OUT std_logic ;
      d_arr_2_20 : OUT std_logic ;
      d_arr_2_19 : OUT std_logic ;
      d_arr_2_18 : OUT std_logic ;
      d_arr_2_17 : OUT std_logic ;
      d_arr_2_16 : OUT std_logic ;
      d_arr_2_15 : OUT std_logic ;
      d_arr_2_14 : OUT std_logic ;
      d_arr_2_13 : OUT std_logic ;
      d_arr_2_12 : OUT std_logic ;
      d_arr_2_11 : OUT std_logic ;
      d_arr_2_10 : OUT std_logic ;
      d_arr_2_9 : OUT std_logic ;
      d_arr_2_8 : OUT std_logic ;
      d_arr_2_7 : OUT std_logic ;
      d_arr_2_6 : OUT std_logic ;
      d_arr_2_5 : OUT std_logic ;
      d_arr_2_4 : OUT std_logic ;
      d_arr_2_3 : OUT std_logic ;
      d_arr_2_2 : OUT std_logic ;
      d_arr_2_1 : OUT std_logic ;
      d_arr_2_0 : OUT std_logic ;
      d_arr_3_31 : OUT std_logic ;
      d_arr_3_30 : OUT std_logic ;
      d_arr_3_29 : OUT std_logic ;
      d_arr_3_28 : OUT std_logic ;
      d_arr_3_27 : OUT std_logic ;
      d_arr_3_26 : OUT std_logic ;
      d_arr_3_25 : OUT std_logic ;
      d_arr_3_24 : OUT std_logic ;
      d_arr_3_23 : OUT std_logic ;
      d_arr_3_22 : OUT std_logic ;
      d_arr_3_21 : OUT std_logic ;
      d_arr_3_20 : OUT std_logic ;
      d_arr_3_19 : OUT std_logic ;
      d_arr_3_18 : OUT std_logic ;
      d_arr_3_17 : OUT std_logic ;
      d_arr_3_16 : OUT std_logic ;
      d_arr_3_15 : OUT std_logic ;
      d_arr_3_14 : OUT std_logic ;
      d_arr_3_13 : OUT std_logic ;
      d_arr_3_12 : OUT std_logic ;
      d_arr_3_11 : OUT std_logic ;
      d_arr_3_10 : OUT std_logic ;
      d_arr_3_9 : OUT std_logic ;
      d_arr_3_8 : OUT std_logic ;
      d_arr_3_7 : OUT std_logic ;
      d_arr_3_6 : OUT std_logic ;
      d_arr_3_5 : OUT std_logic ;
      d_arr_3_4 : OUT std_logic ;
      d_arr_3_3 : OUT std_logic ;
      d_arr_3_2 : OUT std_logic ;
      d_arr_3_1 : OUT std_logic ;
      d_arr_3_0 : OUT std_logic ;
      d_arr_4_31 : OUT std_logic ;
      d_arr_4_30 : OUT std_logic ;
      d_arr_4_29 : OUT std_logic ;
      d_arr_4_28 : OUT std_logic ;
      d_arr_4_27 : OUT std_logic ;
      d_arr_4_26 : OUT std_logic ;
      d_arr_4_25 : OUT std_logic ;
      d_arr_4_24 : OUT std_logic ;
      d_arr_4_23 : OUT std_logic ;
      d_arr_4_22 : OUT std_logic ;
      d_arr_4_21 : OUT std_logic ;
      d_arr_4_20 : OUT std_logic ;
      d_arr_4_19 : OUT std_logic ;
      d_arr_4_18 : OUT std_logic ;
      d_arr_4_17 : OUT std_logic ;
      d_arr_4_16 : OUT std_logic ;
      d_arr_4_15 : OUT std_logic ;
      d_arr_4_14 : OUT std_logic ;
      d_arr_4_13 : OUT std_logic ;
      d_arr_4_12 : OUT std_logic ;
      d_arr_4_11 : OUT std_logic ;
      d_arr_4_10 : OUT std_logic ;
      d_arr_4_9 : OUT std_logic ;
      d_arr_4_8 : OUT std_logic ;
      d_arr_4_7 : OUT std_logic ;
      d_arr_4_6 : OUT std_logic ;
      d_arr_4_5 : OUT std_logic ;
      d_arr_4_4 : OUT std_logic ;
      d_arr_4_3 : OUT std_logic ;
      d_arr_4_2 : OUT std_logic ;
      d_arr_4_1 : OUT std_logic ;
      d_arr_4_0 : OUT std_logic ;
      d_arr_5_31 : OUT std_logic ;
      d_arr_5_30 : OUT std_logic ;
      d_arr_5_29 : OUT std_logic ;
      d_arr_5_28 : OUT std_logic ;
      d_arr_5_27 : OUT std_logic ;
      d_arr_5_26 : OUT std_logic ;
      d_arr_5_25 : OUT std_logic ;
      d_arr_5_24 : OUT std_logic ;
      d_arr_5_23 : OUT std_logic ;
      d_arr_5_22 : OUT std_logic ;
      d_arr_5_21 : OUT std_logic ;
      d_arr_5_20 : OUT std_logic ;
      d_arr_5_19 : OUT std_logic ;
      d_arr_5_18 : OUT std_logic ;
      d_arr_5_17 : OUT std_logic ;
      d_arr_5_16 : OUT std_logic ;
      d_arr_5_15 : OUT std_logic ;
      d_arr_5_14 : OUT std_logic ;
      d_arr_5_13 : OUT std_logic ;
      d_arr_5_12 : OUT std_logic ;
      d_arr_5_11 : OUT std_logic ;
      d_arr_5_10 : OUT std_logic ;
      d_arr_5_9 : OUT std_logic ;
      d_arr_5_8 : OUT std_logic ;
      d_arr_5_7 : OUT std_logic ;
      d_arr_5_6 : OUT std_logic ;
      d_arr_5_5 : OUT std_logic ;
      d_arr_5_4 : OUT std_logic ;
      d_arr_5_3 : OUT std_logic ;
      d_arr_5_2 : OUT std_logic ;
      d_arr_5_1 : OUT std_logic ;
      d_arr_5_0 : OUT std_logic ;
      d_arr_6_31 : OUT std_logic ;
      d_arr_6_30 : OUT std_logic ;
      d_arr_6_29 : OUT std_logic ;
      d_arr_6_28 : OUT std_logic ;
      d_arr_6_27 : OUT std_logic ;
      d_arr_6_26 : OUT std_logic ;
      d_arr_6_25 : OUT std_logic ;
      d_arr_6_24 : OUT std_logic ;
      d_arr_6_23 : OUT std_logic ;
      d_arr_6_22 : OUT std_logic ;
      d_arr_6_21 : OUT std_logic ;
      d_arr_6_20 : OUT std_logic ;
      d_arr_6_19 : OUT std_logic ;
      d_arr_6_18 : OUT std_logic ;
      d_arr_6_17 : OUT std_logic ;
      d_arr_6_16 : OUT std_logic ;
      d_arr_6_15 : OUT std_logic ;
      d_arr_6_14 : OUT std_logic ;
      d_arr_6_13 : OUT std_logic ;
      d_arr_6_12 : OUT std_logic ;
      d_arr_6_11 : OUT std_logic ;
      d_arr_6_10 : OUT std_logic ;
      d_arr_6_9 : OUT std_logic ;
      d_arr_6_8 : OUT std_logic ;
      d_arr_6_7 : OUT std_logic ;
      d_arr_6_6 : OUT std_logic ;
      d_arr_6_5 : OUT std_logic ;
      d_arr_6_4 : OUT std_logic ;
      d_arr_6_3 : OUT std_logic ;
      d_arr_6_2 : OUT std_logic ;
      d_arr_6_1 : OUT std_logic ;
      d_arr_6_0 : OUT std_logic ;
      d_arr_7_31 : OUT std_logic ;
      d_arr_7_30 : OUT std_logic ;
      d_arr_7_29 : OUT std_logic ;
      d_arr_7_28 : OUT std_logic ;
      d_arr_7_27 : OUT std_logic ;
      d_arr_7_26 : OUT std_logic ;
      d_arr_7_25 : OUT std_logic ;
      d_arr_7_24 : OUT std_logic ;
      d_arr_7_23 : OUT std_logic ;
      d_arr_7_22 : OUT std_logic ;
      d_arr_7_21 : OUT std_logic ;
      d_arr_7_20 : OUT std_logic ;
      d_arr_7_19 : OUT std_logic ;
      d_arr_7_18 : OUT std_logic ;
      d_arr_7_17 : OUT std_logic ;
      d_arr_7_16 : OUT std_logic ;
      d_arr_7_15 : OUT std_logic ;
      d_arr_7_14 : OUT std_logic ;
      d_arr_7_13 : OUT std_logic ;
      d_arr_7_12 : OUT std_logic ;
      d_arr_7_11 : OUT std_logic ;
      d_arr_7_10 : OUT std_logic ;
      d_arr_7_9 : OUT std_logic ;
      d_arr_7_8 : OUT std_logic ;
      d_arr_7_7 : OUT std_logic ;
      d_arr_7_6 : OUT std_logic ;
      d_arr_7_5 : OUT std_logic ;
      d_arr_7_4 : OUT std_logic ;
      d_arr_7_3 : OUT std_logic ;
      d_arr_7_2 : OUT std_logic ;
      d_arr_7_1 : OUT std_logic ;
      d_arr_7_0 : OUT std_logic ;
      d_arr_8_31 : OUT std_logic ;
      d_arr_8_30 : OUT std_logic ;
      d_arr_8_29 : OUT std_logic ;
      d_arr_8_28 : OUT std_logic ;
      d_arr_8_27 : OUT std_logic ;
      d_arr_8_26 : OUT std_logic ;
      d_arr_8_25 : OUT std_logic ;
      d_arr_8_24 : OUT std_logic ;
      d_arr_8_23 : OUT std_logic ;
      d_arr_8_22 : OUT std_logic ;
      d_arr_8_21 : OUT std_logic ;
      d_arr_8_20 : OUT std_logic ;
      d_arr_8_19 : OUT std_logic ;
      d_arr_8_18 : OUT std_logic ;
      d_arr_8_17 : OUT std_logic ;
      d_arr_8_16 : OUT std_logic ;
      d_arr_8_15 : OUT std_logic ;
      d_arr_8_14 : OUT std_logic ;
      d_arr_8_13 : OUT std_logic ;
      d_arr_8_12 : OUT std_logic ;
      d_arr_8_11 : OUT std_logic ;
      d_arr_8_10 : OUT std_logic ;
      d_arr_8_9 : OUT std_logic ;
      d_arr_8_8 : OUT std_logic ;
      d_arr_8_7 : OUT std_logic ;
      d_arr_8_6 : OUT std_logic ;
      d_arr_8_5 : OUT std_logic ;
      d_arr_8_4 : OUT std_logic ;
      d_arr_8_3 : OUT std_logic ;
      d_arr_8_2 : OUT std_logic ;
      d_arr_8_1 : OUT std_logic ;
      d_arr_8_0 : OUT std_logic ;
      d_arr_9_31 : OUT std_logic ;
      d_arr_9_30 : OUT std_logic ;
      d_arr_9_29 : OUT std_logic ;
      d_arr_9_28 : OUT std_logic ;
      d_arr_9_27 : OUT std_logic ;
      d_arr_9_26 : OUT std_logic ;
      d_arr_9_25 : OUT std_logic ;
      d_arr_9_24 : OUT std_logic ;
      d_arr_9_23 : OUT std_logic ;
      d_arr_9_22 : OUT std_logic ;
      d_arr_9_21 : OUT std_logic ;
      d_arr_9_20 : OUT std_logic ;
      d_arr_9_19 : OUT std_logic ;
      d_arr_9_18 : OUT std_logic ;
      d_arr_9_17 : OUT std_logic ;
      d_arr_9_16 : OUT std_logic ;
      d_arr_9_15 : OUT std_logic ;
      d_arr_9_14 : OUT std_logic ;
      d_arr_9_13 : OUT std_logic ;
      d_arr_9_12 : OUT std_logic ;
      d_arr_9_11 : OUT std_logic ;
      d_arr_9_10 : OUT std_logic ;
      d_arr_9_9 : OUT std_logic ;
      d_arr_9_8 : OUT std_logic ;
      d_arr_9_7 : OUT std_logic ;
      d_arr_9_6 : OUT std_logic ;
      d_arr_9_5 : OUT std_logic ;
      d_arr_9_4 : OUT std_logic ;
      d_arr_9_3 : OUT std_logic ;
      d_arr_9_2 : OUT std_logic ;
      d_arr_9_1 : OUT std_logic ;
      d_arr_9_0 : OUT std_logic ;
      d_arr_10_31 : OUT std_logic ;
      d_arr_10_30 : OUT std_logic ;
      d_arr_10_29 : OUT std_logic ;
      d_arr_10_28 : OUT std_logic ;
      d_arr_10_27 : OUT std_logic ;
      d_arr_10_26 : OUT std_logic ;
      d_arr_10_25 : OUT std_logic ;
      d_arr_10_24 : OUT std_logic ;
      d_arr_10_23 : OUT std_logic ;
      d_arr_10_22 : OUT std_logic ;
      d_arr_10_21 : OUT std_logic ;
      d_arr_10_20 : OUT std_logic ;
      d_arr_10_19 : OUT std_logic ;
      d_arr_10_18 : OUT std_logic ;
      d_arr_10_17 : OUT std_logic ;
      d_arr_10_16 : OUT std_logic ;
      d_arr_10_15 : OUT std_logic ;
      d_arr_10_14 : OUT std_logic ;
      d_arr_10_13 : OUT std_logic ;
      d_arr_10_12 : OUT std_logic ;
      d_arr_10_11 : OUT std_logic ;
      d_arr_10_10 : OUT std_logic ;
      d_arr_10_9 : OUT std_logic ;
      d_arr_10_8 : OUT std_logic ;
      d_arr_10_7 : OUT std_logic ;
      d_arr_10_6 : OUT std_logic ;
      d_arr_10_5 : OUT std_logic ;
      d_arr_10_4 : OUT std_logic ;
      d_arr_10_3 : OUT std_logic ;
      d_arr_10_2 : OUT std_logic ;
      d_arr_10_1 : OUT std_logic ;
      d_arr_10_0 : OUT std_logic ;
      d_arr_11_31 : OUT std_logic ;
      d_arr_11_30 : OUT std_logic ;
      d_arr_11_29 : OUT std_logic ;
      d_arr_11_28 : OUT std_logic ;
      d_arr_11_27 : OUT std_logic ;
      d_arr_11_26 : OUT std_logic ;
      d_arr_11_25 : OUT std_logic ;
      d_arr_11_24 : OUT std_logic ;
      d_arr_11_23 : OUT std_logic ;
      d_arr_11_22 : OUT std_logic ;
      d_arr_11_21 : OUT std_logic ;
      d_arr_11_20 : OUT std_logic ;
      d_arr_11_19 : OUT std_logic ;
      d_arr_11_18 : OUT std_logic ;
      d_arr_11_17 : OUT std_logic ;
      d_arr_11_16 : OUT std_logic ;
      d_arr_11_15 : OUT std_logic ;
      d_arr_11_14 : OUT std_logic ;
      d_arr_11_13 : OUT std_logic ;
      d_arr_11_12 : OUT std_logic ;
      d_arr_11_11 : OUT std_logic ;
      d_arr_11_10 : OUT std_logic ;
      d_arr_11_9 : OUT std_logic ;
      d_arr_11_8 : OUT std_logic ;
      d_arr_11_7 : OUT std_logic ;
      d_arr_11_6 : OUT std_logic ;
      d_arr_11_5 : OUT std_logic ;
      d_arr_11_4 : OUT std_logic ;
      d_arr_11_3 : OUT std_logic ;
      d_arr_11_2 : OUT std_logic ;
      d_arr_11_1 : OUT std_logic ;
      d_arr_11_0 : OUT std_logic ;
      d_arr_12_31 : OUT std_logic ;
      d_arr_12_30 : OUT std_logic ;
      d_arr_12_29 : OUT std_logic ;
      d_arr_12_28 : OUT std_logic ;
      d_arr_12_27 : OUT std_logic ;
      d_arr_12_26 : OUT std_logic ;
      d_arr_12_25 : OUT std_logic ;
      d_arr_12_24 : OUT std_logic ;
      d_arr_12_23 : OUT std_logic ;
      d_arr_12_22 : OUT std_logic ;
      d_arr_12_21 : OUT std_logic ;
      d_arr_12_20 : OUT std_logic ;
      d_arr_12_19 : OUT std_logic ;
      d_arr_12_18 : OUT std_logic ;
      d_arr_12_17 : OUT std_logic ;
      d_arr_12_16 : OUT std_logic ;
      d_arr_12_15 : OUT std_logic ;
      d_arr_12_14 : OUT std_logic ;
      d_arr_12_13 : OUT std_logic ;
      d_arr_12_12 : OUT std_logic ;
      d_arr_12_11 : OUT std_logic ;
      d_arr_12_10 : OUT std_logic ;
      d_arr_12_9 : OUT std_logic ;
      d_arr_12_8 : OUT std_logic ;
      d_arr_12_7 : OUT std_logic ;
      d_arr_12_6 : OUT std_logic ;
      d_arr_12_5 : OUT std_logic ;
      d_arr_12_4 : OUT std_logic ;
      d_arr_12_3 : OUT std_logic ;
      d_arr_12_2 : OUT std_logic ;
      d_arr_12_1 : OUT std_logic ;
      d_arr_12_0 : OUT std_logic ;
      d_arr_13_31 : OUT std_logic ;
      d_arr_13_30 : OUT std_logic ;
      d_arr_13_29 : OUT std_logic ;
      d_arr_13_28 : OUT std_logic ;
      d_arr_13_27 : OUT std_logic ;
      d_arr_13_26 : OUT std_logic ;
      d_arr_13_25 : OUT std_logic ;
      d_arr_13_24 : OUT std_logic ;
      d_arr_13_23 : OUT std_logic ;
      d_arr_13_22 : OUT std_logic ;
      d_arr_13_21 : OUT std_logic ;
      d_arr_13_20 : OUT std_logic ;
      d_arr_13_19 : OUT std_logic ;
      d_arr_13_18 : OUT std_logic ;
      d_arr_13_17 : OUT std_logic ;
      d_arr_13_16 : OUT std_logic ;
      d_arr_13_15 : OUT std_logic ;
      d_arr_13_14 : OUT std_logic ;
      d_arr_13_13 : OUT std_logic ;
      d_arr_13_12 : OUT std_logic ;
      d_arr_13_11 : OUT std_logic ;
      d_arr_13_10 : OUT std_logic ;
      d_arr_13_9 : OUT std_logic ;
      d_arr_13_8 : OUT std_logic ;
      d_arr_13_7 : OUT std_logic ;
      d_arr_13_6 : OUT std_logic ;
      d_arr_13_5 : OUT std_logic ;
      d_arr_13_4 : OUT std_logic ;
      d_arr_13_3 : OUT std_logic ;
      d_arr_13_2 : OUT std_logic ;
      d_arr_13_1 : OUT std_logic ;
      d_arr_13_0 : OUT std_logic ;
      d_arr_14_31 : OUT std_logic ;
      d_arr_14_30 : OUT std_logic ;
      d_arr_14_29 : OUT std_logic ;
      d_arr_14_28 : OUT std_logic ;
      d_arr_14_27 : OUT std_logic ;
      d_arr_14_26 : OUT std_logic ;
      d_arr_14_25 : OUT std_logic ;
      d_arr_14_24 : OUT std_logic ;
      d_arr_14_23 : OUT std_logic ;
      d_arr_14_22 : OUT std_logic ;
      d_arr_14_21 : OUT std_logic ;
      d_arr_14_20 : OUT std_logic ;
      d_arr_14_19 : OUT std_logic ;
      d_arr_14_18 : OUT std_logic ;
      d_arr_14_17 : OUT std_logic ;
      d_arr_14_16 : OUT std_logic ;
      d_arr_14_15 : OUT std_logic ;
      d_arr_14_14 : OUT std_logic ;
      d_arr_14_13 : OUT std_logic ;
      d_arr_14_12 : OUT std_logic ;
      d_arr_14_11 : OUT std_logic ;
      d_arr_14_10 : OUT std_logic ;
      d_arr_14_9 : OUT std_logic ;
      d_arr_14_8 : OUT std_logic ;
      d_arr_14_7 : OUT std_logic ;
      d_arr_14_6 : OUT std_logic ;
      d_arr_14_5 : OUT std_logic ;
      d_arr_14_4 : OUT std_logic ;
      d_arr_14_3 : OUT std_logic ;
      d_arr_14_2 : OUT std_logic ;
      d_arr_14_1 : OUT std_logic ;
      d_arr_14_0 : OUT std_logic ;
      d_arr_15_31 : OUT std_logic ;
      d_arr_15_30 : OUT std_logic ;
      d_arr_15_29 : OUT std_logic ;
      d_arr_15_28 : OUT std_logic ;
      d_arr_15_27 : OUT std_logic ;
      d_arr_15_26 : OUT std_logic ;
      d_arr_15_25 : OUT std_logic ;
      d_arr_15_24 : OUT std_logic ;
      d_arr_15_23 : OUT std_logic ;
      d_arr_15_22 : OUT std_logic ;
      d_arr_15_21 : OUT std_logic ;
      d_arr_15_20 : OUT std_logic ;
      d_arr_15_19 : OUT std_logic ;
      d_arr_15_18 : OUT std_logic ;
      d_arr_15_17 : OUT std_logic ;
      d_arr_15_16 : OUT std_logic ;
      d_arr_15_15 : OUT std_logic ;
      d_arr_15_14 : OUT std_logic ;
      d_arr_15_13 : OUT std_logic ;
      d_arr_15_12 : OUT std_logic ;
      d_arr_15_11 : OUT std_logic ;
      d_arr_15_10 : OUT std_logic ;
      d_arr_15_9 : OUT std_logic ;
      d_arr_15_8 : OUT std_logic ;
      d_arr_15_7 : OUT std_logic ;
      d_arr_15_6 : OUT std_logic ;
      d_arr_15_5 : OUT std_logic ;
      d_arr_15_4 : OUT std_logic ;
      d_arr_15_3 : OUT std_logic ;
      d_arr_15_2 : OUT std_logic ;
      d_arr_15_1 : OUT std_logic ;
      d_arr_15_0 : OUT std_logic ;
      d_arr_16_31 : OUT std_logic ;
      d_arr_16_30 : OUT std_logic ;
      d_arr_16_29 : OUT std_logic ;
      d_arr_16_28 : OUT std_logic ;
      d_arr_16_27 : OUT std_logic ;
      d_arr_16_26 : OUT std_logic ;
      d_arr_16_25 : OUT std_logic ;
      d_arr_16_24 : OUT std_logic ;
      d_arr_16_23 : OUT std_logic ;
      d_arr_16_22 : OUT std_logic ;
      d_arr_16_21 : OUT std_logic ;
      d_arr_16_20 : OUT std_logic ;
      d_arr_16_19 : OUT std_logic ;
      d_arr_16_18 : OUT std_logic ;
      d_arr_16_17 : OUT std_logic ;
      d_arr_16_16 : OUT std_logic ;
      d_arr_16_15 : OUT std_logic ;
      d_arr_16_14 : OUT std_logic ;
      d_arr_16_13 : OUT std_logic ;
      d_arr_16_12 : OUT std_logic ;
      d_arr_16_11 : OUT std_logic ;
      d_arr_16_10 : OUT std_logic ;
      d_arr_16_9 : OUT std_logic ;
      d_arr_16_8 : OUT std_logic ;
      d_arr_16_7 : OUT std_logic ;
      d_arr_16_6 : OUT std_logic ;
      d_arr_16_5 : OUT std_logic ;
      d_arr_16_4 : OUT std_logic ;
      d_arr_16_3 : OUT std_logic ;
      d_arr_16_2 : OUT std_logic ;
      d_arr_16_1 : OUT std_logic ;
      d_arr_16_0 : OUT std_logic ;
      d_arr_17_31 : OUT std_logic ;
      d_arr_17_30 : OUT std_logic ;
      d_arr_17_29 : OUT std_logic ;
      d_arr_17_28 : OUT std_logic ;
      d_arr_17_27 : OUT std_logic ;
      d_arr_17_26 : OUT std_logic ;
      d_arr_17_25 : OUT std_logic ;
      d_arr_17_24 : OUT std_logic ;
      d_arr_17_23 : OUT std_logic ;
      d_arr_17_22 : OUT std_logic ;
      d_arr_17_21 : OUT std_logic ;
      d_arr_17_20 : OUT std_logic ;
      d_arr_17_19 : OUT std_logic ;
      d_arr_17_18 : OUT std_logic ;
      d_arr_17_17 : OUT std_logic ;
      d_arr_17_16 : OUT std_logic ;
      d_arr_17_15 : OUT std_logic ;
      d_arr_17_14 : OUT std_logic ;
      d_arr_17_13 : OUT std_logic ;
      d_arr_17_12 : OUT std_logic ;
      d_arr_17_11 : OUT std_logic ;
      d_arr_17_10 : OUT std_logic ;
      d_arr_17_9 : OUT std_logic ;
      d_arr_17_8 : OUT std_logic ;
      d_arr_17_7 : OUT std_logic ;
      d_arr_17_6 : OUT std_logic ;
      d_arr_17_5 : OUT std_logic ;
      d_arr_17_4 : OUT std_logic ;
      d_arr_17_3 : OUT std_logic ;
      d_arr_17_2 : OUT std_logic ;
      d_arr_17_1 : OUT std_logic ;
      d_arr_17_0 : OUT std_logic ;
      d_arr_18_31 : OUT std_logic ;
      d_arr_18_30 : OUT std_logic ;
      d_arr_18_29 : OUT std_logic ;
      d_arr_18_28 : OUT std_logic ;
      d_arr_18_27 : OUT std_logic ;
      d_arr_18_26 : OUT std_logic ;
      d_arr_18_25 : OUT std_logic ;
      d_arr_18_24 : OUT std_logic ;
      d_arr_18_23 : OUT std_logic ;
      d_arr_18_22 : OUT std_logic ;
      d_arr_18_21 : OUT std_logic ;
      d_arr_18_20 : OUT std_logic ;
      d_arr_18_19 : OUT std_logic ;
      d_arr_18_18 : OUT std_logic ;
      d_arr_18_17 : OUT std_logic ;
      d_arr_18_16 : OUT std_logic ;
      d_arr_18_15 : OUT std_logic ;
      d_arr_18_14 : OUT std_logic ;
      d_arr_18_13 : OUT std_logic ;
      d_arr_18_12 : OUT std_logic ;
      d_arr_18_11 : OUT std_logic ;
      d_arr_18_10 : OUT std_logic ;
      d_arr_18_9 : OUT std_logic ;
      d_arr_18_8 : OUT std_logic ;
      d_arr_18_7 : OUT std_logic ;
      d_arr_18_6 : OUT std_logic ;
      d_arr_18_5 : OUT std_logic ;
      d_arr_18_4 : OUT std_logic ;
      d_arr_18_3 : OUT std_logic ;
      d_arr_18_2 : OUT std_logic ;
      d_arr_18_1 : OUT std_logic ;
      d_arr_18_0 : OUT std_logic ;
      d_arr_19_31 : OUT std_logic ;
      d_arr_19_30 : OUT std_logic ;
      d_arr_19_29 : OUT std_logic ;
      d_arr_19_28 : OUT std_logic ;
      d_arr_19_27 : OUT std_logic ;
      d_arr_19_26 : OUT std_logic ;
      d_arr_19_25 : OUT std_logic ;
      d_arr_19_24 : OUT std_logic ;
      d_arr_19_23 : OUT std_logic ;
      d_arr_19_22 : OUT std_logic ;
      d_arr_19_21 : OUT std_logic ;
      d_arr_19_20 : OUT std_logic ;
      d_arr_19_19 : OUT std_logic ;
      d_arr_19_18 : OUT std_logic ;
      d_arr_19_17 : OUT std_logic ;
      d_arr_19_16 : OUT std_logic ;
      d_arr_19_15 : OUT std_logic ;
      d_arr_19_14 : OUT std_logic ;
      d_arr_19_13 : OUT std_logic ;
      d_arr_19_12 : OUT std_logic ;
      d_arr_19_11 : OUT std_logic ;
      d_arr_19_10 : OUT std_logic ;
      d_arr_19_9 : OUT std_logic ;
      d_arr_19_8 : OUT std_logic ;
      d_arr_19_7 : OUT std_logic ;
      d_arr_19_6 : OUT std_logic ;
      d_arr_19_5 : OUT std_logic ;
      d_arr_19_4 : OUT std_logic ;
      d_arr_19_3 : OUT std_logic ;
      d_arr_19_2 : OUT std_logic ;
      d_arr_19_1 : OUT std_logic ;
      d_arr_19_0 : OUT std_logic ;
      d_arr_20_31 : OUT std_logic ;
      d_arr_20_30 : OUT std_logic ;
      d_arr_20_29 : OUT std_logic ;
      d_arr_20_28 : OUT std_logic ;
      d_arr_20_27 : OUT std_logic ;
      d_arr_20_26 : OUT std_logic ;
      d_arr_20_25 : OUT std_logic ;
      d_arr_20_24 : OUT std_logic ;
      d_arr_20_23 : OUT std_logic ;
      d_arr_20_22 : OUT std_logic ;
      d_arr_20_21 : OUT std_logic ;
      d_arr_20_20 : OUT std_logic ;
      d_arr_20_19 : OUT std_logic ;
      d_arr_20_18 : OUT std_logic ;
      d_arr_20_17 : OUT std_logic ;
      d_arr_20_16 : OUT std_logic ;
      d_arr_20_15 : OUT std_logic ;
      d_arr_20_14 : OUT std_logic ;
      d_arr_20_13 : OUT std_logic ;
      d_arr_20_12 : OUT std_logic ;
      d_arr_20_11 : OUT std_logic ;
      d_arr_20_10 : OUT std_logic ;
      d_arr_20_9 : OUT std_logic ;
      d_arr_20_8 : OUT std_logic ;
      d_arr_20_7 : OUT std_logic ;
      d_arr_20_6 : OUT std_logic ;
      d_arr_20_5 : OUT std_logic ;
      d_arr_20_4 : OUT std_logic ;
      d_arr_20_3 : OUT std_logic ;
      d_arr_20_2 : OUT std_logic ;
      d_arr_20_1 : OUT std_logic ;
      d_arr_20_0 : OUT std_logic ;
      d_arr_21_31 : OUT std_logic ;
      d_arr_21_30 : OUT std_logic ;
      d_arr_21_29 : OUT std_logic ;
      d_arr_21_28 : OUT std_logic ;
      d_arr_21_27 : OUT std_logic ;
      d_arr_21_26 : OUT std_logic ;
      d_arr_21_25 : OUT std_logic ;
      d_arr_21_24 : OUT std_logic ;
      d_arr_21_23 : OUT std_logic ;
      d_arr_21_22 : OUT std_logic ;
      d_arr_21_21 : OUT std_logic ;
      d_arr_21_20 : OUT std_logic ;
      d_arr_21_19 : OUT std_logic ;
      d_arr_21_18 : OUT std_logic ;
      d_arr_21_17 : OUT std_logic ;
      d_arr_21_16 : OUT std_logic ;
      d_arr_21_15 : OUT std_logic ;
      d_arr_21_14 : OUT std_logic ;
      d_arr_21_13 : OUT std_logic ;
      d_arr_21_12 : OUT std_logic ;
      d_arr_21_11 : OUT std_logic ;
      d_arr_21_10 : OUT std_logic ;
      d_arr_21_9 : OUT std_logic ;
      d_arr_21_8 : OUT std_logic ;
      d_arr_21_7 : OUT std_logic ;
      d_arr_21_6 : OUT std_logic ;
      d_arr_21_5 : OUT std_logic ;
      d_arr_21_4 : OUT std_logic ;
      d_arr_21_3 : OUT std_logic ;
      d_arr_21_2 : OUT std_logic ;
      d_arr_21_1 : OUT std_logic ;
      d_arr_21_0 : OUT std_logic ;
      d_arr_22_31 : OUT std_logic ;
      d_arr_22_30 : OUT std_logic ;
      d_arr_22_29 : OUT std_logic ;
      d_arr_22_28 : OUT std_logic ;
      d_arr_22_27 : OUT std_logic ;
      d_arr_22_26 : OUT std_logic ;
      d_arr_22_25 : OUT std_logic ;
      d_arr_22_24 : OUT std_logic ;
      d_arr_22_23 : OUT std_logic ;
      d_arr_22_22 : OUT std_logic ;
      d_arr_22_21 : OUT std_logic ;
      d_arr_22_20 : OUT std_logic ;
      d_arr_22_19 : OUT std_logic ;
      d_arr_22_18 : OUT std_logic ;
      d_arr_22_17 : OUT std_logic ;
      d_arr_22_16 : OUT std_logic ;
      d_arr_22_15 : OUT std_logic ;
      d_arr_22_14 : OUT std_logic ;
      d_arr_22_13 : OUT std_logic ;
      d_arr_22_12 : OUT std_logic ;
      d_arr_22_11 : OUT std_logic ;
      d_arr_22_10 : OUT std_logic ;
      d_arr_22_9 : OUT std_logic ;
      d_arr_22_8 : OUT std_logic ;
      d_arr_22_7 : OUT std_logic ;
      d_arr_22_6 : OUT std_logic ;
      d_arr_22_5 : OUT std_logic ;
      d_arr_22_4 : OUT std_logic ;
      d_arr_22_3 : OUT std_logic ;
      d_arr_22_2 : OUT std_logic ;
      d_arr_22_1 : OUT std_logic ;
      d_arr_22_0 : OUT std_logic ;
      d_arr_23_31 : OUT std_logic ;
      d_arr_23_30 : OUT std_logic ;
      d_arr_23_29 : OUT std_logic ;
      d_arr_23_28 : OUT std_logic ;
      d_arr_23_27 : OUT std_logic ;
      d_arr_23_26 : OUT std_logic ;
      d_arr_23_25 : OUT std_logic ;
      d_arr_23_24 : OUT std_logic ;
      d_arr_23_23 : OUT std_logic ;
      d_arr_23_22 : OUT std_logic ;
      d_arr_23_21 : OUT std_logic ;
      d_arr_23_20 : OUT std_logic ;
      d_arr_23_19 : OUT std_logic ;
      d_arr_23_18 : OUT std_logic ;
      d_arr_23_17 : OUT std_logic ;
      d_arr_23_16 : OUT std_logic ;
      d_arr_23_15 : OUT std_logic ;
      d_arr_23_14 : OUT std_logic ;
      d_arr_23_13 : OUT std_logic ;
      d_arr_23_12 : OUT std_logic ;
      d_arr_23_11 : OUT std_logic ;
      d_arr_23_10 : OUT std_logic ;
      d_arr_23_9 : OUT std_logic ;
      d_arr_23_8 : OUT std_logic ;
      d_arr_23_7 : OUT std_logic ;
      d_arr_23_6 : OUT std_logic ;
      d_arr_23_5 : OUT std_logic ;
      d_arr_23_4 : OUT std_logic ;
      d_arr_23_3 : OUT std_logic ;
      d_arr_23_2 : OUT std_logic ;
      d_arr_23_1 : OUT std_logic ;
      d_arr_23_0 : OUT std_logic ;
      d_arr_24_31 : OUT std_logic ;
      d_arr_24_30 : OUT std_logic ;
      d_arr_24_29 : OUT std_logic ;
      d_arr_24_28 : OUT std_logic ;
      d_arr_24_27 : OUT std_logic ;
      d_arr_24_26 : OUT std_logic ;
      d_arr_24_25 : OUT std_logic ;
      d_arr_24_24 : OUT std_logic ;
      d_arr_24_23 : OUT std_logic ;
      d_arr_24_22 : OUT std_logic ;
      d_arr_24_21 : OUT std_logic ;
      d_arr_24_20 : OUT std_logic ;
      d_arr_24_19 : OUT std_logic ;
      d_arr_24_18 : OUT std_logic ;
      d_arr_24_17 : OUT std_logic ;
      d_arr_24_16 : OUT std_logic ;
      d_arr_24_15 : OUT std_logic ;
      d_arr_24_14 : OUT std_logic ;
      d_arr_24_13 : OUT std_logic ;
      d_arr_24_12 : OUT std_logic ;
      d_arr_24_11 : OUT std_logic ;
      d_arr_24_10 : OUT std_logic ;
      d_arr_24_9 : OUT std_logic ;
      d_arr_24_8 : OUT std_logic ;
      d_arr_24_7 : OUT std_logic ;
      d_arr_24_6 : OUT std_logic ;
      d_arr_24_5 : OUT std_logic ;
      d_arr_24_4 : OUT std_logic ;
      d_arr_24_3 : OUT std_logic ;
      d_arr_24_2 : OUT std_logic ;
      d_arr_24_1 : OUT std_logic ;
      d_arr_24_0 : OUT std_logic ;
      q_arr_0_31 : IN std_logic ;
      q_arr_0_30 : IN std_logic ;
      q_arr_0_29 : IN std_logic ;
      q_arr_0_28 : IN std_logic ;
      q_arr_0_27 : IN std_logic ;
      q_arr_0_26 : IN std_logic ;
      q_arr_0_25 : IN std_logic ;
      q_arr_0_24 : IN std_logic ;
      q_arr_0_23 : IN std_logic ;
      q_arr_0_22 : IN std_logic ;
      q_arr_0_21 : IN std_logic ;
      q_arr_0_20 : IN std_logic ;
      q_arr_0_19 : IN std_logic ;
      q_arr_0_18 : IN std_logic ;
      q_arr_0_17 : IN std_logic ;
      q_arr_0_16 : IN std_logic ;
      q_arr_0_15 : IN std_logic ;
      q_arr_0_14 : IN std_logic ;
      q_arr_0_13 : IN std_logic ;
      q_arr_0_12 : IN std_logic ;
      q_arr_0_11 : IN std_logic ;
      q_arr_0_10 : IN std_logic ;
      q_arr_0_9 : IN std_logic ;
      q_arr_0_8 : IN std_logic ;
      q_arr_0_7 : IN std_logic ;
      q_arr_0_6 : IN std_logic ;
      q_arr_0_5 : IN std_logic ;
      q_arr_0_4 : IN std_logic ;
      q_arr_0_3 : IN std_logic ;
      q_arr_0_2 : IN std_logic ;
      q_arr_0_1 : IN std_logic ;
      q_arr_0_0 : IN std_logic ;
      q_arr_1_31 : IN std_logic ;
      q_arr_1_30 : IN std_logic ;
      q_arr_1_29 : IN std_logic ;
      q_arr_1_28 : IN std_logic ;
      q_arr_1_27 : IN std_logic ;
      q_arr_1_26 : IN std_logic ;
      q_arr_1_25 : IN std_logic ;
      q_arr_1_24 : IN std_logic ;
      q_arr_1_23 : IN std_logic ;
      q_arr_1_22 : IN std_logic ;
      q_arr_1_21 : IN std_logic ;
      q_arr_1_20 : IN std_logic ;
      q_arr_1_19 : IN std_logic ;
      q_arr_1_18 : IN std_logic ;
      q_arr_1_17 : IN std_logic ;
      q_arr_1_16 : IN std_logic ;
      q_arr_1_15 : IN std_logic ;
      q_arr_1_14 : IN std_logic ;
      q_arr_1_13 : IN std_logic ;
      q_arr_1_12 : IN std_logic ;
      q_arr_1_11 : IN std_logic ;
      q_arr_1_10 : IN std_logic ;
      q_arr_1_9 : IN std_logic ;
      q_arr_1_8 : IN std_logic ;
      q_arr_1_7 : IN std_logic ;
      q_arr_1_6 : IN std_logic ;
      q_arr_1_5 : IN std_logic ;
      q_arr_1_4 : IN std_logic ;
      q_arr_1_3 : IN std_logic ;
      q_arr_1_2 : IN std_logic ;
      q_arr_1_1 : IN std_logic ;
      q_arr_1_0 : IN std_logic ;
      q_arr_2_31 : IN std_logic ;
      q_arr_2_30 : IN std_logic ;
      q_arr_2_29 : IN std_logic ;
      q_arr_2_28 : IN std_logic ;
      q_arr_2_27 : IN std_logic ;
      q_arr_2_26 : IN std_logic ;
      q_arr_2_25 : IN std_logic ;
      q_arr_2_24 : IN std_logic ;
      q_arr_2_23 : IN std_logic ;
      q_arr_2_22 : IN std_logic ;
      q_arr_2_21 : IN std_logic ;
      q_arr_2_20 : IN std_logic ;
      q_arr_2_19 : IN std_logic ;
      q_arr_2_18 : IN std_logic ;
      q_arr_2_17 : IN std_logic ;
      q_arr_2_16 : IN std_logic ;
      q_arr_2_15 : IN std_logic ;
      q_arr_2_14 : IN std_logic ;
      q_arr_2_13 : IN std_logic ;
      q_arr_2_12 : IN std_logic ;
      q_arr_2_11 : IN std_logic ;
      q_arr_2_10 : IN std_logic ;
      q_arr_2_9 : IN std_logic ;
      q_arr_2_8 : IN std_logic ;
      q_arr_2_7 : IN std_logic ;
      q_arr_2_6 : IN std_logic ;
      q_arr_2_5 : IN std_logic ;
      q_arr_2_4 : IN std_logic ;
      q_arr_2_3 : IN std_logic ;
      q_arr_2_2 : IN std_logic ;
      q_arr_2_1 : IN std_logic ;
      q_arr_2_0 : IN std_logic ;
      q_arr_3_31 : IN std_logic ;
      q_arr_3_30 : IN std_logic ;
      q_arr_3_29 : IN std_logic ;
      q_arr_3_28 : IN std_logic ;
      q_arr_3_27 : IN std_logic ;
      q_arr_3_26 : IN std_logic ;
      q_arr_3_25 : IN std_logic ;
      q_arr_3_24 : IN std_logic ;
      q_arr_3_23 : IN std_logic ;
      q_arr_3_22 : IN std_logic ;
      q_arr_3_21 : IN std_logic ;
      q_arr_3_20 : IN std_logic ;
      q_arr_3_19 : IN std_logic ;
      q_arr_3_18 : IN std_logic ;
      q_arr_3_17 : IN std_logic ;
      q_arr_3_16 : IN std_logic ;
      q_arr_3_15 : IN std_logic ;
      q_arr_3_14 : IN std_logic ;
      q_arr_3_13 : IN std_logic ;
      q_arr_3_12 : IN std_logic ;
      q_arr_3_11 : IN std_logic ;
      q_arr_3_10 : IN std_logic ;
      q_arr_3_9 : IN std_logic ;
      q_arr_3_8 : IN std_logic ;
      q_arr_3_7 : IN std_logic ;
      q_arr_3_6 : IN std_logic ;
      q_arr_3_5 : IN std_logic ;
      q_arr_3_4 : IN std_logic ;
      q_arr_3_3 : IN std_logic ;
      q_arr_3_2 : IN std_logic ;
      q_arr_3_1 : IN std_logic ;
      q_arr_3_0 : IN std_logic ;
      q_arr_4_31 : IN std_logic ;
      q_arr_4_30 : IN std_logic ;
      q_arr_4_29 : IN std_logic ;
      q_arr_4_28 : IN std_logic ;
      q_arr_4_27 : IN std_logic ;
      q_arr_4_26 : IN std_logic ;
      q_arr_4_25 : IN std_logic ;
      q_arr_4_24 : IN std_logic ;
      q_arr_4_23 : IN std_logic ;
      q_arr_4_22 : IN std_logic ;
      q_arr_4_21 : IN std_logic ;
      q_arr_4_20 : IN std_logic ;
      q_arr_4_19 : IN std_logic ;
      q_arr_4_18 : IN std_logic ;
      q_arr_4_17 : IN std_logic ;
      q_arr_4_16 : IN std_logic ;
      q_arr_4_15 : IN std_logic ;
      q_arr_4_14 : IN std_logic ;
      q_arr_4_13 : IN std_logic ;
      q_arr_4_12 : IN std_logic ;
      q_arr_4_11 : IN std_logic ;
      q_arr_4_10 : IN std_logic ;
      q_arr_4_9 : IN std_logic ;
      q_arr_4_8 : IN std_logic ;
      q_arr_4_7 : IN std_logic ;
      q_arr_4_6 : IN std_logic ;
      q_arr_4_5 : IN std_logic ;
      q_arr_4_4 : IN std_logic ;
      q_arr_4_3 : IN std_logic ;
      q_arr_4_2 : IN std_logic ;
      q_arr_4_1 : IN std_logic ;
      q_arr_4_0 : IN std_logic ;
      q_arr_5_31 : IN std_logic ;
      q_arr_5_30 : IN std_logic ;
      q_arr_5_29 : IN std_logic ;
      q_arr_5_28 : IN std_logic ;
      q_arr_5_27 : IN std_logic ;
      q_arr_5_26 : IN std_logic ;
      q_arr_5_25 : IN std_logic ;
      q_arr_5_24 : IN std_logic ;
      q_arr_5_23 : IN std_logic ;
      q_arr_5_22 : IN std_logic ;
      q_arr_5_21 : IN std_logic ;
      q_arr_5_20 : IN std_logic ;
      q_arr_5_19 : IN std_logic ;
      q_arr_5_18 : IN std_logic ;
      q_arr_5_17 : IN std_logic ;
      q_arr_5_16 : IN std_logic ;
      q_arr_5_15 : IN std_logic ;
      q_arr_5_14 : IN std_logic ;
      q_arr_5_13 : IN std_logic ;
      q_arr_5_12 : IN std_logic ;
      q_arr_5_11 : IN std_logic ;
      q_arr_5_10 : IN std_logic ;
      q_arr_5_9 : IN std_logic ;
      q_arr_5_8 : IN std_logic ;
      q_arr_5_7 : IN std_logic ;
      q_arr_5_6 : IN std_logic ;
      q_arr_5_5 : IN std_logic ;
      q_arr_5_4 : IN std_logic ;
      q_arr_5_3 : IN std_logic ;
      q_arr_5_2 : IN std_logic ;
      q_arr_5_1 : IN std_logic ;
      q_arr_5_0 : IN std_logic ;
      q_arr_6_31 : IN std_logic ;
      q_arr_6_30 : IN std_logic ;
      q_arr_6_29 : IN std_logic ;
      q_arr_6_28 : IN std_logic ;
      q_arr_6_27 : IN std_logic ;
      q_arr_6_26 : IN std_logic ;
      q_arr_6_25 : IN std_logic ;
      q_arr_6_24 : IN std_logic ;
      q_arr_6_23 : IN std_logic ;
      q_arr_6_22 : IN std_logic ;
      q_arr_6_21 : IN std_logic ;
      q_arr_6_20 : IN std_logic ;
      q_arr_6_19 : IN std_logic ;
      q_arr_6_18 : IN std_logic ;
      q_arr_6_17 : IN std_logic ;
      q_arr_6_16 : IN std_logic ;
      q_arr_6_15 : IN std_logic ;
      q_arr_6_14 : IN std_logic ;
      q_arr_6_13 : IN std_logic ;
      q_arr_6_12 : IN std_logic ;
      q_arr_6_11 : IN std_logic ;
      q_arr_6_10 : IN std_logic ;
      q_arr_6_9 : IN std_logic ;
      q_arr_6_8 : IN std_logic ;
      q_arr_6_7 : IN std_logic ;
      q_arr_6_6 : IN std_logic ;
      q_arr_6_5 : IN std_logic ;
      q_arr_6_4 : IN std_logic ;
      q_arr_6_3 : IN std_logic ;
      q_arr_6_2 : IN std_logic ;
      q_arr_6_1 : IN std_logic ;
      q_arr_6_0 : IN std_logic ;
      q_arr_7_31 : IN std_logic ;
      q_arr_7_30 : IN std_logic ;
      q_arr_7_29 : IN std_logic ;
      q_arr_7_28 : IN std_logic ;
      q_arr_7_27 : IN std_logic ;
      q_arr_7_26 : IN std_logic ;
      q_arr_7_25 : IN std_logic ;
      q_arr_7_24 : IN std_logic ;
      q_arr_7_23 : IN std_logic ;
      q_arr_7_22 : IN std_logic ;
      q_arr_7_21 : IN std_logic ;
      q_arr_7_20 : IN std_logic ;
      q_arr_7_19 : IN std_logic ;
      q_arr_7_18 : IN std_logic ;
      q_arr_7_17 : IN std_logic ;
      q_arr_7_16 : IN std_logic ;
      q_arr_7_15 : IN std_logic ;
      q_arr_7_14 : IN std_logic ;
      q_arr_7_13 : IN std_logic ;
      q_arr_7_12 : IN std_logic ;
      q_arr_7_11 : IN std_logic ;
      q_arr_7_10 : IN std_logic ;
      q_arr_7_9 : IN std_logic ;
      q_arr_7_8 : IN std_logic ;
      q_arr_7_7 : IN std_logic ;
      q_arr_7_6 : IN std_logic ;
      q_arr_7_5 : IN std_logic ;
      q_arr_7_4 : IN std_logic ;
      q_arr_7_3 : IN std_logic ;
      q_arr_7_2 : IN std_logic ;
      q_arr_7_1 : IN std_logic ;
      q_arr_7_0 : IN std_logic ;
      q_arr_8_31 : IN std_logic ;
      q_arr_8_30 : IN std_logic ;
      q_arr_8_29 : IN std_logic ;
      q_arr_8_28 : IN std_logic ;
      q_arr_8_27 : IN std_logic ;
      q_arr_8_26 : IN std_logic ;
      q_arr_8_25 : IN std_logic ;
      q_arr_8_24 : IN std_logic ;
      q_arr_8_23 : IN std_logic ;
      q_arr_8_22 : IN std_logic ;
      q_arr_8_21 : IN std_logic ;
      q_arr_8_20 : IN std_logic ;
      q_arr_8_19 : IN std_logic ;
      q_arr_8_18 : IN std_logic ;
      q_arr_8_17 : IN std_logic ;
      q_arr_8_16 : IN std_logic ;
      q_arr_8_15 : IN std_logic ;
      q_arr_8_14 : IN std_logic ;
      q_arr_8_13 : IN std_logic ;
      q_arr_8_12 : IN std_logic ;
      q_arr_8_11 : IN std_logic ;
      q_arr_8_10 : IN std_logic ;
      q_arr_8_9 : IN std_logic ;
      q_arr_8_8 : IN std_logic ;
      q_arr_8_7 : IN std_logic ;
      q_arr_8_6 : IN std_logic ;
      q_arr_8_5 : IN std_logic ;
      q_arr_8_4 : IN std_logic ;
      q_arr_8_3 : IN std_logic ;
      q_arr_8_2 : IN std_logic ;
      q_arr_8_1 : IN std_logic ;
      q_arr_8_0 : IN std_logic ;
      q_arr_9_31 : IN std_logic ;
      q_arr_9_30 : IN std_logic ;
      q_arr_9_29 : IN std_logic ;
      q_arr_9_28 : IN std_logic ;
      q_arr_9_27 : IN std_logic ;
      q_arr_9_26 : IN std_logic ;
      q_arr_9_25 : IN std_logic ;
      q_arr_9_24 : IN std_logic ;
      q_arr_9_23 : IN std_logic ;
      q_arr_9_22 : IN std_logic ;
      q_arr_9_21 : IN std_logic ;
      q_arr_9_20 : IN std_logic ;
      q_arr_9_19 : IN std_logic ;
      q_arr_9_18 : IN std_logic ;
      q_arr_9_17 : IN std_logic ;
      q_arr_9_16 : IN std_logic ;
      q_arr_9_15 : IN std_logic ;
      q_arr_9_14 : IN std_logic ;
      q_arr_9_13 : IN std_logic ;
      q_arr_9_12 : IN std_logic ;
      q_arr_9_11 : IN std_logic ;
      q_arr_9_10 : IN std_logic ;
      q_arr_9_9 : IN std_logic ;
      q_arr_9_8 : IN std_logic ;
      q_arr_9_7 : IN std_logic ;
      q_arr_9_6 : IN std_logic ;
      q_arr_9_5 : IN std_logic ;
      q_arr_9_4 : IN std_logic ;
      q_arr_9_3 : IN std_logic ;
      q_arr_9_2 : IN std_logic ;
      q_arr_9_1 : IN std_logic ;
      q_arr_9_0 : IN std_logic ;
      q_arr_10_31 : IN std_logic ;
      q_arr_10_30 : IN std_logic ;
      q_arr_10_29 : IN std_logic ;
      q_arr_10_28 : IN std_logic ;
      q_arr_10_27 : IN std_logic ;
      q_arr_10_26 : IN std_logic ;
      q_arr_10_25 : IN std_logic ;
      q_arr_10_24 : IN std_logic ;
      q_arr_10_23 : IN std_logic ;
      q_arr_10_22 : IN std_logic ;
      q_arr_10_21 : IN std_logic ;
      q_arr_10_20 : IN std_logic ;
      q_arr_10_19 : IN std_logic ;
      q_arr_10_18 : IN std_logic ;
      q_arr_10_17 : IN std_logic ;
      q_arr_10_16 : IN std_logic ;
      q_arr_10_15 : IN std_logic ;
      q_arr_10_14 : IN std_logic ;
      q_arr_10_13 : IN std_logic ;
      q_arr_10_12 : IN std_logic ;
      q_arr_10_11 : IN std_logic ;
      q_arr_10_10 : IN std_logic ;
      q_arr_10_9 : IN std_logic ;
      q_arr_10_8 : IN std_logic ;
      q_arr_10_7 : IN std_logic ;
      q_arr_10_6 : IN std_logic ;
      q_arr_10_5 : IN std_logic ;
      q_arr_10_4 : IN std_logic ;
      q_arr_10_3 : IN std_logic ;
      q_arr_10_2 : IN std_logic ;
      q_arr_10_1 : IN std_logic ;
      q_arr_10_0 : IN std_logic ;
      q_arr_11_31 : IN std_logic ;
      q_arr_11_30 : IN std_logic ;
      q_arr_11_29 : IN std_logic ;
      q_arr_11_28 : IN std_logic ;
      q_arr_11_27 : IN std_logic ;
      q_arr_11_26 : IN std_logic ;
      q_arr_11_25 : IN std_logic ;
      q_arr_11_24 : IN std_logic ;
      q_arr_11_23 : IN std_logic ;
      q_arr_11_22 : IN std_logic ;
      q_arr_11_21 : IN std_logic ;
      q_arr_11_20 : IN std_logic ;
      q_arr_11_19 : IN std_logic ;
      q_arr_11_18 : IN std_logic ;
      q_arr_11_17 : IN std_logic ;
      q_arr_11_16 : IN std_logic ;
      q_arr_11_15 : IN std_logic ;
      q_arr_11_14 : IN std_logic ;
      q_arr_11_13 : IN std_logic ;
      q_arr_11_12 : IN std_logic ;
      q_arr_11_11 : IN std_logic ;
      q_arr_11_10 : IN std_logic ;
      q_arr_11_9 : IN std_logic ;
      q_arr_11_8 : IN std_logic ;
      q_arr_11_7 : IN std_logic ;
      q_arr_11_6 : IN std_logic ;
      q_arr_11_5 : IN std_logic ;
      q_arr_11_4 : IN std_logic ;
      q_arr_11_3 : IN std_logic ;
      q_arr_11_2 : IN std_logic ;
      q_arr_11_1 : IN std_logic ;
      q_arr_11_0 : IN std_logic ;
      q_arr_12_31 : IN std_logic ;
      q_arr_12_30 : IN std_logic ;
      q_arr_12_29 : IN std_logic ;
      q_arr_12_28 : IN std_logic ;
      q_arr_12_27 : IN std_logic ;
      q_arr_12_26 : IN std_logic ;
      q_arr_12_25 : IN std_logic ;
      q_arr_12_24 : IN std_logic ;
      q_arr_12_23 : IN std_logic ;
      q_arr_12_22 : IN std_logic ;
      q_arr_12_21 : IN std_logic ;
      q_arr_12_20 : IN std_logic ;
      q_arr_12_19 : IN std_logic ;
      q_arr_12_18 : IN std_logic ;
      q_arr_12_17 : IN std_logic ;
      q_arr_12_16 : IN std_logic ;
      q_arr_12_15 : IN std_logic ;
      q_arr_12_14 : IN std_logic ;
      q_arr_12_13 : IN std_logic ;
      q_arr_12_12 : IN std_logic ;
      q_arr_12_11 : IN std_logic ;
      q_arr_12_10 : IN std_logic ;
      q_arr_12_9 : IN std_logic ;
      q_arr_12_8 : IN std_logic ;
      q_arr_12_7 : IN std_logic ;
      q_arr_12_6 : IN std_logic ;
      q_arr_12_5 : IN std_logic ;
      q_arr_12_4 : IN std_logic ;
      q_arr_12_3 : IN std_logic ;
      q_arr_12_2 : IN std_logic ;
      q_arr_12_1 : IN std_logic ;
      q_arr_12_0 : IN std_logic ;
      q_arr_13_31 : IN std_logic ;
      q_arr_13_30 : IN std_logic ;
      q_arr_13_29 : IN std_logic ;
      q_arr_13_28 : IN std_logic ;
      q_arr_13_27 : IN std_logic ;
      q_arr_13_26 : IN std_logic ;
      q_arr_13_25 : IN std_logic ;
      q_arr_13_24 : IN std_logic ;
      q_arr_13_23 : IN std_logic ;
      q_arr_13_22 : IN std_logic ;
      q_arr_13_21 : IN std_logic ;
      q_arr_13_20 : IN std_logic ;
      q_arr_13_19 : IN std_logic ;
      q_arr_13_18 : IN std_logic ;
      q_arr_13_17 : IN std_logic ;
      q_arr_13_16 : IN std_logic ;
      q_arr_13_15 : IN std_logic ;
      q_arr_13_14 : IN std_logic ;
      q_arr_13_13 : IN std_logic ;
      q_arr_13_12 : IN std_logic ;
      q_arr_13_11 : IN std_logic ;
      q_arr_13_10 : IN std_logic ;
      q_arr_13_9 : IN std_logic ;
      q_arr_13_8 : IN std_logic ;
      q_arr_13_7 : IN std_logic ;
      q_arr_13_6 : IN std_logic ;
      q_arr_13_5 : IN std_logic ;
      q_arr_13_4 : IN std_logic ;
      q_arr_13_3 : IN std_logic ;
      q_arr_13_2 : IN std_logic ;
      q_arr_13_1 : IN std_logic ;
      q_arr_13_0 : IN std_logic ;
      q_arr_14_31 : IN std_logic ;
      q_arr_14_30 : IN std_logic ;
      q_arr_14_29 : IN std_logic ;
      q_arr_14_28 : IN std_logic ;
      q_arr_14_27 : IN std_logic ;
      q_arr_14_26 : IN std_logic ;
      q_arr_14_25 : IN std_logic ;
      q_arr_14_24 : IN std_logic ;
      q_arr_14_23 : IN std_logic ;
      q_arr_14_22 : IN std_logic ;
      q_arr_14_21 : IN std_logic ;
      q_arr_14_20 : IN std_logic ;
      q_arr_14_19 : IN std_logic ;
      q_arr_14_18 : IN std_logic ;
      q_arr_14_17 : IN std_logic ;
      q_arr_14_16 : IN std_logic ;
      q_arr_14_15 : IN std_logic ;
      q_arr_14_14 : IN std_logic ;
      q_arr_14_13 : IN std_logic ;
      q_arr_14_12 : IN std_logic ;
      q_arr_14_11 : IN std_logic ;
      q_arr_14_10 : IN std_logic ;
      q_arr_14_9 : IN std_logic ;
      q_arr_14_8 : IN std_logic ;
      q_arr_14_7 : IN std_logic ;
      q_arr_14_6 : IN std_logic ;
      q_arr_14_5 : IN std_logic ;
      q_arr_14_4 : IN std_logic ;
      q_arr_14_3 : IN std_logic ;
      q_arr_14_2 : IN std_logic ;
      q_arr_14_1 : IN std_logic ;
      q_arr_14_0 : IN std_logic ;
      q_arr_15_31 : IN std_logic ;
      q_arr_15_30 : IN std_logic ;
      q_arr_15_29 : IN std_logic ;
      q_arr_15_28 : IN std_logic ;
      q_arr_15_27 : IN std_logic ;
      q_arr_15_26 : IN std_logic ;
      q_arr_15_25 : IN std_logic ;
      q_arr_15_24 : IN std_logic ;
      q_arr_15_23 : IN std_logic ;
      q_arr_15_22 : IN std_logic ;
      q_arr_15_21 : IN std_logic ;
      q_arr_15_20 : IN std_logic ;
      q_arr_15_19 : IN std_logic ;
      q_arr_15_18 : IN std_logic ;
      q_arr_15_17 : IN std_logic ;
      q_arr_15_16 : IN std_logic ;
      q_arr_15_15 : IN std_logic ;
      q_arr_15_14 : IN std_logic ;
      q_arr_15_13 : IN std_logic ;
      q_arr_15_12 : IN std_logic ;
      q_arr_15_11 : IN std_logic ;
      q_arr_15_10 : IN std_logic ;
      q_arr_15_9 : IN std_logic ;
      q_arr_15_8 : IN std_logic ;
      q_arr_15_7 : IN std_logic ;
      q_arr_15_6 : IN std_logic ;
      q_arr_15_5 : IN std_logic ;
      q_arr_15_4 : IN std_logic ;
      q_arr_15_3 : IN std_logic ;
      q_arr_15_2 : IN std_logic ;
      q_arr_15_1 : IN std_logic ;
      q_arr_15_0 : IN std_logic ;
      q_arr_16_31 : IN std_logic ;
      q_arr_16_30 : IN std_logic ;
      q_arr_16_29 : IN std_logic ;
      q_arr_16_28 : IN std_logic ;
      q_arr_16_27 : IN std_logic ;
      q_arr_16_26 : IN std_logic ;
      q_arr_16_25 : IN std_logic ;
      q_arr_16_24 : IN std_logic ;
      q_arr_16_23 : IN std_logic ;
      q_arr_16_22 : IN std_logic ;
      q_arr_16_21 : IN std_logic ;
      q_arr_16_20 : IN std_logic ;
      q_arr_16_19 : IN std_logic ;
      q_arr_16_18 : IN std_logic ;
      q_arr_16_17 : IN std_logic ;
      q_arr_16_16 : IN std_logic ;
      q_arr_16_15 : IN std_logic ;
      q_arr_16_14 : IN std_logic ;
      q_arr_16_13 : IN std_logic ;
      q_arr_16_12 : IN std_logic ;
      q_arr_16_11 : IN std_logic ;
      q_arr_16_10 : IN std_logic ;
      q_arr_16_9 : IN std_logic ;
      q_arr_16_8 : IN std_logic ;
      q_arr_16_7 : IN std_logic ;
      q_arr_16_6 : IN std_logic ;
      q_arr_16_5 : IN std_logic ;
      q_arr_16_4 : IN std_logic ;
      q_arr_16_3 : IN std_logic ;
      q_arr_16_2 : IN std_logic ;
      q_arr_16_1 : IN std_logic ;
      q_arr_16_0 : IN std_logic ;
      q_arr_17_31 : IN std_logic ;
      q_arr_17_30 : IN std_logic ;
      q_arr_17_29 : IN std_logic ;
      q_arr_17_28 : IN std_logic ;
      q_arr_17_27 : IN std_logic ;
      q_arr_17_26 : IN std_logic ;
      q_arr_17_25 : IN std_logic ;
      q_arr_17_24 : IN std_logic ;
      q_arr_17_23 : IN std_logic ;
      q_arr_17_22 : IN std_logic ;
      q_arr_17_21 : IN std_logic ;
      q_arr_17_20 : IN std_logic ;
      q_arr_17_19 : IN std_logic ;
      q_arr_17_18 : IN std_logic ;
      q_arr_17_17 : IN std_logic ;
      q_arr_17_16 : IN std_logic ;
      q_arr_17_15 : IN std_logic ;
      q_arr_17_14 : IN std_logic ;
      q_arr_17_13 : IN std_logic ;
      q_arr_17_12 : IN std_logic ;
      q_arr_17_11 : IN std_logic ;
      q_arr_17_10 : IN std_logic ;
      q_arr_17_9 : IN std_logic ;
      q_arr_17_8 : IN std_logic ;
      q_arr_17_7 : IN std_logic ;
      q_arr_17_6 : IN std_logic ;
      q_arr_17_5 : IN std_logic ;
      q_arr_17_4 : IN std_logic ;
      q_arr_17_3 : IN std_logic ;
      q_arr_17_2 : IN std_logic ;
      q_arr_17_1 : IN std_logic ;
      q_arr_17_0 : IN std_logic ;
      q_arr_18_31 : IN std_logic ;
      q_arr_18_30 : IN std_logic ;
      q_arr_18_29 : IN std_logic ;
      q_arr_18_28 : IN std_logic ;
      q_arr_18_27 : IN std_logic ;
      q_arr_18_26 : IN std_logic ;
      q_arr_18_25 : IN std_logic ;
      q_arr_18_24 : IN std_logic ;
      q_arr_18_23 : IN std_logic ;
      q_arr_18_22 : IN std_logic ;
      q_arr_18_21 : IN std_logic ;
      q_arr_18_20 : IN std_logic ;
      q_arr_18_19 : IN std_logic ;
      q_arr_18_18 : IN std_logic ;
      q_arr_18_17 : IN std_logic ;
      q_arr_18_16 : IN std_logic ;
      q_arr_18_15 : IN std_logic ;
      q_arr_18_14 : IN std_logic ;
      q_arr_18_13 : IN std_logic ;
      q_arr_18_12 : IN std_logic ;
      q_arr_18_11 : IN std_logic ;
      q_arr_18_10 : IN std_logic ;
      q_arr_18_9 : IN std_logic ;
      q_arr_18_8 : IN std_logic ;
      q_arr_18_7 : IN std_logic ;
      q_arr_18_6 : IN std_logic ;
      q_arr_18_5 : IN std_logic ;
      q_arr_18_4 : IN std_logic ;
      q_arr_18_3 : IN std_logic ;
      q_arr_18_2 : IN std_logic ;
      q_arr_18_1 : IN std_logic ;
      q_arr_18_0 : IN std_logic ;
      q_arr_19_31 : IN std_logic ;
      q_arr_19_30 : IN std_logic ;
      q_arr_19_29 : IN std_logic ;
      q_arr_19_28 : IN std_logic ;
      q_arr_19_27 : IN std_logic ;
      q_arr_19_26 : IN std_logic ;
      q_arr_19_25 : IN std_logic ;
      q_arr_19_24 : IN std_logic ;
      q_arr_19_23 : IN std_logic ;
      q_arr_19_22 : IN std_logic ;
      q_arr_19_21 : IN std_logic ;
      q_arr_19_20 : IN std_logic ;
      q_arr_19_19 : IN std_logic ;
      q_arr_19_18 : IN std_logic ;
      q_arr_19_17 : IN std_logic ;
      q_arr_19_16 : IN std_logic ;
      q_arr_19_15 : IN std_logic ;
      q_arr_19_14 : IN std_logic ;
      q_arr_19_13 : IN std_logic ;
      q_arr_19_12 : IN std_logic ;
      q_arr_19_11 : IN std_logic ;
      q_arr_19_10 : IN std_logic ;
      q_arr_19_9 : IN std_logic ;
      q_arr_19_8 : IN std_logic ;
      q_arr_19_7 : IN std_logic ;
      q_arr_19_6 : IN std_logic ;
      q_arr_19_5 : IN std_logic ;
      q_arr_19_4 : IN std_logic ;
      q_arr_19_3 : IN std_logic ;
      q_arr_19_2 : IN std_logic ;
      q_arr_19_1 : IN std_logic ;
      q_arr_19_0 : IN std_logic ;
      q_arr_20_31 : IN std_logic ;
      q_arr_20_30 : IN std_logic ;
      q_arr_20_29 : IN std_logic ;
      q_arr_20_28 : IN std_logic ;
      q_arr_20_27 : IN std_logic ;
      q_arr_20_26 : IN std_logic ;
      q_arr_20_25 : IN std_logic ;
      q_arr_20_24 : IN std_logic ;
      q_arr_20_23 : IN std_logic ;
      q_arr_20_22 : IN std_logic ;
      q_arr_20_21 : IN std_logic ;
      q_arr_20_20 : IN std_logic ;
      q_arr_20_19 : IN std_logic ;
      q_arr_20_18 : IN std_logic ;
      q_arr_20_17 : IN std_logic ;
      q_arr_20_16 : IN std_logic ;
      q_arr_20_15 : IN std_logic ;
      q_arr_20_14 : IN std_logic ;
      q_arr_20_13 : IN std_logic ;
      q_arr_20_12 : IN std_logic ;
      q_arr_20_11 : IN std_logic ;
      q_arr_20_10 : IN std_logic ;
      q_arr_20_9 : IN std_logic ;
      q_arr_20_8 : IN std_logic ;
      q_arr_20_7 : IN std_logic ;
      q_arr_20_6 : IN std_logic ;
      q_arr_20_5 : IN std_logic ;
      q_arr_20_4 : IN std_logic ;
      q_arr_20_3 : IN std_logic ;
      q_arr_20_2 : IN std_logic ;
      q_arr_20_1 : IN std_logic ;
      q_arr_20_0 : IN std_logic ;
      q_arr_21_31 : IN std_logic ;
      q_arr_21_30 : IN std_logic ;
      q_arr_21_29 : IN std_logic ;
      q_arr_21_28 : IN std_logic ;
      q_arr_21_27 : IN std_logic ;
      q_arr_21_26 : IN std_logic ;
      q_arr_21_25 : IN std_logic ;
      q_arr_21_24 : IN std_logic ;
      q_arr_21_23 : IN std_logic ;
      q_arr_21_22 : IN std_logic ;
      q_arr_21_21 : IN std_logic ;
      q_arr_21_20 : IN std_logic ;
      q_arr_21_19 : IN std_logic ;
      q_arr_21_18 : IN std_logic ;
      q_arr_21_17 : IN std_logic ;
      q_arr_21_16 : IN std_logic ;
      q_arr_21_15 : IN std_logic ;
      q_arr_21_14 : IN std_logic ;
      q_arr_21_13 : IN std_logic ;
      q_arr_21_12 : IN std_logic ;
      q_arr_21_11 : IN std_logic ;
      q_arr_21_10 : IN std_logic ;
      q_arr_21_9 : IN std_logic ;
      q_arr_21_8 : IN std_logic ;
      q_arr_21_7 : IN std_logic ;
      q_arr_21_6 : IN std_logic ;
      q_arr_21_5 : IN std_logic ;
      q_arr_21_4 : IN std_logic ;
      q_arr_21_3 : IN std_logic ;
      q_arr_21_2 : IN std_logic ;
      q_arr_21_1 : IN std_logic ;
      q_arr_21_0 : IN std_logic ;
      q_arr_22_31 : IN std_logic ;
      q_arr_22_30 : IN std_logic ;
      q_arr_22_29 : IN std_logic ;
      q_arr_22_28 : IN std_logic ;
      q_arr_22_27 : IN std_logic ;
      q_arr_22_26 : IN std_logic ;
      q_arr_22_25 : IN std_logic ;
      q_arr_22_24 : IN std_logic ;
      q_arr_22_23 : IN std_logic ;
      q_arr_22_22 : IN std_logic ;
      q_arr_22_21 : IN std_logic ;
      q_arr_22_20 : IN std_logic ;
      q_arr_22_19 : IN std_logic ;
      q_arr_22_18 : IN std_logic ;
      q_arr_22_17 : IN std_logic ;
      q_arr_22_16 : IN std_logic ;
      q_arr_22_15 : IN std_logic ;
      q_arr_22_14 : IN std_logic ;
      q_arr_22_13 : IN std_logic ;
      q_arr_22_12 : IN std_logic ;
      q_arr_22_11 : IN std_logic ;
      q_arr_22_10 : IN std_logic ;
      q_arr_22_9 : IN std_logic ;
      q_arr_22_8 : IN std_logic ;
      q_arr_22_7 : IN std_logic ;
      q_arr_22_6 : IN std_logic ;
      q_arr_22_5 : IN std_logic ;
      q_arr_22_4 : IN std_logic ;
      q_arr_22_3 : IN std_logic ;
      q_arr_22_2 : IN std_logic ;
      q_arr_22_1 : IN std_logic ;
      q_arr_22_0 : IN std_logic ;
      q_arr_23_31 : IN std_logic ;
      q_arr_23_30 : IN std_logic ;
      q_arr_23_29 : IN std_logic ;
      q_arr_23_28 : IN std_logic ;
      q_arr_23_27 : IN std_logic ;
      q_arr_23_26 : IN std_logic ;
      q_arr_23_25 : IN std_logic ;
      q_arr_23_24 : IN std_logic ;
      q_arr_23_23 : IN std_logic ;
      q_arr_23_22 : IN std_logic ;
      q_arr_23_21 : IN std_logic ;
      q_arr_23_20 : IN std_logic ;
      q_arr_23_19 : IN std_logic ;
      q_arr_23_18 : IN std_logic ;
      q_arr_23_17 : IN std_logic ;
      q_arr_23_16 : IN std_logic ;
      q_arr_23_15 : IN std_logic ;
      q_arr_23_14 : IN std_logic ;
      q_arr_23_13 : IN std_logic ;
      q_arr_23_12 : IN std_logic ;
      q_arr_23_11 : IN std_logic ;
      q_arr_23_10 : IN std_logic ;
      q_arr_23_9 : IN std_logic ;
      q_arr_23_8 : IN std_logic ;
      q_arr_23_7 : IN std_logic ;
      q_arr_23_6 : IN std_logic ;
      q_arr_23_5 : IN std_logic ;
      q_arr_23_4 : IN std_logic ;
      q_arr_23_3 : IN std_logic ;
      q_arr_23_2 : IN std_logic ;
      q_arr_23_1 : IN std_logic ;
      q_arr_23_0 : IN std_logic ;
      q_arr_24_31 : IN std_logic ;
      q_arr_24_30 : IN std_logic ;
      q_arr_24_29 : IN std_logic ;
      q_arr_24_28 : IN std_logic ;
      q_arr_24_27 : IN std_logic ;
      q_arr_24_26 : IN std_logic ;
      q_arr_24_25 : IN std_logic ;
      q_arr_24_24 : IN std_logic ;
      q_arr_24_23 : IN std_logic ;
      q_arr_24_22 : IN std_logic ;
      q_arr_24_21 : IN std_logic ;
      q_arr_24_20 : IN std_logic ;
      q_arr_24_19 : IN std_logic ;
      q_arr_24_18 : IN std_logic ;
      q_arr_24_17 : IN std_logic ;
      q_arr_24_16 : IN std_logic ;
      q_arr_24_15 : IN std_logic ;
      q_arr_24_14 : IN std_logic ;
      q_arr_24_13 : IN std_logic ;
      q_arr_24_12 : IN std_logic ;
      q_arr_24_11 : IN std_logic ;
      q_arr_24_10 : IN std_logic ;
      q_arr_24_9 : IN std_logic ;
      q_arr_24_8 : IN std_logic ;
      q_arr_24_7 : IN std_logic ;
      q_arr_24_6 : IN std_logic ;
      q_arr_24_5 : IN std_logic ;
      q_arr_24_4 : IN std_logic ;
      q_arr_24_3 : IN std_logic ;
      q_arr_24_2 : IN std_logic ;
      q_arr_24_1 : IN std_logic ;
      q_arr_24_0 : IN std_logic) ;
end ReluLayer ;

architecture Structural_unfold_3309_0 of ReluLayer is
   signal d_arr_24_0_EXMPLR, nx205, nx207, nx209, nx211, nx213, nx215, nx217, 
      nx219, nx221, nx223, nx225, nx227: std_logic ;

begin
   d_arr_0_15 <= d_arr_24_0_EXMPLR ;
   d_arr_1_15 <= d_arr_24_0_EXMPLR ;
   d_arr_2_31 <= d_arr_24_0_EXMPLR ;
   d_arr_2_30 <= d_arr_24_0_EXMPLR ;
   d_arr_2_29 <= d_arr_24_0_EXMPLR ;
   d_arr_2_28 <= d_arr_24_0_EXMPLR ;
   d_arr_2_27 <= d_arr_24_0_EXMPLR ;
   d_arr_2_26 <= d_arr_24_0_EXMPLR ;
   d_arr_2_25 <= d_arr_24_0_EXMPLR ;
   d_arr_2_24 <= d_arr_24_0_EXMPLR ;
   d_arr_2_23 <= d_arr_24_0_EXMPLR ;
   d_arr_2_22 <= d_arr_24_0_EXMPLR ;
   d_arr_2_21 <= d_arr_24_0_EXMPLR ;
   d_arr_2_20 <= d_arr_24_0_EXMPLR ;
   d_arr_2_19 <= d_arr_24_0_EXMPLR ;
   d_arr_2_18 <= d_arr_24_0_EXMPLR ;
   d_arr_2_17 <= d_arr_24_0_EXMPLR ;
   d_arr_2_16 <= d_arr_24_0_EXMPLR ;
   d_arr_2_15 <= d_arr_24_0_EXMPLR ;
   d_arr_2_14 <= d_arr_24_0_EXMPLR ;
   d_arr_2_13 <= d_arr_24_0_EXMPLR ;
   d_arr_2_12 <= d_arr_24_0_EXMPLR ;
   d_arr_2_11 <= d_arr_24_0_EXMPLR ;
   d_arr_2_10 <= d_arr_24_0_EXMPLR ;
   d_arr_2_9 <= d_arr_24_0_EXMPLR ;
   d_arr_2_8 <= d_arr_24_0_EXMPLR ;
   d_arr_2_7 <= d_arr_24_0_EXMPLR ;
   d_arr_2_6 <= d_arr_24_0_EXMPLR ;
   d_arr_2_5 <= d_arr_24_0_EXMPLR ;
   d_arr_2_4 <= d_arr_24_0_EXMPLR ;
   d_arr_2_3 <= d_arr_24_0_EXMPLR ;
   d_arr_2_2 <= d_arr_24_0_EXMPLR ;
   d_arr_2_1 <= d_arr_24_0_EXMPLR ;
   d_arr_2_0 <= d_arr_24_0_EXMPLR ;
   d_arr_3_31 <= d_arr_24_0_EXMPLR ;
   d_arr_3_30 <= d_arr_24_0_EXMPLR ;
   d_arr_3_29 <= d_arr_24_0_EXMPLR ;
   d_arr_3_28 <= d_arr_24_0_EXMPLR ;
   d_arr_3_27 <= d_arr_24_0_EXMPLR ;
   d_arr_3_26 <= d_arr_24_0_EXMPLR ;
   d_arr_3_25 <= d_arr_24_0_EXMPLR ;
   d_arr_3_24 <= d_arr_24_0_EXMPLR ;
   d_arr_3_23 <= d_arr_24_0_EXMPLR ;
   d_arr_3_22 <= d_arr_24_0_EXMPLR ;
   d_arr_3_21 <= d_arr_24_0_EXMPLR ;
   d_arr_3_20 <= d_arr_24_0_EXMPLR ;
   d_arr_3_19 <= d_arr_24_0_EXMPLR ;
   d_arr_3_18 <= d_arr_24_0_EXMPLR ;
   d_arr_3_17 <= d_arr_24_0_EXMPLR ;
   d_arr_3_16 <= d_arr_24_0_EXMPLR ;
   d_arr_3_15 <= d_arr_24_0_EXMPLR ;
   d_arr_3_14 <= d_arr_24_0_EXMPLR ;
   d_arr_3_13 <= d_arr_24_0_EXMPLR ;
   d_arr_3_12 <= d_arr_24_0_EXMPLR ;
   d_arr_3_11 <= d_arr_24_0_EXMPLR ;
   d_arr_3_10 <= d_arr_24_0_EXMPLR ;
   d_arr_3_9 <= d_arr_24_0_EXMPLR ;
   d_arr_3_8 <= d_arr_24_0_EXMPLR ;
   d_arr_3_7 <= d_arr_24_0_EXMPLR ;
   d_arr_3_6 <= d_arr_24_0_EXMPLR ;
   d_arr_3_5 <= d_arr_24_0_EXMPLR ;
   d_arr_3_4 <= d_arr_24_0_EXMPLR ;
   d_arr_3_3 <= d_arr_24_0_EXMPLR ;
   d_arr_3_2 <= d_arr_24_0_EXMPLR ;
   d_arr_3_1 <= d_arr_24_0_EXMPLR ;
   d_arr_3_0 <= d_arr_24_0_EXMPLR ;
   d_arr_4_31 <= d_arr_24_0_EXMPLR ;
   d_arr_4_30 <= d_arr_24_0_EXMPLR ;
   d_arr_4_29 <= d_arr_24_0_EXMPLR ;
   d_arr_4_28 <= d_arr_24_0_EXMPLR ;
   d_arr_4_27 <= d_arr_24_0_EXMPLR ;
   d_arr_4_26 <= d_arr_24_0_EXMPLR ;
   d_arr_4_25 <= d_arr_24_0_EXMPLR ;
   d_arr_4_24 <= d_arr_24_0_EXMPLR ;
   d_arr_4_23 <= d_arr_24_0_EXMPLR ;
   d_arr_4_22 <= d_arr_24_0_EXMPLR ;
   d_arr_4_21 <= d_arr_24_0_EXMPLR ;
   d_arr_4_20 <= d_arr_24_0_EXMPLR ;
   d_arr_4_19 <= d_arr_24_0_EXMPLR ;
   d_arr_4_18 <= d_arr_24_0_EXMPLR ;
   d_arr_4_17 <= d_arr_24_0_EXMPLR ;
   d_arr_4_16 <= d_arr_24_0_EXMPLR ;
   d_arr_4_15 <= d_arr_24_0_EXMPLR ;
   d_arr_4_14 <= d_arr_24_0_EXMPLR ;
   d_arr_4_13 <= d_arr_24_0_EXMPLR ;
   d_arr_4_12 <= d_arr_24_0_EXMPLR ;
   d_arr_4_11 <= d_arr_24_0_EXMPLR ;
   d_arr_4_10 <= d_arr_24_0_EXMPLR ;
   d_arr_4_9 <= d_arr_24_0_EXMPLR ;
   d_arr_4_8 <= d_arr_24_0_EXMPLR ;
   d_arr_4_7 <= d_arr_24_0_EXMPLR ;
   d_arr_4_6 <= d_arr_24_0_EXMPLR ;
   d_arr_4_5 <= d_arr_24_0_EXMPLR ;
   d_arr_4_4 <= d_arr_24_0_EXMPLR ;
   d_arr_4_3 <= d_arr_24_0_EXMPLR ;
   d_arr_4_2 <= d_arr_24_0_EXMPLR ;
   d_arr_4_1 <= d_arr_24_0_EXMPLR ;
   d_arr_4_0 <= d_arr_24_0_EXMPLR ;
   d_arr_5_31 <= d_arr_24_0_EXMPLR ;
   d_arr_5_30 <= d_arr_24_0_EXMPLR ;
   d_arr_5_29 <= d_arr_24_0_EXMPLR ;
   d_arr_5_28 <= d_arr_24_0_EXMPLR ;
   d_arr_5_27 <= d_arr_24_0_EXMPLR ;
   d_arr_5_26 <= d_arr_24_0_EXMPLR ;
   d_arr_5_25 <= d_arr_24_0_EXMPLR ;
   d_arr_5_24 <= d_arr_24_0_EXMPLR ;
   d_arr_5_23 <= d_arr_24_0_EXMPLR ;
   d_arr_5_22 <= d_arr_24_0_EXMPLR ;
   d_arr_5_21 <= d_arr_24_0_EXMPLR ;
   d_arr_5_20 <= d_arr_24_0_EXMPLR ;
   d_arr_5_19 <= d_arr_24_0_EXMPLR ;
   d_arr_5_18 <= d_arr_24_0_EXMPLR ;
   d_arr_5_17 <= d_arr_24_0_EXMPLR ;
   d_arr_5_16 <= d_arr_24_0_EXMPLR ;
   d_arr_5_15 <= d_arr_24_0_EXMPLR ;
   d_arr_5_14 <= d_arr_24_0_EXMPLR ;
   d_arr_5_13 <= d_arr_24_0_EXMPLR ;
   d_arr_5_12 <= d_arr_24_0_EXMPLR ;
   d_arr_5_11 <= d_arr_24_0_EXMPLR ;
   d_arr_5_10 <= d_arr_24_0_EXMPLR ;
   d_arr_5_9 <= d_arr_24_0_EXMPLR ;
   d_arr_5_8 <= d_arr_24_0_EXMPLR ;
   d_arr_5_7 <= d_arr_24_0_EXMPLR ;
   d_arr_5_6 <= d_arr_24_0_EXMPLR ;
   d_arr_5_5 <= d_arr_24_0_EXMPLR ;
   d_arr_5_4 <= d_arr_24_0_EXMPLR ;
   d_arr_5_3 <= d_arr_24_0_EXMPLR ;
   d_arr_5_2 <= d_arr_24_0_EXMPLR ;
   d_arr_5_1 <= d_arr_24_0_EXMPLR ;
   d_arr_5_0 <= d_arr_24_0_EXMPLR ;
   d_arr_6_31 <= d_arr_24_0_EXMPLR ;
   d_arr_6_30 <= d_arr_24_0_EXMPLR ;
   d_arr_6_29 <= d_arr_24_0_EXMPLR ;
   d_arr_6_28 <= d_arr_24_0_EXMPLR ;
   d_arr_6_27 <= d_arr_24_0_EXMPLR ;
   d_arr_6_26 <= d_arr_24_0_EXMPLR ;
   d_arr_6_25 <= d_arr_24_0_EXMPLR ;
   d_arr_6_24 <= d_arr_24_0_EXMPLR ;
   d_arr_6_23 <= d_arr_24_0_EXMPLR ;
   d_arr_6_22 <= d_arr_24_0_EXMPLR ;
   d_arr_6_21 <= d_arr_24_0_EXMPLR ;
   d_arr_6_20 <= d_arr_24_0_EXMPLR ;
   d_arr_6_19 <= d_arr_24_0_EXMPLR ;
   d_arr_6_18 <= d_arr_24_0_EXMPLR ;
   d_arr_6_17 <= d_arr_24_0_EXMPLR ;
   d_arr_6_16 <= d_arr_24_0_EXMPLR ;
   d_arr_6_15 <= d_arr_24_0_EXMPLR ;
   d_arr_6_14 <= d_arr_24_0_EXMPLR ;
   d_arr_6_13 <= d_arr_24_0_EXMPLR ;
   d_arr_6_12 <= d_arr_24_0_EXMPLR ;
   d_arr_6_11 <= d_arr_24_0_EXMPLR ;
   d_arr_6_10 <= d_arr_24_0_EXMPLR ;
   d_arr_6_9 <= d_arr_24_0_EXMPLR ;
   d_arr_6_8 <= d_arr_24_0_EXMPLR ;
   d_arr_6_7 <= d_arr_24_0_EXMPLR ;
   d_arr_6_6 <= d_arr_24_0_EXMPLR ;
   d_arr_6_5 <= d_arr_24_0_EXMPLR ;
   d_arr_6_4 <= d_arr_24_0_EXMPLR ;
   d_arr_6_3 <= d_arr_24_0_EXMPLR ;
   d_arr_6_2 <= d_arr_24_0_EXMPLR ;
   d_arr_6_1 <= d_arr_24_0_EXMPLR ;
   d_arr_6_0 <= d_arr_24_0_EXMPLR ;
   d_arr_7_31 <= d_arr_24_0_EXMPLR ;
   d_arr_7_30 <= d_arr_24_0_EXMPLR ;
   d_arr_7_29 <= d_arr_24_0_EXMPLR ;
   d_arr_7_28 <= d_arr_24_0_EXMPLR ;
   d_arr_7_27 <= d_arr_24_0_EXMPLR ;
   d_arr_7_26 <= d_arr_24_0_EXMPLR ;
   d_arr_7_25 <= d_arr_24_0_EXMPLR ;
   d_arr_7_24 <= d_arr_24_0_EXMPLR ;
   d_arr_7_23 <= d_arr_24_0_EXMPLR ;
   d_arr_7_22 <= d_arr_24_0_EXMPLR ;
   d_arr_7_21 <= d_arr_24_0_EXMPLR ;
   d_arr_7_20 <= d_arr_24_0_EXMPLR ;
   d_arr_7_19 <= d_arr_24_0_EXMPLR ;
   d_arr_7_18 <= d_arr_24_0_EXMPLR ;
   d_arr_7_17 <= d_arr_24_0_EXMPLR ;
   d_arr_7_16 <= d_arr_24_0_EXMPLR ;
   d_arr_7_15 <= d_arr_24_0_EXMPLR ;
   d_arr_7_14 <= d_arr_24_0_EXMPLR ;
   d_arr_7_13 <= d_arr_24_0_EXMPLR ;
   d_arr_7_12 <= d_arr_24_0_EXMPLR ;
   d_arr_7_11 <= d_arr_24_0_EXMPLR ;
   d_arr_7_10 <= d_arr_24_0_EXMPLR ;
   d_arr_7_9 <= d_arr_24_0_EXMPLR ;
   d_arr_7_8 <= d_arr_24_0_EXMPLR ;
   d_arr_7_7 <= d_arr_24_0_EXMPLR ;
   d_arr_7_6 <= d_arr_24_0_EXMPLR ;
   d_arr_7_5 <= d_arr_24_0_EXMPLR ;
   d_arr_7_4 <= d_arr_24_0_EXMPLR ;
   d_arr_7_3 <= d_arr_24_0_EXMPLR ;
   d_arr_7_2 <= d_arr_24_0_EXMPLR ;
   d_arr_7_1 <= d_arr_24_0_EXMPLR ;
   d_arr_7_0 <= d_arr_24_0_EXMPLR ;
   d_arr_8_31 <= d_arr_24_0_EXMPLR ;
   d_arr_8_30 <= d_arr_24_0_EXMPLR ;
   d_arr_8_29 <= d_arr_24_0_EXMPLR ;
   d_arr_8_28 <= d_arr_24_0_EXMPLR ;
   d_arr_8_27 <= d_arr_24_0_EXMPLR ;
   d_arr_8_26 <= d_arr_24_0_EXMPLR ;
   d_arr_8_25 <= d_arr_24_0_EXMPLR ;
   d_arr_8_24 <= d_arr_24_0_EXMPLR ;
   d_arr_8_23 <= d_arr_24_0_EXMPLR ;
   d_arr_8_22 <= d_arr_24_0_EXMPLR ;
   d_arr_8_21 <= d_arr_24_0_EXMPLR ;
   d_arr_8_20 <= d_arr_24_0_EXMPLR ;
   d_arr_8_19 <= d_arr_24_0_EXMPLR ;
   d_arr_8_18 <= d_arr_24_0_EXMPLR ;
   d_arr_8_17 <= d_arr_24_0_EXMPLR ;
   d_arr_8_16 <= d_arr_24_0_EXMPLR ;
   d_arr_8_15 <= d_arr_24_0_EXMPLR ;
   d_arr_8_14 <= d_arr_24_0_EXMPLR ;
   d_arr_8_13 <= d_arr_24_0_EXMPLR ;
   d_arr_8_12 <= d_arr_24_0_EXMPLR ;
   d_arr_8_11 <= d_arr_24_0_EXMPLR ;
   d_arr_8_10 <= d_arr_24_0_EXMPLR ;
   d_arr_8_9 <= d_arr_24_0_EXMPLR ;
   d_arr_8_8 <= d_arr_24_0_EXMPLR ;
   d_arr_8_7 <= d_arr_24_0_EXMPLR ;
   d_arr_8_6 <= d_arr_24_0_EXMPLR ;
   d_arr_8_5 <= d_arr_24_0_EXMPLR ;
   d_arr_8_4 <= d_arr_24_0_EXMPLR ;
   d_arr_8_3 <= d_arr_24_0_EXMPLR ;
   d_arr_8_2 <= d_arr_24_0_EXMPLR ;
   d_arr_8_1 <= d_arr_24_0_EXMPLR ;
   d_arr_8_0 <= d_arr_24_0_EXMPLR ;
   d_arr_9_31 <= d_arr_24_0_EXMPLR ;
   d_arr_9_30 <= d_arr_24_0_EXMPLR ;
   d_arr_9_29 <= d_arr_24_0_EXMPLR ;
   d_arr_9_28 <= d_arr_24_0_EXMPLR ;
   d_arr_9_27 <= d_arr_24_0_EXMPLR ;
   d_arr_9_26 <= d_arr_24_0_EXMPLR ;
   d_arr_9_25 <= d_arr_24_0_EXMPLR ;
   d_arr_9_24 <= d_arr_24_0_EXMPLR ;
   d_arr_9_23 <= d_arr_24_0_EXMPLR ;
   d_arr_9_22 <= d_arr_24_0_EXMPLR ;
   d_arr_9_21 <= d_arr_24_0_EXMPLR ;
   d_arr_9_20 <= d_arr_24_0_EXMPLR ;
   d_arr_9_19 <= d_arr_24_0_EXMPLR ;
   d_arr_9_18 <= d_arr_24_0_EXMPLR ;
   d_arr_9_17 <= d_arr_24_0_EXMPLR ;
   d_arr_9_16 <= d_arr_24_0_EXMPLR ;
   d_arr_9_15 <= d_arr_24_0_EXMPLR ;
   d_arr_9_14 <= d_arr_24_0_EXMPLR ;
   d_arr_9_13 <= d_arr_24_0_EXMPLR ;
   d_arr_9_12 <= d_arr_24_0_EXMPLR ;
   d_arr_9_11 <= d_arr_24_0_EXMPLR ;
   d_arr_9_10 <= d_arr_24_0_EXMPLR ;
   d_arr_9_9 <= d_arr_24_0_EXMPLR ;
   d_arr_9_8 <= d_arr_24_0_EXMPLR ;
   d_arr_9_7 <= d_arr_24_0_EXMPLR ;
   d_arr_9_6 <= d_arr_24_0_EXMPLR ;
   d_arr_9_5 <= d_arr_24_0_EXMPLR ;
   d_arr_9_4 <= d_arr_24_0_EXMPLR ;
   d_arr_9_3 <= d_arr_24_0_EXMPLR ;
   d_arr_9_2 <= d_arr_24_0_EXMPLR ;
   d_arr_9_1 <= d_arr_24_0_EXMPLR ;
   d_arr_9_0 <= d_arr_24_0_EXMPLR ;
   d_arr_10_31 <= d_arr_24_0_EXMPLR ;
   d_arr_10_30 <= d_arr_24_0_EXMPLR ;
   d_arr_10_29 <= d_arr_24_0_EXMPLR ;
   d_arr_10_28 <= d_arr_24_0_EXMPLR ;
   d_arr_10_27 <= d_arr_24_0_EXMPLR ;
   d_arr_10_26 <= d_arr_24_0_EXMPLR ;
   d_arr_10_25 <= d_arr_24_0_EXMPLR ;
   d_arr_10_24 <= d_arr_24_0_EXMPLR ;
   d_arr_10_23 <= d_arr_24_0_EXMPLR ;
   d_arr_10_22 <= d_arr_24_0_EXMPLR ;
   d_arr_10_21 <= d_arr_24_0_EXMPLR ;
   d_arr_10_20 <= d_arr_24_0_EXMPLR ;
   d_arr_10_19 <= d_arr_24_0_EXMPLR ;
   d_arr_10_18 <= d_arr_24_0_EXMPLR ;
   d_arr_10_17 <= d_arr_24_0_EXMPLR ;
   d_arr_10_16 <= d_arr_24_0_EXMPLR ;
   d_arr_10_15 <= d_arr_24_0_EXMPLR ;
   d_arr_10_14 <= d_arr_24_0_EXMPLR ;
   d_arr_10_13 <= d_arr_24_0_EXMPLR ;
   d_arr_10_12 <= d_arr_24_0_EXMPLR ;
   d_arr_10_11 <= d_arr_24_0_EXMPLR ;
   d_arr_10_10 <= d_arr_24_0_EXMPLR ;
   d_arr_10_9 <= d_arr_24_0_EXMPLR ;
   d_arr_10_8 <= d_arr_24_0_EXMPLR ;
   d_arr_10_7 <= d_arr_24_0_EXMPLR ;
   d_arr_10_6 <= d_arr_24_0_EXMPLR ;
   d_arr_10_5 <= d_arr_24_0_EXMPLR ;
   d_arr_10_4 <= d_arr_24_0_EXMPLR ;
   d_arr_10_3 <= d_arr_24_0_EXMPLR ;
   d_arr_10_2 <= d_arr_24_0_EXMPLR ;
   d_arr_10_1 <= d_arr_24_0_EXMPLR ;
   d_arr_10_0 <= d_arr_24_0_EXMPLR ;
   d_arr_11_31 <= d_arr_24_0_EXMPLR ;
   d_arr_11_30 <= d_arr_24_0_EXMPLR ;
   d_arr_11_29 <= d_arr_24_0_EXMPLR ;
   d_arr_11_28 <= d_arr_24_0_EXMPLR ;
   d_arr_11_27 <= d_arr_24_0_EXMPLR ;
   d_arr_11_26 <= d_arr_24_0_EXMPLR ;
   d_arr_11_25 <= d_arr_24_0_EXMPLR ;
   d_arr_11_24 <= d_arr_24_0_EXMPLR ;
   d_arr_11_23 <= d_arr_24_0_EXMPLR ;
   d_arr_11_22 <= d_arr_24_0_EXMPLR ;
   d_arr_11_21 <= d_arr_24_0_EXMPLR ;
   d_arr_11_20 <= d_arr_24_0_EXMPLR ;
   d_arr_11_19 <= d_arr_24_0_EXMPLR ;
   d_arr_11_18 <= d_arr_24_0_EXMPLR ;
   d_arr_11_17 <= d_arr_24_0_EXMPLR ;
   d_arr_11_16 <= d_arr_24_0_EXMPLR ;
   d_arr_11_15 <= d_arr_24_0_EXMPLR ;
   d_arr_11_14 <= d_arr_24_0_EXMPLR ;
   d_arr_11_13 <= d_arr_24_0_EXMPLR ;
   d_arr_11_12 <= d_arr_24_0_EXMPLR ;
   d_arr_11_11 <= d_arr_24_0_EXMPLR ;
   d_arr_11_10 <= d_arr_24_0_EXMPLR ;
   d_arr_11_9 <= d_arr_24_0_EXMPLR ;
   d_arr_11_8 <= d_arr_24_0_EXMPLR ;
   d_arr_11_7 <= d_arr_24_0_EXMPLR ;
   d_arr_11_6 <= d_arr_24_0_EXMPLR ;
   d_arr_11_5 <= d_arr_24_0_EXMPLR ;
   d_arr_11_4 <= d_arr_24_0_EXMPLR ;
   d_arr_11_3 <= d_arr_24_0_EXMPLR ;
   d_arr_11_2 <= d_arr_24_0_EXMPLR ;
   d_arr_11_1 <= d_arr_24_0_EXMPLR ;
   d_arr_11_0 <= d_arr_24_0_EXMPLR ;
   d_arr_12_31 <= d_arr_24_0_EXMPLR ;
   d_arr_12_30 <= d_arr_24_0_EXMPLR ;
   d_arr_12_29 <= d_arr_24_0_EXMPLR ;
   d_arr_12_28 <= d_arr_24_0_EXMPLR ;
   d_arr_12_27 <= d_arr_24_0_EXMPLR ;
   d_arr_12_26 <= d_arr_24_0_EXMPLR ;
   d_arr_12_25 <= d_arr_24_0_EXMPLR ;
   d_arr_12_24 <= d_arr_24_0_EXMPLR ;
   d_arr_12_23 <= d_arr_24_0_EXMPLR ;
   d_arr_12_22 <= d_arr_24_0_EXMPLR ;
   d_arr_12_21 <= d_arr_24_0_EXMPLR ;
   d_arr_12_20 <= d_arr_24_0_EXMPLR ;
   d_arr_12_19 <= d_arr_24_0_EXMPLR ;
   d_arr_12_18 <= d_arr_24_0_EXMPLR ;
   d_arr_12_17 <= d_arr_24_0_EXMPLR ;
   d_arr_12_16 <= d_arr_24_0_EXMPLR ;
   d_arr_12_15 <= d_arr_24_0_EXMPLR ;
   d_arr_12_14 <= d_arr_24_0_EXMPLR ;
   d_arr_12_13 <= d_arr_24_0_EXMPLR ;
   d_arr_12_12 <= d_arr_24_0_EXMPLR ;
   d_arr_12_11 <= d_arr_24_0_EXMPLR ;
   d_arr_12_10 <= d_arr_24_0_EXMPLR ;
   d_arr_12_9 <= d_arr_24_0_EXMPLR ;
   d_arr_12_8 <= d_arr_24_0_EXMPLR ;
   d_arr_12_7 <= d_arr_24_0_EXMPLR ;
   d_arr_12_6 <= d_arr_24_0_EXMPLR ;
   d_arr_12_5 <= d_arr_24_0_EXMPLR ;
   d_arr_12_4 <= d_arr_24_0_EXMPLR ;
   d_arr_12_3 <= d_arr_24_0_EXMPLR ;
   d_arr_12_2 <= d_arr_24_0_EXMPLR ;
   d_arr_12_1 <= d_arr_24_0_EXMPLR ;
   d_arr_12_0 <= d_arr_24_0_EXMPLR ;
   d_arr_13_31 <= d_arr_24_0_EXMPLR ;
   d_arr_13_30 <= d_arr_24_0_EXMPLR ;
   d_arr_13_29 <= d_arr_24_0_EXMPLR ;
   d_arr_13_28 <= d_arr_24_0_EXMPLR ;
   d_arr_13_27 <= d_arr_24_0_EXMPLR ;
   d_arr_13_26 <= d_arr_24_0_EXMPLR ;
   d_arr_13_25 <= d_arr_24_0_EXMPLR ;
   d_arr_13_24 <= d_arr_24_0_EXMPLR ;
   d_arr_13_23 <= d_arr_24_0_EXMPLR ;
   d_arr_13_22 <= d_arr_24_0_EXMPLR ;
   d_arr_13_21 <= d_arr_24_0_EXMPLR ;
   d_arr_13_20 <= d_arr_24_0_EXMPLR ;
   d_arr_13_19 <= d_arr_24_0_EXMPLR ;
   d_arr_13_18 <= d_arr_24_0_EXMPLR ;
   d_arr_13_17 <= d_arr_24_0_EXMPLR ;
   d_arr_13_16 <= d_arr_24_0_EXMPLR ;
   d_arr_13_15 <= d_arr_24_0_EXMPLR ;
   d_arr_13_14 <= d_arr_24_0_EXMPLR ;
   d_arr_13_13 <= d_arr_24_0_EXMPLR ;
   d_arr_13_12 <= d_arr_24_0_EXMPLR ;
   d_arr_13_11 <= d_arr_24_0_EXMPLR ;
   d_arr_13_10 <= d_arr_24_0_EXMPLR ;
   d_arr_13_9 <= d_arr_24_0_EXMPLR ;
   d_arr_13_8 <= d_arr_24_0_EXMPLR ;
   d_arr_13_7 <= d_arr_24_0_EXMPLR ;
   d_arr_13_6 <= d_arr_24_0_EXMPLR ;
   d_arr_13_5 <= d_arr_24_0_EXMPLR ;
   d_arr_13_4 <= d_arr_24_0_EXMPLR ;
   d_arr_13_3 <= d_arr_24_0_EXMPLR ;
   d_arr_13_2 <= d_arr_24_0_EXMPLR ;
   d_arr_13_1 <= d_arr_24_0_EXMPLR ;
   d_arr_13_0 <= d_arr_24_0_EXMPLR ;
   d_arr_14_31 <= d_arr_24_0_EXMPLR ;
   d_arr_14_30 <= d_arr_24_0_EXMPLR ;
   d_arr_14_29 <= d_arr_24_0_EXMPLR ;
   d_arr_14_28 <= d_arr_24_0_EXMPLR ;
   d_arr_14_27 <= d_arr_24_0_EXMPLR ;
   d_arr_14_26 <= d_arr_24_0_EXMPLR ;
   d_arr_14_25 <= d_arr_24_0_EXMPLR ;
   d_arr_14_24 <= d_arr_24_0_EXMPLR ;
   d_arr_14_23 <= d_arr_24_0_EXMPLR ;
   d_arr_14_22 <= d_arr_24_0_EXMPLR ;
   d_arr_14_21 <= d_arr_24_0_EXMPLR ;
   d_arr_14_20 <= d_arr_24_0_EXMPLR ;
   d_arr_14_19 <= d_arr_24_0_EXMPLR ;
   d_arr_14_18 <= d_arr_24_0_EXMPLR ;
   d_arr_14_17 <= d_arr_24_0_EXMPLR ;
   d_arr_14_16 <= d_arr_24_0_EXMPLR ;
   d_arr_14_15 <= d_arr_24_0_EXMPLR ;
   d_arr_14_14 <= d_arr_24_0_EXMPLR ;
   d_arr_14_13 <= d_arr_24_0_EXMPLR ;
   d_arr_14_12 <= d_arr_24_0_EXMPLR ;
   d_arr_14_11 <= d_arr_24_0_EXMPLR ;
   d_arr_14_10 <= d_arr_24_0_EXMPLR ;
   d_arr_14_9 <= d_arr_24_0_EXMPLR ;
   d_arr_14_8 <= d_arr_24_0_EXMPLR ;
   d_arr_14_7 <= d_arr_24_0_EXMPLR ;
   d_arr_14_6 <= d_arr_24_0_EXMPLR ;
   d_arr_14_5 <= d_arr_24_0_EXMPLR ;
   d_arr_14_4 <= d_arr_24_0_EXMPLR ;
   d_arr_14_3 <= d_arr_24_0_EXMPLR ;
   d_arr_14_2 <= d_arr_24_0_EXMPLR ;
   d_arr_14_1 <= d_arr_24_0_EXMPLR ;
   d_arr_14_0 <= d_arr_24_0_EXMPLR ;
   d_arr_15_31 <= d_arr_24_0_EXMPLR ;
   d_arr_15_30 <= d_arr_24_0_EXMPLR ;
   d_arr_15_29 <= d_arr_24_0_EXMPLR ;
   d_arr_15_28 <= d_arr_24_0_EXMPLR ;
   d_arr_15_27 <= d_arr_24_0_EXMPLR ;
   d_arr_15_26 <= d_arr_24_0_EXMPLR ;
   d_arr_15_25 <= d_arr_24_0_EXMPLR ;
   d_arr_15_24 <= d_arr_24_0_EXMPLR ;
   d_arr_15_23 <= d_arr_24_0_EXMPLR ;
   d_arr_15_22 <= d_arr_24_0_EXMPLR ;
   d_arr_15_21 <= d_arr_24_0_EXMPLR ;
   d_arr_15_20 <= d_arr_24_0_EXMPLR ;
   d_arr_15_19 <= d_arr_24_0_EXMPLR ;
   d_arr_15_18 <= d_arr_24_0_EXMPLR ;
   d_arr_15_17 <= d_arr_24_0_EXMPLR ;
   d_arr_15_16 <= d_arr_24_0_EXMPLR ;
   d_arr_15_15 <= d_arr_24_0_EXMPLR ;
   d_arr_15_14 <= d_arr_24_0_EXMPLR ;
   d_arr_15_13 <= d_arr_24_0_EXMPLR ;
   d_arr_15_12 <= d_arr_24_0_EXMPLR ;
   d_arr_15_11 <= d_arr_24_0_EXMPLR ;
   d_arr_15_10 <= d_arr_24_0_EXMPLR ;
   d_arr_15_9 <= d_arr_24_0_EXMPLR ;
   d_arr_15_8 <= d_arr_24_0_EXMPLR ;
   d_arr_15_7 <= d_arr_24_0_EXMPLR ;
   d_arr_15_6 <= d_arr_24_0_EXMPLR ;
   d_arr_15_5 <= d_arr_24_0_EXMPLR ;
   d_arr_15_4 <= d_arr_24_0_EXMPLR ;
   d_arr_15_3 <= d_arr_24_0_EXMPLR ;
   d_arr_15_2 <= d_arr_24_0_EXMPLR ;
   d_arr_15_1 <= d_arr_24_0_EXMPLR ;
   d_arr_15_0 <= d_arr_24_0_EXMPLR ;
   d_arr_16_31 <= d_arr_24_0_EXMPLR ;
   d_arr_16_30 <= d_arr_24_0_EXMPLR ;
   d_arr_16_29 <= d_arr_24_0_EXMPLR ;
   d_arr_16_28 <= d_arr_24_0_EXMPLR ;
   d_arr_16_27 <= d_arr_24_0_EXMPLR ;
   d_arr_16_26 <= d_arr_24_0_EXMPLR ;
   d_arr_16_25 <= d_arr_24_0_EXMPLR ;
   d_arr_16_24 <= d_arr_24_0_EXMPLR ;
   d_arr_16_23 <= d_arr_24_0_EXMPLR ;
   d_arr_16_22 <= d_arr_24_0_EXMPLR ;
   d_arr_16_21 <= d_arr_24_0_EXMPLR ;
   d_arr_16_20 <= d_arr_24_0_EXMPLR ;
   d_arr_16_19 <= d_arr_24_0_EXMPLR ;
   d_arr_16_18 <= d_arr_24_0_EXMPLR ;
   d_arr_16_17 <= d_arr_24_0_EXMPLR ;
   d_arr_16_16 <= d_arr_24_0_EXMPLR ;
   d_arr_16_15 <= d_arr_24_0_EXMPLR ;
   d_arr_16_14 <= d_arr_24_0_EXMPLR ;
   d_arr_16_13 <= d_arr_24_0_EXMPLR ;
   d_arr_16_12 <= d_arr_24_0_EXMPLR ;
   d_arr_16_11 <= d_arr_24_0_EXMPLR ;
   d_arr_16_10 <= d_arr_24_0_EXMPLR ;
   d_arr_16_9 <= d_arr_24_0_EXMPLR ;
   d_arr_16_8 <= d_arr_24_0_EXMPLR ;
   d_arr_16_7 <= d_arr_24_0_EXMPLR ;
   d_arr_16_6 <= d_arr_24_0_EXMPLR ;
   d_arr_16_5 <= d_arr_24_0_EXMPLR ;
   d_arr_16_4 <= d_arr_24_0_EXMPLR ;
   d_arr_16_3 <= d_arr_24_0_EXMPLR ;
   d_arr_16_2 <= d_arr_24_0_EXMPLR ;
   d_arr_16_1 <= d_arr_24_0_EXMPLR ;
   d_arr_16_0 <= d_arr_24_0_EXMPLR ;
   d_arr_17_31 <= d_arr_24_0_EXMPLR ;
   d_arr_17_30 <= d_arr_24_0_EXMPLR ;
   d_arr_17_29 <= d_arr_24_0_EXMPLR ;
   d_arr_17_28 <= d_arr_24_0_EXMPLR ;
   d_arr_17_27 <= d_arr_24_0_EXMPLR ;
   d_arr_17_26 <= d_arr_24_0_EXMPLR ;
   d_arr_17_25 <= d_arr_24_0_EXMPLR ;
   d_arr_17_24 <= d_arr_24_0_EXMPLR ;
   d_arr_17_23 <= d_arr_24_0_EXMPLR ;
   d_arr_17_22 <= d_arr_24_0_EXMPLR ;
   d_arr_17_21 <= d_arr_24_0_EXMPLR ;
   d_arr_17_20 <= d_arr_24_0_EXMPLR ;
   d_arr_17_19 <= d_arr_24_0_EXMPLR ;
   d_arr_17_18 <= d_arr_24_0_EXMPLR ;
   d_arr_17_17 <= d_arr_24_0_EXMPLR ;
   d_arr_17_16 <= d_arr_24_0_EXMPLR ;
   d_arr_17_15 <= d_arr_24_0_EXMPLR ;
   d_arr_17_14 <= d_arr_24_0_EXMPLR ;
   d_arr_17_13 <= d_arr_24_0_EXMPLR ;
   d_arr_17_12 <= d_arr_24_0_EXMPLR ;
   d_arr_17_11 <= d_arr_24_0_EXMPLR ;
   d_arr_17_10 <= d_arr_24_0_EXMPLR ;
   d_arr_17_9 <= d_arr_24_0_EXMPLR ;
   d_arr_17_8 <= d_arr_24_0_EXMPLR ;
   d_arr_17_7 <= d_arr_24_0_EXMPLR ;
   d_arr_17_6 <= d_arr_24_0_EXMPLR ;
   d_arr_17_5 <= d_arr_24_0_EXMPLR ;
   d_arr_17_4 <= d_arr_24_0_EXMPLR ;
   d_arr_17_3 <= d_arr_24_0_EXMPLR ;
   d_arr_17_2 <= d_arr_24_0_EXMPLR ;
   d_arr_17_1 <= d_arr_24_0_EXMPLR ;
   d_arr_17_0 <= d_arr_24_0_EXMPLR ;
   d_arr_18_31 <= d_arr_24_0_EXMPLR ;
   d_arr_18_30 <= d_arr_24_0_EXMPLR ;
   d_arr_18_29 <= d_arr_24_0_EXMPLR ;
   d_arr_18_28 <= d_arr_24_0_EXMPLR ;
   d_arr_18_27 <= d_arr_24_0_EXMPLR ;
   d_arr_18_26 <= d_arr_24_0_EXMPLR ;
   d_arr_18_25 <= d_arr_24_0_EXMPLR ;
   d_arr_18_24 <= d_arr_24_0_EXMPLR ;
   d_arr_18_23 <= d_arr_24_0_EXMPLR ;
   d_arr_18_22 <= d_arr_24_0_EXMPLR ;
   d_arr_18_21 <= d_arr_24_0_EXMPLR ;
   d_arr_18_20 <= d_arr_24_0_EXMPLR ;
   d_arr_18_19 <= d_arr_24_0_EXMPLR ;
   d_arr_18_18 <= d_arr_24_0_EXMPLR ;
   d_arr_18_17 <= d_arr_24_0_EXMPLR ;
   d_arr_18_16 <= d_arr_24_0_EXMPLR ;
   d_arr_18_15 <= d_arr_24_0_EXMPLR ;
   d_arr_18_14 <= d_arr_24_0_EXMPLR ;
   d_arr_18_13 <= d_arr_24_0_EXMPLR ;
   d_arr_18_12 <= d_arr_24_0_EXMPLR ;
   d_arr_18_11 <= d_arr_24_0_EXMPLR ;
   d_arr_18_10 <= d_arr_24_0_EXMPLR ;
   d_arr_18_9 <= d_arr_24_0_EXMPLR ;
   d_arr_18_8 <= d_arr_24_0_EXMPLR ;
   d_arr_18_7 <= d_arr_24_0_EXMPLR ;
   d_arr_18_6 <= d_arr_24_0_EXMPLR ;
   d_arr_18_5 <= d_arr_24_0_EXMPLR ;
   d_arr_18_4 <= d_arr_24_0_EXMPLR ;
   d_arr_18_3 <= d_arr_24_0_EXMPLR ;
   d_arr_18_2 <= d_arr_24_0_EXMPLR ;
   d_arr_18_1 <= d_arr_24_0_EXMPLR ;
   d_arr_18_0 <= d_arr_24_0_EXMPLR ;
   d_arr_19_31 <= d_arr_24_0_EXMPLR ;
   d_arr_19_30 <= d_arr_24_0_EXMPLR ;
   d_arr_19_29 <= d_arr_24_0_EXMPLR ;
   d_arr_19_28 <= d_arr_24_0_EXMPLR ;
   d_arr_19_27 <= d_arr_24_0_EXMPLR ;
   d_arr_19_26 <= d_arr_24_0_EXMPLR ;
   d_arr_19_25 <= d_arr_24_0_EXMPLR ;
   d_arr_19_24 <= d_arr_24_0_EXMPLR ;
   d_arr_19_23 <= d_arr_24_0_EXMPLR ;
   d_arr_19_22 <= d_arr_24_0_EXMPLR ;
   d_arr_19_21 <= d_arr_24_0_EXMPLR ;
   d_arr_19_20 <= d_arr_24_0_EXMPLR ;
   d_arr_19_19 <= d_arr_24_0_EXMPLR ;
   d_arr_19_18 <= d_arr_24_0_EXMPLR ;
   d_arr_19_17 <= d_arr_24_0_EXMPLR ;
   d_arr_19_16 <= d_arr_24_0_EXMPLR ;
   d_arr_19_15 <= d_arr_24_0_EXMPLR ;
   d_arr_19_14 <= d_arr_24_0_EXMPLR ;
   d_arr_19_13 <= d_arr_24_0_EXMPLR ;
   d_arr_19_12 <= d_arr_24_0_EXMPLR ;
   d_arr_19_11 <= d_arr_24_0_EXMPLR ;
   d_arr_19_10 <= d_arr_24_0_EXMPLR ;
   d_arr_19_9 <= d_arr_24_0_EXMPLR ;
   d_arr_19_8 <= d_arr_24_0_EXMPLR ;
   d_arr_19_7 <= d_arr_24_0_EXMPLR ;
   d_arr_19_6 <= d_arr_24_0_EXMPLR ;
   d_arr_19_5 <= d_arr_24_0_EXMPLR ;
   d_arr_19_4 <= d_arr_24_0_EXMPLR ;
   d_arr_19_3 <= d_arr_24_0_EXMPLR ;
   d_arr_19_2 <= d_arr_24_0_EXMPLR ;
   d_arr_19_1 <= d_arr_24_0_EXMPLR ;
   d_arr_19_0 <= d_arr_24_0_EXMPLR ;
   d_arr_20_31 <= d_arr_24_0_EXMPLR ;
   d_arr_20_30 <= d_arr_24_0_EXMPLR ;
   d_arr_20_29 <= d_arr_24_0_EXMPLR ;
   d_arr_20_28 <= d_arr_24_0_EXMPLR ;
   d_arr_20_27 <= d_arr_24_0_EXMPLR ;
   d_arr_20_26 <= d_arr_24_0_EXMPLR ;
   d_arr_20_25 <= d_arr_24_0_EXMPLR ;
   d_arr_20_24 <= d_arr_24_0_EXMPLR ;
   d_arr_20_23 <= d_arr_24_0_EXMPLR ;
   d_arr_20_22 <= d_arr_24_0_EXMPLR ;
   d_arr_20_21 <= d_arr_24_0_EXMPLR ;
   d_arr_20_20 <= d_arr_24_0_EXMPLR ;
   d_arr_20_19 <= d_arr_24_0_EXMPLR ;
   d_arr_20_18 <= d_arr_24_0_EXMPLR ;
   d_arr_20_17 <= d_arr_24_0_EXMPLR ;
   d_arr_20_16 <= d_arr_24_0_EXMPLR ;
   d_arr_20_15 <= d_arr_24_0_EXMPLR ;
   d_arr_20_14 <= d_arr_24_0_EXMPLR ;
   d_arr_20_13 <= d_arr_24_0_EXMPLR ;
   d_arr_20_12 <= d_arr_24_0_EXMPLR ;
   d_arr_20_11 <= d_arr_24_0_EXMPLR ;
   d_arr_20_10 <= d_arr_24_0_EXMPLR ;
   d_arr_20_9 <= d_arr_24_0_EXMPLR ;
   d_arr_20_8 <= d_arr_24_0_EXMPLR ;
   d_arr_20_7 <= d_arr_24_0_EXMPLR ;
   d_arr_20_6 <= d_arr_24_0_EXMPLR ;
   d_arr_20_5 <= d_arr_24_0_EXMPLR ;
   d_arr_20_4 <= d_arr_24_0_EXMPLR ;
   d_arr_20_3 <= d_arr_24_0_EXMPLR ;
   d_arr_20_2 <= d_arr_24_0_EXMPLR ;
   d_arr_20_1 <= d_arr_24_0_EXMPLR ;
   d_arr_20_0 <= d_arr_24_0_EXMPLR ;
   d_arr_21_31 <= d_arr_24_0_EXMPLR ;
   d_arr_21_30 <= d_arr_24_0_EXMPLR ;
   d_arr_21_29 <= d_arr_24_0_EXMPLR ;
   d_arr_21_28 <= d_arr_24_0_EXMPLR ;
   d_arr_21_27 <= d_arr_24_0_EXMPLR ;
   d_arr_21_26 <= d_arr_24_0_EXMPLR ;
   d_arr_21_25 <= d_arr_24_0_EXMPLR ;
   d_arr_21_24 <= d_arr_24_0_EXMPLR ;
   d_arr_21_23 <= d_arr_24_0_EXMPLR ;
   d_arr_21_22 <= d_arr_24_0_EXMPLR ;
   d_arr_21_21 <= d_arr_24_0_EXMPLR ;
   d_arr_21_20 <= d_arr_24_0_EXMPLR ;
   d_arr_21_19 <= d_arr_24_0_EXMPLR ;
   d_arr_21_18 <= d_arr_24_0_EXMPLR ;
   d_arr_21_17 <= d_arr_24_0_EXMPLR ;
   d_arr_21_16 <= d_arr_24_0_EXMPLR ;
   d_arr_21_15 <= d_arr_24_0_EXMPLR ;
   d_arr_21_14 <= d_arr_24_0_EXMPLR ;
   d_arr_21_13 <= d_arr_24_0_EXMPLR ;
   d_arr_21_12 <= d_arr_24_0_EXMPLR ;
   d_arr_21_11 <= d_arr_24_0_EXMPLR ;
   d_arr_21_10 <= d_arr_24_0_EXMPLR ;
   d_arr_21_9 <= d_arr_24_0_EXMPLR ;
   d_arr_21_8 <= d_arr_24_0_EXMPLR ;
   d_arr_21_7 <= d_arr_24_0_EXMPLR ;
   d_arr_21_6 <= d_arr_24_0_EXMPLR ;
   d_arr_21_5 <= d_arr_24_0_EXMPLR ;
   d_arr_21_4 <= d_arr_24_0_EXMPLR ;
   d_arr_21_3 <= d_arr_24_0_EXMPLR ;
   d_arr_21_2 <= d_arr_24_0_EXMPLR ;
   d_arr_21_1 <= d_arr_24_0_EXMPLR ;
   d_arr_21_0 <= d_arr_24_0_EXMPLR ;
   d_arr_22_31 <= d_arr_24_0_EXMPLR ;
   d_arr_22_30 <= d_arr_24_0_EXMPLR ;
   d_arr_22_29 <= d_arr_24_0_EXMPLR ;
   d_arr_22_28 <= d_arr_24_0_EXMPLR ;
   d_arr_22_27 <= d_arr_24_0_EXMPLR ;
   d_arr_22_26 <= d_arr_24_0_EXMPLR ;
   d_arr_22_25 <= d_arr_24_0_EXMPLR ;
   d_arr_22_24 <= d_arr_24_0_EXMPLR ;
   d_arr_22_23 <= d_arr_24_0_EXMPLR ;
   d_arr_22_22 <= d_arr_24_0_EXMPLR ;
   d_arr_22_21 <= d_arr_24_0_EXMPLR ;
   d_arr_22_20 <= d_arr_24_0_EXMPLR ;
   d_arr_22_19 <= d_arr_24_0_EXMPLR ;
   d_arr_22_18 <= d_arr_24_0_EXMPLR ;
   d_arr_22_17 <= d_arr_24_0_EXMPLR ;
   d_arr_22_16 <= d_arr_24_0_EXMPLR ;
   d_arr_22_15 <= d_arr_24_0_EXMPLR ;
   d_arr_22_14 <= d_arr_24_0_EXMPLR ;
   d_arr_22_13 <= d_arr_24_0_EXMPLR ;
   d_arr_22_12 <= d_arr_24_0_EXMPLR ;
   d_arr_22_11 <= d_arr_24_0_EXMPLR ;
   d_arr_22_10 <= d_arr_24_0_EXMPLR ;
   d_arr_22_9 <= d_arr_24_0_EXMPLR ;
   d_arr_22_8 <= d_arr_24_0_EXMPLR ;
   d_arr_22_7 <= d_arr_24_0_EXMPLR ;
   d_arr_22_6 <= d_arr_24_0_EXMPLR ;
   d_arr_22_5 <= d_arr_24_0_EXMPLR ;
   d_arr_22_4 <= d_arr_24_0_EXMPLR ;
   d_arr_22_3 <= d_arr_24_0_EXMPLR ;
   d_arr_22_2 <= d_arr_24_0_EXMPLR ;
   d_arr_22_1 <= d_arr_24_0_EXMPLR ;
   d_arr_22_0 <= d_arr_24_0_EXMPLR ;
   d_arr_23_31 <= d_arr_24_0_EXMPLR ;
   d_arr_23_30 <= d_arr_24_0_EXMPLR ;
   d_arr_23_29 <= d_arr_24_0_EXMPLR ;
   d_arr_23_28 <= d_arr_24_0_EXMPLR ;
   d_arr_23_27 <= d_arr_24_0_EXMPLR ;
   d_arr_23_26 <= d_arr_24_0_EXMPLR ;
   d_arr_23_25 <= d_arr_24_0_EXMPLR ;
   d_arr_23_24 <= d_arr_24_0_EXMPLR ;
   d_arr_23_23 <= d_arr_24_0_EXMPLR ;
   d_arr_23_22 <= d_arr_24_0_EXMPLR ;
   d_arr_23_21 <= d_arr_24_0_EXMPLR ;
   d_arr_23_20 <= d_arr_24_0_EXMPLR ;
   d_arr_23_19 <= d_arr_24_0_EXMPLR ;
   d_arr_23_18 <= d_arr_24_0_EXMPLR ;
   d_arr_23_17 <= d_arr_24_0_EXMPLR ;
   d_arr_23_16 <= d_arr_24_0_EXMPLR ;
   d_arr_23_15 <= d_arr_24_0_EXMPLR ;
   d_arr_23_14 <= d_arr_24_0_EXMPLR ;
   d_arr_23_13 <= d_arr_24_0_EXMPLR ;
   d_arr_23_12 <= d_arr_24_0_EXMPLR ;
   d_arr_23_11 <= d_arr_24_0_EXMPLR ;
   d_arr_23_10 <= d_arr_24_0_EXMPLR ;
   d_arr_23_9 <= d_arr_24_0_EXMPLR ;
   d_arr_23_8 <= d_arr_24_0_EXMPLR ;
   d_arr_23_7 <= d_arr_24_0_EXMPLR ;
   d_arr_23_6 <= d_arr_24_0_EXMPLR ;
   d_arr_23_5 <= d_arr_24_0_EXMPLR ;
   d_arr_23_4 <= d_arr_24_0_EXMPLR ;
   d_arr_23_3 <= d_arr_24_0_EXMPLR ;
   d_arr_23_2 <= d_arr_24_0_EXMPLR ;
   d_arr_23_1 <= d_arr_24_0_EXMPLR ;
   d_arr_23_0 <= d_arr_24_0_EXMPLR ;
   d_arr_24_31 <= d_arr_24_0_EXMPLR ;
   d_arr_24_30 <= d_arr_24_0_EXMPLR ;
   d_arr_24_29 <= d_arr_24_0_EXMPLR ;
   d_arr_24_28 <= d_arr_24_0_EXMPLR ;
   d_arr_24_27 <= d_arr_24_0_EXMPLR ;
   d_arr_24_26 <= d_arr_24_0_EXMPLR ;
   d_arr_24_25 <= d_arr_24_0_EXMPLR ;
   d_arr_24_24 <= d_arr_24_0_EXMPLR ;
   d_arr_24_23 <= d_arr_24_0_EXMPLR ;
   d_arr_24_22 <= d_arr_24_0_EXMPLR ;
   d_arr_24_21 <= d_arr_24_0_EXMPLR ;
   d_arr_24_20 <= d_arr_24_0_EXMPLR ;
   d_arr_24_19 <= d_arr_24_0_EXMPLR ;
   d_arr_24_18 <= d_arr_24_0_EXMPLR ;
   d_arr_24_17 <= d_arr_24_0_EXMPLR ;
   d_arr_24_16 <= d_arr_24_0_EXMPLR ;
   d_arr_24_15 <= d_arr_24_0_EXMPLR ;
   d_arr_24_14 <= d_arr_24_0_EXMPLR ;
   d_arr_24_13 <= d_arr_24_0_EXMPLR ;
   d_arr_24_12 <= d_arr_24_0_EXMPLR ;
   d_arr_24_11 <= d_arr_24_0_EXMPLR ;
   d_arr_24_10 <= d_arr_24_0_EXMPLR ;
   d_arr_24_9 <= d_arr_24_0_EXMPLR ;
   d_arr_24_8 <= d_arr_24_0_EXMPLR ;
   d_arr_24_7 <= d_arr_24_0_EXMPLR ;
   d_arr_24_6 <= d_arr_24_0_EXMPLR ;
   d_arr_24_5 <= d_arr_24_0_EXMPLR ;
   d_arr_24_4 <= d_arr_24_0_EXMPLR ;
   d_arr_24_3 <= d_arr_24_0_EXMPLR ;
   d_arr_24_2 <= d_arr_24_0_EXMPLR ;
   d_arr_24_1 <= d_arr_24_0_EXMPLR ;
   d_arr_24_0 <= d_arr_24_0_EXMPLR ;
   ix42 : fake_gnd port map ( Y=>d_arr_24_0_EXMPLR);
   ix3 : nor02ii port map ( Y=>d_arr_1_0, A0=>nx219, A1=>q_arr_1_0);
   ix7 : nor02ii port map ( Y=>d_arr_1_1, A0=>nx219, A1=>q_arr_1_1);
   ix11 : nor02ii port map ( Y=>d_arr_1_2, A0=>nx219, A1=>q_arr_1_2);
   ix15 : nor02ii port map ( Y=>d_arr_1_3, A0=>nx219, A1=>q_arr_1_3);
   ix19 : nor02ii port map ( Y=>d_arr_1_4, A0=>nx219, A1=>q_arr_1_4);
   ix23 : nor02ii port map ( Y=>d_arr_1_5, A0=>nx219, A1=>q_arr_1_5);
   ix27 : nor02ii port map ( Y=>d_arr_1_6, A0=>nx219, A1=>q_arr_1_6);
   ix31 : nor02ii port map ( Y=>d_arr_1_7, A0=>nx221, A1=>q_arr_1_7);
   ix35 : nor02ii port map ( Y=>d_arr_1_8, A0=>nx221, A1=>q_arr_1_8);
   ix39 : nor02ii port map ( Y=>d_arr_1_9, A0=>nx221, A1=>q_arr_1_9);
   ix43 : nor02ii port map ( Y=>d_arr_1_10, A0=>nx221, A1=>q_arr_1_10);
   ix47 : nor02ii port map ( Y=>d_arr_1_11, A0=>nx221, A1=>q_arr_1_11);
   ix51 : nor02ii port map ( Y=>d_arr_1_12, A0=>nx221, A1=>q_arr_1_12);
   ix55 : nor02ii port map ( Y=>d_arr_1_13, A0=>nx221, A1=>q_arr_1_13);
   ix59 : nor02ii port map ( Y=>d_arr_1_14, A0=>nx223, A1=>q_arr_1_14);
   ix63 : nor02ii port map ( Y=>d_arr_1_16, A0=>nx223, A1=>q_arr_1_16);
   ix67 : nor02ii port map ( Y=>d_arr_1_17, A0=>nx223, A1=>q_arr_1_17);
   ix71 : nor02ii port map ( Y=>d_arr_1_18, A0=>nx223, A1=>q_arr_1_18);
   ix75 : nor02ii port map ( Y=>d_arr_1_19, A0=>nx223, A1=>q_arr_1_19);
   ix79 : nor02ii port map ( Y=>d_arr_1_20, A0=>nx223, A1=>q_arr_1_20);
   ix83 : nor02ii port map ( Y=>d_arr_1_21, A0=>nx223, A1=>q_arr_1_21);
   ix87 : nor02ii port map ( Y=>d_arr_1_22, A0=>nx225, A1=>q_arr_1_22);
   ix91 : nor02ii port map ( Y=>d_arr_1_23, A0=>nx225, A1=>q_arr_1_23);
   ix95 : nor02ii port map ( Y=>d_arr_1_24, A0=>nx225, A1=>q_arr_1_24);
   ix99 : nor02ii port map ( Y=>d_arr_1_25, A0=>nx225, A1=>q_arr_1_25);
   ix103 : nor02ii port map ( Y=>d_arr_1_26, A0=>nx225, A1=>q_arr_1_26);
   ix107 : nor02ii port map ( Y=>d_arr_1_27, A0=>nx225, A1=>q_arr_1_27);
   ix111 : nor02ii port map ( Y=>d_arr_1_28, A0=>nx225, A1=>q_arr_1_28);
   ix115 : nor02ii port map ( Y=>d_arr_1_29, A0=>nx227, A1=>q_arr_1_29);
   ix119 : nor02ii port map ( Y=>d_arr_1_30, A0=>nx227, A1=>q_arr_1_30);
   ix123 : nor02ii port map ( Y=>d_arr_1_31, A0=>nx227, A1=>q_arr_1_31);
   ix127 : nor02ii port map ( Y=>d_arr_0_0, A0=>nx207, A1=>q_arr_0_0);
   ix131 : nor02ii port map ( Y=>d_arr_0_1, A0=>nx207, A1=>q_arr_0_1);
   ix135 : nor02ii port map ( Y=>d_arr_0_2, A0=>nx207, A1=>q_arr_0_2);
   ix139 : nor02ii port map ( Y=>d_arr_0_3, A0=>nx207, A1=>q_arr_0_3);
   ix143 : nor02ii port map ( Y=>d_arr_0_4, A0=>nx207, A1=>q_arr_0_4);
   ix147 : nor02ii port map ( Y=>d_arr_0_5, A0=>nx207, A1=>q_arr_0_5);
   ix151 : nor02ii port map ( Y=>d_arr_0_6, A0=>nx207, A1=>q_arr_0_6);
   ix155 : nor02ii port map ( Y=>d_arr_0_7, A0=>nx209, A1=>q_arr_0_7);
   ix159 : nor02ii port map ( Y=>d_arr_0_8, A0=>nx209, A1=>q_arr_0_8);
   ix163 : nor02ii port map ( Y=>d_arr_0_9, A0=>nx209, A1=>q_arr_0_9);
   ix167 : nor02ii port map ( Y=>d_arr_0_10, A0=>nx209, A1=>q_arr_0_10);
   ix171 : nor02ii port map ( Y=>d_arr_0_11, A0=>nx209, A1=>q_arr_0_11);
   ix175 : nor02ii port map ( Y=>d_arr_0_12, A0=>nx209, A1=>q_arr_0_12);
   ix179 : nor02ii port map ( Y=>d_arr_0_13, A0=>nx209, A1=>q_arr_0_13);
   ix183 : nor02ii port map ( Y=>d_arr_0_14, A0=>nx211, A1=>q_arr_0_14);
   ix187 : nor02ii port map ( Y=>d_arr_0_16, A0=>nx211, A1=>q_arr_0_16);
   ix191 : nor02ii port map ( Y=>d_arr_0_17, A0=>nx211, A1=>q_arr_0_17);
   ix195 : nor02ii port map ( Y=>d_arr_0_18, A0=>nx211, A1=>q_arr_0_18);
   ix199 : nor02ii port map ( Y=>d_arr_0_19, A0=>nx211, A1=>q_arr_0_19);
   ix203 : nor02ii port map ( Y=>d_arr_0_20, A0=>nx211, A1=>q_arr_0_20);
   ix207 : nor02ii port map ( Y=>d_arr_0_21, A0=>nx211, A1=>q_arr_0_21);
   ix211 : nor02ii port map ( Y=>d_arr_0_22, A0=>nx213, A1=>q_arr_0_22);
   ix215 : nor02ii port map ( Y=>d_arr_0_23, A0=>nx213, A1=>q_arr_0_23);
   ix219 : nor02ii port map ( Y=>d_arr_0_24, A0=>nx213, A1=>q_arr_0_24);
   ix223 : nor02ii port map ( Y=>d_arr_0_25, A0=>nx213, A1=>q_arr_0_25);
   ix227 : nor02ii port map ( Y=>d_arr_0_26, A0=>nx213, A1=>q_arr_0_26);
   ix231 : nor02ii port map ( Y=>d_arr_0_27, A0=>nx213, A1=>q_arr_0_27);
   ix235 : nor02ii port map ( Y=>d_arr_0_28, A0=>nx213, A1=>q_arr_0_28);
   ix239 : nor02ii port map ( Y=>d_arr_0_29, A0=>nx215, A1=>q_arr_0_29);
   ix243 : nor02ii port map ( Y=>d_arr_0_30, A0=>nx215, A1=>q_arr_0_30);
   ix247 : nor02ii port map ( Y=>d_arr_0_31, A0=>nx215, A1=>q_arr_0_31);
   ix204 : inv01 port map ( Y=>nx205, A=>q_arr_0_15);
   ix206 : inv01 port map ( Y=>nx207, A=>nx205);
   ix208 : inv01 port map ( Y=>nx209, A=>nx205);
   ix210 : inv01 port map ( Y=>nx211, A=>nx205);
   ix212 : inv01 port map ( Y=>nx213, A=>nx205);
   ix214 : inv01 port map ( Y=>nx215, A=>nx205);
   ix216 : inv01 port map ( Y=>nx217, A=>q_arr_1_15);
   ix218 : inv01 port map ( Y=>nx219, A=>nx217);
   ix220 : inv01 port map ( Y=>nx221, A=>nx217);
   ix222 : inv01 port map ( Y=>nx223, A=>nx217);
   ix224 : inv01 port map ( Y=>nx225, A=>nx217);
   ix226 : inv01 port map ( Y=>nx227, A=>nx217);
end Structural_unfold_3309_0 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity ModifiedBoothMultiplier is
   port (
      M : IN std_logic_vector (15 DOWNTO 0) ;
      R : IN std_logic_vector (15 DOWNTO 0) ;
      cnt_enable : IN std_logic ;
      product : OUT std_logic_vector (31 DOWNTO 0) ;
      clk : IN std_logic) ;
end ModifiedBoothMultiplier ;

architecture ModifiedBoothMultiplierWorkFlow of ModifiedBoothMultiplier is
   signal aux_product_0, shifting_R_0, shifting_R_4, shifting_R_6, 
      shifting_R_8, shifting_R_10, shifting_R_12, shifting_R_14, 
      shifting_R_16, nx30, nx40, nx50, nx60, nx70, nx80, nx90, nx100, nx108, 
      shifting_R_1, shifting_R_3, shifting_R_5, shifting_R_7, shifting_R_9, 
      shifting_R_11, shifting_R_13, shifting_R_15, nx146, nx156, nx166, 
      nx176, nx186, nx196, nx206, nx216, nx228, nx254, positive_2M_1, nx258, 
      nx268, nx270, aux_product_1, negative_M_1, nx296, nx306, nx310, 
      positive_M_1, nx338, nx350, nx354, nx370, aux_product_2, positive_M_2, 
      nx398, nx406, nx426, negative_M_2, nx442, nx464, aux_product_3, 
      positive_M_3, nx500, nx508, nx520, negative_M_3, nx536, nx552, nx558, 
      aux_product_4, positive_M_4, nx614, negative_M_4, nx630, nx646, nx652, 
      aux_product_5, positive_M_5, nx708, negative_M_5, nx724, nx740, nx746, 
      aux_product_6, positive_M_6, nx802, negative_M_6, nx818, nx834, nx840, 
      aux_product_7, positive_M_7, nx896, negative_M_7, nx912, nx934, 
      aux_product_8, positive_M_8, nx990, negative_M_8, nx1006, nx1028, 
      aux_product_9, positive_M_9, nx1084, negative_M_9, nx1100, nx1122, 
      aux_product_10, positive_M_10, nx1150, nx1178, negative_M_10, nx1194, 
      nx1216, aux_product_11, positive_M_11, nx1272, negative_M_11, nx1288, 
      nx1308, nx1310, aux_product_12, positive_M_12, nx1366, negative_M_12, 
      nx1382, nx1404, aux_product_13, positive_M_13, nx1460, negative_M_13, 
      nx1476, nx1498, aux_product_14, positive_M_14, nx1526, nx1554, 
      negative_M_14, nx1570, nx1592, aux_product_15, positive_M_15, nx1616, 
      nx1624, negative_M_15, nx1640, nx1656, nx1660, nx1662, aux_product_16, 
      positive_M_16, nx1694, negative_M_16, nx1710, nx1726, nx1732, 
      aux_product_17, positive_M_17, nx1758, negative_M_17, nx1770, nx1792, 
      aux_product_18, positive_M_18, nx1818, negative_M_18, nx1830, nx1852, 
      aux_product_19, positive_M_19, nx1878, negative_M_19, nx1890, nx1906, 
      nx1912, aux_product_20, positive_M_20, nx1938, negative_M_20, nx1950, 
      nx1966, nx1972, aux_product_21, positive_M_21, nx1998, negative_M_21, 
      nx2010, nx2026, nx2032, aux_product_22, positive_M_22, nx2058, 
      negative_M_22, nx2070, nx2090, nx2092, aux_product_23, positive_M_23, 
      nx2118, negative_M_23, nx2130, aux_product_24, positive_M_24, nx2178, 
      negative_M_24, nx2190, nx2206, nx2210, aux_product_25, positive_M_25, 
      nx2238, negative_M_25, nx2250, nx2272, aux_product_26, positive_M_26, 
      nx2298, negative_M_26, nx2310, aux_product_27, positive_M_27, nx2358, 
      negative_M_27, nx2370, nx2386, nx2390, aux_product_28, positive_M_28, 
      nx2418, negative_M_28, nx2430, nx2446, aux_product_29, positive_M_29, 
      nx2478, negative_M_29, nx2490, nx2506, nx2510, aux_product_30, 
      positive_2M_31, nx2538, negative_2M_31, nx2550, nx2566, nx2570, 
      aux_product_31, positive_M_31, nx2598, negative_M_31, nx2610, nx2626, 
      nx2630, nx3098, nx3108, nx3118, nx3128, nx3138, nx3148, nx3158, nx3168, 
      nx3178, nx3188, nx3198, nx3208, nx3218, nx3228, nx3238, nx3248, nx3258, 
      nx3268, nx3278, nx3288, nx3298, nx3308, nx3318, nx3348, nx3368, nx3398, 
      nx3421, nx3483, nx3487, nx3498, nx3500, nx3508, nx3521, nx3523, nx3534, 
      nx3540, nx3544, nx3550, nx3552, nx3566, nx3568, nx3574, nx3576, nx3582, 
      nx3591, nx3597, nx3601, nx3607, nx3609, nx3615, nx3624, nx3627, nx3629, 
      nx3635, nx3637, nx3643, nx3652, nx3655, nx3657, nx3663, nx3665, nx3680, 
      nx3683, nx3685, nx3691, nx3693, nx3708, nx3711, nx3713, nx3719, nx3721, 
      nx3736, nx3739, nx3741, nx3747, nx3749, nx3764, nx3767, nx3769, nx3775, 
      nx3777, nx3792, nx3795, nx3797, nx3803, nx3805, nx3820, nx3823, nx3825, 
      nx3831, nx3833, nx3848, nx3851, nx3853, nx3859, nx3861, nx3873, nx3876, 
      nx3879, nx3887, nx3889, nx3895, nx3901, nx3904, nx3912, nx3914, nx3920, 
      nx3924, nx3926, nx3928, nx3931, nx3933, nx3943, nx3945, nx3955, nx3964, 
      nx3966, nx3976, nx3985, nx3987, nx3993, nx3997, nx4006, nx4008, nx4014, 
      nx4018, nx4027, nx4029, nx4035, nx4039, nx4048, nx4050, nx4060, nx4069, 
      nx4081, nx4090, nx4098, nx4102, nx4111, nx4113, nx4123, nx4132, nx4144, 
      nx4153, nx4161, nx4165, nx4174, nx4182, nx4186, nx4195, nx4203, nx4207, 
      nx4216, nx4224, nx4237, nx4245, nx4262, nx4268, nx4270, nx4272, nx4280, 
      nx4284, nx4286, nx4288, nx4290, nx4292, nx4294, nx4296, nx4298, nx4308, 
      nx4310, nx4312, nx4314, nx4316, nx4318, nx4320, nx4332, nx4348, nx4350, 
      nx4352, nx4354, nx4376, nx4380, nx4382, nx4384, nx4396, nx4398, nx4400, 
      nx4402, nx4406, nx4410, nx4412, nx4414, nx4416, nx4418, nx4420, nx4436, 
      nx4438, nx4440, nx4442, nx4444, nx4446, nx4448, nx4450, nx4456, nx4458, 
      nx4460, nx4466, nx4468, nx4470, nx4476, nx4480, nx4482, nx4484, nx4486, 
      nx4488, nx4490, nx236, nx4322_XX0_XREP40, nx4274, shifting_R_2, nx3454, 
      nx3424, nx4274_XX0_XREP44, nx884, nx790, nx4322, nx4478_XX0_XREP64, 
      nx4580, nx4581, nx4582, nx4583, nx4584, nx4585, nx4586, nx4587, nx4588, 
      nx4589, nx4590, nx4591, nx4592, nx4593, nx4594, nx4218, nx4595, nx4596, 
      nx4597, nx4598, nx4599, nx4600, nx4601, nx4602, nx4603, nx4604, nx4454, 
      nx4605, nx4606, nx4607, nx4608, nx4609, nx4610, nx4611, nx4612, nx4613, 
      nx4614, nx4615, nx4616, nx4617, nx4618, nx4619, nx4620, nx4304, nx4621, 
      nx4622, nx4623, nx4624, nx4625, nx4626, nx4627, nx4628, nx4629, nx4630, 
      nx4631, nx4632, nx4633, nx4634, nx4635, nx4074, nx4636, nx4637, nx4638, 
      nx4639, nx4640, nx4641, nx4642, nx4643, nx4644, nx4645, nx4646, nx4647, 
      nx4648, nx4649, nx4650, nx4651, nx4652, nx4653, nx3526, nx3492, nx4654, 
      nx368, nx4655, nx4656, nx4657, nx4658, nx4158, nx4659, nx4032, nx4660, 
      nx4661, nx4137, nx4662, nx3358, nx4663, nx4664, nx458, nx3529, nx4665, 
      nx462, nx4472, nx4462, nx4666, nx4667, nx4668, nx4669, nx4670, nx4671, 
      nx4672, nx4673, nx4674, nx4675, nx4676, nx4677, nx3990, nx3969, nx4678, 
      nx4679, nx4680, nx4681, nx4682, nx4683, nx3917, nx4684, nx4685, nx4686, 
      nx4687, nx3555, nx4688, nx4689, nx4690, nx4691, nx4692, nx4693, nx4694, 
      nx4695, nx4696, nx4697, nx4698, nx4699, nx4700, nx4701, nx4702, nx4703, 
      nx4704, nx4705, nx4706, nx4707, nx4708, nx3892, nx4709, nx3864, nx4710, 
      nx4711, nx4712, nx4713, nx4714, nx3579, nx4715, nx4716, nx556, nx4717, 
      nx4718, nx4719, nx4720, nx4721, nx4722, nx3948, nx4723, nx4724, nx4725, 
      nx4726, nx4727, nx4728, nx4729, nx4730, nx4731, nx4732, nx4733, nx4734, 
      nx4735, nx4736, nx4737, nx4738, nx4739, nx4740, nx4741, nx3808, nx3780, 
      nx4742, nx4743, nx4744, nx3612, nx4745, nx4746, nx4747, nx3752, nx4748, 
      nx4749, nx4750, nx4751, nx3724, nx3696, nx3668, nx4752, nx492, nx4753, 
      nx4754, nx4755, nx4756, nx4757, nx4758, nx4759, nx4760, nx4761, nx4762, 
      nx4763, nx4764, nx4765, nx4766, nx4767, nx4768, nx4769, nx876, nx4770, 
      nx782, nx4771, nx4772, nx696, nx688, nx4773, nx594, nx4774, nx4775, 
      nx4776, nx4777, nx4276, nx4264, nx4778, nx4779, nx928, nx3671, nx4780, 
      nx4781, nx4782, nx4783, nx4784, nx4785, nx4786, nx4787, nx3951, nx4788, 
      nx4789, nx1790, nx4790, nx4791, nx4792, nx4793, nx4794, nx4795, nx1850, 
      nx4796, nx4797, nx4798, nx4799, nx4800, nx4801, nx4802, nx4803, nx4804, 
      nx4805, nx4806, nx4807, nx4808, nx1910, nx4809, nx4810, nx4811, nx4812, 
      nx4813, nx4814, nx4815, nx4816, nx4817, nx4818, nx4819, nx4820, nx4821, 
      nx4822, nx4823, nx4824, nx4825, nx744, nx4826, nx650, nx838, nx4827, 
      nx4828, nx4829, nx4830, nx4831, nx602, nx4832, nx4833, nx4834, nx4835, 
      nx4836, nx4837, nx4838, nx1166, nx4839, nx4840, nx4841, nx1158, nx4842, 
      nx4843, nx4844, nx4845, nx4846, nx1072, nx4847, nx1064, nx4848, nx978, 
      nx4849, nx970, nx4850, nx4851, nx4852, nx4853, nx4854, nx4855, nx4856, 
      nx4857, nx4858, nx4859, nx4861, nx4862, nx1542, nx4863, nx4864, nx4865, 
      nx4866, nx4867, nx1534, nx4868, nx4869, nx1448, nx4870, nx1432, nx4871, 
      nx4872, nx1440, nx4873, nx4874, nx4875, nx1354, nx1346, nx4876, nx1260, 
      nx1252, nx4877, nx4878, nx1846, nx3972, nx4282, nx4478, nx4879, nx4880, 
      nx4881, nx4882, nx4883, nx4884, nx2270, nx4885, nx4886, nx4887, nx4888, 
      nx4053, nx4889, nx4890, nx4891, nx4892, nx4893, nx4894, nx4895, nx4896, 
      nx4897, nx4898, nx4899, nx4900, nx4901, nx4902, nx4903, nx4904, nx4905, 
      nx4906, nx4907, nx4908, nx4909, nx4910, nx4911, nx4221, nx4912, nx4913, 
      nx4914, nx4915, nx4916, nx4917, nx4918, nx4919, nx4920, nx4921, nx4922, 
      nx4923, nx4924, nx4925, nx4926, nx4927, nx1970, nx4928, nx4929, nx4930, 
      nx2030, nx4931, nx4932, nx4933, nx4934, nx4935, nx4936, nx4937, nx4938, 
      nx4939, nx4940, nx4941, nx4942, nx4943, nx4944, nx4945, nx4946, nx4947, 
      nx4948, nx3836, nx2326, nx4140, nx4949, nx4950, nx1210, nx3755, nx4951, 
      nx4952, nx4953, nx4954, nx1214, nx4955, nx4956, nx4957, nx4958, nx4959, 
      nx4960, nx4961, nx4962, nx4963, nx4964, nx4965, nx4966, nx4967, nx4968, 
      nx4011, nx4969, nx4970, nx4971, nx4155, nx4972, nx4973, nx4974, nx4975, 
      nx1056, nx4976, nx868, nx4977, nx4978, nx4979, nx4980, nx4981, nx4982, 
      nx4983, nx4984, nx4985, nx4986, nx4987, nx4988, nx3378, nx2146, nx4077, 
      nx3408, nx4989, nx4266, nx4990, nx4991, nx1398, nx3811, nx4992, nx4993, 
      nx4994, nx4995, nx1402, nx4996, nx4997, nx4998, nx4999, nx4474, nx4464, 
      nx4278, nx5000, nx1116, nx5001, nx5002, nx5003, nx5004, nx5005, nx5006, 
      nx5007, nx3699, nx5008, nx1026, nx5009, nx5010, nx5011, nx5012, nx5013, 
      nx5014, nx5015, nx1120, nx5016, nx5017, nx5018, nx5019, nx5020, nx2150, 
      nx5021, nx5022, nx5023, nx5024, nx5025, nx5026, nx5027, nx5028, nx5029, 
      nx5030, nx5031, nx5032, nx5033, nx5034, nx5035, nx5036, nx5037, nx5038, 
      nx5039, nx5040, nx5041, nx5042, nx5043, nx1022, nx5044, nx5045, nx5046, 
      nx5047, nx5048, nx5049, nx5050, nx5051, nx5052, nx5053, nx4119, nx5054, 
      nx5055, nx5056, nx5057, nx5058, nx5059, nx5060, nx5061, nx5062, nx932, 
      nx5063, nx1586, nx3867, nx5064, nx5065, nx5066, nx5067, nx1492, nx3839, 
      nx5068, nx5069, nx5070, nx5071, nx5072, nx1590, nx5073, nx5074, nx1496, 
      nx5075, nx5076, nx5077, nx5078, nx1304, nx5079, nx3640, nx5080, nx5081, 
      nx5082, nx5083, nx5084, nx5085, nx5086, nx3388, nx5087, nx5088, nx5089, 
      nx5090, nx5091, nx5092, nx5093, nx5094, nx5095, nx3783, nx5096, nx5097, 
      nx5098, nx5099, nx5100, nx5101, nx5102, nx5103, nx5104, nx5105, nx5106, 
      nx5107, nx5108, nx5109, nx5110, nx5111, nx5112, nx5113, nx5114, nx5115, 
      nx5116, nx5117, nx5118, nx5119, nx5120, nx5121, nx5122, nx3328, nx5123, 
      nx5124, nx5125, nx5126, nx5127, nx5128, nx5129, nx5130, nx5131, nx5132, 
      nx5133, nx5134, nx5135, nx5136, nx5137, nx5138, nx5139, nx5140, nx5141, 
      nx5142, nx5143, nx5144, nx5145, nx5146, nx5147, nx5148, nx5149, nx5150, 
      nx5151, nx5152, nx2450, nx1786, nx5153, nx4116, nx5154, nx5155, nx5156, 
      nx5157, nx5158, nx5159, nx5160, nx4302, nx5161, nx5162, nx5163, nx3338, 
      nx4452, nx5164, nx5165, nx5166, nx5167, nx5168, nx5169, nx5170, nx5171, 
      nx5172, nx5173, nx5174, nx5175, nx5176, nx5177, nx2330, nx5178, nx5179, 
      nx5180, nx2086, nx4056, nx5181, nx5182, nx5183, nx1730, nx5184, nx5185, 
      nx5186, nx5187, nx5188, nx5189, nx5190, nx5191, nx5192, nx5193, nx5194, 
      nx5195, nx5196, nx5197, nx5198, nx5199, nx5200, nx5201, nx5202, nx5203, 
      nx5204, nx5205, nx5206, nx5207, nx5208, nx5209, nx5210, nx5211, nx5212, 
      nx5213, nx5214, nx5215, nx5216, nx5217, nx5218, nx5219, nx5220, nx5221, 
      nx5222, nx5223, nx5224, nx5225, nx5226, nx5227, nx5228, nx5229, nx5230, 
      nx5231, nx5232, nx5233, nx5234, nx5235, nx5236, nx5237, nx5238, nx5239, 
      nx5240, nx5241, nx5905, nx5907, nx5909, nx5911, nx5913, nx5915, nx5917, 
      nx5919, nx5921, nx5923, nx5925, nx5927, nx5929, nx5931, nx5933, nx5935, 
      nx5937, nx5939, nx5941, nx5943, nx5945, nx5947, nx5949, nx5951, nx5953, 
      nx5955, nx5957, nx5959, nx5961, nx5971, nx5973, nx5975, nx5977, nx5979, 
      nx5981, nx5983, nx5985, nx5987, nx5989, nx5991, nx5993, nx5995, nx5997, 
      nx5999, nx6001, nx6003, nx6005, nx6007, nx6009: std_logic ;

begin
   reg_product_0 : dff port map ( Q=>product(0), QB=>OPEN, D=>aux_product_0, 
      CLK=>clk);
   ix3099 : oai21 port map ( Y=>nx3098, A0=>nx3421, A1=>nx4288, B0=>nx3483);
   reg_aux_product_0 : dff port map ( Q=>aux_product_0, QB=>nx3421, D=>
      nx3098, CLK=>clk);
   ix255 : nand04 port map ( Y=>nx254, A0=>nx3424, A1=>nx4322, A2=>nx4440, 
      A3=>nx5208);
   reg_shifting_R_1 : dff port map ( Q=>shifting_R_1, QB=>OPEN, D=>nx216, 
      CLK=>clk);
   ix217 : mux21_ni port map ( Y=>nx216, A0=>R(0), A1=>shifting_R_3, S0=>
      nx4438);
   reg_shifting_R_3 : dff port map ( Q=>shifting_R_3, QB=>OPEN, D=>nx206, 
      CLK=>clk);
   ix207 : mux21_ni port map ( Y=>nx206, A0=>R(2), A1=>shifting_R_5, S0=>
      nx4436);
   reg_shifting_R_5 : dff port map ( Q=>shifting_R_5, QB=>OPEN, D=>nx196, 
      CLK=>clk);
   ix197 : mux21_ni port map ( Y=>nx196, A0=>R(4), A1=>shifting_R_7, S0=>
      nx4436);
   reg_shifting_R_7 : dff port map ( Q=>shifting_R_7, QB=>OPEN, D=>nx186, 
      CLK=>clk);
   ix187 : mux21_ni port map ( Y=>nx186, A0=>R(6), A1=>shifting_R_9, S0=>
      nx4436);
   reg_shifting_R_9 : dff port map ( Q=>shifting_R_9, QB=>OPEN, D=>nx176, 
      CLK=>clk);
   ix177 : mux21_ni port map ( Y=>nx176, A0=>R(8), A1=>shifting_R_11, S0=>
      nx4436);
   reg_shifting_R_11 : dff port map ( Q=>shifting_R_11, QB=>OPEN, D=>nx166, 
      CLK=>clk);
   ix167 : mux21_ni port map ( Y=>nx166, A0=>R(10), A1=>shifting_R_13, S0=>
      nx4436);
   reg_shifting_R_13 : dff port map ( Q=>shifting_R_13, QB=>OPEN, D=>nx156, 
      CLK=>clk);
   ix157 : mux21_ni port map ( Y=>nx156, A0=>R(12), A1=>shifting_R_15, S0=>
      nx4436);
   reg_shifting_R_15 : dff port map ( Q=>shifting_R_15, QB=>OPEN, D=>nx146, 
      CLK=>clk);
   ix147 : nor02ii port map ( Y=>nx146, A0=>nx4436, A1=>R(14));
   reg_shifting_R_0 : dff port map ( Q=>shifting_R_0, QB=>OPEN, D=>nx108, 
      CLK=>clk);
   ix101 : mux21_ni port map ( Y=>nx100, A0=>R(1), A1=>shifting_R_4, S0=>
      nx4440);
   reg_shifting_R_4 : dff port map ( Q=>shifting_R_4, QB=>OPEN, D=>nx90, CLK
      =>clk);
   ix91 : mux21_ni port map ( Y=>nx90, A0=>R(3), A1=>shifting_R_6, S0=>
      nx4440);
   reg_shifting_R_6 : dff port map ( Q=>shifting_R_6, QB=>OPEN, D=>nx80, CLK
      =>clk);
   ix81 : mux21_ni port map ( Y=>nx80, A0=>R(5), A1=>shifting_R_8, S0=>
      nx4438);
   reg_shifting_R_8 : dff port map ( Q=>shifting_R_8, QB=>OPEN, D=>nx70, CLK
      =>clk);
   ix71 : mux21_ni port map ( Y=>nx70, A0=>R(7), A1=>shifting_R_10, S0=>
      nx4438);
   reg_shifting_R_10 : dff port map ( Q=>shifting_R_10, QB=>OPEN, D=>nx60, 
      CLK=>clk);
   ix61 : mux21_ni port map ( Y=>nx60, A0=>R(9), A1=>shifting_R_12, S0=>
      nx4438);
   reg_shifting_R_12 : dff port map ( Q=>shifting_R_12, QB=>OPEN, D=>nx50, 
      CLK=>clk);
   ix51 : mux21_ni port map ( Y=>nx50, A0=>R(11), A1=>shifting_R_14, S0=>
      nx4438);
   reg_shifting_R_14 : dff port map ( Q=>shifting_R_14, QB=>OPEN, D=>nx40, 
      CLK=>clk);
   ix41 : mux21_ni port map ( Y=>nx40, A0=>R(13), A1=>shifting_R_16, S0=>
      nx4438);
   reg_shifting_R_16 : dff port map ( Q=>shifting_R_16, QB=>OPEN, D=>nx30, 
      CLK=>clk);
   ix31 : nor02ii port map ( Y=>nx30, A0=>nx4438, A1=>R(15));
   ix3484 : nand04 port map ( Y=>nx3483, A0=>nx270, A1=>nx4440, A2=>nx3492, 
      A3=>nx4288);
   ix271 : or02 port map ( Y=>nx270, A0=>nx268, A1=>aux_product_0);
   reg_positive_2M_1 : dff port map ( Q=>positive_2M_1, QB=>nx3487, D=>nx258, 
      CLK=>clk);
   reg_product_1 : dff port map ( Q=>product(1), QB=>OPEN, D=>aux_product_1, 
      CLK=>clk);
   ix3109 : oai21 port map ( Y=>nx3108, A0=>nx3498, A1=>nx4288, B0=>nx3500);
   reg_aux_product_1 : dff port map ( Q=>aux_product_1, QB=>nx3498, D=>
      nx3108, CLK=>clk);
   ix3501 : nand03 port map ( Y=>nx3500, A0=>nx4440, A1=>nx370, A2=>nx4288);
   ix371 : xnor2 port map ( Y=>nx370, A0=>nx3492, A1=>nx368);
   reg_positive_M_1 : dff port map ( Q=>positive_M_1, QB=>nx3508, D=>nx354, 
      CLK=>clk);
   ix355 : nor02ii port map ( Y=>nx354, A0=>nx4440, A1=>nx6003);
   reg_negative_M_1 : dff port map ( Q=>negative_M_1, QB=>OPEN, D=>nx310, 
      CLK=>clk);
   ix311 : nor02ii port map ( Y=>nx310, A0=>nx4440, A1=>nx306);
   ix307 : aoi21 port map ( Y=>nx306, A0=>nx6003, A1=>nx6007, B0=>nx296);
   ix297 : nor02_2x port map ( Y=>nx296, A0=>nx6007, A1=>nx6003);
   reg_product_2 : dff port map ( Q=>product(2), QB=>OPEN, D=>aux_product_2, 
      CLK=>clk);
   ix3119 : oai21 port map ( Y=>nx3118, A0=>nx3521, A1=>nx4288, B0=>nx3523);
   reg_aux_product_2 : dff port map ( Q=>aux_product_2, QB=>nx3521, D=>
      nx3118, CLK=>clk);
   ix3524 : nand03 port map ( Y=>nx3523, A0=>nx4442, A1=>nx464, A2=>nx4288);
   ix465 : xnor2 port map ( Y=>nx464, A0=>nx3526, A1=>nx462);
   reg_negative_M_2 : dff port map ( Q=>negative_M_2, QB=>OPEN, D=>nx442, 
      CLK=>clk);
   ix443 : mux21_ni port map ( Y=>nx442, A0=>nx406, A1=>positive_2M_1, S0=>
      nx4442);
   ix407 : aoi21 port map ( Y=>nx406, A0=>nx3534, A1=>nx5999, B0=>nx398);
   ix399 : nor03_2x port map ( Y=>nx398, A0=>nx5999, A1=>nx6007, A2=>nx6003
   );
   reg_positive_M_2 : dff port map ( Q=>positive_M_2, QB=>nx3544, D=>nx426, 
      CLK=>clk);
   ix427 : oai21 port map ( Y=>nx426, A0=>nx4484, A1=>nx3487, B0=>nx3540);
   ix3541 : oai21 port map ( Y=>nx3540, A0=>nx350, A1=>nx4482, B0=>nx5999);
   ix351 : nor02_2x port map ( Y=>nx350, A0=>M(15), A1=>nx4442);
   reg_product_3 : dff port map ( Q=>product(3), QB=>OPEN, D=>aux_product_3, 
      CLK=>clk);
   ix3129 : oai21 port map ( Y=>nx3128, A0=>nx3550, A1=>nx4288, B0=>nx3552);
   reg_aux_product_3 : dff port map ( Q=>aux_product_3, QB=>nx3550, D=>
      nx3128, CLK=>clk);
   ix3553 : nand03 port map ( Y=>nx3552, A0=>nx4442, A1=>nx558, A2=>nx4290);
   ix559 : xnor2 port map ( Y=>nx558, A0=>nx3555, A1=>nx556);
   reg_negative_M_3 : dff port map ( Q=>negative_M_3, QB=>OPEN, D=>nx536, 
      CLK=>clk);
   ix537 : mux21_ni port map ( Y=>nx536, A0=>nx500, A1=>negative_M_1, S0=>
      nx4442);
   ix501 : xnor2 port map ( Y=>nx500, A0=>nx5997, A1=>nx398);
   reg_positive_M_3 : dff port map ( Q=>positive_M_3, QB=>nx3568, D=>nx520, 
      CLK=>clk);
   ix521 : oai21 port map ( Y=>nx520, A0=>nx4484, A1=>nx3508, B0=>nx3566);
   ix3567 : oai21 port map ( Y=>nx3566, A0=>nx350, A1=>nx4482, B0=>nx5997);
   reg_product_4 : dff port map ( Q=>product(4), QB=>OPEN, D=>aux_product_4, 
      CLK=>clk);
   ix3139 : oai21 port map ( Y=>nx3138, A0=>nx3574, A1=>nx4290, B0=>nx3576);
   reg_aux_product_4 : dff port map ( Q=>aux_product_4, QB=>nx3574, D=>
      nx3138, CLK=>clk);
   ix3577 : nand03 port map ( Y=>nx3576, A0=>nx4442, A1=>nx652, A2=>nx4290);
   ix653 : xnor2 port map ( Y=>nx652, A0=>nx3579, A1=>nx650);
   ix3583 : aoi221 port map ( Y=>nx3582, A0=>negative_M_4, A1=>nx4264, B0=>
      positive_M_4, B1=>nx4276, C0=>nx646);
   reg_negative_M_4 : dff port map ( Q=>negative_M_4, QB=>OPEN, D=>nx630, 
      CLK=>clk);
   ix631 : mux21_ni port map ( Y=>nx630, A0=>nx594, A1=>negative_M_2, S0=>
      nx4442);
   reg_positive_M_4 : dff port map ( Q=>positive_M_4, QB=>nx3601, D=>nx614, 
      CLK=>clk);
   ix615 : oai322 port map ( Y=>nx614, A0=>nx3591, A1=>nx5210, A2=>nx4348, 
      B0=>nx3597, B1=>nx4352, C0=>nx4484, C1=>nx3544);
   ix3592 : nor02ii port map ( Y=>nx3591, A0=>nx508, A1=>nx594);
   ix509 : nor04 port map ( Y=>nx508, A0=>nx5997, A1=>nx5999, A2=>nx6007, A3
      =>nx6003);
   ix3598 : inv01 port map ( Y=>nx3597, A=>M(4));
   reg_product_5 : dff port map ( Q=>product(5), QB=>OPEN, D=>aux_product_5, 
      CLK=>clk);
   ix3149 : oai21 port map ( Y=>nx3148, A0=>nx3607, A1=>nx4290, B0=>nx3609);
   reg_aux_product_5 : dff port map ( Q=>aux_product_5, QB=>nx3607, D=>
      nx3148, CLK=>clk);
   ix3610 : nand03 port map ( Y=>nx3609, A0=>nx4444, A1=>nx746, A2=>nx4290);
   ix747 : xnor2 port map ( Y=>nx746, A0=>nx3612, A1=>nx744);
   ix3616 : aoi221 port map ( Y=>nx3615, A0=>negative_M_5, A1=>nx4264, B0=>
      positive_M_5, B1=>nx4276, C0=>nx740);
   reg_negative_M_5 : dff port map ( Q=>negative_M_5, QB=>OPEN, D=>nx724, 
      CLK=>clk);
   ix725 : mux21_ni port map ( Y=>nx724, A0=>nx688, A1=>negative_M_3, S0=>
      nx4444);
   reg_positive_M_5 : dff port map ( Q=>positive_M_5, QB=>nx3629, D=>nx708, 
      CLK=>clk);
   ix709 : oai322 port map ( Y=>nx708, A0=>nx3624, A1=>nx696, A2=>nx4348, B0
      =>nx3627, B1=>nx4352, C0=>nx4484, C1=>nx3568);
   ix3625 : nor02ii port map ( Y=>nx3624, A0=>nx5210, A1=>nx4773);
   ix3628 : inv01 port map ( Y=>nx3627, A=>M(5));
   reg_product_6 : dff port map ( Q=>product(6), QB=>OPEN, D=>aux_product_6, 
      CLK=>clk);
   ix3159 : oai21 port map ( Y=>nx3158, A0=>nx3635, A1=>nx4290, B0=>nx3637);
   reg_aux_product_6 : dff port map ( Q=>aux_product_6, QB=>nx3635, D=>
      nx3158, CLK=>clk);
   ix3638 : nand03 port map ( Y=>nx3637, A0=>nx4444, A1=>nx840, A2=>nx4290);
   ix841 : xnor2 port map ( Y=>nx840, A0=>nx3640, A1=>nx838);
   ix3644 : aoi221 port map ( Y=>nx3643, A0=>negative_M_6, A1=>nx4264, B0=>
      positive_M_6, B1=>nx4276, C0=>nx834);
   reg_negative_M_6 : dff port map ( Q=>negative_M_6, QB=>OPEN, D=>nx818, 
      CLK=>clk);
   ix819 : mux21_ni port map ( Y=>nx818, A0=>nx782, A1=>negative_M_4, S0=>
      nx4444);
   reg_positive_M_6 : dff port map ( Q=>positive_M_6, QB=>nx3657, D=>nx802, 
      CLK=>clk);
   ix803 : oai322 port map ( Y=>nx802, A0=>nx3652, A1=>nx790, A2=>nx4348, B0
      =>nx3655, B1=>nx4352, C0=>nx4484, C1=>nx3601);
   ix3653 : nor02ii port map ( Y=>nx3652, A0=>nx696, A1=>nx4771);
   ix3656 : inv01 port map ( Y=>nx3655, A=>M(6));
   reg_product_7 : dff port map ( Q=>product(7), QB=>OPEN, D=>aux_product_7, 
      CLK=>clk);
   ix3169 : oai21 port map ( Y=>nx3168, A0=>nx3663, A1=>nx4292, B0=>nx3665);
   reg_aux_product_7 : dff port map ( Q=>aux_product_7, QB=>nx3663, D=>
      nx3168, CLK=>clk);
   ix3666 : nand03 port map ( Y=>nx3665, A0=>nx4444, A1=>nx934, A2=>nx4292);
   ix935 : xnor2 port map ( Y=>nx934, A0=>nx3668, A1=>nx932);
   reg_negative_M_7 : dff port map ( Q=>negative_M_7, QB=>OPEN, D=>nx912, 
      CLK=>clk);
   ix913 : mux21_ni port map ( Y=>nx912, A0=>nx4580, A1=>negative_M_5, S0=>
      nx4444);
   reg_positive_M_7 : dff port map ( Q=>positive_M_7, QB=>nx3685, D=>nx896, 
      CLK=>clk);
   ix897 : oai322 port map ( Y=>nx896, A0=>nx3680, A1=>nx884, A2=>nx4348, B0
      =>nx3683, B1=>nx4352, C0=>nx4310, C1=>nx3629);
   ix3681 : nor02ii port map ( Y=>nx3680, A0=>nx790, A1=>nx4580);
   ix3684 : inv01 port map ( Y=>nx3683, A=>M(7));
   reg_product_8 : dff port map ( Q=>product(8), QB=>OPEN, D=>aux_product_8, 
      CLK=>clk);
   ix3179 : oai21 port map ( Y=>nx3178, A0=>nx3691, A1=>nx4292, B0=>nx3693);
   reg_aux_product_8 : dff port map ( Q=>aux_product_8, QB=>nx3691, D=>
      nx3178, CLK=>clk);
   ix3694 : nand03 port map ( Y=>nx3693, A0=>nx4444, A1=>nx1028, A2=>nx4292
   );
   ix1029 : xnor2 port map ( Y=>nx1028, A0=>nx5921, A1=>nx1026);
   reg_negative_M_8 : dff port map ( Q=>negative_M_8, QB=>OPEN, D=>nx1006, 
      CLK=>clk);
   ix1007 : mux21_ni port map ( Y=>nx1006, A0=>nx970, A1=>negative_M_6, S0=>
      nx4446);
   reg_positive_M_8 : dff port map ( Q=>positive_M_8, QB=>nx3713, D=>nx990, 
      CLK=>clk);
   ix991 : oai322 port map ( Y=>nx990, A0=>nx3708, A1=>nx978, A2=>nx4348, B0
      =>nx3711, B1=>nx4352, C0=>nx4310, C1=>nx3657);
   ix3709 : nor02ii port map ( Y=>nx3708, A0=>nx884, A1=>nx970);
   ix3712 : inv01 port map ( Y=>nx3711, A=>M(8));
   reg_product_9 : dff port map ( Q=>product(9), QB=>OPEN, D=>aux_product_9, 
      CLK=>clk);
   ix3189 : oai21 port map ( Y=>nx3188, A0=>nx3719, A1=>nx4292, B0=>nx3721);
   reg_aux_product_9 : dff port map ( Q=>aux_product_9, QB=>nx3719, D=>
      nx3188, CLK=>clk);
   ix3722 : nand03 port map ( Y=>nx3721, A0=>nx4446, A1=>nx1122, A2=>nx4292
   );
   ix1123 : xnor2 port map ( Y=>nx1122, A0=>nx3724, A1=>nx1120);
   reg_negative_M_9 : dff port map ( Q=>negative_M_9, QB=>OPEN, D=>nx1100, 
      CLK=>clk);
   ix1101 : mux21_ni port map ( Y=>nx1100, A0=>nx1064, A1=>negative_M_7, S0
      =>nx4446);
   reg_positive_M_9 : dff port map ( Q=>positive_M_9, QB=>nx3741, D=>nx1084, 
      CLK=>clk);
   ix1085 : oai322 port map ( Y=>nx1084, A0=>nx3736, A1=>nx1072, A2=>nx4348, 
      B0=>nx3739, B1=>nx4352, C0=>nx4310, C1=>nx3685);
   ix3737 : nor02ii port map ( Y=>nx3736, A0=>nx4849, A1=>nx1064);
   ix3740 : inv01 port map ( Y=>nx3739, A=>M(9));
   reg_product_10 : dff port map ( Q=>product(10), QB=>OPEN, D=>
      aux_product_10, CLK=>clk);
   ix3199 : oai21 port map ( Y=>nx3198, A0=>nx3747, A1=>nx4292, B0=>nx3749);
   reg_aux_product_10 : dff port map ( Q=>aux_product_10, QB=>nx3747, D=>
      nx3198, CLK=>clk);
   ix3750 : nand03 port map ( Y=>nx3749, A0=>nx4446, A1=>nx1216, A2=>nx4294
   );
   ix1217 : xnor2 port map ( Y=>nx1216, A0=>nx3752, A1=>nx1214);
   reg_negative_M_10 : dff port map ( Q=>negative_M_10, QB=>OPEN, D=>nx1194, 
      CLK=>clk);
   ix1195 : mux21_ni port map ( Y=>nx1194, A0=>nx1158, A1=>negative_M_8, S0
      =>nx4446);
   reg_positive_M_10 : dff port map ( Q=>positive_M_10, QB=>nx3769, D=>
      nx1178, CLK=>clk);
   ix1179 : oai322 port map ( Y=>nx1178, A0=>nx3764, A1=>nx1166, A2=>nx4348, 
      B0=>nx3767, B1=>nx4352, C0=>nx4310, C1=>nx3713);
   ix3765 : nor02ii port map ( Y=>nx3764, A0=>nx4847, A1=>nx4842);
   ix3768 : inv01 port map ( Y=>nx3767, A=>M(10));
   reg_product_11 : dff port map ( Q=>product(11), QB=>OPEN, D=>
      aux_product_11, CLK=>clk);
   ix3209 : oai21 port map ( Y=>nx3208, A0=>nx3775, A1=>nx4294, B0=>nx3777);
   reg_aux_product_11 : dff port map ( Q=>aux_product_11, QB=>nx3775, D=>
      nx3208, CLK=>clk);
   ix3778 : nand03 port map ( Y=>nx3777, A0=>nx4446, A1=>nx1310, A2=>nx4294
   );
   ix1311 : xnor2 port map ( Y=>nx1310, A0=>nx3780, A1=>nx5905);
   reg_negative_M_11 : dff port map ( Q=>negative_M_11, QB=>OPEN, D=>nx1288, 
      CLK=>clk);
   ix1289 : mux21_ni port map ( Y=>nx1288, A0=>nx1252, A1=>negative_M_9, S0
      =>nx4446);
   ix1151 : nor02ii port map ( Y=>nx1150, A0=>M(10), A1=>nx1056);
   reg_positive_M_11 : dff port map ( Q=>positive_M_11, QB=>nx3797, D=>
      nx1272, CLK=>clk);
   ix1273 : oai322 port map ( Y=>nx1272, A0=>nx3792, A1=>nx1260, A2=>nx4350, 
      B0=>nx3795, B1=>nx4354, C0=>nx4310, C1=>nx3741);
   ix3793 : nor02ii port map ( Y=>nx3792, A0=>nx4839, A1=>nx1252);
   ix3796 : inv01 port map ( Y=>nx3795, A=>M(11));
   reg_product_12 : dff port map ( Q=>product(12), QB=>OPEN, D=>
      aux_product_12, CLK=>clk);
   ix3219 : oai21 port map ( Y=>nx3218, A0=>nx3803, A1=>nx4294, B0=>nx3805);
   reg_aux_product_12 : dff port map ( Q=>aux_product_12, QB=>nx3803, D=>
      nx3218, CLK=>clk);
   ix3806 : nand03 port map ( Y=>nx3805, A0=>nx4448, A1=>nx1404, A2=>nx4294
   );
   ix1405 : xnor2 port map ( Y=>nx1404, A0=>nx3808, A1=>nx1402);
   reg_negative_M_12 : dff port map ( Q=>negative_M_12, QB=>OPEN, D=>nx1382, 
      CLK=>clk);
   ix1383 : mux21_ni port map ( Y=>nx1382, A0=>nx1346, A1=>negative_M_10, S0
      =>nx4448);
   reg_positive_M_12 : dff port map ( Q=>positive_M_12, QB=>nx3825, D=>
      nx1366, CLK=>clk);
   ix1367 : oai322 port map ( Y=>nx1366, A0=>nx3820, A1=>nx1354, A2=>nx4350, 
      B0=>nx3823, B1=>nx4354, C0=>nx4310, C1=>nx3769);
   ix3821 : nor02ii port map ( Y=>nx3820, A0=>nx1260, A1=>nx1346);
   ix3824 : inv01 port map ( Y=>nx3823, A=>M(12));
   reg_product_13 : dff port map ( Q=>product(13), QB=>OPEN, D=>
      aux_product_13, CLK=>clk);
   ix3229 : oai21 port map ( Y=>nx3228, A0=>nx3831, A1=>nx4294, B0=>nx3833);
   reg_aux_product_13 : dff port map ( Q=>aux_product_13, QB=>nx3831, D=>
      nx3228, CLK=>clk);
   ix3834 : nand03 port map ( Y=>nx3833, A0=>nx4448, A1=>nx1498, A2=>nx4294
   );
   ix1499 : xnor2 port map ( Y=>nx1498, A0=>nx3836, A1=>nx1496);
   reg_negative_M_13 : dff port map ( Q=>negative_M_13, QB=>OPEN, D=>nx1476, 
      CLK=>clk);
   ix1477 : mux21_ni port map ( Y=>nx1476, A0=>nx1440, A1=>negative_M_11, S0
      =>nx4448);
   reg_positive_M_13 : dff port map ( Q=>positive_M_13, QB=>nx3853, D=>
      nx1460, CLK=>clk);
   ix1461 : oai322 port map ( Y=>nx1460, A0=>nx3848, A1=>nx1448, A2=>nx4350, 
      B0=>nx3851, B1=>nx4354, C0=>nx4310, C1=>nx3797);
   ix3849 : nor02ii port map ( Y=>nx3848, A0=>nx1354, A1=>nx4873);
   ix3852 : inv01 port map ( Y=>nx3851, A=>M(13));
   reg_product_14 : dff port map ( Q=>product(14), QB=>OPEN, D=>
      aux_product_14, CLK=>clk);
   ix3239 : oai21 port map ( Y=>nx3238, A0=>nx3859, A1=>nx4296, B0=>nx3861);
   reg_aux_product_14 : dff port map ( Q=>aux_product_14, QB=>nx3859, D=>
      nx3238, CLK=>clk);
   ix3862 : nand03 port map ( Y=>nx3861, A0=>nx4448, A1=>nx1592, A2=>nx4296
   );
   ix1593 : xnor2 port map ( Y=>nx1592, A0=>nx3864, A1=>nx1590);
   reg_negative_M_14 : dff port map ( Q=>negative_M_14, QB=>nx3873, D=>
      nx1570, CLK=>clk);
   ix1571 : mux21_ni port map ( Y=>nx1570, A0=>nx1534, A1=>negative_M_12, S0
      =>nx4448);
   reg_positive_M_14 : dff port map ( Q=>positive_M_14, QB=>OPEN, D=>nx1554, 
      CLK=>clk);
   ix1555 : oai322 port map ( Y=>nx1554, A0=>nx3876, A1=>nx1542, A2=>nx4350, 
      B0=>nx3879, B1=>nx4354, C0=>nx4312, C1=>nx3825);
   ix3877 : nor02ii port map ( Y=>nx3876, A0=>nx1448, A1=>nx4868);
   ix3880 : inv01 port map ( Y=>nx3879, A=>M(14));
   reg_product_15 : dff port map ( Q=>product(15), QB=>OPEN, D=>
      aux_product_15, CLK=>clk);
   ix3249 : oai21 port map ( Y=>nx3248, A0=>nx3887, A1=>nx4296, B0=>nx3889);
   reg_aux_product_15 : dff port map ( Q=>aux_product_15, QB=>nx3887, D=>
      nx3248, CLK=>clk);
   ix3890 : nand03 port map ( Y=>nx3889, A0=>nx4448, A1=>nx1662, A2=>nx4296
   );
   ix1663 : xnor2 port map ( Y=>nx1662, A0=>nx3892, A1=>nx1660);
   ix3896 : aoi221 port map ( Y=>nx3895, A0=>negative_M_15, A1=>nx4268, B0=>
      positive_M_15, B1=>nx4280, C0=>nx1656);
   reg_negative_M_15 : dff port map ( Q=>negative_M_15, QB=>nx3901, D=>
      nx1640, CLK=>clk);
   ix1641 : mux21_ni port map ( Y=>nx1640, A0=>nx1616, A1=>negative_M_13, S0
      =>nx4450);
   ix1617 : xnor2 port map ( Y=>nx1616, A0=>M(15), A1=>nx1526);
   ix1527 : nor02ii port map ( Y=>nx1526, A0=>M(14), A1=>nx1432);
   reg_positive_M_15 : dff port map ( Q=>positive_M_15, QB=>OPEN, D=>nx1624, 
      CLK=>clk);
   ix1625 : oai22 port map ( Y=>nx1624, A0=>nx3904, A1=>nx4350, B0=>nx4312, 
      B1=>nx3853);
   ix3905 : xor2 port map ( Y=>nx3904, A0=>nx1616, A1=>nx1542);
   reg_product_16 : dff port map ( Q=>product(16), QB=>OPEN, D=>
      aux_product_16, CLK=>clk);
   ix3259 : oai21 port map ( Y=>nx3258, A0=>nx3912, A1=>nx4296, B0=>nx3914);
   reg_aux_product_16 : dff port map ( Q=>aux_product_16, QB=>nx3912, D=>
      nx3258, CLK=>clk);
   ix3915 : nand03 port map ( Y=>nx3914, A0=>nx4450, A1=>nx1732, A2=>nx4296
   );
   ix1733 : xnor2 port map ( Y=>nx1732, A0=>nx3917, A1=>nx1730);
   ix3921 : aoi221 port map ( Y=>nx3920, A0=>negative_M_16, A1=>nx4268, B0=>
      positive_M_16, B1=>nx4280, C0=>nx1726);
   reg_negative_M_16 : dff port map ( Q=>negative_M_16, QB=>nx3928, D=>
      nx1710, CLK=>clk);
   ix1711 : oai21 port map ( Y=>nx1710, A0=>nx4312, A1=>nx3873, B0=>nx4380);
   ix3925 : nand02 port map ( Y=>nx3924, A0=>nx3926, A1=>nx350);
   reg_positive_M_16 : dff port map ( Q=>positive_M_16, QB=>OPEN, D=>nx1694, 
      CLK=>clk);
   ix3932 : oai21 port map ( Y=>nx3931, A0=>nx3933, A1=>nx1616, B0=>nx4482);
   reg_product_17 : dff port map ( Q=>product(17), QB=>OPEN, D=>
      aux_product_17, CLK=>clk);
   ix3269 : oai21 port map ( Y=>nx3268, A0=>nx3943, A1=>nx4296, B0=>nx3945);
   reg_aux_product_17 : dff port map ( Q=>aux_product_17, QB=>nx3943, D=>
      nx3268, CLK=>clk);
   ix3946 : nand03 port map ( Y=>nx3945, A0=>nx4450, A1=>nx1792, A2=>nx4298
   );
   ix1793 : xnor2 port map ( Y=>nx1792, A0=>nx3948, A1=>nx1790);
   reg_negative_M_17 : dff port map ( Q=>negative_M_17, QB=>nx3955, D=>
      nx1770, CLK=>clk);
   ix1771 : oai21 port map ( Y=>nx1770, A0=>nx4312, A1=>nx3901, B0=>nx4380);
   reg_positive_M_17 : dff port map ( Q=>positive_M_17, QB=>OPEN, D=>nx1758, 
      CLK=>clk);
   reg_product_18 : dff port map ( Q=>product(18), QB=>OPEN, D=>
      aux_product_18, CLK=>clk);
   ix3279 : oai21 port map ( Y=>nx3278, A0=>nx3964, A1=>nx4298, B0=>nx3966);
   reg_aux_product_18 : dff port map ( Q=>aux_product_18, QB=>nx3964, D=>
      nx3278, CLK=>clk);
   ix3967 : nand03 port map ( Y=>nx3966, A0=>nx4450, A1=>nx1852, A2=>nx4298
   );
   ix1853 : xnor2 port map ( Y=>nx1852, A0=>nx3969, A1=>nx5220);
   reg_negative_M_18 : dff port map ( Q=>negative_M_18, QB=>nx3976, D=>
      nx1830, CLK=>clk);
   ix1831 : oai21 port map ( Y=>nx1830, A0=>nx4312, A1=>nx3928, B0=>nx4380);
   reg_positive_M_18 : dff port map ( Q=>positive_M_18, QB=>OPEN, D=>nx1818, 
      CLK=>clk);
   reg_product_19 : dff port map ( Q=>product(19), QB=>OPEN, D=>
      aux_product_19, CLK=>clk);
   ix3289 : oai21 port map ( Y=>nx3288, A0=>nx3985, A1=>nx4298, B0=>nx3987);
   reg_aux_product_19 : dff port map ( Q=>aux_product_19, QB=>nx3985, D=>
      nx3288, CLK=>clk);
   ix3988 : nand03 port map ( Y=>nx3987, A0=>nx4450, A1=>nx1912, A2=>nx4298
   );
   ix1913 : xnor2 port map ( Y=>nx1912, A0=>nx3990, A1=>nx1910);
   ix3994 : aoi221 port map ( Y=>nx3993, A0=>negative_M_19, A1=>nx4268, B0=>
      positive_M_19, B1=>nx4280, C0=>nx1906);
   reg_negative_M_19 : dff port map ( Q=>negative_M_19, QB=>nx3997, D=>
      nx1890, CLK=>clk);
   ix1891 : oai21 port map ( Y=>nx1890, A0=>nx4314, A1=>nx3955, B0=>nx4380);
   reg_positive_M_19 : dff port map ( Q=>positive_M_19, QB=>OPEN, D=>nx1878, 
      CLK=>clk);
   reg_product_20 : dff port map ( Q=>product(20), QB=>OPEN, D=>
      aux_product_20, CLK=>clk);
   ix3299 : oai21 port map ( Y=>nx3298, A0=>nx4006, A1=>nx4298, B0=>nx4008);
   reg_aux_product_20 : dff port map ( Q=>aux_product_20, QB=>nx4006, D=>
      nx3298, CLK=>clk);
   ix4009 : nand03 port map ( Y=>nx4008, A0=>nx4450, A1=>nx1972, A2=>nx4298
   );
   ix1973 : xnor2 port map ( Y=>nx1972, A0=>nx4011, A1=>nx1970);
   ix4015 : aoi221 port map ( Y=>nx4014, A0=>negative_M_20, A1=>nx4268, B0=>
      positive_M_20, B1=>nx4280, C0=>nx1966);
   reg_negative_M_20 : dff port map ( Q=>negative_M_20, QB=>nx4018, D=>
      nx1950, CLK=>clk);
   ix1951 : oai21 port map ( Y=>nx1950, A0=>nx4314, A1=>nx3976, B0=>nx4380);
   reg_positive_M_20 : dff port map ( Q=>positive_M_20, QB=>OPEN, D=>nx1938, 
      CLK=>clk);
   reg_product_21 : dff port map ( Q=>product(21), QB=>OPEN, D=>
      aux_product_21, CLK=>clk);
   ix3309 : oai21 port map ( Y=>nx3308, A0=>nx4027, A1=>nx5228, B0=>nx4029);
   reg_aux_product_21 : dff port map ( Q=>aux_product_21, QB=>nx4027, D=>
      nx3308, CLK=>clk);
   ix4030 : nand03 port map ( Y=>nx4029, A0=>nx4450, A1=>nx2032, A2=>nx5228
   );
   ix2033 : xnor2 port map ( Y=>nx2032, A0=>nx4032, A1=>nx2030);
   ix4036 : aoi221 port map ( Y=>nx4035, A0=>negative_M_21, A1=>nx4268, B0=>
      positive_M_21, B1=>nx4280, C0=>nx2026);
   reg_negative_M_21 : dff port map ( Q=>negative_M_21, QB=>nx4039, D=>
      nx2010, CLK=>clk);
   ix2011 : oai21 port map ( Y=>nx2010, A0=>nx4314, A1=>nx3997, B0=>nx4380);
   reg_positive_M_21 : dff port map ( Q=>positive_M_21, QB=>OPEN, D=>nx1998, 
      CLK=>clk);
   reg_product_22 : dff port map ( Q=>product(22), QB=>OPEN, D=>
      aux_product_22, CLK=>clk);
   ix3319 : oai21 port map ( Y=>nx3318, A0=>nx4048, A1=>nx5228, B0=>nx4050);
   reg_aux_product_22 : dff port map ( Q=>aux_product_22, QB=>nx4048, D=>
      nx3318, CLK=>clk);
   ix4051 : nand03 port map ( Y=>nx4050, A0=>nx4452, A1=>nx2092, A2=>nx5228
   );
   ix2093 : xnor2 port map ( Y=>nx2092, A0=>nx4053, A1=>nx5234);
   reg_negative_M_22 : dff port map ( Q=>negative_M_22, QB=>nx4060, D=>
      nx2070, CLK=>clk);
   ix2071 : oai21 port map ( Y=>nx2070, A0=>nx4316, A1=>nx4018, B0=>nx4380);
   reg_positive_M_22 : dff port map ( Q=>positive_M_22, QB=>OPEN, D=>nx2058, 
      CLK=>clk);
   reg_product_23 : dff port map ( Q=>product(23), QB=>OPEN, D=>
      aux_product_23, CLK=>clk);
   reg_aux_product_23 : dff port map ( Q=>aux_product_23, QB=>nx4069, D=>
      nx3328, CLK=>clk);
   reg_negative_M_23 : dff port map ( Q=>negative_M_23, QB=>nx4081, D=>
      nx2130, CLK=>clk);
   ix2131 : oai21 port map ( Y=>nx2130, A0=>nx4316, A1=>nx4039, B0=>nx4382);
   reg_positive_M_23 : dff port map ( Q=>positive_M_23, QB=>OPEN, D=>nx2118, 
      CLK=>clk);
   reg_product_24 : dff port map ( Q=>product(24), QB=>OPEN, D=>
      aux_product_24, CLK=>clk);
   reg_aux_product_24 : dff port map ( Q=>aux_product_24, QB=>nx4090, D=>
      nx3338, CLK=>clk);
   ix4099 : aoi221 port map ( Y=>nx4098, A0=>negative_M_24, A1=>nx4270, B0=>
      positive_M_24, B1=>nx4282, C0=>nx2206);
   reg_negative_M_24 : dff port map ( Q=>negative_M_24, QB=>nx4102, D=>
      nx2190, CLK=>clk);
   ix2191 : oai21 port map ( Y=>nx2190, A0=>nx4316, A1=>nx4060, B0=>nx4382);
   reg_positive_M_24 : dff port map ( Q=>positive_M_24, QB=>OPEN, D=>nx2178, 
      CLK=>clk);
   reg_product_25 : dff port map ( Q=>product(25), QB=>OPEN, D=>
      aux_product_25, CLK=>clk);
   ix3349 : oai21 port map ( Y=>nx3348, A0=>nx4111, A1=>nx5228, B0=>nx4113);
   reg_aux_product_25 : dff port map ( Q=>aux_product_25, QB=>nx4111, D=>
      nx3348, CLK=>clk);
   ix4114 : nand03 port map ( Y=>nx4113, A0=>nx4452, A1=>nx2272, A2=>nx5228
   );
   ix2273 : xnor2 port map ( Y=>nx2272, A0=>nx4116, A1=>nx2270);
   reg_negative_M_25 : dff port map ( Q=>negative_M_25, QB=>nx4123, D=>
      nx2250, CLK=>clk);
   ix2251 : oai21 port map ( Y=>nx2250, A0=>nx4316, A1=>nx4081, B0=>nx4382);
   reg_positive_M_25 : dff port map ( Q=>positive_M_25, QB=>OPEN, D=>nx2238, 
      CLK=>clk);
   reg_product_26 : dff port map ( Q=>product(26), QB=>OPEN, D=>
      aux_product_26, CLK=>clk);
   reg_aux_product_26 : dff port map ( Q=>aux_product_26, QB=>nx4132, D=>
      nx3358, CLK=>clk);
   reg_negative_M_26 : dff port map ( Q=>negative_M_26, QB=>nx4144, D=>
      nx2310, CLK=>clk);
   ix2311 : oai21 port map ( Y=>nx2310, A0=>nx4318, A1=>nx4102, B0=>nx4382);
   reg_positive_M_26 : dff port map ( Q=>positive_M_26, QB=>OPEN, D=>nx2298, 
      CLK=>clk);
   reg_product_27 : dff port map ( Q=>product(27), QB=>OPEN, D=>
      aux_product_27, CLK=>clk);
   ix3369 : oai21 port map ( Y=>nx3368, A0=>nx4153, A1=>nx5228, B0=>nx4155);
   reg_aux_product_27 : dff port map ( Q=>aux_product_27, QB=>nx4153, D=>
      nx3368, CLK=>clk);
   ix4162 : aoi221 port map ( Y=>nx4161, A0=>negative_M_27, A1=>nx4270, B0=>
      positive_M_27, B1=>nx4282, C0=>nx2386);
   reg_negative_M_27 : dff port map ( Q=>negative_M_27, QB=>nx4165, D=>
      nx2370, CLK=>clk);
   ix2371 : oai21 port map ( Y=>nx2370, A0=>nx4318, A1=>nx4123, B0=>nx4382);
   reg_positive_M_27 : dff port map ( Q=>positive_M_27, QB=>OPEN, D=>nx2358, 
      CLK=>clk);
   reg_product_28 : dff port map ( Q=>product(28), QB=>OPEN, D=>
      aux_product_28, CLK=>clk);
   reg_aux_product_28 : dff port map ( Q=>aux_product_28, QB=>nx4174, D=>
      nx3378, CLK=>clk);
   ix4183 : aoi221 port map ( Y=>nx4182, A0=>negative_M_28, A1=>nx4270, B0=>
      positive_M_28, B1=>nx4282, C0=>nx2446);
   reg_negative_M_28 : dff port map ( Q=>negative_M_28, QB=>nx4186, D=>
      nx2430, CLK=>clk);
   ix2431 : oai21 port map ( Y=>nx2430, A0=>nx4318, A1=>nx4144, B0=>nx4382);
   reg_positive_M_28 : dff port map ( Q=>positive_M_28, QB=>OPEN, D=>nx2418, 
      CLK=>clk);
   reg_product_29 : dff port map ( Q=>product(29), QB=>OPEN, D=>
      aux_product_29, CLK=>clk);
   reg_aux_product_29 : dff port map ( Q=>aux_product_29, QB=>nx4195, D=>
      nx3388, CLK=>clk);
   ix4204 : aoi221 port map ( Y=>nx4203, A0=>negative_M_29, A1=>nx4272, B0=>
      positive_M_29, B1=>nx4284, C0=>nx2506);
   reg_negative_M_29 : dff port map ( Q=>negative_M_29, QB=>nx4207, D=>
      nx2490, CLK=>clk);
   ix2491 : oai21 port map ( Y=>nx2490, A0=>nx4320, A1=>nx4165, B0=>nx4382);
   reg_positive_M_29 : dff port map ( Q=>positive_M_29, QB=>OPEN, D=>nx2478, 
      CLK=>clk);
   reg_product_30 : dff port map ( Q=>product(30), QB=>OPEN, D=>
      aux_product_30, CLK=>clk);
   ix3399 : oai21 port map ( Y=>nx3398, A0=>nx4216, A1=>nx4304, B0=>nx4218);
   reg_aux_product_30 : dff port map ( Q=>aux_product_30, QB=>nx4216, D=>
      nx3398, CLK=>clk);
   ix4225 : aoi221 port map ( Y=>nx4224, A0=>negative_2M_31, A1=>nx4272, B0
      =>positive_2M_31, B1=>nx4284, C0=>nx2566);
   reg_negative_2M_31 : dff port map ( Q=>negative_2M_31, QB=>OPEN, D=>
      nx2550, CLK=>clk);
   ix2551 : oai21 port map ( Y=>nx2550, A0=>nx4320, A1=>nx4186, B0=>nx3924);
   reg_positive_2M_31 : dff port map ( Q=>positive_2M_31, QB=>OPEN, D=>
      nx2538, CLK=>clk);
   reg_product_31 : dff port map ( Q=>product(31), QB=>OPEN, D=>
      aux_product_31, CLK=>clk);
   reg_aux_product_31 : dff port map ( Q=>aux_product_31, QB=>nx4237, D=>
      nx3408, CLK=>clk);
   ix4246 : aoi221 port map ( Y=>nx4245, A0=>negative_M_31, A1=>nx4272, B0=>
      positive_M_31, B1=>nx4284, C0=>nx2626);
   reg_negative_M_31 : dff port map ( Q=>negative_M_31, QB=>OPEN, D=>nx2610, 
      CLK=>clk);
   ix2611 : oai21 port map ( Y=>nx2610, A0=>nx4320, A1=>nx4207, B0=>nx3924);
   reg_positive_M_31 : dff port map ( Q=>positive_M_31, QB=>OPEN, D=>nx2598, 
      CLK=>clk);
   ix2627 : ao22 port map ( Y=>nx2626, A0=>negative_2M_31, A1=>nx4472, B0=>
      positive_2M_31, B1=>nx4462);
   ix3934 : inv01 port map ( Y=>nx3933, A=>nx1542);
   ix3927 : inv01 port map ( Y=>nx3926, A=>nx1526);
   ix3535 : inv01 port map ( Y=>nx3534, A=>nx296);
   ix4267 : inv02 port map ( Y=>nx4268, A=>nx4262);
   ix4269 : inv02 port map ( Y=>nx4270, A=>nx4262);
   ix4271 : inv02 port map ( Y=>nx4272, A=>nx4262);
   ix4279 : inv02 port map ( Y=>nx4280, A=>nx4274);
   ix4283 : inv02 port map ( Y=>nx4284, A=>nx4274);
   ix4285 : inv01 port map ( Y=>nx4286, A=>nx254);
   ix4287 : inv02 port map ( Y=>nx4288, A=>nx4420);
   ix4289 : inv02 port map ( Y=>nx4290, A=>nx4420);
   ix4291 : inv02 port map ( Y=>nx4292, A=>nx4420);
   ix4293 : inv02 port map ( Y=>nx4294, A=>nx4420);
   ix4295 : inv02 port map ( Y=>nx4296, A=>nx4420);
   ix4297 : inv02 port map ( Y=>nx4298, A=>nx5226);
   ix4307 : inv02 port map ( Y=>nx4308, A=>cnt_enable);
   ix4309 : inv02 port map ( Y=>nx4310, A=>nx4454);
   ix4311 : inv02 port map ( Y=>nx4312, A=>nx4454);
   ix4313 : inv02 port map ( Y=>nx4314, A=>nx4454);
   ix4315 : inv02 port map ( Y=>nx4316, A=>nx4454);
   ix4317 : inv02 port map ( Y=>nx4318, A=>nx4456);
   ix4319 : inv02 port map ( Y=>nx4320, A=>nx4456);
   ix4331 : inv02 port map ( Y=>nx4332, A=>nx228);
   ix4347 : inv04 port map ( Y=>nx4348, A=>nx338);
   ix4349 : inv04 port map ( Y=>nx4350, A=>nx4482);
   ix4351 : inv02 port map ( Y=>nx4352, A=>nx350);
   ix4353 : inv02 port map ( Y=>nx4354, A=>nx350);
   ix4375 : buf02 port map ( Y=>nx4376, A=>nx3895);
   ix4379 : nand02 port map ( Y=>nx4380, A0=>nx3926, A1=>nx350);
   ix4381 : nand02 port map ( Y=>nx4382, A0=>nx3926, A1=>nx350);
   ix4383 : inv01 port map ( Y=>nx4384, A=>nx3931);
   ix4395 : buf02 port map ( Y=>nx4396, A=>nx3993);
   ix4397 : buf02 port map ( Y=>nx4398, A=>nx4014);
   ix4399 : buf02 port map ( Y=>nx4400, A=>nx4035);
   ix4401 : buf02 port map ( Y=>nx4402, A=>nx4056);
   ix4405 : buf02 port map ( Y=>nx4406, A=>nx4098);
   ix4409 : buf02 port map ( Y=>nx4410, A=>nx4140);
   ix4411 : buf02 port map ( Y=>nx4412, A=>nx4161);
   ix4413 : buf02 port map ( Y=>nx4414, A=>nx4182);
   ix4415 : buf02 port map ( Y=>nx4416, A=>nx4203);
   ix4417 : buf02 port map ( Y=>nx4418, A=>nx4224);
   ix4419 : inv01 port map ( Y=>nx4420, A=>nx254);
   ix109 : and02 port map ( Y=>nx108, A0=>nx4456, A1=>shifting_R_2);
   ix3482 : and03 port map ( Y=>nx228, A0=>shifting_R_0, A1=>nx3454, A2=>
      shifting_R_1);
   ix269 : nor02ii port map ( Y=>nx268, A0=>nx3424, A1=>positive_2M_1);
   ix259 : nor02ii port map ( Y=>nx258, A0=>nx4456, A1=>nx6007);
   ix247 : or02 port map ( Y=>nx4262, A0=>nx3454, A1=>nx3424);
   ix553 : ao22 port map ( Y=>nx552, A0=>negative_M_2, A1=>nx4472, B0=>
      positive_M_2, B1=>nx4462);
   ix3596 : nor02ii port map ( Y=>nx338, A0=>nx4456, A1=>M(15));
   ix647 : ao22 port map ( Y=>nx646, A0=>negative_M_3, A1=>nx4472, B0=>
      positive_M_3, B1=>nx4462);
   ix741 : ao22 port map ( Y=>nx740, A0=>negative_M_4, A1=>nx4472, B0=>
      positive_M_4, B1=>nx4462);
   ix835 : ao22 port map ( Y=>nx834, A0=>negative_M_5, A1=>nx4472, B0=>
      positive_M_5, B1=>nx4462);
   ix1309 : xor2 port map ( Y=>nx1308, A0=>nx3775, A1=>nx5953);
   ix1661 : xor2 port map ( Y=>nx1660, A0=>nx3887, A1=>nx4376);
   ix1657 : ao22 port map ( Y=>nx1656, A0=>negative_M_14, A1=>nx4476, B0=>
      positive_M_14, B1=>nx4466);
   ix1695 : ao21 port map ( Y=>nx1694, A0=>nx4456, A1=>positive_M_14, B0=>
      nx4488);
   ix1727 : ao22 port map ( Y=>nx1726, A0=>negative_M_15, A1=>nx4476, B0=>
      positive_M_15, B1=>nx4466);
   ix1759 : ao21 port map ( Y=>nx1758, A0=>nx4456, A1=>positive_M_15, B0=>
      nx4488);
   ix1819 : ao21 port map ( Y=>nx1818, A0=>nx4458, A1=>positive_M_16, B0=>
      nx4488);
   ix1879 : ao21 port map ( Y=>nx1878, A0=>nx4458, A1=>positive_M_17, B0=>
      nx4488);
   ix1907 : ao22 port map ( Y=>nx1906, A0=>negative_M_18, A1=>nx4476, B0=>
      positive_M_18, B1=>nx4466);
   ix1939 : ao21 port map ( Y=>nx1938, A0=>nx4458, A1=>positive_M_18, B0=>
      nx4488);
   ix1967 : ao22 port map ( Y=>nx1966, A0=>negative_M_19, A1=>nx4476, B0=>
      positive_M_19, B1=>nx4466);
   ix1999 : ao21 port map ( Y=>nx1998, A0=>nx4458, A1=>positive_M_19, B0=>
      nx4488);
   ix2027 : ao22 port map ( Y=>nx2026, A0=>negative_M_20, A1=>
      nx4478_XX0_XREP64, B0=>positive_M_20, B1=>nx4468);
   ix2091 : xor2 port map ( Y=>nx2090, A0=>nx4048, A1=>nx4402);
   ix2059 : ao21 port map ( Y=>nx2058, A0=>nx4458, A1=>positive_M_20, B0=>
      nx4488);
   ix2119 : ao21 port map ( Y=>nx2118, A0=>nx4458, A1=>positive_M_21, B0=>
      nx4490);
   ix2211 : xor2_2x port map ( Y=>nx2210, A0=>nx4090, A1=>nx4406);
   ix2179 : ao21 port map ( Y=>nx2178, A0=>nx4458, A1=>positive_M_22, B0=>
      nx4490);
   ix2207 : ao22 port map ( Y=>nx2206, A0=>negative_M_23, A1=>nx4478, B0=>
      positive_M_23, B1=>nx4468);
   ix2239 : ao21 port map ( Y=>nx2238, A0=>nx4460, A1=>positive_M_23, B0=>
      nx4490);
   ix2299 : ao21 port map ( Y=>nx2298, A0=>nx4460, A1=>positive_M_24, B0=>
      nx4490);
   ix2391 : xor2 port map ( Y=>nx2390, A0=>nx4153, A1=>nx4412);
   ix2359 : ao21 port map ( Y=>nx2358, A0=>nx4460, A1=>positive_M_25, B0=>
      nx4490);
   ix2387 : ao22 port map ( Y=>nx2386, A0=>negative_M_26, A1=>nx4478, B0=>
      positive_M_26, B1=>nx4468);
   ix2419 : ao21 port map ( Y=>nx2418, A0=>nx4460, A1=>positive_M_26, B0=>
      nx4490);
   ix2447 : ao22 port map ( Y=>nx2446, A0=>negative_M_27, A1=>nx4480, B0=>
      positive_M_27, B1=>nx4470);
   ix2511 : xor2 port map ( Y=>nx2510, A0=>nx4195, A1=>nx4416);
   ix2479 : ao21 port map ( Y=>nx2478, A0=>nx4460, A1=>positive_M_27, B0=>
      nx4490);
   ix2507 : ao22 port map ( Y=>nx2506, A0=>negative_M_28, A1=>nx4480, B0=>
      positive_M_28, B1=>nx4470);
   ix2571 : xor2 port map ( Y=>nx2570, A0=>nx4216, A1=>nx4418);
   ix2539 : ao21 port map ( Y=>nx2538, A0=>nx4460, A1=>positive_M_28, B0=>
      nx4384);
   ix2567 : ao22 port map ( Y=>nx2566, A0=>negative_M_29, A1=>nx4480, B0=>
      positive_M_29, B1=>nx4470);
   ix2631 : xor2 port map ( Y=>nx2630, A0=>nx4237, A1=>nx4245);
   ix2599 : ao21 port map ( Y=>nx2598, A0=>nx4460, A1=>positive_M_29, B0=>
      nx4384);
   ix4435 : inv02 port map ( Y=>nx4436, A=>nx4484);
   ix4437 : inv02 port map ( Y=>nx4438, A=>nx4484);
   ix4439 : inv02 port map ( Y=>nx4440, A=>nx5232);
   ix4441 : inv02 port map ( Y=>nx4442, A=>nx5232);
   ix4443 : inv02 port map ( Y=>nx4444, A=>nx5232);
   ix4445 : inv02 port map ( Y=>nx4446, A=>nx5232);
   ix4447 : inv02 port map ( Y=>nx4448, A=>nx5232);
   ix4449 : inv02 port map ( Y=>nx4450, A=>nx5233);
   ix4455 : inv02 port map ( Y=>nx4456, A=>nx4308);
   ix4457 : inv02 port map ( Y=>nx4458, A=>nx4308);
   ix4459 : inv02 port map ( Y=>nx4460, A=>nx4308);
   ix4465 : inv02 port map ( Y=>nx4466, A=>nx5208);
   ix4467 : inv02 port map ( Y=>nx4468, A=>nx5208);
   ix4469 : inv02 port map ( Y=>nx4470, A=>nx5208);
   ix4475 : inv02 port map ( Y=>nx4476, A=>nx4322_XX0_XREP40);
   ix4479 : inv02 port map ( Y=>nx4480, A=>nx4322);
   ix4481 : inv02 port map ( Y=>nx4482, A=>nx4348);
   ix4483 : inv02 port map ( Y=>nx4484, A=>cnt_enable);
   ix4485 : inv02 port map ( Y=>nx4486, A=>cnt_enable);
   ix4487 : inv01 port map ( Y=>nx4488, A=>nx3931);
   ix4489 : inv01 port map ( Y=>nx4490, A=>nx3931);
   ix237 : nor03_2x port map ( Y=>nx236, A0=>shifting_R_0, A1=>nx3454, A2=>
      shifting_R_1);
   ix4321_0_XREP40 : inv02 port map ( Y=>nx4322_XX0_XREP40, A=>nx236);
   ix251 : or02 port map ( Y=>nx4274, A0=>shifting_R_2, A1=>nx3424);
   reg_shifting_R_2 : dff port map ( Q=>shifting_R_2, QB=>nx3454, D=>nx100, 
      CLK=>clk);
   ix3425 : xnor2 port map ( Y=>nx3424, A0=>shifting_R_1, A1=>shifting_R_0);
   ix251_0_XREP44 : or02 port map ( Y=>nx4274_XX0_XREP44, A0=>shifting_R_2, 
      A1=>nx3424);
   ix885 : nor02ii port map ( Y=>nx884, A0=>nx4580, A1=>nx790);
   ix791 : nor02ii port map ( Y=>nx790, A0=>nx4772, A1=>nx696);
   ix4321 : inv02 port map ( Y=>nx4322, A=>nx236);
   ix4477_0_XREP64 : inv02 port map ( Y=>nx4478_XX0_XREP64, A=>nx4322);
   ix5242 : buf04 port map ( Y=>nx4580, A=>nx876);
   ix5243 : inv01 port map ( Y=>nx4581, A=>nx2510);
   ix5244 : inv02 port map ( Y=>nx4582, A=>nx2570);
   ix5245 : nor04_2x port map ( Y=>nx4583, A0=>nx4582, A1=>nx2630, A2=>
      nx5226, A3=>nx4308);
   ix5246 : inv02 port map ( Y=>nx4584, A=>nx2630);
   ix5247 : inv01 port map ( Y=>nx4585, A=>nx4418);
   ix5248 : aoi22 port map ( Y=>nx4586, A0=>nx2630, A1=>nx4418, B0=>nx4584, 
      B1=>nx4585);
   ix5249 : nor02_2x port map ( Y=>nx4587, A0=>nx5226, A1=>nx4308);
   ix5250 : nand03_2x port map ( Y=>nx4588, A0=>nx4587, A1=>nx2630, A2=>
      nx2570);
   ix5251 : inv02 port map ( Y=>nx4589, A=>nx2570);
   ix5252 : and02 port map ( Y=>nx4590, A0=>nx4416, A1=>nx4581);
   ix5253 : inv01 port map ( Y=>nx4591, A=>nx4414);
   ix5254 : nand02_2x port map ( Y=>nx4592, A0=>nx5152, A1=>nx4591);
   ix5255 : aoi22 port map ( Y=>nx4593, A0=>nx4416, A1=>nx4581, B0=>nx2510, 
      B1=>nx4592);
   ix5256 : nand02_2x port map ( Y=>nx4594, A0=>nx4589, A1=>nx4221);
   reg_nx4218 : nand04_2x port map ( Y=>nx4218, A0=>nx4594, A1=>nx4614, A2=>
      nx4454, A3=>nx4304);
   ix5257 : inv01 port map ( Y=>nx4595, A=>nx5240);
   ix5258 : nor03_2x port map ( Y=>nx4596, A0=>nx4595, A1=>nx4588, A2=>
      nx4593);
   ix5259 : nor02ii port map ( Y=>nx4597, A0=>nx5240, A1=>nx4412);
   ix5260 : nor03_2x port map ( Y=>nx4598, A0=>nx4597, A1=>nx5152, A2=>
      nx4590);
   ix5261 : inv01 port map ( Y=>nx4599, A=>nx5226);
   ix5262 : inv02 port map ( Y=>nx4600, A=>nx4308);
   ix5263 : nand02_2x port map ( Y=>nx4601, A0=>nx4599, A1=>nx4600);
   ix5264 : oai332 port map ( Y=>nx4602, A0=>nx4598, A1=>nx4588, A2=>nx4593, 
      B0=>nx4586, B1=>nx2570, B2=>nx4601, C0=>nx4304, C1=>nx4237);
   ix5265 : inv01 port map ( Y=>nx4603, A=>nx4593);
   ix5266 : inv01 port map ( Y=>nx4604, A=>nx4598);
   reg_nx4454 : inv02 port map ( Y=>nx4454, A=>nx4308);
   ix5267 : nand03_2x port map ( Y=>nx4605, A0=>nx2510, A1=>nx4304, A2=>
      nx4454);
   ix5268 : inv02 port map ( Y=>nx4606, A=>nx2510);
   ix5269 : nor02_2x port map ( Y=>nx4607, A0=>nx5226, A1=>nx4308);
   ix5270 : and02 port map ( Y=>nx4608, A0=>nx5240, A1=>nx4603);
   ix5271 : nand04_2x port map ( Y=>nx4609, A0=>nx4116, A1=>nx4608, A2=>
      nx2330, A3=>nx4885);
   ix5272 : inv01 port map ( Y=>nx4610, A=>nx5236);
   ix5273 : inv01 port map ( Y=>nx4611, A=>nx5238);
   ix5274 : oai32 port map ( Y=>nx4612, A0=>nx4886, A1=>nx5959, A2=>nx4610, 
      B0=>nx4611, B1=>nx5178);
   ix5275 : aoi321 port map ( Y=>nx4613, A0=>nx4612, A1=>nx5240, A2=>nx4603, 
      B0=>nx4603, B1=>nx4604, C0=>nx4589);
   ix5276 : nand02_2x port map ( Y=>nx4614, A0=>nx4609, A1=>nx4613);
   ix5277 : inv01 port map ( Y=>nx4615, A=>nx4604);
   ix5278 : oai321 port map ( Y=>nx4616, A0=>nx5959, A1=>nx4887, A2=>nx5236, 
      B0=>nx5179, B1=>nx5238, C0=>nx5240);
   ix5279 : inv01 port map ( Y=>nx4617, A=>nx4603);
   ix5280 : inv01 port map ( Y=>nx4618, A=>nx2450);
   ix5281 : inv01 port map ( Y=>nx4619, A=>nx4412);
   ix5282 : inv01 port map ( Y=>nx4620, A=>nx4595);
   reg_nx4304 : inv02 port map ( Y=>nx4304, A=>nx5227);
   ix5283 : nand03_2x port map ( Y=>nx4621, A0=>nx4618, A1=>nx4304, A2=>
      nx4452);
   ix5284 : inv01 port map ( Y=>nx4622, A=>nx5236);
   ix5285 : inv01 port map ( Y=>nx4623, A=>nx5238);
   ix5286 : inv01 port map ( Y=>nx4624, A=>nx5234);
   ix5287 : nor02ii port map ( Y=>nx4625, A0=>nx5022, A1=>nx5941);
   ix5288 : inv01 port map ( Y=>nx4626, A=>nx2210);
   ix5289 : aoi422 port map ( Y=>nx4627, A0=>nx2210, A1=>nx4624, A2=>nx5023, 
      A3=>nx4402, B0=>nx2210, B1=>nx4625, C0=>nx4406, C1=>nx4626);
   ix5290 : oai322 port map ( Y=>nx4628, A0=>nx5129, A1=>nx5143, A2=>nx4622, 
      B0=>nx4623, B1=>nx5139, C0=>nx5174, C1=>nx4627);
   ix5291 : inv01 port map ( Y=>nx4629, A=>nx4402);
   ix5292 : inv01 port map ( Y=>nx4630, A=>nx4077);
   ix5293 : oai32 port map ( Y=>nx4631, A0=>nx5029, A1=>nx4629, A2=>nx5234, 
      B0=>nx4630, B1=>nx5024);
   ix5294 : nor02_2x port map ( Y=>nx4632, A0=>nx5959, A1=>nx5236);
   ix5295 : nor02_2x port map ( Y=>nx4633, A0=>nx5959, A1=>nx5052);
   ix5296 : nor02_2x port map ( Y=>nx4634, A0=>nx4629, A1=>nx5234);
   ix5297 : aoi22 port map ( Y=>nx4635, A0=>nx5941, A1=>nx5029, B0=>nx5026, 
      B1=>nx4634);
   reg_nx4074 : ao22 port map ( Y=>nx4074, A0=>nx4402, A1=>nx4624, B0=>
      nx4053, B1=>nx5235);
   ix5298 : nor02_2x port map ( Y=>nx4636, A0=>nx4632, A1=>nx4633);
   ix5299 : nor02_2x port map ( Y=>nx4637, A0=>nx4619, A1=>nx4620);
   ix5300 : nand03_2x port map ( Y=>nx4638, A0=>nx4905, A1=>nx4907, A2=>
      nx4909);
   ix5301 : nand02_2x port map ( Y=>nx4639, A0=>nx4904, A1=>nx4638);
   ix5302 : ao21 port map ( Y=>nx4640, A0=>nx5027, A1=>nx5235, B0=>nx4631);
   ix5303 : aoi22 port map ( Y=>nx4641, A0=>nx2210, A1=>nx4640, B0=>nx4406, 
      B1=>nx4626);
   ix5304 : and02 port map ( Y=>nx4642, A0=>nx4406, A1=>nx4626);
   ix5305 : inv02 port map ( Y=>nx4643, A=>positive_M_1);
   ix5306 : nor02_2x port map ( Y=>nx4644, A0=>nx4643, A1=>nx4274_XX0_XREP44
   );
   ix5307 : inv02 port map ( Y=>nx4645, A=>negative_M_1);
   ix5308 : nor02_2x port map ( Y=>nx4646, A0=>nx4645, A1=>nx4262);
   ix5309 : nor04_2x port map ( Y=>nx4647, A0=>nx4644, A1=>nx4646, A2=>
      nx4462, A3=>nx4472);
   ix5310 : inv01 port map ( Y=>nx4648, A=>positive_2M_1);
   ix5311 : aoi22 port map ( Y=>nx4649, A0=>nx4645, A1=>nx4648, B0=>nx4262, 
      B1=>nx4648);
   ix5312 : nor02_2x port map ( Y=>nx4650, A0=>nx4649, A1=>nx4644);
   ix5313 : inv01 port map ( Y=>nx4651, A=>nx3498);
   ix5314 : and03 port map ( Y=>nx4652, A0=>nx268, A1=>aux_product_0, A2=>
      nx4651);
   ix5315 : and02 port map ( Y=>nx4653, A0=>aux_product_0, A1=>nx268);
   reg_nx3526 : inv02 port map ( Y=>nx3526, A=>nx4690);
   reg_nx3492 : nand02_2x port map ( Y=>nx3492, A0=>aux_product_0, A1=>nx268
   );
   ix5316 : nor02_2x port map ( Y=>nx4654, A0=>nx4711, A1=>nx3498);
   reg_nx368 : ao21 port map ( Y=>nx368, A0=>nx3498, A1=>nx4711, B0=>nx4654
   );
   ix5317 : and02 port map ( Y=>nx4655, A0=>nx4931, A1=>nx1970);
   ix5318 : oai32 port map ( Y=>nx4656, A0=>nx1970, A1=>nx4922, A2=>nx5224, 
      B0=>nx4932, B1=>nx5230);
   ix5319 : inv01 port map ( Y=>nx4657, A=>nx4641);
   ix5320 : nand02_2x port map ( Y=>nx4658, A0=>nx4639, A1=>nx4657);
   reg_nx4158 : aoi322 port map ( Y=>nx4158, A0=>nx4683, A1=>nx4898, A2=>
      nx4655, B0=>nx4656, B1=>nx4898, C0=>nx4658, C1=>nx4895);
   ix5321 : inv01 port map ( Y=>nx4659, A=>nx1970);
   reg_nx4032 : ao22 port map ( Y=>nx4032, A0=>nx5224, A1=>nx4659, B0=>
      nx4011, B1=>nx1970);
   ix5322 : aoi22 port map ( Y=>nx4660, A0=>nx5236, A1=>nx4880, B0=>nx4888, 
      B1=>nx4116);
   ix5323 : inv01 port map ( Y=>nx4661, A=>nx5236);
   reg_nx4137 : oai22 port map ( Y=>nx4137, A0=>nx4661, A1=>nx5129, B0=>
      nx4884, B1=>nx5154);
   ix5324 : nand03_2x port map ( Y=>nx4662, A0=>nx5144, A1=>nx5229, A2=>
      nx4452);
   reg_nx3358 : oai422 port map ( Y=>nx3358, A0=>nx4660, A1=>nx5145, A2=>
      nx5227, A3=>nx5233, B0=>nx4137, B1=>nx4662, C0=>nx5229, C1=>nx4132);
   ix5325 : inv02 port map ( Y=>nx4663, A=>negative_M_1);
   ix5326 : inv02 port map ( Y=>nx4664, A=>positive_M_1);
   reg_nx458 : oai22 port map ( Y=>nx458, A0=>nx4663, A1=>nx4322_XX0_XREP40, 
      B0=>nx4664, B1=>nx5208);
   reg_nx3529 : aoi221 port map ( Y=>nx3529, A0=>positive_M_2, A1=>nx4276, 
      B0=>negative_M_2, B1=>nx4264, C0=>nx458);
   ix5327 : inv02 port map ( Y=>nx4665, A=>nx3521);
   reg_nx462 : inv01 port map ( Y=>nx462, A=>nx4692);
   reg_nx4472 : inv02 port map ( Y=>nx4472, A=>nx4322_XX0_XREP40);
   reg_nx4462 : inv02 port map ( Y=>nx4462, A=>nx5209);
   ix5328 : nor02_2x port map ( Y=>nx4666, A0=>nx4808, A1=>nx4919);
   ix5329 : and02 port map ( Y=>nx4667, A0=>nx5220, A1=>nx4790);
   ix5330 : oai32 port map ( Y=>nx4668, A0=>nx4791, A1=>nx4786, A2=>nx5200, 
      B0=>nx5220, B1=>nx5931);
   ix5331 : inv01 port map ( Y=>nx4669, A=>nx5222);
   ix5332 : inv01 port map ( Y=>nx4670, A=>nx4655);
   ix5333 : aoi21 port map ( Y=>nx4671, A0=>nx4808, A1=>nx4669, B0=>nx4670);
   ix5334 : nor02_2x port map ( Y=>nx4672, A0=>nx4617, A1=>nx4616);
   ix5335 : oai21 port map ( Y=>nx4673, A0=>nx5169, A1=>nx4616, B0=>nx4615);
   ix5336 : inv01 port map ( Y=>nx4674, A=>nx4617);
   ix5337 : nand03_2x port map ( Y=>nx4675, A0=>nx4723, A1=>nx5220, A2=>
      nx4792);
   ix5338 : nor02_2x port map ( Y=>nx4676, A0=>nx3951, A1=>nx4793);
   ix5339 : aoi22 port map ( Y=>nx4677, A0=>nx5931, A1=>nx4787, B0=>nx5221, 
      B1=>nx4676);
   reg_nx3990 : nand02_2x port map ( Y=>nx3990, A0=>nx4675, A1=>nx4677);
   reg_nx3969 : ao22 port map ( Y=>nx3969, A0=>nx5200, A1=>nx4804, B0=>
      nx4724, B1=>nx4794);
   ix5340 : inv01 port map ( Y=>nx4678, A=>nx1660);
   ix5341 : and02 port map ( Y=>nx4679, A0=>nx5222, A1=>nx4808);
   ix5342 : nor02_2x port map ( Y=>nx4680, A0=>nx4679, A1=>nx4783);
   ix5343 : inv01 port map ( Y=>nx4681, A=>nx5230);
   ix5344 : nand02_2x port map ( Y=>nx4682, A0=>nx4930, A1=>nx4681);
   ix5345 : inv01 port map ( Y=>nx4683, A=>nx4011);
   reg_nx3917 : ao22 port map ( Y=>nx3917, A0=>nx4376, A1=>nx4678, B0=>
      nx4709, B1=>nx1660);
   ix5346 : inv01 port map ( Y=>nx4684, A=>nx4653);
   ix5347 : inv02 port map ( Y=>nx4685, A=>nx4651);
   ix5348 : inv02 port map ( Y=>nx4686, A=>nx4665);
   ix5349 : oai21 port map ( Y=>nx4687, A0=>nx4653, A1=>nx4651, B0=>nx4665);
   reg_nx3555 : inv02 port map ( Y=>nx3555, A=>nx4816);
   ix5350 : nor02_2x port map ( Y=>nx4688, A0=>nx4653, A1=>nx4651);
   ix5351 : nor02_2x port map ( Y=>nx4689, A0=>nx4711, A1=>nx4652);
   ix5352 : nor02_2x port map ( Y=>nx4690, A0=>nx4688, A1=>nx4689);
   ix5353 : inv01 port map ( Y=>nx4691, A=>nx3529);
   ix5354 : oai22 port map ( Y=>nx4692, A0=>nx4686, A1=>nx5915, B0=>nx4691, 
      B1=>nx4665);
   ix5355 : inv01 port map ( Y=>nx4693, A=>nx1660);
   ix5356 : nor03_2x port map ( Y=>nx4694, A0=>nx4693, A1=>nx5218, A2=>
      nx4806);
   ix5357 : inv01 port map ( Y=>nx4695, A=>nx3839);
   ix5358 : inv01 port map ( Y=>nx4696, A=>nx3867);
   ix5359 : oai32 port map ( Y=>nx4697, A0=>nx5075, A1=>nx5067, A2=>nx4695, 
      B0=>nx4696, B1=>nx5073);
   ix5360 : nor02_2x port map ( Y=>nx4698, A0=>nx5218, A1=>nx5925);
   ix5361 : inv01 port map ( Y=>nx4699, A=>nx3920);
   ix5362 : oai21 port map ( Y=>nx4700, A0=>nx4699, A1=>nx5184, B0=>nx4680);
   ix5363 : aoi322 port map ( Y=>nx4701, A0=>nx5074, A1=>nx5951, A2=>nx5071, 
      B0=>nx5949, B1=>nx5067, C0=>nx4944, C1=>nx5072);
   ix5364 : inv01 port map ( Y=>nx4702, A=>nx4678);
   ix5365 : inv01 port map ( Y=>nx4703, A=>nx4376);
   ix5366 : nor02_2x port map ( Y=>nx4704, A0=>nx4376, A1=>nx5911);
   ix5367 : aoi33 port map ( Y=>nx4705, A0=>nx5186, A1=>nx4693, A2=>nx4703, 
      B0=>nx5185, B1=>nx4693, B2=>nx4702);
   ix5368 : aoi33 port map ( Y=>nx4706, A0=>nx4693, A1=>nx4703, A2=>nx4699, 
      B0=>nx4702, B1=>nx4693, B2=>nx4699);
   ix5369 : aoi22 port map ( Y=>nx4707, A0=>nx5218, A1=>nx4699, B0=>nx5218, 
      B1=>nx5187);
   ix5370 : nand03_2x port map ( Y=>nx4708, A0=>nx4705, A1=>nx4706, A2=>
      nx4707);
   reg_nx3892 : inv01 port map ( Y=>nx3892, A=>nx4701);
   ix5371 : inv01 port map ( Y=>nx4709, A=>nx4701);
   reg_nx3864 : ao22 port map ( Y=>nx3864, A0=>nx5951, A1=>nx5071, B0=>
      nx3836, B1=>nx5076);
   ix5372 : aoi221 port map ( Y=>nx4710, A0=>negative_M_3, A1=>nx4264, B0=>
      positive_M_3, B1=>nx4276, C0=>nx552);
   ix5373 : nor02_2x port map ( Y=>nx4711, A0=>nx4647, A1=>nx4650);
   ix5374 : inv01 port map ( Y=>nx4712, A=>nx4652);
   ix5375 : aoi22 port map ( Y=>nx4713, A0=>nx4686, A1=>nx4712, B0=>nx5915, 
      B1=>nx4712);
   ix5376 : nor02_2x port map ( Y=>nx4714, A0=>nx4711, A1=>nx4713);
   reg_nx3579 : inv02 port map ( Y=>nx3579, A=>nx4745);
   ix5377 : inv02 port map ( Y=>nx4715, A=>nx3550);
   ix5378 : nand02_2x port map ( Y=>nx4716, A0=>nx4715, A1=>nx5917);
   reg_nx556 : oai21 port map ( Y=>nx556, A0=>nx4715, A1=>nx5917, B0=>nx4716
   );
   ix5379 : nand02_2x port map ( Y=>nx4717, A0=>nx4673, A1=>nx4674);
   ix5380 : and02 port map ( Y=>nx4718, A0=>nx4703, A1=>nx5188);
   ix5381 : oai22 port map ( Y=>nx4719, A0=>nx4718, A1=>nx4702, B0=>nx4699, 
      B1=>nx5189);
   ix5382 : nor02ii port map ( Y=>nx4720, A0=>nx4704, A1=>nx4719);
   ix5383 : inv01 port map ( Y=>nx4721, A=>nx4708);
   ix5384 : aoi22 port map ( Y=>nx4722, A0=>nx4912, A1=>nx4721, B0=>nx4720, 
      B1=>nx4721);
   reg_nx3948 : inv01 port map ( Y=>nx3948, A=>nx4722);
   ix5385 : inv01 port map ( Y=>nx4723, A=>nx4722);
   ix5386 : inv01 port map ( Y=>nx4724, A=>nx4722);
   ix5387 : inv01 port map ( Y=>nx4725, A=>nx1308);
   ix5388 : and02 port map ( Y=>nx4726, A0=>nx5905, A1=>nx4955);
   ix5389 : aoi322 port map ( Y=>nx4727, A0=>nx5905, A1=>nx5935, A2=>nx5214, 
      B0=>nx5953, B1=>nx4725, C0=>nx4748, C1=>nx4726);
   ix5390 : nand02_2x port map ( Y=>nx4728, A0=>nx5072, A1=>nx4996);
   ix5391 : inv01 port map ( Y=>nx4729, A=>nx3811);
   ix5392 : nor02_2x port map ( Y=>nx4730, A0=>nx4729, A1=>nx4997);
   ix5393 : aoi21 port map ( Y=>nx4731, A0=>nx5072, A1=>nx4730, B0=>nx4697);
   ix5394 : nand02_2x port map ( Y=>nx4732, A0=>nx5905, A1=>nx4956);
   ix5395 : inv01 port map ( Y=>nx4733, A=>nx3755);
   ix5396 : inv01 port map ( Y=>nx4734, A=>nx3783);
   ix5397 : aoi32 port map ( Y=>nx4735, A0=>nx5905, A1=>nx5214, A2=>nx4733, 
      B0=>nx4725, B1=>nx4734);
   ix5398 : inv01 port map ( Y=>nx4736, A=>nx5072);
   ix5399 : aoi21 port map ( Y=>nx4737, A0=>nx4729, A1=>nx5216, B0=>nx4736);
   ix5400 : inv01 port map ( Y=>nx4738, A=>nx4697);
   ix5401 : and02 port map ( Y=>nx4739, A0=>nx4998, A1=>nx5905);
   ix5402 : nor02_2x port map ( Y=>nx4740, A0=>nx4733, A1=>nx4957);
   ix5403 : oai32 port map ( Y=>nx4741, A0=>nx5905, A1=>nx5216, A2=>nx4734, 
      B0=>nx4729, B1=>nx4999);
   reg_nx3808 : inv01 port map ( Y=>nx3808, A=>nx4727);
   reg_nx3780 : ao22 port map ( Y=>nx3780, A0=>nx5935, A1=>nx5214, B0=>
      nx4749, B1=>nx4958);
   ix5404 : inv01 port map ( Y=>nx4742, A=>nx3582);
   ix5405 : nor02_2x port map ( Y=>nx4743, A0=>nx4816, A1=>nx4814);
   ix5406 : nor02_2x port map ( Y=>nx4744, A0=>nx4743, A1=>nx4831);
   reg_nx3612 : oai22 port map ( Y=>nx3612, A0=>nx4742, A1=>nx650, B0=>
      nx4826, B1=>nx4744);
   ix5407 : ao22 port map ( Y=>nx4745, A0=>nx4816, A1=>nx4830, B0=>nx4814, 
      B1=>nx4830);
   ix5408 : inv01 port map ( Y=>nx4746, A=>nx3643);
   ix5409 : inv01 port map ( Y=>nx4747, A=>nx3671);
   reg_nx3752 : inv02 port map ( Y=>nx3752, A=>nx5102);
   ix5410 : inv01 port map ( Y=>nx4748, A=>nx5957);
   ix5411 : inv01 port map ( Y=>nx4749, A=>nx5957);
   ix5412 : nor02_2x port map ( Y=>nx4750, A0=>nx4746, A1=>nx4827);
   ix5413 : aoi22 port map ( Y=>nx4751, A0=>nx3671, A1=>nx5057, B0=>nx932, 
      B1=>nx4750);
   reg_nx3724 : oai422 port map ( Y=>nx3724, A0=>nx5945, A1=>nx4822, A2=>
      nx5058, A3=>nx4825, B0=>nx5012, B1=>nx5009, C0=>nx5945, C1=>nx4751);
   reg_nx3696 : oai332 port map ( Y=>nx3696, A0=>nx5060, A1=>nx4825, A2=>
      nx4823, B0=>nx5059, B1=>nx4746, B2=>nx4828, C0=>nx4747, C1=>nx932);
   reg_nx3668 : oai22 port map ( Y=>nx3668, A0=>nx4746, A1=>nx4829, B0=>
      nx4825, B1=>nx4824);
   ix5414 : or02 port map ( Y=>nx4752, A0=>nx5995, A1=>nx5997);
   reg_nx492 : nor04_2x port map ( Y=>nx492, A0=>nx5997, A1=>nx5999, A2=>
      nx6007, A3=>nx6003);
   ix5415 : inv01 port map ( Y=>nx4753, A=>nx4752);
   ix5416 : nor02_2x port map ( Y=>nx4754, A0=>nx5999, A1=>nx6007);
   ix5417 : inv01 port map ( Y=>nx4755, A=>M(1));
   ix5418 : or03 port map ( Y=>nx4756, A0=>nx6003, A1=>nx5999, A2=>nx6009);
   ix5419 : inv02 port map ( Y=>nx4757, A=>nx5993);
   ix5420 : aoi422 port map ( Y=>nx4758, A0=>nx4753, A1=>nx4754, A2=>nx5993, 
      A3=>nx4755, B0=>nx4756, B1=>nx4757, C0=>nx4752, C1=>nx4757);
   ix5421 : inv02 port map ( Y=>nx4759, A=>nx5989);
   ix5422 : nand02_2x port map ( Y=>nx4760, A0=>nx5989, A1=>nx5991);
   ix5423 : nand04_2x port map ( Y=>nx4761, A0=>nx4978, A1=>nx4979, A2=>
      nx4759, A3=>nx4980);
   ix5424 : oai321 port map ( Y=>nx4762, A0=>nx4979, A1=>nx4759, A2=>nx4980, 
      B0=>nx4978, B1=>nx4760, C0=>nx4761);
   ix5425 : inv02 port map ( Y=>nx4763, A=>nx508);
   ix5426 : inv02 port map ( Y=>nx4764, A=>nx5995);
   ix5427 : inv01 port map ( Y=>nx4765, A=>nx492);
   ix5428 : aoi22 port map ( Y=>nx4766, A0=>nx492, A1=>nx4764, B0=>nx5995, 
      B1=>nx4765);
   ix5429 : inv02 port map ( Y=>nx4767, A=>nx4978);
   ix5430 : inv01 port map ( Y=>nx4768, A=>nx4979);
   ix5431 : and02 port map ( Y=>nx4769, A0=>nx4979, A1=>nx4980);
   reg_nx876 : oai422 port map ( Y=>nx876, A0=>nx4767, A1=>nx4768, A2=>
      nx4759, A3=>nx5991, B0=>nx4769, B1=>nx5989, C0=>nx4978, C1=>nx5989);
   ix5432 : aoi322 port map ( Y=>nx4770, A0=>nx4978, A1=>nx5991, A2=>nx4979, 
      B0=>nx4767, B1=>nx4980, C0=>nx4768, C1=>nx4980);
   reg_nx782 : inv01 port map ( Y=>nx782, A=>nx4770);
   ix5433 : inv01 port map ( Y=>nx4771, A=>nx4770);
   ix5434 : inv01 port map ( Y=>nx4772, A=>nx4770);
   reg_nx696 : and02 port map ( Y=>nx696, A0=>nx5210, A1=>nx5212);
   reg_nx688 : inv02 port map ( Y=>nx688, A=>nx5212);
   ix5435 : inv02 port map ( Y=>nx4773, A=>nx5212);
   reg_nx594 : oai22 port map ( Y=>nx594, A0=>nx4764, A1=>nx4765, B0=>nx5995, 
      B1=>nx492);
   ix5436 : inv01 port map ( Y=>nx4774, A=>nx4659);
   ix5437 : nand02_2x port map ( Y=>nx4775, A0=>nx5933, A1=>nx4774);
   ix5438 : inv01 port map ( Y=>nx4776, A=>nx5097);
   ix5439 : and02 port map ( Y=>nx4777, A0=>nx5224, A1=>nx4659);
   reg_nx4276 : inv01 port map ( Y=>nx4276, A=>nx4274_XX0_XREP44);
   reg_nx4264 : inv01 port map ( Y=>nx4264, A=>nx4262);
   ix5440 : inv02 port map ( Y=>nx4778, A=>negative_M_6);
   ix5441 : inv02 port map ( Y=>nx4779, A=>positive_M_6);
   reg_nx928 : oai22 port map ( Y=>nx928, A0=>nx4778, A1=>nx4322_XX0_XREP40, 
      B0=>nx4779, B1=>nx5209);
   reg_nx3671 : aoi221 port map ( Y=>nx3671, A0=>positive_M_7, A1=>nx4276, 
      B0=>negative_M_7, B1=>nx4264, C0=>nx928);
   ix5442 : inv02 port map ( Y=>nx4780, A=>nx3663);
   ix5443 : and02 port map ( Y=>nx4781, A0=>nx3964, A1=>nx3943);
   ix5444 : aoi322 port map ( Y=>nx4782, A0=>nx5200, A1=>nx3943, A2=>nx5931, 
      B0=>nx5200, B1=>nx4781, C0=>nx5931, C1=>nx3964);
   ix5445 : inv01 port map ( Y=>nx4783, A=>nx4782);
   ix5446 : inv02 port map ( Y=>nx4784, A=>nx3964);
   ix5447 : nor02_2x port map ( Y=>nx4785, A0=>nx5931, A1=>nx3964);
   ix5448 : inv01 port map ( Y=>nx4786, A=>nx5221);
   ix5449 : inv02 port map ( Y=>nx4787, A=>nx5221);
   reg_nx3951 : inv02 port map ( Y=>nx3951, A=>nx5200);
   ix5450 : inv02 port map ( Y=>nx4788, A=>nx3943);
   ix5451 : and02 port map ( Y=>nx4789, A0=>nx5200, A1=>nx4788);
   reg_nx1790 : inv02 port map ( Y=>nx1790, A=>nx4804);
   ix5452 : inv01 port map ( Y=>nx4790, A=>nx4804);
   ix5453 : inv01 port map ( Y=>nx4791, A=>nx4804);
   ix5454 : inv02 port map ( Y=>nx4792, A=>nx4804);
   ix5455 : inv02 port map ( Y=>nx4793, A=>nx4804);
   ix5456 : inv02 port map ( Y=>nx4794, A=>nx4804);
   ix5457 : or02 port map ( Y=>nx4795, A0=>nx4784, A1=>nx5931);
   reg_nx1850 : aoi21 port map ( Y=>nx1850, A0=>nx3964, A1=>nx4795, B0=>
      nx4785);
   ix5458 : inv01 port map ( Y=>nx4796, A=>nx4782);
   ix5459 : and02 port map ( Y=>nx4797, A0=>nx5222, A1=>nx3985);
   ix5460 : inv01 port map ( Y=>nx4798, A=>nx5222);
   ix5461 : inv02 port map ( Y=>nx4799, A=>nx3985);
   ix5462 : oai21 port map ( Y=>nx4800, A0=>nx4798, A1=>nx4799, B0=>nx4782);
   ix5463 : oai332 port map ( Y=>nx4801, A0=>nx5221, A1=>nx4796, A2=>nx4797, 
      B0=>nx4800, B1=>nx4789, B2=>nx5196, C0=>nx5223, C1=>nx3985);
   ix5464 : nor02_2x port map ( Y=>nx4802, A0=>nx5223, A1=>nx3985);
   ix5465 : inv01 port map ( Y=>nx4803, A=>nx4802);
   ix5466 : nor02_2x port map ( Y=>nx4804, A0=>nx4789, A1=>nx5197);
   ix5467 : nor02_2x port map ( Y=>nx4805, A0=>nx4804, A1=>nx4802);
   ix5468 : aoi222 port map ( Y=>nx4806, A0=>nx5223, A1=>nx3985, B0=>nx4803, 
      B1=>nx4796, C0=>nx5221, C1=>nx4805);
   ix5469 : inv01 port map ( Y=>nx4807, A=>nx4806);
   ix5470 : ao21 port map ( Y=>nx4808, A0=>nx5223, A1=>nx3985, B0=>nx4802);
   reg_nx1910 : oai22 port map ( Y=>nx1910, A0=>nx4798, A1=>nx3985, B0=>
      nx4799, B1=>nx5223);
   ix5471 : inv01 port map ( Y=>nx4809, A=>nx3615);
   ix5472 : inv02 port map ( Y=>nx4810, A=>nx3607);
   ix5473 : aoi22 port map ( Y=>nx4811, A0=>nx3615, A1=>nx4810, B0=>nx3607, 
      B1=>nx4809);
   ix5474 : inv01 port map ( Y=>nx4812, A=>nx5907);
   ix5475 : inv02 port map ( Y=>nx4813, A=>nx3574);
   ix5476 : nor02_2x port map ( Y=>nx4814, A0=>nx5917, A1=>nx3550);
   ix5477 : aoi22 port map ( Y=>nx4815, A0=>nx5917, A1=>nx3550, B0=>nx5907, 
      B1=>nx3574);
   ix5478 : aoi321 port map ( Y=>nx4816, A0=>nx4684, A1=>nx4685, A2=>nx4686, 
      B0=>nx5915, B1=>nx4687, C0=>nx4714);
   ix5479 : aoi222 port map ( Y=>nx4817, A0=>nx4812, A1=>nx4813, B0=>nx4814, 
      B1=>nx4815, C0=>nx4816, C1=>nx4815);
   ix5480 : inv02 port map ( Y=>nx4818, A=>nx3635);
   ix5481 : inv01 port map ( Y=>nx4819, A=>nx5909);
   ix5482 : aoi22 port map ( Y=>nx4820, A0=>nx5909, A1=>nx4818, B0=>nx3635, 
      B1=>nx4819);
   ix5483 : nor02_2x port map ( Y=>nx4821, A0=>nx5061, A1=>nx4820);
   ix5484 : inv01 port map ( Y=>nx4822, A=>nx3640);
   ix5485 : inv01 port map ( Y=>nx4823, A=>nx3640);
   ix5486 : inv01 port map ( Y=>nx4824, A=>nx3640);
   ix5487 : oai22 port map ( Y=>nx4825, A0=>nx4818, A1=>nx4819, B0=>nx3635, 
      B1=>nx5909);
   reg_nx744 : oai22 port map ( Y=>nx744, A0=>nx4809, A1=>nx3607, B0=>nx4810, 
      B1=>nx3615);
   ix5488 : oai22 port map ( Y=>nx4826, A0=>nx4812, A1=>nx4813, B0=>nx5907, 
      B1=>nx3574);
   reg_nx650 : oai22 port map ( Y=>nx650, A0=>nx4813, A1=>nx5907, B0=>nx4812, 
      B1=>nx3574);
   reg_nx838 : inv01 port map ( Y=>nx838, A=>nx4820);
   ix5489 : inv01 port map ( Y=>nx4827, A=>nx4820);
   ix5490 : inv01 port map ( Y=>nx4828, A=>nx4820);
   ix5491 : inv01 port map ( Y=>nx4829, A=>nx4820);
   ix5492 : nand02_2x port map ( Y=>nx4830, A0=>nx5917, A1=>nx3550);
   ix5493 : and02 port map ( Y=>nx4831, A0=>nx5917, A1=>nx3550);
   reg_nx602 : nor02_2x port map ( Y=>nx602, A0=>nx4763, A1=>nx4766);
   ix5494 : inv02 port map ( Y=>nx4832, A=>nx5985);
   ix5495 : inv02 port map ( Y=>nx4833, A=>M(10));
   ix5496 : inv02 port map ( Y=>nx4834, A=>nx5981);
   ix5497 : and04 port map ( Y=>nx4835, A0=>nx5212, A1=>nx4832, A2=>nx4833, 
      A3=>nx4834);
   ix5498 : and04 port map ( Y=>nx4836, A0=>nx5213, A1=>nx5985, A2=>M(10), 
      A3=>nx5981);
   ix5499 : inv02 port map ( Y=>nx4837, A=>nx868);
   ix5500 : aoi44 port map ( Y=>nx4838, A0=>nx5211, A1=>nx4835, A2=>nx5939, 
      A3=>nx4762, B0=>nx5210, B1=>nx4836, B2=>nx4762, B3=>nx4837);
   reg_nx1166 : inv02 port map ( Y=>nx1166, A=>nx4838);
   ix5501 : inv02 port map ( Y=>nx4839, A=>nx4838);
   ix5502 : or02 port map ( Y=>nx4840, A0=>nx5985, A1=>nx5981);
   ix5503 : aoi422 port map ( Y=>nx4841, A0=>nx5939, A1=>nx4832, A2=>M(10), 
      A3=>nx4834, B0=>nx4840, B1=>nx4833, C0=>nx4833, C1=>nx4837);
   reg_nx1158 : inv02 port map ( Y=>nx1158, A=>nx4841);
   ix5504 : inv02 port map ( Y=>nx4842, A=>nx4841);
   ix5505 : and02 port map ( Y=>nx4843, A0=>nx5939, A1=>nx4762);
   ix5506 : nor02ii port map ( Y=>nx4844, A0=>nx5939, A1=>nx4762);
   ix5507 : and02 port map ( Y=>nx4845, A0=>nx5981, A1=>nx5985);
   ix5508 : aoi44 port map ( Y=>nx4846, A0=>nx4843, A1=>nx5211, A2=>nx5213, 
      A3=>nx4977, B0=>nx4844, B1=>nx5211, B2=>nx5213, B3=>nx4845);
   reg_nx1072 : inv02 port map ( Y=>nx1072, A=>nx4846);
   ix5509 : inv02 port map ( Y=>nx4847, A=>nx4846);
   reg_nx1064 : oai322 port map ( Y=>nx1064, A0=>nx4837, A1=>nx4834, A2=>
      nx5985, B0=>nx5981, B1=>nx5939, C0=>nx4832, C1=>nx5981);
   ix5510 : aoi44 port map ( Y=>nx4848, A0=>nx4843, A1=>nx5211, A2=>nx5213, 
      A3=>nx4832, B0=>nx4844, B1=>nx5211, B2=>nx5985, B3=>nx5213);
   reg_nx978 : inv02 port map ( Y=>nx978, A=>nx4848);
   ix5511 : inv02 port map ( Y=>nx4849, A=>nx4848);
   reg_nx970 : oai22 port map ( Y=>nx970, A0=>nx4832, A1=>nx4837, B0=>nx5985, 
      B1=>nx5939);
   ix5512 : oai21 port map ( Y=>nx4850, A0=>nx5216, A1=>nx4735, B0=>nx4737);
   ix5513 : nor02_2x port map ( Y=>nx4851, A0=>nx5216, A1=>nx4732);
   ix5514 : and02 port map ( Y=>nx4852, A0=>nx4738, A1=>nx4851);
   ix5515 : inv01 port map ( Y=>nx4853, A=>nx4694);
   ix5516 : nor02_2x port map ( Y=>nx4854, A0=>nx5216, A1=>nx4735);
   ix5517 : nor02ii port map ( Y=>nx4855, A0=>nx4854, A1=>nx4737);
   ix5518 : nand02_2x port map ( Y=>nx4856, A0=>nx5101, A1=>nx4855);
   ix5519 : nor02_2x port map ( Y=>nx4857, A0=>M(14), A1=>nx5971);
   ix5520 : inv02 port map ( Y=>nx4858, A=>nx5973);
   ix5521 : inv02 port map ( Y=>nx4859, A=>nx5977);
   ix5523 : and02 port map ( Y=>nx4861, A0=>M(14), A1=>nx5971);
   ix5524 : aoi44 port map ( Y=>nx4862, A0=>nx4877, A1=>nx4857, A2=>nx4858, 
      A3=>nx4859, B0=>nx5927, B1=>nx4861, B2=>nx5973, B3=>nx5977);
   reg_nx1542 : nor02_2x port map ( Y=>nx1542, A0=>nx4862, A1=>nx4838);
   ix5525 : nor02_2x port map ( Y=>nx4863, A0=>nx5973, A1=>nx5977);
   ix5526 : inv02 port map ( Y=>nx4864, A=>nx5971);
   ix5527 : or03 port map ( Y=>nx4865, A0=>nx5977, A1=>nx5971, A2=>nx5973);
   ix5528 : inv02 port map ( Y=>nx4866, A=>M(14));
   ix5529 : aoi422 port map ( Y=>nx4867, A0=>nx4877, A1=>nx4863, A2=>M(14), 
      A3=>nx4864, B0=>nx4865, B1=>nx4866, C0=>nx5927, C1=>nx4866);
   reg_nx1534 : inv02 port map ( Y=>nx1534, A=>nx4867);
   ix5530 : inv02 port map ( Y=>nx4868, A=>nx4867);
   ix5531 : aoi44 port map ( Y=>nx4869, A0=>nx4877, A1=>nx4859, A2=>nx4864, 
      A3=>nx4858, B0=>nx5927, B1=>nx5977, B2=>nx5971, B3=>nx5973);
   reg_nx1448 : nor02_2x port map ( Y=>nx1448, A0=>nx4869, A1=>nx4838);
   ix5532 : nor03_2x port map ( Y=>nx4870, A0=>nx5977, A1=>nx5971, A2=>
      nx5973);
   reg_nx1432 : and02 port map ( Y=>nx1432, A0=>nx4877, A1=>nx4870);
   ix5533 : inv02 port map ( Y=>nx4871, A=>nx4863);
   ix5534 : aoi422 port map ( Y=>nx4872, A0=>nx4878, A1=>nx4859, A2=>nx5971, 
      A3=>nx4858, B0=>nx4871, B1=>nx4864, C0=>nx5927, C1=>nx4864);
   reg_nx1440 : inv02 port map ( Y=>nx1440, A=>nx4872);
   ix5535 : inv02 port map ( Y=>nx4873, A=>nx4872);
   ix5536 : and02 port map ( Y=>nx4874, A0=>nx5973, A1=>nx5977);
   ix5537 : aoi22 port map ( Y=>nx4875, A0=>nx4878, A1=>nx4863, B0=>nx5927, 
      B1=>nx4874);
   reg_nx1354 : nor02_2x port map ( Y=>nx1354, A0=>nx4875, A1=>nx4838);
   reg_nx1346 : oai322 port map ( Y=>nx1346, A0=>nx5927, A1=>nx4858, A2=>
      nx5979, B0=>nx4878, B1=>nx5975, C0=>nx4859, C1=>nx5975);
   ix5538 : aoi22 port map ( Y=>nx4876, A0=>nx4878, A1=>nx4859, B0=>nx5979, 
      B1=>nx5927);
   reg_nx1260 : nor02_2x port map ( Y=>nx1260, A0=>nx4876, A1=>nx4838);
   reg_nx1252 : oai22 port map ( Y=>nx1252, A0=>nx4859, A1=>nx5929, B0=>
      nx4878, B1=>nx5979);
   ix5539 : buf04 port map ( Y=>nx4877, A=>nx1150);
   ix5540 : buf04 port map ( Y=>nx4878, A=>nx1150);
   reg_nx1846 : ao22 port map ( Y=>nx1846, A0=>negative_M_17, A1=>nx4476, B0
      =>positive_M_17, B1=>nx4466);
   reg_nx3972 : aoi221 port map ( Y=>nx3972, A0=>positive_M_18, A1=>nx4280, 
      B0=>negative_M_18, B1=>nx4268, C0=>nx1846);
   reg_nx4282 : inv01 port map ( Y=>nx4282, A=>nx4274);
   reg_nx4478 : inv01 port map ( Y=>nx4478, A=>nx4322);
   ix5541 : nor02_2x port map ( Y=>nx4879, A0=>nx5237, A1=>nx4111);
   ix5542 : inv02 port map ( Y=>nx4880, A=>nx5129);
   ix5543 : inv02 port map ( Y=>nx4881, A=>nx4111);
   ix5544 : and02 port map ( Y=>nx4882, A0=>nx5237, A1=>nx4881);
   ix5545 : nor02_2x port map ( Y=>nx4883, A0=>nx4881, A1=>nx5237);
   ix5546 : nor02_2x port map ( Y=>nx4884, A0=>nx4882, A1=>nx4883);
   reg_nx2270 : inv02 port map ( Y=>nx2270, A=>nx4884);
   ix5547 : inv02 port map ( Y=>nx4885, A=>nx4884);
   ix5548 : inv02 port map ( Y=>nx4886, A=>nx4884);
   ix5549 : inv01 port map ( Y=>nx4887, A=>nx4884);
   ix5550 : inv02 port map ( Y=>nx4888, A=>nx4884);
   reg_nx4053 : nor04_2x port map ( Y=>nx4053, A0=>nx5937, A1=>nx4966, A2=>
      nx5043, A3=>nx4964);
   ix5551 : and02 port map ( Y=>nx4889, A0=>nx4623, A1=>nx5129);
   ix5552 : oai22 port map ( Y=>nx4890, A0=>nx4889, A1=>nx5146, B0=>nx4623, 
      B1=>nx5140);
   ix5553 : and02 port map ( Y=>nx4891, A0=>nx4636, A1=>nx5132);
   ix5554 : inv01 port map ( Y=>nx4892, A=>nx4633);
   ix5555 : nor02_2x port map ( Y=>nx4893, A0=>nx4632, A1=>nx5124);
   ix5556 : nand02_2x port map ( Y=>nx4894, A0=>nx4623, A1=>nx5147);
   ix5557 : aoi44 port map ( Y=>nx4895, A0=>nx4890, A1=>nx4891, A2=>nx4892, 
      A3=>nx4893, B0=>nx4894, B1=>nx5169, B2=>nx4636, B3=>nx5136);
   ix5558 : inv01 port map ( Y=>nx4896, A=>nx4642);
   ix5559 : inv01 port map ( Y=>nx4897, A=>nx4631);
   ix5560 : and03 port map ( Y=>nx4898, A0=>nx4895, A1=>nx4896, A2=>nx4897);
   ix5561 : aoi21 port map ( Y=>nx4899, A0=>nx5148, A1=>nx5141, B0=>nx4632);
   ix5562 : nor02_2x port map ( Y=>nx4900, A0=>nx5169, A1=>nx4899);
   ix5563 : nor02_2x port map ( Y=>nx4901, A0=>nx4889, A1=>nx4633);
   ix5564 : nor02_2x port map ( Y=>nx4902, A0=>nx5169, A1=>nx4901);
   ix5565 : nand02_2x port map ( Y=>nx4903, A0=>nx4636, A1=>nx5136);
   ix5566 : or04 port map ( Y=>nx4904, A0=>nx4900, A1=>nx5171, A2=>nx4902, 
      A3=>nx4903);
   ix5567 : oai21 port map ( Y=>nx4905, A0=>nx4889, A1=>nx4633, B0=>nx5175);
   ix5568 : ao21 port map ( Y=>nx4906, A0=>nx5961, A1=>nx5142, B0=>nx4632);
   ix5569 : nand02_2x port map ( Y=>nx4907, A0=>nx5176, A1=>nx4906);
   ix5570 : and02 port map ( Y=>nx4908, A0=>nx4623, A1=>nx5961);
   ix5571 : oai21 port map ( Y=>nx4909, A0=>nx4908, A1=>nx5124, B0=>nx5177);
   ix5572 : nor02ii port map ( Y=>nx4910, A0=>nx5155, A1=>nx4717);
   ix5573 : nor02ii port map ( Y=>nx4911, A0=>nx4720, A1=>nx4701);
   reg_nx4221 : oai22 port map ( Y=>nx4221, A0=>nx4910, A1=>nx5206, B0=>
      nx4911, B1=>nx5205);
   ix5574 : inv01 port map ( Y=>nx4912, A=>nx4701);
   ix5575 : and02 port map ( Y=>nx4913, A0=>nx5230, A1=>nx4027);
   ix5576 : nor02_2x port map ( Y=>nx4914, A0=>nx5230, A1=>nx4027);
   ix5577 : inv01 port map ( Y=>nx4915, A=>nx5224);
   ix5578 : inv02 port map ( Y=>nx4916, A=>nx4006);
   ix5579 : nor03_2x port map ( Y=>nx4917, A0=>nx4914, A1=>nx4915, A2=>
      nx4916);
   ix5580 : nor04_2x port map ( Y=>nx4918, A0=>nx4913, A1=>nx4631, A2=>
      nx4917, A3=>nx4642);
   ix5581 : inv01 port map ( Y=>nx4919, A=>nx4918);
   ix5582 : inv01 port map ( Y=>nx4920, A=>nx4918);
   ix5583 : aoi21 port map ( Y=>nx4921, A0=>nx5230, A1=>nx4027, B0=>nx4914);
   ix5584 : inv01 port map ( Y=>nx4922, A=>nx4921);
   ix5585 : inv01 port map ( Y=>nx4923, A=>nx5933);
   ix5586 : inv01 port map ( Y=>nx4924, A=>nx5933);
   ix5587 : inv01 port map ( Y=>nx4925, A=>nx5933);
   ix5588 : inv01 port map ( Y=>nx4926, A=>nx5933);
   ix5589 : inv01 port map ( Y=>nx4927, A=>nx5933);
   reg_nx1970 : oai22 port map ( Y=>nx1970, A0=>nx4915, A1=>nx4006, B0=>
      nx4916, B1=>nx5224);
   ix5590 : inv02 port map ( Y=>nx4928, A=>nx4027);
   ix5591 : inv01 port map ( Y=>nx4929, A=>nx5231);
   ix5592 : aoi22 port map ( Y=>nx4930, A0=>nx5231, A1=>nx4928, B0=>nx4027, 
      B1=>nx4929);
   reg_nx2030 : inv01 port map ( Y=>nx2030, A=>nx4930);
   ix5593 : inv01 port map ( Y=>nx4931, A=>nx4930);
   ix5594 : inv01 port map ( Y=>nx4932, A=>nx4930);
   ix5595 : inv01 port map ( Y=>nx4933, A=>nx4930);
   ix5596 : inv01 port map ( Y=>nx4934, A=>nx4930);
   ix5597 : inv01 port map ( Y=>nx4935, A=>nx4930);
   ix5598 : inv02 port map ( Y=>nx4936, A=>nx3719);
   ix5599 : nor02ii port map ( Y=>nx4937, A0=>nx5079, A1=>nx4821);
   ix5600 : nand02_2x port map ( Y=>nx4938, A0=>nx4809, A1=>nx4811);
   ix5601 : and02 port map ( Y=>nx4939, A0=>nx5016, A1=>nx5010);
   ix5602 : aoi321 port map ( Y=>nx4940, A0=>nx4937, A1=>nx5063, A2=>nx4938, 
      B0=>nx5192, B1=>nx4939, C0=>nx5005);
   ix5603 : inv01 port map ( Y=>nx4941, A=>nx4739);
   ix5604 : inv01 port map ( Y=>nx4942, A=>nx4740);
   ix5605 : inv01 port map ( Y=>nx4943, A=>nx4741);
   ix5606 : oai321 port map ( Y=>nx4944, A0=>nx4940, A1=>nx5214, A2=>nx4941, 
      B0=>nx4941, B1=>nx4942, C0=>nx4943);
   ix5607 : and02 port map ( Y=>nx4945, A0=>nx4809, A1=>nx4811);
   ix5608 : ao21 port map ( Y=>nx4946, A0=>nx5017, A1=>nx5011, B0=>nx5006);
   ix5609 : or02 port map ( Y=>nx4947, A0=>nx5007, A1=>nx5192);
   ix5610 : oai21 port map ( Y=>nx4948, A0=>nx4740, A1=>nx4959, B0=>nx4739);
   reg_nx3836 : aoi32 port map ( Y=>nx3836, A0=>nx5957, A1=>nx4943, A2=>
      nx4942, B0=>nx4948, B1=>nx4943);
   reg_nx2326 : ao22 port map ( Y=>nx2326, A0=>negative_M_25, A1=>nx4478, B0
      =>positive_M_25, B1=>nx4468);
   reg_nx4140 : aoi221 port map ( Y=>nx4140, A0=>positive_M_26, A1=>nx4282, 
      B0=>negative_M_26, B1=>nx4270, C0=>nx2326);
   ix5611 : inv02 port map ( Y=>nx4949, A=>negative_M_9);
   ix5612 : inv02 port map ( Y=>nx4950, A=>positive_M_9);
   reg_nx1210 : oai22 port map ( Y=>nx1210, A0=>nx4949, A1=>
      nx4322_XX0_XREP40, B0=>nx4950, B1=>nx5209);
   reg_nx3755 : aoi221 port map ( Y=>nx3755, A0=>positive_M_10, A1=>nx4278, 
      B0=>negative_M_10, B1=>nx4266, C0=>nx1210);
   ix5613 : inv02 port map ( Y=>nx4951, A=>nx3747);
   ix5614 : and02 port map ( Y=>nx4952, A0=>nx5935, A1=>nx4951);
   ix5615 : nor02_2x port map ( Y=>nx4953, A0=>nx4951, A1=>nx5935);
   ix5616 : nor02_2x port map ( Y=>nx4954, A0=>nx4952, A1=>nx4953);
   reg_nx1214 : inv02 port map ( Y=>nx1214, A=>nx5214);
   ix5617 : inv01 port map ( Y=>nx4955, A=>nx5215);
   ix5618 : inv01 port map ( Y=>nx4956, A=>nx5215);
   ix5619 : inv01 port map ( Y=>nx4957, A=>nx5215);
   ix5620 : inv02 port map ( Y=>nx4958, A=>nx5215);
   ix5621 : inv02 port map ( Y=>nx4959, A=>nx5215);
   ix5622 : nand02_2x port map ( Y=>nx4960, A0=>nx4727, A1=>nx5919);
   ix5623 : nand02_2x port map ( Y=>nx4961, A0=>nx4728, A1=>nx5919);
   ix5624 : inv01 port map ( Y=>nx4962, A=>nx4853);
   ix5625 : inv01 port map ( Y=>nx4963, A=>nx5955);
   ix5626 : aoi321 port map ( Y=>nx4964, A0=>nx4960, A1=>nx4961, A2=>nx4962, 
      B0=>nx4682, B1=>nx4775, C0=>nx4963);
   ix5627 : aoi21 port map ( Y=>nx4965, A0=>nx4856, A1=>nx4738, B0=>nx4853);
   ix5628 : nor04_2x port map ( Y=>nx4966, A0=>nx4965, A1=>nx4776, A2=>
      nx4777, A3=>nx5231);
   ix5629 : oai22 port map ( Y=>nx4967, A0=>nx4924, A1=>nx4933, B0=>nx5225, 
      B1=>nx4923);
   ix5630 : nor02ii port map ( Y=>nx4968, A0=>nx5098, A1=>nx4967);
   reg_nx4011 : oai321 port map ( Y=>nx4011, A0=>nx4727, A1=>nx4853, A2=>
      nx4728, B0=>nx4853, B1=>nx5919, C0=>nx5955);
   ix5631 : inv01 port map ( Y=>nx4969, A=>nx4158);
   ix5632 : inv02 port map ( Y=>nx4970, A=>nx5241);
   ix5633 : and02 port map ( Y=>nx4971, A0=>nx5229, A1=>nx4452);
   reg_nx4155 : oai221 port map ( Y=>nx4155, A0=>nx4969, A1=>nx5241, B0=>
      nx4970, B1=>nx4158, C0=>nx4971);
   ix5634 : nor02_2x port map ( Y=>nx4972, A0=>nx5995, A1=>nx5997);
   ix5635 : nor02_2x port map ( Y=>nx4973, A0=>nx6005, A1=>nx5993);
   ix5636 : nor02_2x port map ( Y=>nx4974, A0=>nx5991, A1=>nx6001);
   ix5637 : nor04_2x port map ( Y=>nx4975, A0=>nx5981, A1=>nx6009, A2=>
      nx5989, A3=>nx5987);
   reg_nx1056 : and04 port map ( Y=>nx1056, A0=>nx4972, A1=>nx4973, A2=>
      nx4974, A3=>nx4975);
   ix5638 : nor02_2x port map ( Y=>nx4976, A0=>nx6009, A1=>nx5989);
   reg_nx868 : and04 port map ( Y=>nx868, A0=>nx4972, A1=>nx4974, A2=>nx4973, 
      A3=>nx4976);
   ix5639 : nor02_2x port map ( Y=>nx4977, A0=>nx5983, A1=>nx5987);
   ix5640 : nor02_2x port map ( Y=>nx4978, A0=>nx6005, A1=>nx6009);
   ix5641 : nor04_2x port map ( Y=>nx4979, A0=>nx5997, A1=>nx6001, A2=>
      nx5995, A3=>nx5993);
   ix5642 : inv02 port map ( Y=>nx4980, A=>nx5991);
   ix5643 : nor03_2x port map ( Y=>nx4981, A0=>nx4618, A1=>nx5227, A2=>
      nx5233);
   ix5644 : inv01 port map ( Y=>nx4982, A=>nx4158);
   ix5645 : nor02_2x port map ( Y=>nx4983, A0=>nx4621, A1=>nx4637);
   ix5646 : aoi32 port map ( Y=>nx4984, A0=>nx4158, A1=>nx5241, A2=>nx4981, 
      B0=>nx4982, B1=>nx4983);
   ix5647 : inv02 port map ( Y=>nx4985, A=>nx4304);
   ix5648 : inv02 port map ( Y=>nx4986, A=>nx4174);
   ix5649 : inv02 port map ( Y=>nx4987, A=>nx5241);
   ix5650 : aoi322 port map ( Y=>nx4988, A0=>nx4981, A1=>nx4412, A2=>nx4595, 
      B0=>nx4985, B1=>nx4986, C0=>nx4983, C1=>nx4987);
   reg_nx3378 : nand02_2x port map ( Y=>nx3378, A0=>nx4984, A1=>nx4988);
   reg_nx2146 : ao22 port map ( Y=>nx2146, A0=>negative_M_22, A1=>
      nx4478_XX0_XREP64, B0=>positive_M_22, B1=>nx4468);
   reg_nx4077 : aoi221 port map ( Y=>nx4077, A0=>positive_M_23, A1=>nx4282, 
      B0=>negative_M_23, B1=>nx4270, C0=>nx2146);
   reg_nx3408 : ao221 port map ( Y=>nx3408, A0=>nx4158, A1=>nx4596, B0=>
      nx4583, B1=>nx5045, C0=>nx5913);
   ix5651 : inv02 port map ( Y=>nx4989, A=>nx4132);
   reg_nx4266 : inv01 port map ( Y=>nx4266, A=>nx4262);
   ix5652 : inv02 port map ( Y=>nx4990, A=>negative_M_11);
   ix5653 : inv02 port map ( Y=>nx4991, A=>positive_M_11);
   reg_nx1398 : oai22 port map ( Y=>nx1398, A0=>nx4990, A1=>
      nx4322_XX0_XREP40, B0=>nx4991, B1=>nx5209);
   reg_nx3811 : aoi221 port map ( Y=>nx3811, A0=>positive_M_12, A1=>nx4278, 
      B0=>negative_M_12, B1=>nx4266, C0=>nx1398);
   ix5654 : inv02 port map ( Y=>nx4992, A=>nx3803);
   ix5655 : and02 port map ( Y=>nx4993, A0=>nx3811, A1=>nx4992);
   ix5656 : nor02_2x port map ( Y=>nx4994, A0=>nx4992, A1=>nx3811);
   ix5657 : nor02_2x port map ( Y=>nx4995, A0=>nx4993, A1=>nx4994);
   reg_nx1402 : inv02 port map ( Y=>nx1402, A=>nx5217);
   ix5658 : inv02 port map ( Y=>nx4996, A=>nx5217);
   ix5659 : inv01 port map ( Y=>nx4997, A=>nx5217);
   ix5660 : inv01 port map ( Y=>nx4998, A=>nx5217);
   ix5661 : inv01 port map ( Y=>nx4999, A=>nx5217);
   reg_nx4474 : inv01 port map ( Y=>nx4474, A=>nx4322_XX0_XREP40);
   reg_nx4464 : inv01 port map ( Y=>nx4464, A=>nx5209);
   reg_nx4278 : inv01 port map ( Y=>nx4278, A=>nx4274_XX0_XREP44);
   ix5662 : ao21 port map ( Y=>nx5000, A0=>nx3691, A1=>nx5947, B0=>nx3719);
   reg_nx1116 : ao22 port map ( Y=>nx1116, A0=>negative_M_8, A1=>nx4474, B0
      =>positive_M_8, B1=>nx4464);
   ix5663 : aoi221 port map ( Y=>nx5001, A0=>positive_M_9, A1=>nx4278, B0=>
      negative_M_9, B1=>nx4266, C0=>nx1116);
   ix5664 : inv02 port map ( Y=>nx5002, A=>nx3691);
   ix5665 : nor02_2x port map ( Y=>nx5003, A0=>nx5002, A1=>nx4936);
   ix5666 : aoi22 port map ( Y=>nx5004, A0=>nx5000, A1=>nx5943, B0=>nx5947, 
      B1=>nx5003);
   ix5667 : inv01 port map ( Y=>nx5005, A=>nx5004);
   ix5668 : inv01 port map ( Y=>nx5006, A=>nx5004);
   ix5669 : inv01 port map ( Y=>nx5007, A=>nx5004);
   reg_nx3699 : inv01 port map ( Y=>nx3699, A=>nx5044);
   ix5670 : aoi22 port map ( Y=>nx5008, A0=>nx3691, A1=>nx3699, B0=>nx5947, 
      B1=>nx5002);
   reg_nx1026 : inv01 port map ( Y=>nx1026, A=>nx5008);
   ix5671 : inv01 port map ( Y=>nx5009, A=>nx5945);
   ix5672 : inv01 port map ( Y=>nx5010, A=>nx5945);
   ix5673 : inv01 port map ( Y=>nx5011, A=>nx5945);
   ix5674 : inv01 port map ( Y=>nx5012, A=>nx5947);
   ix5675 : inv02 port map ( Y=>nx5013, A=>nx3719);
   ix5676 : nor02_2x port map ( Y=>nx5014, A0=>nx5943, A1=>nx4936);
   ix5677 : aoi21 port map ( Y=>nx5015, A0=>nx5943, A1=>nx5013, B0=>nx5014);
   reg_nx1120 : inv01 port map ( Y=>nx1120, A=>nx5015);
   ix5678 : inv01 port map ( Y=>nx5016, A=>nx5015);
   ix5679 : inv01 port map ( Y=>nx5017, A=>nx5015);
   ix5680 : inv02 port map ( Y=>nx5018, A=>nx4069);
   ix5681 : inv01 port map ( Y=>nx5019, A=>nx5941);
   ix5682 : aoi22 port map ( Y=>nx5020, A0=>nx5941, A1=>nx5018, B0=>nx4069, 
      B1=>nx5019);
   reg_nx2150 : inv01 port map ( Y=>nx2150, A=>nx5028);
   ix5683 : inv01 port map ( Y=>nx5021, A=>nx5028);
   ix5684 : inv01 port map ( Y=>nx5022, A=>nx5028);
   ix5685 : inv01 port map ( Y=>nx5023, A=>nx5028);
   ix5686 : inv01 port map ( Y=>nx5024, A=>nx5029);
   ix5687 : inv01 port map ( Y=>nx5025, A=>nx5029);
   ix5688 : inv01 port map ( Y=>nx5026, A=>nx5029);
   ix5689 : inv01 port map ( Y=>nx5027, A=>nx5029);
   ix5690 : buf02 port map ( Y=>nx5028, A=>nx5020);
   ix5691 : buf02 port map ( Y=>nx5029, A=>nx5020);
   ix5692 : inv01 port map ( Y=>nx5030, A=>nx4655);
   ix5693 : nor02_2x port map ( Y=>nx5031, A0=>nx5225, A1=>nx4926);
   ix5694 : nor02_2x port map ( Y=>nx5032, A0=>nx4927, A1=>nx4934);
   ix5695 : nand02_2x port map ( Y=>nx5033, A0=>nx5225, A1=>nx4935);
   ix5696 : inv01 port map ( Y=>nx5034, A=>nx5231);
   ix5697 : inv01 port map ( Y=>nx5035, A=>nx4659);
   ix5698 : ao21 port map ( Y=>nx5036, A0=>nx5033, A1=>nx5034, B0=>nx5035);
   ix5699 : aoi21 port map ( Y=>nx5037, A0=>nx5231, A1=>nx4925, B0=>nx4655);
   ix5700 : aoi222 port map ( Y=>nx5038, A0=>nx5030, A1=>nx5031, B0=>nx5030, 
      B1=>nx5032, C0=>nx5036, C1=>nx5037);
   ix5701 : and04 port map ( Y=>nx5039, A0=>nx5021, A1=>nx5169, A2=>nx2210, 
      A3=>nx5235);
   ix5702 : nand02_2x port map ( Y=>nx5040, A0=>nx5038, A1=>nx5039);
   ix5703 : nand03_2x port map ( Y=>nx5041, A0=>nx4935, A1=>nx4659, A2=>
      nx5225);
   ix5704 : oai222 port map ( Y=>nx5042, A0=>nx4659, A1=>nx4925, B0=>nx5225, 
      B1=>nx4926, C0=>nx4927, C1=>nx4934);
   ix5705 : ao32 port map ( Y=>nx5043, A0=>nx5041, A1=>nx5030, A2=>nx5034, 
      B0=>nx5042, B1=>nx5030);
   reg_nx1022 : ao22 port map ( Y=>nx1022, A0=>negative_M_7, A1=>nx4474, B0
      =>positive_M_7, B1=>nx4464);
   ix5706 : aoi221 port map ( Y=>nx5044, A0=>positive_M_8, A1=>nx4278, B0=>
      nx4266, B1=>negative_M_8, C0=>nx1022);
   ix5707 : inv01 port map ( Y=>nx5045, A=>nx4221);
   ix5708 : and02 port map ( Y=>nx5046, A0=>positive_M_24, A1=>nx4468);
   ix5709 : and02 port map ( Y=>nx5047, A0=>positive_M_25, A1=>nx4282);
   ix5710 : and02 port map ( Y=>nx5048, A0=>negative_M_25, A1=>nx4270);
   ix5711 : inv02 port map ( Y=>nx5049, A=>nx4111);
   ix5712 : ao21 port map ( Y=>nx5050, A0=>negative_M_24, A1=>nx4478, B0=>
      nx5049);
   ix5713 : nor04_2x port map ( Y=>nx5051, A0=>nx5046, A1=>nx5047, A2=>
      nx5048, A3=>nx5050);
   ix5714 : inv01 port map ( Y=>nx5052, A=>nx5129);
   ix5715 : and02 port map ( Y=>nx5053, A0=>negative_M_24, A1=>nx4478);
   reg_nx4119 : nor04_2x port map ( Y=>nx4119, A0=>nx5046, A1=>nx5053, A2=>
      nx5048, A3=>nx5047);
   ix5716 : inv01 port map ( Y=>nx5054, A=>nx3671);
   ix5717 : inv02 port map ( Y=>nx5055, A=>nx4780);
   ix5718 : aoi22 port map ( Y=>nx5056, A0=>nx4780, A1=>nx5054, B0=>nx3671, 
      B1=>nx5055);
   ix5719 : inv01 port map ( Y=>nx5057, A=>nx5062);
   ix5720 : inv01 port map ( Y=>nx5058, A=>nx5062);
   ix5721 : inv01 port map ( Y=>nx5059, A=>nx5062);
   ix5722 : inv01 port map ( Y=>nx5060, A=>nx5062);
   ix5723 : inv01 port map ( Y=>nx5061, A=>nx932);
   ix5724 : buf02 port map ( Y=>nx5062, A=>nx5056);
   reg_nx932 : buf02 port map ( Y=>nx932, A=>nx5056);
   ix5725 : nor02_2x port map ( Y=>nx5063, A0=>nx5015, A1=>nx5945);
   reg_nx1586 : ao22 port map ( Y=>nx1586, A0=>negative_M_13, A1=>nx4476, B0
      =>positive_M_13, B1=>nx4466);
   reg_nx3867 : aoi221 port map ( Y=>nx3867, A0=>positive_M_14, A1=>nx4278, 
      B0=>negative_M_14, B1=>nx4266, C0=>nx1586);
   ix5726 : inv02 port map ( Y=>nx5064, A=>nx3859);
   ix5727 : and02 port map ( Y=>nx5065, A0=>nx5949, A1=>nx5064);
   ix5728 : nor02_2x port map ( Y=>nx5066, A0=>nx5064, A1=>nx5949);
   ix5729 : nor02_2x port map ( Y=>nx5067, A0=>nx5065, A1=>nx5066);
   reg_nx1492 : ao22 port map ( Y=>nx1492, A0=>negative_M_12, A1=>nx4474, B0
      =>positive_M_12, B1=>nx4464);
   reg_nx3839 : aoi221 port map ( Y=>nx3839, A0=>nx4278, A1=>positive_M_13, 
      B0=>nx4266, B1=>negative_M_13, C0=>nx1492);
   ix5730 : inv02 port map ( Y=>nx5068, A=>nx3831);
   ix5731 : and02 port map ( Y=>nx5069, A0=>nx5951, A1=>nx5068);
   ix5732 : nor02_2x port map ( Y=>nx5070, A0=>nx5068, A1=>nx5951);
   ix5733 : nor02_2x port map ( Y=>nx5071, A0=>nx5069, A1=>nx5070);
   ix5734 : nor02_2x port map ( Y=>nx5072, A0=>nx5067, A1=>nx5071);
   reg_nx1590 : inv02 port map ( Y=>nx1590, A=>nx5067);
   ix5735 : inv01 port map ( Y=>nx5073, A=>nx5067);
   ix5736 : inv01 port map ( Y=>nx5074, A=>nx5067);
   reg_nx1496 : inv02 port map ( Y=>nx1496, A=>nx5071);
   ix5737 : inv01 port map ( Y=>nx5075, A=>nx5071);
   ix5738 : inv02 port map ( Y=>nx5076, A=>nx5071);
   ix5739 : inv02 port map ( Y=>nx5077, A=>nx5229);
   ix5740 : inv02 port map ( Y=>nx5078, A=>nx4069);
   reg_nx1304 : ao22 port map ( Y=>nx1304, A0=>negative_M_10, A1=>nx4474, B0
      =>positive_M_10, B1=>nx4464);
   ix5741 : nor02_2x port map ( Y=>nx5079, A0=>nx4811, A1=>nx4817);
   reg_nx3640 : nor02_2x port map ( Y=>nx3640, A0=>nx5079, A1=>nx4945);
   ix5742 : inv01 port map ( Y=>nx5080, A=>nx2450);
   ix5743 : inv02 port map ( Y=>nx5081, A=>nx5241);
   ix5744 : or04 port map ( Y=>nx5082, A0=>nx5117, A1=>nx4605, A2=>nx5080, 
      A3=>nx5081);
   ix5745 : ao32 port map ( Y=>nx5083, A0=>nx4595, A1=>nx2450, A2=>nx4412, 
      B0=>nx4414, B1=>nx5152);
   ix5746 : inv02 port map ( Y=>nx5084, A=>nx4605);
   ix5747 : nand02_2x port map ( Y=>nx5085, A0=>nx5083, A1=>nx5084);
   ix5748 : or02 port map ( Y=>nx5086, A0=>nx4304, A1=>nx4195);
   reg_nx3388 : nand04_2x port map ( Y=>nx3388, A0=>nx5082, A1=>nx5085, A2=>
      nx5114, A3=>nx5086);
   ix5749 : inv01 port map ( Y=>nx5087, A=>nx5152);
   ix5750 : inv01 port map ( Y=>nx5088, A=>nx4412);
   ix5751 : inv01 port map ( Y=>nx5089, A=>nx4414);
   ix5752 : inv01 port map ( Y=>nx5090, A=>nx4595);
   ix5753 : nor02_2x port map ( Y=>nx5091, A0=>nx4414, A1=>nx4412);
   ix5754 : nor02_2x port map ( Y=>nx5092, A0=>nx4414, A1=>nx5241);
   ix5755 : aoi332 port map ( Y=>nx5093, A0=>nx5081, A1=>nx5089, A2=>nx5088, 
      B0=>nx5090, B1=>nx5087, B2=>nx5081, C0=>nx5090, C1=>nx5092);
   ix5756 : aoi322 port map ( Y=>nx5094, A0=>nx5087, A1=>nx5088, A2=>nx5081, 
      B0=>nx5087, B1=>nx5080, C0=>nx5089, C1=>nx5080);
   ix5757 : nand02_2x port map ( Y=>nx5095, A0=>nx5093, A1=>nx5094);
   reg_nx3783 : aoi221 port map ( Y=>nx3783, A0=>negative_M_11, A1=>nx4266, 
      B0=>positive_M_11, B1=>nx4278, C0=>nx1304);
   ix5758 : ao221 port map ( Y=>nx5096, A0=>nx4738, A1=>nx4850, B0=>nx5957, 
      B1=>nx4852, C0=>nx4853);
   ix5759 : aoi32 port map ( Y=>nx5097, A0=>nx4698, A1=>nx4376, A2=>nx4678, 
      B0=>nx4700, B1=>nx4807);
   ix5760 : nand02_2x port map ( Y=>nx5098, A0=>nx5096, A1=>nx5955);
   ix5761 : nand03_2x port map ( Y=>nx5099, A0=>nx4821, A1=>nx3640, A2=>
      nx5063);
   ix5762 : nand02_2x port map ( Y=>nx5100, A0=>nx4946, A1=>nx4947);
   ix5763 : nand03_2x port map ( Y=>nx5101, A0=>nx5099, A1=>nx4851, A2=>
      nx5100);
   ix5764 : aoi32 port map ( Y=>nx5102, A0=>nx4821, A1=>nx3640, A2=>nx5063, 
      B0=>nx4946, B1=>nx4947);
   ix5765 : inv02 port map ( Y=>nx5103, A=>nx5095);
   ix5766 : inv01 port map ( Y=>nx5104, A=>nx4628);
   ix5767 : or03 port map ( Y=>nx5105, A0=>nx5040, A1=>nx5937, A2=>nx4964);
   ix5768 : aoi22 port map ( Y=>nx5106, A0=>nx4966, A1=>nx5104, B0=>nx5105, 
      B1=>nx5104);
   ix5769 : nand02_2x port map ( Y=>nx5107, A0=>nx5103, A1=>nx5106);
   ix5770 : nand02_2x port map ( Y=>nx5108, A0=>nx5087, A1=>nx5088);
   ix5771 : inv02 port map ( Y=>nx5109, A=>nx5090);
   ix5772 : inv02 port map ( Y=>nx5110, A=>nx5087);
   ix5773 : inv02 port map ( Y=>nx5111, A=>nx5089);
   ix5774 : aoi22 port map ( Y=>nx5112, A0=>nx5108, A1=>nx5109, B0=>nx5110, 
      B1=>nx5111);
   ix5775 : or03 port map ( Y=>nx5113, A0=>nx5095, A1=>nx5112, A2=>nx5091);
   ix5776 : nand04_2x port map ( Y=>nx5114, A0=>nx5107, A1=>nx5113, A2=>
      nx4606, A3=>nx4607);
   ix5777 : inv01 port map ( Y=>nx5115, A=>nx4966);
   ix5778 : nor03_2x port map ( Y=>nx5116, A0=>nx5040, A1=>nx5937, A2=>
      nx4964);
   ix5779 : oai22 port map ( Y=>nx5117, A0=>nx5115, A1=>nx4628, B0=>nx5116, 
      B1=>nx4628);
   ix5780 : inv02 port map ( Y=>nx5118, A=>nx5229);
   ix5781 : inv02 port map ( Y=>nx5119, A=>nx4452);
   ix5782 : or03 port map ( Y=>nx5120, A0=>nx2150, A1=>nx5118, A2=>nx5119);
   ix5783 : and02 port map ( Y=>nx5121, A0=>nx5229, A1=>nx4452);
   ix5784 : aoi32 port map ( Y=>nx5122, A0=>nx4074, A1=>nx2150, A2=>nx5121, 
      B0=>nx5077, B1=>nx5078);
   reg_nx3328 : oai21 port map ( Y=>nx3328, A0=>nx4074, A1=>nx5120, B0=>
      nx5122);
   ix5785 : inv01 port map ( Y=>nx5123, A=>nx5237);
   ix5786 : nor02_2x port map ( Y=>nx5124, A0=>nx5237, A1=>nx5238);
   ix5787 : inv02 port map ( Y=>nx5125, A=>nx4989);
   ix5788 : nor02_2x port map ( Y=>nx5126, A0=>nx5125, A1=>nx5123);
   ix5789 : and02 port map ( Y=>nx5127, A0=>nx4132, A1=>nx5237);
   ix5790 : nor02_2x port map ( Y=>nx5128, A0=>nx5126, A1=>nx5127);
   ix5791 : nor02_2x port map ( Y=>nx5129, A0=>nx5051, A1=>nx4879);
   ix5792 : inv01 port map ( Y=>nx5130, A=>nx5239);
   ix5793 : nor02_2x port map ( Y=>nx5131, A0=>nx4132, A1=>nx4989);
   ix5794 : oai22 port map ( Y=>nx5132, A0=>nx5128, A1=>nx5129, B0=>nx5130, 
      B1=>nx5131);
   ix5795 : inv01 port map ( Y=>nx5133, A=>nx5123);
   ix5796 : oai22 port map ( Y=>nx5134, A0=>nx5133, A1=>nx5127, B0=>nx5051, 
      B1=>nx4879);
   ix5797 : oai21 port map ( Y=>nx5135, A0=>nx5239, A1=>nx5237, B0=>nx4132);
   ix5798 : aoi22 port map ( Y=>nx5136, A0=>nx5134, A1=>nx5130, B0=>nx5135, 
      B1=>nx5125);
   ix5799 : inv02 port map ( Y=>nx5137, A=>nx4132);
   ix5800 : aoi222 port map ( Y=>nx5138, A0=>nx5137, A1=>nx5125, B0=>nx5239, 
      B1=>nx5137, C0=>nx5130, C1=>nx5125);
   ix5801 : inv02 port map ( Y=>nx5139, A=>nx5138);
   ix5802 : inv01 port map ( Y=>nx5140, A=>nx5959);
   ix5803 : inv01 port map ( Y=>nx5141, A=>nx5959);
   ix5804 : inv01 port map ( Y=>nx5142, A=>nx5959);
   ix5805 : inv01 port map ( Y=>nx5143, A=>nx5149);
   ix5806 : inv02 port map ( Y=>nx5144, A=>nx5149);
   ix5807 : inv02 port map ( Y=>nx5145, A=>nx5149);
   ix5808 : inv01 port map ( Y=>nx5146, A=>nx5149);
   ix5809 : inv01 port map ( Y=>nx5147, A=>nx5149);
   ix5810 : inv01 port map ( Y=>nx5148, A=>nx5149);
   ix5811 : buf02 port map ( Y=>nx5149, A=>nx5180);
   ix5812 : inv02 port map ( Y=>nx5150, A=>nx4174);
   ix5813 : inv01 port map ( Y=>nx5151, A=>nx4414);
   ix5814 : oai22 port map ( Y=>nx5152, A0=>nx5150, A1=>nx5151, B0=>nx4174, 
      B1=>nx4414);
   reg_nx2450 : oai22 port map ( Y=>nx2450, A0=>nx5151, A1=>nx4174, B0=>
      nx5150, B1=>nx4414);
   reg_nx1786 : ao22 port map ( Y=>nx1786, A0=>negative_M_16, A1=>nx4476, B0
      =>positive_M_16, B1=>nx4466);
   ix5815 : ao21 port map ( Y=>nx5153, A0=>nx4708, A1=>nx4667, B0=>nx4668);
   reg_nx4116 : aoi321 port map ( Y=>nx4116, A0=>nx4666, A1=>nx4911, A2=>
      nx4667, B0=>nx4666, B1=>nx5153, C0=>nx5207);
   ix5816 : inv01 port map ( Y=>nx5154, A=>nx4116);
   ix5817 : oai32 port map ( Y=>nx5155, A0=>nx5207, A1=>nx4668, A2=>nx4667, 
      B0=>nx4666, B1=>nx5207);
   ix5818 : nor02_2x port map ( Y=>nx5156, A0=>nx5233, A1=>nx5227);
   ix5819 : and04 port map ( Y=>nx5157, A0=>nx5025, A1=>nx5235, A2=>nx2210, 
      A3=>nx5156);
   ix5820 : inv01 port map ( Y=>nx5158, A=>nx4053);
   ix5821 : inv02 port map ( Y=>nx5159, A=>nx2210);
   ix5822 : and03 port map ( Y=>nx5160, A0=>nx4635, A1=>nx5159, A2=>nx5156);
   reg_nx4302 : inv02 port map ( Y=>nx4302, A=>nx5227);
   ix5823 : and02 port map ( Y=>nx5161, A0=>nx5025, A1=>nx5235);
   ix5824 : nand03_2x port map ( Y=>nx5162, A0=>nx4635, A1=>nx5159, A2=>
      nx5156);
   ix5825 : oai422 port map ( Y=>nx5163, A0=>nx4635, A1=>nx5159, A2=>nx5233, 
      A3=>nx5227, B0=>nx5229, B1=>nx4090, C0=>nx5161, C1=>nx5162);
   reg_nx3338 : ao221 port map ( Y=>nx3338, A0=>nx4053, A1=>nx5157, B0=>
      nx5158, B1=>nx5160, C0=>nx5163);
   reg_nx4452 : inv02 port map ( Y=>nx4452, A=>nx5233);
   ix5826 : inv01 port map ( Y=>nx5164, A=>nx5125);
   ix5827 : inv01 port map ( Y=>nx5165, A=>nx5130);
   ix5828 : nand02_2x port map ( Y=>nx5166, A0=>nx5125, A1=>nx5239);
   ix5829 : inv02 port map ( Y=>nx5167, A=>nx5137);
   ix5830 : aoi22 port map ( Y=>nx5168, A0=>nx5164, A1=>nx5165, B0=>nx5166, 
      B1=>nx5167);
   ix5831 : nor02_2x port map ( Y=>nx5169, A0=>nx5961, A1=>nx4884);
   ix5832 : aoi21 port map ( Y=>nx5170, A0=>nx4623, A1=>nx5961, B0=>nx5124);
   ix5833 : nor02_2x port map ( Y=>nx5171, A0=>nx5169, A1=>nx5170);
   ix5834 : or02 port map ( Y=>nx5172, A0=>nx5137, A1=>nx5239);
   ix5835 : aoi221 port map ( Y=>nx5173, A0=>nx5125, A1=>nx5172, B0=>nx5130, 
      B1=>nx5137, C0=>nx4884);
   ix5836 : inv01 port map ( Y=>nx5174, A=>nx5173);
   ix5837 : inv01 port map ( Y=>nx5175, A=>nx5173);
   ix5838 : inv01 port map ( Y=>nx5176, A=>nx5173);
   ix5839 : inv01 port map ( Y=>nx5177, A=>nx5173);
   reg_nx2330 : inv01 port map ( Y=>nx2330, A=>nx5168);
   ix5840 : inv01 port map ( Y=>nx5178, A=>nx5961);
   ix5841 : inv01 port map ( Y=>nx5179, A=>nx5961);
   ix5842 : inv01 port map ( Y=>nx5180, A=>nx5961);
   reg_nx2086 : ao22 port map ( Y=>nx2086, A0=>negative_M_21, A1=>
      nx4478_XX0_XREP64, B0=>positive_M_21, B1=>nx4468);
   reg_nx4056 : aoi221 port map ( Y=>nx4056, A0=>positive_M_22, A1=>nx4282, 
      B0=>negative_M_22, B1=>nx4270, C0=>nx2086);
   ix5843 : inv02 port map ( Y=>nx5181, A=>nx3912);
   ix5844 : inv01 port map ( Y=>nx5182, A=>nx5911);
   ix5845 : aoi22 port map ( Y=>nx5183, A0=>nx5911, A1=>nx5181, B0=>nx3912, 
      B1=>nx5182);
   reg_nx1730 : inv01 port map ( Y=>nx1730, A=>nx5218);
   ix5846 : inv01 port map ( Y=>nx5184, A=>nx5219);
   ix5847 : inv01 port map ( Y=>nx5185, A=>nx5219);
   ix5848 : inv01 port map ( Y=>nx5186, A=>nx5219);
   ix5849 : inv01 port map ( Y=>nx5187, A=>nx5219);
   ix5850 : inv01 port map ( Y=>nx5188, A=>nx5219);
   ix5851 : inv01 port map ( Y=>nx5189, A=>nx5219);
   ix5852 : inv01 port map ( Y=>nx5190, A=>nx5062);
   ix5853 : inv01 port map ( Y=>nx5191, A=>nx4820);
   ix5854 : oai32 port map ( Y=>nx5192, A0=>nx5190, A1=>nx5191, A2=>nx4746, 
      B0=>nx4747, B1=>nx932);
   ix5855 : inv02 port map ( Y=>nx5193, A=>nx4788);
   ix5856 : ao22 port map ( Y=>nx5194, A0=>nx4280, A1=>positive_M_17, B0=>
      nx4268, B1=>negative_M_17);
   ix5857 : aoi22 port map ( Y=>nx5195, A0=>nx1786, A1=>nx5193, B0=>nx5194, 
      B1=>nx5193);
   ix5858 : inv01 port map ( Y=>nx5196, A=>nx5195);
   ix5859 : inv01 port map ( Y=>nx5197, A=>nx5195);
   ix5860 : and02 port map ( Y=>nx5198, A0=>nx4268, A1=>negative_M_17);
   ix5861 : and02 port map ( Y=>nx5199, A0=>nx4280, A1=>positive_M_17);
   ix5862 : nor03_2x port map ( Y=>nx5200, A0=>nx5198, A1=>nx5199, A2=>
      nx1786);
   ix5863 : ao21 port map ( Y=>nx5201, A0=>nx4673, A1=>nx4674, B0=>nx4672);
   ix5864 : nor02_2x port map ( Y=>nx5202, A0=>nx4671, A1=>nx4920);
   ix5865 : inv01 port map ( Y=>nx5203, A=>nx4657);
   ix5866 : nor04_2x port map ( Y=>nx5204, A0=>nx5202, A1=>nx5203, A2=>
      nx4708, A3=>nx4668);
   ix5867 : nand02_2x port map ( Y=>nx5205, A0=>nx5201, A1=>nx5204);
   ix5868 : oai22 port map ( Y=>nx5206, A0=>nx4672, A1=>nx4673, B0=>nx4672, 
      B1=>nx4674);
   ix5869 : oai21 port map ( Y=>nx5207, A0=>nx4671, A1=>nx4920, B0=>nx4657);
   ix5870 : buf16 port map ( Y=>nx5208, A=>nx4332);
   ix5871 : buf16 port map ( Y=>nx5209, A=>nx4332);
   ix5872 : buf16 port map ( Y=>nx5210, A=>nx602);
   ix5873 : buf16 port map ( Y=>nx5211, A=>nx602);
   ix5874 : buf16 port map ( Y=>nx5212, A=>nx4758);
   ix5875 : buf16 port map ( Y=>nx5213, A=>nx4758);
   ix5876 : buf16 port map ( Y=>nx5214, A=>nx4954);
   ix5877 : buf16 port map ( Y=>nx5215, A=>nx4954);
   ix5878 : buf16 port map ( Y=>nx5216, A=>nx4995);
   ix5879 : buf16 port map ( Y=>nx5217, A=>nx4995);
   ix5880 : buf16 port map ( Y=>nx5218, A=>nx5183);
   ix5881 : buf16 port map ( Y=>nx5219, A=>nx5183);
   ix5882 : buf16 port map ( Y=>nx5220, A=>nx5923);
   ix5883 : buf16 port map ( Y=>nx5221, A=>nx5923);
   ix5884 : buf16 port map ( Y=>nx5222, A=>nx4396);
   ix5885 : buf16 port map ( Y=>nx5223, A=>nx4396);
   ix5886 : buf16 port map ( Y=>nx5224, A=>nx4398);
   ix5887 : buf16 port map ( Y=>nx5225, A=>nx4398);
   ix5888 : buf16 port map ( Y=>nx5226, A=>nx4286);
   ix5889 : buf16 port map ( Y=>nx5227, A=>nx4286);
   ix5890 : buf16 port map ( Y=>nx5228, A=>nx4302);
   ix5891 : buf16 port map ( Y=>nx5229, A=>nx4302);
   ix5892 : buf16 port map ( Y=>nx5230, A=>nx4400);
   ix5893 : buf16 port map ( Y=>nx5231, A=>nx4400);
   ix5894 : buf16 port map ( Y=>nx5232, A=>nx4486);
   ix5895 : buf16 port map ( Y=>nx5233, A=>nx4486);
   ix5896 : buf16 port map ( Y=>nx5234, A=>nx2090);
   ix5897 : buf16 port map ( Y=>nx5235, A=>nx2090);
   ix5898 : buf16 port map ( Y=>nx5236, A=>nx4119);
   ix5899 : buf16 port map ( Y=>nx5237, A=>nx4119);
   ix5900 : buf16 port map ( Y=>nx5238, A=>nx4410);
   ix5901 : buf16 port map ( Y=>nx5239, A=>nx4410);
   ix5902 : buf16 port map ( Y=>nx5240, A=>nx2390);
   ix5903 : buf16 port map ( Y=>nx5241, A=>nx2390);
   ix5904 : inv02 port map ( Y=>nx5905, A=>nx4725);
   ix5906 : inv01 port map ( Y=>nx5907, A=>nx4742);
   ix5908 : inv01 port map ( Y=>nx5909, A=>nx4746);
   ix5910 : inv01 port map ( Y=>nx5911, A=>nx4699);
   ix5912 : buf02 port map ( Y=>nx5913, A=>nx4602);
   ix5914 : inv01 port map ( Y=>nx5915, A=>nx4691);
   ix5916 : buf02 port map ( Y=>nx5917, A=>nx4710);
   ix5918 : buf02 port map ( Y=>nx5919, A=>nx4731);
   ix5920 : buf02 port map ( Y=>nx5921, A=>nx3696);
   ix5922 : buf02 port map ( Y=>nx5923, A=>nx1850);
   ix5924 : buf02 port map ( Y=>nx5925, A=>nx4801);
   ix5926 : inv02 port map ( Y=>nx5927, A=>nx4877);
   ix5928 : inv02 port map ( Y=>nx5929, A=>nx4877);
   ix5930 : buf02 port map ( Y=>nx5931, A=>nx3972);
   ix5932 : inv01 port map ( Y=>nx5933, A=>nx4922);
   ix5934 : inv01 port map ( Y=>nx5935, A=>nx4733);
   ix5936 : buf02 port map ( Y=>nx5937, A=>nx4968);
   ix5938 : inv02 port map ( Y=>nx5939, A=>nx4837);
   ix5940 : inv01 port map ( Y=>nx5941, A=>nx4630);
   ix5942 : buf02 port map ( Y=>nx5943, A=>nx5001);
   ix5944 : inv02 port map ( Y=>nx5945, A=>nx1026);
   ix5946 : inv01 port map ( Y=>nx5947, A=>nx3699);
   ix5948 : inv01 port map ( Y=>nx5949, A=>nx4696);
   ix5950 : inv01 port map ( Y=>nx5951, A=>nx4695);
   ix5952 : inv01 port map ( Y=>nx5953, A=>nx4734);
   ix5954 : inv01 port map ( Y=>nx5955, A=>nx4776);
   ix5956 : inv01 port map ( Y=>nx5957, A=>nx3752);
   ix5958 : inv02 port map ( Y=>nx5959, A=>nx5139);
   ix5960 : inv01 port map ( Y=>nx5961, A=>nx2330);
   ix5970 : inv02 port map ( Y=>nx5971, A=>nx3851);
   ix5972 : inv02 port map ( Y=>nx5973, A=>nx3823);
   ix5974 : inv02 port map ( Y=>nx5975, A=>nx3823);
   ix5976 : inv02 port map ( Y=>nx5977, A=>nx3795);
   ix5978 : inv02 port map ( Y=>nx5979, A=>nx3795);
   ix5980 : inv02 port map ( Y=>nx5981, A=>nx3739);
   ix5982 : inv02 port map ( Y=>nx5983, A=>nx3739);
   ix5984 : inv02 port map ( Y=>nx5985, A=>nx3711);
   ix5986 : inv02 port map ( Y=>nx5987, A=>nx3711);
   ix5988 : inv02 port map ( Y=>nx5989, A=>nx3683);
   ix5990 : inv02 port map ( Y=>nx5991, A=>nx3655);
   ix5992 : inv02 port map ( Y=>nx5993, A=>nx3627);
   ix5994 : inv02 port map ( Y=>nx5995, A=>nx3597);
   ix5996 : buf02 port map ( Y=>nx5997, A=>M(3));
   ix5998 : buf02 port map ( Y=>nx5999, A=>M(2));
   ix6000 : buf02 port map ( Y=>nx6001, A=>M(2));
   ix6002 : inv02 port map ( Y=>nx6003, A=>nx4755);
   ix6004 : inv02 port map ( Y=>nx6005, A=>nx4755);
   ix6006 : buf02 port map ( Y=>nx6007, A=>M(0));
   ix6008 : buf02 port map ( Y=>nx6009, A=>M(0));
end ModifiedBoothMultiplierWorkFlow ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity NAdder_32_unfolded0 is
   port (
      a : IN std_logic_vector (31 DOWNTO 0) ;
      b : IN std_logic_vector (31 DOWNTO 0) ;
      cin : IN std_logic ;
      s : OUT std_logic_vector (31 DOWNTO 0) ;
      cout : OUT std_logic) ;
end NAdder_32_unfolded0 ;

architecture DataFlow_unfold_2009_1 of NAdder_32_unfolded0 is
   signal nx131, nx149, nx165, nx181, nx197, nx213, nx229, nx245, nx263, 
      nx275, nx287, nx331, nx340, nx341, nx342, nx343, nx344, nx345, nx346, 
      nx347, nx348, nx349, nx350, nx351, nx352, nx353, nx354, nx355, nx356, 
      nx357, nx358, nx359, nx360, nx361, nx362, nx363, nx364, nx365, nx366, 
      nx367, nx160, nx368, nx16, nx369, nx141, nx133, nx370, nx371, nx372, 
      nx373, nx374, s_27_EXMPLR, nx375, nx376, nx377, nx378, nx379, nx380, 
      nx329, nx381, nx382, nx383, nx384, nx385, nx386, nx387, nx311, nx388, 
      nx389, nx144, nx390, nx391, nx392, nx393, nx394, nx395, nx396, nx397, 
      nx398, nx399, nx400, nx401, nx402, nx403, nx404, nx327, nx405, nx406, 
      nx407, nx408, nx409, nx410, nx411, nx412, nx413, nx414, nx415, nx416, 
      nx417, nx329_XX0_XREP70, nx418, nx419, nx420, nx421, nx422, nx423, 
      nx424, nx425, nx128, nx426, nx427, nx249, nx255, nx112, nx237, nx428, 
      nx429, nx430, nx431, nx432, nx433, nx434, nx435, nx436, nx437, nx438, 
      nx439, nx440, nx441, nx266, nx442, nx443, nx444, nx445, nx446, nx447, 
      nx448, nx449, nx450, nx169, nx157, nx451, nx452, nx453, nx454, nx455, 
      nx456, nx457, nx458, nx459, nx460, nx461, nx462, nx233, nx463, nx464, 
      nx465, nx466, nx467, nx468, nx469, nx470, nx471, nx96, nx472, nx473, 
      nx474, nx475, nx476, nx477, nx478, nx201, nx205, nx479, nx480, nx481, 
      nx482, nx483, nx484, nx485, nx64, nx486, nx189, nx487, nx488, nx489, 
      nx490, nx491, nx492, nx493, nx494, nx495, nx185, nx496, nx173, nx497, 
      nx498, nx499, nx500, nx501, nx502, nx503, nx504, nx505, nx290, nx506, 
      nx507, nx508, nx509, nx510, nx511, nx512, nx513, nx514, nx515, nx299, 
      nx516, nx517, nx518, nx519, NOT_nx278, nx520, nx521, nx522, nx523, 
      nx524, nx525, nx526, nx527, nx528, nx529, nx530, nx531, nx32, nx532, 
      nx533, nx153, nx534, nx535, nx536, nx537, nx538, nx539, nx540, nx541, 
      nx542, nx543, nx544, nx545, nx546, nx547, nx548, nx549, nx550, nx551, 
      nx552, nx553, nx554, nx555, nx48, nx556, nx557, nx558, nx559, nx560, 
      nx561, nx562, nx563, nx564, nx565, nx566, NOT_nx302, nx567, nx568, 
      nx569, nx570, nx571, nx572, nx573, nx574, nx575, nx576, nx577, nx578, 
      nx579, nx580, nx581, nx582, nx583, nx584, nx585, nx586, nx587, nx588, 
      nx589, nx590, nx591, nx592, nx80, nx593, nx594, nx595, nx596, nx597, 
      nx598, nx137, nx599, nx600, nx601, nx602, nx603, nx604, nx605, nx606, 
      nx607, nx608, nx609, nx610, nx611, nx612, nx613, nx614, nx615, nx616, 
      nx617, nx618, nx619, nx620, nx621, nx622, nx623, nx909, nx911, nx913, 
      nx915, nx917, nx919, nx921, nx923, nx925, nx931, nx933, nx935, nx937, 
      nx939, nx941: std_logic ;

begin
   s(31) <= s_27_EXMPLR ;
   s(30) <= s_27_EXMPLR ;
   s(29) <= s_27_EXMPLR ;
   s(28) <= s_27_EXMPLR ;
   s(27) <= s_27_EXMPLR ;
   ix73 : fake_gnd port map ( Y=>cout);
   ix259 : xor2 port map ( Y=>s(0), A0=>a(0), A1=>b(0));
   ix257 : xor2 port map ( Y=>s(1), A0=>nx131, A1=>nx133);
   ix132 : nand02 port map ( Y=>nx131, A0=>b(0), A1=>a(0));
   ix255 : xor2 port map ( Y=>s(2), A0=>nx925, A1=>nx141);
   ix253 : xnor2 port map ( Y=>s(3), A0=>nx16, A1=>nx149);
   ix150 : xnor2_2x port map ( Y=>nx149, A0=>a(3), A1=>b(3));
   ix251 : xor2 port map ( Y=>s(4), A0=>nx153, A1=>nx157);
   ix249 : xnor2 port map ( Y=>s(5), A0=>nx32, A1=>nx165);
   ix166 : xnor2 port map ( Y=>nx165, A0=>a(5), A1=>b(5));
   ix247 : xor2 port map ( Y=>s(6), A0=>nx169, A1=>nx173);
   ix245 : xnor2 port map ( Y=>s(7), A0=>nx48, A1=>nx181);
   ix182 : xnor2 port map ( Y=>nx181, A0=>a(7), A1=>b(7));
   ix243 : xor2 port map ( Y=>s(8), A0=>nx185, A1=>nx189);
   ix241 : xnor2 port map ( Y=>s(9), A0=>nx64, A1=>nx197);
   ix198 : xnor2 port map ( Y=>nx197, A0=>a(9), A1=>b(9));
   ix239 : xor2 port map ( Y=>s(10), A0=>nx201, A1=>nx205);
   ix237 : xnor2 port map ( Y=>s(11), A0=>nx80, A1=>nx213);
   ix214 : xnor2 port map ( Y=>nx213, A0=>a(11), A1=>b(11));
   ix233 : xnor2 port map ( Y=>s(13), A0=>nx96, A1=>nx229);
   ix230 : xnor2 port map ( Y=>nx229, A0=>a(13), A1=>b(13));
   ix231 : xor2 port map ( Y=>s(14), A0=>nx233, A1=>nx237);
   ix229 : xnor2 port map ( Y=>s(15), A0=>nx112, A1=>nx245);
   ix246 : xnor2 port map ( Y=>nx245, A0=>a(15), A1=>nx935);
   ix227 : xor2 port map ( Y=>s(16), A0=>nx249, A1=>nx255);
   ix225 : xnor2 port map ( Y=>s(17), A0=>nx128, A1=>nx263);
   ix264 : xnor2 port map ( Y=>nx263, A0=>a(17), A1=>nx935);
   ix221 : xnor2 port map ( Y=>s(19), A0=>nx144, A1=>nx275);
   ix276 : xnor2 port map ( Y=>nx275, A0=>a(19), A1=>nx935);
   ix217 : xnor2 port map ( Y=>s(21), A0=>nx160, A1=>nx287);
   ix288 : xnor2 port map ( Y=>nx287, A0=>a(21), A1=>nx935);
   ix330 : inv02 port map ( Y=>nx331, A=>b(31));
   ix624 : aoi21 port map ( Y=>nx340, A0=>nx933, A1=>nx618, B0=>nx311);
   ix625 : nor03_2x port map ( Y=>nx341, A0=>nx340, A1=>nx620, A2=>nx931);
   ix626 : nand02_2x port map ( Y=>nx342, A0=>a(23), A1=>nx935);
   ix627 : inv02 port map ( Y=>nx343, A=>a(22));
   ix628 : oai21 port map ( Y=>nx344, A0=>a(23), A1=>a(22), B0=>nx935);
   ix629 : inv02 port map ( Y=>nx345, A=>a(24));
   ix630 : inv02 port map ( Y=>nx346, A=>a(25));
   ix631 : aoi22 port map ( Y=>nx347, A0=>nx620, A1=>nx618, B0=>nx345, B1=>
      nx346);
   ix632 : nand02_2x port map ( Y=>nx348, A0=>nx622, A1=>nx931);
   ix633 : aoi422 port map ( Y=>nx349, A0=>nx618, A1=>nx622, A2=>nx933, A3=>
      nx346, B0=>nx620, B1=>nx345, C0=>nx311, C1=>nx348);
   ix634 : oai22 port map ( Y=>nx350, A0=>nx622, A1=>nx345, B0=>nx620, B1=>
      nx933);
   ix635 : nor02_2x port map ( Y=>nx351, A0=>nx935, A1=>a(22));
   ix636 : inv02 port map ( Y=>nx352, A=>a(21));
   ix637 : inv02 port map ( Y=>nx353, A=>nx287);
   ix638 : nand02_2x port map ( Y=>nx354, A0=>a(20), A1=>nx353);
   ix639 : oai21 port map ( Y=>nx355, A0=>a(20), A1=>a(21), B0=>nx937);
   ix640 : aoi22 port map ( Y=>nx356, A0=>nx299, A1=>nx342, B0=>nx343, B1=>
      nx618);
   ix641 : inv02 port map ( Y=>nx357, A=>nx343);
   ix642 : nor02_2x port map ( Y=>nx358, A0=>nx357, A1=>nx937);
   ix643 : and02 port map ( Y=>nx359, A0=>nx516, A1=>nx342);
   ix644 : nor03_2x port map ( Y=>nx360, A0=>nx358, A1=>nx359, A2=>nx344);
   ix645 : inv02 port map ( Y=>nx361, A=>nx621);
   ix646 : inv02 port map ( Y=>nx362, A=>nx345);
   ix647 : inv02 port map ( Y=>nx363, A=>nx622);
   ix648 : inv02 port map ( Y=>nx364, A=>nx933);
   ix649 : aoi22 port map ( Y=>nx365, A0=>nx361, A1=>nx362, B0=>nx363, B1=>
      nx364);
   reg_s_24 : oai21 port map ( Y=>s(24), A0=>nx447, A1=>nx365, B0=>nx431);
   ix650 : nor02_2x port map ( Y=>nx366, A0=>nx937, A1=>a(20));
   ix651 : inv02 port map ( Y=>nx367, A=>a(20));
   reg_nx160 : oai22 port map ( Y=>nx160, A0=>nx366, A1=>NOT_nx278, B0=>
      nx618, B1=>nx367);
   ix652 : nand02_2x port map ( Y=>nx368, A0=>b(3), A1=>a(3));
   reg_nx16 : inv01 port map ( Y=>nx16, A=>nx451);
   ix653 : nor02_2x port map ( Y=>nx369, A0=>a(2), A1=>b(2));
   reg_nx141 : ao21 port map ( Y=>nx141, A0=>a(2), A1=>b(2), B0=>nx369);
   reg_nx133 : ao21 port map ( Y=>nx133, A0=>b(1), A1=>a(1), B0=>nx615);
   ix654 : inv02 port map ( Y=>nx370, A=>nx341);
   ix655 : nand02_2x port map ( Y=>nx371, A0=>nx618, A1=>nx354);
   ix656 : nand02_2x port map ( Y=>nx372, A0=>nx287, A1=>nx352);
   ix657 : nand03_2x port map ( Y=>nx373, A0=>nx371, A1=>nx356, A2=>nx372);
   ix658 : or03 port map ( Y=>nx374, A0=>nx931, A1=>nx933, A2=>nx621);
   s_31_EXMPLR : aoi22 port map ( Y=>s_27_EXMPLR, A0=>nx370, A1=>nx921, B0=>
      nx374, B1=>nx370);
   ix659 : aoi22 port map ( Y=>nx375, A0=>nx287, A1=>nx352, B0=>nx619, B1=>
      nx354);
   ix660 : inv02 port map ( Y=>nx376, A=>a(18));
   ix661 : inv02 port map ( Y=>nx377, A=>nx937);
   ix662 : aoi22 port map ( Y=>nx378, A0=>nx937, A1=>nx376, B0=>a(18), B1=>
      nx377);
   ix663 : nand02_2x port map ( Y=>nx379, A0=>nx937, A1=>a(19));
   ix664 : aoi21 port map ( Y=>nx380, A0=>nx355, A1=>nx379, B0=>nx373);
   reg_nx329 : inv02 port map ( Y=>nx329, A=>nx937);
   ix665 : nor04_2x port map ( Y=>nx381, A0=>nx373, A1=>nx275, A2=>nx619, A3
      =>nx376);
   ix666 : inv02 port map ( Y=>nx382, A=>nx350);
   ix667 : inv02 port map ( Y=>nx383, A=>nx931);
   ix668 : inv02 port map ( Y=>nx384, A=>nx623);
   ix669 : aoi22 port map ( Y=>nx385, A0=>nx931, A1=>nx623, B0=>nx383, B1=>
      nx384);
   ix670 : or02 port map ( Y=>nx386, A0=>nx382, A1=>nx385);
   ix671 : aoi222 port map ( Y=>nx387, A0=>nx931, A1=>nx623, B0=>nx383, B1=>
      nx384, C0=>nx933, C1=>nx939);
   reg_nx311 : oai22 port map ( Y=>nx311, A0=>nx383, A1=>nx384, B0=>nx931, 
      B1=>nx623);
   ix672 : and02 port map ( Y=>nx388, A0=>nx933, A1=>nx939);
   reg_s_25 : oai21 port map ( Y=>s(25), A0=>nx448, A1=>nx386, B0=>nx411);
   ix673 : and02 port map ( Y=>nx389, A0=>nx939, A1=>a(18));
   reg_nx144 : oai22 port map ( Y=>nx144, A0=>nx378, A1=>nx397, B0=>nx619, 
      B1=>nx376);
   ix674 : inv02 port map ( Y=>nx390, A=>nx263);
   ix675 : nor02_2x port map ( Y=>nx391, A0=>nx275, A1=>nx378);
   ix676 : nor02ii port map ( Y=>nx392, A0=>nx329_XX0_XREP70, A1=>a(17));
   ix677 : inv02 port map ( Y=>nx393, A=>nx275);
   ix678 : nand02_2x port map ( Y=>nx394, A0=>nx389, A1=>nx393);
   ix679 : nand02_2x port map ( Y=>nx395, A0=>nx379, A1=>nx394);
   ix680 : inv01 port map ( Y=>nx396, A=>nx375);
   ix681 : inv02 port map ( Y=>nx397, A=>nx442);
   ix682 : nor03_2x port map ( Y=>nx398, A0=>nx380, A1=>nx360, A2=>nx381);
   ix683 : inv02 port map ( Y=>nx399, A=>nx373);
   ix684 : inv01 port map ( Y=>nx400, A=>nx378);
   ix685 : inv02 port map ( Y=>nx401, A=>nx275);
   ix686 : nand03_2x port map ( Y=>nx402, A0=>nx399, A1=>nx400, A2=>nx401);
   ix687 : or02 port map ( Y=>nx403, A0=>nx621, A1=>nx347);
   ix688 : and02 port map ( Y=>nx404, A0=>nx621, A1=>nx349);
   reg_nx327 : inv02 port map ( Y=>nx327, A=>nx621);
   ix689 : inv02 port map ( Y=>nx405, A=>nx349);
   reg_s_26 : oai21 port map ( Y=>s(26), A0=>nx921, A1=>nx403, B0=>nx446);
   ix690 : inv02 port map ( Y=>nx406, A=>nx382);
   ix691 : inv02 port map ( Y=>nx407, A=>nx311);
   ix692 : inv02 port map ( Y=>nx408, A=>nx388);
   ix693 : aoi22 port map ( Y=>nx409, A0=>nx406, A1=>nx407, B0=>nx406, B1=>
      nx408);
   ix694 : ao21 port map ( Y=>nx410, A0=>nx311, A1=>nx388, B0=>nx387);
   ix695 : oai321 port map ( Y=>nx411, A0=>nx266, A1=>nx409, A2=>nx402, B0=>
      nx409, B1=>nx398, C0=>nx410);
   ix696 : nor02ii port map ( Y=>nx412, A0=>nx396, A1=>nx391);
   ix697 : inv02 port map ( Y=>nx413, A=>nx395);
   ix698 : nand02_2x port map ( Y=>nx414, A0=>nx355, A1=>nx413);
   ix699 : inv02 port map ( Y=>nx415, A=>nx396);
   ix700 : inv02 port map ( Y=>nx416, A=>a(15));
   ix701 : inv02 port map ( Y=>nx417, A=>a(16));
   reg_nx329_XX0_XREP70 : inv02 port map ( Y=>nx329_XX0_XREP70, A=>nx939);
   ix702 : aoi21 port map ( Y=>nx418, A0=>nx416, A1=>nx417, B0=>
      nx329_XX0_XREP70);
   ix703 : nor02_2x port map ( Y=>nx419, A0=>a(14), A1=>b(14));
   ix704 : and02 port map ( Y=>nx420, A0=>a(14), A1=>b(14));
   ix705 : nor02_2x port map ( Y=>nx421, A0=>nx939, A1=>a(16));
   ix706 : inv02 port map ( Y=>nx422, A=>nx390);
   ix707 : inv02 port map ( Y=>nx423, A=>nx391);
   ix708 : inv01 port map ( Y=>nx424, A=>nx392);
   ix709 : oai21 port map ( Y=>nx425, A0=>nx392, A1=>nx390, B0=>nx391);
   reg_nx128 : inv02 port map ( Y=>nx128, A=>nx527);
   ix710 : and02 port map ( Y=>nx426, A0=>a(15), A1=>nx939);
   ix711 : inv02 port map ( Y=>nx427, A=>nx245);
   reg_nx249 : oai32 port map ( Y=>nx249, A0=>nx426, A1=>nx462, A2=>nx420, 
      B0=>nx427, B1=>nx426);
   reg_nx255 : oai22 port map ( Y=>nx255, A0=>nx417, A1=>nx329_XX0_XREP70, 
      B0=>nx939, B1=>a(16));
   reg_nx112 : inv01 port map ( Y=>nx112, A=>nx459);
   reg_nx237 : ao21 port map ( Y=>nx237, A0=>a(14), A1=>b(14), B0=>nx419);
   ix712 : inv02 port map ( Y=>nx428, A=>nx390);
   ix713 : inv02 port map ( Y=>nx429, A=>nx392);
   ix714 : and02 port map ( Y=>nx430, A0=>nx365, A1=>nx398);
   ix715 : oai321 port map ( Y=>nx431, A0=>nx527, A1=>nx428, A2=>nx402, B0=>
      nx429, B1=>nx402, C0=>nx430);
   ix716 : inv01 port map ( Y=>nx432, A=>nx418);
   ix717 : aoi32 port map ( Y=>nx433, A0=>nx923, A1=>nx429, A2=>nx432, B0=>
      nx429, B1=>nx428);
   ix718 : oai22 port map ( Y=>nx434, A0=>nx376, A1=>nx377, B0=>a(18), B1=>
      nx941);
   ix719 : inv02 port map ( Y=>nx435, A=>nx376);
   ix720 : inv02 port map ( Y=>nx436, A=>nx377);
   ix721 : inv02 port map ( Y=>nx437, A=>a(18));
   ix722 : inv02 port map ( Y=>nx438, A=>nx941);
   ix723 : aoi22 port map ( Y=>nx439, A0=>nx435, A1=>nx436, B0=>nx437, B1=>
      nx438);
   ix724 : inv02 port map ( Y=>nx440, A=>nx429);
   ix725 : inv02 port map ( Y=>nx441, A=>nx428);
   reg_nx266 : oai32 port map ( Y=>nx266, A0=>nx482, A1=>nx440, A2=>nx909, 
      B0=>nx440, B1=>nx441);
   reg_s_18 : oai22 port map ( Y=>s(18), A0=>nx433, A1=>nx434, B0=>nx439, B1
      =>nx266);
   ix726 : ao221 port map ( Y=>nx442, A0=>nx909, A1=>nx441, B0=>nx483, B1=>
      nx441, C0=>nx440);
   ix727 : or02 port map ( Y=>nx443, A0=>nx428, A1=>nx402);
   ix728 : nor02_2x port map ( Y=>nx444, A0=>nx545, A1=>nx546);
   ix729 : and02 port map ( Y=>nx445, A0=>nx623, A1=>nx405);
   ix730 : oai32 port map ( Y=>nx446, A0=>nx921, A1=>nx445, A2=>nx347, B0=>
      nx445, B1=>nx404);
   ix731 : inv01 port map ( Y=>nx447, A=>NOT_nx302);
   ix732 : inv01 port map ( Y=>nx448, A=>nx921);
   ix733 : nand02_2x port map ( Y=>nx449, A0=>b(5), A1=>a(5));
   ix734 : nor02_2x port map ( Y=>nx450, A0=>a(4), A1=>b(4));
   reg_nx169 : inv02 port map ( Y=>nx169, A=>nx497);
   reg_nx157 : ao21 port map ( Y=>nx157, A0=>a(4), A1=>b(4), B0=>nx450);
   ix735 : aoi22 port map ( Y=>nx451, A0=>a(2), A1=>b(2), B0=>nx609, B1=>
      nx612);
   ix736 : inv01 port map ( Y=>nx452, A=>nx909);
   ix737 : inv02 port map ( Y=>nx453, A=>nx229);
   ix738 : nor03_2x port map ( Y=>nx454, A0=>nx419, A1=>nx421, A2=>nx245);
   ix739 : nor02_2x port map ( Y=>nx455, A0=>nx421, A1=>nx245);
   ix740 : and02 port map ( Y=>nx456, A0=>b(13), A1=>a(13));
   ix741 : nor02_2x port map ( Y=>nx457, A0=>nx453, A1=>nx911);
   ix742 : nor02_2x port map ( Y=>nx458, A0=>nx457, A1=>nx419);
   ix743 : oai32 port map ( Y=>nx459, A0=>nx472, A1=>nx911, A2=>nx420, B0=>
      nx458, B1=>nx420);
   ix744 : inv02 port map ( Y=>nx460, A=>nx419);
   ix745 : nor02_2x port map ( Y=>nx461, A0=>nx229, A1=>nx419);
   ix746 : ao22 port map ( Y=>nx462, A0=>nx460, A1=>nx911, B0=>nx473, B1=>
      nx461);
   reg_nx233 : oai22 port map ( Y=>nx233, A0=>nx911, A1=>nx474, B0=>nx453, 
      B1=>nx911);
   ix747 : or02 port map ( Y=>nx463, A0=>a(12), A1=>b(12));
   ix748 : or02 port map ( Y=>nx464, A0=>a(10), A1=>b(10));
   ix749 : and02 port map ( Y=>nx465, A0=>b(9), A1=>a(9));
   ix750 : nor02_2x port map ( Y=>nx466, A0=>a(10), A1=>b(10));
   ix751 : nor02_2x port map ( Y=>nx467, A0=>nx466, A1=>nx197);
   ix752 : nor02_2x port map ( Y=>nx468, A0=>a(12), A1=>b(12));
   ix753 : aoi21 port map ( Y=>nx469, A0=>nx420, A1=>nx455, B0=>nx911);
   ix754 : nand02_2x port map ( Y=>nx470, A0=>nx420, A1=>nx455);
   ix755 : oai21 port map ( Y=>nx471, A0=>nx453, A1=>nx911, B0=>nx454);
   reg_nx96 : inv01 port map ( Y=>nx96, A=>nx551);
   ix756 : inv01 port map ( Y=>nx472, A=>nx551);
   ix757 : inv01 port map ( Y=>nx473, A=>nx551);
   ix758 : inv01 port map ( Y=>nx474, A=>nx551);
   ix759 : nand02_2x port map ( Y=>nx475, A0=>b(11), A1=>a(11));
   ix760 : inv02 port map ( Y=>nx476, A=>nx213);
   ix761 : aoi21 port map ( Y=>nx477, A0=>b(11), A1=>a(11), B0=>nx476);
   ix762 : inv02 port map ( Y=>nx478, A=>nx197);
   reg_nx201 : oai22 port map ( Y=>nx201, A0=>nx465, A1=>nx486, B0=>nx478, 
      B1=>nx465);
   reg_nx205 : ao21 port map ( Y=>nx205, A0=>a(10), A1=>b(10), B0=>nx466);
   ix763 : or02 port map ( Y=>nx479, A0=>nx468, A1=>nx213);
   ix764 : nor02_2x port map ( Y=>nx480, A0=>a(8), A1=>b(8));
   ix765 : and02 port map ( Y=>nx481, A0=>nx470, A1=>nx471);
   ix766 : inv02 port map ( Y=>nx482, A=>nx597);
   ix767 : inv02 port map ( Y=>nx483, A=>nx923);
   ix768 : aoi22 port map ( Y=>nx484, A0=>a(10), A1=>b(10), B0=>nx464, B1=>
      nx465);
   ix769 : and02 port map ( Y=>nx485, A0=>a(8), A1=>b(8));
   reg_nx64 : inv01 port map ( Y=>nx64, A=>nx565);
   ix770 : inv01 port map ( Y=>nx486, A=>nx565);
   reg_nx189 : ao21 port map ( Y=>nx189, A0=>a(8), A1=>b(8), B0=>nx480);
   ix771 : inv02 port map ( Y=>nx487, A=>b(6));
   ix772 : nand02_2x port map ( Y=>nx488, A0=>nx449, A1=>nx487);
   ix773 : inv02 port map ( Y=>nx489, A=>nx449);
   ix774 : nor02_2x port map ( Y=>nx490, A0=>b(6), A1=>a(6));
   ix775 : nor02_2x port map ( Y=>nx491, A0=>nx490, A1=>nx165);
   ix776 : inv02 port map ( Y=>nx492, A=>nx181);
   ix777 : inv02 port map ( Y=>nx493, A=>nx468);
   ix778 : inv02 port map ( Y=>nx494, A=>nx213);
   ix779 : nand02_2x port map ( Y=>nx495, A0=>b(7), A1=>a(7));
   reg_nx185 : inv02 port map ( Y=>nx185, A=>nx595);
   ix780 : inv02 port map ( Y=>nx496, A=>a(6));
   reg_nx173 : oai22 port map ( Y=>nx173, A0=>nx496, A1=>nx487, B0=>b(6), B1
      =>a(6));
   ix781 : oai21 port map ( Y=>nx497, A0=>nx532, A1=>nx165, B0=>nx449);
   ix782 : inv02 port map ( Y=>nx498, A=>nx619);
   ix783 : inv02 port map ( Y=>nx499, A=>nx343);
   ix784 : inv02 port map ( Y=>nx500, A=>nx941);
   ix785 : inv02 port map ( Y=>nx501, A=>a(22));
   ix786 : aoi22 port map ( Y=>nx502, A0=>nx498, A1=>nx499, B0=>nx500, B1=>
      nx501);
   ix787 : nor02_2x port map ( Y=>nx503, A0=>nx290, A1=>nx502);
   reg_s_22 : ao21 port map ( Y=>s(22), A0=>nx290, A1=>nx502, B0=>nx503);
   ix788 : nand02_2x port map ( Y=>nx504, A0=>nx452, A1=>nx923);
   ix789 : nor03_2x port map ( Y=>nx505, A0=>nx423, A1=>nx422, A2=>nx396);
   reg_nx290 : aoi222 port map ( Y=>nx290, A0=>nx414, A1=>nx415, B0=>nx392, 
      B1=>nx412, C0=>nx504, C1=>nx505);
   ix790 : inv02 port map ( Y=>nx506, A=>nx619);
   ix791 : inv02 port map ( Y=>nx507, A=>nx343);
   ix792 : nand02_2x port map ( Y=>nx508, A0=>nx506, A1=>nx507);
   ix793 : inv02 port map ( Y=>nx509, A=>a(23));
   ix794 : inv02 port map ( Y=>nx510, A=>nx941);
   ix795 : aoi22 port map ( Y=>nx511, A0=>a(23), A1=>nx941, B0=>nx509, B1=>
      nx510);
   ix796 : nand03_2x port map ( Y=>nx512, A0=>nx290, A1=>nx508, A2=>nx917);
   ix797 : or03 port map ( Y=>nx513, A0=>nx290, A1=>nx917, A2=>nx351);
   ix798 : nand03_2x port map ( Y=>nx514, A0=>nx917, A1=>nx351, A2=>nx508);
   ix799 : or03 port map ( Y=>nx515, A0=>nx917, A1=>nx619, A2=>nx343);
   reg_s_23 : nand04_2x port map ( Y=>s(23), A0=>nx512, A1=>nx513, A2=>nx514, 
      A3=>nx515);
   reg_nx299 : inv01 port map ( Y=>nx299, A=>nx511);
   ix800 : inv01 port map ( Y=>nx516, A=>nx917);
   ix801 : inv02 port map ( Y=>nx517, A=>nx425);
   ix802 : ao21 port map ( Y=>nx518, A0=>nx424, A1=>nx452, B0=>nx425);
   ix803 : nand02_2x port map ( Y=>nx519, A0=>nx413, A1=>nx518);
   reg_NOT_nx278 : aoi21 port map ( Y=>NOT_nx278, A0=>nx547, A1=>nx517, B0=>
      nx519);
   ix804 : inv02 port map ( Y=>nx520, A=>nx941);
   ix805 : inv02 port map ( Y=>nx521, A=>a(20));
   ix806 : inv02 port map ( Y=>nx522, A=>nx619);
   ix807 : inv02 port map ( Y=>nx523, A=>nx367);
   ix808 : aoi22 port map ( Y=>nx524, A0=>nx520, A1=>nx521, B0=>nx522, B1=>
      nx523);
   ix809 : nand02_2x port map ( Y=>nx525, A0=>NOT_nx278, A1=>nx524);
   reg_s_20 : oai21 port map ( Y=>s(20), A0=>NOT_nx278, A1=>nx524, B0=>nx525
   );
   ix810 : inv02 port map ( Y=>nx526, A=>nx452);
   ix811 : nor02_2x port map ( Y=>nx527, A0=>nx526, A1=>nx548);
   ix812 : nand02_2x port map ( Y=>nx528, A0=>nx610, A1=>nx613);
   ix813 : inv02 port map ( Y=>nx529, A=>nx608);
   ix814 : inv02 port map ( Y=>nx530, A=>nx368);
   ix815 : nor02_2x port map ( Y=>nx531, A0=>nx530, A1=>nx617);
   reg_nx32 : aoi422 port map ( Y=>nx32, A0=>nx528, A1=>nx529, A2=>nx368, A3
      =>nx616, B0=>nx450, B1=>nx616, C0=>nx149, C1=>nx531);
   ix816 : inv02 port map ( Y=>nx532, A=>nx32);
   ix817 : inv02 port map ( Y=>nx533, A=>nx149);
   reg_nx153 : oai32 port map ( Y=>nx153, A0=>nx557, A1=>nx530, A2=>nx608, 
      B0=>nx533, B1=>nx530);
   ix818 : inv02 port map ( Y=>nx534, A=>nx481);
   ix819 : inv02 port map ( Y=>nx535, A=>nx463);
   ix820 : inv02 port map ( Y=>nx536, A=>b(11));
   ix821 : inv02 port map ( Y=>nx537, A=>a(11));
   ix822 : inv02 port map ( Y=>nx538, A=>a(12));
   ix823 : inv02 port map ( Y=>nx539, A=>b(12));
   ix824 : oai321 port map ( Y=>nx540, A0=>nx535, A1=>nx536, A2=>nx537, B0=>
      nx538, B1=>nx539, C0=>nx469);
   ix825 : inv02 port map ( Y=>nx541, A=>nx429);
   ix826 : inv02 port map ( Y=>nx542, A=>nx402);
   ix827 : nand02_2x port map ( Y=>nx543, A0=>nx541, A1=>nx542);
   ix828 : inv01 port map ( Y=>nx544, A=>nx909);
   ix829 : inv02 port map ( Y=>nx545, A=>nx398);
   ix830 : nor02_2x port map ( Y=>nx546, A0=>nx429, A1=>nx402);
   ix831 : inv02 port map ( Y=>nx547, A=>nx923);
   ix832 : inv02 port map ( Y=>nx548, A=>nx923);
   ix833 : and03 port map ( Y=>nx549, A0=>nx463, A1=>b(11), A2=>a(11));
   ix834 : and02 port map ( Y=>nx550, A0=>a(12), A1=>b(12));
   ix835 : nor03_2x port map ( Y=>nx551, A0=>nx549, A1=>nx550, A2=>nx554);
   ix836 : nand02_2x port map ( Y=>nx552, A0=>b(7), A1=>a(7));
   ix837 : inv02 port map ( Y=>nx553, A=>nx480);
   ix838 : inv01 port map ( Y=>nx554, A=>nx582);
   ix839 : inv02 port map ( Y=>nx555, A=>nx491);
   reg_nx48 : aoi22 port map ( Y=>nx48, A0=>nx555, A1=>nx567, B0=>nx606, B1
      =>nx567);
   ix840 : inv02 port map ( Y=>nx556, A=>nx48);
   ix841 : and02 port map ( Y=>nx557, A0=>nx611, A1=>nx614);
   ix842 : inv02 port map ( Y=>nx558, A=>nx571);
   ix843 : inv02 port map ( Y=>nx559, A=>nx484);
   ix844 : aoi21 port map ( Y=>nx560, A0=>a(12), A1=>b(12), B0=>nx468);
   ix845 : nand03_2x port map ( Y=>nx561, A0=>nx593, A1=>nx475, A2=>nx919);
   ix846 : inv02 port map ( Y=>nx562, A=>nx475);
   ix847 : nor02_2x port map ( Y=>nx563, A0=>nx919, A1=>nx913);
   ix848 : aoi22 port map ( Y=>nx564, A0=>nx562, A1=>nx563, B0=>nx913, B1=>
      nx919);
   reg_s_12 : nand03_2x port map ( Y=>s(12), A0=>nx561, A1=>nx589, A2=>nx564
   );
   ix849 : nor02_2x port map ( Y=>nx565, A0=>nx594, A1=>nx915);
   ix850 : and02 port map ( Y=>nx566, A0=>nx398, A1=>nx544);
   reg_NOT_nx302 : aoi32 port map ( Y=>NOT_nx302, A0=>nx566, A1=>nx923, A2=>
      nx543, B0=>nx443, B1=>nx444);
   ix851 : aoi22 port map ( Y=>nx567, A0=>a(6), A1=>nx488, B0=>b(6), B1=>
      nx489);
   ix852 : nand02_2x port map ( Y=>nx568, A0=>nx553, A1=>nx492);
   ix853 : oai22 port map ( Y=>nx569, A0=>nx480, A1=>nx552, B0=>nx567, B1=>
      nx568);
   ix854 : inv02 port map ( Y=>nx570, A=>nx479);
   ix855 : inv02 port map ( Y=>nx571, A=>nx467);
   ix856 : inv02 port map ( Y=>nx572, A=>a(8));
   ix857 : inv02 port map ( Y=>nx573, A=>b(8));
   ix858 : inv02 port map ( Y=>nx574, A=>a(10));
   ix859 : inv02 port map ( Y=>nx575, A=>b(10));
   ix860 : inv02 port map ( Y=>nx576, A=>nx464);
   ix861 : inv02 port map ( Y=>nx577, A=>nx465);
   ix862 : oai322 port map ( Y=>nx578, A0=>nx571, A1=>nx572, A2=>nx573, B0=>
      nx574, B1=>nx575, C0=>nx576, C1=>nx577);
   ix863 : nand02_2x port map ( Y=>nx579, A0=>nx491, A1=>nx467);
   ix864 : inv02 port map ( Y=>nx580, A=>nx492);
   ix865 : nor04_2x port map ( Y=>nx581, A0=>nx579, A1=>nx479, A2=>nx580, A3
      =>nx480);
   ix866 : aoi332 port map ( Y=>nx582, A0=>nx569, A1=>nx467, A2=>nx570, B0=>
      nx578, B1=>nx493, B2=>nx494, C0=>nx607, C1=>nx581);
   ix867 : nor02_2x port map ( Y=>nx583, A0=>nx559, A1=>nx915);
   ix868 : nand03_2x port map ( Y=>nx584, A0=>nx583, A1=>nx495, A2=>nx556);
   ix869 : aoi21 port map ( Y=>nx585, A0=>nx495, A1=>nx181, B0=>nx480);
   ix870 : nor03_2x port map ( Y=>nx586, A0=>nx585, A1=>nx559, A2=>nx915);
   ix871 : nor02_2x port map ( Y=>nx587, A0=>nx558, A1=>nx559);
   ix872 : nor04_2x port map ( Y=>nx588, A0=>nx586, A1=>nx587, A2=>nx919, A3
      =>nx913);
   ix873 : nand02_2x port map ( Y=>nx589, A0=>nx584, A1=>nx588);
   ix874 : inv02 port map ( Y=>nx590, A=>nx495);
   ix875 : inv01 port map ( Y=>nx591, A=>nx556);
   ix876 : nor04_2x port map ( Y=>nx592, A0=>nx559, A1=>nx915, A2=>nx590, A3
      =>nx591);
   reg_nx80 : nor03_2x port map ( Y=>nx80, A0=>nx592, A1=>nx586, A2=>nx587);
   ix877 : inv02 port map ( Y=>nx593, A=>nx80);
   ix878 : oai32 port map ( Y=>nx594, A0=>nx556, A1=>nx480, A2=>nx181, B0=>
      nx480, B1=>nx495);
   ix879 : oai21 port map ( Y=>nx595, A0=>nx181, A1=>nx556, B0=>nx495);
   ix880 : inv01 port map ( Y=>nx596, A=>nx582);
   ix881 : oai21 port map ( Y=>nx597, A0=>nx596, A1=>nx540, B0=>nx534);
   ix882 : or02 port map ( Y=>nx598, A0=>b(1), A1=>a(1));
   reg_nx137 : aoi32 port map ( Y=>nx137, A0=>nx598, A1=>b(0), A2=>a(0), B0
      =>b(1), B1=>a(1));
   ix883 : nor02_2x port map ( Y=>nx599, A0=>a(2), A1=>b(2));
   ix884 : nor04_2x port map ( Y=>nx600, A0=>nx925, A1=>nx599, A2=>nx450, A3
      =>nx149);
   ix885 : inv02 port map ( Y=>nx601, A=>a(2));
   ix886 : inv02 port map ( Y=>nx602, A=>b(2));
   ix887 : inv02 port map ( Y=>nx603, A=>a(4));
   ix888 : inv02 port map ( Y=>nx604, A=>b(4));
   ix889 : oai422 port map ( Y=>nx605, A0=>nx601, A1=>nx602, A2=>nx450, A3=>
      nx149, B0=>nx368, B1=>nx450, C0=>nx603, C1=>nx604);
   ix890 : nor02_2x port map ( Y=>nx606, A0=>nx600, A1=>nx605);
   ix891 : inv01 port map ( Y=>nx607, A=>nx606);
   ix892 : and02 port map ( Y=>nx608, A0=>a(2), A1=>b(2));
   ix893 : inv02 port map ( Y=>nx609, A=>nx599);
   ix894 : inv02 port map ( Y=>nx610, A=>nx599);
   ix895 : inv02 port map ( Y=>nx611, A=>nx599);
   ix896 : inv01 port map ( Y=>nx612, A=>nx137);
   ix897 : inv01 port map ( Y=>nx613, A=>nx925);
   ix898 : inv01 port map ( Y=>nx614, A=>nx925);
   ix899 : nor02_2x port map ( Y=>nx615, A0=>b(1), A1=>a(1));
   ix900 : nand02_2x port map ( Y=>nx616, A0=>a(4), A1=>b(4));
   ix901 : and02 port map ( Y=>nx617, A0=>a(4), A1=>b(4));
   ix902 : buf16 port map ( Y=>nx618, A=>nx329);
   ix903 : buf16 port map ( Y=>nx619, A=>nx329);
   ix904 : buf16 port map ( Y=>nx620, A=>nx331);
   ix905 : buf16 port map ( Y=>nx621, A=>nx331);
   ix906 : buf16 port map ( Y=>nx622, A=>nx327);
   ix907 : buf16 port map ( Y=>nx623, A=>nx327);
   ix908 : inv01 port map ( Y=>nx909, A=>nx432);
   ix910 : buf02 port map ( Y=>nx911, A=>nx456);
   ix912 : buf02 port map ( Y=>nx913, A=>nx477);
   ix914 : buf02 port map ( Y=>nx915, A=>nx485);
   ix916 : inv01 port map ( Y=>nx917, A=>nx299);
   ix918 : buf02 port map ( Y=>nx919, A=>nx560);
   ix920 : inv01 port map ( Y=>nx921, A=>nx447);
   ix922 : inv02 port map ( Y=>nx923, A=>nx482);
   ix924 : inv02 port map ( Y=>nx925, A=>nx612);
   ix930 : inv02 port map ( Y=>nx931, A=>nx346);
   ix932 : inv02 port map ( Y=>nx933, A=>nx345);
   ix934 : inv02 port map ( Y=>nx935, A=>nx331);
   ix936 : inv02 port map ( Y=>nx937, A=>nx331);
   ix938 : inv02 port map ( Y=>nx939, A=>nx331);
   ix940 : inv02 port map ( Y=>nx941, A=>nx331);
end DataFlow_unfold_2009_1 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity ComputationPipeline is
   port (
      img_data_0_15 : IN std_logic ;
      img_data_0_14 : IN std_logic ;
      img_data_0_13 : IN std_logic ;
      img_data_0_12 : IN std_logic ;
      img_data_0_11 : IN std_logic ;
      img_data_0_10 : IN std_logic ;
      img_data_0_9 : IN std_logic ;
      img_data_0_8 : IN std_logic ;
      img_data_0_7 : IN std_logic ;
      img_data_0_6 : IN std_logic ;
      img_data_0_5 : IN std_logic ;
      img_data_0_4 : IN std_logic ;
      img_data_0_3 : IN std_logic ;
      img_data_0_2 : IN std_logic ;
      img_data_0_1 : IN std_logic ;
      img_data_0_0 : IN std_logic ;
      img_data_1_15 : IN std_logic ;
      img_data_1_14 : IN std_logic ;
      img_data_1_13 : IN std_logic ;
      img_data_1_12 : IN std_logic ;
      img_data_1_11 : IN std_logic ;
      img_data_1_10 : IN std_logic ;
      img_data_1_9 : IN std_logic ;
      img_data_1_8 : IN std_logic ;
      img_data_1_7 : IN std_logic ;
      img_data_1_6 : IN std_logic ;
      img_data_1_5 : IN std_logic ;
      img_data_1_4 : IN std_logic ;
      img_data_1_3 : IN std_logic ;
      img_data_1_2 : IN std_logic ;
      img_data_1_1 : IN std_logic ;
      img_data_1_0 : IN std_logic ;
      img_data_2_15 : IN std_logic ;
      img_data_2_14 : IN std_logic ;
      img_data_2_13 : IN std_logic ;
      img_data_2_12 : IN std_logic ;
      img_data_2_11 : IN std_logic ;
      img_data_2_10 : IN std_logic ;
      img_data_2_9 : IN std_logic ;
      img_data_2_8 : IN std_logic ;
      img_data_2_7 : IN std_logic ;
      img_data_2_6 : IN std_logic ;
      img_data_2_5 : IN std_logic ;
      img_data_2_4 : IN std_logic ;
      img_data_2_3 : IN std_logic ;
      img_data_2_2 : IN std_logic ;
      img_data_2_1 : IN std_logic ;
      img_data_2_0 : IN std_logic ;
      img_data_3_15 : IN std_logic ;
      img_data_3_14 : IN std_logic ;
      img_data_3_13 : IN std_logic ;
      img_data_3_12 : IN std_logic ;
      img_data_3_11 : IN std_logic ;
      img_data_3_10 : IN std_logic ;
      img_data_3_9 : IN std_logic ;
      img_data_3_8 : IN std_logic ;
      img_data_3_7 : IN std_logic ;
      img_data_3_6 : IN std_logic ;
      img_data_3_5 : IN std_logic ;
      img_data_3_4 : IN std_logic ;
      img_data_3_3 : IN std_logic ;
      img_data_3_2 : IN std_logic ;
      img_data_3_1 : IN std_logic ;
      img_data_3_0 : IN std_logic ;
      img_data_4_15 : IN std_logic ;
      img_data_4_14 : IN std_logic ;
      img_data_4_13 : IN std_logic ;
      img_data_4_12 : IN std_logic ;
      img_data_4_11 : IN std_logic ;
      img_data_4_10 : IN std_logic ;
      img_data_4_9 : IN std_logic ;
      img_data_4_8 : IN std_logic ;
      img_data_4_7 : IN std_logic ;
      img_data_4_6 : IN std_logic ;
      img_data_4_5 : IN std_logic ;
      img_data_4_4 : IN std_logic ;
      img_data_4_3 : IN std_logic ;
      img_data_4_2 : IN std_logic ;
      img_data_4_1 : IN std_logic ;
      img_data_4_0 : IN std_logic ;
      img_data_5_15 : IN std_logic ;
      img_data_5_14 : IN std_logic ;
      img_data_5_13 : IN std_logic ;
      img_data_5_12 : IN std_logic ;
      img_data_5_11 : IN std_logic ;
      img_data_5_10 : IN std_logic ;
      img_data_5_9 : IN std_logic ;
      img_data_5_8 : IN std_logic ;
      img_data_5_7 : IN std_logic ;
      img_data_5_6 : IN std_logic ;
      img_data_5_5 : IN std_logic ;
      img_data_5_4 : IN std_logic ;
      img_data_5_3 : IN std_logic ;
      img_data_5_2 : IN std_logic ;
      img_data_5_1 : IN std_logic ;
      img_data_5_0 : IN std_logic ;
      img_data_6_15 : IN std_logic ;
      img_data_6_14 : IN std_logic ;
      img_data_6_13 : IN std_logic ;
      img_data_6_12 : IN std_logic ;
      img_data_6_11 : IN std_logic ;
      img_data_6_10 : IN std_logic ;
      img_data_6_9 : IN std_logic ;
      img_data_6_8 : IN std_logic ;
      img_data_6_7 : IN std_logic ;
      img_data_6_6 : IN std_logic ;
      img_data_6_5 : IN std_logic ;
      img_data_6_4 : IN std_logic ;
      img_data_6_3 : IN std_logic ;
      img_data_6_2 : IN std_logic ;
      img_data_6_1 : IN std_logic ;
      img_data_6_0 : IN std_logic ;
      img_data_7_15 : IN std_logic ;
      img_data_7_14 : IN std_logic ;
      img_data_7_13 : IN std_logic ;
      img_data_7_12 : IN std_logic ;
      img_data_7_11 : IN std_logic ;
      img_data_7_10 : IN std_logic ;
      img_data_7_9 : IN std_logic ;
      img_data_7_8 : IN std_logic ;
      img_data_7_7 : IN std_logic ;
      img_data_7_6 : IN std_logic ;
      img_data_7_5 : IN std_logic ;
      img_data_7_4 : IN std_logic ;
      img_data_7_3 : IN std_logic ;
      img_data_7_2 : IN std_logic ;
      img_data_7_1 : IN std_logic ;
      img_data_7_0 : IN std_logic ;
      img_data_8_15 : IN std_logic ;
      img_data_8_14 : IN std_logic ;
      img_data_8_13 : IN std_logic ;
      img_data_8_12 : IN std_logic ;
      img_data_8_11 : IN std_logic ;
      img_data_8_10 : IN std_logic ;
      img_data_8_9 : IN std_logic ;
      img_data_8_8 : IN std_logic ;
      img_data_8_7 : IN std_logic ;
      img_data_8_6 : IN std_logic ;
      img_data_8_5 : IN std_logic ;
      img_data_8_4 : IN std_logic ;
      img_data_8_3 : IN std_logic ;
      img_data_8_2 : IN std_logic ;
      img_data_8_1 : IN std_logic ;
      img_data_8_0 : IN std_logic ;
      img_data_9_15 : IN std_logic ;
      img_data_9_14 : IN std_logic ;
      img_data_9_13 : IN std_logic ;
      img_data_9_12 : IN std_logic ;
      img_data_9_11 : IN std_logic ;
      img_data_9_10 : IN std_logic ;
      img_data_9_9 : IN std_logic ;
      img_data_9_8 : IN std_logic ;
      img_data_9_7 : IN std_logic ;
      img_data_9_6 : IN std_logic ;
      img_data_9_5 : IN std_logic ;
      img_data_9_4 : IN std_logic ;
      img_data_9_3 : IN std_logic ;
      img_data_9_2 : IN std_logic ;
      img_data_9_1 : IN std_logic ;
      img_data_9_0 : IN std_logic ;
      img_data_10_15 : IN std_logic ;
      img_data_10_14 : IN std_logic ;
      img_data_10_13 : IN std_logic ;
      img_data_10_12 : IN std_logic ;
      img_data_10_11 : IN std_logic ;
      img_data_10_10 : IN std_logic ;
      img_data_10_9 : IN std_logic ;
      img_data_10_8 : IN std_logic ;
      img_data_10_7 : IN std_logic ;
      img_data_10_6 : IN std_logic ;
      img_data_10_5 : IN std_logic ;
      img_data_10_4 : IN std_logic ;
      img_data_10_3 : IN std_logic ;
      img_data_10_2 : IN std_logic ;
      img_data_10_1 : IN std_logic ;
      img_data_10_0 : IN std_logic ;
      img_data_11_15 : IN std_logic ;
      img_data_11_14 : IN std_logic ;
      img_data_11_13 : IN std_logic ;
      img_data_11_12 : IN std_logic ;
      img_data_11_11 : IN std_logic ;
      img_data_11_10 : IN std_logic ;
      img_data_11_9 : IN std_logic ;
      img_data_11_8 : IN std_logic ;
      img_data_11_7 : IN std_logic ;
      img_data_11_6 : IN std_logic ;
      img_data_11_5 : IN std_logic ;
      img_data_11_4 : IN std_logic ;
      img_data_11_3 : IN std_logic ;
      img_data_11_2 : IN std_logic ;
      img_data_11_1 : IN std_logic ;
      img_data_11_0 : IN std_logic ;
      img_data_12_15 : IN std_logic ;
      img_data_12_14 : IN std_logic ;
      img_data_12_13 : IN std_logic ;
      img_data_12_12 : IN std_logic ;
      img_data_12_11 : IN std_logic ;
      img_data_12_10 : IN std_logic ;
      img_data_12_9 : IN std_logic ;
      img_data_12_8 : IN std_logic ;
      img_data_12_7 : IN std_logic ;
      img_data_12_6 : IN std_logic ;
      img_data_12_5 : IN std_logic ;
      img_data_12_4 : IN std_logic ;
      img_data_12_3 : IN std_logic ;
      img_data_12_2 : IN std_logic ;
      img_data_12_1 : IN std_logic ;
      img_data_12_0 : IN std_logic ;
      img_data_13_15 : IN std_logic ;
      img_data_13_14 : IN std_logic ;
      img_data_13_13 : IN std_logic ;
      img_data_13_12 : IN std_logic ;
      img_data_13_11 : IN std_logic ;
      img_data_13_10 : IN std_logic ;
      img_data_13_9 : IN std_logic ;
      img_data_13_8 : IN std_logic ;
      img_data_13_7 : IN std_logic ;
      img_data_13_6 : IN std_logic ;
      img_data_13_5 : IN std_logic ;
      img_data_13_4 : IN std_logic ;
      img_data_13_3 : IN std_logic ;
      img_data_13_2 : IN std_logic ;
      img_data_13_1 : IN std_logic ;
      img_data_13_0 : IN std_logic ;
      img_data_14_15 : IN std_logic ;
      img_data_14_14 : IN std_logic ;
      img_data_14_13 : IN std_logic ;
      img_data_14_12 : IN std_logic ;
      img_data_14_11 : IN std_logic ;
      img_data_14_10 : IN std_logic ;
      img_data_14_9 : IN std_logic ;
      img_data_14_8 : IN std_logic ;
      img_data_14_7 : IN std_logic ;
      img_data_14_6 : IN std_logic ;
      img_data_14_5 : IN std_logic ;
      img_data_14_4 : IN std_logic ;
      img_data_14_3 : IN std_logic ;
      img_data_14_2 : IN std_logic ;
      img_data_14_1 : IN std_logic ;
      img_data_14_0 : IN std_logic ;
      img_data_15_15 : IN std_logic ;
      img_data_15_14 : IN std_logic ;
      img_data_15_13 : IN std_logic ;
      img_data_15_12 : IN std_logic ;
      img_data_15_11 : IN std_logic ;
      img_data_15_10 : IN std_logic ;
      img_data_15_9 : IN std_logic ;
      img_data_15_8 : IN std_logic ;
      img_data_15_7 : IN std_logic ;
      img_data_15_6 : IN std_logic ;
      img_data_15_5 : IN std_logic ;
      img_data_15_4 : IN std_logic ;
      img_data_15_3 : IN std_logic ;
      img_data_15_2 : IN std_logic ;
      img_data_15_1 : IN std_logic ;
      img_data_15_0 : IN std_logic ;
      img_data_16_15 : IN std_logic ;
      img_data_16_14 : IN std_logic ;
      img_data_16_13 : IN std_logic ;
      img_data_16_12 : IN std_logic ;
      img_data_16_11 : IN std_logic ;
      img_data_16_10 : IN std_logic ;
      img_data_16_9 : IN std_logic ;
      img_data_16_8 : IN std_logic ;
      img_data_16_7 : IN std_logic ;
      img_data_16_6 : IN std_logic ;
      img_data_16_5 : IN std_logic ;
      img_data_16_4 : IN std_logic ;
      img_data_16_3 : IN std_logic ;
      img_data_16_2 : IN std_logic ;
      img_data_16_1 : IN std_logic ;
      img_data_16_0 : IN std_logic ;
      img_data_17_15 : IN std_logic ;
      img_data_17_14 : IN std_logic ;
      img_data_17_13 : IN std_logic ;
      img_data_17_12 : IN std_logic ;
      img_data_17_11 : IN std_logic ;
      img_data_17_10 : IN std_logic ;
      img_data_17_9 : IN std_logic ;
      img_data_17_8 : IN std_logic ;
      img_data_17_7 : IN std_logic ;
      img_data_17_6 : IN std_logic ;
      img_data_17_5 : IN std_logic ;
      img_data_17_4 : IN std_logic ;
      img_data_17_3 : IN std_logic ;
      img_data_17_2 : IN std_logic ;
      img_data_17_1 : IN std_logic ;
      img_data_17_0 : IN std_logic ;
      img_data_18_15 : IN std_logic ;
      img_data_18_14 : IN std_logic ;
      img_data_18_13 : IN std_logic ;
      img_data_18_12 : IN std_logic ;
      img_data_18_11 : IN std_logic ;
      img_data_18_10 : IN std_logic ;
      img_data_18_9 : IN std_logic ;
      img_data_18_8 : IN std_logic ;
      img_data_18_7 : IN std_logic ;
      img_data_18_6 : IN std_logic ;
      img_data_18_5 : IN std_logic ;
      img_data_18_4 : IN std_logic ;
      img_data_18_3 : IN std_logic ;
      img_data_18_2 : IN std_logic ;
      img_data_18_1 : IN std_logic ;
      img_data_18_0 : IN std_logic ;
      img_data_19_15 : IN std_logic ;
      img_data_19_14 : IN std_logic ;
      img_data_19_13 : IN std_logic ;
      img_data_19_12 : IN std_logic ;
      img_data_19_11 : IN std_logic ;
      img_data_19_10 : IN std_logic ;
      img_data_19_9 : IN std_logic ;
      img_data_19_8 : IN std_logic ;
      img_data_19_7 : IN std_logic ;
      img_data_19_6 : IN std_logic ;
      img_data_19_5 : IN std_logic ;
      img_data_19_4 : IN std_logic ;
      img_data_19_3 : IN std_logic ;
      img_data_19_2 : IN std_logic ;
      img_data_19_1 : IN std_logic ;
      img_data_19_0 : IN std_logic ;
      img_data_20_15 : IN std_logic ;
      img_data_20_14 : IN std_logic ;
      img_data_20_13 : IN std_logic ;
      img_data_20_12 : IN std_logic ;
      img_data_20_11 : IN std_logic ;
      img_data_20_10 : IN std_logic ;
      img_data_20_9 : IN std_logic ;
      img_data_20_8 : IN std_logic ;
      img_data_20_7 : IN std_logic ;
      img_data_20_6 : IN std_logic ;
      img_data_20_5 : IN std_logic ;
      img_data_20_4 : IN std_logic ;
      img_data_20_3 : IN std_logic ;
      img_data_20_2 : IN std_logic ;
      img_data_20_1 : IN std_logic ;
      img_data_20_0 : IN std_logic ;
      img_data_21_15 : IN std_logic ;
      img_data_21_14 : IN std_logic ;
      img_data_21_13 : IN std_logic ;
      img_data_21_12 : IN std_logic ;
      img_data_21_11 : IN std_logic ;
      img_data_21_10 : IN std_logic ;
      img_data_21_9 : IN std_logic ;
      img_data_21_8 : IN std_logic ;
      img_data_21_7 : IN std_logic ;
      img_data_21_6 : IN std_logic ;
      img_data_21_5 : IN std_logic ;
      img_data_21_4 : IN std_logic ;
      img_data_21_3 : IN std_logic ;
      img_data_21_2 : IN std_logic ;
      img_data_21_1 : IN std_logic ;
      img_data_21_0 : IN std_logic ;
      img_data_22_15 : IN std_logic ;
      img_data_22_14 : IN std_logic ;
      img_data_22_13 : IN std_logic ;
      img_data_22_12 : IN std_logic ;
      img_data_22_11 : IN std_logic ;
      img_data_22_10 : IN std_logic ;
      img_data_22_9 : IN std_logic ;
      img_data_22_8 : IN std_logic ;
      img_data_22_7 : IN std_logic ;
      img_data_22_6 : IN std_logic ;
      img_data_22_5 : IN std_logic ;
      img_data_22_4 : IN std_logic ;
      img_data_22_3 : IN std_logic ;
      img_data_22_2 : IN std_logic ;
      img_data_22_1 : IN std_logic ;
      img_data_22_0 : IN std_logic ;
      img_data_23_15 : IN std_logic ;
      img_data_23_14 : IN std_logic ;
      img_data_23_13 : IN std_logic ;
      img_data_23_12 : IN std_logic ;
      img_data_23_11 : IN std_logic ;
      img_data_23_10 : IN std_logic ;
      img_data_23_9 : IN std_logic ;
      img_data_23_8 : IN std_logic ;
      img_data_23_7 : IN std_logic ;
      img_data_23_6 : IN std_logic ;
      img_data_23_5 : IN std_logic ;
      img_data_23_4 : IN std_logic ;
      img_data_23_3 : IN std_logic ;
      img_data_23_2 : IN std_logic ;
      img_data_23_1 : IN std_logic ;
      img_data_23_0 : IN std_logic ;
      img_data_24_15 : IN std_logic ;
      img_data_24_14 : IN std_logic ;
      img_data_24_13 : IN std_logic ;
      img_data_24_12 : IN std_logic ;
      img_data_24_11 : IN std_logic ;
      img_data_24_10 : IN std_logic ;
      img_data_24_9 : IN std_logic ;
      img_data_24_8 : IN std_logic ;
      img_data_24_7 : IN std_logic ;
      img_data_24_6 : IN std_logic ;
      img_data_24_5 : IN std_logic ;
      img_data_24_4 : IN std_logic ;
      img_data_24_3 : IN std_logic ;
      img_data_24_2 : IN std_logic ;
      img_data_24_1 : IN std_logic ;
      img_data_24_0 : IN std_logic ;
      filter_data_0_15 : IN std_logic ;
      filter_data_0_14 : IN std_logic ;
      filter_data_0_13 : IN std_logic ;
      filter_data_0_12 : IN std_logic ;
      filter_data_0_11 : IN std_logic ;
      filter_data_0_10 : IN std_logic ;
      filter_data_0_9 : IN std_logic ;
      filter_data_0_8 : IN std_logic ;
      filter_data_0_7 : IN std_logic ;
      filter_data_0_6 : IN std_logic ;
      filter_data_0_5 : IN std_logic ;
      filter_data_0_4 : IN std_logic ;
      filter_data_0_3 : IN std_logic ;
      filter_data_0_2 : IN std_logic ;
      filter_data_0_1 : IN std_logic ;
      filter_data_0_0 : IN std_logic ;
      filter_data_1_15 : IN std_logic ;
      filter_data_1_14 : IN std_logic ;
      filter_data_1_13 : IN std_logic ;
      filter_data_1_12 : IN std_logic ;
      filter_data_1_11 : IN std_logic ;
      filter_data_1_10 : IN std_logic ;
      filter_data_1_9 : IN std_logic ;
      filter_data_1_8 : IN std_logic ;
      filter_data_1_7 : IN std_logic ;
      filter_data_1_6 : IN std_logic ;
      filter_data_1_5 : IN std_logic ;
      filter_data_1_4 : IN std_logic ;
      filter_data_1_3 : IN std_logic ;
      filter_data_1_2 : IN std_logic ;
      filter_data_1_1 : IN std_logic ;
      filter_data_1_0 : IN std_logic ;
      filter_data_2_15 : IN std_logic ;
      filter_data_2_14 : IN std_logic ;
      filter_data_2_13 : IN std_logic ;
      filter_data_2_12 : IN std_logic ;
      filter_data_2_11 : IN std_logic ;
      filter_data_2_10 : IN std_logic ;
      filter_data_2_9 : IN std_logic ;
      filter_data_2_8 : IN std_logic ;
      filter_data_2_7 : IN std_logic ;
      filter_data_2_6 : IN std_logic ;
      filter_data_2_5 : IN std_logic ;
      filter_data_2_4 : IN std_logic ;
      filter_data_2_3 : IN std_logic ;
      filter_data_2_2 : IN std_logic ;
      filter_data_2_1 : IN std_logic ;
      filter_data_2_0 : IN std_logic ;
      filter_data_3_15 : IN std_logic ;
      filter_data_3_14 : IN std_logic ;
      filter_data_3_13 : IN std_logic ;
      filter_data_3_12 : IN std_logic ;
      filter_data_3_11 : IN std_logic ;
      filter_data_3_10 : IN std_logic ;
      filter_data_3_9 : IN std_logic ;
      filter_data_3_8 : IN std_logic ;
      filter_data_3_7 : IN std_logic ;
      filter_data_3_6 : IN std_logic ;
      filter_data_3_5 : IN std_logic ;
      filter_data_3_4 : IN std_logic ;
      filter_data_3_3 : IN std_logic ;
      filter_data_3_2 : IN std_logic ;
      filter_data_3_1 : IN std_logic ;
      filter_data_3_0 : IN std_logic ;
      filter_data_4_15 : IN std_logic ;
      filter_data_4_14 : IN std_logic ;
      filter_data_4_13 : IN std_logic ;
      filter_data_4_12 : IN std_logic ;
      filter_data_4_11 : IN std_logic ;
      filter_data_4_10 : IN std_logic ;
      filter_data_4_9 : IN std_logic ;
      filter_data_4_8 : IN std_logic ;
      filter_data_4_7 : IN std_logic ;
      filter_data_4_6 : IN std_logic ;
      filter_data_4_5 : IN std_logic ;
      filter_data_4_4 : IN std_logic ;
      filter_data_4_3 : IN std_logic ;
      filter_data_4_2 : IN std_logic ;
      filter_data_4_1 : IN std_logic ;
      filter_data_4_0 : IN std_logic ;
      filter_data_5_15 : IN std_logic ;
      filter_data_5_14 : IN std_logic ;
      filter_data_5_13 : IN std_logic ;
      filter_data_5_12 : IN std_logic ;
      filter_data_5_11 : IN std_logic ;
      filter_data_5_10 : IN std_logic ;
      filter_data_5_9 : IN std_logic ;
      filter_data_5_8 : IN std_logic ;
      filter_data_5_7 : IN std_logic ;
      filter_data_5_6 : IN std_logic ;
      filter_data_5_5 : IN std_logic ;
      filter_data_5_4 : IN std_logic ;
      filter_data_5_3 : IN std_logic ;
      filter_data_5_2 : IN std_logic ;
      filter_data_5_1 : IN std_logic ;
      filter_data_5_0 : IN std_logic ;
      filter_data_6_15 : IN std_logic ;
      filter_data_6_14 : IN std_logic ;
      filter_data_6_13 : IN std_logic ;
      filter_data_6_12 : IN std_logic ;
      filter_data_6_11 : IN std_logic ;
      filter_data_6_10 : IN std_logic ;
      filter_data_6_9 : IN std_logic ;
      filter_data_6_8 : IN std_logic ;
      filter_data_6_7 : IN std_logic ;
      filter_data_6_6 : IN std_logic ;
      filter_data_6_5 : IN std_logic ;
      filter_data_6_4 : IN std_logic ;
      filter_data_6_3 : IN std_logic ;
      filter_data_6_2 : IN std_logic ;
      filter_data_6_1 : IN std_logic ;
      filter_data_6_0 : IN std_logic ;
      filter_data_7_15 : IN std_logic ;
      filter_data_7_14 : IN std_logic ;
      filter_data_7_13 : IN std_logic ;
      filter_data_7_12 : IN std_logic ;
      filter_data_7_11 : IN std_logic ;
      filter_data_7_10 : IN std_logic ;
      filter_data_7_9 : IN std_logic ;
      filter_data_7_8 : IN std_logic ;
      filter_data_7_7 : IN std_logic ;
      filter_data_7_6 : IN std_logic ;
      filter_data_7_5 : IN std_logic ;
      filter_data_7_4 : IN std_logic ;
      filter_data_7_3 : IN std_logic ;
      filter_data_7_2 : IN std_logic ;
      filter_data_7_1 : IN std_logic ;
      filter_data_7_0 : IN std_logic ;
      filter_data_8_15 : IN std_logic ;
      filter_data_8_14 : IN std_logic ;
      filter_data_8_13 : IN std_logic ;
      filter_data_8_12 : IN std_logic ;
      filter_data_8_11 : IN std_logic ;
      filter_data_8_10 : IN std_logic ;
      filter_data_8_9 : IN std_logic ;
      filter_data_8_8 : IN std_logic ;
      filter_data_8_7 : IN std_logic ;
      filter_data_8_6 : IN std_logic ;
      filter_data_8_5 : IN std_logic ;
      filter_data_8_4 : IN std_logic ;
      filter_data_8_3 : IN std_logic ;
      filter_data_8_2 : IN std_logic ;
      filter_data_8_1 : IN std_logic ;
      filter_data_8_0 : IN std_logic ;
      filter_data_9_15 : IN std_logic ;
      filter_data_9_14 : IN std_logic ;
      filter_data_9_13 : IN std_logic ;
      filter_data_9_12 : IN std_logic ;
      filter_data_9_11 : IN std_logic ;
      filter_data_9_10 : IN std_logic ;
      filter_data_9_9 : IN std_logic ;
      filter_data_9_8 : IN std_logic ;
      filter_data_9_7 : IN std_logic ;
      filter_data_9_6 : IN std_logic ;
      filter_data_9_5 : IN std_logic ;
      filter_data_9_4 : IN std_logic ;
      filter_data_9_3 : IN std_logic ;
      filter_data_9_2 : IN std_logic ;
      filter_data_9_1 : IN std_logic ;
      filter_data_9_0 : IN std_logic ;
      filter_data_10_15 : IN std_logic ;
      filter_data_10_14 : IN std_logic ;
      filter_data_10_13 : IN std_logic ;
      filter_data_10_12 : IN std_logic ;
      filter_data_10_11 : IN std_logic ;
      filter_data_10_10 : IN std_logic ;
      filter_data_10_9 : IN std_logic ;
      filter_data_10_8 : IN std_logic ;
      filter_data_10_7 : IN std_logic ;
      filter_data_10_6 : IN std_logic ;
      filter_data_10_5 : IN std_logic ;
      filter_data_10_4 : IN std_logic ;
      filter_data_10_3 : IN std_logic ;
      filter_data_10_2 : IN std_logic ;
      filter_data_10_1 : IN std_logic ;
      filter_data_10_0 : IN std_logic ;
      filter_data_11_15 : IN std_logic ;
      filter_data_11_14 : IN std_logic ;
      filter_data_11_13 : IN std_logic ;
      filter_data_11_12 : IN std_logic ;
      filter_data_11_11 : IN std_logic ;
      filter_data_11_10 : IN std_logic ;
      filter_data_11_9 : IN std_logic ;
      filter_data_11_8 : IN std_logic ;
      filter_data_11_7 : IN std_logic ;
      filter_data_11_6 : IN std_logic ;
      filter_data_11_5 : IN std_logic ;
      filter_data_11_4 : IN std_logic ;
      filter_data_11_3 : IN std_logic ;
      filter_data_11_2 : IN std_logic ;
      filter_data_11_1 : IN std_logic ;
      filter_data_11_0 : IN std_logic ;
      filter_data_12_15 : IN std_logic ;
      filter_data_12_14 : IN std_logic ;
      filter_data_12_13 : IN std_logic ;
      filter_data_12_12 : IN std_logic ;
      filter_data_12_11 : IN std_logic ;
      filter_data_12_10 : IN std_logic ;
      filter_data_12_9 : IN std_logic ;
      filter_data_12_8 : IN std_logic ;
      filter_data_12_7 : IN std_logic ;
      filter_data_12_6 : IN std_logic ;
      filter_data_12_5 : IN std_logic ;
      filter_data_12_4 : IN std_logic ;
      filter_data_12_3 : IN std_logic ;
      filter_data_12_2 : IN std_logic ;
      filter_data_12_1 : IN std_logic ;
      filter_data_12_0 : IN std_logic ;
      filter_data_13_15 : IN std_logic ;
      filter_data_13_14 : IN std_logic ;
      filter_data_13_13 : IN std_logic ;
      filter_data_13_12 : IN std_logic ;
      filter_data_13_11 : IN std_logic ;
      filter_data_13_10 : IN std_logic ;
      filter_data_13_9 : IN std_logic ;
      filter_data_13_8 : IN std_logic ;
      filter_data_13_7 : IN std_logic ;
      filter_data_13_6 : IN std_logic ;
      filter_data_13_5 : IN std_logic ;
      filter_data_13_4 : IN std_logic ;
      filter_data_13_3 : IN std_logic ;
      filter_data_13_2 : IN std_logic ;
      filter_data_13_1 : IN std_logic ;
      filter_data_13_0 : IN std_logic ;
      filter_data_14_15 : IN std_logic ;
      filter_data_14_14 : IN std_logic ;
      filter_data_14_13 : IN std_logic ;
      filter_data_14_12 : IN std_logic ;
      filter_data_14_11 : IN std_logic ;
      filter_data_14_10 : IN std_logic ;
      filter_data_14_9 : IN std_logic ;
      filter_data_14_8 : IN std_logic ;
      filter_data_14_7 : IN std_logic ;
      filter_data_14_6 : IN std_logic ;
      filter_data_14_5 : IN std_logic ;
      filter_data_14_4 : IN std_logic ;
      filter_data_14_3 : IN std_logic ;
      filter_data_14_2 : IN std_logic ;
      filter_data_14_1 : IN std_logic ;
      filter_data_14_0 : IN std_logic ;
      filter_data_15_15 : IN std_logic ;
      filter_data_15_14 : IN std_logic ;
      filter_data_15_13 : IN std_logic ;
      filter_data_15_12 : IN std_logic ;
      filter_data_15_11 : IN std_logic ;
      filter_data_15_10 : IN std_logic ;
      filter_data_15_9 : IN std_logic ;
      filter_data_15_8 : IN std_logic ;
      filter_data_15_7 : IN std_logic ;
      filter_data_15_6 : IN std_logic ;
      filter_data_15_5 : IN std_logic ;
      filter_data_15_4 : IN std_logic ;
      filter_data_15_3 : IN std_logic ;
      filter_data_15_2 : IN std_logic ;
      filter_data_15_1 : IN std_logic ;
      filter_data_15_0 : IN std_logic ;
      filter_data_16_15 : IN std_logic ;
      filter_data_16_14 : IN std_logic ;
      filter_data_16_13 : IN std_logic ;
      filter_data_16_12 : IN std_logic ;
      filter_data_16_11 : IN std_logic ;
      filter_data_16_10 : IN std_logic ;
      filter_data_16_9 : IN std_logic ;
      filter_data_16_8 : IN std_logic ;
      filter_data_16_7 : IN std_logic ;
      filter_data_16_6 : IN std_logic ;
      filter_data_16_5 : IN std_logic ;
      filter_data_16_4 : IN std_logic ;
      filter_data_16_3 : IN std_logic ;
      filter_data_16_2 : IN std_logic ;
      filter_data_16_1 : IN std_logic ;
      filter_data_16_0 : IN std_logic ;
      filter_data_17_15 : IN std_logic ;
      filter_data_17_14 : IN std_logic ;
      filter_data_17_13 : IN std_logic ;
      filter_data_17_12 : IN std_logic ;
      filter_data_17_11 : IN std_logic ;
      filter_data_17_10 : IN std_logic ;
      filter_data_17_9 : IN std_logic ;
      filter_data_17_8 : IN std_logic ;
      filter_data_17_7 : IN std_logic ;
      filter_data_17_6 : IN std_logic ;
      filter_data_17_5 : IN std_logic ;
      filter_data_17_4 : IN std_logic ;
      filter_data_17_3 : IN std_logic ;
      filter_data_17_2 : IN std_logic ;
      filter_data_17_1 : IN std_logic ;
      filter_data_17_0 : IN std_logic ;
      filter_data_18_15 : IN std_logic ;
      filter_data_18_14 : IN std_logic ;
      filter_data_18_13 : IN std_logic ;
      filter_data_18_12 : IN std_logic ;
      filter_data_18_11 : IN std_logic ;
      filter_data_18_10 : IN std_logic ;
      filter_data_18_9 : IN std_logic ;
      filter_data_18_8 : IN std_logic ;
      filter_data_18_7 : IN std_logic ;
      filter_data_18_6 : IN std_logic ;
      filter_data_18_5 : IN std_logic ;
      filter_data_18_4 : IN std_logic ;
      filter_data_18_3 : IN std_logic ;
      filter_data_18_2 : IN std_logic ;
      filter_data_18_1 : IN std_logic ;
      filter_data_18_0 : IN std_logic ;
      filter_data_19_15 : IN std_logic ;
      filter_data_19_14 : IN std_logic ;
      filter_data_19_13 : IN std_logic ;
      filter_data_19_12 : IN std_logic ;
      filter_data_19_11 : IN std_logic ;
      filter_data_19_10 : IN std_logic ;
      filter_data_19_9 : IN std_logic ;
      filter_data_19_8 : IN std_logic ;
      filter_data_19_7 : IN std_logic ;
      filter_data_19_6 : IN std_logic ;
      filter_data_19_5 : IN std_logic ;
      filter_data_19_4 : IN std_logic ;
      filter_data_19_3 : IN std_logic ;
      filter_data_19_2 : IN std_logic ;
      filter_data_19_1 : IN std_logic ;
      filter_data_19_0 : IN std_logic ;
      filter_data_20_15 : IN std_logic ;
      filter_data_20_14 : IN std_logic ;
      filter_data_20_13 : IN std_logic ;
      filter_data_20_12 : IN std_logic ;
      filter_data_20_11 : IN std_logic ;
      filter_data_20_10 : IN std_logic ;
      filter_data_20_9 : IN std_logic ;
      filter_data_20_8 : IN std_logic ;
      filter_data_20_7 : IN std_logic ;
      filter_data_20_6 : IN std_logic ;
      filter_data_20_5 : IN std_logic ;
      filter_data_20_4 : IN std_logic ;
      filter_data_20_3 : IN std_logic ;
      filter_data_20_2 : IN std_logic ;
      filter_data_20_1 : IN std_logic ;
      filter_data_20_0 : IN std_logic ;
      filter_data_21_15 : IN std_logic ;
      filter_data_21_14 : IN std_logic ;
      filter_data_21_13 : IN std_logic ;
      filter_data_21_12 : IN std_logic ;
      filter_data_21_11 : IN std_logic ;
      filter_data_21_10 : IN std_logic ;
      filter_data_21_9 : IN std_logic ;
      filter_data_21_8 : IN std_logic ;
      filter_data_21_7 : IN std_logic ;
      filter_data_21_6 : IN std_logic ;
      filter_data_21_5 : IN std_logic ;
      filter_data_21_4 : IN std_logic ;
      filter_data_21_3 : IN std_logic ;
      filter_data_21_2 : IN std_logic ;
      filter_data_21_1 : IN std_logic ;
      filter_data_21_0 : IN std_logic ;
      filter_data_22_15 : IN std_logic ;
      filter_data_22_14 : IN std_logic ;
      filter_data_22_13 : IN std_logic ;
      filter_data_22_12 : IN std_logic ;
      filter_data_22_11 : IN std_logic ;
      filter_data_22_10 : IN std_logic ;
      filter_data_22_9 : IN std_logic ;
      filter_data_22_8 : IN std_logic ;
      filter_data_22_7 : IN std_logic ;
      filter_data_22_6 : IN std_logic ;
      filter_data_22_5 : IN std_logic ;
      filter_data_22_4 : IN std_logic ;
      filter_data_22_3 : IN std_logic ;
      filter_data_22_2 : IN std_logic ;
      filter_data_22_1 : IN std_logic ;
      filter_data_22_0 : IN std_logic ;
      filter_data_23_15 : IN std_logic ;
      filter_data_23_14 : IN std_logic ;
      filter_data_23_13 : IN std_logic ;
      filter_data_23_12 : IN std_logic ;
      filter_data_23_11 : IN std_logic ;
      filter_data_23_10 : IN std_logic ;
      filter_data_23_9 : IN std_logic ;
      filter_data_23_8 : IN std_logic ;
      filter_data_23_7 : IN std_logic ;
      filter_data_23_6 : IN std_logic ;
      filter_data_23_5 : IN std_logic ;
      filter_data_23_4 : IN std_logic ;
      filter_data_23_3 : IN std_logic ;
      filter_data_23_2 : IN std_logic ;
      filter_data_23_1 : IN std_logic ;
      filter_data_23_0 : IN std_logic ;
      filter_data_24_15 : IN std_logic ;
      filter_data_24_14 : IN std_logic ;
      filter_data_24_13 : IN std_logic ;
      filter_data_24_12 : IN std_logic ;
      filter_data_24_11 : IN std_logic ;
      filter_data_24_10 : IN std_logic ;
      filter_data_24_9 : IN std_logic ;
      filter_data_24_8 : IN std_logic ;
      filter_data_24_7 : IN std_logic ;
      filter_data_24_6 : IN std_logic ;
      filter_data_24_5 : IN std_logic ;
      filter_data_24_4 : IN std_logic ;
      filter_data_24_3 : IN std_logic ;
      filter_data_24_2 : IN std_logic ;
      filter_data_24_1 : IN std_logic ;
      filter_data_24_0 : IN std_logic ;
      d_arr_0_31 : OUT std_logic ;
      d_arr_0_30 : OUT std_logic ;
      d_arr_0_29 : OUT std_logic ;
      d_arr_0_28 : OUT std_logic ;
      d_arr_0_27 : OUT std_logic ;
      d_arr_0_26 : OUT std_logic ;
      d_arr_0_25 : OUT std_logic ;
      d_arr_0_24 : OUT std_logic ;
      d_arr_0_23 : OUT std_logic ;
      d_arr_0_22 : OUT std_logic ;
      d_arr_0_21 : OUT std_logic ;
      d_arr_0_20 : OUT std_logic ;
      d_arr_0_19 : OUT std_logic ;
      d_arr_0_18 : OUT std_logic ;
      d_arr_0_17 : OUT std_logic ;
      d_arr_0_16 : OUT std_logic ;
      d_arr_0_15 : OUT std_logic ;
      d_arr_0_14 : OUT std_logic ;
      d_arr_0_13 : OUT std_logic ;
      d_arr_0_12 : OUT std_logic ;
      d_arr_0_11 : OUT std_logic ;
      d_arr_0_10 : OUT std_logic ;
      d_arr_0_9 : OUT std_logic ;
      d_arr_0_8 : OUT std_logic ;
      d_arr_0_7 : OUT std_logic ;
      d_arr_0_6 : OUT std_logic ;
      d_arr_0_5 : OUT std_logic ;
      d_arr_0_4 : OUT std_logic ;
      d_arr_0_3 : OUT std_logic ;
      d_arr_0_2 : OUT std_logic ;
      d_arr_0_1 : OUT std_logic ;
      d_arr_0_0 : OUT std_logic ;
      d_arr_1_31 : OUT std_logic ;
      d_arr_1_30 : OUT std_logic ;
      d_arr_1_29 : OUT std_logic ;
      d_arr_1_28 : OUT std_logic ;
      d_arr_1_27 : OUT std_logic ;
      d_arr_1_26 : OUT std_logic ;
      d_arr_1_25 : OUT std_logic ;
      d_arr_1_24 : OUT std_logic ;
      d_arr_1_23 : OUT std_logic ;
      d_arr_1_22 : OUT std_logic ;
      d_arr_1_21 : OUT std_logic ;
      d_arr_1_20 : OUT std_logic ;
      d_arr_1_19 : OUT std_logic ;
      d_arr_1_18 : OUT std_logic ;
      d_arr_1_17 : OUT std_logic ;
      d_arr_1_16 : OUT std_logic ;
      d_arr_1_15 : OUT std_logic ;
      d_arr_1_14 : OUT std_logic ;
      d_arr_1_13 : OUT std_logic ;
      d_arr_1_12 : OUT std_logic ;
      d_arr_1_11 : OUT std_logic ;
      d_arr_1_10 : OUT std_logic ;
      d_arr_1_9 : OUT std_logic ;
      d_arr_1_8 : OUT std_logic ;
      d_arr_1_7 : OUT std_logic ;
      d_arr_1_6 : OUT std_logic ;
      d_arr_1_5 : OUT std_logic ;
      d_arr_1_4 : OUT std_logic ;
      d_arr_1_3 : OUT std_logic ;
      d_arr_1_2 : OUT std_logic ;
      d_arr_1_1 : OUT std_logic ;
      d_arr_1_0 : OUT std_logic ;
      d_arr_2_31 : OUT std_logic ;
      d_arr_2_30 : OUT std_logic ;
      d_arr_2_29 : OUT std_logic ;
      d_arr_2_28 : OUT std_logic ;
      d_arr_2_27 : OUT std_logic ;
      d_arr_2_26 : OUT std_logic ;
      d_arr_2_25 : OUT std_logic ;
      d_arr_2_24 : OUT std_logic ;
      d_arr_2_23 : OUT std_logic ;
      d_arr_2_22 : OUT std_logic ;
      d_arr_2_21 : OUT std_logic ;
      d_arr_2_20 : OUT std_logic ;
      d_arr_2_19 : OUT std_logic ;
      d_arr_2_18 : OUT std_logic ;
      d_arr_2_17 : OUT std_logic ;
      d_arr_2_16 : OUT std_logic ;
      d_arr_2_15 : OUT std_logic ;
      d_arr_2_14 : OUT std_logic ;
      d_arr_2_13 : OUT std_logic ;
      d_arr_2_12 : OUT std_logic ;
      d_arr_2_11 : OUT std_logic ;
      d_arr_2_10 : OUT std_logic ;
      d_arr_2_9 : OUT std_logic ;
      d_arr_2_8 : OUT std_logic ;
      d_arr_2_7 : OUT std_logic ;
      d_arr_2_6 : OUT std_logic ;
      d_arr_2_5 : OUT std_logic ;
      d_arr_2_4 : OUT std_logic ;
      d_arr_2_3 : OUT std_logic ;
      d_arr_2_2 : OUT std_logic ;
      d_arr_2_1 : OUT std_logic ;
      d_arr_2_0 : OUT std_logic ;
      d_arr_3_31 : OUT std_logic ;
      d_arr_3_30 : OUT std_logic ;
      d_arr_3_29 : OUT std_logic ;
      d_arr_3_28 : OUT std_logic ;
      d_arr_3_27 : OUT std_logic ;
      d_arr_3_26 : OUT std_logic ;
      d_arr_3_25 : OUT std_logic ;
      d_arr_3_24 : OUT std_logic ;
      d_arr_3_23 : OUT std_logic ;
      d_arr_3_22 : OUT std_logic ;
      d_arr_3_21 : OUT std_logic ;
      d_arr_3_20 : OUT std_logic ;
      d_arr_3_19 : OUT std_logic ;
      d_arr_3_18 : OUT std_logic ;
      d_arr_3_17 : OUT std_logic ;
      d_arr_3_16 : OUT std_logic ;
      d_arr_3_15 : OUT std_logic ;
      d_arr_3_14 : OUT std_logic ;
      d_arr_3_13 : OUT std_logic ;
      d_arr_3_12 : OUT std_logic ;
      d_arr_3_11 : OUT std_logic ;
      d_arr_3_10 : OUT std_logic ;
      d_arr_3_9 : OUT std_logic ;
      d_arr_3_8 : OUT std_logic ;
      d_arr_3_7 : OUT std_logic ;
      d_arr_3_6 : OUT std_logic ;
      d_arr_3_5 : OUT std_logic ;
      d_arr_3_4 : OUT std_logic ;
      d_arr_3_3 : OUT std_logic ;
      d_arr_3_2 : OUT std_logic ;
      d_arr_3_1 : OUT std_logic ;
      d_arr_3_0 : OUT std_logic ;
      d_arr_4_31 : OUT std_logic ;
      d_arr_4_30 : OUT std_logic ;
      d_arr_4_29 : OUT std_logic ;
      d_arr_4_28 : OUT std_logic ;
      d_arr_4_27 : OUT std_logic ;
      d_arr_4_26 : OUT std_logic ;
      d_arr_4_25 : OUT std_logic ;
      d_arr_4_24 : OUT std_logic ;
      d_arr_4_23 : OUT std_logic ;
      d_arr_4_22 : OUT std_logic ;
      d_arr_4_21 : OUT std_logic ;
      d_arr_4_20 : OUT std_logic ;
      d_arr_4_19 : OUT std_logic ;
      d_arr_4_18 : OUT std_logic ;
      d_arr_4_17 : OUT std_logic ;
      d_arr_4_16 : OUT std_logic ;
      d_arr_4_15 : OUT std_logic ;
      d_arr_4_14 : OUT std_logic ;
      d_arr_4_13 : OUT std_logic ;
      d_arr_4_12 : OUT std_logic ;
      d_arr_4_11 : OUT std_logic ;
      d_arr_4_10 : OUT std_logic ;
      d_arr_4_9 : OUT std_logic ;
      d_arr_4_8 : OUT std_logic ;
      d_arr_4_7 : OUT std_logic ;
      d_arr_4_6 : OUT std_logic ;
      d_arr_4_5 : OUT std_logic ;
      d_arr_4_4 : OUT std_logic ;
      d_arr_4_3 : OUT std_logic ;
      d_arr_4_2 : OUT std_logic ;
      d_arr_4_1 : OUT std_logic ;
      d_arr_4_0 : OUT std_logic ;
      d_arr_5_31 : OUT std_logic ;
      d_arr_5_30 : OUT std_logic ;
      d_arr_5_29 : OUT std_logic ;
      d_arr_5_28 : OUT std_logic ;
      d_arr_5_27 : OUT std_logic ;
      d_arr_5_26 : OUT std_logic ;
      d_arr_5_25 : OUT std_logic ;
      d_arr_5_24 : OUT std_logic ;
      d_arr_5_23 : OUT std_logic ;
      d_arr_5_22 : OUT std_logic ;
      d_arr_5_21 : OUT std_logic ;
      d_arr_5_20 : OUT std_logic ;
      d_arr_5_19 : OUT std_logic ;
      d_arr_5_18 : OUT std_logic ;
      d_arr_5_17 : OUT std_logic ;
      d_arr_5_16 : OUT std_logic ;
      d_arr_5_15 : OUT std_logic ;
      d_arr_5_14 : OUT std_logic ;
      d_arr_5_13 : OUT std_logic ;
      d_arr_5_12 : OUT std_logic ;
      d_arr_5_11 : OUT std_logic ;
      d_arr_5_10 : OUT std_logic ;
      d_arr_5_9 : OUT std_logic ;
      d_arr_5_8 : OUT std_logic ;
      d_arr_5_7 : OUT std_logic ;
      d_arr_5_6 : OUT std_logic ;
      d_arr_5_5 : OUT std_logic ;
      d_arr_5_4 : OUT std_logic ;
      d_arr_5_3 : OUT std_logic ;
      d_arr_5_2 : OUT std_logic ;
      d_arr_5_1 : OUT std_logic ;
      d_arr_5_0 : OUT std_logic ;
      d_arr_6_31 : OUT std_logic ;
      d_arr_6_30 : OUT std_logic ;
      d_arr_6_29 : OUT std_logic ;
      d_arr_6_28 : OUT std_logic ;
      d_arr_6_27 : OUT std_logic ;
      d_arr_6_26 : OUT std_logic ;
      d_arr_6_25 : OUT std_logic ;
      d_arr_6_24 : OUT std_logic ;
      d_arr_6_23 : OUT std_logic ;
      d_arr_6_22 : OUT std_logic ;
      d_arr_6_21 : OUT std_logic ;
      d_arr_6_20 : OUT std_logic ;
      d_arr_6_19 : OUT std_logic ;
      d_arr_6_18 : OUT std_logic ;
      d_arr_6_17 : OUT std_logic ;
      d_arr_6_16 : OUT std_logic ;
      d_arr_6_15 : OUT std_logic ;
      d_arr_6_14 : OUT std_logic ;
      d_arr_6_13 : OUT std_logic ;
      d_arr_6_12 : OUT std_logic ;
      d_arr_6_11 : OUT std_logic ;
      d_arr_6_10 : OUT std_logic ;
      d_arr_6_9 : OUT std_logic ;
      d_arr_6_8 : OUT std_logic ;
      d_arr_6_7 : OUT std_logic ;
      d_arr_6_6 : OUT std_logic ;
      d_arr_6_5 : OUT std_logic ;
      d_arr_6_4 : OUT std_logic ;
      d_arr_6_3 : OUT std_logic ;
      d_arr_6_2 : OUT std_logic ;
      d_arr_6_1 : OUT std_logic ;
      d_arr_6_0 : OUT std_logic ;
      d_arr_7_31 : OUT std_logic ;
      d_arr_7_30 : OUT std_logic ;
      d_arr_7_29 : OUT std_logic ;
      d_arr_7_28 : OUT std_logic ;
      d_arr_7_27 : OUT std_logic ;
      d_arr_7_26 : OUT std_logic ;
      d_arr_7_25 : OUT std_logic ;
      d_arr_7_24 : OUT std_logic ;
      d_arr_7_23 : OUT std_logic ;
      d_arr_7_22 : OUT std_logic ;
      d_arr_7_21 : OUT std_logic ;
      d_arr_7_20 : OUT std_logic ;
      d_arr_7_19 : OUT std_logic ;
      d_arr_7_18 : OUT std_logic ;
      d_arr_7_17 : OUT std_logic ;
      d_arr_7_16 : OUT std_logic ;
      d_arr_7_15 : OUT std_logic ;
      d_arr_7_14 : OUT std_logic ;
      d_arr_7_13 : OUT std_logic ;
      d_arr_7_12 : OUT std_logic ;
      d_arr_7_11 : OUT std_logic ;
      d_arr_7_10 : OUT std_logic ;
      d_arr_7_9 : OUT std_logic ;
      d_arr_7_8 : OUT std_logic ;
      d_arr_7_7 : OUT std_logic ;
      d_arr_7_6 : OUT std_logic ;
      d_arr_7_5 : OUT std_logic ;
      d_arr_7_4 : OUT std_logic ;
      d_arr_7_3 : OUT std_logic ;
      d_arr_7_2 : OUT std_logic ;
      d_arr_7_1 : OUT std_logic ;
      d_arr_7_0 : OUT std_logic ;
      d_arr_8_31 : OUT std_logic ;
      d_arr_8_30 : OUT std_logic ;
      d_arr_8_29 : OUT std_logic ;
      d_arr_8_28 : OUT std_logic ;
      d_arr_8_27 : OUT std_logic ;
      d_arr_8_26 : OUT std_logic ;
      d_arr_8_25 : OUT std_logic ;
      d_arr_8_24 : OUT std_logic ;
      d_arr_8_23 : OUT std_logic ;
      d_arr_8_22 : OUT std_logic ;
      d_arr_8_21 : OUT std_logic ;
      d_arr_8_20 : OUT std_logic ;
      d_arr_8_19 : OUT std_logic ;
      d_arr_8_18 : OUT std_logic ;
      d_arr_8_17 : OUT std_logic ;
      d_arr_8_16 : OUT std_logic ;
      d_arr_8_15 : OUT std_logic ;
      d_arr_8_14 : OUT std_logic ;
      d_arr_8_13 : OUT std_logic ;
      d_arr_8_12 : OUT std_logic ;
      d_arr_8_11 : OUT std_logic ;
      d_arr_8_10 : OUT std_logic ;
      d_arr_8_9 : OUT std_logic ;
      d_arr_8_8 : OUT std_logic ;
      d_arr_8_7 : OUT std_logic ;
      d_arr_8_6 : OUT std_logic ;
      d_arr_8_5 : OUT std_logic ;
      d_arr_8_4 : OUT std_logic ;
      d_arr_8_3 : OUT std_logic ;
      d_arr_8_2 : OUT std_logic ;
      d_arr_8_1 : OUT std_logic ;
      d_arr_8_0 : OUT std_logic ;
      d_arr_9_31 : OUT std_logic ;
      d_arr_9_30 : OUT std_logic ;
      d_arr_9_29 : OUT std_logic ;
      d_arr_9_28 : OUT std_logic ;
      d_arr_9_27 : OUT std_logic ;
      d_arr_9_26 : OUT std_logic ;
      d_arr_9_25 : OUT std_logic ;
      d_arr_9_24 : OUT std_logic ;
      d_arr_9_23 : OUT std_logic ;
      d_arr_9_22 : OUT std_logic ;
      d_arr_9_21 : OUT std_logic ;
      d_arr_9_20 : OUT std_logic ;
      d_arr_9_19 : OUT std_logic ;
      d_arr_9_18 : OUT std_logic ;
      d_arr_9_17 : OUT std_logic ;
      d_arr_9_16 : OUT std_logic ;
      d_arr_9_15 : OUT std_logic ;
      d_arr_9_14 : OUT std_logic ;
      d_arr_9_13 : OUT std_logic ;
      d_arr_9_12 : OUT std_logic ;
      d_arr_9_11 : OUT std_logic ;
      d_arr_9_10 : OUT std_logic ;
      d_arr_9_9 : OUT std_logic ;
      d_arr_9_8 : OUT std_logic ;
      d_arr_9_7 : OUT std_logic ;
      d_arr_9_6 : OUT std_logic ;
      d_arr_9_5 : OUT std_logic ;
      d_arr_9_4 : OUT std_logic ;
      d_arr_9_3 : OUT std_logic ;
      d_arr_9_2 : OUT std_logic ;
      d_arr_9_1 : OUT std_logic ;
      d_arr_9_0 : OUT std_logic ;
      d_arr_10_31 : OUT std_logic ;
      d_arr_10_30 : OUT std_logic ;
      d_arr_10_29 : OUT std_logic ;
      d_arr_10_28 : OUT std_logic ;
      d_arr_10_27 : OUT std_logic ;
      d_arr_10_26 : OUT std_logic ;
      d_arr_10_25 : OUT std_logic ;
      d_arr_10_24 : OUT std_logic ;
      d_arr_10_23 : OUT std_logic ;
      d_arr_10_22 : OUT std_logic ;
      d_arr_10_21 : OUT std_logic ;
      d_arr_10_20 : OUT std_logic ;
      d_arr_10_19 : OUT std_logic ;
      d_arr_10_18 : OUT std_logic ;
      d_arr_10_17 : OUT std_logic ;
      d_arr_10_16 : OUT std_logic ;
      d_arr_10_15 : OUT std_logic ;
      d_arr_10_14 : OUT std_logic ;
      d_arr_10_13 : OUT std_logic ;
      d_arr_10_12 : OUT std_logic ;
      d_arr_10_11 : OUT std_logic ;
      d_arr_10_10 : OUT std_logic ;
      d_arr_10_9 : OUT std_logic ;
      d_arr_10_8 : OUT std_logic ;
      d_arr_10_7 : OUT std_logic ;
      d_arr_10_6 : OUT std_logic ;
      d_arr_10_5 : OUT std_logic ;
      d_arr_10_4 : OUT std_logic ;
      d_arr_10_3 : OUT std_logic ;
      d_arr_10_2 : OUT std_logic ;
      d_arr_10_1 : OUT std_logic ;
      d_arr_10_0 : OUT std_logic ;
      d_arr_11_31 : OUT std_logic ;
      d_arr_11_30 : OUT std_logic ;
      d_arr_11_29 : OUT std_logic ;
      d_arr_11_28 : OUT std_logic ;
      d_arr_11_27 : OUT std_logic ;
      d_arr_11_26 : OUT std_logic ;
      d_arr_11_25 : OUT std_logic ;
      d_arr_11_24 : OUT std_logic ;
      d_arr_11_23 : OUT std_logic ;
      d_arr_11_22 : OUT std_logic ;
      d_arr_11_21 : OUT std_logic ;
      d_arr_11_20 : OUT std_logic ;
      d_arr_11_19 : OUT std_logic ;
      d_arr_11_18 : OUT std_logic ;
      d_arr_11_17 : OUT std_logic ;
      d_arr_11_16 : OUT std_logic ;
      d_arr_11_15 : OUT std_logic ;
      d_arr_11_14 : OUT std_logic ;
      d_arr_11_13 : OUT std_logic ;
      d_arr_11_12 : OUT std_logic ;
      d_arr_11_11 : OUT std_logic ;
      d_arr_11_10 : OUT std_logic ;
      d_arr_11_9 : OUT std_logic ;
      d_arr_11_8 : OUT std_logic ;
      d_arr_11_7 : OUT std_logic ;
      d_arr_11_6 : OUT std_logic ;
      d_arr_11_5 : OUT std_logic ;
      d_arr_11_4 : OUT std_logic ;
      d_arr_11_3 : OUT std_logic ;
      d_arr_11_2 : OUT std_logic ;
      d_arr_11_1 : OUT std_logic ;
      d_arr_11_0 : OUT std_logic ;
      d_arr_12_31 : OUT std_logic ;
      d_arr_12_30 : OUT std_logic ;
      d_arr_12_29 : OUT std_logic ;
      d_arr_12_28 : OUT std_logic ;
      d_arr_12_27 : OUT std_logic ;
      d_arr_12_26 : OUT std_logic ;
      d_arr_12_25 : OUT std_logic ;
      d_arr_12_24 : OUT std_logic ;
      d_arr_12_23 : OUT std_logic ;
      d_arr_12_22 : OUT std_logic ;
      d_arr_12_21 : OUT std_logic ;
      d_arr_12_20 : OUT std_logic ;
      d_arr_12_19 : OUT std_logic ;
      d_arr_12_18 : OUT std_logic ;
      d_arr_12_17 : OUT std_logic ;
      d_arr_12_16 : OUT std_logic ;
      d_arr_12_15 : OUT std_logic ;
      d_arr_12_14 : OUT std_logic ;
      d_arr_12_13 : OUT std_logic ;
      d_arr_12_12 : OUT std_logic ;
      d_arr_12_11 : OUT std_logic ;
      d_arr_12_10 : OUT std_logic ;
      d_arr_12_9 : OUT std_logic ;
      d_arr_12_8 : OUT std_logic ;
      d_arr_12_7 : OUT std_logic ;
      d_arr_12_6 : OUT std_logic ;
      d_arr_12_5 : OUT std_logic ;
      d_arr_12_4 : OUT std_logic ;
      d_arr_12_3 : OUT std_logic ;
      d_arr_12_2 : OUT std_logic ;
      d_arr_12_1 : OUT std_logic ;
      d_arr_12_0 : OUT std_logic ;
      d_arr_13_31 : OUT std_logic ;
      d_arr_13_30 : OUT std_logic ;
      d_arr_13_29 : OUT std_logic ;
      d_arr_13_28 : OUT std_logic ;
      d_arr_13_27 : OUT std_logic ;
      d_arr_13_26 : OUT std_logic ;
      d_arr_13_25 : OUT std_logic ;
      d_arr_13_24 : OUT std_logic ;
      d_arr_13_23 : OUT std_logic ;
      d_arr_13_22 : OUT std_logic ;
      d_arr_13_21 : OUT std_logic ;
      d_arr_13_20 : OUT std_logic ;
      d_arr_13_19 : OUT std_logic ;
      d_arr_13_18 : OUT std_logic ;
      d_arr_13_17 : OUT std_logic ;
      d_arr_13_16 : OUT std_logic ;
      d_arr_13_15 : OUT std_logic ;
      d_arr_13_14 : OUT std_logic ;
      d_arr_13_13 : OUT std_logic ;
      d_arr_13_12 : OUT std_logic ;
      d_arr_13_11 : OUT std_logic ;
      d_arr_13_10 : OUT std_logic ;
      d_arr_13_9 : OUT std_logic ;
      d_arr_13_8 : OUT std_logic ;
      d_arr_13_7 : OUT std_logic ;
      d_arr_13_6 : OUT std_logic ;
      d_arr_13_5 : OUT std_logic ;
      d_arr_13_4 : OUT std_logic ;
      d_arr_13_3 : OUT std_logic ;
      d_arr_13_2 : OUT std_logic ;
      d_arr_13_1 : OUT std_logic ;
      d_arr_13_0 : OUT std_logic ;
      d_arr_14_31 : OUT std_logic ;
      d_arr_14_30 : OUT std_logic ;
      d_arr_14_29 : OUT std_logic ;
      d_arr_14_28 : OUT std_logic ;
      d_arr_14_27 : OUT std_logic ;
      d_arr_14_26 : OUT std_logic ;
      d_arr_14_25 : OUT std_logic ;
      d_arr_14_24 : OUT std_logic ;
      d_arr_14_23 : OUT std_logic ;
      d_arr_14_22 : OUT std_logic ;
      d_arr_14_21 : OUT std_logic ;
      d_arr_14_20 : OUT std_logic ;
      d_arr_14_19 : OUT std_logic ;
      d_arr_14_18 : OUT std_logic ;
      d_arr_14_17 : OUT std_logic ;
      d_arr_14_16 : OUT std_logic ;
      d_arr_14_15 : OUT std_logic ;
      d_arr_14_14 : OUT std_logic ;
      d_arr_14_13 : OUT std_logic ;
      d_arr_14_12 : OUT std_logic ;
      d_arr_14_11 : OUT std_logic ;
      d_arr_14_10 : OUT std_logic ;
      d_arr_14_9 : OUT std_logic ;
      d_arr_14_8 : OUT std_logic ;
      d_arr_14_7 : OUT std_logic ;
      d_arr_14_6 : OUT std_logic ;
      d_arr_14_5 : OUT std_logic ;
      d_arr_14_4 : OUT std_logic ;
      d_arr_14_3 : OUT std_logic ;
      d_arr_14_2 : OUT std_logic ;
      d_arr_14_1 : OUT std_logic ;
      d_arr_14_0 : OUT std_logic ;
      d_arr_15_31 : OUT std_logic ;
      d_arr_15_30 : OUT std_logic ;
      d_arr_15_29 : OUT std_logic ;
      d_arr_15_28 : OUT std_logic ;
      d_arr_15_27 : OUT std_logic ;
      d_arr_15_26 : OUT std_logic ;
      d_arr_15_25 : OUT std_logic ;
      d_arr_15_24 : OUT std_logic ;
      d_arr_15_23 : OUT std_logic ;
      d_arr_15_22 : OUT std_logic ;
      d_arr_15_21 : OUT std_logic ;
      d_arr_15_20 : OUT std_logic ;
      d_arr_15_19 : OUT std_logic ;
      d_arr_15_18 : OUT std_logic ;
      d_arr_15_17 : OUT std_logic ;
      d_arr_15_16 : OUT std_logic ;
      d_arr_15_15 : OUT std_logic ;
      d_arr_15_14 : OUT std_logic ;
      d_arr_15_13 : OUT std_logic ;
      d_arr_15_12 : OUT std_logic ;
      d_arr_15_11 : OUT std_logic ;
      d_arr_15_10 : OUT std_logic ;
      d_arr_15_9 : OUT std_logic ;
      d_arr_15_8 : OUT std_logic ;
      d_arr_15_7 : OUT std_logic ;
      d_arr_15_6 : OUT std_logic ;
      d_arr_15_5 : OUT std_logic ;
      d_arr_15_4 : OUT std_logic ;
      d_arr_15_3 : OUT std_logic ;
      d_arr_15_2 : OUT std_logic ;
      d_arr_15_1 : OUT std_logic ;
      d_arr_15_0 : OUT std_logic ;
      d_arr_16_31 : OUT std_logic ;
      d_arr_16_30 : OUT std_logic ;
      d_arr_16_29 : OUT std_logic ;
      d_arr_16_28 : OUT std_logic ;
      d_arr_16_27 : OUT std_logic ;
      d_arr_16_26 : OUT std_logic ;
      d_arr_16_25 : OUT std_logic ;
      d_arr_16_24 : OUT std_logic ;
      d_arr_16_23 : OUT std_logic ;
      d_arr_16_22 : OUT std_logic ;
      d_arr_16_21 : OUT std_logic ;
      d_arr_16_20 : OUT std_logic ;
      d_arr_16_19 : OUT std_logic ;
      d_arr_16_18 : OUT std_logic ;
      d_arr_16_17 : OUT std_logic ;
      d_arr_16_16 : OUT std_logic ;
      d_arr_16_15 : OUT std_logic ;
      d_arr_16_14 : OUT std_logic ;
      d_arr_16_13 : OUT std_logic ;
      d_arr_16_12 : OUT std_logic ;
      d_arr_16_11 : OUT std_logic ;
      d_arr_16_10 : OUT std_logic ;
      d_arr_16_9 : OUT std_logic ;
      d_arr_16_8 : OUT std_logic ;
      d_arr_16_7 : OUT std_logic ;
      d_arr_16_6 : OUT std_logic ;
      d_arr_16_5 : OUT std_logic ;
      d_arr_16_4 : OUT std_logic ;
      d_arr_16_3 : OUT std_logic ;
      d_arr_16_2 : OUT std_logic ;
      d_arr_16_1 : OUT std_logic ;
      d_arr_16_0 : OUT std_logic ;
      d_arr_17_31 : OUT std_logic ;
      d_arr_17_30 : OUT std_logic ;
      d_arr_17_29 : OUT std_logic ;
      d_arr_17_28 : OUT std_logic ;
      d_arr_17_27 : OUT std_logic ;
      d_arr_17_26 : OUT std_logic ;
      d_arr_17_25 : OUT std_logic ;
      d_arr_17_24 : OUT std_logic ;
      d_arr_17_23 : OUT std_logic ;
      d_arr_17_22 : OUT std_logic ;
      d_arr_17_21 : OUT std_logic ;
      d_arr_17_20 : OUT std_logic ;
      d_arr_17_19 : OUT std_logic ;
      d_arr_17_18 : OUT std_logic ;
      d_arr_17_17 : OUT std_logic ;
      d_arr_17_16 : OUT std_logic ;
      d_arr_17_15 : OUT std_logic ;
      d_arr_17_14 : OUT std_logic ;
      d_arr_17_13 : OUT std_logic ;
      d_arr_17_12 : OUT std_logic ;
      d_arr_17_11 : OUT std_logic ;
      d_arr_17_10 : OUT std_logic ;
      d_arr_17_9 : OUT std_logic ;
      d_arr_17_8 : OUT std_logic ;
      d_arr_17_7 : OUT std_logic ;
      d_arr_17_6 : OUT std_logic ;
      d_arr_17_5 : OUT std_logic ;
      d_arr_17_4 : OUT std_logic ;
      d_arr_17_3 : OUT std_logic ;
      d_arr_17_2 : OUT std_logic ;
      d_arr_17_1 : OUT std_logic ;
      d_arr_17_0 : OUT std_logic ;
      d_arr_18_31 : OUT std_logic ;
      d_arr_18_30 : OUT std_logic ;
      d_arr_18_29 : OUT std_logic ;
      d_arr_18_28 : OUT std_logic ;
      d_arr_18_27 : OUT std_logic ;
      d_arr_18_26 : OUT std_logic ;
      d_arr_18_25 : OUT std_logic ;
      d_arr_18_24 : OUT std_logic ;
      d_arr_18_23 : OUT std_logic ;
      d_arr_18_22 : OUT std_logic ;
      d_arr_18_21 : OUT std_logic ;
      d_arr_18_20 : OUT std_logic ;
      d_arr_18_19 : OUT std_logic ;
      d_arr_18_18 : OUT std_logic ;
      d_arr_18_17 : OUT std_logic ;
      d_arr_18_16 : OUT std_logic ;
      d_arr_18_15 : OUT std_logic ;
      d_arr_18_14 : OUT std_logic ;
      d_arr_18_13 : OUT std_logic ;
      d_arr_18_12 : OUT std_logic ;
      d_arr_18_11 : OUT std_logic ;
      d_arr_18_10 : OUT std_logic ;
      d_arr_18_9 : OUT std_logic ;
      d_arr_18_8 : OUT std_logic ;
      d_arr_18_7 : OUT std_logic ;
      d_arr_18_6 : OUT std_logic ;
      d_arr_18_5 : OUT std_logic ;
      d_arr_18_4 : OUT std_logic ;
      d_arr_18_3 : OUT std_logic ;
      d_arr_18_2 : OUT std_logic ;
      d_arr_18_1 : OUT std_logic ;
      d_arr_18_0 : OUT std_logic ;
      d_arr_19_31 : OUT std_logic ;
      d_arr_19_30 : OUT std_logic ;
      d_arr_19_29 : OUT std_logic ;
      d_arr_19_28 : OUT std_logic ;
      d_arr_19_27 : OUT std_logic ;
      d_arr_19_26 : OUT std_logic ;
      d_arr_19_25 : OUT std_logic ;
      d_arr_19_24 : OUT std_logic ;
      d_arr_19_23 : OUT std_logic ;
      d_arr_19_22 : OUT std_logic ;
      d_arr_19_21 : OUT std_logic ;
      d_arr_19_20 : OUT std_logic ;
      d_arr_19_19 : OUT std_logic ;
      d_arr_19_18 : OUT std_logic ;
      d_arr_19_17 : OUT std_logic ;
      d_arr_19_16 : OUT std_logic ;
      d_arr_19_15 : OUT std_logic ;
      d_arr_19_14 : OUT std_logic ;
      d_arr_19_13 : OUT std_logic ;
      d_arr_19_12 : OUT std_logic ;
      d_arr_19_11 : OUT std_logic ;
      d_arr_19_10 : OUT std_logic ;
      d_arr_19_9 : OUT std_logic ;
      d_arr_19_8 : OUT std_logic ;
      d_arr_19_7 : OUT std_logic ;
      d_arr_19_6 : OUT std_logic ;
      d_arr_19_5 : OUT std_logic ;
      d_arr_19_4 : OUT std_logic ;
      d_arr_19_3 : OUT std_logic ;
      d_arr_19_2 : OUT std_logic ;
      d_arr_19_1 : OUT std_logic ;
      d_arr_19_0 : OUT std_logic ;
      d_arr_20_31 : OUT std_logic ;
      d_arr_20_30 : OUT std_logic ;
      d_arr_20_29 : OUT std_logic ;
      d_arr_20_28 : OUT std_logic ;
      d_arr_20_27 : OUT std_logic ;
      d_arr_20_26 : OUT std_logic ;
      d_arr_20_25 : OUT std_logic ;
      d_arr_20_24 : OUT std_logic ;
      d_arr_20_23 : OUT std_logic ;
      d_arr_20_22 : OUT std_logic ;
      d_arr_20_21 : OUT std_logic ;
      d_arr_20_20 : OUT std_logic ;
      d_arr_20_19 : OUT std_logic ;
      d_arr_20_18 : OUT std_logic ;
      d_arr_20_17 : OUT std_logic ;
      d_arr_20_16 : OUT std_logic ;
      d_arr_20_15 : OUT std_logic ;
      d_arr_20_14 : OUT std_logic ;
      d_arr_20_13 : OUT std_logic ;
      d_arr_20_12 : OUT std_logic ;
      d_arr_20_11 : OUT std_logic ;
      d_arr_20_10 : OUT std_logic ;
      d_arr_20_9 : OUT std_logic ;
      d_arr_20_8 : OUT std_logic ;
      d_arr_20_7 : OUT std_logic ;
      d_arr_20_6 : OUT std_logic ;
      d_arr_20_5 : OUT std_logic ;
      d_arr_20_4 : OUT std_logic ;
      d_arr_20_3 : OUT std_logic ;
      d_arr_20_2 : OUT std_logic ;
      d_arr_20_1 : OUT std_logic ;
      d_arr_20_0 : OUT std_logic ;
      d_arr_21_31 : OUT std_logic ;
      d_arr_21_30 : OUT std_logic ;
      d_arr_21_29 : OUT std_logic ;
      d_arr_21_28 : OUT std_logic ;
      d_arr_21_27 : OUT std_logic ;
      d_arr_21_26 : OUT std_logic ;
      d_arr_21_25 : OUT std_logic ;
      d_arr_21_24 : OUT std_logic ;
      d_arr_21_23 : OUT std_logic ;
      d_arr_21_22 : OUT std_logic ;
      d_arr_21_21 : OUT std_logic ;
      d_arr_21_20 : OUT std_logic ;
      d_arr_21_19 : OUT std_logic ;
      d_arr_21_18 : OUT std_logic ;
      d_arr_21_17 : OUT std_logic ;
      d_arr_21_16 : OUT std_logic ;
      d_arr_21_15 : OUT std_logic ;
      d_arr_21_14 : OUT std_logic ;
      d_arr_21_13 : OUT std_logic ;
      d_arr_21_12 : OUT std_logic ;
      d_arr_21_11 : OUT std_logic ;
      d_arr_21_10 : OUT std_logic ;
      d_arr_21_9 : OUT std_logic ;
      d_arr_21_8 : OUT std_logic ;
      d_arr_21_7 : OUT std_logic ;
      d_arr_21_6 : OUT std_logic ;
      d_arr_21_5 : OUT std_logic ;
      d_arr_21_4 : OUT std_logic ;
      d_arr_21_3 : OUT std_logic ;
      d_arr_21_2 : OUT std_logic ;
      d_arr_21_1 : OUT std_logic ;
      d_arr_21_0 : OUT std_logic ;
      d_arr_22_31 : OUT std_logic ;
      d_arr_22_30 : OUT std_logic ;
      d_arr_22_29 : OUT std_logic ;
      d_arr_22_28 : OUT std_logic ;
      d_arr_22_27 : OUT std_logic ;
      d_arr_22_26 : OUT std_logic ;
      d_arr_22_25 : OUT std_logic ;
      d_arr_22_24 : OUT std_logic ;
      d_arr_22_23 : OUT std_logic ;
      d_arr_22_22 : OUT std_logic ;
      d_arr_22_21 : OUT std_logic ;
      d_arr_22_20 : OUT std_logic ;
      d_arr_22_19 : OUT std_logic ;
      d_arr_22_18 : OUT std_logic ;
      d_arr_22_17 : OUT std_logic ;
      d_arr_22_16 : OUT std_logic ;
      d_arr_22_15 : OUT std_logic ;
      d_arr_22_14 : OUT std_logic ;
      d_arr_22_13 : OUT std_logic ;
      d_arr_22_12 : OUT std_logic ;
      d_arr_22_11 : OUT std_logic ;
      d_arr_22_10 : OUT std_logic ;
      d_arr_22_9 : OUT std_logic ;
      d_arr_22_8 : OUT std_logic ;
      d_arr_22_7 : OUT std_logic ;
      d_arr_22_6 : OUT std_logic ;
      d_arr_22_5 : OUT std_logic ;
      d_arr_22_4 : OUT std_logic ;
      d_arr_22_3 : OUT std_logic ;
      d_arr_22_2 : OUT std_logic ;
      d_arr_22_1 : OUT std_logic ;
      d_arr_22_0 : OUT std_logic ;
      d_arr_23_31 : OUT std_logic ;
      d_arr_23_30 : OUT std_logic ;
      d_arr_23_29 : OUT std_logic ;
      d_arr_23_28 : OUT std_logic ;
      d_arr_23_27 : OUT std_logic ;
      d_arr_23_26 : OUT std_logic ;
      d_arr_23_25 : OUT std_logic ;
      d_arr_23_24 : OUT std_logic ;
      d_arr_23_23 : OUT std_logic ;
      d_arr_23_22 : OUT std_logic ;
      d_arr_23_21 : OUT std_logic ;
      d_arr_23_20 : OUT std_logic ;
      d_arr_23_19 : OUT std_logic ;
      d_arr_23_18 : OUT std_logic ;
      d_arr_23_17 : OUT std_logic ;
      d_arr_23_16 : OUT std_logic ;
      d_arr_23_15 : OUT std_logic ;
      d_arr_23_14 : OUT std_logic ;
      d_arr_23_13 : OUT std_logic ;
      d_arr_23_12 : OUT std_logic ;
      d_arr_23_11 : OUT std_logic ;
      d_arr_23_10 : OUT std_logic ;
      d_arr_23_9 : OUT std_logic ;
      d_arr_23_8 : OUT std_logic ;
      d_arr_23_7 : OUT std_logic ;
      d_arr_23_6 : OUT std_logic ;
      d_arr_23_5 : OUT std_logic ;
      d_arr_23_4 : OUT std_logic ;
      d_arr_23_3 : OUT std_logic ;
      d_arr_23_2 : OUT std_logic ;
      d_arr_23_1 : OUT std_logic ;
      d_arr_23_0 : OUT std_logic ;
      d_arr_24_31 : OUT std_logic ;
      d_arr_24_30 : OUT std_logic ;
      d_arr_24_29 : OUT std_logic ;
      d_arr_24_28 : OUT std_logic ;
      d_arr_24_27 : OUT std_logic ;
      d_arr_24_26 : OUT std_logic ;
      d_arr_24_25 : OUT std_logic ;
      d_arr_24_24 : OUT std_logic ;
      d_arr_24_23 : OUT std_logic ;
      d_arr_24_22 : OUT std_logic ;
      d_arr_24_21 : OUT std_logic ;
      d_arr_24_20 : OUT std_logic ;
      d_arr_24_19 : OUT std_logic ;
      d_arr_24_18 : OUT std_logic ;
      d_arr_24_17 : OUT std_logic ;
      d_arr_24_16 : OUT std_logic ;
      d_arr_24_15 : OUT std_logic ;
      d_arr_24_14 : OUT std_logic ;
      d_arr_24_13 : OUT std_logic ;
      d_arr_24_12 : OUT std_logic ;
      d_arr_24_11 : OUT std_logic ;
      d_arr_24_10 : OUT std_logic ;
      d_arr_24_9 : OUT std_logic ;
      d_arr_24_8 : OUT std_logic ;
      d_arr_24_7 : OUT std_logic ;
      d_arr_24_6 : OUT std_logic ;
      d_arr_24_5 : OUT std_logic ;
      d_arr_24_4 : OUT std_logic ;
      d_arr_24_3 : OUT std_logic ;
      d_arr_24_2 : OUT std_logic ;
      d_arr_24_1 : OUT std_logic ;
      d_arr_24_0 : OUT std_logic ;
      q_arr_0_31 : IN std_logic ;
      q_arr_0_30 : IN std_logic ;
      q_arr_0_29 : IN std_logic ;
      q_arr_0_28 : IN std_logic ;
      q_arr_0_27 : IN std_logic ;
      q_arr_0_26 : IN std_logic ;
      q_arr_0_25 : IN std_logic ;
      q_arr_0_24 : IN std_logic ;
      q_arr_0_23 : IN std_logic ;
      q_arr_0_22 : IN std_logic ;
      q_arr_0_21 : IN std_logic ;
      q_arr_0_20 : IN std_logic ;
      q_arr_0_19 : IN std_logic ;
      q_arr_0_18 : IN std_logic ;
      q_arr_0_17 : IN std_logic ;
      q_arr_0_16 : IN std_logic ;
      q_arr_0_15 : IN std_logic ;
      q_arr_0_14 : IN std_logic ;
      q_arr_0_13 : IN std_logic ;
      q_arr_0_12 : IN std_logic ;
      q_arr_0_11 : IN std_logic ;
      q_arr_0_10 : IN std_logic ;
      q_arr_0_9 : IN std_logic ;
      q_arr_0_8 : IN std_logic ;
      q_arr_0_7 : IN std_logic ;
      q_arr_0_6 : IN std_logic ;
      q_arr_0_5 : IN std_logic ;
      q_arr_0_4 : IN std_logic ;
      q_arr_0_3 : IN std_logic ;
      q_arr_0_2 : IN std_logic ;
      q_arr_0_1 : IN std_logic ;
      q_arr_0_0 : IN std_logic ;
      q_arr_1_31 : IN std_logic ;
      q_arr_1_30 : IN std_logic ;
      q_arr_1_29 : IN std_logic ;
      q_arr_1_28 : IN std_logic ;
      q_arr_1_27 : IN std_logic ;
      q_arr_1_26 : IN std_logic ;
      q_arr_1_25 : IN std_logic ;
      q_arr_1_24 : IN std_logic ;
      q_arr_1_23 : IN std_logic ;
      q_arr_1_22 : IN std_logic ;
      q_arr_1_21 : IN std_logic ;
      q_arr_1_20 : IN std_logic ;
      q_arr_1_19 : IN std_logic ;
      q_arr_1_18 : IN std_logic ;
      q_arr_1_17 : IN std_logic ;
      q_arr_1_16 : IN std_logic ;
      q_arr_1_15 : IN std_logic ;
      q_arr_1_14 : IN std_logic ;
      q_arr_1_13 : IN std_logic ;
      q_arr_1_12 : IN std_logic ;
      q_arr_1_11 : IN std_logic ;
      q_arr_1_10 : IN std_logic ;
      q_arr_1_9 : IN std_logic ;
      q_arr_1_8 : IN std_logic ;
      q_arr_1_7 : IN std_logic ;
      q_arr_1_6 : IN std_logic ;
      q_arr_1_5 : IN std_logic ;
      q_arr_1_4 : IN std_logic ;
      q_arr_1_3 : IN std_logic ;
      q_arr_1_2 : IN std_logic ;
      q_arr_1_1 : IN std_logic ;
      q_arr_1_0 : IN std_logic ;
      q_arr_2_31 : IN std_logic ;
      q_arr_2_30 : IN std_logic ;
      q_arr_2_29 : IN std_logic ;
      q_arr_2_28 : IN std_logic ;
      q_arr_2_27 : IN std_logic ;
      q_arr_2_26 : IN std_logic ;
      q_arr_2_25 : IN std_logic ;
      q_arr_2_24 : IN std_logic ;
      q_arr_2_23 : IN std_logic ;
      q_arr_2_22 : IN std_logic ;
      q_arr_2_21 : IN std_logic ;
      q_arr_2_20 : IN std_logic ;
      q_arr_2_19 : IN std_logic ;
      q_arr_2_18 : IN std_logic ;
      q_arr_2_17 : IN std_logic ;
      q_arr_2_16 : IN std_logic ;
      q_arr_2_15 : IN std_logic ;
      q_arr_2_14 : IN std_logic ;
      q_arr_2_13 : IN std_logic ;
      q_arr_2_12 : IN std_logic ;
      q_arr_2_11 : IN std_logic ;
      q_arr_2_10 : IN std_logic ;
      q_arr_2_9 : IN std_logic ;
      q_arr_2_8 : IN std_logic ;
      q_arr_2_7 : IN std_logic ;
      q_arr_2_6 : IN std_logic ;
      q_arr_2_5 : IN std_logic ;
      q_arr_2_4 : IN std_logic ;
      q_arr_2_3 : IN std_logic ;
      q_arr_2_2 : IN std_logic ;
      q_arr_2_1 : IN std_logic ;
      q_arr_2_0 : IN std_logic ;
      q_arr_3_31 : IN std_logic ;
      q_arr_3_30 : IN std_logic ;
      q_arr_3_29 : IN std_logic ;
      q_arr_3_28 : IN std_logic ;
      q_arr_3_27 : IN std_logic ;
      q_arr_3_26 : IN std_logic ;
      q_arr_3_25 : IN std_logic ;
      q_arr_3_24 : IN std_logic ;
      q_arr_3_23 : IN std_logic ;
      q_arr_3_22 : IN std_logic ;
      q_arr_3_21 : IN std_logic ;
      q_arr_3_20 : IN std_logic ;
      q_arr_3_19 : IN std_logic ;
      q_arr_3_18 : IN std_logic ;
      q_arr_3_17 : IN std_logic ;
      q_arr_3_16 : IN std_logic ;
      q_arr_3_15 : IN std_logic ;
      q_arr_3_14 : IN std_logic ;
      q_arr_3_13 : IN std_logic ;
      q_arr_3_12 : IN std_logic ;
      q_arr_3_11 : IN std_logic ;
      q_arr_3_10 : IN std_logic ;
      q_arr_3_9 : IN std_logic ;
      q_arr_3_8 : IN std_logic ;
      q_arr_3_7 : IN std_logic ;
      q_arr_3_6 : IN std_logic ;
      q_arr_3_5 : IN std_logic ;
      q_arr_3_4 : IN std_logic ;
      q_arr_3_3 : IN std_logic ;
      q_arr_3_2 : IN std_logic ;
      q_arr_3_1 : IN std_logic ;
      q_arr_3_0 : IN std_logic ;
      q_arr_4_31 : IN std_logic ;
      q_arr_4_30 : IN std_logic ;
      q_arr_4_29 : IN std_logic ;
      q_arr_4_28 : IN std_logic ;
      q_arr_4_27 : IN std_logic ;
      q_arr_4_26 : IN std_logic ;
      q_arr_4_25 : IN std_logic ;
      q_arr_4_24 : IN std_logic ;
      q_arr_4_23 : IN std_logic ;
      q_arr_4_22 : IN std_logic ;
      q_arr_4_21 : IN std_logic ;
      q_arr_4_20 : IN std_logic ;
      q_arr_4_19 : IN std_logic ;
      q_arr_4_18 : IN std_logic ;
      q_arr_4_17 : IN std_logic ;
      q_arr_4_16 : IN std_logic ;
      q_arr_4_15 : IN std_logic ;
      q_arr_4_14 : IN std_logic ;
      q_arr_4_13 : IN std_logic ;
      q_arr_4_12 : IN std_logic ;
      q_arr_4_11 : IN std_logic ;
      q_arr_4_10 : IN std_logic ;
      q_arr_4_9 : IN std_logic ;
      q_arr_4_8 : IN std_logic ;
      q_arr_4_7 : IN std_logic ;
      q_arr_4_6 : IN std_logic ;
      q_arr_4_5 : IN std_logic ;
      q_arr_4_4 : IN std_logic ;
      q_arr_4_3 : IN std_logic ;
      q_arr_4_2 : IN std_logic ;
      q_arr_4_1 : IN std_logic ;
      q_arr_4_0 : IN std_logic ;
      q_arr_5_31 : IN std_logic ;
      q_arr_5_30 : IN std_logic ;
      q_arr_5_29 : IN std_logic ;
      q_arr_5_28 : IN std_logic ;
      q_arr_5_27 : IN std_logic ;
      q_arr_5_26 : IN std_logic ;
      q_arr_5_25 : IN std_logic ;
      q_arr_5_24 : IN std_logic ;
      q_arr_5_23 : IN std_logic ;
      q_arr_5_22 : IN std_logic ;
      q_arr_5_21 : IN std_logic ;
      q_arr_5_20 : IN std_logic ;
      q_arr_5_19 : IN std_logic ;
      q_arr_5_18 : IN std_logic ;
      q_arr_5_17 : IN std_logic ;
      q_arr_5_16 : IN std_logic ;
      q_arr_5_15 : IN std_logic ;
      q_arr_5_14 : IN std_logic ;
      q_arr_5_13 : IN std_logic ;
      q_arr_5_12 : IN std_logic ;
      q_arr_5_11 : IN std_logic ;
      q_arr_5_10 : IN std_logic ;
      q_arr_5_9 : IN std_logic ;
      q_arr_5_8 : IN std_logic ;
      q_arr_5_7 : IN std_logic ;
      q_arr_5_6 : IN std_logic ;
      q_arr_5_5 : IN std_logic ;
      q_arr_5_4 : IN std_logic ;
      q_arr_5_3 : IN std_logic ;
      q_arr_5_2 : IN std_logic ;
      q_arr_5_1 : IN std_logic ;
      q_arr_5_0 : IN std_logic ;
      q_arr_6_31 : IN std_logic ;
      q_arr_6_30 : IN std_logic ;
      q_arr_6_29 : IN std_logic ;
      q_arr_6_28 : IN std_logic ;
      q_arr_6_27 : IN std_logic ;
      q_arr_6_26 : IN std_logic ;
      q_arr_6_25 : IN std_logic ;
      q_arr_6_24 : IN std_logic ;
      q_arr_6_23 : IN std_logic ;
      q_arr_6_22 : IN std_logic ;
      q_arr_6_21 : IN std_logic ;
      q_arr_6_20 : IN std_logic ;
      q_arr_6_19 : IN std_logic ;
      q_arr_6_18 : IN std_logic ;
      q_arr_6_17 : IN std_logic ;
      q_arr_6_16 : IN std_logic ;
      q_arr_6_15 : IN std_logic ;
      q_arr_6_14 : IN std_logic ;
      q_arr_6_13 : IN std_logic ;
      q_arr_6_12 : IN std_logic ;
      q_arr_6_11 : IN std_logic ;
      q_arr_6_10 : IN std_logic ;
      q_arr_6_9 : IN std_logic ;
      q_arr_6_8 : IN std_logic ;
      q_arr_6_7 : IN std_logic ;
      q_arr_6_6 : IN std_logic ;
      q_arr_6_5 : IN std_logic ;
      q_arr_6_4 : IN std_logic ;
      q_arr_6_3 : IN std_logic ;
      q_arr_6_2 : IN std_logic ;
      q_arr_6_1 : IN std_logic ;
      q_arr_6_0 : IN std_logic ;
      q_arr_7_31 : IN std_logic ;
      q_arr_7_30 : IN std_logic ;
      q_arr_7_29 : IN std_logic ;
      q_arr_7_28 : IN std_logic ;
      q_arr_7_27 : IN std_logic ;
      q_arr_7_26 : IN std_logic ;
      q_arr_7_25 : IN std_logic ;
      q_arr_7_24 : IN std_logic ;
      q_arr_7_23 : IN std_logic ;
      q_arr_7_22 : IN std_logic ;
      q_arr_7_21 : IN std_logic ;
      q_arr_7_20 : IN std_logic ;
      q_arr_7_19 : IN std_logic ;
      q_arr_7_18 : IN std_logic ;
      q_arr_7_17 : IN std_logic ;
      q_arr_7_16 : IN std_logic ;
      q_arr_7_15 : IN std_logic ;
      q_arr_7_14 : IN std_logic ;
      q_arr_7_13 : IN std_logic ;
      q_arr_7_12 : IN std_logic ;
      q_arr_7_11 : IN std_logic ;
      q_arr_7_10 : IN std_logic ;
      q_arr_7_9 : IN std_logic ;
      q_arr_7_8 : IN std_logic ;
      q_arr_7_7 : IN std_logic ;
      q_arr_7_6 : IN std_logic ;
      q_arr_7_5 : IN std_logic ;
      q_arr_7_4 : IN std_logic ;
      q_arr_7_3 : IN std_logic ;
      q_arr_7_2 : IN std_logic ;
      q_arr_7_1 : IN std_logic ;
      q_arr_7_0 : IN std_logic ;
      q_arr_8_31 : IN std_logic ;
      q_arr_8_30 : IN std_logic ;
      q_arr_8_29 : IN std_logic ;
      q_arr_8_28 : IN std_logic ;
      q_arr_8_27 : IN std_logic ;
      q_arr_8_26 : IN std_logic ;
      q_arr_8_25 : IN std_logic ;
      q_arr_8_24 : IN std_logic ;
      q_arr_8_23 : IN std_logic ;
      q_arr_8_22 : IN std_logic ;
      q_arr_8_21 : IN std_logic ;
      q_arr_8_20 : IN std_logic ;
      q_arr_8_19 : IN std_logic ;
      q_arr_8_18 : IN std_logic ;
      q_arr_8_17 : IN std_logic ;
      q_arr_8_16 : IN std_logic ;
      q_arr_8_15 : IN std_logic ;
      q_arr_8_14 : IN std_logic ;
      q_arr_8_13 : IN std_logic ;
      q_arr_8_12 : IN std_logic ;
      q_arr_8_11 : IN std_logic ;
      q_arr_8_10 : IN std_logic ;
      q_arr_8_9 : IN std_logic ;
      q_arr_8_8 : IN std_logic ;
      q_arr_8_7 : IN std_logic ;
      q_arr_8_6 : IN std_logic ;
      q_arr_8_5 : IN std_logic ;
      q_arr_8_4 : IN std_logic ;
      q_arr_8_3 : IN std_logic ;
      q_arr_8_2 : IN std_logic ;
      q_arr_8_1 : IN std_logic ;
      q_arr_8_0 : IN std_logic ;
      q_arr_9_31 : IN std_logic ;
      q_arr_9_30 : IN std_logic ;
      q_arr_9_29 : IN std_logic ;
      q_arr_9_28 : IN std_logic ;
      q_arr_9_27 : IN std_logic ;
      q_arr_9_26 : IN std_logic ;
      q_arr_9_25 : IN std_logic ;
      q_arr_9_24 : IN std_logic ;
      q_arr_9_23 : IN std_logic ;
      q_arr_9_22 : IN std_logic ;
      q_arr_9_21 : IN std_logic ;
      q_arr_9_20 : IN std_logic ;
      q_arr_9_19 : IN std_logic ;
      q_arr_9_18 : IN std_logic ;
      q_arr_9_17 : IN std_logic ;
      q_arr_9_16 : IN std_logic ;
      q_arr_9_15 : IN std_logic ;
      q_arr_9_14 : IN std_logic ;
      q_arr_9_13 : IN std_logic ;
      q_arr_9_12 : IN std_logic ;
      q_arr_9_11 : IN std_logic ;
      q_arr_9_10 : IN std_logic ;
      q_arr_9_9 : IN std_logic ;
      q_arr_9_8 : IN std_logic ;
      q_arr_9_7 : IN std_logic ;
      q_arr_9_6 : IN std_logic ;
      q_arr_9_5 : IN std_logic ;
      q_arr_9_4 : IN std_logic ;
      q_arr_9_3 : IN std_logic ;
      q_arr_9_2 : IN std_logic ;
      q_arr_9_1 : IN std_logic ;
      q_arr_9_0 : IN std_logic ;
      q_arr_10_31 : IN std_logic ;
      q_arr_10_30 : IN std_logic ;
      q_arr_10_29 : IN std_logic ;
      q_arr_10_28 : IN std_logic ;
      q_arr_10_27 : IN std_logic ;
      q_arr_10_26 : IN std_logic ;
      q_arr_10_25 : IN std_logic ;
      q_arr_10_24 : IN std_logic ;
      q_arr_10_23 : IN std_logic ;
      q_arr_10_22 : IN std_logic ;
      q_arr_10_21 : IN std_logic ;
      q_arr_10_20 : IN std_logic ;
      q_arr_10_19 : IN std_logic ;
      q_arr_10_18 : IN std_logic ;
      q_arr_10_17 : IN std_logic ;
      q_arr_10_16 : IN std_logic ;
      q_arr_10_15 : IN std_logic ;
      q_arr_10_14 : IN std_logic ;
      q_arr_10_13 : IN std_logic ;
      q_arr_10_12 : IN std_logic ;
      q_arr_10_11 : IN std_logic ;
      q_arr_10_10 : IN std_logic ;
      q_arr_10_9 : IN std_logic ;
      q_arr_10_8 : IN std_logic ;
      q_arr_10_7 : IN std_logic ;
      q_arr_10_6 : IN std_logic ;
      q_arr_10_5 : IN std_logic ;
      q_arr_10_4 : IN std_logic ;
      q_arr_10_3 : IN std_logic ;
      q_arr_10_2 : IN std_logic ;
      q_arr_10_1 : IN std_logic ;
      q_arr_10_0 : IN std_logic ;
      q_arr_11_31 : IN std_logic ;
      q_arr_11_30 : IN std_logic ;
      q_arr_11_29 : IN std_logic ;
      q_arr_11_28 : IN std_logic ;
      q_arr_11_27 : IN std_logic ;
      q_arr_11_26 : IN std_logic ;
      q_arr_11_25 : IN std_logic ;
      q_arr_11_24 : IN std_logic ;
      q_arr_11_23 : IN std_logic ;
      q_arr_11_22 : IN std_logic ;
      q_arr_11_21 : IN std_logic ;
      q_arr_11_20 : IN std_logic ;
      q_arr_11_19 : IN std_logic ;
      q_arr_11_18 : IN std_logic ;
      q_arr_11_17 : IN std_logic ;
      q_arr_11_16 : IN std_logic ;
      q_arr_11_15 : IN std_logic ;
      q_arr_11_14 : IN std_logic ;
      q_arr_11_13 : IN std_logic ;
      q_arr_11_12 : IN std_logic ;
      q_arr_11_11 : IN std_logic ;
      q_arr_11_10 : IN std_logic ;
      q_arr_11_9 : IN std_logic ;
      q_arr_11_8 : IN std_logic ;
      q_arr_11_7 : IN std_logic ;
      q_arr_11_6 : IN std_logic ;
      q_arr_11_5 : IN std_logic ;
      q_arr_11_4 : IN std_logic ;
      q_arr_11_3 : IN std_logic ;
      q_arr_11_2 : IN std_logic ;
      q_arr_11_1 : IN std_logic ;
      q_arr_11_0 : IN std_logic ;
      q_arr_12_31 : IN std_logic ;
      q_arr_12_30 : IN std_logic ;
      q_arr_12_29 : IN std_logic ;
      q_arr_12_28 : IN std_logic ;
      q_arr_12_27 : IN std_logic ;
      q_arr_12_26 : IN std_logic ;
      q_arr_12_25 : IN std_logic ;
      q_arr_12_24 : IN std_logic ;
      q_arr_12_23 : IN std_logic ;
      q_arr_12_22 : IN std_logic ;
      q_arr_12_21 : IN std_logic ;
      q_arr_12_20 : IN std_logic ;
      q_arr_12_19 : IN std_logic ;
      q_arr_12_18 : IN std_logic ;
      q_arr_12_17 : IN std_logic ;
      q_arr_12_16 : IN std_logic ;
      q_arr_12_15 : IN std_logic ;
      q_arr_12_14 : IN std_logic ;
      q_arr_12_13 : IN std_logic ;
      q_arr_12_12 : IN std_logic ;
      q_arr_12_11 : IN std_logic ;
      q_arr_12_10 : IN std_logic ;
      q_arr_12_9 : IN std_logic ;
      q_arr_12_8 : IN std_logic ;
      q_arr_12_7 : IN std_logic ;
      q_arr_12_6 : IN std_logic ;
      q_arr_12_5 : IN std_logic ;
      q_arr_12_4 : IN std_logic ;
      q_arr_12_3 : IN std_logic ;
      q_arr_12_2 : IN std_logic ;
      q_arr_12_1 : IN std_logic ;
      q_arr_12_0 : IN std_logic ;
      q_arr_13_31 : IN std_logic ;
      q_arr_13_30 : IN std_logic ;
      q_arr_13_29 : IN std_logic ;
      q_arr_13_28 : IN std_logic ;
      q_arr_13_27 : IN std_logic ;
      q_arr_13_26 : IN std_logic ;
      q_arr_13_25 : IN std_logic ;
      q_arr_13_24 : IN std_logic ;
      q_arr_13_23 : IN std_logic ;
      q_arr_13_22 : IN std_logic ;
      q_arr_13_21 : IN std_logic ;
      q_arr_13_20 : IN std_logic ;
      q_arr_13_19 : IN std_logic ;
      q_arr_13_18 : IN std_logic ;
      q_arr_13_17 : IN std_logic ;
      q_arr_13_16 : IN std_logic ;
      q_arr_13_15 : IN std_logic ;
      q_arr_13_14 : IN std_logic ;
      q_arr_13_13 : IN std_logic ;
      q_arr_13_12 : IN std_logic ;
      q_arr_13_11 : IN std_logic ;
      q_arr_13_10 : IN std_logic ;
      q_arr_13_9 : IN std_logic ;
      q_arr_13_8 : IN std_logic ;
      q_arr_13_7 : IN std_logic ;
      q_arr_13_6 : IN std_logic ;
      q_arr_13_5 : IN std_logic ;
      q_arr_13_4 : IN std_logic ;
      q_arr_13_3 : IN std_logic ;
      q_arr_13_2 : IN std_logic ;
      q_arr_13_1 : IN std_logic ;
      q_arr_13_0 : IN std_logic ;
      q_arr_14_31 : IN std_logic ;
      q_arr_14_30 : IN std_logic ;
      q_arr_14_29 : IN std_logic ;
      q_arr_14_28 : IN std_logic ;
      q_arr_14_27 : IN std_logic ;
      q_arr_14_26 : IN std_logic ;
      q_arr_14_25 : IN std_logic ;
      q_arr_14_24 : IN std_logic ;
      q_arr_14_23 : IN std_logic ;
      q_arr_14_22 : IN std_logic ;
      q_arr_14_21 : IN std_logic ;
      q_arr_14_20 : IN std_logic ;
      q_arr_14_19 : IN std_logic ;
      q_arr_14_18 : IN std_logic ;
      q_arr_14_17 : IN std_logic ;
      q_arr_14_16 : IN std_logic ;
      q_arr_14_15 : IN std_logic ;
      q_arr_14_14 : IN std_logic ;
      q_arr_14_13 : IN std_logic ;
      q_arr_14_12 : IN std_logic ;
      q_arr_14_11 : IN std_logic ;
      q_arr_14_10 : IN std_logic ;
      q_arr_14_9 : IN std_logic ;
      q_arr_14_8 : IN std_logic ;
      q_arr_14_7 : IN std_logic ;
      q_arr_14_6 : IN std_logic ;
      q_arr_14_5 : IN std_logic ;
      q_arr_14_4 : IN std_logic ;
      q_arr_14_3 : IN std_logic ;
      q_arr_14_2 : IN std_logic ;
      q_arr_14_1 : IN std_logic ;
      q_arr_14_0 : IN std_logic ;
      q_arr_15_31 : IN std_logic ;
      q_arr_15_30 : IN std_logic ;
      q_arr_15_29 : IN std_logic ;
      q_arr_15_28 : IN std_logic ;
      q_arr_15_27 : IN std_logic ;
      q_arr_15_26 : IN std_logic ;
      q_arr_15_25 : IN std_logic ;
      q_arr_15_24 : IN std_logic ;
      q_arr_15_23 : IN std_logic ;
      q_arr_15_22 : IN std_logic ;
      q_arr_15_21 : IN std_logic ;
      q_arr_15_20 : IN std_logic ;
      q_arr_15_19 : IN std_logic ;
      q_arr_15_18 : IN std_logic ;
      q_arr_15_17 : IN std_logic ;
      q_arr_15_16 : IN std_logic ;
      q_arr_15_15 : IN std_logic ;
      q_arr_15_14 : IN std_logic ;
      q_arr_15_13 : IN std_logic ;
      q_arr_15_12 : IN std_logic ;
      q_arr_15_11 : IN std_logic ;
      q_arr_15_10 : IN std_logic ;
      q_arr_15_9 : IN std_logic ;
      q_arr_15_8 : IN std_logic ;
      q_arr_15_7 : IN std_logic ;
      q_arr_15_6 : IN std_logic ;
      q_arr_15_5 : IN std_logic ;
      q_arr_15_4 : IN std_logic ;
      q_arr_15_3 : IN std_logic ;
      q_arr_15_2 : IN std_logic ;
      q_arr_15_1 : IN std_logic ;
      q_arr_15_0 : IN std_logic ;
      q_arr_16_31 : IN std_logic ;
      q_arr_16_30 : IN std_logic ;
      q_arr_16_29 : IN std_logic ;
      q_arr_16_28 : IN std_logic ;
      q_arr_16_27 : IN std_logic ;
      q_arr_16_26 : IN std_logic ;
      q_arr_16_25 : IN std_logic ;
      q_arr_16_24 : IN std_logic ;
      q_arr_16_23 : IN std_logic ;
      q_arr_16_22 : IN std_logic ;
      q_arr_16_21 : IN std_logic ;
      q_arr_16_20 : IN std_logic ;
      q_arr_16_19 : IN std_logic ;
      q_arr_16_18 : IN std_logic ;
      q_arr_16_17 : IN std_logic ;
      q_arr_16_16 : IN std_logic ;
      q_arr_16_15 : IN std_logic ;
      q_arr_16_14 : IN std_logic ;
      q_arr_16_13 : IN std_logic ;
      q_arr_16_12 : IN std_logic ;
      q_arr_16_11 : IN std_logic ;
      q_arr_16_10 : IN std_logic ;
      q_arr_16_9 : IN std_logic ;
      q_arr_16_8 : IN std_logic ;
      q_arr_16_7 : IN std_logic ;
      q_arr_16_6 : IN std_logic ;
      q_arr_16_5 : IN std_logic ;
      q_arr_16_4 : IN std_logic ;
      q_arr_16_3 : IN std_logic ;
      q_arr_16_2 : IN std_logic ;
      q_arr_16_1 : IN std_logic ;
      q_arr_16_0 : IN std_logic ;
      q_arr_17_31 : IN std_logic ;
      q_arr_17_30 : IN std_logic ;
      q_arr_17_29 : IN std_logic ;
      q_arr_17_28 : IN std_logic ;
      q_arr_17_27 : IN std_logic ;
      q_arr_17_26 : IN std_logic ;
      q_arr_17_25 : IN std_logic ;
      q_arr_17_24 : IN std_logic ;
      q_arr_17_23 : IN std_logic ;
      q_arr_17_22 : IN std_logic ;
      q_arr_17_21 : IN std_logic ;
      q_arr_17_20 : IN std_logic ;
      q_arr_17_19 : IN std_logic ;
      q_arr_17_18 : IN std_logic ;
      q_arr_17_17 : IN std_logic ;
      q_arr_17_16 : IN std_logic ;
      q_arr_17_15 : IN std_logic ;
      q_arr_17_14 : IN std_logic ;
      q_arr_17_13 : IN std_logic ;
      q_arr_17_12 : IN std_logic ;
      q_arr_17_11 : IN std_logic ;
      q_arr_17_10 : IN std_logic ;
      q_arr_17_9 : IN std_logic ;
      q_arr_17_8 : IN std_logic ;
      q_arr_17_7 : IN std_logic ;
      q_arr_17_6 : IN std_logic ;
      q_arr_17_5 : IN std_logic ;
      q_arr_17_4 : IN std_logic ;
      q_arr_17_3 : IN std_logic ;
      q_arr_17_2 : IN std_logic ;
      q_arr_17_1 : IN std_logic ;
      q_arr_17_0 : IN std_logic ;
      q_arr_18_31 : IN std_logic ;
      q_arr_18_30 : IN std_logic ;
      q_arr_18_29 : IN std_logic ;
      q_arr_18_28 : IN std_logic ;
      q_arr_18_27 : IN std_logic ;
      q_arr_18_26 : IN std_logic ;
      q_arr_18_25 : IN std_logic ;
      q_arr_18_24 : IN std_logic ;
      q_arr_18_23 : IN std_logic ;
      q_arr_18_22 : IN std_logic ;
      q_arr_18_21 : IN std_logic ;
      q_arr_18_20 : IN std_logic ;
      q_arr_18_19 : IN std_logic ;
      q_arr_18_18 : IN std_logic ;
      q_arr_18_17 : IN std_logic ;
      q_arr_18_16 : IN std_logic ;
      q_arr_18_15 : IN std_logic ;
      q_arr_18_14 : IN std_logic ;
      q_arr_18_13 : IN std_logic ;
      q_arr_18_12 : IN std_logic ;
      q_arr_18_11 : IN std_logic ;
      q_arr_18_10 : IN std_logic ;
      q_arr_18_9 : IN std_logic ;
      q_arr_18_8 : IN std_logic ;
      q_arr_18_7 : IN std_logic ;
      q_arr_18_6 : IN std_logic ;
      q_arr_18_5 : IN std_logic ;
      q_arr_18_4 : IN std_logic ;
      q_arr_18_3 : IN std_logic ;
      q_arr_18_2 : IN std_logic ;
      q_arr_18_1 : IN std_logic ;
      q_arr_18_0 : IN std_logic ;
      q_arr_19_31 : IN std_logic ;
      q_arr_19_30 : IN std_logic ;
      q_arr_19_29 : IN std_logic ;
      q_arr_19_28 : IN std_logic ;
      q_arr_19_27 : IN std_logic ;
      q_arr_19_26 : IN std_logic ;
      q_arr_19_25 : IN std_logic ;
      q_arr_19_24 : IN std_logic ;
      q_arr_19_23 : IN std_logic ;
      q_arr_19_22 : IN std_logic ;
      q_arr_19_21 : IN std_logic ;
      q_arr_19_20 : IN std_logic ;
      q_arr_19_19 : IN std_logic ;
      q_arr_19_18 : IN std_logic ;
      q_arr_19_17 : IN std_logic ;
      q_arr_19_16 : IN std_logic ;
      q_arr_19_15 : IN std_logic ;
      q_arr_19_14 : IN std_logic ;
      q_arr_19_13 : IN std_logic ;
      q_arr_19_12 : IN std_logic ;
      q_arr_19_11 : IN std_logic ;
      q_arr_19_10 : IN std_logic ;
      q_arr_19_9 : IN std_logic ;
      q_arr_19_8 : IN std_logic ;
      q_arr_19_7 : IN std_logic ;
      q_arr_19_6 : IN std_logic ;
      q_arr_19_5 : IN std_logic ;
      q_arr_19_4 : IN std_logic ;
      q_arr_19_3 : IN std_logic ;
      q_arr_19_2 : IN std_logic ;
      q_arr_19_1 : IN std_logic ;
      q_arr_19_0 : IN std_logic ;
      q_arr_20_31 : IN std_logic ;
      q_arr_20_30 : IN std_logic ;
      q_arr_20_29 : IN std_logic ;
      q_arr_20_28 : IN std_logic ;
      q_arr_20_27 : IN std_logic ;
      q_arr_20_26 : IN std_logic ;
      q_arr_20_25 : IN std_logic ;
      q_arr_20_24 : IN std_logic ;
      q_arr_20_23 : IN std_logic ;
      q_arr_20_22 : IN std_logic ;
      q_arr_20_21 : IN std_logic ;
      q_arr_20_20 : IN std_logic ;
      q_arr_20_19 : IN std_logic ;
      q_arr_20_18 : IN std_logic ;
      q_arr_20_17 : IN std_logic ;
      q_arr_20_16 : IN std_logic ;
      q_arr_20_15 : IN std_logic ;
      q_arr_20_14 : IN std_logic ;
      q_arr_20_13 : IN std_logic ;
      q_arr_20_12 : IN std_logic ;
      q_arr_20_11 : IN std_logic ;
      q_arr_20_10 : IN std_logic ;
      q_arr_20_9 : IN std_logic ;
      q_arr_20_8 : IN std_logic ;
      q_arr_20_7 : IN std_logic ;
      q_arr_20_6 : IN std_logic ;
      q_arr_20_5 : IN std_logic ;
      q_arr_20_4 : IN std_logic ;
      q_arr_20_3 : IN std_logic ;
      q_arr_20_2 : IN std_logic ;
      q_arr_20_1 : IN std_logic ;
      q_arr_20_0 : IN std_logic ;
      q_arr_21_31 : IN std_logic ;
      q_arr_21_30 : IN std_logic ;
      q_arr_21_29 : IN std_logic ;
      q_arr_21_28 : IN std_logic ;
      q_arr_21_27 : IN std_logic ;
      q_arr_21_26 : IN std_logic ;
      q_arr_21_25 : IN std_logic ;
      q_arr_21_24 : IN std_logic ;
      q_arr_21_23 : IN std_logic ;
      q_arr_21_22 : IN std_logic ;
      q_arr_21_21 : IN std_logic ;
      q_arr_21_20 : IN std_logic ;
      q_arr_21_19 : IN std_logic ;
      q_arr_21_18 : IN std_logic ;
      q_arr_21_17 : IN std_logic ;
      q_arr_21_16 : IN std_logic ;
      q_arr_21_15 : IN std_logic ;
      q_arr_21_14 : IN std_logic ;
      q_arr_21_13 : IN std_logic ;
      q_arr_21_12 : IN std_logic ;
      q_arr_21_11 : IN std_logic ;
      q_arr_21_10 : IN std_logic ;
      q_arr_21_9 : IN std_logic ;
      q_arr_21_8 : IN std_logic ;
      q_arr_21_7 : IN std_logic ;
      q_arr_21_6 : IN std_logic ;
      q_arr_21_5 : IN std_logic ;
      q_arr_21_4 : IN std_logic ;
      q_arr_21_3 : IN std_logic ;
      q_arr_21_2 : IN std_logic ;
      q_arr_21_1 : IN std_logic ;
      q_arr_21_0 : IN std_logic ;
      q_arr_22_31 : IN std_logic ;
      q_arr_22_30 : IN std_logic ;
      q_arr_22_29 : IN std_logic ;
      q_arr_22_28 : IN std_logic ;
      q_arr_22_27 : IN std_logic ;
      q_arr_22_26 : IN std_logic ;
      q_arr_22_25 : IN std_logic ;
      q_arr_22_24 : IN std_logic ;
      q_arr_22_23 : IN std_logic ;
      q_arr_22_22 : IN std_logic ;
      q_arr_22_21 : IN std_logic ;
      q_arr_22_20 : IN std_logic ;
      q_arr_22_19 : IN std_logic ;
      q_arr_22_18 : IN std_logic ;
      q_arr_22_17 : IN std_logic ;
      q_arr_22_16 : IN std_logic ;
      q_arr_22_15 : IN std_logic ;
      q_arr_22_14 : IN std_logic ;
      q_arr_22_13 : IN std_logic ;
      q_arr_22_12 : IN std_logic ;
      q_arr_22_11 : IN std_logic ;
      q_arr_22_10 : IN std_logic ;
      q_arr_22_9 : IN std_logic ;
      q_arr_22_8 : IN std_logic ;
      q_arr_22_7 : IN std_logic ;
      q_arr_22_6 : IN std_logic ;
      q_arr_22_5 : IN std_logic ;
      q_arr_22_4 : IN std_logic ;
      q_arr_22_3 : IN std_logic ;
      q_arr_22_2 : IN std_logic ;
      q_arr_22_1 : IN std_logic ;
      q_arr_22_0 : IN std_logic ;
      q_arr_23_31 : IN std_logic ;
      q_arr_23_30 : IN std_logic ;
      q_arr_23_29 : IN std_logic ;
      q_arr_23_28 : IN std_logic ;
      q_arr_23_27 : IN std_logic ;
      q_arr_23_26 : IN std_logic ;
      q_arr_23_25 : IN std_logic ;
      q_arr_23_24 : IN std_logic ;
      q_arr_23_23 : IN std_logic ;
      q_arr_23_22 : IN std_logic ;
      q_arr_23_21 : IN std_logic ;
      q_arr_23_20 : IN std_logic ;
      q_arr_23_19 : IN std_logic ;
      q_arr_23_18 : IN std_logic ;
      q_arr_23_17 : IN std_logic ;
      q_arr_23_16 : IN std_logic ;
      q_arr_23_15 : IN std_logic ;
      q_arr_23_14 : IN std_logic ;
      q_arr_23_13 : IN std_logic ;
      q_arr_23_12 : IN std_logic ;
      q_arr_23_11 : IN std_logic ;
      q_arr_23_10 : IN std_logic ;
      q_arr_23_9 : IN std_logic ;
      q_arr_23_8 : IN std_logic ;
      q_arr_23_7 : IN std_logic ;
      q_arr_23_6 : IN std_logic ;
      q_arr_23_5 : IN std_logic ;
      q_arr_23_4 : IN std_logic ;
      q_arr_23_3 : IN std_logic ;
      q_arr_23_2 : IN std_logic ;
      q_arr_23_1 : IN std_logic ;
      q_arr_23_0 : IN std_logic ;
      q_arr_24_31 : IN std_logic ;
      q_arr_24_30 : IN std_logic ;
      q_arr_24_29 : IN std_logic ;
      q_arr_24_28 : IN std_logic ;
      q_arr_24_27 : IN std_logic ;
      q_arr_24_26 : IN std_logic ;
      q_arr_24_25 : IN std_logic ;
      q_arr_24_24 : IN std_logic ;
      q_arr_24_23 : IN std_logic ;
      q_arr_24_22 : IN std_logic ;
      q_arr_24_21 : IN std_logic ;
      q_arr_24_20 : IN std_logic ;
      q_arr_24_19 : IN std_logic ;
      q_arr_24_18 : IN std_logic ;
      q_arr_24_17 : IN std_logic ;
      q_arr_24_16 : IN std_logic ;
      q_arr_24_15 : IN std_logic ;
      q_arr_24_14 : IN std_logic ;
      q_arr_24_13 : IN std_logic ;
      q_arr_24_12 : IN std_logic ;
      q_arr_24_11 : IN std_logic ;
      q_arr_24_10 : IN std_logic ;
      q_arr_24_9 : IN std_logic ;
      q_arr_24_8 : IN std_logic ;
      q_arr_24_7 : IN std_logic ;
      q_arr_24_6 : IN std_logic ;
      q_arr_24_5 : IN std_logic ;
      q_arr_24_4 : IN std_logic ;
      q_arr_24_3 : IN std_logic ;
      q_arr_24_2 : IN std_logic ;
      q_arr_24_1 : IN std_logic ;
      q_arr_24_0 : IN std_logic ;
      output1_init : IN std_logic_vector (15 DOWNTO 0) ;
      output2_init : IN std_logic_vector (15 DOWNTO 0) ;
      filter_size : IN std_logic ;
      operation : IN std_logic ;
      compute_relu : IN std_logic ;
      clk : IN std_logic ;
      en : IN std_logic ;
      reset : IN std_logic ;
      buffer_ready : OUT std_logic ;
      semi_ready : OUT std_logic ;
      ready : OUT std_logic) ;
end ComputationPipeline ;

architecture Behavioral of ComputationPipeline is
   component CacheMuxer
      port (
         d_arr_mux_0_31 : IN std_logic ;
         d_arr_mux_0_30 : IN std_logic ;
         d_arr_mux_0_29 : IN std_logic ;
         d_arr_mux_0_28 : IN std_logic ;
         d_arr_mux_0_27 : IN std_logic ;
         d_arr_mux_0_26 : IN std_logic ;
         d_arr_mux_0_25 : IN std_logic ;
         d_arr_mux_0_24 : IN std_logic ;
         d_arr_mux_0_23 : IN std_logic ;
         d_arr_mux_0_22 : IN std_logic ;
         d_arr_mux_0_21 : IN std_logic ;
         d_arr_mux_0_20 : IN std_logic ;
         d_arr_mux_0_19 : IN std_logic ;
         d_arr_mux_0_18 : IN std_logic ;
         d_arr_mux_0_17 : IN std_logic ;
         d_arr_mux_0_16 : IN std_logic ;
         d_arr_mux_0_15 : IN std_logic ;
         d_arr_mux_0_14 : IN std_logic ;
         d_arr_mux_0_13 : IN std_logic ;
         d_arr_mux_0_12 : IN std_logic ;
         d_arr_mux_0_11 : IN std_logic ;
         d_arr_mux_0_10 : IN std_logic ;
         d_arr_mux_0_9 : IN std_logic ;
         d_arr_mux_0_8 : IN std_logic ;
         d_arr_mux_0_7 : IN std_logic ;
         d_arr_mux_0_6 : IN std_logic ;
         d_arr_mux_0_5 : IN std_logic ;
         d_arr_mux_0_4 : IN std_logic ;
         d_arr_mux_0_3 : IN std_logic ;
         d_arr_mux_0_2 : IN std_logic ;
         d_arr_mux_0_1 : IN std_logic ;
         d_arr_mux_0_0 : IN std_logic ;
         d_arr_mux_1_31 : IN std_logic ;
         d_arr_mux_1_30 : IN std_logic ;
         d_arr_mux_1_29 : IN std_logic ;
         d_arr_mux_1_28 : IN std_logic ;
         d_arr_mux_1_27 : IN std_logic ;
         d_arr_mux_1_26 : IN std_logic ;
         d_arr_mux_1_25 : IN std_logic ;
         d_arr_mux_1_24 : IN std_logic ;
         d_arr_mux_1_23 : IN std_logic ;
         d_arr_mux_1_22 : IN std_logic ;
         d_arr_mux_1_21 : IN std_logic ;
         d_arr_mux_1_20 : IN std_logic ;
         d_arr_mux_1_19 : IN std_logic ;
         d_arr_mux_1_18 : IN std_logic ;
         d_arr_mux_1_17 : IN std_logic ;
         d_arr_mux_1_16 : IN std_logic ;
         d_arr_mux_1_15 : IN std_logic ;
         d_arr_mux_1_14 : IN std_logic ;
         d_arr_mux_1_13 : IN std_logic ;
         d_arr_mux_1_12 : IN std_logic ;
         d_arr_mux_1_11 : IN std_logic ;
         d_arr_mux_1_10 : IN std_logic ;
         d_arr_mux_1_9 : IN std_logic ;
         d_arr_mux_1_8 : IN std_logic ;
         d_arr_mux_1_7 : IN std_logic ;
         d_arr_mux_1_6 : IN std_logic ;
         d_arr_mux_1_5 : IN std_logic ;
         d_arr_mux_1_4 : IN std_logic ;
         d_arr_mux_1_3 : IN std_logic ;
         d_arr_mux_1_2 : IN std_logic ;
         d_arr_mux_1_1 : IN std_logic ;
         d_arr_mux_1_0 : IN std_logic ;
         d_arr_mux_2_31 : IN std_logic ;
         d_arr_mux_2_30 : IN std_logic ;
         d_arr_mux_2_29 : IN std_logic ;
         d_arr_mux_2_28 : IN std_logic ;
         d_arr_mux_2_27 : IN std_logic ;
         d_arr_mux_2_26 : IN std_logic ;
         d_arr_mux_2_25 : IN std_logic ;
         d_arr_mux_2_24 : IN std_logic ;
         d_arr_mux_2_23 : IN std_logic ;
         d_arr_mux_2_22 : IN std_logic ;
         d_arr_mux_2_21 : IN std_logic ;
         d_arr_mux_2_20 : IN std_logic ;
         d_arr_mux_2_19 : IN std_logic ;
         d_arr_mux_2_18 : IN std_logic ;
         d_arr_mux_2_17 : IN std_logic ;
         d_arr_mux_2_16 : IN std_logic ;
         d_arr_mux_2_15 : IN std_logic ;
         d_arr_mux_2_14 : IN std_logic ;
         d_arr_mux_2_13 : IN std_logic ;
         d_arr_mux_2_12 : IN std_logic ;
         d_arr_mux_2_11 : IN std_logic ;
         d_arr_mux_2_10 : IN std_logic ;
         d_arr_mux_2_9 : IN std_logic ;
         d_arr_mux_2_8 : IN std_logic ;
         d_arr_mux_2_7 : IN std_logic ;
         d_arr_mux_2_6 : IN std_logic ;
         d_arr_mux_2_5 : IN std_logic ;
         d_arr_mux_2_4 : IN std_logic ;
         d_arr_mux_2_3 : IN std_logic ;
         d_arr_mux_2_2 : IN std_logic ;
         d_arr_mux_2_1 : IN std_logic ;
         d_arr_mux_2_0 : IN std_logic ;
         d_arr_mux_3_31 : IN std_logic ;
         d_arr_mux_3_30 : IN std_logic ;
         d_arr_mux_3_29 : IN std_logic ;
         d_arr_mux_3_28 : IN std_logic ;
         d_arr_mux_3_27 : IN std_logic ;
         d_arr_mux_3_26 : IN std_logic ;
         d_arr_mux_3_25 : IN std_logic ;
         d_arr_mux_3_24 : IN std_logic ;
         d_arr_mux_3_23 : IN std_logic ;
         d_arr_mux_3_22 : IN std_logic ;
         d_arr_mux_3_21 : IN std_logic ;
         d_arr_mux_3_20 : IN std_logic ;
         d_arr_mux_3_19 : IN std_logic ;
         d_arr_mux_3_18 : IN std_logic ;
         d_arr_mux_3_17 : IN std_logic ;
         d_arr_mux_3_16 : IN std_logic ;
         d_arr_mux_3_15 : IN std_logic ;
         d_arr_mux_3_14 : IN std_logic ;
         d_arr_mux_3_13 : IN std_logic ;
         d_arr_mux_3_12 : IN std_logic ;
         d_arr_mux_3_11 : IN std_logic ;
         d_arr_mux_3_10 : IN std_logic ;
         d_arr_mux_3_9 : IN std_logic ;
         d_arr_mux_3_8 : IN std_logic ;
         d_arr_mux_3_7 : IN std_logic ;
         d_arr_mux_3_6 : IN std_logic ;
         d_arr_mux_3_5 : IN std_logic ;
         d_arr_mux_3_4 : IN std_logic ;
         d_arr_mux_3_3 : IN std_logic ;
         d_arr_mux_3_2 : IN std_logic ;
         d_arr_mux_3_1 : IN std_logic ;
         d_arr_mux_3_0 : IN std_logic ;
         d_arr_mux_4_31 : IN std_logic ;
         d_arr_mux_4_30 : IN std_logic ;
         d_arr_mux_4_29 : IN std_logic ;
         d_arr_mux_4_28 : IN std_logic ;
         d_arr_mux_4_27 : IN std_logic ;
         d_arr_mux_4_26 : IN std_logic ;
         d_arr_mux_4_25 : IN std_logic ;
         d_arr_mux_4_24 : IN std_logic ;
         d_arr_mux_4_23 : IN std_logic ;
         d_arr_mux_4_22 : IN std_logic ;
         d_arr_mux_4_21 : IN std_logic ;
         d_arr_mux_4_20 : IN std_logic ;
         d_arr_mux_4_19 : IN std_logic ;
         d_arr_mux_4_18 : IN std_logic ;
         d_arr_mux_4_17 : IN std_logic ;
         d_arr_mux_4_16 : IN std_logic ;
         d_arr_mux_4_15 : IN std_logic ;
         d_arr_mux_4_14 : IN std_logic ;
         d_arr_mux_4_13 : IN std_logic ;
         d_arr_mux_4_12 : IN std_logic ;
         d_arr_mux_4_11 : IN std_logic ;
         d_arr_mux_4_10 : IN std_logic ;
         d_arr_mux_4_9 : IN std_logic ;
         d_arr_mux_4_8 : IN std_logic ;
         d_arr_mux_4_7 : IN std_logic ;
         d_arr_mux_4_6 : IN std_logic ;
         d_arr_mux_4_5 : IN std_logic ;
         d_arr_mux_4_4 : IN std_logic ;
         d_arr_mux_4_3 : IN std_logic ;
         d_arr_mux_4_2 : IN std_logic ;
         d_arr_mux_4_1 : IN std_logic ;
         d_arr_mux_4_0 : IN std_logic ;
         d_arr_mux_5_31 : IN std_logic ;
         d_arr_mux_5_30 : IN std_logic ;
         d_arr_mux_5_29 : IN std_logic ;
         d_arr_mux_5_28 : IN std_logic ;
         d_arr_mux_5_27 : IN std_logic ;
         d_arr_mux_5_26 : IN std_logic ;
         d_arr_mux_5_25 : IN std_logic ;
         d_arr_mux_5_24 : IN std_logic ;
         d_arr_mux_5_23 : IN std_logic ;
         d_arr_mux_5_22 : IN std_logic ;
         d_arr_mux_5_21 : IN std_logic ;
         d_arr_mux_5_20 : IN std_logic ;
         d_arr_mux_5_19 : IN std_logic ;
         d_arr_mux_5_18 : IN std_logic ;
         d_arr_mux_5_17 : IN std_logic ;
         d_arr_mux_5_16 : IN std_logic ;
         d_arr_mux_5_15 : IN std_logic ;
         d_arr_mux_5_14 : IN std_logic ;
         d_arr_mux_5_13 : IN std_logic ;
         d_arr_mux_5_12 : IN std_logic ;
         d_arr_mux_5_11 : IN std_logic ;
         d_arr_mux_5_10 : IN std_logic ;
         d_arr_mux_5_9 : IN std_logic ;
         d_arr_mux_5_8 : IN std_logic ;
         d_arr_mux_5_7 : IN std_logic ;
         d_arr_mux_5_6 : IN std_logic ;
         d_arr_mux_5_5 : IN std_logic ;
         d_arr_mux_5_4 : IN std_logic ;
         d_arr_mux_5_3 : IN std_logic ;
         d_arr_mux_5_2 : IN std_logic ;
         d_arr_mux_5_1 : IN std_logic ;
         d_arr_mux_5_0 : IN std_logic ;
         d_arr_mux_6_31 : IN std_logic ;
         d_arr_mux_6_30 : IN std_logic ;
         d_arr_mux_6_29 : IN std_logic ;
         d_arr_mux_6_28 : IN std_logic ;
         d_arr_mux_6_27 : IN std_logic ;
         d_arr_mux_6_26 : IN std_logic ;
         d_arr_mux_6_25 : IN std_logic ;
         d_arr_mux_6_24 : IN std_logic ;
         d_arr_mux_6_23 : IN std_logic ;
         d_arr_mux_6_22 : IN std_logic ;
         d_arr_mux_6_21 : IN std_logic ;
         d_arr_mux_6_20 : IN std_logic ;
         d_arr_mux_6_19 : IN std_logic ;
         d_arr_mux_6_18 : IN std_logic ;
         d_arr_mux_6_17 : IN std_logic ;
         d_arr_mux_6_16 : IN std_logic ;
         d_arr_mux_6_15 : IN std_logic ;
         d_arr_mux_6_14 : IN std_logic ;
         d_arr_mux_6_13 : IN std_logic ;
         d_arr_mux_6_12 : IN std_logic ;
         d_arr_mux_6_11 : IN std_logic ;
         d_arr_mux_6_10 : IN std_logic ;
         d_arr_mux_6_9 : IN std_logic ;
         d_arr_mux_6_8 : IN std_logic ;
         d_arr_mux_6_7 : IN std_logic ;
         d_arr_mux_6_6 : IN std_logic ;
         d_arr_mux_6_5 : IN std_logic ;
         d_arr_mux_6_4 : IN std_logic ;
         d_arr_mux_6_3 : IN std_logic ;
         d_arr_mux_6_2 : IN std_logic ;
         d_arr_mux_6_1 : IN std_logic ;
         d_arr_mux_6_0 : IN std_logic ;
         d_arr_mux_7_31 : IN std_logic ;
         d_arr_mux_7_30 : IN std_logic ;
         d_arr_mux_7_29 : IN std_logic ;
         d_arr_mux_7_28 : IN std_logic ;
         d_arr_mux_7_27 : IN std_logic ;
         d_arr_mux_7_26 : IN std_logic ;
         d_arr_mux_7_25 : IN std_logic ;
         d_arr_mux_7_24 : IN std_logic ;
         d_arr_mux_7_23 : IN std_logic ;
         d_arr_mux_7_22 : IN std_logic ;
         d_arr_mux_7_21 : IN std_logic ;
         d_arr_mux_7_20 : IN std_logic ;
         d_arr_mux_7_19 : IN std_logic ;
         d_arr_mux_7_18 : IN std_logic ;
         d_arr_mux_7_17 : IN std_logic ;
         d_arr_mux_7_16 : IN std_logic ;
         d_arr_mux_7_15 : IN std_logic ;
         d_arr_mux_7_14 : IN std_logic ;
         d_arr_mux_7_13 : IN std_logic ;
         d_arr_mux_7_12 : IN std_logic ;
         d_arr_mux_7_11 : IN std_logic ;
         d_arr_mux_7_10 : IN std_logic ;
         d_arr_mux_7_9 : IN std_logic ;
         d_arr_mux_7_8 : IN std_logic ;
         d_arr_mux_7_7 : IN std_logic ;
         d_arr_mux_7_6 : IN std_logic ;
         d_arr_mux_7_5 : IN std_logic ;
         d_arr_mux_7_4 : IN std_logic ;
         d_arr_mux_7_3 : IN std_logic ;
         d_arr_mux_7_2 : IN std_logic ;
         d_arr_mux_7_1 : IN std_logic ;
         d_arr_mux_7_0 : IN std_logic ;
         d_arr_mux_8_31 : IN std_logic ;
         d_arr_mux_8_30 : IN std_logic ;
         d_arr_mux_8_29 : IN std_logic ;
         d_arr_mux_8_28 : IN std_logic ;
         d_arr_mux_8_27 : IN std_logic ;
         d_arr_mux_8_26 : IN std_logic ;
         d_arr_mux_8_25 : IN std_logic ;
         d_arr_mux_8_24 : IN std_logic ;
         d_arr_mux_8_23 : IN std_logic ;
         d_arr_mux_8_22 : IN std_logic ;
         d_arr_mux_8_21 : IN std_logic ;
         d_arr_mux_8_20 : IN std_logic ;
         d_arr_mux_8_19 : IN std_logic ;
         d_arr_mux_8_18 : IN std_logic ;
         d_arr_mux_8_17 : IN std_logic ;
         d_arr_mux_8_16 : IN std_logic ;
         d_arr_mux_8_15 : IN std_logic ;
         d_arr_mux_8_14 : IN std_logic ;
         d_arr_mux_8_13 : IN std_logic ;
         d_arr_mux_8_12 : IN std_logic ;
         d_arr_mux_8_11 : IN std_logic ;
         d_arr_mux_8_10 : IN std_logic ;
         d_arr_mux_8_9 : IN std_logic ;
         d_arr_mux_8_8 : IN std_logic ;
         d_arr_mux_8_7 : IN std_logic ;
         d_arr_mux_8_6 : IN std_logic ;
         d_arr_mux_8_5 : IN std_logic ;
         d_arr_mux_8_4 : IN std_logic ;
         d_arr_mux_8_3 : IN std_logic ;
         d_arr_mux_8_2 : IN std_logic ;
         d_arr_mux_8_1 : IN std_logic ;
         d_arr_mux_8_0 : IN std_logic ;
         d_arr_mux_9_31 : IN std_logic ;
         d_arr_mux_9_30 : IN std_logic ;
         d_arr_mux_9_29 : IN std_logic ;
         d_arr_mux_9_28 : IN std_logic ;
         d_arr_mux_9_27 : IN std_logic ;
         d_arr_mux_9_26 : IN std_logic ;
         d_arr_mux_9_25 : IN std_logic ;
         d_arr_mux_9_24 : IN std_logic ;
         d_arr_mux_9_23 : IN std_logic ;
         d_arr_mux_9_22 : IN std_logic ;
         d_arr_mux_9_21 : IN std_logic ;
         d_arr_mux_9_20 : IN std_logic ;
         d_arr_mux_9_19 : IN std_logic ;
         d_arr_mux_9_18 : IN std_logic ;
         d_arr_mux_9_17 : IN std_logic ;
         d_arr_mux_9_16 : IN std_logic ;
         d_arr_mux_9_15 : IN std_logic ;
         d_arr_mux_9_14 : IN std_logic ;
         d_arr_mux_9_13 : IN std_logic ;
         d_arr_mux_9_12 : IN std_logic ;
         d_arr_mux_9_11 : IN std_logic ;
         d_arr_mux_9_10 : IN std_logic ;
         d_arr_mux_9_9 : IN std_logic ;
         d_arr_mux_9_8 : IN std_logic ;
         d_arr_mux_9_7 : IN std_logic ;
         d_arr_mux_9_6 : IN std_logic ;
         d_arr_mux_9_5 : IN std_logic ;
         d_arr_mux_9_4 : IN std_logic ;
         d_arr_mux_9_3 : IN std_logic ;
         d_arr_mux_9_2 : IN std_logic ;
         d_arr_mux_9_1 : IN std_logic ;
         d_arr_mux_9_0 : IN std_logic ;
         d_arr_mux_10_31 : IN std_logic ;
         d_arr_mux_10_30 : IN std_logic ;
         d_arr_mux_10_29 : IN std_logic ;
         d_arr_mux_10_28 : IN std_logic ;
         d_arr_mux_10_27 : IN std_logic ;
         d_arr_mux_10_26 : IN std_logic ;
         d_arr_mux_10_25 : IN std_logic ;
         d_arr_mux_10_24 : IN std_logic ;
         d_arr_mux_10_23 : IN std_logic ;
         d_arr_mux_10_22 : IN std_logic ;
         d_arr_mux_10_21 : IN std_logic ;
         d_arr_mux_10_20 : IN std_logic ;
         d_arr_mux_10_19 : IN std_logic ;
         d_arr_mux_10_18 : IN std_logic ;
         d_arr_mux_10_17 : IN std_logic ;
         d_arr_mux_10_16 : IN std_logic ;
         d_arr_mux_10_15 : IN std_logic ;
         d_arr_mux_10_14 : IN std_logic ;
         d_arr_mux_10_13 : IN std_logic ;
         d_arr_mux_10_12 : IN std_logic ;
         d_arr_mux_10_11 : IN std_logic ;
         d_arr_mux_10_10 : IN std_logic ;
         d_arr_mux_10_9 : IN std_logic ;
         d_arr_mux_10_8 : IN std_logic ;
         d_arr_mux_10_7 : IN std_logic ;
         d_arr_mux_10_6 : IN std_logic ;
         d_arr_mux_10_5 : IN std_logic ;
         d_arr_mux_10_4 : IN std_logic ;
         d_arr_mux_10_3 : IN std_logic ;
         d_arr_mux_10_2 : IN std_logic ;
         d_arr_mux_10_1 : IN std_logic ;
         d_arr_mux_10_0 : IN std_logic ;
         d_arr_mux_11_31 : IN std_logic ;
         d_arr_mux_11_30 : IN std_logic ;
         d_arr_mux_11_29 : IN std_logic ;
         d_arr_mux_11_28 : IN std_logic ;
         d_arr_mux_11_27 : IN std_logic ;
         d_arr_mux_11_26 : IN std_logic ;
         d_arr_mux_11_25 : IN std_logic ;
         d_arr_mux_11_24 : IN std_logic ;
         d_arr_mux_11_23 : IN std_logic ;
         d_arr_mux_11_22 : IN std_logic ;
         d_arr_mux_11_21 : IN std_logic ;
         d_arr_mux_11_20 : IN std_logic ;
         d_arr_mux_11_19 : IN std_logic ;
         d_arr_mux_11_18 : IN std_logic ;
         d_arr_mux_11_17 : IN std_logic ;
         d_arr_mux_11_16 : IN std_logic ;
         d_arr_mux_11_15 : IN std_logic ;
         d_arr_mux_11_14 : IN std_logic ;
         d_arr_mux_11_13 : IN std_logic ;
         d_arr_mux_11_12 : IN std_logic ;
         d_arr_mux_11_11 : IN std_logic ;
         d_arr_mux_11_10 : IN std_logic ;
         d_arr_mux_11_9 : IN std_logic ;
         d_arr_mux_11_8 : IN std_logic ;
         d_arr_mux_11_7 : IN std_logic ;
         d_arr_mux_11_6 : IN std_logic ;
         d_arr_mux_11_5 : IN std_logic ;
         d_arr_mux_11_4 : IN std_logic ;
         d_arr_mux_11_3 : IN std_logic ;
         d_arr_mux_11_2 : IN std_logic ;
         d_arr_mux_11_1 : IN std_logic ;
         d_arr_mux_11_0 : IN std_logic ;
         d_arr_mux_12_31 : IN std_logic ;
         d_arr_mux_12_30 : IN std_logic ;
         d_arr_mux_12_29 : IN std_logic ;
         d_arr_mux_12_28 : IN std_logic ;
         d_arr_mux_12_27 : IN std_logic ;
         d_arr_mux_12_26 : IN std_logic ;
         d_arr_mux_12_25 : IN std_logic ;
         d_arr_mux_12_24 : IN std_logic ;
         d_arr_mux_12_23 : IN std_logic ;
         d_arr_mux_12_22 : IN std_logic ;
         d_arr_mux_12_21 : IN std_logic ;
         d_arr_mux_12_20 : IN std_logic ;
         d_arr_mux_12_19 : IN std_logic ;
         d_arr_mux_12_18 : IN std_logic ;
         d_arr_mux_12_17 : IN std_logic ;
         d_arr_mux_12_16 : IN std_logic ;
         d_arr_mux_12_15 : IN std_logic ;
         d_arr_mux_12_14 : IN std_logic ;
         d_arr_mux_12_13 : IN std_logic ;
         d_arr_mux_12_12 : IN std_logic ;
         d_arr_mux_12_11 : IN std_logic ;
         d_arr_mux_12_10 : IN std_logic ;
         d_arr_mux_12_9 : IN std_logic ;
         d_arr_mux_12_8 : IN std_logic ;
         d_arr_mux_12_7 : IN std_logic ;
         d_arr_mux_12_6 : IN std_logic ;
         d_arr_mux_12_5 : IN std_logic ;
         d_arr_mux_12_4 : IN std_logic ;
         d_arr_mux_12_3 : IN std_logic ;
         d_arr_mux_12_2 : IN std_logic ;
         d_arr_mux_12_1 : IN std_logic ;
         d_arr_mux_12_0 : IN std_logic ;
         d_arr_mux_13_31 : IN std_logic ;
         d_arr_mux_13_30 : IN std_logic ;
         d_arr_mux_13_29 : IN std_logic ;
         d_arr_mux_13_28 : IN std_logic ;
         d_arr_mux_13_27 : IN std_logic ;
         d_arr_mux_13_26 : IN std_logic ;
         d_arr_mux_13_25 : IN std_logic ;
         d_arr_mux_13_24 : IN std_logic ;
         d_arr_mux_13_23 : IN std_logic ;
         d_arr_mux_13_22 : IN std_logic ;
         d_arr_mux_13_21 : IN std_logic ;
         d_arr_mux_13_20 : IN std_logic ;
         d_arr_mux_13_19 : IN std_logic ;
         d_arr_mux_13_18 : IN std_logic ;
         d_arr_mux_13_17 : IN std_logic ;
         d_arr_mux_13_16 : IN std_logic ;
         d_arr_mux_13_15 : IN std_logic ;
         d_arr_mux_13_14 : IN std_logic ;
         d_arr_mux_13_13 : IN std_logic ;
         d_arr_mux_13_12 : IN std_logic ;
         d_arr_mux_13_11 : IN std_logic ;
         d_arr_mux_13_10 : IN std_logic ;
         d_arr_mux_13_9 : IN std_logic ;
         d_arr_mux_13_8 : IN std_logic ;
         d_arr_mux_13_7 : IN std_logic ;
         d_arr_mux_13_6 : IN std_logic ;
         d_arr_mux_13_5 : IN std_logic ;
         d_arr_mux_13_4 : IN std_logic ;
         d_arr_mux_13_3 : IN std_logic ;
         d_arr_mux_13_2 : IN std_logic ;
         d_arr_mux_13_1 : IN std_logic ;
         d_arr_mux_13_0 : IN std_logic ;
         d_arr_mux_14_31 : IN std_logic ;
         d_arr_mux_14_30 : IN std_logic ;
         d_arr_mux_14_29 : IN std_logic ;
         d_arr_mux_14_28 : IN std_logic ;
         d_arr_mux_14_27 : IN std_logic ;
         d_arr_mux_14_26 : IN std_logic ;
         d_arr_mux_14_25 : IN std_logic ;
         d_arr_mux_14_24 : IN std_logic ;
         d_arr_mux_14_23 : IN std_logic ;
         d_arr_mux_14_22 : IN std_logic ;
         d_arr_mux_14_21 : IN std_logic ;
         d_arr_mux_14_20 : IN std_logic ;
         d_arr_mux_14_19 : IN std_logic ;
         d_arr_mux_14_18 : IN std_logic ;
         d_arr_mux_14_17 : IN std_logic ;
         d_arr_mux_14_16 : IN std_logic ;
         d_arr_mux_14_15 : IN std_logic ;
         d_arr_mux_14_14 : IN std_logic ;
         d_arr_mux_14_13 : IN std_logic ;
         d_arr_mux_14_12 : IN std_logic ;
         d_arr_mux_14_11 : IN std_logic ;
         d_arr_mux_14_10 : IN std_logic ;
         d_arr_mux_14_9 : IN std_logic ;
         d_arr_mux_14_8 : IN std_logic ;
         d_arr_mux_14_7 : IN std_logic ;
         d_arr_mux_14_6 : IN std_logic ;
         d_arr_mux_14_5 : IN std_logic ;
         d_arr_mux_14_4 : IN std_logic ;
         d_arr_mux_14_3 : IN std_logic ;
         d_arr_mux_14_2 : IN std_logic ;
         d_arr_mux_14_1 : IN std_logic ;
         d_arr_mux_14_0 : IN std_logic ;
         d_arr_mux_15_31 : IN std_logic ;
         d_arr_mux_15_30 : IN std_logic ;
         d_arr_mux_15_29 : IN std_logic ;
         d_arr_mux_15_28 : IN std_logic ;
         d_arr_mux_15_27 : IN std_logic ;
         d_arr_mux_15_26 : IN std_logic ;
         d_arr_mux_15_25 : IN std_logic ;
         d_arr_mux_15_24 : IN std_logic ;
         d_arr_mux_15_23 : IN std_logic ;
         d_arr_mux_15_22 : IN std_logic ;
         d_arr_mux_15_21 : IN std_logic ;
         d_arr_mux_15_20 : IN std_logic ;
         d_arr_mux_15_19 : IN std_logic ;
         d_arr_mux_15_18 : IN std_logic ;
         d_arr_mux_15_17 : IN std_logic ;
         d_arr_mux_15_16 : IN std_logic ;
         d_arr_mux_15_15 : IN std_logic ;
         d_arr_mux_15_14 : IN std_logic ;
         d_arr_mux_15_13 : IN std_logic ;
         d_arr_mux_15_12 : IN std_logic ;
         d_arr_mux_15_11 : IN std_logic ;
         d_arr_mux_15_10 : IN std_logic ;
         d_arr_mux_15_9 : IN std_logic ;
         d_arr_mux_15_8 : IN std_logic ;
         d_arr_mux_15_7 : IN std_logic ;
         d_arr_mux_15_6 : IN std_logic ;
         d_arr_mux_15_5 : IN std_logic ;
         d_arr_mux_15_4 : IN std_logic ;
         d_arr_mux_15_3 : IN std_logic ;
         d_arr_mux_15_2 : IN std_logic ;
         d_arr_mux_15_1 : IN std_logic ;
         d_arr_mux_15_0 : IN std_logic ;
         d_arr_mux_16_31 : IN std_logic ;
         d_arr_mux_16_30 : IN std_logic ;
         d_arr_mux_16_29 : IN std_logic ;
         d_arr_mux_16_28 : IN std_logic ;
         d_arr_mux_16_27 : IN std_logic ;
         d_arr_mux_16_26 : IN std_logic ;
         d_arr_mux_16_25 : IN std_logic ;
         d_arr_mux_16_24 : IN std_logic ;
         d_arr_mux_16_23 : IN std_logic ;
         d_arr_mux_16_22 : IN std_logic ;
         d_arr_mux_16_21 : IN std_logic ;
         d_arr_mux_16_20 : IN std_logic ;
         d_arr_mux_16_19 : IN std_logic ;
         d_arr_mux_16_18 : IN std_logic ;
         d_arr_mux_16_17 : IN std_logic ;
         d_arr_mux_16_16 : IN std_logic ;
         d_arr_mux_16_15 : IN std_logic ;
         d_arr_mux_16_14 : IN std_logic ;
         d_arr_mux_16_13 : IN std_logic ;
         d_arr_mux_16_12 : IN std_logic ;
         d_arr_mux_16_11 : IN std_logic ;
         d_arr_mux_16_10 : IN std_logic ;
         d_arr_mux_16_9 : IN std_logic ;
         d_arr_mux_16_8 : IN std_logic ;
         d_arr_mux_16_7 : IN std_logic ;
         d_arr_mux_16_6 : IN std_logic ;
         d_arr_mux_16_5 : IN std_logic ;
         d_arr_mux_16_4 : IN std_logic ;
         d_arr_mux_16_3 : IN std_logic ;
         d_arr_mux_16_2 : IN std_logic ;
         d_arr_mux_16_1 : IN std_logic ;
         d_arr_mux_16_0 : IN std_logic ;
         d_arr_mux_17_31 : IN std_logic ;
         d_arr_mux_17_30 : IN std_logic ;
         d_arr_mux_17_29 : IN std_logic ;
         d_arr_mux_17_28 : IN std_logic ;
         d_arr_mux_17_27 : IN std_logic ;
         d_arr_mux_17_26 : IN std_logic ;
         d_arr_mux_17_25 : IN std_logic ;
         d_arr_mux_17_24 : IN std_logic ;
         d_arr_mux_17_23 : IN std_logic ;
         d_arr_mux_17_22 : IN std_logic ;
         d_arr_mux_17_21 : IN std_logic ;
         d_arr_mux_17_20 : IN std_logic ;
         d_arr_mux_17_19 : IN std_logic ;
         d_arr_mux_17_18 : IN std_logic ;
         d_arr_mux_17_17 : IN std_logic ;
         d_arr_mux_17_16 : IN std_logic ;
         d_arr_mux_17_15 : IN std_logic ;
         d_arr_mux_17_14 : IN std_logic ;
         d_arr_mux_17_13 : IN std_logic ;
         d_arr_mux_17_12 : IN std_logic ;
         d_arr_mux_17_11 : IN std_logic ;
         d_arr_mux_17_10 : IN std_logic ;
         d_arr_mux_17_9 : IN std_logic ;
         d_arr_mux_17_8 : IN std_logic ;
         d_arr_mux_17_7 : IN std_logic ;
         d_arr_mux_17_6 : IN std_logic ;
         d_arr_mux_17_5 : IN std_logic ;
         d_arr_mux_17_4 : IN std_logic ;
         d_arr_mux_17_3 : IN std_logic ;
         d_arr_mux_17_2 : IN std_logic ;
         d_arr_mux_17_1 : IN std_logic ;
         d_arr_mux_17_0 : IN std_logic ;
         d_arr_mux_18_31 : IN std_logic ;
         d_arr_mux_18_30 : IN std_logic ;
         d_arr_mux_18_29 : IN std_logic ;
         d_arr_mux_18_28 : IN std_logic ;
         d_arr_mux_18_27 : IN std_logic ;
         d_arr_mux_18_26 : IN std_logic ;
         d_arr_mux_18_25 : IN std_logic ;
         d_arr_mux_18_24 : IN std_logic ;
         d_arr_mux_18_23 : IN std_logic ;
         d_arr_mux_18_22 : IN std_logic ;
         d_arr_mux_18_21 : IN std_logic ;
         d_arr_mux_18_20 : IN std_logic ;
         d_arr_mux_18_19 : IN std_logic ;
         d_arr_mux_18_18 : IN std_logic ;
         d_arr_mux_18_17 : IN std_logic ;
         d_arr_mux_18_16 : IN std_logic ;
         d_arr_mux_18_15 : IN std_logic ;
         d_arr_mux_18_14 : IN std_logic ;
         d_arr_mux_18_13 : IN std_logic ;
         d_arr_mux_18_12 : IN std_logic ;
         d_arr_mux_18_11 : IN std_logic ;
         d_arr_mux_18_10 : IN std_logic ;
         d_arr_mux_18_9 : IN std_logic ;
         d_arr_mux_18_8 : IN std_logic ;
         d_arr_mux_18_7 : IN std_logic ;
         d_arr_mux_18_6 : IN std_logic ;
         d_arr_mux_18_5 : IN std_logic ;
         d_arr_mux_18_4 : IN std_logic ;
         d_arr_mux_18_3 : IN std_logic ;
         d_arr_mux_18_2 : IN std_logic ;
         d_arr_mux_18_1 : IN std_logic ;
         d_arr_mux_18_0 : IN std_logic ;
         d_arr_mux_19_31 : IN std_logic ;
         d_arr_mux_19_30 : IN std_logic ;
         d_arr_mux_19_29 : IN std_logic ;
         d_arr_mux_19_28 : IN std_logic ;
         d_arr_mux_19_27 : IN std_logic ;
         d_arr_mux_19_26 : IN std_logic ;
         d_arr_mux_19_25 : IN std_logic ;
         d_arr_mux_19_24 : IN std_logic ;
         d_arr_mux_19_23 : IN std_logic ;
         d_arr_mux_19_22 : IN std_logic ;
         d_arr_mux_19_21 : IN std_logic ;
         d_arr_mux_19_20 : IN std_logic ;
         d_arr_mux_19_19 : IN std_logic ;
         d_arr_mux_19_18 : IN std_logic ;
         d_arr_mux_19_17 : IN std_logic ;
         d_arr_mux_19_16 : IN std_logic ;
         d_arr_mux_19_15 : IN std_logic ;
         d_arr_mux_19_14 : IN std_logic ;
         d_arr_mux_19_13 : IN std_logic ;
         d_arr_mux_19_12 : IN std_logic ;
         d_arr_mux_19_11 : IN std_logic ;
         d_arr_mux_19_10 : IN std_logic ;
         d_arr_mux_19_9 : IN std_logic ;
         d_arr_mux_19_8 : IN std_logic ;
         d_arr_mux_19_7 : IN std_logic ;
         d_arr_mux_19_6 : IN std_logic ;
         d_arr_mux_19_5 : IN std_logic ;
         d_arr_mux_19_4 : IN std_logic ;
         d_arr_mux_19_3 : IN std_logic ;
         d_arr_mux_19_2 : IN std_logic ;
         d_arr_mux_19_1 : IN std_logic ;
         d_arr_mux_19_0 : IN std_logic ;
         d_arr_mux_20_31 : IN std_logic ;
         d_arr_mux_20_30 : IN std_logic ;
         d_arr_mux_20_29 : IN std_logic ;
         d_arr_mux_20_28 : IN std_logic ;
         d_arr_mux_20_27 : IN std_logic ;
         d_arr_mux_20_26 : IN std_logic ;
         d_arr_mux_20_25 : IN std_logic ;
         d_arr_mux_20_24 : IN std_logic ;
         d_arr_mux_20_23 : IN std_logic ;
         d_arr_mux_20_22 : IN std_logic ;
         d_arr_mux_20_21 : IN std_logic ;
         d_arr_mux_20_20 : IN std_logic ;
         d_arr_mux_20_19 : IN std_logic ;
         d_arr_mux_20_18 : IN std_logic ;
         d_arr_mux_20_17 : IN std_logic ;
         d_arr_mux_20_16 : IN std_logic ;
         d_arr_mux_20_15 : IN std_logic ;
         d_arr_mux_20_14 : IN std_logic ;
         d_arr_mux_20_13 : IN std_logic ;
         d_arr_mux_20_12 : IN std_logic ;
         d_arr_mux_20_11 : IN std_logic ;
         d_arr_mux_20_10 : IN std_logic ;
         d_arr_mux_20_9 : IN std_logic ;
         d_arr_mux_20_8 : IN std_logic ;
         d_arr_mux_20_7 : IN std_logic ;
         d_arr_mux_20_6 : IN std_logic ;
         d_arr_mux_20_5 : IN std_logic ;
         d_arr_mux_20_4 : IN std_logic ;
         d_arr_mux_20_3 : IN std_logic ;
         d_arr_mux_20_2 : IN std_logic ;
         d_arr_mux_20_1 : IN std_logic ;
         d_arr_mux_20_0 : IN std_logic ;
         d_arr_mux_21_31 : IN std_logic ;
         d_arr_mux_21_30 : IN std_logic ;
         d_arr_mux_21_29 : IN std_logic ;
         d_arr_mux_21_28 : IN std_logic ;
         d_arr_mux_21_27 : IN std_logic ;
         d_arr_mux_21_26 : IN std_logic ;
         d_arr_mux_21_25 : IN std_logic ;
         d_arr_mux_21_24 : IN std_logic ;
         d_arr_mux_21_23 : IN std_logic ;
         d_arr_mux_21_22 : IN std_logic ;
         d_arr_mux_21_21 : IN std_logic ;
         d_arr_mux_21_20 : IN std_logic ;
         d_arr_mux_21_19 : IN std_logic ;
         d_arr_mux_21_18 : IN std_logic ;
         d_arr_mux_21_17 : IN std_logic ;
         d_arr_mux_21_16 : IN std_logic ;
         d_arr_mux_21_15 : IN std_logic ;
         d_arr_mux_21_14 : IN std_logic ;
         d_arr_mux_21_13 : IN std_logic ;
         d_arr_mux_21_12 : IN std_logic ;
         d_arr_mux_21_11 : IN std_logic ;
         d_arr_mux_21_10 : IN std_logic ;
         d_arr_mux_21_9 : IN std_logic ;
         d_arr_mux_21_8 : IN std_logic ;
         d_arr_mux_21_7 : IN std_logic ;
         d_arr_mux_21_6 : IN std_logic ;
         d_arr_mux_21_5 : IN std_logic ;
         d_arr_mux_21_4 : IN std_logic ;
         d_arr_mux_21_3 : IN std_logic ;
         d_arr_mux_21_2 : IN std_logic ;
         d_arr_mux_21_1 : IN std_logic ;
         d_arr_mux_21_0 : IN std_logic ;
         d_arr_mux_22_31 : IN std_logic ;
         d_arr_mux_22_30 : IN std_logic ;
         d_arr_mux_22_29 : IN std_logic ;
         d_arr_mux_22_28 : IN std_logic ;
         d_arr_mux_22_27 : IN std_logic ;
         d_arr_mux_22_26 : IN std_logic ;
         d_arr_mux_22_25 : IN std_logic ;
         d_arr_mux_22_24 : IN std_logic ;
         d_arr_mux_22_23 : IN std_logic ;
         d_arr_mux_22_22 : IN std_logic ;
         d_arr_mux_22_21 : IN std_logic ;
         d_arr_mux_22_20 : IN std_logic ;
         d_arr_mux_22_19 : IN std_logic ;
         d_arr_mux_22_18 : IN std_logic ;
         d_arr_mux_22_17 : IN std_logic ;
         d_arr_mux_22_16 : IN std_logic ;
         d_arr_mux_22_15 : IN std_logic ;
         d_arr_mux_22_14 : IN std_logic ;
         d_arr_mux_22_13 : IN std_logic ;
         d_arr_mux_22_12 : IN std_logic ;
         d_arr_mux_22_11 : IN std_logic ;
         d_arr_mux_22_10 : IN std_logic ;
         d_arr_mux_22_9 : IN std_logic ;
         d_arr_mux_22_8 : IN std_logic ;
         d_arr_mux_22_7 : IN std_logic ;
         d_arr_mux_22_6 : IN std_logic ;
         d_arr_mux_22_5 : IN std_logic ;
         d_arr_mux_22_4 : IN std_logic ;
         d_arr_mux_22_3 : IN std_logic ;
         d_arr_mux_22_2 : IN std_logic ;
         d_arr_mux_22_1 : IN std_logic ;
         d_arr_mux_22_0 : IN std_logic ;
         d_arr_mux_23_31 : IN std_logic ;
         d_arr_mux_23_30 : IN std_logic ;
         d_arr_mux_23_29 : IN std_logic ;
         d_arr_mux_23_28 : IN std_logic ;
         d_arr_mux_23_27 : IN std_logic ;
         d_arr_mux_23_26 : IN std_logic ;
         d_arr_mux_23_25 : IN std_logic ;
         d_arr_mux_23_24 : IN std_logic ;
         d_arr_mux_23_23 : IN std_logic ;
         d_arr_mux_23_22 : IN std_logic ;
         d_arr_mux_23_21 : IN std_logic ;
         d_arr_mux_23_20 : IN std_logic ;
         d_arr_mux_23_19 : IN std_logic ;
         d_arr_mux_23_18 : IN std_logic ;
         d_arr_mux_23_17 : IN std_logic ;
         d_arr_mux_23_16 : IN std_logic ;
         d_arr_mux_23_15 : IN std_logic ;
         d_arr_mux_23_14 : IN std_logic ;
         d_arr_mux_23_13 : IN std_logic ;
         d_arr_mux_23_12 : IN std_logic ;
         d_arr_mux_23_11 : IN std_logic ;
         d_arr_mux_23_10 : IN std_logic ;
         d_arr_mux_23_9 : IN std_logic ;
         d_arr_mux_23_8 : IN std_logic ;
         d_arr_mux_23_7 : IN std_logic ;
         d_arr_mux_23_6 : IN std_logic ;
         d_arr_mux_23_5 : IN std_logic ;
         d_arr_mux_23_4 : IN std_logic ;
         d_arr_mux_23_3 : IN std_logic ;
         d_arr_mux_23_2 : IN std_logic ;
         d_arr_mux_23_1 : IN std_logic ;
         d_arr_mux_23_0 : IN std_logic ;
         d_arr_mux_24_31 : IN std_logic ;
         d_arr_mux_24_30 : IN std_logic ;
         d_arr_mux_24_29 : IN std_logic ;
         d_arr_mux_24_28 : IN std_logic ;
         d_arr_mux_24_27 : IN std_logic ;
         d_arr_mux_24_26 : IN std_logic ;
         d_arr_mux_24_25 : IN std_logic ;
         d_arr_mux_24_24 : IN std_logic ;
         d_arr_mux_24_23 : IN std_logic ;
         d_arr_mux_24_22 : IN std_logic ;
         d_arr_mux_24_21 : IN std_logic ;
         d_arr_mux_24_20 : IN std_logic ;
         d_arr_mux_24_19 : IN std_logic ;
         d_arr_mux_24_18 : IN std_logic ;
         d_arr_mux_24_17 : IN std_logic ;
         d_arr_mux_24_16 : IN std_logic ;
         d_arr_mux_24_15 : IN std_logic ;
         d_arr_mux_24_14 : IN std_logic ;
         d_arr_mux_24_13 : IN std_logic ;
         d_arr_mux_24_12 : IN std_logic ;
         d_arr_mux_24_11 : IN std_logic ;
         d_arr_mux_24_10 : IN std_logic ;
         d_arr_mux_24_9 : IN std_logic ;
         d_arr_mux_24_8 : IN std_logic ;
         d_arr_mux_24_7 : IN std_logic ;
         d_arr_mux_24_6 : IN std_logic ;
         d_arr_mux_24_5 : IN std_logic ;
         d_arr_mux_24_4 : IN std_logic ;
         d_arr_mux_24_3 : IN std_logic ;
         d_arr_mux_24_2 : IN std_logic ;
         d_arr_mux_24_1 : IN std_logic ;
         d_arr_mux_24_0 : IN std_logic ;
         d_arr_mul_0_31 : IN std_logic ;
         d_arr_mul_0_30 : IN std_logic ;
         d_arr_mul_0_29 : IN std_logic ;
         d_arr_mul_0_28 : IN std_logic ;
         d_arr_mul_0_27 : IN std_logic ;
         d_arr_mul_0_26 : IN std_logic ;
         d_arr_mul_0_25 : IN std_logic ;
         d_arr_mul_0_24 : IN std_logic ;
         d_arr_mul_0_23 : IN std_logic ;
         d_arr_mul_0_22 : IN std_logic ;
         d_arr_mul_0_21 : IN std_logic ;
         d_arr_mul_0_20 : IN std_logic ;
         d_arr_mul_0_19 : IN std_logic ;
         d_arr_mul_0_18 : IN std_logic ;
         d_arr_mul_0_17 : IN std_logic ;
         d_arr_mul_0_16 : IN std_logic ;
         d_arr_mul_0_15 : IN std_logic ;
         d_arr_mul_0_14 : IN std_logic ;
         d_arr_mul_0_13 : IN std_logic ;
         d_arr_mul_0_12 : IN std_logic ;
         d_arr_mul_0_11 : IN std_logic ;
         d_arr_mul_0_10 : IN std_logic ;
         d_arr_mul_0_9 : IN std_logic ;
         d_arr_mul_0_8 : IN std_logic ;
         d_arr_mul_0_7 : IN std_logic ;
         d_arr_mul_0_6 : IN std_logic ;
         d_arr_mul_0_5 : IN std_logic ;
         d_arr_mul_0_4 : IN std_logic ;
         d_arr_mul_0_3 : IN std_logic ;
         d_arr_mul_0_2 : IN std_logic ;
         d_arr_mul_0_1 : IN std_logic ;
         d_arr_mul_0_0 : IN std_logic ;
         d_arr_mul_1_31 : IN std_logic ;
         d_arr_mul_1_30 : IN std_logic ;
         d_arr_mul_1_29 : IN std_logic ;
         d_arr_mul_1_28 : IN std_logic ;
         d_arr_mul_1_27 : IN std_logic ;
         d_arr_mul_1_26 : IN std_logic ;
         d_arr_mul_1_25 : IN std_logic ;
         d_arr_mul_1_24 : IN std_logic ;
         d_arr_mul_1_23 : IN std_logic ;
         d_arr_mul_1_22 : IN std_logic ;
         d_arr_mul_1_21 : IN std_logic ;
         d_arr_mul_1_20 : IN std_logic ;
         d_arr_mul_1_19 : IN std_logic ;
         d_arr_mul_1_18 : IN std_logic ;
         d_arr_mul_1_17 : IN std_logic ;
         d_arr_mul_1_16 : IN std_logic ;
         d_arr_mul_1_15 : IN std_logic ;
         d_arr_mul_1_14 : IN std_logic ;
         d_arr_mul_1_13 : IN std_logic ;
         d_arr_mul_1_12 : IN std_logic ;
         d_arr_mul_1_11 : IN std_logic ;
         d_arr_mul_1_10 : IN std_logic ;
         d_arr_mul_1_9 : IN std_logic ;
         d_arr_mul_1_8 : IN std_logic ;
         d_arr_mul_1_7 : IN std_logic ;
         d_arr_mul_1_6 : IN std_logic ;
         d_arr_mul_1_5 : IN std_logic ;
         d_arr_mul_1_4 : IN std_logic ;
         d_arr_mul_1_3 : IN std_logic ;
         d_arr_mul_1_2 : IN std_logic ;
         d_arr_mul_1_1 : IN std_logic ;
         d_arr_mul_1_0 : IN std_logic ;
         d_arr_mul_2_31 : IN std_logic ;
         d_arr_mul_2_30 : IN std_logic ;
         d_arr_mul_2_29 : IN std_logic ;
         d_arr_mul_2_28 : IN std_logic ;
         d_arr_mul_2_27 : IN std_logic ;
         d_arr_mul_2_26 : IN std_logic ;
         d_arr_mul_2_25 : IN std_logic ;
         d_arr_mul_2_24 : IN std_logic ;
         d_arr_mul_2_23 : IN std_logic ;
         d_arr_mul_2_22 : IN std_logic ;
         d_arr_mul_2_21 : IN std_logic ;
         d_arr_mul_2_20 : IN std_logic ;
         d_arr_mul_2_19 : IN std_logic ;
         d_arr_mul_2_18 : IN std_logic ;
         d_arr_mul_2_17 : IN std_logic ;
         d_arr_mul_2_16 : IN std_logic ;
         d_arr_mul_2_15 : IN std_logic ;
         d_arr_mul_2_14 : IN std_logic ;
         d_arr_mul_2_13 : IN std_logic ;
         d_arr_mul_2_12 : IN std_logic ;
         d_arr_mul_2_11 : IN std_logic ;
         d_arr_mul_2_10 : IN std_logic ;
         d_arr_mul_2_9 : IN std_logic ;
         d_arr_mul_2_8 : IN std_logic ;
         d_arr_mul_2_7 : IN std_logic ;
         d_arr_mul_2_6 : IN std_logic ;
         d_arr_mul_2_5 : IN std_logic ;
         d_arr_mul_2_4 : IN std_logic ;
         d_arr_mul_2_3 : IN std_logic ;
         d_arr_mul_2_2 : IN std_logic ;
         d_arr_mul_2_1 : IN std_logic ;
         d_arr_mul_2_0 : IN std_logic ;
         d_arr_mul_3_31 : IN std_logic ;
         d_arr_mul_3_30 : IN std_logic ;
         d_arr_mul_3_29 : IN std_logic ;
         d_arr_mul_3_28 : IN std_logic ;
         d_arr_mul_3_27 : IN std_logic ;
         d_arr_mul_3_26 : IN std_logic ;
         d_arr_mul_3_25 : IN std_logic ;
         d_arr_mul_3_24 : IN std_logic ;
         d_arr_mul_3_23 : IN std_logic ;
         d_arr_mul_3_22 : IN std_logic ;
         d_arr_mul_3_21 : IN std_logic ;
         d_arr_mul_3_20 : IN std_logic ;
         d_arr_mul_3_19 : IN std_logic ;
         d_arr_mul_3_18 : IN std_logic ;
         d_arr_mul_3_17 : IN std_logic ;
         d_arr_mul_3_16 : IN std_logic ;
         d_arr_mul_3_15 : IN std_logic ;
         d_arr_mul_3_14 : IN std_logic ;
         d_arr_mul_3_13 : IN std_logic ;
         d_arr_mul_3_12 : IN std_logic ;
         d_arr_mul_3_11 : IN std_logic ;
         d_arr_mul_3_10 : IN std_logic ;
         d_arr_mul_3_9 : IN std_logic ;
         d_arr_mul_3_8 : IN std_logic ;
         d_arr_mul_3_7 : IN std_logic ;
         d_arr_mul_3_6 : IN std_logic ;
         d_arr_mul_3_5 : IN std_logic ;
         d_arr_mul_3_4 : IN std_logic ;
         d_arr_mul_3_3 : IN std_logic ;
         d_arr_mul_3_2 : IN std_logic ;
         d_arr_mul_3_1 : IN std_logic ;
         d_arr_mul_3_0 : IN std_logic ;
         d_arr_mul_4_31 : IN std_logic ;
         d_arr_mul_4_30 : IN std_logic ;
         d_arr_mul_4_29 : IN std_logic ;
         d_arr_mul_4_28 : IN std_logic ;
         d_arr_mul_4_27 : IN std_logic ;
         d_arr_mul_4_26 : IN std_logic ;
         d_arr_mul_4_25 : IN std_logic ;
         d_arr_mul_4_24 : IN std_logic ;
         d_arr_mul_4_23 : IN std_logic ;
         d_arr_mul_4_22 : IN std_logic ;
         d_arr_mul_4_21 : IN std_logic ;
         d_arr_mul_4_20 : IN std_logic ;
         d_arr_mul_4_19 : IN std_logic ;
         d_arr_mul_4_18 : IN std_logic ;
         d_arr_mul_4_17 : IN std_logic ;
         d_arr_mul_4_16 : IN std_logic ;
         d_arr_mul_4_15 : IN std_logic ;
         d_arr_mul_4_14 : IN std_logic ;
         d_arr_mul_4_13 : IN std_logic ;
         d_arr_mul_4_12 : IN std_logic ;
         d_arr_mul_4_11 : IN std_logic ;
         d_arr_mul_4_10 : IN std_logic ;
         d_arr_mul_4_9 : IN std_logic ;
         d_arr_mul_4_8 : IN std_logic ;
         d_arr_mul_4_7 : IN std_logic ;
         d_arr_mul_4_6 : IN std_logic ;
         d_arr_mul_4_5 : IN std_logic ;
         d_arr_mul_4_4 : IN std_logic ;
         d_arr_mul_4_3 : IN std_logic ;
         d_arr_mul_4_2 : IN std_logic ;
         d_arr_mul_4_1 : IN std_logic ;
         d_arr_mul_4_0 : IN std_logic ;
         d_arr_mul_5_31 : IN std_logic ;
         d_arr_mul_5_30 : IN std_logic ;
         d_arr_mul_5_29 : IN std_logic ;
         d_arr_mul_5_28 : IN std_logic ;
         d_arr_mul_5_27 : IN std_logic ;
         d_arr_mul_5_26 : IN std_logic ;
         d_arr_mul_5_25 : IN std_logic ;
         d_arr_mul_5_24 : IN std_logic ;
         d_arr_mul_5_23 : IN std_logic ;
         d_arr_mul_5_22 : IN std_logic ;
         d_arr_mul_5_21 : IN std_logic ;
         d_arr_mul_5_20 : IN std_logic ;
         d_arr_mul_5_19 : IN std_logic ;
         d_arr_mul_5_18 : IN std_logic ;
         d_arr_mul_5_17 : IN std_logic ;
         d_arr_mul_5_16 : IN std_logic ;
         d_arr_mul_5_15 : IN std_logic ;
         d_arr_mul_5_14 : IN std_logic ;
         d_arr_mul_5_13 : IN std_logic ;
         d_arr_mul_5_12 : IN std_logic ;
         d_arr_mul_5_11 : IN std_logic ;
         d_arr_mul_5_10 : IN std_logic ;
         d_arr_mul_5_9 : IN std_logic ;
         d_arr_mul_5_8 : IN std_logic ;
         d_arr_mul_5_7 : IN std_logic ;
         d_arr_mul_5_6 : IN std_logic ;
         d_arr_mul_5_5 : IN std_logic ;
         d_arr_mul_5_4 : IN std_logic ;
         d_arr_mul_5_3 : IN std_logic ;
         d_arr_mul_5_2 : IN std_logic ;
         d_arr_mul_5_1 : IN std_logic ;
         d_arr_mul_5_0 : IN std_logic ;
         d_arr_mul_6_31 : IN std_logic ;
         d_arr_mul_6_30 : IN std_logic ;
         d_arr_mul_6_29 : IN std_logic ;
         d_arr_mul_6_28 : IN std_logic ;
         d_arr_mul_6_27 : IN std_logic ;
         d_arr_mul_6_26 : IN std_logic ;
         d_arr_mul_6_25 : IN std_logic ;
         d_arr_mul_6_24 : IN std_logic ;
         d_arr_mul_6_23 : IN std_logic ;
         d_arr_mul_6_22 : IN std_logic ;
         d_arr_mul_6_21 : IN std_logic ;
         d_arr_mul_6_20 : IN std_logic ;
         d_arr_mul_6_19 : IN std_logic ;
         d_arr_mul_6_18 : IN std_logic ;
         d_arr_mul_6_17 : IN std_logic ;
         d_arr_mul_6_16 : IN std_logic ;
         d_arr_mul_6_15 : IN std_logic ;
         d_arr_mul_6_14 : IN std_logic ;
         d_arr_mul_6_13 : IN std_logic ;
         d_arr_mul_6_12 : IN std_logic ;
         d_arr_mul_6_11 : IN std_logic ;
         d_arr_mul_6_10 : IN std_logic ;
         d_arr_mul_6_9 : IN std_logic ;
         d_arr_mul_6_8 : IN std_logic ;
         d_arr_mul_6_7 : IN std_logic ;
         d_arr_mul_6_6 : IN std_logic ;
         d_arr_mul_6_5 : IN std_logic ;
         d_arr_mul_6_4 : IN std_logic ;
         d_arr_mul_6_3 : IN std_logic ;
         d_arr_mul_6_2 : IN std_logic ;
         d_arr_mul_6_1 : IN std_logic ;
         d_arr_mul_6_0 : IN std_logic ;
         d_arr_mul_7_31 : IN std_logic ;
         d_arr_mul_7_30 : IN std_logic ;
         d_arr_mul_7_29 : IN std_logic ;
         d_arr_mul_7_28 : IN std_logic ;
         d_arr_mul_7_27 : IN std_logic ;
         d_arr_mul_7_26 : IN std_logic ;
         d_arr_mul_7_25 : IN std_logic ;
         d_arr_mul_7_24 : IN std_logic ;
         d_arr_mul_7_23 : IN std_logic ;
         d_arr_mul_7_22 : IN std_logic ;
         d_arr_mul_7_21 : IN std_logic ;
         d_arr_mul_7_20 : IN std_logic ;
         d_arr_mul_7_19 : IN std_logic ;
         d_arr_mul_7_18 : IN std_logic ;
         d_arr_mul_7_17 : IN std_logic ;
         d_arr_mul_7_16 : IN std_logic ;
         d_arr_mul_7_15 : IN std_logic ;
         d_arr_mul_7_14 : IN std_logic ;
         d_arr_mul_7_13 : IN std_logic ;
         d_arr_mul_7_12 : IN std_logic ;
         d_arr_mul_7_11 : IN std_logic ;
         d_arr_mul_7_10 : IN std_logic ;
         d_arr_mul_7_9 : IN std_logic ;
         d_arr_mul_7_8 : IN std_logic ;
         d_arr_mul_7_7 : IN std_logic ;
         d_arr_mul_7_6 : IN std_logic ;
         d_arr_mul_7_5 : IN std_logic ;
         d_arr_mul_7_4 : IN std_logic ;
         d_arr_mul_7_3 : IN std_logic ;
         d_arr_mul_7_2 : IN std_logic ;
         d_arr_mul_7_1 : IN std_logic ;
         d_arr_mul_7_0 : IN std_logic ;
         d_arr_mul_8_31 : IN std_logic ;
         d_arr_mul_8_30 : IN std_logic ;
         d_arr_mul_8_29 : IN std_logic ;
         d_arr_mul_8_28 : IN std_logic ;
         d_arr_mul_8_27 : IN std_logic ;
         d_arr_mul_8_26 : IN std_logic ;
         d_arr_mul_8_25 : IN std_logic ;
         d_arr_mul_8_24 : IN std_logic ;
         d_arr_mul_8_23 : IN std_logic ;
         d_arr_mul_8_22 : IN std_logic ;
         d_arr_mul_8_21 : IN std_logic ;
         d_arr_mul_8_20 : IN std_logic ;
         d_arr_mul_8_19 : IN std_logic ;
         d_arr_mul_8_18 : IN std_logic ;
         d_arr_mul_8_17 : IN std_logic ;
         d_arr_mul_8_16 : IN std_logic ;
         d_arr_mul_8_15 : IN std_logic ;
         d_arr_mul_8_14 : IN std_logic ;
         d_arr_mul_8_13 : IN std_logic ;
         d_arr_mul_8_12 : IN std_logic ;
         d_arr_mul_8_11 : IN std_logic ;
         d_arr_mul_8_10 : IN std_logic ;
         d_arr_mul_8_9 : IN std_logic ;
         d_arr_mul_8_8 : IN std_logic ;
         d_arr_mul_8_7 : IN std_logic ;
         d_arr_mul_8_6 : IN std_logic ;
         d_arr_mul_8_5 : IN std_logic ;
         d_arr_mul_8_4 : IN std_logic ;
         d_arr_mul_8_3 : IN std_logic ;
         d_arr_mul_8_2 : IN std_logic ;
         d_arr_mul_8_1 : IN std_logic ;
         d_arr_mul_8_0 : IN std_logic ;
         d_arr_mul_9_31 : IN std_logic ;
         d_arr_mul_9_30 : IN std_logic ;
         d_arr_mul_9_29 : IN std_logic ;
         d_arr_mul_9_28 : IN std_logic ;
         d_arr_mul_9_27 : IN std_logic ;
         d_arr_mul_9_26 : IN std_logic ;
         d_arr_mul_9_25 : IN std_logic ;
         d_arr_mul_9_24 : IN std_logic ;
         d_arr_mul_9_23 : IN std_logic ;
         d_arr_mul_9_22 : IN std_logic ;
         d_arr_mul_9_21 : IN std_logic ;
         d_arr_mul_9_20 : IN std_logic ;
         d_arr_mul_9_19 : IN std_logic ;
         d_arr_mul_9_18 : IN std_logic ;
         d_arr_mul_9_17 : IN std_logic ;
         d_arr_mul_9_16 : IN std_logic ;
         d_arr_mul_9_15 : IN std_logic ;
         d_arr_mul_9_14 : IN std_logic ;
         d_arr_mul_9_13 : IN std_logic ;
         d_arr_mul_9_12 : IN std_logic ;
         d_arr_mul_9_11 : IN std_logic ;
         d_arr_mul_9_10 : IN std_logic ;
         d_arr_mul_9_9 : IN std_logic ;
         d_arr_mul_9_8 : IN std_logic ;
         d_arr_mul_9_7 : IN std_logic ;
         d_arr_mul_9_6 : IN std_logic ;
         d_arr_mul_9_5 : IN std_logic ;
         d_arr_mul_9_4 : IN std_logic ;
         d_arr_mul_9_3 : IN std_logic ;
         d_arr_mul_9_2 : IN std_logic ;
         d_arr_mul_9_1 : IN std_logic ;
         d_arr_mul_9_0 : IN std_logic ;
         d_arr_mul_10_31 : IN std_logic ;
         d_arr_mul_10_30 : IN std_logic ;
         d_arr_mul_10_29 : IN std_logic ;
         d_arr_mul_10_28 : IN std_logic ;
         d_arr_mul_10_27 : IN std_logic ;
         d_arr_mul_10_26 : IN std_logic ;
         d_arr_mul_10_25 : IN std_logic ;
         d_arr_mul_10_24 : IN std_logic ;
         d_arr_mul_10_23 : IN std_logic ;
         d_arr_mul_10_22 : IN std_logic ;
         d_arr_mul_10_21 : IN std_logic ;
         d_arr_mul_10_20 : IN std_logic ;
         d_arr_mul_10_19 : IN std_logic ;
         d_arr_mul_10_18 : IN std_logic ;
         d_arr_mul_10_17 : IN std_logic ;
         d_arr_mul_10_16 : IN std_logic ;
         d_arr_mul_10_15 : IN std_logic ;
         d_arr_mul_10_14 : IN std_logic ;
         d_arr_mul_10_13 : IN std_logic ;
         d_arr_mul_10_12 : IN std_logic ;
         d_arr_mul_10_11 : IN std_logic ;
         d_arr_mul_10_10 : IN std_logic ;
         d_arr_mul_10_9 : IN std_logic ;
         d_arr_mul_10_8 : IN std_logic ;
         d_arr_mul_10_7 : IN std_logic ;
         d_arr_mul_10_6 : IN std_logic ;
         d_arr_mul_10_5 : IN std_logic ;
         d_arr_mul_10_4 : IN std_logic ;
         d_arr_mul_10_3 : IN std_logic ;
         d_arr_mul_10_2 : IN std_logic ;
         d_arr_mul_10_1 : IN std_logic ;
         d_arr_mul_10_0 : IN std_logic ;
         d_arr_mul_11_31 : IN std_logic ;
         d_arr_mul_11_30 : IN std_logic ;
         d_arr_mul_11_29 : IN std_logic ;
         d_arr_mul_11_28 : IN std_logic ;
         d_arr_mul_11_27 : IN std_logic ;
         d_arr_mul_11_26 : IN std_logic ;
         d_arr_mul_11_25 : IN std_logic ;
         d_arr_mul_11_24 : IN std_logic ;
         d_arr_mul_11_23 : IN std_logic ;
         d_arr_mul_11_22 : IN std_logic ;
         d_arr_mul_11_21 : IN std_logic ;
         d_arr_mul_11_20 : IN std_logic ;
         d_arr_mul_11_19 : IN std_logic ;
         d_arr_mul_11_18 : IN std_logic ;
         d_arr_mul_11_17 : IN std_logic ;
         d_arr_mul_11_16 : IN std_logic ;
         d_arr_mul_11_15 : IN std_logic ;
         d_arr_mul_11_14 : IN std_logic ;
         d_arr_mul_11_13 : IN std_logic ;
         d_arr_mul_11_12 : IN std_logic ;
         d_arr_mul_11_11 : IN std_logic ;
         d_arr_mul_11_10 : IN std_logic ;
         d_arr_mul_11_9 : IN std_logic ;
         d_arr_mul_11_8 : IN std_logic ;
         d_arr_mul_11_7 : IN std_logic ;
         d_arr_mul_11_6 : IN std_logic ;
         d_arr_mul_11_5 : IN std_logic ;
         d_arr_mul_11_4 : IN std_logic ;
         d_arr_mul_11_3 : IN std_logic ;
         d_arr_mul_11_2 : IN std_logic ;
         d_arr_mul_11_1 : IN std_logic ;
         d_arr_mul_11_0 : IN std_logic ;
         d_arr_mul_12_31 : IN std_logic ;
         d_arr_mul_12_30 : IN std_logic ;
         d_arr_mul_12_29 : IN std_logic ;
         d_arr_mul_12_28 : IN std_logic ;
         d_arr_mul_12_27 : IN std_logic ;
         d_arr_mul_12_26 : IN std_logic ;
         d_arr_mul_12_25 : IN std_logic ;
         d_arr_mul_12_24 : IN std_logic ;
         d_arr_mul_12_23 : IN std_logic ;
         d_arr_mul_12_22 : IN std_logic ;
         d_arr_mul_12_21 : IN std_logic ;
         d_arr_mul_12_20 : IN std_logic ;
         d_arr_mul_12_19 : IN std_logic ;
         d_arr_mul_12_18 : IN std_logic ;
         d_arr_mul_12_17 : IN std_logic ;
         d_arr_mul_12_16 : IN std_logic ;
         d_arr_mul_12_15 : IN std_logic ;
         d_arr_mul_12_14 : IN std_logic ;
         d_arr_mul_12_13 : IN std_logic ;
         d_arr_mul_12_12 : IN std_logic ;
         d_arr_mul_12_11 : IN std_logic ;
         d_arr_mul_12_10 : IN std_logic ;
         d_arr_mul_12_9 : IN std_logic ;
         d_arr_mul_12_8 : IN std_logic ;
         d_arr_mul_12_7 : IN std_logic ;
         d_arr_mul_12_6 : IN std_logic ;
         d_arr_mul_12_5 : IN std_logic ;
         d_arr_mul_12_4 : IN std_logic ;
         d_arr_mul_12_3 : IN std_logic ;
         d_arr_mul_12_2 : IN std_logic ;
         d_arr_mul_12_1 : IN std_logic ;
         d_arr_mul_12_0 : IN std_logic ;
         d_arr_mul_13_31 : IN std_logic ;
         d_arr_mul_13_30 : IN std_logic ;
         d_arr_mul_13_29 : IN std_logic ;
         d_arr_mul_13_28 : IN std_logic ;
         d_arr_mul_13_27 : IN std_logic ;
         d_arr_mul_13_26 : IN std_logic ;
         d_arr_mul_13_25 : IN std_logic ;
         d_arr_mul_13_24 : IN std_logic ;
         d_arr_mul_13_23 : IN std_logic ;
         d_arr_mul_13_22 : IN std_logic ;
         d_arr_mul_13_21 : IN std_logic ;
         d_arr_mul_13_20 : IN std_logic ;
         d_arr_mul_13_19 : IN std_logic ;
         d_arr_mul_13_18 : IN std_logic ;
         d_arr_mul_13_17 : IN std_logic ;
         d_arr_mul_13_16 : IN std_logic ;
         d_arr_mul_13_15 : IN std_logic ;
         d_arr_mul_13_14 : IN std_logic ;
         d_arr_mul_13_13 : IN std_logic ;
         d_arr_mul_13_12 : IN std_logic ;
         d_arr_mul_13_11 : IN std_logic ;
         d_arr_mul_13_10 : IN std_logic ;
         d_arr_mul_13_9 : IN std_logic ;
         d_arr_mul_13_8 : IN std_logic ;
         d_arr_mul_13_7 : IN std_logic ;
         d_arr_mul_13_6 : IN std_logic ;
         d_arr_mul_13_5 : IN std_logic ;
         d_arr_mul_13_4 : IN std_logic ;
         d_arr_mul_13_3 : IN std_logic ;
         d_arr_mul_13_2 : IN std_logic ;
         d_arr_mul_13_1 : IN std_logic ;
         d_arr_mul_13_0 : IN std_logic ;
         d_arr_mul_14_31 : IN std_logic ;
         d_arr_mul_14_30 : IN std_logic ;
         d_arr_mul_14_29 : IN std_logic ;
         d_arr_mul_14_28 : IN std_logic ;
         d_arr_mul_14_27 : IN std_logic ;
         d_arr_mul_14_26 : IN std_logic ;
         d_arr_mul_14_25 : IN std_logic ;
         d_arr_mul_14_24 : IN std_logic ;
         d_arr_mul_14_23 : IN std_logic ;
         d_arr_mul_14_22 : IN std_logic ;
         d_arr_mul_14_21 : IN std_logic ;
         d_arr_mul_14_20 : IN std_logic ;
         d_arr_mul_14_19 : IN std_logic ;
         d_arr_mul_14_18 : IN std_logic ;
         d_arr_mul_14_17 : IN std_logic ;
         d_arr_mul_14_16 : IN std_logic ;
         d_arr_mul_14_15 : IN std_logic ;
         d_arr_mul_14_14 : IN std_logic ;
         d_arr_mul_14_13 : IN std_logic ;
         d_arr_mul_14_12 : IN std_logic ;
         d_arr_mul_14_11 : IN std_logic ;
         d_arr_mul_14_10 : IN std_logic ;
         d_arr_mul_14_9 : IN std_logic ;
         d_arr_mul_14_8 : IN std_logic ;
         d_arr_mul_14_7 : IN std_logic ;
         d_arr_mul_14_6 : IN std_logic ;
         d_arr_mul_14_5 : IN std_logic ;
         d_arr_mul_14_4 : IN std_logic ;
         d_arr_mul_14_3 : IN std_logic ;
         d_arr_mul_14_2 : IN std_logic ;
         d_arr_mul_14_1 : IN std_logic ;
         d_arr_mul_14_0 : IN std_logic ;
         d_arr_mul_15_31 : IN std_logic ;
         d_arr_mul_15_30 : IN std_logic ;
         d_arr_mul_15_29 : IN std_logic ;
         d_arr_mul_15_28 : IN std_logic ;
         d_arr_mul_15_27 : IN std_logic ;
         d_arr_mul_15_26 : IN std_logic ;
         d_arr_mul_15_25 : IN std_logic ;
         d_arr_mul_15_24 : IN std_logic ;
         d_arr_mul_15_23 : IN std_logic ;
         d_arr_mul_15_22 : IN std_logic ;
         d_arr_mul_15_21 : IN std_logic ;
         d_arr_mul_15_20 : IN std_logic ;
         d_arr_mul_15_19 : IN std_logic ;
         d_arr_mul_15_18 : IN std_logic ;
         d_arr_mul_15_17 : IN std_logic ;
         d_arr_mul_15_16 : IN std_logic ;
         d_arr_mul_15_15 : IN std_logic ;
         d_arr_mul_15_14 : IN std_logic ;
         d_arr_mul_15_13 : IN std_logic ;
         d_arr_mul_15_12 : IN std_logic ;
         d_arr_mul_15_11 : IN std_logic ;
         d_arr_mul_15_10 : IN std_logic ;
         d_arr_mul_15_9 : IN std_logic ;
         d_arr_mul_15_8 : IN std_logic ;
         d_arr_mul_15_7 : IN std_logic ;
         d_arr_mul_15_6 : IN std_logic ;
         d_arr_mul_15_5 : IN std_logic ;
         d_arr_mul_15_4 : IN std_logic ;
         d_arr_mul_15_3 : IN std_logic ;
         d_arr_mul_15_2 : IN std_logic ;
         d_arr_mul_15_1 : IN std_logic ;
         d_arr_mul_15_0 : IN std_logic ;
         d_arr_mul_16_31 : IN std_logic ;
         d_arr_mul_16_30 : IN std_logic ;
         d_arr_mul_16_29 : IN std_logic ;
         d_arr_mul_16_28 : IN std_logic ;
         d_arr_mul_16_27 : IN std_logic ;
         d_arr_mul_16_26 : IN std_logic ;
         d_arr_mul_16_25 : IN std_logic ;
         d_arr_mul_16_24 : IN std_logic ;
         d_arr_mul_16_23 : IN std_logic ;
         d_arr_mul_16_22 : IN std_logic ;
         d_arr_mul_16_21 : IN std_logic ;
         d_arr_mul_16_20 : IN std_logic ;
         d_arr_mul_16_19 : IN std_logic ;
         d_arr_mul_16_18 : IN std_logic ;
         d_arr_mul_16_17 : IN std_logic ;
         d_arr_mul_16_16 : IN std_logic ;
         d_arr_mul_16_15 : IN std_logic ;
         d_arr_mul_16_14 : IN std_logic ;
         d_arr_mul_16_13 : IN std_logic ;
         d_arr_mul_16_12 : IN std_logic ;
         d_arr_mul_16_11 : IN std_logic ;
         d_arr_mul_16_10 : IN std_logic ;
         d_arr_mul_16_9 : IN std_logic ;
         d_arr_mul_16_8 : IN std_logic ;
         d_arr_mul_16_7 : IN std_logic ;
         d_arr_mul_16_6 : IN std_logic ;
         d_arr_mul_16_5 : IN std_logic ;
         d_arr_mul_16_4 : IN std_logic ;
         d_arr_mul_16_3 : IN std_logic ;
         d_arr_mul_16_2 : IN std_logic ;
         d_arr_mul_16_1 : IN std_logic ;
         d_arr_mul_16_0 : IN std_logic ;
         d_arr_mul_17_31 : IN std_logic ;
         d_arr_mul_17_30 : IN std_logic ;
         d_arr_mul_17_29 : IN std_logic ;
         d_arr_mul_17_28 : IN std_logic ;
         d_arr_mul_17_27 : IN std_logic ;
         d_arr_mul_17_26 : IN std_logic ;
         d_arr_mul_17_25 : IN std_logic ;
         d_arr_mul_17_24 : IN std_logic ;
         d_arr_mul_17_23 : IN std_logic ;
         d_arr_mul_17_22 : IN std_logic ;
         d_arr_mul_17_21 : IN std_logic ;
         d_arr_mul_17_20 : IN std_logic ;
         d_arr_mul_17_19 : IN std_logic ;
         d_arr_mul_17_18 : IN std_logic ;
         d_arr_mul_17_17 : IN std_logic ;
         d_arr_mul_17_16 : IN std_logic ;
         d_arr_mul_17_15 : IN std_logic ;
         d_arr_mul_17_14 : IN std_logic ;
         d_arr_mul_17_13 : IN std_logic ;
         d_arr_mul_17_12 : IN std_logic ;
         d_arr_mul_17_11 : IN std_logic ;
         d_arr_mul_17_10 : IN std_logic ;
         d_arr_mul_17_9 : IN std_logic ;
         d_arr_mul_17_8 : IN std_logic ;
         d_arr_mul_17_7 : IN std_logic ;
         d_arr_mul_17_6 : IN std_logic ;
         d_arr_mul_17_5 : IN std_logic ;
         d_arr_mul_17_4 : IN std_logic ;
         d_arr_mul_17_3 : IN std_logic ;
         d_arr_mul_17_2 : IN std_logic ;
         d_arr_mul_17_1 : IN std_logic ;
         d_arr_mul_17_0 : IN std_logic ;
         d_arr_mul_18_31 : IN std_logic ;
         d_arr_mul_18_30 : IN std_logic ;
         d_arr_mul_18_29 : IN std_logic ;
         d_arr_mul_18_28 : IN std_logic ;
         d_arr_mul_18_27 : IN std_logic ;
         d_arr_mul_18_26 : IN std_logic ;
         d_arr_mul_18_25 : IN std_logic ;
         d_arr_mul_18_24 : IN std_logic ;
         d_arr_mul_18_23 : IN std_logic ;
         d_arr_mul_18_22 : IN std_logic ;
         d_arr_mul_18_21 : IN std_logic ;
         d_arr_mul_18_20 : IN std_logic ;
         d_arr_mul_18_19 : IN std_logic ;
         d_arr_mul_18_18 : IN std_logic ;
         d_arr_mul_18_17 : IN std_logic ;
         d_arr_mul_18_16 : IN std_logic ;
         d_arr_mul_18_15 : IN std_logic ;
         d_arr_mul_18_14 : IN std_logic ;
         d_arr_mul_18_13 : IN std_logic ;
         d_arr_mul_18_12 : IN std_logic ;
         d_arr_mul_18_11 : IN std_logic ;
         d_arr_mul_18_10 : IN std_logic ;
         d_arr_mul_18_9 : IN std_logic ;
         d_arr_mul_18_8 : IN std_logic ;
         d_arr_mul_18_7 : IN std_logic ;
         d_arr_mul_18_6 : IN std_logic ;
         d_arr_mul_18_5 : IN std_logic ;
         d_arr_mul_18_4 : IN std_logic ;
         d_arr_mul_18_3 : IN std_logic ;
         d_arr_mul_18_2 : IN std_logic ;
         d_arr_mul_18_1 : IN std_logic ;
         d_arr_mul_18_0 : IN std_logic ;
         d_arr_mul_19_31 : IN std_logic ;
         d_arr_mul_19_30 : IN std_logic ;
         d_arr_mul_19_29 : IN std_logic ;
         d_arr_mul_19_28 : IN std_logic ;
         d_arr_mul_19_27 : IN std_logic ;
         d_arr_mul_19_26 : IN std_logic ;
         d_arr_mul_19_25 : IN std_logic ;
         d_arr_mul_19_24 : IN std_logic ;
         d_arr_mul_19_23 : IN std_logic ;
         d_arr_mul_19_22 : IN std_logic ;
         d_arr_mul_19_21 : IN std_logic ;
         d_arr_mul_19_20 : IN std_logic ;
         d_arr_mul_19_19 : IN std_logic ;
         d_arr_mul_19_18 : IN std_logic ;
         d_arr_mul_19_17 : IN std_logic ;
         d_arr_mul_19_16 : IN std_logic ;
         d_arr_mul_19_15 : IN std_logic ;
         d_arr_mul_19_14 : IN std_logic ;
         d_arr_mul_19_13 : IN std_logic ;
         d_arr_mul_19_12 : IN std_logic ;
         d_arr_mul_19_11 : IN std_logic ;
         d_arr_mul_19_10 : IN std_logic ;
         d_arr_mul_19_9 : IN std_logic ;
         d_arr_mul_19_8 : IN std_logic ;
         d_arr_mul_19_7 : IN std_logic ;
         d_arr_mul_19_6 : IN std_logic ;
         d_arr_mul_19_5 : IN std_logic ;
         d_arr_mul_19_4 : IN std_logic ;
         d_arr_mul_19_3 : IN std_logic ;
         d_arr_mul_19_2 : IN std_logic ;
         d_arr_mul_19_1 : IN std_logic ;
         d_arr_mul_19_0 : IN std_logic ;
         d_arr_mul_20_31 : IN std_logic ;
         d_arr_mul_20_30 : IN std_logic ;
         d_arr_mul_20_29 : IN std_logic ;
         d_arr_mul_20_28 : IN std_logic ;
         d_arr_mul_20_27 : IN std_logic ;
         d_arr_mul_20_26 : IN std_logic ;
         d_arr_mul_20_25 : IN std_logic ;
         d_arr_mul_20_24 : IN std_logic ;
         d_arr_mul_20_23 : IN std_logic ;
         d_arr_mul_20_22 : IN std_logic ;
         d_arr_mul_20_21 : IN std_logic ;
         d_arr_mul_20_20 : IN std_logic ;
         d_arr_mul_20_19 : IN std_logic ;
         d_arr_mul_20_18 : IN std_logic ;
         d_arr_mul_20_17 : IN std_logic ;
         d_arr_mul_20_16 : IN std_logic ;
         d_arr_mul_20_15 : IN std_logic ;
         d_arr_mul_20_14 : IN std_logic ;
         d_arr_mul_20_13 : IN std_logic ;
         d_arr_mul_20_12 : IN std_logic ;
         d_arr_mul_20_11 : IN std_logic ;
         d_arr_mul_20_10 : IN std_logic ;
         d_arr_mul_20_9 : IN std_logic ;
         d_arr_mul_20_8 : IN std_logic ;
         d_arr_mul_20_7 : IN std_logic ;
         d_arr_mul_20_6 : IN std_logic ;
         d_arr_mul_20_5 : IN std_logic ;
         d_arr_mul_20_4 : IN std_logic ;
         d_arr_mul_20_3 : IN std_logic ;
         d_arr_mul_20_2 : IN std_logic ;
         d_arr_mul_20_1 : IN std_logic ;
         d_arr_mul_20_0 : IN std_logic ;
         d_arr_mul_21_31 : IN std_logic ;
         d_arr_mul_21_30 : IN std_logic ;
         d_arr_mul_21_29 : IN std_logic ;
         d_arr_mul_21_28 : IN std_logic ;
         d_arr_mul_21_27 : IN std_logic ;
         d_arr_mul_21_26 : IN std_logic ;
         d_arr_mul_21_25 : IN std_logic ;
         d_arr_mul_21_24 : IN std_logic ;
         d_arr_mul_21_23 : IN std_logic ;
         d_arr_mul_21_22 : IN std_logic ;
         d_arr_mul_21_21 : IN std_logic ;
         d_arr_mul_21_20 : IN std_logic ;
         d_arr_mul_21_19 : IN std_logic ;
         d_arr_mul_21_18 : IN std_logic ;
         d_arr_mul_21_17 : IN std_logic ;
         d_arr_mul_21_16 : IN std_logic ;
         d_arr_mul_21_15 : IN std_logic ;
         d_arr_mul_21_14 : IN std_logic ;
         d_arr_mul_21_13 : IN std_logic ;
         d_arr_mul_21_12 : IN std_logic ;
         d_arr_mul_21_11 : IN std_logic ;
         d_arr_mul_21_10 : IN std_logic ;
         d_arr_mul_21_9 : IN std_logic ;
         d_arr_mul_21_8 : IN std_logic ;
         d_arr_mul_21_7 : IN std_logic ;
         d_arr_mul_21_6 : IN std_logic ;
         d_arr_mul_21_5 : IN std_logic ;
         d_arr_mul_21_4 : IN std_logic ;
         d_arr_mul_21_3 : IN std_logic ;
         d_arr_mul_21_2 : IN std_logic ;
         d_arr_mul_21_1 : IN std_logic ;
         d_arr_mul_21_0 : IN std_logic ;
         d_arr_mul_22_31 : IN std_logic ;
         d_arr_mul_22_30 : IN std_logic ;
         d_arr_mul_22_29 : IN std_logic ;
         d_arr_mul_22_28 : IN std_logic ;
         d_arr_mul_22_27 : IN std_logic ;
         d_arr_mul_22_26 : IN std_logic ;
         d_arr_mul_22_25 : IN std_logic ;
         d_arr_mul_22_24 : IN std_logic ;
         d_arr_mul_22_23 : IN std_logic ;
         d_arr_mul_22_22 : IN std_logic ;
         d_arr_mul_22_21 : IN std_logic ;
         d_arr_mul_22_20 : IN std_logic ;
         d_arr_mul_22_19 : IN std_logic ;
         d_arr_mul_22_18 : IN std_logic ;
         d_arr_mul_22_17 : IN std_logic ;
         d_arr_mul_22_16 : IN std_logic ;
         d_arr_mul_22_15 : IN std_logic ;
         d_arr_mul_22_14 : IN std_logic ;
         d_arr_mul_22_13 : IN std_logic ;
         d_arr_mul_22_12 : IN std_logic ;
         d_arr_mul_22_11 : IN std_logic ;
         d_arr_mul_22_10 : IN std_logic ;
         d_arr_mul_22_9 : IN std_logic ;
         d_arr_mul_22_8 : IN std_logic ;
         d_arr_mul_22_7 : IN std_logic ;
         d_arr_mul_22_6 : IN std_logic ;
         d_arr_mul_22_5 : IN std_logic ;
         d_arr_mul_22_4 : IN std_logic ;
         d_arr_mul_22_3 : IN std_logic ;
         d_arr_mul_22_2 : IN std_logic ;
         d_arr_mul_22_1 : IN std_logic ;
         d_arr_mul_22_0 : IN std_logic ;
         d_arr_mul_23_31 : IN std_logic ;
         d_arr_mul_23_30 : IN std_logic ;
         d_arr_mul_23_29 : IN std_logic ;
         d_arr_mul_23_28 : IN std_logic ;
         d_arr_mul_23_27 : IN std_logic ;
         d_arr_mul_23_26 : IN std_logic ;
         d_arr_mul_23_25 : IN std_logic ;
         d_arr_mul_23_24 : IN std_logic ;
         d_arr_mul_23_23 : IN std_logic ;
         d_arr_mul_23_22 : IN std_logic ;
         d_arr_mul_23_21 : IN std_logic ;
         d_arr_mul_23_20 : IN std_logic ;
         d_arr_mul_23_19 : IN std_logic ;
         d_arr_mul_23_18 : IN std_logic ;
         d_arr_mul_23_17 : IN std_logic ;
         d_arr_mul_23_16 : IN std_logic ;
         d_arr_mul_23_15 : IN std_logic ;
         d_arr_mul_23_14 : IN std_logic ;
         d_arr_mul_23_13 : IN std_logic ;
         d_arr_mul_23_12 : IN std_logic ;
         d_arr_mul_23_11 : IN std_logic ;
         d_arr_mul_23_10 : IN std_logic ;
         d_arr_mul_23_9 : IN std_logic ;
         d_arr_mul_23_8 : IN std_logic ;
         d_arr_mul_23_7 : IN std_logic ;
         d_arr_mul_23_6 : IN std_logic ;
         d_arr_mul_23_5 : IN std_logic ;
         d_arr_mul_23_4 : IN std_logic ;
         d_arr_mul_23_3 : IN std_logic ;
         d_arr_mul_23_2 : IN std_logic ;
         d_arr_mul_23_1 : IN std_logic ;
         d_arr_mul_23_0 : IN std_logic ;
         d_arr_mul_24_31 : IN std_logic ;
         d_arr_mul_24_30 : IN std_logic ;
         d_arr_mul_24_29 : IN std_logic ;
         d_arr_mul_24_28 : IN std_logic ;
         d_arr_mul_24_27 : IN std_logic ;
         d_arr_mul_24_26 : IN std_logic ;
         d_arr_mul_24_25 : IN std_logic ;
         d_arr_mul_24_24 : IN std_logic ;
         d_arr_mul_24_23 : IN std_logic ;
         d_arr_mul_24_22 : IN std_logic ;
         d_arr_mul_24_21 : IN std_logic ;
         d_arr_mul_24_20 : IN std_logic ;
         d_arr_mul_24_19 : IN std_logic ;
         d_arr_mul_24_18 : IN std_logic ;
         d_arr_mul_24_17 : IN std_logic ;
         d_arr_mul_24_16 : IN std_logic ;
         d_arr_mul_24_15 : IN std_logic ;
         d_arr_mul_24_14 : IN std_logic ;
         d_arr_mul_24_13 : IN std_logic ;
         d_arr_mul_24_12 : IN std_logic ;
         d_arr_mul_24_11 : IN std_logic ;
         d_arr_mul_24_10 : IN std_logic ;
         d_arr_mul_24_9 : IN std_logic ;
         d_arr_mul_24_8 : IN std_logic ;
         d_arr_mul_24_7 : IN std_logic ;
         d_arr_mul_24_6 : IN std_logic ;
         d_arr_mul_24_5 : IN std_logic ;
         d_arr_mul_24_4 : IN std_logic ;
         d_arr_mul_24_3 : IN std_logic ;
         d_arr_mul_24_2 : IN std_logic ;
         d_arr_mul_24_1 : IN std_logic ;
         d_arr_mul_24_0 : IN std_logic ;
         d_arr_add_0_31 : IN std_logic ;
         d_arr_add_0_30 : IN std_logic ;
         d_arr_add_0_29 : IN std_logic ;
         d_arr_add_0_28 : IN std_logic ;
         d_arr_add_0_27 : IN std_logic ;
         d_arr_add_0_26 : IN std_logic ;
         d_arr_add_0_25 : IN std_logic ;
         d_arr_add_0_24 : IN std_logic ;
         d_arr_add_0_23 : IN std_logic ;
         d_arr_add_0_22 : IN std_logic ;
         d_arr_add_0_21 : IN std_logic ;
         d_arr_add_0_20 : IN std_logic ;
         d_arr_add_0_19 : IN std_logic ;
         d_arr_add_0_18 : IN std_logic ;
         d_arr_add_0_17 : IN std_logic ;
         d_arr_add_0_16 : IN std_logic ;
         d_arr_add_0_15 : IN std_logic ;
         d_arr_add_0_14 : IN std_logic ;
         d_arr_add_0_13 : IN std_logic ;
         d_arr_add_0_12 : IN std_logic ;
         d_arr_add_0_11 : IN std_logic ;
         d_arr_add_0_10 : IN std_logic ;
         d_arr_add_0_9 : IN std_logic ;
         d_arr_add_0_8 : IN std_logic ;
         d_arr_add_0_7 : IN std_logic ;
         d_arr_add_0_6 : IN std_logic ;
         d_arr_add_0_5 : IN std_logic ;
         d_arr_add_0_4 : IN std_logic ;
         d_arr_add_0_3 : IN std_logic ;
         d_arr_add_0_2 : IN std_logic ;
         d_arr_add_0_1 : IN std_logic ;
         d_arr_add_0_0 : IN std_logic ;
         d_arr_add_1_31 : IN std_logic ;
         d_arr_add_1_30 : IN std_logic ;
         d_arr_add_1_29 : IN std_logic ;
         d_arr_add_1_28 : IN std_logic ;
         d_arr_add_1_27 : IN std_logic ;
         d_arr_add_1_26 : IN std_logic ;
         d_arr_add_1_25 : IN std_logic ;
         d_arr_add_1_24 : IN std_logic ;
         d_arr_add_1_23 : IN std_logic ;
         d_arr_add_1_22 : IN std_logic ;
         d_arr_add_1_21 : IN std_logic ;
         d_arr_add_1_20 : IN std_logic ;
         d_arr_add_1_19 : IN std_logic ;
         d_arr_add_1_18 : IN std_logic ;
         d_arr_add_1_17 : IN std_logic ;
         d_arr_add_1_16 : IN std_logic ;
         d_arr_add_1_15 : IN std_logic ;
         d_arr_add_1_14 : IN std_logic ;
         d_arr_add_1_13 : IN std_logic ;
         d_arr_add_1_12 : IN std_logic ;
         d_arr_add_1_11 : IN std_logic ;
         d_arr_add_1_10 : IN std_logic ;
         d_arr_add_1_9 : IN std_logic ;
         d_arr_add_1_8 : IN std_logic ;
         d_arr_add_1_7 : IN std_logic ;
         d_arr_add_1_6 : IN std_logic ;
         d_arr_add_1_5 : IN std_logic ;
         d_arr_add_1_4 : IN std_logic ;
         d_arr_add_1_3 : IN std_logic ;
         d_arr_add_1_2 : IN std_logic ;
         d_arr_add_1_1 : IN std_logic ;
         d_arr_add_1_0 : IN std_logic ;
         d_arr_add_2_31 : IN std_logic ;
         d_arr_add_2_30 : IN std_logic ;
         d_arr_add_2_29 : IN std_logic ;
         d_arr_add_2_28 : IN std_logic ;
         d_arr_add_2_27 : IN std_logic ;
         d_arr_add_2_26 : IN std_logic ;
         d_arr_add_2_25 : IN std_logic ;
         d_arr_add_2_24 : IN std_logic ;
         d_arr_add_2_23 : IN std_logic ;
         d_arr_add_2_22 : IN std_logic ;
         d_arr_add_2_21 : IN std_logic ;
         d_arr_add_2_20 : IN std_logic ;
         d_arr_add_2_19 : IN std_logic ;
         d_arr_add_2_18 : IN std_logic ;
         d_arr_add_2_17 : IN std_logic ;
         d_arr_add_2_16 : IN std_logic ;
         d_arr_add_2_15 : IN std_logic ;
         d_arr_add_2_14 : IN std_logic ;
         d_arr_add_2_13 : IN std_logic ;
         d_arr_add_2_12 : IN std_logic ;
         d_arr_add_2_11 : IN std_logic ;
         d_arr_add_2_10 : IN std_logic ;
         d_arr_add_2_9 : IN std_logic ;
         d_arr_add_2_8 : IN std_logic ;
         d_arr_add_2_7 : IN std_logic ;
         d_arr_add_2_6 : IN std_logic ;
         d_arr_add_2_5 : IN std_logic ;
         d_arr_add_2_4 : IN std_logic ;
         d_arr_add_2_3 : IN std_logic ;
         d_arr_add_2_2 : IN std_logic ;
         d_arr_add_2_1 : IN std_logic ;
         d_arr_add_2_0 : IN std_logic ;
         d_arr_add_3_31 : IN std_logic ;
         d_arr_add_3_30 : IN std_logic ;
         d_arr_add_3_29 : IN std_logic ;
         d_arr_add_3_28 : IN std_logic ;
         d_arr_add_3_27 : IN std_logic ;
         d_arr_add_3_26 : IN std_logic ;
         d_arr_add_3_25 : IN std_logic ;
         d_arr_add_3_24 : IN std_logic ;
         d_arr_add_3_23 : IN std_logic ;
         d_arr_add_3_22 : IN std_logic ;
         d_arr_add_3_21 : IN std_logic ;
         d_arr_add_3_20 : IN std_logic ;
         d_arr_add_3_19 : IN std_logic ;
         d_arr_add_3_18 : IN std_logic ;
         d_arr_add_3_17 : IN std_logic ;
         d_arr_add_3_16 : IN std_logic ;
         d_arr_add_3_15 : IN std_logic ;
         d_arr_add_3_14 : IN std_logic ;
         d_arr_add_3_13 : IN std_logic ;
         d_arr_add_3_12 : IN std_logic ;
         d_arr_add_3_11 : IN std_logic ;
         d_arr_add_3_10 : IN std_logic ;
         d_arr_add_3_9 : IN std_logic ;
         d_arr_add_3_8 : IN std_logic ;
         d_arr_add_3_7 : IN std_logic ;
         d_arr_add_3_6 : IN std_logic ;
         d_arr_add_3_5 : IN std_logic ;
         d_arr_add_3_4 : IN std_logic ;
         d_arr_add_3_3 : IN std_logic ;
         d_arr_add_3_2 : IN std_logic ;
         d_arr_add_3_1 : IN std_logic ;
         d_arr_add_3_0 : IN std_logic ;
         d_arr_add_4_31 : IN std_logic ;
         d_arr_add_4_30 : IN std_logic ;
         d_arr_add_4_29 : IN std_logic ;
         d_arr_add_4_28 : IN std_logic ;
         d_arr_add_4_27 : IN std_logic ;
         d_arr_add_4_26 : IN std_logic ;
         d_arr_add_4_25 : IN std_logic ;
         d_arr_add_4_24 : IN std_logic ;
         d_arr_add_4_23 : IN std_logic ;
         d_arr_add_4_22 : IN std_logic ;
         d_arr_add_4_21 : IN std_logic ;
         d_arr_add_4_20 : IN std_logic ;
         d_arr_add_4_19 : IN std_logic ;
         d_arr_add_4_18 : IN std_logic ;
         d_arr_add_4_17 : IN std_logic ;
         d_arr_add_4_16 : IN std_logic ;
         d_arr_add_4_15 : IN std_logic ;
         d_arr_add_4_14 : IN std_logic ;
         d_arr_add_4_13 : IN std_logic ;
         d_arr_add_4_12 : IN std_logic ;
         d_arr_add_4_11 : IN std_logic ;
         d_arr_add_4_10 : IN std_logic ;
         d_arr_add_4_9 : IN std_logic ;
         d_arr_add_4_8 : IN std_logic ;
         d_arr_add_4_7 : IN std_logic ;
         d_arr_add_4_6 : IN std_logic ;
         d_arr_add_4_5 : IN std_logic ;
         d_arr_add_4_4 : IN std_logic ;
         d_arr_add_4_3 : IN std_logic ;
         d_arr_add_4_2 : IN std_logic ;
         d_arr_add_4_1 : IN std_logic ;
         d_arr_add_4_0 : IN std_logic ;
         d_arr_add_5_31 : IN std_logic ;
         d_arr_add_5_30 : IN std_logic ;
         d_arr_add_5_29 : IN std_logic ;
         d_arr_add_5_28 : IN std_logic ;
         d_arr_add_5_27 : IN std_logic ;
         d_arr_add_5_26 : IN std_logic ;
         d_arr_add_5_25 : IN std_logic ;
         d_arr_add_5_24 : IN std_logic ;
         d_arr_add_5_23 : IN std_logic ;
         d_arr_add_5_22 : IN std_logic ;
         d_arr_add_5_21 : IN std_logic ;
         d_arr_add_5_20 : IN std_logic ;
         d_arr_add_5_19 : IN std_logic ;
         d_arr_add_5_18 : IN std_logic ;
         d_arr_add_5_17 : IN std_logic ;
         d_arr_add_5_16 : IN std_logic ;
         d_arr_add_5_15 : IN std_logic ;
         d_arr_add_5_14 : IN std_logic ;
         d_arr_add_5_13 : IN std_logic ;
         d_arr_add_5_12 : IN std_logic ;
         d_arr_add_5_11 : IN std_logic ;
         d_arr_add_5_10 : IN std_logic ;
         d_arr_add_5_9 : IN std_logic ;
         d_arr_add_5_8 : IN std_logic ;
         d_arr_add_5_7 : IN std_logic ;
         d_arr_add_5_6 : IN std_logic ;
         d_arr_add_5_5 : IN std_logic ;
         d_arr_add_5_4 : IN std_logic ;
         d_arr_add_5_3 : IN std_logic ;
         d_arr_add_5_2 : IN std_logic ;
         d_arr_add_5_1 : IN std_logic ;
         d_arr_add_5_0 : IN std_logic ;
         d_arr_add_6_31 : IN std_logic ;
         d_arr_add_6_30 : IN std_logic ;
         d_arr_add_6_29 : IN std_logic ;
         d_arr_add_6_28 : IN std_logic ;
         d_arr_add_6_27 : IN std_logic ;
         d_arr_add_6_26 : IN std_logic ;
         d_arr_add_6_25 : IN std_logic ;
         d_arr_add_6_24 : IN std_logic ;
         d_arr_add_6_23 : IN std_logic ;
         d_arr_add_6_22 : IN std_logic ;
         d_arr_add_6_21 : IN std_logic ;
         d_arr_add_6_20 : IN std_logic ;
         d_arr_add_6_19 : IN std_logic ;
         d_arr_add_6_18 : IN std_logic ;
         d_arr_add_6_17 : IN std_logic ;
         d_arr_add_6_16 : IN std_logic ;
         d_arr_add_6_15 : IN std_logic ;
         d_arr_add_6_14 : IN std_logic ;
         d_arr_add_6_13 : IN std_logic ;
         d_arr_add_6_12 : IN std_logic ;
         d_arr_add_6_11 : IN std_logic ;
         d_arr_add_6_10 : IN std_logic ;
         d_arr_add_6_9 : IN std_logic ;
         d_arr_add_6_8 : IN std_logic ;
         d_arr_add_6_7 : IN std_logic ;
         d_arr_add_6_6 : IN std_logic ;
         d_arr_add_6_5 : IN std_logic ;
         d_arr_add_6_4 : IN std_logic ;
         d_arr_add_6_3 : IN std_logic ;
         d_arr_add_6_2 : IN std_logic ;
         d_arr_add_6_1 : IN std_logic ;
         d_arr_add_6_0 : IN std_logic ;
         d_arr_add_7_31 : IN std_logic ;
         d_arr_add_7_30 : IN std_logic ;
         d_arr_add_7_29 : IN std_logic ;
         d_arr_add_7_28 : IN std_logic ;
         d_arr_add_7_27 : IN std_logic ;
         d_arr_add_7_26 : IN std_logic ;
         d_arr_add_7_25 : IN std_logic ;
         d_arr_add_7_24 : IN std_logic ;
         d_arr_add_7_23 : IN std_logic ;
         d_arr_add_7_22 : IN std_logic ;
         d_arr_add_7_21 : IN std_logic ;
         d_arr_add_7_20 : IN std_logic ;
         d_arr_add_7_19 : IN std_logic ;
         d_arr_add_7_18 : IN std_logic ;
         d_arr_add_7_17 : IN std_logic ;
         d_arr_add_7_16 : IN std_logic ;
         d_arr_add_7_15 : IN std_logic ;
         d_arr_add_7_14 : IN std_logic ;
         d_arr_add_7_13 : IN std_logic ;
         d_arr_add_7_12 : IN std_logic ;
         d_arr_add_7_11 : IN std_logic ;
         d_arr_add_7_10 : IN std_logic ;
         d_arr_add_7_9 : IN std_logic ;
         d_arr_add_7_8 : IN std_logic ;
         d_arr_add_7_7 : IN std_logic ;
         d_arr_add_7_6 : IN std_logic ;
         d_arr_add_7_5 : IN std_logic ;
         d_arr_add_7_4 : IN std_logic ;
         d_arr_add_7_3 : IN std_logic ;
         d_arr_add_7_2 : IN std_logic ;
         d_arr_add_7_1 : IN std_logic ;
         d_arr_add_7_0 : IN std_logic ;
         d_arr_add_8_31 : IN std_logic ;
         d_arr_add_8_30 : IN std_logic ;
         d_arr_add_8_29 : IN std_logic ;
         d_arr_add_8_28 : IN std_logic ;
         d_arr_add_8_27 : IN std_logic ;
         d_arr_add_8_26 : IN std_logic ;
         d_arr_add_8_25 : IN std_logic ;
         d_arr_add_8_24 : IN std_logic ;
         d_arr_add_8_23 : IN std_logic ;
         d_arr_add_8_22 : IN std_logic ;
         d_arr_add_8_21 : IN std_logic ;
         d_arr_add_8_20 : IN std_logic ;
         d_arr_add_8_19 : IN std_logic ;
         d_arr_add_8_18 : IN std_logic ;
         d_arr_add_8_17 : IN std_logic ;
         d_arr_add_8_16 : IN std_logic ;
         d_arr_add_8_15 : IN std_logic ;
         d_arr_add_8_14 : IN std_logic ;
         d_arr_add_8_13 : IN std_logic ;
         d_arr_add_8_12 : IN std_logic ;
         d_arr_add_8_11 : IN std_logic ;
         d_arr_add_8_10 : IN std_logic ;
         d_arr_add_8_9 : IN std_logic ;
         d_arr_add_8_8 : IN std_logic ;
         d_arr_add_8_7 : IN std_logic ;
         d_arr_add_8_6 : IN std_logic ;
         d_arr_add_8_5 : IN std_logic ;
         d_arr_add_8_4 : IN std_logic ;
         d_arr_add_8_3 : IN std_logic ;
         d_arr_add_8_2 : IN std_logic ;
         d_arr_add_8_1 : IN std_logic ;
         d_arr_add_8_0 : IN std_logic ;
         d_arr_add_9_31 : IN std_logic ;
         d_arr_add_9_30 : IN std_logic ;
         d_arr_add_9_29 : IN std_logic ;
         d_arr_add_9_28 : IN std_logic ;
         d_arr_add_9_27 : IN std_logic ;
         d_arr_add_9_26 : IN std_logic ;
         d_arr_add_9_25 : IN std_logic ;
         d_arr_add_9_24 : IN std_logic ;
         d_arr_add_9_23 : IN std_logic ;
         d_arr_add_9_22 : IN std_logic ;
         d_arr_add_9_21 : IN std_logic ;
         d_arr_add_9_20 : IN std_logic ;
         d_arr_add_9_19 : IN std_logic ;
         d_arr_add_9_18 : IN std_logic ;
         d_arr_add_9_17 : IN std_logic ;
         d_arr_add_9_16 : IN std_logic ;
         d_arr_add_9_15 : IN std_logic ;
         d_arr_add_9_14 : IN std_logic ;
         d_arr_add_9_13 : IN std_logic ;
         d_arr_add_9_12 : IN std_logic ;
         d_arr_add_9_11 : IN std_logic ;
         d_arr_add_9_10 : IN std_logic ;
         d_arr_add_9_9 : IN std_logic ;
         d_arr_add_9_8 : IN std_logic ;
         d_arr_add_9_7 : IN std_logic ;
         d_arr_add_9_6 : IN std_logic ;
         d_arr_add_9_5 : IN std_logic ;
         d_arr_add_9_4 : IN std_logic ;
         d_arr_add_9_3 : IN std_logic ;
         d_arr_add_9_2 : IN std_logic ;
         d_arr_add_9_1 : IN std_logic ;
         d_arr_add_9_0 : IN std_logic ;
         d_arr_add_10_31 : IN std_logic ;
         d_arr_add_10_30 : IN std_logic ;
         d_arr_add_10_29 : IN std_logic ;
         d_arr_add_10_28 : IN std_logic ;
         d_arr_add_10_27 : IN std_logic ;
         d_arr_add_10_26 : IN std_logic ;
         d_arr_add_10_25 : IN std_logic ;
         d_arr_add_10_24 : IN std_logic ;
         d_arr_add_10_23 : IN std_logic ;
         d_arr_add_10_22 : IN std_logic ;
         d_arr_add_10_21 : IN std_logic ;
         d_arr_add_10_20 : IN std_logic ;
         d_arr_add_10_19 : IN std_logic ;
         d_arr_add_10_18 : IN std_logic ;
         d_arr_add_10_17 : IN std_logic ;
         d_arr_add_10_16 : IN std_logic ;
         d_arr_add_10_15 : IN std_logic ;
         d_arr_add_10_14 : IN std_logic ;
         d_arr_add_10_13 : IN std_logic ;
         d_arr_add_10_12 : IN std_logic ;
         d_arr_add_10_11 : IN std_logic ;
         d_arr_add_10_10 : IN std_logic ;
         d_arr_add_10_9 : IN std_logic ;
         d_arr_add_10_8 : IN std_logic ;
         d_arr_add_10_7 : IN std_logic ;
         d_arr_add_10_6 : IN std_logic ;
         d_arr_add_10_5 : IN std_logic ;
         d_arr_add_10_4 : IN std_logic ;
         d_arr_add_10_3 : IN std_logic ;
         d_arr_add_10_2 : IN std_logic ;
         d_arr_add_10_1 : IN std_logic ;
         d_arr_add_10_0 : IN std_logic ;
         d_arr_add_11_31 : IN std_logic ;
         d_arr_add_11_30 : IN std_logic ;
         d_arr_add_11_29 : IN std_logic ;
         d_arr_add_11_28 : IN std_logic ;
         d_arr_add_11_27 : IN std_logic ;
         d_arr_add_11_26 : IN std_logic ;
         d_arr_add_11_25 : IN std_logic ;
         d_arr_add_11_24 : IN std_logic ;
         d_arr_add_11_23 : IN std_logic ;
         d_arr_add_11_22 : IN std_logic ;
         d_arr_add_11_21 : IN std_logic ;
         d_arr_add_11_20 : IN std_logic ;
         d_arr_add_11_19 : IN std_logic ;
         d_arr_add_11_18 : IN std_logic ;
         d_arr_add_11_17 : IN std_logic ;
         d_arr_add_11_16 : IN std_logic ;
         d_arr_add_11_15 : IN std_logic ;
         d_arr_add_11_14 : IN std_logic ;
         d_arr_add_11_13 : IN std_logic ;
         d_arr_add_11_12 : IN std_logic ;
         d_arr_add_11_11 : IN std_logic ;
         d_arr_add_11_10 : IN std_logic ;
         d_arr_add_11_9 : IN std_logic ;
         d_arr_add_11_8 : IN std_logic ;
         d_arr_add_11_7 : IN std_logic ;
         d_arr_add_11_6 : IN std_logic ;
         d_arr_add_11_5 : IN std_logic ;
         d_arr_add_11_4 : IN std_logic ;
         d_arr_add_11_3 : IN std_logic ;
         d_arr_add_11_2 : IN std_logic ;
         d_arr_add_11_1 : IN std_logic ;
         d_arr_add_11_0 : IN std_logic ;
         d_arr_add_12_31 : IN std_logic ;
         d_arr_add_12_30 : IN std_logic ;
         d_arr_add_12_29 : IN std_logic ;
         d_arr_add_12_28 : IN std_logic ;
         d_arr_add_12_27 : IN std_logic ;
         d_arr_add_12_26 : IN std_logic ;
         d_arr_add_12_25 : IN std_logic ;
         d_arr_add_12_24 : IN std_logic ;
         d_arr_add_12_23 : IN std_logic ;
         d_arr_add_12_22 : IN std_logic ;
         d_arr_add_12_21 : IN std_logic ;
         d_arr_add_12_20 : IN std_logic ;
         d_arr_add_12_19 : IN std_logic ;
         d_arr_add_12_18 : IN std_logic ;
         d_arr_add_12_17 : IN std_logic ;
         d_arr_add_12_16 : IN std_logic ;
         d_arr_add_12_15 : IN std_logic ;
         d_arr_add_12_14 : IN std_logic ;
         d_arr_add_12_13 : IN std_logic ;
         d_arr_add_12_12 : IN std_logic ;
         d_arr_add_12_11 : IN std_logic ;
         d_arr_add_12_10 : IN std_logic ;
         d_arr_add_12_9 : IN std_logic ;
         d_arr_add_12_8 : IN std_logic ;
         d_arr_add_12_7 : IN std_logic ;
         d_arr_add_12_6 : IN std_logic ;
         d_arr_add_12_5 : IN std_logic ;
         d_arr_add_12_4 : IN std_logic ;
         d_arr_add_12_3 : IN std_logic ;
         d_arr_add_12_2 : IN std_logic ;
         d_arr_add_12_1 : IN std_logic ;
         d_arr_add_12_0 : IN std_logic ;
         d_arr_add_13_31 : IN std_logic ;
         d_arr_add_13_30 : IN std_logic ;
         d_arr_add_13_29 : IN std_logic ;
         d_arr_add_13_28 : IN std_logic ;
         d_arr_add_13_27 : IN std_logic ;
         d_arr_add_13_26 : IN std_logic ;
         d_arr_add_13_25 : IN std_logic ;
         d_arr_add_13_24 : IN std_logic ;
         d_arr_add_13_23 : IN std_logic ;
         d_arr_add_13_22 : IN std_logic ;
         d_arr_add_13_21 : IN std_logic ;
         d_arr_add_13_20 : IN std_logic ;
         d_arr_add_13_19 : IN std_logic ;
         d_arr_add_13_18 : IN std_logic ;
         d_arr_add_13_17 : IN std_logic ;
         d_arr_add_13_16 : IN std_logic ;
         d_arr_add_13_15 : IN std_logic ;
         d_arr_add_13_14 : IN std_logic ;
         d_arr_add_13_13 : IN std_logic ;
         d_arr_add_13_12 : IN std_logic ;
         d_arr_add_13_11 : IN std_logic ;
         d_arr_add_13_10 : IN std_logic ;
         d_arr_add_13_9 : IN std_logic ;
         d_arr_add_13_8 : IN std_logic ;
         d_arr_add_13_7 : IN std_logic ;
         d_arr_add_13_6 : IN std_logic ;
         d_arr_add_13_5 : IN std_logic ;
         d_arr_add_13_4 : IN std_logic ;
         d_arr_add_13_3 : IN std_logic ;
         d_arr_add_13_2 : IN std_logic ;
         d_arr_add_13_1 : IN std_logic ;
         d_arr_add_13_0 : IN std_logic ;
         d_arr_add_14_31 : IN std_logic ;
         d_arr_add_14_30 : IN std_logic ;
         d_arr_add_14_29 : IN std_logic ;
         d_arr_add_14_28 : IN std_logic ;
         d_arr_add_14_27 : IN std_logic ;
         d_arr_add_14_26 : IN std_logic ;
         d_arr_add_14_25 : IN std_logic ;
         d_arr_add_14_24 : IN std_logic ;
         d_arr_add_14_23 : IN std_logic ;
         d_arr_add_14_22 : IN std_logic ;
         d_arr_add_14_21 : IN std_logic ;
         d_arr_add_14_20 : IN std_logic ;
         d_arr_add_14_19 : IN std_logic ;
         d_arr_add_14_18 : IN std_logic ;
         d_arr_add_14_17 : IN std_logic ;
         d_arr_add_14_16 : IN std_logic ;
         d_arr_add_14_15 : IN std_logic ;
         d_arr_add_14_14 : IN std_logic ;
         d_arr_add_14_13 : IN std_logic ;
         d_arr_add_14_12 : IN std_logic ;
         d_arr_add_14_11 : IN std_logic ;
         d_arr_add_14_10 : IN std_logic ;
         d_arr_add_14_9 : IN std_logic ;
         d_arr_add_14_8 : IN std_logic ;
         d_arr_add_14_7 : IN std_logic ;
         d_arr_add_14_6 : IN std_logic ;
         d_arr_add_14_5 : IN std_logic ;
         d_arr_add_14_4 : IN std_logic ;
         d_arr_add_14_3 : IN std_logic ;
         d_arr_add_14_2 : IN std_logic ;
         d_arr_add_14_1 : IN std_logic ;
         d_arr_add_14_0 : IN std_logic ;
         d_arr_add_15_31 : IN std_logic ;
         d_arr_add_15_30 : IN std_logic ;
         d_arr_add_15_29 : IN std_logic ;
         d_arr_add_15_28 : IN std_logic ;
         d_arr_add_15_27 : IN std_logic ;
         d_arr_add_15_26 : IN std_logic ;
         d_arr_add_15_25 : IN std_logic ;
         d_arr_add_15_24 : IN std_logic ;
         d_arr_add_15_23 : IN std_logic ;
         d_arr_add_15_22 : IN std_logic ;
         d_arr_add_15_21 : IN std_logic ;
         d_arr_add_15_20 : IN std_logic ;
         d_arr_add_15_19 : IN std_logic ;
         d_arr_add_15_18 : IN std_logic ;
         d_arr_add_15_17 : IN std_logic ;
         d_arr_add_15_16 : IN std_logic ;
         d_arr_add_15_15 : IN std_logic ;
         d_arr_add_15_14 : IN std_logic ;
         d_arr_add_15_13 : IN std_logic ;
         d_arr_add_15_12 : IN std_logic ;
         d_arr_add_15_11 : IN std_logic ;
         d_arr_add_15_10 : IN std_logic ;
         d_arr_add_15_9 : IN std_logic ;
         d_arr_add_15_8 : IN std_logic ;
         d_arr_add_15_7 : IN std_logic ;
         d_arr_add_15_6 : IN std_logic ;
         d_arr_add_15_5 : IN std_logic ;
         d_arr_add_15_4 : IN std_logic ;
         d_arr_add_15_3 : IN std_logic ;
         d_arr_add_15_2 : IN std_logic ;
         d_arr_add_15_1 : IN std_logic ;
         d_arr_add_15_0 : IN std_logic ;
         d_arr_add_16_31 : IN std_logic ;
         d_arr_add_16_30 : IN std_logic ;
         d_arr_add_16_29 : IN std_logic ;
         d_arr_add_16_28 : IN std_logic ;
         d_arr_add_16_27 : IN std_logic ;
         d_arr_add_16_26 : IN std_logic ;
         d_arr_add_16_25 : IN std_logic ;
         d_arr_add_16_24 : IN std_logic ;
         d_arr_add_16_23 : IN std_logic ;
         d_arr_add_16_22 : IN std_logic ;
         d_arr_add_16_21 : IN std_logic ;
         d_arr_add_16_20 : IN std_logic ;
         d_arr_add_16_19 : IN std_logic ;
         d_arr_add_16_18 : IN std_logic ;
         d_arr_add_16_17 : IN std_logic ;
         d_arr_add_16_16 : IN std_logic ;
         d_arr_add_16_15 : IN std_logic ;
         d_arr_add_16_14 : IN std_logic ;
         d_arr_add_16_13 : IN std_logic ;
         d_arr_add_16_12 : IN std_logic ;
         d_arr_add_16_11 : IN std_logic ;
         d_arr_add_16_10 : IN std_logic ;
         d_arr_add_16_9 : IN std_logic ;
         d_arr_add_16_8 : IN std_logic ;
         d_arr_add_16_7 : IN std_logic ;
         d_arr_add_16_6 : IN std_logic ;
         d_arr_add_16_5 : IN std_logic ;
         d_arr_add_16_4 : IN std_logic ;
         d_arr_add_16_3 : IN std_logic ;
         d_arr_add_16_2 : IN std_logic ;
         d_arr_add_16_1 : IN std_logic ;
         d_arr_add_16_0 : IN std_logic ;
         d_arr_add_17_31 : IN std_logic ;
         d_arr_add_17_30 : IN std_logic ;
         d_arr_add_17_29 : IN std_logic ;
         d_arr_add_17_28 : IN std_logic ;
         d_arr_add_17_27 : IN std_logic ;
         d_arr_add_17_26 : IN std_logic ;
         d_arr_add_17_25 : IN std_logic ;
         d_arr_add_17_24 : IN std_logic ;
         d_arr_add_17_23 : IN std_logic ;
         d_arr_add_17_22 : IN std_logic ;
         d_arr_add_17_21 : IN std_logic ;
         d_arr_add_17_20 : IN std_logic ;
         d_arr_add_17_19 : IN std_logic ;
         d_arr_add_17_18 : IN std_logic ;
         d_arr_add_17_17 : IN std_logic ;
         d_arr_add_17_16 : IN std_logic ;
         d_arr_add_17_15 : IN std_logic ;
         d_arr_add_17_14 : IN std_logic ;
         d_arr_add_17_13 : IN std_logic ;
         d_arr_add_17_12 : IN std_logic ;
         d_arr_add_17_11 : IN std_logic ;
         d_arr_add_17_10 : IN std_logic ;
         d_arr_add_17_9 : IN std_logic ;
         d_arr_add_17_8 : IN std_logic ;
         d_arr_add_17_7 : IN std_logic ;
         d_arr_add_17_6 : IN std_logic ;
         d_arr_add_17_5 : IN std_logic ;
         d_arr_add_17_4 : IN std_logic ;
         d_arr_add_17_3 : IN std_logic ;
         d_arr_add_17_2 : IN std_logic ;
         d_arr_add_17_1 : IN std_logic ;
         d_arr_add_17_0 : IN std_logic ;
         d_arr_add_18_31 : IN std_logic ;
         d_arr_add_18_30 : IN std_logic ;
         d_arr_add_18_29 : IN std_logic ;
         d_arr_add_18_28 : IN std_logic ;
         d_arr_add_18_27 : IN std_logic ;
         d_arr_add_18_26 : IN std_logic ;
         d_arr_add_18_25 : IN std_logic ;
         d_arr_add_18_24 : IN std_logic ;
         d_arr_add_18_23 : IN std_logic ;
         d_arr_add_18_22 : IN std_logic ;
         d_arr_add_18_21 : IN std_logic ;
         d_arr_add_18_20 : IN std_logic ;
         d_arr_add_18_19 : IN std_logic ;
         d_arr_add_18_18 : IN std_logic ;
         d_arr_add_18_17 : IN std_logic ;
         d_arr_add_18_16 : IN std_logic ;
         d_arr_add_18_15 : IN std_logic ;
         d_arr_add_18_14 : IN std_logic ;
         d_arr_add_18_13 : IN std_logic ;
         d_arr_add_18_12 : IN std_logic ;
         d_arr_add_18_11 : IN std_logic ;
         d_arr_add_18_10 : IN std_logic ;
         d_arr_add_18_9 : IN std_logic ;
         d_arr_add_18_8 : IN std_logic ;
         d_arr_add_18_7 : IN std_logic ;
         d_arr_add_18_6 : IN std_logic ;
         d_arr_add_18_5 : IN std_logic ;
         d_arr_add_18_4 : IN std_logic ;
         d_arr_add_18_3 : IN std_logic ;
         d_arr_add_18_2 : IN std_logic ;
         d_arr_add_18_1 : IN std_logic ;
         d_arr_add_18_0 : IN std_logic ;
         d_arr_add_19_31 : IN std_logic ;
         d_arr_add_19_30 : IN std_logic ;
         d_arr_add_19_29 : IN std_logic ;
         d_arr_add_19_28 : IN std_logic ;
         d_arr_add_19_27 : IN std_logic ;
         d_arr_add_19_26 : IN std_logic ;
         d_arr_add_19_25 : IN std_logic ;
         d_arr_add_19_24 : IN std_logic ;
         d_arr_add_19_23 : IN std_logic ;
         d_arr_add_19_22 : IN std_logic ;
         d_arr_add_19_21 : IN std_logic ;
         d_arr_add_19_20 : IN std_logic ;
         d_arr_add_19_19 : IN std_logic ;
         d_arr_add_19_18 : IN std_logic ;
         d_arr_add_19_17 : IN std_logic ;
         d_arr_add_19_16 : IN std_logic ;
         d_arr_add_19_15 : IN std_logic ;
         d_arr_add_19_14 : IN std_logic ;
         d_arr_add_19_13 : IN std_logic ;
         d_arr_add_19_12 : IN std_logic ;
         d_arr_add_19_11 : IN std_logic ;
         d_arr_add_19_10 : IN std_logic ;
         d_arr_add_19_9 : IN std_logic ;
         d_arr_add_19_8 : IN std_logic ;
         d_arr_add_19_7 : IN std_logic ;
         d_arr_add_19_6 : IN std_logic ;
         d_arr_add_19_5 : IN std_logic ;
         d_arr_add_19_4 : IN std_logic ;
         d_arr_add_19_3 : IN std_logic ;
         d_arr_add_19_2 : IN std_logic ;
         d_arr_add_19_1 : IN std_logic ;
         d_arr_add_19_0 : IN std_logic ;
         d_arr_add_20_31 : IN std_logic ;
         d_arr_add_20_30 : IN std_logic ;
         d_arr_add_20_29 : IN std_logic ;
         d_arr_add_20_28 : IN std_logic ;
         d_arr_add_20_27 : IN std_logic ;
         d_arr_add_20_26 : IN std_logic ;
         d_arr_add_20_25 : IN std_logic ;
         d_arr_add_20_24 : IN std_logic ;
         d_arr_add_20_23 : IN std_logic ;
         d_arr_add_20_22 : IN std_logic ;
         d_arr_add_20_21 : IN std_logic ;
         d_arr_add_20_20 : IN std_logic ;
         d_arr_add_20_19 : IN std_logic ;
         d_arr_add_20_18 : IN std_logic ;
         d_arr_add_20_17 : IN std_logic ;
         d_arr_add_20_16 : IN std_logic ;
         d_arr_add_20_15 : IN std_logic ;
         d_arr_add_20_14 : IN std_logic ;
         d_arr_add_20_13 : IN std_logic ;
         d_arr_add_20_12 : IN std_logic ;
         d_arr_add_20_11 : IN std_logic ;
         d_arr_add_20_10 : IN std_logic ;
         d_arr_add_20_9 : IN std_logic ;
         d_arr_add_20_8 : IN std_logic ;
         d_arr_add_20_7 : IN std_logic ;
         d_arr_add_20_6 : IN std_logic ;
         d_arr_add_20_5 : IN std_logic ;
         d_arr_add_20_4 : IN std_logic ;
         d_arr_add_20_3 : IN std_logic ;
         d_arr_add_20_2 : IN std_logic ;
         d_arr_add_20_1 : IN std_logic ;
         d_arr_add_20_0 : IN std_logic ;
         d_arr_add_21_31 : IN std_logic ;
         d_arr_add_21_30 : IN std_logic ;
         d_arr_add_21_29 : IN std_logic ;
         d_arr_add_21_28 : IN std_logic ;
         d_arr_add_21_27 : IN std_logic ;
         d_arr_add_21_26 : IN std_logic ;
         d_arr_add_21_25 : IN std_logic ;
         d_arr_add_21_24 : IN std_logic ;
         d_arr_add_21_23 : IN std_logic ;
         d_arr_add_21_22 : IN std_logic ;
         d_arr_add_21_21 : IN std_logic ;
         d_arr_add_21_20 : IN std_logic ;
         d_arr_add_21_19 : IN std_logic ;
         d_arr_add_21_18 : IN std_logic ;
         d_arr_add_21_17 : IN std_logic ;
         d_arr_add_21_16 : IN std_logic ;
         d_arr_add_21_15 : IN std_logic ;
         d_arr_add_21_14 : IN std_logic ;
         d_arr_add_21_13 : IN std_logic ;
         d_arr_add_21_12 : IN std_logic ;
         d_arr_add_21_11 : IN std_logic ;
         d_arr_add_21_10 : IN std_logic ;
         d_arr_add_21_9 : IN std_logic ;
         d_arr_add_21_8 : IN std_logic ;
         d_arr_add_21_7 : IN std_logic ;
         d_arr_add_21_6 : IN std_logic ;
         d_arr_add_21_5 : IN std_logic ;
         d_arr_add_21_4 : IN std_logic ;
         d_arr_add_21_3 : IN std_logic ;
         d_arr_add_21_2 : IN std_logic ;
         d_arr_add_21_1 : IN std_logic ;
         d_arr_add_21_0 : IN std_logic ;
         d_arr_add_22_31 : IN std_logic ;
         d_arr_add_22_30 : IN std_logic ;
         d_arr_add_22_29 : IN std_logic ;
         d_arr_add_22_28 : IN std_logic ;
         d_arr_add_22_27 : IN std_logic ;
         d_arr_add_22_26 : IN std_logic ;
         d_arr_add_22_25 : IN std_logic ;
         d_arr_add_22_24 : IN std_logic ;
         d_arr_add_22_23 : IN std_logic ;
         d_arr_add_22_22 : IN std_logic ;
         d_arr_add_22_21 : IN std_logic ;
         d_arr_add_22_20 : IN std_logic ;
         d_arr_add_22_19 : IN std_logic ;
         d_arr_add_22_18 : IN std_logic ;
         d_arr_add_22_17 : IN std_logic ;
         d_arr_add_22_16 : IN std_logic ;
         d_arr_add_22_15 : IN std_logic ;
         d_arr_add_22_14 : IN std_logic ;
         d_arr_add_22_13 : IN std_logic ;
         d_arr_add_22_12 : IN std_logic ;
         d_arr_add_22_11 : IN std_logic ;
         d_arr_add_22_10 : IN std_logic ;
         d_arr_add_22_9 : IN std_logic ;
         d_arr_add_22_8 : IN std_logic ;
         d_arr_add_22_7 : IN std_logic ;
         d_arr_add_22_6 : IN std_logic ;
         d_arr_add_22_5 : IN std_logic ;
         d_arr_add_22_4 : IN std_logic ;
         d_arr_add_22_3 : IN std_logic ;
         d_arr_add_22_2 : IN std_logic ;
         d_arr_add_22_1 : IN std_logic ;
         d_arr_add_22_0 : IN std_logic ;
         d_arr_add_23_31 : IN std_logic ;
         d_arr_add_23_30 : IN std_logic ;
         d_arr_add_23_29 : IN std_logic ;
         d_arr_add_23_28 : IN std_logic ;
         d_arr_add_23_27 : IN std_logic ;
         d_arr_add_23_26 : IN std_logic ;
         d_arr_add_23_25 : IN std_logic ;
         d_arr_add_23_24 : IN std_logic ;
         d_arr_add_23_23 : IN std_logic ;
         d_arr_add_23_22 : IN std_logic ;
         d_arr_add_23_21 : IN std_logic ;
         d_arr_add_23_20 : IN std_logic ;
         d_arr_add_23_19 : IN std_logic ;
         d_arr_add_23_18 : IN std_logic ;
         d_arr_add_23_17 : IN std_logic ;
         d_arr_add_23_16 : IN std_logic ;
         d_arr_add_23_15 : IN std_logic ;
         d_arr_add_23_14 : IN std_logic ;
         d_arr_add_23_13 : IN std_logic ;
         d_arr_add_23_12 : IN std_logic ;
         d_arr_add_23_11 : IN std_logic ;
         d_arr_add_23_10 : IN std_logic ;
         d_arr_add_23_9 : IN std_logic ;
         d_arr_add_23_8 : IN std_logic ;
         d_arr_add_23_7 : IN std_logic ;
         d_arr_add_23_6 : IN std_logic ;
         d_arr_add_23_5 : IN std_logic ;
         d_arr_add_23_4 : IN std_logic ;
         d_arr_add_23_3 : IN std_logic ;
         d_arr_add_23_2 : IN std_logic ;
         d_arr_add_23_1 : IN std_logic ;
         d_arr_add_23_0 : IN std_logic ;
         d_arr_add_24_31 : IN std_logic ;
         d_arr_add_24_30 : IN std_logic ;
         d_arr_add_24_29 : IN std_logic ;
         d_arr_add_24_28 : IN std_logic ;
         d_arr_add_24_27 : IN std_logic ;
         d_arr_add_24_26 : IN std_logic ;
         d_arr_add_24_25 : IN std_logic ;
         d_arr_add_24_24 : IN std_logic ;
         d_arr_add_24_23 : IN std_logic ;
         d_arr_add_24_22 : IN std_logic ;
         d_arr_add_24_21 : IN std_logic ;
         d_arr_add_24_20 : IN std_logic ;
         d_arr_add_24_19 : IN std_logic ;
         d_arr_add_24_18 : IN std_logic ;
         d_arr_add_24_17 : IN std_logic ;
         d_arr_add_24_16 : IN std_logic ;
         d_arr_add_24_15 : IN std_logic ;
         d_arr_add_24_14 : IN std_logic ;
         d_arr_add_24_13 : IN std_logic ;
         d_arr_add_24_12 : IN std_logic ;
         d_arr_add_24_11 : IN std_logic ;
         d_arr_add_24_10 : IN std_logic ;
         d_arr_add_24_9 : IN std_logic ;
         d_arr_add_24_8 : IN std_logic ;
         d_arr_add_24_7 : IN std_logic ;
         d_arr_add_24_6 : IN std_logic ;
         d_arr_add_24_5 : IN std_logic ;
         d_arr_add_24_4 : IN std_logic ;
         d_arr_add_24_3 : IN std_logic ;
         d_arr_add_24_2 : IN std_logic ;
         d_arr_add_24_1 : IN std_logic ;
         d_arr_add_24_0 : IN std_logic ;
         d_arr_merge1_0_31 : IN std_logic ;
         d_arr_merge1_0_30 : IN std_logic ;
         d_arr_merge1_0_29 : IN std_logic ;
         d_arr_merge1_0_28 : IN std_logic ;
         d_arr_merge1_0_27 : IN std_logic ;
         d_arr_merge1_0_26 : IN std_logic ;
         d_arr_merge1_0_25 : IN std_logic ;
         d_arr_merge1_0_24 : IN std_logic ;
         d_arr_merge1_0_23 : IN std_logic ;
         d_arr_merge1_0_22 : IN std_logic ;
         d_arr_merge1_0_21 : IN std_logic ;
         d_arr_merge1_0_20 : IN std_logic ;
         d_arr_merge1_0_19 : IN std_logic ;
         d_arr_merge1_0_18 : IN std_logic ;
         d_arr_merge1_0_17 : IN std_logic ;
         d_arr_merge1_0_16 : IN std_logic ;
         d_arr_merge1_0_15 : IN std_logic ;
         d_arr_merge1_0_14 : IN std_logic ;
         d_arr_merge1_0_13 : IN std_logic ;
         d_arr_merge1_0_12 : IN std_logic ;
         d_arr_merge1_0_11 : IN std_logic ;
         d_arr_merge1_0_10 : IN std_logic ;
         d_arr_merge1_0_9 : IN std_logic ;
         d_arr_merge1_0_8 : IN std_logic ;
         d_arr_merge1_0_7 : IN std_logic ;
         d_arr_merge1_0_6 : IN std_logic ;
         d_arr_merge1_0_5 : IN std_logic ;
         d_arr_merge1_0_4 : IN std_logic ;
         d_arr_merge1_0_3 : IN std_logic ;
         d_arr_merge1_0_2 : IN std_logic ;
         d_arr_merge1_0_1 : IN std_logic ;
         d_arr_merge1_0_0 : IN std_logic ;
         d_arr_merge1_1_31 : IN std_logic ;
         d_arr_merge1_1_30 : IN std_logic ;
         d_arr_merge1_1_29 : IN std_logic ;
         d_arr_merge1_1_28 : IN std_logic ;
         d_arr_merge1_1_27 : IN std_logic ;
         d_arr_merge1_1_26 : IN std_logic ;
         d_arr_merge1_1_25 : IN std_logic ;
         d_arr_merge1_1_24 : IN std_logic ;
         d_arr_merge1_1_23 : IN std_logic ;
         d_arr_merge1_1_22 : IN std_logic ;
         d_arr_merge1_1_21 : IN std_logic ;
         d_arr_merge1_1_20 : IN std_logic ;
         d_arr_merge1_1_19 : IN std_logic ;
         d_arr_merge1_1_18 : IN std_logic ;
         d_arr_merge1_1_17 : IN std_logic ;
         d_arr_merge1_1_16 : IN std_logic ;
         d_arr_merge1_1_15 : IN std_logic ;
         d_arr_merge1_1_14 : IN std_logic ;
         d_arr_merge1_1_13 : IN std_logic ;
         d_arr_merge1_1_12 : IN std_logic ;
         d_arr_merge1_1_11 : IN std_logic ;
         d_arr_merge1_1_10 : IN std_logic ;
         d_arr_merge1_1_9 : IN std_logic ;
         d_arr_merge1_1_8 : IN std_logic ;
         d_arr_merge1_1_7 : IN std_logic ;
         d_arr_merge1_1_6 : IN std_logic ;
         d_arr_merge1_1_5 : IN std_logic ;
         d_arr_merge1_1_4 : IN std_logic ;
         d_arr_merge1_1_3 : IN std_logic ;
         d_arr_merge1_1_2 : IN std_logic ;
         d_arr_merge1_1_1 : IN std_logic ;
         d_arr_merge1_1_0 : IN std_logic ;
         d_arr_merge1_2_31 : IN std_logic ;
         d_arr_merge1_2_30 : IN std_logic ;
         d_arr_merge1_2_29 : IN std_logic ;
         d_arr_merge1_2_28 : IN std_logic ;
         d_arr_merge1_2_27 : IN std_logic ;
         d_arr_merge1_2_26 : IN std_logic ;
         d_arr_merge1_2_25 : IN std_logic ;
         d_arr_merge1_2_24 : IN std_logic ;
         d_arr_merge1_2_23 : IN std_logic ;
         d_arr_merge1_2_22 : IN std_logic ;
         d_arr_merge1_2_21 : IN std_logic ;
         d_arr_merge1_2_20 : IN std_logic ;
         d_arr_merge1_2_19 : IN std_logic ;
         d_arr_merge1_2_18 : IN std_logic ;
         d_arr_merge1_2_17 : IN std_logic ;
         d_arr_merge1_2_16 : IN std_logic ;
         d_arr_merge1_2_15 : IN std_logic ;
         d_arr_merge1_2_14 : IN std_logic ;
         d_arr_merge1_2_13 : IN std_logic ;
         d_arr_merge1_2_12 : IN std_logic ;
         d_arr_merge1_2_11 : IN std_logic ;
         d_arr_merge1_2_10 : IN std_logic ;
         d_arr_merge1_2_9 : IN std_logic ;
         d_arr_merge1_2_8 : IN std_logic ;
         d_arr_merge1_2_7 : IN std_logic ;
         d_arr_merge1_2_6 : IN std_logic ;
         d_arr_merge1_2_5 : IN std_logic ;
         d_arr_merge1_2_4 : IN std_logic ;
         d_arr_merge1_2_3 : IN std_logic ;
         d_arr_merge1_2_2 : IN std_logic ;
         d_arr_merge1_2_1 : IN std_logic ;
         d_arr_merge1_2_0 : IN std_logic ;
         d_arr_merge1_3_31 : IN std_logic ;
         d_arr_merge1_3_30 : IN std_logic ;
         d_arr_merge1_3_29 : IN std_logic ;
         d_arr_merge1_3_28 : IN std_logic ;
         d_arr_merge1_3_27 : IN std_logic ;
         d_arr_merge1_3_26 : IN std_logic ;
         d_arr_merge1_3_25 : IN std_logic ;
         d_arr_merge1_3_24 : IN std_logic ;
         d_arr_merge1_3_23 : IN std_logic ;
         d_arr_merge1_3_22 : IN std_logic ;
         d_arr_merge1_3_21 : IN std_logic ;
         d_arr_merge1_3_20 : IN std_logic ;
         d_arr_merge1_3_19 : IN std_logic ;
         d_arr_merge1_3_18 : IN std_logic ;
         d_arr_merge1_3_17 : IN std_logic ;
         d_arr_merge1_3_16 : IN std_logic ;
         d_arr_merge1_3_15 : IN std_logic ;
         d_arr_merge1_3_14 : IN std_logic ;
         d_arr_merge1_3_13 : IN std_logic ;
         d_arr_merge1_3_12 : IN std_logic ;
         d_arr_merge1_3_11 : IN std_logic ;
         d_arr_merge1_3_10 : IN std_logic ;
         d_arr_merge1_3_9 : IN std_logic ;
         d_arr_merge1_3_8 : IN std_logic ;
         d_arr_merge1_3_7 : IN std_logic ;
         d_arr_merge1_3_6 : IN std_logic ;
         d_arr_merge1_3_5 : IN std_logic ;
         d_arr_merge1_3_4 : IN std_logic ;
         d_arr_merge1_3_3 : IN std_logic ;
         d_arr_merge1_3_2 : IN std_logic ;
         d_arr_merge1_3_1 : IN std_logic ;
         d_arr_merge1_3_0 : IN std_logic ;
         d_arr_merge1_4_31 : IN std_logic ;
         d_arr_merge1_4_30 : IN std_logic ;
         d_arr_merge1_4_29 : IN std_logic ;
         d_arr_merge1_4_28 : IN std_logic ;
         d_arr_merge1_4_27 : IN std_logic ;
         d_arr_merge1_4_26 : IN std_logic ;
         d_arr_merge1_4_25 : IN std_logic ;
         d_arr_merge1_4_24 : IN std_logic ;
         d_arr_merge1_4_23 : IN std_logic ;
         d_arr_merge1_4_22 : IN std_logic ;
         d_arr_merge1_4_21 : IN std_logic ;
         d_arr_merge1_4_20 : IN std_logic ;
         d_arr_merge1_4_19 : IN std_logic ;
         d_arr_merge1_4_18 : IN std_logic ;
         d_arr_merge1_4_17 : IN std_logic ;
         d_arr_merge1_4_16 : IN std_logic ;
         d_arr_merge1_4_15 : IN std_logic ;
         d_arr_merge1_4_14 : IN std_logic ;
         d_arr_merge1_4_13 : IN std_logic ;
         d_arr_merge1_4_12 : IN std_logic ;
         d_arr_merge1_4_11 : IN std_logic ;
         d_arr_merge1_4_10 : IN std_logic ;
         d_arr_merge1_4_9 : IN std_logic ;
         d_arr_merge1_4_8 : IN std_logic ;
         d_arr_merge1_4_7 : IN std_logic ;
         d_arr_merge1_4_6 : IN std_logic ;
         d_arr_merge1_4_5 : IN std_logic ;
         d_arr_merge1_4_4 : IN std_logic ;
         d_arr_merge1_4_3 : IN std_logic ;
         d_arr_merge1_4_2 : IN std_logic ;
         d_arr_merge1_4_1 : IN std_logic ;
         d_arr_merge1_4_0 : IN std_logic ;
         d_arr_merge1_5_31 : IN std_logic ;
         d_arr_merge1_5_30 : IN std_logic ;
         d_arr_merge1_5_29 : IN std_logic ;
         d_arr_merge1_5_28 : IN std_logic ;
         d_arr_merge1_5_27 : IN std_logic ;
         d_arr_merge1_5_26 : IN std_logic ;
         d_arr_merge1_5_25 : IN std_logic ;
         d_arr_merge1_5_24 : IN std_logic ;
         d_arr_merge1_5_23 : IN std_logic ;
         d_arr_merge1_5_22 : IN std_logic ;
         d_arr_merge1_5_21 : IN std_logic ;
         d_arr_merge1_5_20 : IN std_logic ;
         d_arr_merge1_5_19 : IN std_logic ;
         d_arr_merge1_5_18 : IN std_logic ;
         d_arr_merge1_5_17 : IN std_logic ;
         d_arr_merge1_5_16 : IN std_logic ;
         d_arr_merge1_5_15 : IN std_logic ;
         d_arr_merge1_5_14 : IN std_logic ;
         d_arr_merge1_5_13 : IN std_logic ;
         d_arr_merge1_5_12 : IN std_logic ;
         d_arr_merge1_5_11 : IN std_logic ;
         d_arr_merge1_5_10 : IN std_logic ;
         d_arr_merge1_5_9 : IN std_logic ;
         d_arr_merge1_5_8 : IN std_logic ;
         d_arr_merge1_5_7 : IN std_logic ;
         d_arr_merge1_5_6 : IN std_logic ;
         d_arr_merge1_5_5 : IN std_logic ;
         d_arr_merge1_5_4 : IN std_logic ;
         d_arr_merge1_5_3 : IN std_logic ;
         d_arr_merge1_5_2 : IN std_logic ;
         d_arr_merge1_5_1 : IN std_logic ;
         d_arr_merge1_5_0 : IN std_logic ;
         d_arr_merge1_6_31 : IN std_logic ;
         d_arr_merge1_6_30 : IN std_logic ;
         d_arr_merge1_6_29 : IN std_logic ;
         d_arr_merge1_6_28 : IN std_logic ;
         d_arr_merge1_6_27 : IN std_logic ;
         d_arr_merge1_6_26 : IN std_logic ;
         d_arr_merge1_6_25 : IN std_logic ;
         d_arr_merge1_6_24 : IN std_logic ;
         d_arr_merge1_6_23 : IN std_logic ;
         d_arr_merge1_6_22 : IN std_logic ;
         d_arr_merge1_6_21 : IN std_logic ;
         d_arr_merge1_6_20 : IN std_logic ;
         d_arr_merge1_6_19 : IN std_logic ;
         d_arr_merge1_6_18 : IN std_logic ;
         d_arr_merge1_6_17 : IN std_logic ;
         d_arr_merge1_6_16 : IN std_logic ;
         d_arr_merge1_6_15 : IN std_logic ;
         d_arr_merge1_6_14 : IN std_logic ;
         d_arr_merge1_6_13 : IN std_logic ;
         d_arr_merge1_6_12 : IN std_logic ;
         d_arr_merge1_6_11 : IN std_logic ;
         d_arr_merge1_6_10 : IN std_logic ;
         d_arr_merge1_6_9 : IN std_logic ;
         d_arr_merge1_6_8 : IN std_logic ;
         d_arr_merge1_6_7 : IN std_logic ;
         d_arr_merge1_6_6 : IN std_logic ;
         d_arr_merge1_6_5 : IN std_logic ;
         d_arr_merge1_6_4 : IN std_logic ;
         d_arr_merge1_6_3 : IN std_logic ;
         d_arr_merge1_6_2 : IN std_logic ;
         d_arr_merge1_6_1 : IN std_logic ;
         d_arr_merge1_6_0 : IN std_logic ;
         d_arr_merge1_7_31 : IN std_logic ;
         d_arr_merge1_7_30 : IN std_logic ;
         d_arr_merge1_7_29 : IN std_logic ;
         d_arr_merge1_7_28 : IN std_logic ;
         d_arr_merge1_7_27 : IN std_logic ;
         d_arr_merge1_7_26 : IN std_logic ;
         d_arr_merge1_7_25 : IN std_logic ;
         d_arr_merge1_7_24 : IN std_logic ;
         d_arr_merge1_7_23 : IN std_logic ;
         d_arr_merge1_7_22 : IN std_logic ;
         d_arr_merge1_7_21 : IN std_logic ;
         d_arr_merge1_7_20 : IN std_logic ;
         d_arr_merge1_7_19 : IN std_logic ;
         d_arr_merge1_7_18 : IN std_logic ;
         d_arr_merge1_7_17 : IN std_logic ;
         d_arr_merge1_7_16 : IN std_logic ;
         d_arr_merge1_7_15 : IN std_logic ;
         d_arr_merge1_7_14 : IN std_logic ;
         d_arr_merge1_7_13 : IN std_logic ;
         d_arr_merge1_7_12 : IN std_logic ;
         d_arr_merge1_7_11 : IN std_logic ;
         d_arr_merge1_7_10 : IN std_logic ;
         d_arr_merge1_7_9 : IN std_logic ;
         d_arr_merge1_7_8 : IN std_logic ;
         d_arr_merge1_7_7 : IN std_logic ;
         d_arr_merge1_7_6 : IN std_logic ;
         d_arr_merge1_7_5 : IN std_logic ;
         d_arr_merge1_7_4 : IN std_logic ;
         d_arr_merge1_7_3 : IN std_logic ;
         d_arr_merge1_7_2 : IN std_logic ;
         d_arr_merge1_7_1 : IN std_logic ;
         d_arr_merge1_7_0 : IN std_logic ;
         d_arr_merge1_8_31 : IN std_logic ;
         d_arr_merge1_8_30 : IN std_logic ;
         d_arr_merge1_8_29 : IN std_logic ;
         d_arr_merge1_8_28 : IN std_logic ;
         d_arr_merge1_8_27 : IN std_logic ;
         d_arr_merge1_8_26 : IN std_logic ;
         d_arr_merge1_8_25 : IN std_logic ;
         d_arr_merge1_8_24 : IN std_logic ;
         d_arr_merge1_8_23 : IN std_logic ;
         d_arr_merge1_8_22 : IN std_logic ;
         d_arr_merge1_8_21 : IN std_logic ;
         d_arr_merge1_8_20 : IN std_logic ;
         d_arr_merge1_8_19 : IN std_logic ;
         d_arr_merge1_8_18 : IN std_logic ;
         d_arr_merge1_8_17 : IN std_logic ;
         d_arr_merge1_8_16 : IN std_logic ;
         d_arr_merge1_8_15 : IN std_logic ;
         d_arr_merge1_8_14 : IN std_logic ;
         d_arr_merge1_8_13 : IN std_logic ;
         d_arr_merge1_8_12 : IN std_logic ;
         d_arr_merge1_8_11 : IN std_logic ;
         d_arr_merge1_8_10 : IN std_logic ;
         d_arr_merge1_8_9 : IN std_logic ;
         d_arr_merge1_8_8 : IN std_logic ;
         d_arr_merge1_8_7 : IN std_logic ;
         d_arr_merge1_8_6 : IN std_logic ;
         d_arr_merge1_8_5 : IN std_logic ;
         d_arr_merge1_8_4 : IN std_logic ;
         d_arr_merge1_8_3 : IN std_logic ;
         d_arr_merge1_8_2 : IN std_logic ;
         d_arr_merge1_8_1 : IN std_logic ;
         d_arr_merge1_8_0 : IN std_logic ;
         d_arr_merge1_9_31 : IN std_logic ;
         d_arr_merge1_9_30 : IN std_logic ;
         d_arr_merge1_9_29 : IN std_logic ;
         d_arr_merge1_9_28 : IN std_logic ;
         d_arr_merge1_9_27 : IN std_logic ;
         d_arr_merge1_9_26 : IN std_logic ;
         d_arr_merge1_9_25 : IN std_logic ;
         d_arr_merge1_9_24 : IN std_logic ;
         d_arr_merge1_9_23 : IN std_logic ;
         d_arr_merge1_9_22 : IN std_logic ;
         d_arr_merge1_9_21 : IN std_logic ;
         d_arr_merge1_9_20 : IN std_logic ;
         d_arr_merge1_9_19 : IN std_logic ;
         d_arr_merge1_9_18 : IN std_logic ;
         d_arr_merge1_9_17 : IN std_logic ;
         d_arr_merge1_9_16 : IN std_logic ;
         d_arr_merge1_9_15 : IN std_logic ;
         d_arr_merge1_9_14 : IN std_logic ;
         d_arr_merge1_9_13 : IN std_logic ;
         d_arr_merge1_9_12 : IN std_logic ;
         d_arr_merge1_9_11 : IN std_logic ;
         d_arr_merge1_9_10 : IN std_logic ;
         d_arr_merge1_9_9 : IN std_logic ;
         d_arr_merge1_9_8 : IN std_logic ;
         d_arr_merge1_9_7 : IN std_logic ;
         d_arr_merge1_9_6 : IN std_logic ;
         d_arr_merge1_9_5 : IN std_logic ;
         d_arr_merge1_9_4 : IN std_logic ;
         d_arr_merge1_9_3 : IN std_logic ;
         d_arr_merge1_9_2 : IN std_logic ;
         d_arr_merge1_9_1 : IN std_logic ;
         d_arr_merge1_9_0 : IN std_logic ;
         d_arr_merge1_10_31 : IN std_logic ;
         d_arr_merge1_10_30 : IN std_logic ;
         d_arr_merge1_10_29 : IN std_logic ;
         d_arr_merge1_10_28 : IN std_logic ;
         d_arr_merge1_10_27 : IN std_logic ;
         d_arr_merge1_10_26 : IN std_logic ;
         d_arr_merge1_10_25 : IN std_logic ;
         d_arr_merge1_10_24 : IN std_logic ;
         d_arr_merge1_10_23 : IN std_logic ;
         d_arr_merge1_10_22 : IN std_logic ;
         d_arr_merge1_10_21 : IN std_logic ;
         d_arr_merge1_10_20 : IN std_logic ;
         d_arr_merge1_10_19 : IN std_logic ;
         d_arr_merge1_10_18 : IN std_logic ;
         d_arr_merge1_10_17 : IN std_logic ;
         d_arr_merge1_10_16 : IN std_logic ;
         d_arr_merge1_10_15 : IN std_logic ;
         d_arr_merge1_10_14 : IN std_logic ;
         d_arr_merge1_10_13 : IN std_logic ;
         d_arr_merge1_10_12 : IN std_logic ;
         d_arr_merge1_10_11 : IN std_logic ;
         d_arr_merge1_10_10 : IN std_logic ;
         d_arr_merge1_10_9 : IN std_logic ;
         d_arr_merge1_10_8 : IN std_logic ;
         d_arr_merge1_10_7 : IN std_logic ;
         d_arr_merge1_10_6 : IN std_logic ;
         d_arr_merge1_10_5 : IN std_logic ;
         d_arr_merge1_10_4 : IN std_logic ;
         d_arr_merge1_10_3 : IN std_logic ;
         d_arr_merge1_10_2 : IN std_logic ;
         d_arr_merge1_10_1 : IN std_logic ;
         d_arr_merge1_10_0 : IN std_logic ;
         d_arr_merge1_11_31 : IN std_logic ;
         d_arr_merge1_11_30 : IN std_logic ;
         d_arr_merge1_11_29 : IN std_logic ;
         d_arr_merge1_11_28 : IN std_logic ;
         d_arr_merge1_11_27 : IN std_logic ;
         d_arr_merge1_11_26 : IN std_logic ;
         d_arr_merge1_11_25 : IN std_logic ;
         d_arr_merge1_11_24 : IN std_logic ;
         d_arr_merge1_11_23 : IN std_logic ;
         d_arr_merge1_11_22 : IN std_logic ;
         d_arr_merge1_11_21 : IN std_logic ;
         d_arr_merge1_11_20 : IN std_logic ;
         d_arr_merge1_11_19 : IN std_logic ;
         d_arr_merge1_11_18 : IN std_logic ;
         d_arr_merge1_11_17 : IN std_logic ;
         d_arr_merge1_11_16 : IN std_logic ;
         d_arr_merge1_11_15 : IN std_logic ;
         d_arr_merge1_11_14 : IN std_logic ;
         d_arr_merge1_11_13 : IN std_logic ;
         d_arr_merge1_11_12 : IN std_logic ;
         d_arr_merge1_11_11 : IN std_logic ;
         d_arr_merge1_11_10 : IN std_logic ;
         d_arr_merge1_11_9 : IN std_logic ;
         d_arr_merge1_11_8 : IN std_logic ;
         d_arr_merge1_11_7 : IN std_logic ;
         d_arr_merge1_11_6 : IN std_logic ;
         d_arr_merge1_11_5 : IN std_logic ;
         d_arr_merge1_11_4 : IN std_logic ;
         d_arr_merge1_11_3 : IN std_logic ;
         d_arr_merge1_11_2 : IN std_logic ;
         d_arr_merge1_11_1 : IN std_logic ;
         d_arr_merge1_11_0 : IN std_logic ;
         d_arr_merge1_12_31 : IN std_logic ;
         d_arr_merge1_12_30 : IN std_logic ;
         d_arr_merge1_12_29 : IN std_logic ;
         d_arr_merge1_12_28 : IN std_logic ;
         d_arr_merge1_12_27 : IN std_logic ;
         d_arr_merge1_12_26 : IN std_logic ;
         d_arr_merge1_12_25 : IN std_logic ;
         d_arr_merge1_12_24 : IN std_logic ;
         d_arr_merge1_12_23 : IN std_logic ;
         d_arr_merge1_12_22 : IN std_logic ;
         d_arr_merge1_12_21 : IN std_logic ;
         d_arr_merge1_12_20 : IN std_logic ;
         d_arr_merge1_12_19 : IN std_logic ;
         d_arr_merge1_12_18 : IN std_logic ;
         d_arr_merge1_12_17 : IN std_logic ;
         d_arr_merge1_12_16 : IN std_logic ;
         d_arr_merge1_12_15 : IN std_logic ;
         d_arr_merge1_12_14 : IN std_logic ;
         d_arr_merge1_12_13 : IN std_logic ;
         d_arr_merge1_12_12 : IN std_logic ;
         d_arr_merge1_12_11 : IN std_logic ;
         d_arr_merge1_12_10 : IN std_logic ;
         d_arr_merge1_12_9 : IN std_logic ;
         d_arr_merge1_12_8 : IN std_logic ;
         d_arr_merge1_12_7 : IN std_logic ;
         d_arr_merge1_12_6 : IN std_logic ;
         d_arr_merge1_12_5 : IN std_logic ;
         d_arr_merge1_12_4 : IN std_logic ;
         d_arr_merge1_12_3 : IN std_logic ;
         d_arr_merge1_12_2 : IN std_logic ;
         d_arr_merge1_12_1 : IN std_logic ;
         d_arr_merge1_12_0 : IN std_logic ;
         d_arr_merge1_13_31 : IN std_logic ;
         d_arr_merge1_13_30 : IN std_logic ;
         d_arr_merge1_13_29 : IN std_logic ;
         d_arr_merge1_13_28 : IN std_logic ;
         d_arr_merge1_13_27 : IN std_logic ;
         d_arr_merge1_13_26 : IN std_logic ;
         d_arr_merge1_13_25 : IN std_logic ;
         d_arr_merge1_13_24 : IN std_logic ;
         d_arr_merge1_13_23 : IN std_logic ;
         d_arr_merge1_13_22 : IN std_logic ;
         d_arr_merge1_13_21 : IN std_logic ;
         d_arr_merge1_13_20 : IN std_logic ;
         d_arr_merge1_13_19 : IN std_logic ;
         d_arr_merge1_13_18 : IN std_logic ;
         d_arr_merge1_13_17 : IN std_logic ;
         d_arr_merge1_13_16 : IN std_logic ;
         d_arr_merge1_13_15 : IN std_logic ;
         d_arr_merge1_13_14 : IN std_logic ;
         d_arr_merge1_13_13 : IN std_logic ;
         d_arr_merge1_13_12 : IN std_logic ;
         d_arr_merge1_13_11 : IN std_logic ;
         d_arr_merge1_13_10 : IN std_logic ;
         d_arr_merge1_13_9 : IN std_logic ;
         d_arr_merge1_13_8 : IN std_logic ;
         d_arr_merge1_13_7 : IN std_logic ;
         d_arr_merge1_13_6 : IN std_logic ;
         d_arr_merge1_13_5 : IN std_logic ;
         d_arr_merge1_13_4 : IN std_logic ;
         d_arr_merge1_13_3 : IN std_logic ;
         d_arr_merge1_13_2 : IN std_logic ;
         d_arr_merge1_13_1 : IN std_logic ;
         d_arr_merge1_13_0 : IN std_logic ;
         d_arr_merge1_14_31 : IN std_logic ;
         d_arr_merge1_14_30 : IN std_logic ;
         d_arr_merge1_14_29 : IN std_logic ;
         d_arr_merge1_14_28 : IN std_logic ;
         d_arr_merge1_14_27 : IN std_logic ;
         d_arr_merge1_14_26 : IN std_logic ;
         d_arr_merge1_14_25 : IN std_logic ;
         d_arr_merge1_14_24 : IN std_logic ;
         d_arr_merge1_14_23 : IN std_logic ;
         d_arr_merge1_14_22 : IN std_logic ;
         d_arr_merge1_14_21 : IN std_logic ;
         d_arr_merge1_14_20 : IN std_logic ;
         d_arr_merge1_14_19 : IN std_logic ;
         d_arr_merge1_14_18 : IN std_logic ;
         d_arr_merge1_14_17 : IN std_logic ;
         d_arr_merge1_14_16 : IN std_logic ;
         d_arr_merge1_14_15 : IN std_logic ;
         d_arr_merge1_14_14 : IN std_logic ;
         d_arr_merge1_14_13 : IN std_logic ;
         d_arr_merge1_14_12 : IN std_logic ;
         d_arr_merge1_14_11 : IN std_logic ;
         d_arr_merge1_14_10 : IN std_logic ;
         d_arr_merge1_14_9 : IN std_logic ;
         d_arr_merge1_14_8 : IN std_logic ;
         d_arr_merge1_14_7 : IN std_logic ;
         d_arr_merge1_14_6 : IN std_logic ;
         d_arr_merge1_14_5 : IN std_logic ;
         d_arr_merge1_14_4 : IN std_logic ;
         d_arr_merge1_14_3 : IN std_logic ;
         d_arr_merge1_14_2 : IN std_logic ;
         d_arr_merge1_14_1 : IN std_logic ;
         d_arr_merge1_14_0 : IN std_logic ;
         d_arr_merge1_15_31 : IN std_logic ;
         d_arr_merge1_15_30 : IN std_logic ;
         d_arr_merge1_15_29 : IN std_logic ;
         d_arr_merge1_15_28 : IN std_logic ;
         d_arr_merge1_15_27 : IN std_logic ;
         d_arr_merge1_15_26 : IN std_logic ;
         d_arr_merge1_15_25 : IN std_logic ;
         d_arr_merge1_15_24 : IN std_logic ;
         d_arr_merge1_15_23 : IN std_logic ;
         d_arr_merge1_15_22 : IN std_logic ;
         d_arr_merge1_15_21 : IN std_logic ;
         d_arr_merge1_15_20 : IN std_logic ;
         d_arr_merge1_15_19 : IN std_logic ;
         d_arr_merge1_15_18 : IN std_logic ;
         d_arr_merge1_15_17 : IN std_logic ;
         d_arr_merge1_15_16 : IN std_logic ;
         d_arr_merge1_15_15 : IN std_logic ;
         d_arr_merge1_15_14 : IN std_logic ;
         d_arr_merge1_15_13 : IN std_logic ;
         d_arr_merge1_15_12 : IN std_logic ;
         d_arr_merge1_15_11 : IN std_logic ;
         d_arr_merge1_15_10 : IN std_logic ;
         d_arr_merge1_15_9 : IN std_logic ;
         d_arr_merge1_15_8 : IN std_logic ;
         d_arr_merge1_15_7 : IN std_logic ;
         d_arr_merge1_15_6 : IN std_logic ;
         d_arr_merge1_15_5 : IN std_logic ;
         d_arr_merge1_15_4 : IN std_logic ;
         d_arr_merge1_15_3 : IN std_logic ;
         d_arr_merge1_15_2 : IN std_logic ;
         d_arr_merge1_15_1 : IN std_logic ;
         d_arr_merge1_15_0 : IN std_logic ;
         d_arr_merge1_16_31 : IN std_logic ;
         d_arr_merge1_16_30 : IN std_logic ;
         d_arr_merge1_16_29 : IN std_logic ;
         d_arr_merge1_16_28 : IN std_logic ;
         d_arr_merge1_16_27 : IN std_logic ;
         d_arr_merge1_16_26 : IN std_logic ;
         d_arr_merge1_16_25 : IN std_logic ;
         d_arr_merge1_16_24 : IN std_logic ;
         d_arr_merge1_16_23 : IN std_logic ;
         d_arr_merge1_16_22 : IN std_logic ;
         d_arr_merge1_16_21 : IN std_logic ;
         d_arr_merge1_16_20 : IN std_logic ;
         d_arr_merge1_16_19 : IN std_logic ;
         d_arr_merge1_16_18 : IN std_logic ;
         d_arr_merge1_16_17 : IN std_logic ;
         d_arr_merge1_16_16 : IN std_logic ;
         d_arr_merge1_16_15 : IN std_logic ;
         d_arr_merge1_16_14 : IN std_logic ;
         d_arr_merge1_16_13 : IN std_logic ;
         d_arr_merge1_16_12 : IN std_logic ;
         d_arr_merge1_16_11 : IN std_logic ;
         d_arr_merge1_16_10 : IN std_logic ;
         d_arr_merge1_16_9 : IN std_logic ;
         d_arr_merge1_16_8 : IN std_logic ;
         d_arr_merge1_16_7 : IN std_logic ;
         d_arr_merge1_16_6 : IN std_logic ;
         d_arr_merge1_16_5 : IN std_logic ;
         d_arr_merge1_16_4 : IN std_logic ;
         d_arr_merge1_16_3 : IN std_logic ;
         d_arr_merge1_16_2 : IN std_logic ;
         d_arr_merge1_16_1 : IN std_logic ;
         d_arr_merge1_16_0 : IN std_logic ;
         d_arr_merge1_17_31 : IN std_logic ;
         d_arr_merge1_17_30 : IN std_logic ;
         d_arr_merge1_17_29 : IN std_logic ;
         d_arr_merge1_17_28 : IN std_logic ;
         d_arr_merge1_17_27 : IN std_logic ;
         d_arr_merge1_17_26 : IN std_logic ;
         d_arr_merge1_17_25 : IN std_logic ;
         d_arr_merge1_17_24 : IN std_logic ;
         d_arr_merge1_17_23 : IN std_logic ;
         d_arr_merge1_17_22 : IN std_logic ;
         d_arr_merge1_17_21 : IN std_logic ;
         d_arr_merge1_17_20 : IN std_logic ;
         d_arr_merge1_17_19 : IN std_logic ;
         d_arr_merge1_17_18 : IN std_logic ;
         d_arr_merge1_17_17 : IN std_logic ;
         d_arr_merge1_17_16 : IN std_logic ;
         d_arr_merge1_17_15 : IN std_logic ;
         d_arr_merge1_17_14 : IN std_logic ;
         d_arr_merge1_17_13 : IN std_logic ;
         d_arr_merge1_17_12 : IN std_logic ;
         d_arr_merge1_17_11 : IN std_logic ;
         d_arr_merge1_17_10 : IN std_logic ;
         d_arr_merge1_17_9 : IN std_logic ;
         d_arr_merge1_17_8 : IN std_logic ;
         d_arr_merge1_17_7 : IN std_logic ;
         d_arr_merge1_17_6 : IN std_logic ;
         d_arr_merge1_17_5 : IN std_logic ;
         d_arr_merge1_17_4 : IN std_logic ;
         d_arr_merge1_17_3 : IN std_logic ;
         d_arr_merge1_17_2 : IN std_logic ;
         d_arr_merge1_17_1 : IN std_logic ;
         d_arr_merge1_17_0 : IN std_logic ;
         d_arr_merge1_18_31 : IN std_logic ;
         d_arr_merge1_18_30 : IN std_logic ;
         d_arr_merge1_18_29 : IN std_logic ;
         d_arr_merge1_18_28 : IN std_logic ;
         d_arr_merge1_18_27 : IN std_logic ;
         d_arr_merge1_18_26 : IN std_logic ;
         d_arr_merge1_18_25 : IN std_logic ;
         d_arr_merge1_18_24 : IN std_logic ;
         d_arr_merge1_18_23 : IN std_logic ;
         d_arr_merge1_18_22 : IN std_logic ;
         d_arr_merge1_18_21 : IN std_logic ;
         d_arr_merge1_18_20 : IN std_logic ;
         d_arr_merge1_18_19 : IN std_logic ;
         d_arr_merge1_18_18 : IN std_logic ;
         d_arr_merge1_18_17 : IN std_logic ;
         d_arr_merge1_18_16 : IN std_logic ;
         d_arr_merge1_18_15 : IN std_logic ;
         d_arr_merge1_18_14 : IN std_logic ;
         d_arr_merge1_18_13 : IN std_logic ;
         d_arr_merge1_18_12 : IN std_logic ;
         d_arr_merge1_18_11 : IN std_logic ;
         d_arr_merge1_18_10 : IN std_logic ;
         d_arr_merge1_18_9 : IN std_logic ;
         d_arr_merge1_18_8 : IN std_logic ;
         d_arr_merge1_18_7 : IN std_logic ;
         d_arr_merge1_18_6 : IN std_logic ;
         d_arr_merge1_18_5 : IN std_logic ;
         d_arr_merge1_18_4 : IN std_logic ;
         d_arr_merge1_18_3 : IN std_logic ;
         d_arr_merge1_18_2 : IN std_logic ;
         d_arr_merge1_18_1 : IN std_logic ;
         d_arr_merge1_18_0 : IN std_logic ;
         d_arr_merge1_19_31 : IN std_logic ;
         d_arr_merge1_19_30 : IN std_logic ;
         d_arr_merge1_19_29 : IN std_logic ;
         d_arr_merge1_19_28 : IN std_logic ;
         d_arr_merge1_19_27 : IN std_logic ;
         d_arr_merge1_19_26 : IN std_logic ;
         d_arr_merge1_19_25 : IN std_logic ;
         d_arr_merge1_19_24 : IN std_logic ;
         d_arr_merge1_19_23 : IN std_logic ;
         d_arr_merge1_19_22 : IN std_logic ;
         d_arr_merge1_19_21 : IN std_logic ;
         d_arr_merge1_19_20 : IN std_logic ;
         d_arr_merge1_19_19 : IN std_logic ;
         d_arr_merge1_19_18 : IN std_logic ;
         d_arr_merge1_19_17 : IN std_logic ;
         d_arr_merge1_19_16 : IN std_logic ;
         d_arr_merge1_19_15 : IN std_logic ;
         d_arr_merge1_19_14 : IN std_logic ;
         d_arr_merge1_19_13 : IN std_logic ;
         d_arr_merge1_19_12 : IN std_logic ;
         d_arr_merge1_19_11 : IN std_logic ;
         d_arr_merge1_19_10 : IN std_logic ;
         d_arr_merge1_19_9 : IN std_logic ;
         d_arr_merge1_19_8 : IN std_logic ;
         d_arr_merge1_19_7 : IN std_logic ;
         d_arr_merge1_19_6 : IN std_logic ;
         d_arr_merge1_19_5 : IN std_logic ;
         d_arr_merge1_19_4 : IN std_logic ;
         d_arr_merge1_19_3 : IN std_logic ;
         d_arr_merge1_19_2 : IN std_logic ;
         d_arr_merge1_19_1 : IN std_logic ;
         d_arr_merge1_19_0 : IN std_logic ;
         d_arr_merge1_20_31 : IN std_logic ;
         d_arr_merge1_20_30 : IN std_logic ;
         d_arr_merge1_20_29 : IN std_logic ;
         d_arr_merge1_20_28 : IN std_logic ;
         d_arr_merge1_20_27 : IN std_logic ;
         d_arr_merge1_20_26 : IN std_logic ;
         d_arr_merge1_20_25 : IN std_logic ;
         d_arr_merge1_20_24 : IN std_logic ;
         d_arr_merge1_20_23 : IN std_logic ;
         d_arr_merge1_20_22 : IN std_logic ;
         d_arr_merge1_20_21 : IN std_logic ;
         d_arr_merge1_20_20 : IN std_logic ;
         d_arr_merge1_20_19 : IN std_logic ;
         d_arr_merge1_20_18 : IN std_logic ;
         d_arr_merge1_20_17 : IN std_logic ;
         d_arr_merge1_20_16 : IN std_logic ;
         d_arr_merge1_20_15 : IN std_logic ;
         d_arr_merge1_20_14 : IN std_logic ;
         d_arr_merge1_20_13 : IN std_logic ;
         d_arr_merge1_20_12 : IN std_logic ;
         d_arr_merge1_20_11 : IN std_logic ;
         d_arr_merge1_20_10 : IN std_logic ;
         d_arr_merge1_20_9 : IN std_logic ;
         d_arr_merge1_20_8 : IN std_logic ;
         d_arr_merge1_20_7 : IN std_logic ;
         d_arr_merge1_20_6 : IN std_logic ;
         d_arr_merge1_20_5 : IN std_logic ;
         d_arr_merge1_20_4 : IN std_logic ;
         d_arr_merge1_20_3 : IN std_logic ;
         d_arr_merge1_20_2 : IN std_logic ;
         d_arr_merge1_20_1 : IN std_logic ;
         d_arr_merge1_20_0 : IN std_logic ;
         d_arr_merge1_21_31 : IN std_logic ;
         d_arr_merge1_21_30 : IN std_logic ;
         d_arr_merge1_21_29 : IN std_logic ;
         d_arr_merge1_21_28 : IN std_logic ;
         d_arr_merge1_21_27 : IN std_logic ;
         d_arr_merge1_21_26 : IN std_logic ;
         d_arr_merge1_21_25 : IN std_logic ;
         d_arr_merge1_21_24 : IN std_logic ;
         d_arr_merge1_21_23 : IN std_logic ;
         d_arr_merge1_21_22 : IN std_logic ;
         d_arr_merge1_21_21 : IN std_logic ;
         d_arr_merge1_21_20 : IN std_logic ;
         d_arr_merge1_21_19 : IN std_logic ;
         d_arr_merge1_21_18 : IN std_logic ;
         d_arr_merge1_21_17 : IN std_logic ;
         d_arr_merge1_21_16 : IN std_logic ;
         d_arr_merge1_21_15 : IN std_logic ;
         d_arr_merge1_21_14 : IN std_logic ;
         d_arr_merge1_21_13 : IN std_logic ;
         d_arr_merge1_21_12 : IN std_logic ;
         d_arr_merge1_21_11 : IN std_logic ;
         d_arr_merge1_21_10 : IN std_logic ;
         d_arr_merge1_21_9 : IN std_logic ;
         d_arr_merge1_21_8 : IN std_logic ;
         d_arr_merge1_21_7 : IN std_logic ;
         d_arr_merge1_21_6 : IN std_logic ;
         d_arr_merge1_21_5 : IN std_logic ;
         d_arr_merge1_21_4 : IN std_logic ;
         d_arr_merge1_21_3 : IN std_logic ;
         d_arr_merge1_21_2 : IN std_logic ;
         d_arr_merge1_21_1 : IN std_logic ;
         d_arr_merge1_21_0 : IN std_logic ;
         d_arr_merge1_22_31 : IN std_logic ;
         d_arr_merge1_22_30 : IN std_logic ;
         d_arr_merge1_22_29 : IN std_logic ;
         d_arr_merge1_22_28 : IN std_logic ;
         d_arr_merge1_22_27 : IN std_logic ;
         d_arr_merge1_22_26 : IN std_logic ;
         d_arr_merge1_22_25 : IN std_logic ;
         d_arr_merge1_22_24 : IN std_logic ;
         d_arr_merge1_22_23 : IN std_logic ;
         d_arr_merge1_22_22 : IN std_logic ;
         d_arr_merge1_22_21 : IN std_logic ;
         d_arr_merge1_22_20 : IN std_logic ;
         d_arr_merge1_22_19 : IN std_logic ;
         d_arr_merge1_22_18 : IN std_logic ;
         d_arr_merge1_22_17 : IN std_logic ;
         d_arr_merge1_22_16 : IN std_logic ;
         d_arr_merge1_22_15 : IN std_logic ;
         d_arr_merge1_22_14 : IN std_logic ;
         d_arr_merge1_22_13 : IN std_logic ;
         d_arr_merge1_22_12 : IN std_logic ;
         d_arr_merge1_22_11 : IN std_logic ;
         d_arr_merge1_22_10 : IN std_logic ;
         d_arr_merge1_22_9 : IN std_logic ;
         d_arr_merge1_22_8 : IN std_logic ;
         d_arr_merge1_22_7 : IN std_logic ;
         d_arr_merge1_22_6 : IN std_logic ;
         d_arr_merge1_22_5 : IN std_logic ;
         d_arr_merge1_22_4 : IN std_logic ;
         d_arr_merge1_22_3 : IN std_logic ;
         d_arr_merge1_22_2 : IN std_logic ;
         d_arr_merge1_22_1 : IN std_logic ;
         d_arr_merge1_22_0 : IN std_logic ;
         d_arr_merge1_23_31 : IN std_logic ;
         d_arr_merge1_23_30 : IN std_logic ;
         d_arr_merge1_23_29 : IN std_logic ;
         d_arr_merge1_23_28 : IN std_logic ;
         d_arr_merge1_23_27 : IN std_logic ;
         d_arr_merge1_23_26 : IN std_logic ;
         d_arr_merge1_23_25 : IN std_logic ;
         d_arr_merge1_23_24 : IN std_logic ;
         d_arr_merge1_23_23 : IN std_logic ;
         d_arr_merge1_23_22 : IN std_logic ;
         d_arr_merge1_23_21 : IN std_logic ;
         d_arr_merge1_23_20 : IN std_logic ;
         d_arr_merge1_23_19 : IN std_logic ;
         d_arr_merge1_23_18 : IN std_logic ;
         d_arr_merge1_23_17 : IN std_logic ;
         d_arr_merge1_23_16 : IN std_logic ;
         d_arr_merge1_23_15 : IN std_logic ;
         d_arr_merge1_23_14 : IN std_logic ;
         d_arr_merge1_23_13 : IN std_logic ;
         d_arr_merge1_23_12 : IN std_logic ;
         d_arr_merge1_23_11 : IN std_logic ;
         d_arr_merge1_23_10 : IN std_logic ;
         d_arr_merge1_23_9 : IN std_logic ;
         d_arr_merge1_23_8 : IN std_logic ;
         d_arr_merge1_23_7 : IN std_logic ;
         d_arr_merge1_23_6 : IN std_logic ;
         d_arr_merge1_23_5 : IN std_logic ;
         d_arr_merge1_23_4 : IN std_logic ;
         d_arr_merge1_23_3 : IN std_logic ;
         d_arr_merge1_23_2 : IN std_logic ;
         d_arr_merge1_23_1 : IN std_logic ;
         d_arr_merge1_23_0 : IN std_logic ;
         d_arr_merge1_24_31 : IN std_logic ;
         d_arr_merge1_24_30 : IN std_logic ;
         d_arr_merge1_24_29 : IN std_logic ;
         d_arr_merge1_24_28 : IN std_logic ;
         d_arr_merge1_24_27 : IN std_logic ;
         d_arr_merge1_24_26 : IN std_logic ;
         d_arr_merge1_24_25 : IN std_logic ;
         d_arr_merge1_24_24 : IN std_logic ;
         d_arr_merge1_24_23 : IN std_logic ;
         d_arr_merge1_24_22 : IN std_logic ;
         d_arr_merge1_24_21 : IN std_logic ;
         d_arr_merge1_24_20 : IN std_logic ;
         d_arr_merge1_24_19 : IN std_logic ;
         d_arr_merge1_24_18 : IN std_logic ;
         d_arr_merge1_24_17 : IN std_logic ;
         d_arr_merge1_24_16 : IN std_logic ;
         d_arr_merge1_24_15 : IN std_logic ;
         d_arr_merge1_24_14 : IN std_logic ;
         d_arr_merge1_24_13 : IN std_logic ;
         d_arr_merge1_24_12 : IN std_logic ;
         d_arr_merge1_24_11 : IN std_logic ;
         d_arr_merge1_24_10 : IN std_logic ;
         d_arr_merge1_24_9 : IN std_logic ;
         d_arr_merge1_24_8 : IN std_logic ;
         d_arr_merge1_24_7 : IN std_logic ;
         d_arr_merge1_24_6 : IN std_logic ;
         d_arr_merge1_24_5 : IN std_logic ;
         d_arr_merge1_24_4 : IN std_logic ;
         d_arr_merge1_24_3 : IN std_logic ;
         d_arr_merge1_24_2 : IN std_logic ;
         d_arr_merge1_24_1 : IN std_logic ;
         d_arr_merge1_24_0 : IN std_logic ;
         d_arr_merge2_0_31 : IN std_logic ;
         d_arr_merge2_0_30 : IN std_logic ;
         d_arr_merge2_0_29 : IN std_logic ;
         d_arr_merge2_0_28 : IN std_logic ;
         d_arr_merge2_0_27 : IN std_logic ;
         d_arr_merge2_0_26 : IN std_logic ;
         d_arr_merge2_0_25 : IN std_logic ;
         d_arr_merge2_0_24 : IN std_logic ;
         d_arr_merge2_0_23 : IN std_logic ;
         d_arr_merge2_0_22 : IN std_logic ;
         d_arr_merge2_0_21 : IN std_logic ;
         d_arr_merge2_0_20 : IN std_logic ;
         d_arr_merge2_0_19 : IN std_logic ;
         d_arr_merge2_0_18 : IN std_logic ;
         d_arr_merge2_0_17 : IN std_logic ;
         d_arr_merge2_0_16 : IN std_logic ;
         d_arr_merge2_0_15 : IN std_logic ;
         d_arr_merge2_0_14 : IN std_logic ;
         d_arr_merge2_0_13 : IN std_logic ;
         d_arr_merge2_0_12 : IN std_logic ;
         d_arr_merge2_0_11 : IN std_logic ;
         d_arr_merge2_0_10 : IN std_logic ;
         d_arr_merge2_0_9 : IN std_logic ;
         d_arr_merge2_0_8 : IN std_logic ;
         d_arr_merge2_0_7 : IN std_logic ;
         d_arr_merge2_0_6 : IN std_logic ;
         d_arr_merge2_0_5 : IN std_logic ;
         d_arr_merge2_0_4 : IN std_logic ;
         d_arr_merge2_0_3 : IN std_logic ;
         d_arr_merge2_0_2 : IN std_logic ;
         d_arr_merge2_0_1 : IN std_logic ;
         d_arr_merge2_0_0 : IN std_logic ;
         d_arr_merge2_1_31 : IN std_logic ;
         d_arr_merge2_1_30 : IN std_logic ;
         d_arr_merge2_1_29 : IN std_logic ;
         d_arr_merge2_1_28 : IN std_logic ;
         d_arr_merge2_1_27 : IN std_logic ;
         d_arr_merge2_1_26 : IN std_logic ;
         d_arr_merge2_1_25 : IN std_logic ;
         d_arr_merge2_1_24 : IN std_logic ;
         d_arr_merge2_1_23 : IN std_logic ;
         d_arr_merge2_1_22 : IN std_logic ;
         d_arr_merge2_1_21 : IN std_logic ;
         d_arr_merge2_1_20 : IN std_logic ;
         d_arr_merge2_1_19 : IN std_logic ;
         d_arr_merge2_1_18 : IN std_logic ;
         d_arr_merge2_1_17 : IN std_logic ;
         d_arr_merge2_1_16 : IN std_logic ;
         d_arr_merge2_1_15 : IN std_logic ;
         d_arr_merge2_1_14 : IN std_logic ;
         d_arr_merge2_1_13 : IN std_logic ;
         d_arr_merge2_1_12 : IN std_logic ;
         d_arr_merge2_1_11 : IN std_logic ;
         d_arr_merge2_1_10 : IN std_logic ;
         d_arr_merge2_1_9 : IN std_logic ;
         d_arr_merge2_1_8 : IN std_logic ;
         d_arr_merge2_1_7 : IN std_logic ;
         d_arr_merge2_1_6 : IN std_logic ;
         d_arr_merge2_1_5 : IN std_logic ;
         d_arr_merge2_1_4 : IN std_logic ;
         d_arr_merge2_1_3 : IN std_logic ;
         d_arr_merge2_1_2 : IN std_logic ;
         d_arr_merge2_1_1 : IN std_logic ;
         d_arr_merge2_1_0 : IN std_logic ;
         d_arr_merge2_2_31 : IN std_logic ;
         d_arr_merge2_2_30 : IN std_logic ;
         d_arr_merge2_2_29 : IN std_logic ;
         d_arr_merge2_2_28 : IN std_logic ;
         d_arr_merge2_2_27 : IN std_logic ;
         d_arr_merge2_2_26 : IN std_logic ;
         d_arr_merge2_2_25 : IN std_logic ;
         d_arr_merge2_2_24 : IN std_logic ;
         d_arr_merge2_2_23 : IN std_logic ;
         d_arr_merge2_2_22 : IN std_logic ;
         d_arr_merge2_2_21 : IN std_logic ;
         d_arr_merge2_2_20 : IN std_logic ;
         d_arr_merge2_2_19 : IN std_logic ;
         d_arr_merge2_2_18 : IN std_logic ;
         d_arr_merge2_2_17 : IN std_logic ;
         d_arr_merge2_2_16 : IN std_logic ;
         d_arr_merge2_2_15 : IN std_logic ;
         d_arr_merge2_2_14 : IN std_logic ;
         d_arr_merge2_2_13 : IN std_logic ;
         d_arr_merge2_2_12 : IN std_logic ;
         d_arr_merge2_2_11 : IN std_logic ;
         d_arr_merge2_2_10 : IN std_logic ;
         d_arr_merge2_2_9 : IN std_logic ;
         d_arr_merge2_2_8 : IN std_logic ;
         d_arr_merge2_2_7 : IN std_logic ;
         d_arr_merge2_2_6 : IN std_logic ;
         d_arr_merge2_2_5 : IN std_logic ;
         d_arr_merge2_2_4 : IN std_logic ;
         d_arr_merge2_2_3 : IN std_logic ;
         d_arr_merge2_2_2 : IN std_logic ;
         d_arr_merge2_2_1 : IN std_logic ;
         d_arr_merge2_2_0 : IN std_logic ;
         d_arr_merge2_3_31 : IN std_logic ;
         d_arr_merge2_3_30 : IN std_logic ;
         d_arr_merge2_3_29 : IN std_logic ;
         d_arr_merge2_3_28 : IN std_logic ;
         d_arr_merge2_3_27 : IN std_logic ;
         d_arr_merge2_3_26 : IN std_logic ;
         d_arr_merge2_3_25 : IN std_logic ;
         d_arr_merge2_3_24 : IN std_logic ;
         d_arr_merge2_3_23 : IN std_logic ;
         d_arr_merge2_3_22 : IN std_logic ;
         d_arr_merge2_3_21 : IN std_logic ;
         d_arr_merge2_3_20 : IN std_logic ;
         d_arr_merge2_3_19 : IN std_logic ;
         d_arr_merge2_3_18 : IN std_logic ;
         d_arr_merge2_3_17 : IN std_logic ;
         d_arr_merge2_3_16 : IN std_logic ;
         d_arr_merge2_3_15 : IN std_logic ;
         d_arr_merge2_3_14 : IN std_logic ;
         d_arr_merge2_3_13 : IN std_logic ;
         d_arr_merge2_3_12 : IN std_logic ;
         d_arr_merge2_3_11 : IN std_logic ;
         d_arr_merge2_3_10 : IN std_logic ;
         d_arr_merge2_3_9 : IN std_logic ;
         d_arr_merge2_3_8 : IN std_logic ;
         d_arr_merge2_3_7 : IN std_logic ;
         d_arr_merge2_3_6 : IN std_logic ;
         d_arr_merge2_3_5 : IN std_logic ;
         d_arr_merge2_3_4 : IN std_logic ;
         d_arr_merge2_3_3 : IN std_logic ;
         d_arr_merge2_3_2 : IN std_logic ;
         d_arr_merge2_3_1 : IN std_logic ;
         d_arr_merge2_3_0 : IN std_logic ;
         d_arr_merge2_4_31 : IN std_logic ;
         d_arr_merge2_4_30 : IN std_logic ;
         d_arr_merge2_4_29 : IN std_logic ;
         d_arr_merge2_4_28 : IN std_logic ;
         d_arr_merge2_4_27 : IN std_logic ;
         d_arr_merge2_4_26 : IN std_logic ;
         d_arr_merge2_4_25 : IN std_logic ;
         d_arr_merge2_4_24 : IN std_logic ;
         d_arr_merge2_4_23 : IN std_logic ;
         d_arr_merge2_4_22 : IN std_logic ;
         d_arr_merge2_4_21 : IN std_logic ;
         d_arr_merge2_4_20 : IN std_logic ;
         d_arr_merge2_4_19 : IN std_logic ;
         d_arr_merge2_4_18 : IN std_logic ;
         d_arr_merge2_4_17 : IN std_logic ;
         d_arr_merge2_4_16 : IN std_logic ;
         d_arr_merge2_4_15 : IN std_logic ;
         d_arr_merge2_4_14 : IN std_logic ;
         d_arr_merge2_4_13 : IN std_logic ;
         d_arr_merge2_4_12 : IN std_logic ;
         d_arr_merge2_4_11 : IN std_logic ;
         d_arr_merge2_4_10 : IN std_logic ;
         d_arr_merge2_4_9 : IN std_logic ;
         d_arr_merge2_4_8 : IN std_logic ;
         d_arr_merge2_4_7 : IN std_logic ;
         d_arr_merge2_4_6 : IN std_logic ;
         d_arr_merge2_4_5 : IN std_logic ;
         d_arr_merge2_4_4 : IN std_logic ;
         d_arr_merge2_4_3 : IN std_logic ;
         d_arr_merge2_4_2 : IN std_logic ;
         d_arr_merge2_4_1 : IN std_logic ;
         d_arr_merge2_4_0 : IN std_logic ;
         d_arr_merge2_5_31 : IN std_logic ;
         d_arr_merge2_5_30 : IN std_logic ;
         d_arr_merge2_5_29 : IN std_logic ;
         d_arr_merge2_5_28 : IN std_logic ;
         d_arr_merge2_5_27 : IN std_logic ;
         d_arr_merge2_5_26 : IN std_logic ;
         d_arr_merge2_5_25 : IN std_logic ;
         d_arr_merge2_5_24 : IN std_logic ;
         d_arr_merge2_5_23 : IN std_logic ;
         d_arr_merge2_5_22 : IN std_logic ;
         d_arr_merge2_5_21 : IN std_logic ;
         d_arr_merge2_5_20 : IN std_logic ;
         d_arr_merge2_5_19 : IN std_logic ;
         d_arr_merge2_5_18 : IN std_logic ;
         d_arr_merge2_5_17 : IN std_logic ;
         d_arr_merge2_5_16 : IN std_logic ;
         d_arr_merge2_5_15 : IN std_logic ;
         d_arr_merge2_5_14 : IN std_logic ;
         d_arr_merge2_5_13 : IN std_logic ;
         d_arr_merge2_5_12 : IN std_logic ;
         d_arr_merge2_5_11 : IN std_logic ;
         d_arr_merge2_5_10 : IN std_logic ;
         d_arr_merge2_5_9 : IN std_logic ;
         d_arr_merge2_5_8 : IN std_logic ;
         d_arr_merge2_5_7 : IN std_logic ;
         d_arr_merge2_5_6 : IN std_logic ;
         d_arr_merge2_5_5 : IN std_logic ;
         d_arr_merge2_5_4 : IN std_logic ;
         d_arr_merge2_5_3 : IN std_logic ;
         d_arr_merge2_5_2 : IN std_logic ;
         d_arr_merge2_5_1 : IN std_logic ;
         d_arr_merge2_5_0 : IN std_logic ;
         d_arr_merge2_6_31 : IN std_logic ;
         d_arr_merge2_6_30 : IN std_logic ;
         d_arr_merge2_6_29 : IN std_logic ;
         d_arr_merge2_6_28 : IN std_logic ;
         d_arr_merge2_6_27 : IN std_logic ;
         d_arr_merge2_6_26 : IN std_logic ;
         d_arr_merge2_6_25 : IN std_logic ;
         d_arr_merge2_6_24 : IN std_logic ;
         d_arr_merge2_6_23 : IN std_logic ;
         d_arr_merge2_6_22 : IN std_logic ;
         d_arr_merge2_6_21 : IN std_logic ;
         d_arr_merge2_6_20 : IN std_logic ;
         d_arr_merge2_6_19 : IN std_logic ;
         d_arr_merge2_6_18 : IN std_logic ;
         d_arr_merge2_6_17 : IN std_logic ;
         d_arr_merge2_6_16 : IN std_logic ;
         d_arr_merge2_6_15 : IN std_logic ;
         d_arr_merge2_6_14 : IN std_logic ;
         d_arr_merge2_6_13 : IN std_logic ;
         d_arr_merge2_6_12 : IN std_logic ;
         d_arr_merge2_6_11 : IN std_logic ;
         d_arr_merge2_6_10 : IN std_logic ;
         d_arr_merge2_6_9 : IN std_logic ;
         d_arr_merge2_6_8 : IN std_logic ;
         d_arr_merge2_6_7 : IN std_logic ;
         d_arr_merge2_6_6 : IN std_logic ;
         d_arr_merge2_6_5 : IN std_logic ;
         d_arr_merge2_6_4 : IN std_logic ;
         d_arr_merge2_6_3 : IN std_logic ;
         d_arr_merge2_6_2 : IN std_logic ;
         d_arr_merge2_6_1 : IN std_logic ;
         d_arr_merge2_6_0 : IN std_logic ;
         d_arr_merge2_7_31 : IN std_logic ;
         d_arr_merge2_7_30 : IN std_logic ;
         d_arr_merge2_7_29 : IN std_logic ;
         d_arr_merge2_7_28 : IN std_logic ;
         d_arr_merge2_7_27 : IN std_logic ;
         d_arr_merge2_7_26 : IN std_logic ;
         d_arr_merge2_7_25 : IN std_logic ;
         d_arr_merge2_7_24 : IN std_logic ;
         d_arr_merge2_7_23 : IN std_logic ;
         d_arr_merge2_7_22 : IN std_logic ;
         d_arr_merge2_7_21 : IN std_logic ;
         d_arr_merge2_7_20 : IN std_logic ;
         d_arr_merge2_7_19 : IN std_logic ;
         d_arr_merge2_7_18 : IN std_logic ;
         d_arr_merge2_7_17 : IN std_logic ;
         d_arr_merge2_7_16 : IN std_logic ;
         d_arr_merge2_7_15 : IN std_logic ;
         d_arr_merge2_7_14 : IN std_logic ;
         d_arr_merge2_7_13 : IN std_logic ;
         d_arr_merge2_7_12 : IN std_logic ;
         d_arr_merge2_7_11 : IN std_logic ;
         d_arr_merge2_7_10 : IN std_logic ;
         d_arr_merge2_7_9 : IN std_logic ;
         d_arr_merge2_7_8 : IN std_logic ;
         d_arr_merge2_7_7 : IN std_logic ;
         d_arr_merge2_7_6 : IN std_logic ;
         d_arr_merge2_7_5 : IN std_logic ;
         d_arr_merge2_7_4 : IN std_logic ;
         d_arr_merge2_7_3 : IN std_logic ;
         d_arr_merge2_7_2 : IN std_logic ;
         d_arr_merge2_7_1 : IN std_logic ;
         d_arr_merge2_7_0 : IN std_logic ;
         d_arr_merge2_8_31 : IN std_logic ;
         d_arr_merge2_8_30 : IN std_logic ;
         d_arr_merge2_8_29 : IN std_logic ;
         d_arr_merge2_8_28 : IN std_logic ;
         d_arr_merge2_8_27 : IN std_logic ;
         d_arr_merge2_8_26 : IN std_logic ;
         d_arr_merge2_8_25 : IN std_logic ;
         d_arr_merge2_8_24 : IN std_logic ;
         d_arr_merge2_8_23 : IN std_logic ;
         d_arr_merge2_8_22 : IN std_logic ;
         d_arr_merge2_8_21 : IN std_logic ;
         d_arr_merge2_8_20 : IN std_logic ;
         d_arr_merge2_8_19 : IN std_logic ;
         d_arr_merge2_8_18 : IN std_logic ;
         d_arr_merge2_8_17 : IN std_logic ;
         d_arr_merge2_8_16 : IN std_logic ;
         d_arr_merge2_8_15 : IN std_logic ;
         d_arr_merge2_8_14 : IN std_logic ;
         d_arr_merge2_8_13 : IN std_logic ;
         d_arr_merge2_8_12 : IN std_logic ;
         d_arr_merge2_8_11 : IN std_logic ;
         d_arr_merge2_8_10 : IN std_logic ;
         d_arr_merge2_8_9 : IN std_logic ;
         d_arr_merge2_8_8 : IN std_logic ;
         d_arr_merge2_8_7 : IN std_logic ;
         d_arr_merge2_8_6 : IN std_logic ;
         d_arr_merge2_8_5 : IN std_logic ;
         d_arr_merge2_8_4 : IN std_logic ;
         d_arr_merge2_8_3 : IN std_logic ;
         d_arr_merge2_8_2 : IN std_logic ;
         d_arr_merge2_8_1 : IN std_logic ;
         d_arr_merge2_8_0 : IN std_logic ;
         d_arr_merge2_9_31 : IN std_logic ;
         d_arr_merge2_9_30 : IN std_logic ;
         d_arr_merge2_9_29 : IN std_logic ;
         d_arr_merge2_9_28 : IN std_logic ;
         d_arr_merge2_9_27 : IN std_logic ;
         d_arr_merge2_9_26 : IN std_logic ;
         d_arr_merge2_9_25 : IN std_logic ;
         d_arr_merge2_9_24 : IN std_logic ;
         d_arr_merge2_9_23 : IN std_logic ;
         d_arr_merge2_9_22 : IN std_logic ;
         d_arr_merge2_9_21 : IN std_logic ;
         d_arr_merge2_9_20 : IN std_logic ;
         d_arr_merge2_9_19 : IN std_logic ;
         d_arr_merge2_9_18 : IN std_logic ;
         d_arr_merge2_9_17 : IN std_logic ;
         d_arr_merge2_9_16 : IN std_logic ;
         d_arr_merge2_9_15 : IN std_logic ;
         d_arr_merge2_9_14 : IN std_logic ;
         d_arr_merge2_9_13 : IN std_logic ;
         d_arr_merge2_9_12 : IN std_logic ;
         d_arr_merge2_9_11 : IN std_logic ;
         d_arr_merge2_9_10 : IN std_logic ;
         d_arr_merge2_9_9 : IN std_logic ;
         d_arr_merge2_9_8 : IN std_logic ;
         d_arr_merge2_9_7 : IN std_logic ;
         d_arr_merge2_9_6 : IN std_logic ;
         d_arr_merge2_9_5 : IN std_logic ;
         d_arr_merge2_9_4 : IN std_logic ;
         d_arr_merge2_9_3 : IN std_logic ;
         d_arr_merge2_9_2 : IN std_logic ;
         d_arr_merge2_9_1 : IN std_logic ;
         d_arr_merge2_9_0 : IN std_logic ;
         d_arr_merge2_10_31 : IN std_logic ;
         d_arr_merge2_10_30 : IN std_logic ;
         d_arr_merge2_10_29 : IN std_logic ;
         d_arr_merge2_10_28 : IN std_logic ;
         d_arr_merge2_10_27 : IN std_logic ;
         d_arr_merge2_10_26 : IN std_logic ;
         d_arr_merge2_10_25 : IN std_logic ;
         d_arr_merge2_10_24 : IN std_logic ;
         d_arr_merge2_10_23 : IN std_logic ;
         d_arr_merge2_10_22 : IN std_logic ;
         d_arr_merge2_10_21 : IN std_logic ;
         d_arr_merge2_10_20 : IN std_logic ;
         d_arr_merge2_10_19 : IN std_logic ;
         d_arr_merge2_10_18 : IN std_logic ;
         d_arr_merge2_10_17 : IN std_logic ;
         d_arr_merge2_10_16 : IN std_logic ;
         d_arr_merge2_10_15 : IN std_logic ;
         d_arr_merge2_10_14 : IN std_logic ;
         d_arr_merge2_10_13 : IN std_logic ;
         d_arr_merge2_10_12 : IN std_logic ;
         d_arr_merge2_10_11 : IN std_logic ;
         d_arr_merge2_10_10 : IN std_logic ;
         d_arr_merge2_10_9 : IN std_logic ;
         d_arr_merge2_10_8 : IN std_logic ;
         d_arr_merge2_10_7 : IN std_logic ;
         d_arr_merge2_10_6 : IN std_logic ;
         d_arr_merge2_10_5 : IN std_logic ;
         d_arr_merge2_10_4 : IN std_logic ;
         d_arr_merge2_10_3 : IN std_logic ;
         d_arr_merge2_10_2 : IN std_logic ;
         d_arr_merge2_10_1 : IN std_logic ;
         d_arr_merge2_10_0 : IN std_logic ;
         d_arr_merge2_11_31 : IN std_logic ;
         d_arr_merge2_11_30 : IN std_logic ;
         d_arr_merge2_11_29 : IN std_logic ;
         d_arr_merge2_11_28 : IN std_logic ;
         d_arr_merge2_11_27 : IN std_logic ;
         d_arr_merge2_11_26 : IN std_logic ;
         d_arr_merge2_11_25 : IN std_logic ;
         d_arr_merge2_11_24 : IN std_logic ;
         d_arr_merge2_11_23 : IN std_logic ;
         d_arr_merge2_11_22 : IN std_logic ;
         d_arr_merge2_11_21 : IN std_logic ;
         d_arr_merge2_11_20 : IN std_logic ;
         d_arr_merge2_11_19 : IN std_logic ;
         d_arr_merge2_11_18 : IN std_logic ;
         d_arr_merge2_11_17 : IN std_logic ;
         d_arr_merge2_11_16 : IN std_logic ;
         d_arr_merge2_11_15 : IN std_logic ;
         d_arr_merge2_11_14 : IN std_logic ;
         d_arr_merge2_11_13 : IN std_logic ;
         d_arr_merge2_11_12 : IN std_logic ;
         d_arr_merge2_11_11 : IN std_logic ;
         d_arr_merge2_11_10 : IN std_logic ;
         d_arr_merge2_11_9 : IN std_logic ;
         d_arr_merge2_11_8 : IN std_logic ;
         d_arr_merge2_11_7 : IN std_logic ;
         d_arr_merge2_11_6 : IN std_logic ;
         d_arr_merge2_11_5 : IN std_logic ;
         d_arr_merge2_11_4 : IN std_logic ;
         d_arr_merge2_11_3 : IN std_logic ;
         d_arr_merge2_11_2 : IN std_logic ;
         d_arr_merge2_11_1 : IN std_logic ;
         d_arr_merge2_11_0 : IN std_logic ;
         d_arr_merge2_12_31 : IN std_logic ;
         d_arr_merge2_12_30 : IN std_logic ;
         d_arr_merge2_12_29 : IN std_logic ;
         d_arr_merge2_12_28 : IN std_logic ;
         d_arr_merge2_12_27 : IN std_logic ;
         d_arr_merge2_12_26 : IN std_logic ;
         d_arr_merge2_12_25 : IN std_logic ;
         d_arr_merge2_12_24 : IN std_logic ;
         d_arr_merge2_12_23 : IN std_logic ;
         d_arr_merge2_12_22 : IN std_logic ;
         d_arr_merge2_12_21 : IN std_logic ;
         d_arr_merge2_12_20 : IN std_logic ;
         d_arr_merge2_12_19 : IN std_logic ;
         d_arr_merge2_12_18 : IN std_logic ;
         d_arr_merge2_12_17 : IN std_logic ;
         d_arr_merge2_12_16 : IN std_logic ;
         d_arr_merge2_12_15 : IN std_logic ;
         d_arr_merge2_12_14 : IN std_logic ;
         d_arr_merge2_12_13 : IN std_logic ;
         d_arr_merge2_12_12 : IN std_logic ;
         d_arr_merge2_12_11 : IN std_logic ;
         d_arr_merge2_12_10 : IN std_logic ;
         d_arr_merge2_12_9 : IN std_logic ;
         d_arr_merge2_12_8 : IN std_logic ;
         d_arr_merge2_12_7 : IN std_logic ;
         d_arr_merge2_12_6 : IN std_logic ;
         d_arr_merge2_12_5 : IN std_logic ;
         d_arr_merge2_12_4 : IN std_logic ;
         d_arr_merge2_12_3 : IN std_logic ;
         d_arr_merge2_12_2 : IN std_logic ;
         d_arr_merge2_12_1 : IN std_logic ;
         d_arr_merge2_12_0 : IN std_logic ;
         d_arr_merge2_13_31 : IN std_logic ;
         d_arr_merge2_13_30 : IN std_logic ;
         d_arr_merge2_13_29 : IN std_logic ;
         d_arr_merge2_13_28 : IN std_logic ;
         d_arr_merge2_13_27 : IN std_logic ;
         d_arr_merge2_13_26 : IN std_logic ;
         d_arr_merge2_13_25 : IN std_logic ;
         d_arr_merge2_13_24 : IN std_logic ;
         d_arr_merge2_13_23 : IN std_logic ;
         d_arr_merge2_13_22 : IN std_logic ;
         d_arr_merge2_13_21 : IN std_logic ;
         d_arr_merge2_13_20 : IN std_logic ;
         d_arr_merge2_13_19 : IN std_logic ;
         d_arr_merge2_13_18 : IN std_logic ;
         d_arr_merge2_13_17 : IN std_logic ;
         d_arr_merge2_13_16 : IN std_logic ;
         d_arr_merge2_13_15 : IN std_logic ;
         d_arr_merge2_13_14 : IN std_logic ;
         d_arr_merge2_13_13 : IN std_logic ;
         d_arr_merge2_13_12 : IN std_logic ;
         d_arr_merge2_13_11 : IN std_logic ;
         d_arr_merge2_13_10 : IN std_logic ;
         d_arr_merge2_13_9 : IN std_logic ;
         d_arr_merge2_13_8 : IN std_logic ;
         d_arr_merge2_13_7 : IN std_logic ;
         d_arr_merge2_13_6 : IN std_logic ;
         d_arr_merge2_13_5 : IN std_logic ;
         d_arr_merge2_13_4 : IN std_logic ;
         d_arr_merge2_13_3 : IN std_logic ;
         d_arr_merge2_13_2 : IN std_logic ;
         d_arr_merge2_13_1 : IN std_logic ;
         d_arr_merge2_13_0 : IN std_logic ;
         d_arr_merge2_14_31 : IN std_logic ;
         d_arr_merge2_14_30 : IN std_logic ;
         d_arr_merge2_14_29 : IN std_logic ;
         d_arr_merge2_14_28 : IN std_logic ;
         d_arr_merge2_14_27 : IN std_logic ;
         d_arr_merge2_14_26 : IN std_logic ;
         d_arr_merge2_14_25 : IN std_logic ;
         d_arr_merge2_14_24 : IN std_logic ;
         d_arr_merge2_14_23 : IN std_logic ;
         d_arr_merge2_14_22 : IN std_logic ;
         d_arr_merge2_14_21 : IN std_logic ;
         d_arr_merge2_14_20 : IN std_logic ;
         d_arr_merge2_14_19 : IN std_logic ;
         d_arr_merge2_14_18 : IN std_logic ;
         d_arr_merge2_14_17 : IN std_logic ;
         d_arr_merge2_14_16 : IN std_logic ;
         d_arr_merge2_14_15 : IN std_logic ;
         d_arr_merge2_14_14 : IN std_logic ;
         d_arr_merge2_14_13 : IN std_logic ;
         d_arr_merge2_14_12 : IN std_logic ;
         d_arr_merge2_14_11 : IN std_logic ;
         d_arr_merge2_14_10 : IN std_logic ;
         d_arr_merge2_14_9 : IN std_logic ;
         d_arr_merge2_14_8 : IN std_logic ;
         d_arr_merge2_14_7 : IN std_logic ;
         d_arr_merge2_14_6 : IN std_logic ;
         d_arr_merge2_14_5 : IN std_logic ;
         d_arr_merge2_14_4 : IN std_logic ;
         d_arr_merge2_14_3 : IN std_logic ;
         d_arr_merge2_14_2 : IN std_logic ;
         d_arr_merge2_14_1 : IN std_logic ;
         d_arr_merge2_14_0 : IN std_logic ;
         d_arr_merge2_15_31 : IN std_logic ;
         d_arr_merge2_15_30 : IN std_logic ;
         d_arr_merge2_15_29 : IN std_logic ;
         d_arr_merge2_15_28 : IN std_logic ;
         d_arr_merge2_15_27 : IN std_logic ;
         d_arr_merge2_15_26 : IN std_logic ;
         d_arr_merge2_15_25 : IN std_logic ;
         d_arr_merge2_15_24 : IN std_logic ;
         d_arr_merge2_15_23 : IN std_logic ;
         d_arr_merge2_15_22 : IN std_logic ;
         d_arr_merge2_15_21 : IN std_logic ;
         d_arr_merge2_15_20 : IN std_logic ;
         d_arr_merge2_15_19 : IN std_logic ;
         d_arr_merge2_15_18 : IN std_logic ;
         d_arr_merge2_15_17 : IN std_logic ;
         d_arr_merge2_15_16 : IN std_logic ;
         d_arr_merge2_15_15 : IN std_logic ;
         d_arr_merge2_15_14 : IN std_logic ;
         d_arr_merge2_15_13 : IN std_logic ;
         d_arr_merge2_15_12 : IN std_logic ;
         d_arr_merge2_15_11 : IN std_logic ;
         d_arr_merge2_15_10 : IN std_logic ;
         d_arr_merge2_15_9 : IN std_logic ;
         d_arr_merge2_15_8 : IN std_logic ;
         d_arr_merge2_15_7 : IN std_logic ;
         d_arr_merge2_15_6 : IN std_logic ;
         d_arr_merge2_15_5 : IN std_logic ;
         d_arr_merge2_15_4 : IN std_logic ;
         d_arr_merge2_15_3 : IN std_logic ;
         d_arr_merge2_15_2 : IN std_logic ;
         d_arr_merge2_15_1 : IN std_logic ;
         d_arr_merge2_15_0 : IN std_logic ;
         d_arr_merge2_16_31 : IN std_logic ;
         d_arr_merge2_16_30 : IN std_logic ;
         d_arr_merge2_16_29 : IN std_logic ;
         d_arr_merge2_16_28 : IN std_logic ;
         d_arr_merge2_16_27 : IN std_logic ;
         d_arr_merge2_16_26 : IN std_logic ;
         d_arr_merge2_16_25 : IN std_logic ;
         d_arr_merge2_16_24 : IN std_logic ;
         d_arr_merge2_16_23 : IN std_logic ;
         d_arr_merge2_16_22 : IN std_logic ;
         d_arr_merge2_16_21 : IN std_logic ;
         d_arr_merge2_16_20 : IN std_logic ;
         d_arr_merge2_16_19 : IN std_logic ;
         d_arr_merge2_16_18 : IN std_logic ;
         d_arr_merge2_16_17 : IN std_logic ;
         d_arr_merge2_16_16 : IN std_logic ;
         d_arr_merge2_16_15 : IN std_logic ;
         d_arr_merge2_16_14 : IN std_logic ;
         d_arr_merge2_16_13 : IN std_logic ;
         d_arr_merge2_16_12 : IN std_logic ;
         d_arr_merge2_16_11 : IN std_logic ;
         d_arr_merge2_16_10 : IN std_logic ;
         d_arr_merge2_16_9 : IN std_logic ;
         d_arr_merge2_16_8 : IN std_logic ;
         d_arr_merge2_16_7 : IN std_logic ;
         d_arr_merge2_16_6 : IN std_logic ;
         d_arr_merge2_16_5 : IN std_logic ;
         d_arr_merge2_16_4 : IN std_logic ;
         d_arr_merge2_16_3 : IN std_logic ;
         d_arr_merge2_16_2 : IN std_logic ;
         d_arr_merge2_16_1 : IN std_logic ;
         d_arr_merge2_16_0 : IN std_logic ;
         d_arr_merge2_17_31 : IN std_logic ;
         d_arr_merge2_17_30 : IN std_logic ;
         d_arr_merge2_17_29 : IN std_logic ;
         d_arr_merge2_17_28 : IN std_logic ;
         d_arr_merge2_17_27 : IN std_logic ;
         d_arr_merge2_17_26 : IN std_logic ;
         d_arr_merge2_17_25 : IN std_logic ;
         d_arr_merge2_17_24 : IN std_logic ;
         d_arr_merge2_17_23 : IN std_logic ;
         d_arr_merge2_17_22 : IN std_logic ;
         d_arr_merge2_17_21 : IN std_logic ;
         d_arr_merge2_17_20 : IN std_logic ;
         d_arr_merge2_17_19 : IN std_logic ;
         d_arr_merge2_17_18 : IN std_logic ;
         d_arr_merge2_17_17 : IN std_logic ;
         d_arr_merge2_17_16 : IN std_logic ;
         d_arr_merge2_17_15 : IN std_logic ;
         d_arr_merge2_17_14 : IN std_logic ;
         d_arr_merge2_17_13 : IN std_logic ;
         d_arr_merge2_17_12 : IN std_logic ;
         d_arr_merge2_17_11 : IN std_logic ;
         d_arr_merge2_17_10 : IN std_logic ;
         d_arr_merge2_17_9 : IN std_logic ;
         d_arr_merge2_17_8 : IN std_logic ;
         d_arr_merge2_17_7 : IN std_logic ;
         d_arr_merge2_17_6 : IN std_logic ;
         d_arr_merge2_17_5 : IN std_logic ;
         d_arr_merge2_17_4 : IN std_logic ;
         d_arr_merge2_17_3 : IN std_logic ;
         d_arr_merge2_17_2 : IN std_logic ;
         d_arr_merge2_17_1 : IN std_logic ;
         d_arr_merge2_17_0 : IN std_logic ;
         d_arr_merge2_18_31 : IN std_logic ;
         d_arr_merge2_18_30 : IN std_logic ;
         d_arr_merge2_18_29 : IN std_logic ;
         d_arr_merge2_18_28 : IN std_logic ;
         d_arr_merge2_18_27 : IN std_logic ;
         d_arr_merge2_18_26 : IN std_logic ;
         d_arr_merge2_18_25 : IN std_logic ;
         d_arr_merge2_18_24 : IN std_logic ;
         d_arr_merge2_18_23 : IN std_logic ;
         d_arr_merge2_18_22 : IN std_logic ;
         d_arr_merge2_18_21 : IN std_logic ;
         d_arr_merge2_18_20 : IN std_logic ;
         d_arr_merge2_18_19 : IN std_logic ;
         d_arr_merge2_18_18 : IN std_logic ;
         d_arr_merge2_18_17 : IN std_logic ;
         d_arr_merge2_18_16 : IN std_logic ;
         d_arr_merge2_18_15 : IN std_logic ;
         d_arr_merge2_18_14 : IN std_logic ;
         d_arr_merge2_18_13 : IN std_logic ;
         d_arr_merge2_18_12 : IN std_logic ;
         d_arr_merge2_18_11 : IN std_logic ;
         d_arr_merge2_18_10 : IN std_logic ;
         d_arr_merge2_18_9 : IN std_logic ;
         d_arr_merge2_18_8 : IN std_logic ;
         d_arr_merge2_18_7 : IN std_logic ;
         d_arr_merge2_18_6 : IN std_logic ;
         d_arr_merge2_18_5 : IN std_logic ;
         d_arr_merge2_18_4 : IN std_logic ;
         d_arr_merge2_18_3 : IN std_logic ;
         d_arr_merge2_18_2 : IN std_logic ;
         d_arr_merge2_18_1 : IN std_logic ;
         d_arr_merge2_18_0 : IN std_logic ;
         d_arr_merge2_19_31 : IN std_logic ;
         d_arr_merge2_19_30 : IN std_logic ;
         d_arr_merge2_19_29 : IN std_logic ;
         d_arr_merge2_19_28 : IN std_logic ;
         d_arr_merge2_19_27 : IN std_logic ;
         d_arr_merge2_19_26 : IN std_logic ;
         d_arr_merge2_19_25 : IN std_logic ;
         d_arr_merge2_19_24 : IN std_logic ;
         d_arr_merge2_19_23 : IN std_logic ;
         d_arr_merge2_19_22 : IN std_logic ;
         d_arr_merge2_19_21 : IN std_logic ;
         d_arr_merge2_19_20 : IN std_logic ;
         d_arr_merge2_19_19 : IN std_logic ;
         d_arr_merge2_19_18 : IN std_logic ;
         d_arr_merge2_19_17 : IN std_logic ;
         d_arr_merge2_19_16 : IN std_logic ;
         d_arr_merge2_19_15 : IN std_logic ;
         d_arr_merge2_19_14 : IN std_logic ;
         d_arr_merge2_19_13 : IN std_logic ;
         d_arr_merge2_19_12 : IN std_logic ;
         d_arr_merge2_19_11 : IN std_logic ;
         d_arr_merge2_19_10 : IN std_logic ;
         d_arr_merge2_19_9 : IN std_logic ;
         d_arr_merge2_19_8 : IN std_logic ;
         d_arr_merge2_19_7 : IN std_logic ;
         d_arr_merge2_19_6 : IN std_logic ;
         d_arr_merge2_19_5 : IN std_logic ;
         d_arr_merge2_19_4 : IN std_logic ;
         d_arr_merge2_19_3 : IN std_logic ;
         d_arr_merge2_19_2 : IN std_logic ;
         d_arr_merge2_19_1 : IN std_logic ;
         d_arr_merge2_19_0 : IN std_logic ;
         d_arr_merge2_20_31 : IN std_logic ;
         d_arr_merge2_20_30 : IN std_logic ;
         d_arr_merge2_20_29 : IN std_logic ;
         d_arr_merge2_20_28 : IN std_logic ;
         d_arr_merge2_20_27 : IN std_logic ;
         d_arr_merge2_20_26 : IN std_logic ;
         d_arr_merge2_20_25 : IN std_logic ;
         d_arr_merge2_20_24 : IN std_logic ;
         d_arr_merge2_20_23 : IN std_logic ;
         d_arr_merge2_20_22 : IN std_logic ;
         d_arr_merge2_20_21 : IN std_logic ;
         d_arr_merge2_20_20 : IN std_logic ;
         d_arr_merge2_20_19 : IN std_logic ;
         d_arr_merge2_20_18 : IN std_logic ;
         d_arr_merge2_20_17 : IN std_logic ;
         d_arr_merge2_20_16 : IN std_logic ;
         d_arr_merge2_20_15 : IN std_logic ;
         d_arr_merge2_20_14 : IN std_logic ;
         d_arr_merge2_20_13 : IN std_logic ;
         d_arr_merge2_20_12 : IN std_logic ;
         d_arr_merge2_20_11 : IN std_logic ;
         d_arr_merge2_20_10 : IN std_logic ;
         d_arr_merge2_20_9 : IN std_logic ;
         d_arr_merge2_20_8 : IN std_logic ;
         d_arr_merge2_20_7 : IN std_logic ;
         d_arr_merge2_20_6 : IN std_logic ;
         d_arr_merge2_20_5 : IN std_logic ;
         d_arr_merge2_20_4 : IN std_logic ;
         d_arr_merge2_20_3 : IN std_logic ;
         d_arr_merge2_20_2 : IN std_logic ;
         d_arr_merge2_20_1 : IN std_logic ;
         d_arr_merge2_20_0 : IN std_logic ;
         d_arr_merge2_21_31 : IN std_logic ;
         d_arr_merge2_21_30 : IN std_logic ;
         d_arr_merge2_21_29 : IN std_logic ;
         d_arr_merge2_21_28 : IN std_logic ;
         d_arr_merge2_21_27 : IN std_logic ;
         d_arr_merge2_21_26 : IN std_logic ;
         d_arr_merge2_21_25 : IN std_logic ;
         d_arr_merge2_21_24 : IN std_logic ;
         d_arr_merge2_21_23 : IN std_logic ;
         d_arr_merge2_21_22 : IN std_logic ;
         d_arr_merge2_21_21 : IN std_logic ;
         d_arr_merge2_21_20 : IN std_logic ;
         d_arr_merge2_21_19 : IN std_logic ;
         d_arr_merge2_21_18 : IN std_logic ;
         d_arr_merge2_21_17 : IN std_logic ;
         d_arr_merge2_21_16 : IN std_logic ;
         d_arr_merge2_21_15 : IN std_logic ;
         d_arr_merge2_21_14 : IN std_logic ;
         d_arr_merge2_21_13 : IN std_logic ;
         d_arr_merge2_21_12 : IN std_logic ;
         d_arr_merge2_21_11 : IN std_logic ;
         d_arr_merge2_21_10 : IN std_logic ;
         d_arr_merge2_21_9 : IN std_logic ;
         d_arr_merge2_21_8 : IN std_logic ;
         d_arr_merge2_21_7 : IN std_logic ;
         d_arr_merge2_21_6 : IN std_logic ;
         d_arr_merge2_21_5 : IN std_logic ;
         d_arr_merge2_21_4 : IN std_logic ;
         d_arr_merge2_21_3 : IN std_logic ;
         d_arr_merge2_21_2 : IN std_logic ;
         d_arr_merge2_21_1 : IN std_logic ;
         d_arr_merge2_21_0 : IN std_logic ;
         d_arr_merge2_22_31 : IN std_logic ;
         d_arr_merge2_22_30 : IN std_logic ;
         d_arr_merge2_22_29 : IN std_logic ;
         d_arr_merge2_22_28 : IN std_logic ;
         d_arr_merge2_22_27 : IN std_logic ;
         d_arr_merge2_22_26 : IN std_logic ;
         d_arr_merge2_22_25 : IN std_logic ;
         d_arr_merge2_22_24 : IN std_logic ;
         d_arr_merge2_22_23 : IN std_logic ;
         d_arr_merge2_22_22 : IN std_logic ;
         d_arr_merge2_22_21 : IN std_logic ;
         d_arr_merge2_22_20 : IN std_logic ;
         d_arr_merge2_22_19 : IN std_logic ;
         d_arr_merge2_22_18 : IN std_logic ;
         d_arr_merge2_22_17 : IN std_logic ;
         d_arr_merge2_22_16 : IN std_logic ;
         d_arr_merge2_22_15 : IN std_logic ;
         d_arr_merge2_22_14 : IN std_logic ;
         d_arr_merge2_22_13 : IN std_logic ;
         d_arr_merge2_22_12 : IN std_logic ;
         d_arr_merge2_22_11 : IN std_logic ;
         d_arr_merge2_22_10 : IN std_logic ;
         d_arr_merge2_22_9 : IN std_logic ;
         d_arr_merge2_22_8 : IN std_logic ;
         d_arr_merge2_22_7 : IN std_logic ;
         d_arr_merge2_22_6 : IN std_logic ;
         d_arr_merge2_22_5 : IN std_logic ;
         d_arr_merge2_22_4 : IN std_logic ;
         d_arr_merge2_22_3 : IN std_logic ;
         d_arr_merge2_22_2 : IN std_logic ;
         d_arr_merge2_22_1 : IN std_logic ;
         d_arr_merge2_22_0 : IN std_logic ;
         d_arr_merge2_23_31 : IN std_logic ;
         d_arr_merge2_23_30 : IN std_logic ;
         d_arr_merge2_23_29 : IN std_logic ;
         d_arr_merge2_23_28 : IN std_logic ;
         d_arr_merge2_23_27 : IN std_logic ;
         d_arr_merge2_23_26 : IN std_logic ;
         d_arr_merge2_23_25 : IN std_logic ;
         d_arr_merge2_23_24 : IN std_logic ;
         d_arr_merge2_23_23 : IN std_logic ;
         d_arr_merge2_23_22 : IN std_logic ;
         d_arr_merge2_23_21 : IN std_logic ;
         d_arr_merge2_23_20 : IN std_logic ;
         d_arr_merge2_23_19 : IN std_logic ;
         d_arr_merge2_23_18 : IN std_logic ;
         d_arr_merge2_23_17 : IN std_logic ;
         d_arr_merge2_23_16 : IN std_logic ;
         d_arr_merge2_23_15 : IN std_logic ;
         d_arr_merge2_23_14 : IN std_logic ;
         d_arr_merge2_23_13 : IN std_logic ;
         d_arr_merge2_23_12 : IN std_logic ;
         d_arr_merge2_23_11 : IN std_logic ;
         d_arr_merge2_23_10 : IN std_logic ;
         d_arr_merge2_23_9 : IN std_logic ;
         d_arr_merge2_23_8 : IN std_logic ;
         d_arr_merge2_23_7 : IN std_logic ;
         d_arr_merge2_23_6 : IN std_logic ;
         d_arr_merge2_23_5 : IN std_logic ;
         d_arr_merge2_23_4 : IN std_logic ;
         d_arr_merge2_23_3 : IN std_logic ;
         d_arr_merge2_23_2 : IN std_logic ;
         d_arr_merge2_23_1 : IN std_logic ;
         d_arr_merge2_23_0 : IN std_logic ;
         d_arr_merge2_24_31 : IN std_logic ;
         d_arr_merge2_24_30 : IN std_logic ;
         d_arr_merge2_24_29 : IN std_logic ;
         d_arr_merge2_24_28 : IN std_logic ;
         d_arr_merge2_24_27 : IN std_logic ;
         d_arr_merge2_24_26 : IN std_logic ;
         d_arr_merge2_24_25 : IN std_logic ;
         d_arr_merge2_24_24 : IN std_logic ;
         d_arr_merge2_24_23 : IN std_logic ;
         d_arr_merge2_24_22 : IN std_logic ;
         d_arr_merge2_24_21 : IN std_logic ;
         d_arr_merge2_24_20 : IN std_logic ;
         d_arr_merge2_24_19 : IN std_logic ;
         d_arr_merge2_24_18 : IN std_logic ;
         d_arr_merge2_24_17 : IN std_logic ;
         d_arr_merge2_24_16 : IN std_logic ;
         d_arr_merge2_24_15 : IN std_logic ;
         d_arr_merge2_24_14 : IN std_logic ;
         d_arr_merge2_24_13 : IN std_logic ;
         d_arr_merge2_24_12 : IN std_logic ;
         d_arr_merge2_24_11 : IN std_logic ;
         d_arr_merge2_24_10 : IN std_logic ;
         d_arr_merge2_24_9 : IN std_logic ;
         d_arr_merge2_24_8 : IN std_logic ;
         d_arr_merge2_24_7 : IN std_logic ;
         d_arr_merge2_24_6 : IN std_logic ;
         d_arr_merge2_24_5 : IN std_logic ;
         d_arr_merge2_24_4 : IN std_logic ;
         d_arr_merge2_24_3 : IN std_logic ;
         d_arr_merge2_24_2 : IN std_logic ;
         d_arr_merge2_24_1 : IN std_logic ;
         d_arr_merge2_24_0 : IN std_logic ;
         d_arr_relu_0_31 : IN std_logic ;
         d_arr_relu_0_30 : IN std_logic ;
         d_arr_relu_0_29 : IN std_logic ;
         d_arr_relu_0_28 : IN std_logic ;
         d_arr_relu_0_27 : IN std_logic ;
         d_arr_relu_0_26 : IN std_logic ;
         d_arr_relu_0_25 : IN std_logic ;
         d_arr_relu_0_24 : IN std_logic ;
         d_arr_relu_0_23 : IN std_logic ;
         d_arr_relu_0_22 : IN std_logic ;
         d_arr_relu_0_21 : IN std_logic ;
         d_arr_relu_0_20 : IN std_logic ;
         d_arr_relu_0_19 : IN std_logic ;
         d_arr_relu_0_18 : IN std_logic ;
         d_arr_relu_0_17 : IN std_logic ;
         d_arr_relu_0_16 : IN std_logic ;
         d_arr_relu_0_15 : IN std_logic ;
         d_arr_relu_0_14 : IN std_logic ;
         d_arr_relu_0_13 : IN std_logic ;
         d_arr_relu_0_12 : IN std_logic ;
         d_arr_relu_0_11 : IN std_logic ;
         d_arr_relu_0_10 : IN std_logic ;
         d_arr_relu_0_9 : IN std_logic ;
         d_arr_relu_0_8 : IN std_logic ;
         d_arr_relu_0_7 : IN std_logic ;
         d_arr_relu_0_6 : IN std_logic ;
         d_arr_relu_0_5 : IN std_logic ;
         d_arr_relu_0_4 : IN std_logic ;
         d_arr_relu_0_3 : IN std_logic ;
         d_arr_relu_0_2 : IN std_logic ;
         d_arr_relu_0_1 : IN std_logic ;
         d_arr_relu_0_0 : IN std_logic ;
         d_arr_relu_1_31 : IN std_logic ;
         d_arr_relu_1_30 : IN std_logic ;
         d_arr_relu_1_29 : IN std_logic ;
         d_arr_relu_1_28 : IN std_logic ;
         d_arr_relu_1_27 : IN std_logic ;
         d_arr_relu_1_26 : IN std_logic ;
         d_arr_relu_1_25 : IN std_logic ;
         d_arr_relu_1_24 : IN std_logic ;
         d_arr_relu_1_23 : IN std_logic ;
         d_arr_relu_1_22 : IN std_logic ;
         d_arr_relu_1_21 : IN std_logic ;
         d_arr_relu_1_20 : IN std_logic ;
         d_arr_relu_1_19 : IN std_logic ;
         d_arr_relu_1_18 : IN std_logic ;
         d_arr_relu_1_17 : IN std_logic ;
         d_arr_relu_1_16 : IN std_logic ;
         d_arr_relu_1_15 : IN std_logic ;
         d_arr_relu_1_14 : IN std_logic ;
         d_arr_relu_1_13 : IN std_logic ;
         d_arr_relu_1_12 : IN std_logic ;
         d_arr_relu_1_11 : IN std_logic ;
         d_arr_relu_1_10 : IN std_logic ;
         d_arr_relu_1_9 : IN std_logic ;
         d_arr_relu_1_8 : IN std_logic ;
         d_arr_relu_1_7 : IN std_logic ;
         d_arr_relu_1_6 : IN std_logic ;
         d_arr_relu_1_5 : IN std_logic ;
         d_arr_relu_1_4 : IN std_logic ;
         d_arr_relu_1_3 : IN std_logic ;
         d_arr_relu_1_2 : IN std_logic ;
         d_arr_relu_1_1 : IN std_logic ;
         d_arr_relu_1_0 : IN std_logic ;
         d_arr_relu_2_31 : IN std_logic ;
         d_arr_relu_2_30 : IN std_logic ;
         d_arr_relu_2_29 : IN std_logic ;
         d_arr_relu_2_28 : IN std_logic ;
         d_arr_relu_2_27 : IN std_logic ;
         d_arr_relu_2_26 : IN std_logic ;
         d_arr_relu_2_25 : IN std_logic ;
         d_arr_relu_2_24 : IN std_logic ;
         d_arr_relu_2_23 : IN std_logic ;
         d_arr_relu_2_22 : IN std_logic ;
         d_arr_relu_2_21 : IN std_logic ;
         d_arr_relu_2_20 : IN std_logic ;
         d_arr_relu_2_19 : IN std_logic ;
         d_arr_relu_2_18 : IN std_logic ;
         d_arr_relu_2_17 : IN std_logic ;
         d_arr_relu_2_16 : IN std_logic ;
         d_arr_relu_2_15 : IN std_logic ;
         d_arr_relu_2_14 : IN std_logic ;
         d_arr_relu_2_13 : IN std_logic ;
         d_arr_relu_2_12 : IN std_logic ;
         d_arr_relu_2_11 : IN std_logic ;
         d_arr_relu_2_10 : IN std_logic ;
         d_arr_relu_2_9 : IN std_logic ;
         d_arr_relu_2_8 : IN std_logic ;
         d_arr_relu_2_7 : IN std_logic ;
         d_arr_relu_2_6 : IN std_logic ;
         d_arr_relu_2_5 : IN std_logic ;
         d_arr_relu_2_4 : IN std_logic ;
         d_arr_relu_2_3 : IN std_logic ;
         d_arr_relu_2_2 : IN std_logic ;
         d_arr_relu_2_1 : IN std_logic ;
         d_arr_relu_2_0 : IN std_logic ;
         d_arr_relu_3_31 : IN std_logic ;
         d_arr_relu_3_30 : IN std_logic ;
         d_arr_relu_3_29 : IN std_logic ;
         d_arr_relu_3_28 : IN std_logic ;
         d_arr_relu_3_27 : IN std_logic ;
         d_arr_relu_3_26 : IN std_logic ;
         d_arr_relu_3_25 : IN std_logic ;
         d_arr_relu_3_24 : IN std_logic ;
         d_arr_relu_3_23 : IN std_logic ;
         d_arr_relu_3_22 : IN std_logic ;
         d_arr_relu_3_21 : IN std_logic ;
         d_arr_relu_3_20 : IN std_logic ;
         d_arr_relu_3_19 : IN std_logic ;
         d_arr_relu_3_18 : IN std_logic ;
         d_arr_relu_3_17 : IN std_logic ;
         d_arr_relu_3_16 : IN std_logic ;
         d_arr_relu_3_15 : IN std_logic ;
         d_arr_relu_3_14 : IN std_logic ;
         d_arr_relu_3_13 : IN std_logic ;
         d_arr_relu_3_12 : IN std_logic ;
         d_arr_relu_3_11 : IN std_logic ;
         d_arr_relu_3_10 : IN std_logic ;
         d_arr_relu_3_9 : IN std_logic ;
         d_arr_relu_3_8 : IN std_logic ;
         d_arr_relu_3_7 : IN std_logic ;
         d_arr_relu_3_6 : IN std_logic ;
         d_arr_relu_3_5 : IN std_logic ;
         d_arr_relu_3_4 : IN std_logic ;
         d_arr_relu_3_3 : IN std_logic ;
         d_arr_relu_3_2 : IN std_logic ;
         d_arr_relu_3_1 : IN std_logic ;
         d_arr_relu_3_0 : IN std_logic ;
         d_arr_relu_4_31 : IN std_logic ;
         d_arr_relu_4_30 : IN std_logic ;
         d_arr_relu_4_29 : IN std_logic ;
         d_arr_relu_4_28 : IN std_logic ;
         d_arr_relu_4_27 : IN std_logic ;
         d_arr_relu_4_26 : IN std_logic ;
         d_arr_relu_4_25 : IN std_logic ;
         d_arr_relu_4_24 : IN std_logic ;
         d_arr_relu_4_23 : IN std_logic ;
         d_arr_relu_4_22 : IN std_logic ;
         d_arr_relu_4_21 : IN std_logic ;
         d_arr_relu_4_20 : IN std_logic ;
         d_arr_relu_4_19 : IN std_logic ;
         d_arr_relu_4_18 : IN std_logic ;
         d_arr_relu_4_17 : IN std_logic ;
         d_arr_relu_4_16 : IN std_logic ;
         d_arr_relu_4_15 : IN std_logic ;
         d_arr_relu_4_14 : IN std_logic ;
         d_arr_relu_4_13 : IN std_logic ;
         d_arr_relu_4_12 : IN std_logic ;
         d_arr_relu_4_11 : IN std_logic ;
         d_arr_relu_4_10 : IN std_logic ;
         d_arr_relu_4_9 : IN std_logic ;
         d_arr_relu_4_8 : IN std_logic ;
         d_arr_relu_4_7 : IN std_logic ;
         d_arr_relu_4_6 : IN std_logic ;
         d_arr_relu_4_5 : IN std_logic ;
         d_arr_relu_4_4 : IN std_logic ;
         d_arr_relu_4_3 : IN std_logic ;
         d_arr_relu_4_2 : IN std_logic ;
         d_arr_relu_4_1 : IN std_logic ;
         d_arr_relu_4_0 : IN std_logic ;
         d_arr_relu_5_31 : IN std_logic ;
         d_arr_relu_5_30 : IN std_logic ;
         d_arr_relu_5_29 : IN std_logic ;
         d_arr_relu_5_28 : IN std_logic ;
         d_arr_relu_5_27 : IN std_logic ;
         d_arr_relu_5_26 : IN std_logic ;
         d_arr_relu_5_25 : IN std_logic ;
         d_arr_relu_5_24 : IN std_logic ;
         d_arr_relu_5_23 : IN std_logic ;
         d_arr_relu_5_22 : IN std_logic ;
         d_arr_relu_5_21 : IN std_logic ;
         d_arr_relu_5_20 : IN std_logic ;
         d_arr_relu_5_19 : IN std_logic ;
         d_arr_relu_5_18 : IN std_logic ;
         d_arr_relu_5_17 : IN std_logic ;
         d_arr_relu_5_16 : IN std_logic ;
         d_arr_relu_5_15 : IN std_logic ;
         d_arr_relu_5_14 : IN std_logic ;
         d_arr_relu_5_13 : IN std_logic ;
         d_arr_relu_5_12 : IN std_logic ;
         d_arr_relu_5_11 : IN std_logic ;
         d_arr_relu_5_10 : IN std_logic ;
         d_arr_relu_5_9 : IN std_logic ;
         d_arr_relu_5_8 : IN std_logic ;
         d_arr_relu_5_7 : IN std_logic ;
         d_arr_relu_5_6 : IN std_logic ;
         d_arr_relu_5_5 : IN std_logic ;
         d_arr_relu_5_4 : IN std_logic ;
         d_arr_relu_5_3 : IN std_logic ;
         d_arr_relu_5_2 : IN std_logic ;
         d_arr_relu_5_1 : IN std_logic ;
         d_arr_relu_5_0 : IN std_logic ;
         d_arr_relu_6_31 : IN std_logic ;
         d_arr_relu_6_30 : IN std_logic ;
         d_arr_relu_6_29 : IN std_logic ;
         d_arr_relu_6_28 : IN std_logic ;
         d_arr_relu_6_27 : IN std_logic ;
         d_arr_relu_6_26 : IN std_logic ;
         d_arr_relu_6_25 : IN std_logic ;
         d_arr_relu_6_24 : IN std_logic ;
         d_arr_relu_6_23 : IN std_logic ;
         d_arr_relu_6_22 : IN std_logic ;
         d_arr_relu_6_21 : IN std_logic ;
         d_arr_relu_6_20 : IN std_logic ;
         d_arr_relu_6_19 : IN std_logic ;
         d_arr_relu_6_18 : IN std_logic ;
         d_arr_relu_6_17 : IN std_logic ;
         d_arr_relu_6_16 : IN std_logic ;
         d_arr_relu_6_15 : IN std_logic ;
         d_arr_relu_6_14 : IN std_logic ;
         d_arr_relu_6_13 : IN std_logic ;
         d_arr_relu_6_12 : IN std_logic ;
         d_arr_relu_6_11 : IN std_logic ;
         d_arr_relu_6_10 : IN std_logic ;
         d_arr_relu_6_9 : IN std_logic ;
         d_arr_relu_6_8 : IN std_logic ;
         d_arr_relu_6_7 : IN std_logic ;
         d_arr_relu_6_6 : IN std_logic ;
         d_arr_relu_6_5 : IN std_logic ;
         d_arr_relu_6_4 : IN std_logic ;
         d_arr_relu_6_3 : IN std_logic ;
         d_arr_relu_6_2 : IN std_logic ;
         d_arr_relu_6_1 : IN std_logic ;
         d_arr_relu_6_0 : IN std_logic ;
         d_arr_relu_7_31 : IN std_logic ;
         d_arr_relu_7_30 : IN std_logic ;
         d_arr_relu_7_29 : IN std_logic ;
         d_arr_relu_7_28 : IN std_logic ;
         d_arr_relu_7_27 : IN std_logic ;
         d_arr_relu_7_26 : IN std_logic ;
         d_arr_relu_7_25 : IN std_logic ;
         d_arr_relu_7_24 : IN std_logic ;
         d_arr_relu_7_23 : IN std_logic ;
         d_arr_relu_7_22 : IN std_logic ;
         d_arr_relu_7_21 : IN std_logic ;
         d_arr_relu_7_20 : IN std_logic ;
         d_arr_relu_7_19 : IN std_logic ;
         d_arr_relu_7_18 : IN std_logic ;
         d_arr_relu_7_17 : IN std_logic ;
         d_arr_relu_7_16 : IN std_logic ;
         d_arr_relu_7_15 : IN std_logic ;
         d_arr_relu_7_14 : IN std_logic ;
         d_arr_relu_7_13 : IN std_logic ;
         d_arr_relu_7_12 : IN std_logic ;
         d_arr_relu_7_11 : IN std_logic ;
         d_arr_relu_7_10 : IN std_logic ;
         d_arr_relu_7_9 : IN std_logic ;
         d_arr_relu_7_8 : IN std_logic ;
         d_arr_relu_7_7 : IN std_logic ;
         d_arr_relu_7_6 : IN std_logic ;
         d_arr_relu_7_5 : IN std_logic ;
         d_arr_relu_7_4 : IN std_logic ;
         d_arr_relu_7_3 : IN std_logic ;
         d_arr_relu_7_2 : IN std_logic ;
         d_arr_relu_7_1 : IN std_logic ;
         d_arr_relu_7_0 : IN std_logic ;
         d_arr_relu_8_31 : IN std_logic ;
         d_arr_relu_8_30 : IN std_logic ;
         d_arr_relu_8_29 : IN std_logic ;
         d_arr_relu_8_28 : IN std_logic ;
         d_arr_relu_8_27 : IN std_logic ;
         d_arr_relu_8_26 : IN std_logic ;
         d_arr_relu_8_25 : IN std_logic ;
         d_arr_relu_8_24 : IN std_logic ;
         d_arr_relu_8_23 : IN std_logic ;
         d_arr_relu_8_22 : IN std_logic ;
         d_arr_relu_8_21 : IN std_logic ;
         d_arr_relu_8_20 : IN std_logic ;
         d_arr_relu_8_19 : IN std_logic ;
         d_arr_relu_8_18 : IN std_logic ;
         d_arr_relu_8_17 : IN std_logic ;
         d_arr_relu_8_16 : IN std_logic ;
         d_arr_relu_8_15 : IN std_logic ;
         d_arr_relu_8_14 : IN std_logic ;
         d_arr_relu_8_13 : IN std_logic ;
         d_arr_relu_8_12 : IN std_logic ;
         d_arr_relu_8_11 : IN std_logic ;
         d_arr_relu_8_10 : IN std_logic ;
         d_arr_relu_8_9 : IN std_logic ;
         d_arr_relu_8_8 : IN std_logic ;
         d_arr_relu_8_7 : IN std_logic ;
         d_arr_relu_8_6 : IN std_logic ;
         d_arr_relu_8_5 : IN std_logic ;
         d_arr_relu_8_4 : IN std_logic ;
         d_arr_relu_8_3 : IN std_logic ;
         d_arr_relu_8_2 : IN std_logic ;
         d_arr_relu_8_1 : IN std_logic ;
         d_arr_relu_8_0 : IN std_logic ;
         d_arr_relu_9_31 : IN std_logic ;
         d_arr_relu_9_30 : IN std_logic ;
         d_arr_relu_9_29 : IN std_logic ;
         d_arr_relu_9_28 : IN std_logic ;
         d_arr_relu_9_27 : IN std_logic ;
         d_arr_relu_9_26 : IN std_logic ;
         d_arr_relu_9_25 : IN std_logic ;
         d_arr_relu_9_24 : IN std_logic ;
         d_arr_relu_9_23 : IN std_logic ;
         d_arr_relu_9_22 : IN std_logic ;
         d_arr_relu_9_21 : IN std_logic ;
         d_arr_relu_9_20 : IN std_logic ;
         d_arr_relu_9_19 : IN std_logic ;
         d_arr_relu_9_18 : IN std_logic ;
         d_arr_relu_9_17 : IN std_logic ;
         d_arr_relu_9_16 : IN std_logic ;
         d_arr_relu_9_15 : IN std_logic ;
         d_arr_relu_9_14 : IN std_logic ;
         d_arr_relu_9_13 : IN std_logic ;
         d_arr_relu_9_12 : IN std_logic ;
         d_arr_relu_9_11 : IN std_logic ;
         d_arr_relu_9_10 : IN std_logic ;
         d_arr_relu_9_9 : IN std_logic ;
         d_arr_relu_9_8 : IN std_logic ;
         d_arr_relu_9_7 : IN std_logic ;
         d_arr_relu_9_6 : IN std_logic ;
         d_arr_relu_9_5 : IN std_logic ;
         d_arr_relu_9_4 : IN std_logic ;
         d_arr_relu_9_3 : IN std_logic ;
         d_arr_relu_9_2 : IN std_logic ;
         d_arr_relu_9_1 : IN std_logic ;
         d_arr_relu_9_0 : IN std_logic ;
         d_arr_relu_10_31 : IN std_logic ;
         d_arr_relu_10_30 : IN std_logic ;
         d_arr_relu_10_29 : IN std_logic ;
         d_arr_relu_10_28 : IN std_logic ;
         d_arr_relu_10_27 : IN std_logic ;
         d_arr_relu_10_26 : IN std_logic ;
         d_arr_relu_10_25 : IN std_logic ;
         d_arr_relu_10_24 : IN std_logic ;
         d_arr_relu_10_23 : IN std_logic ;
         d_arr_relu_10_22 : IN std_logic ;
         d_arr_relu_10_21 : IN std_logic ;
         d_arr_relu_10_20 : IN std_logic ;
         d_arr_relu_10_19 : IN std_logic ;
         d_arr_relu_10_18 : IN std_logic ;
         d_arr_relu_10_17 : IN std_logic ;
         d_arr_relu_10_16 : IN std_logic ;
         d_arr_relu_10_15 : IN std_logic ;
         d_arr_relu_10_14 : IN std_logic ;
         d_arr_relu_10_13 : IN std_logic ;
         d_arr_relu_10_12 : IN std_logic ;
         d_arr_relu_10_11 : IN std_logic ;
         d_arr_relu_10_10 : IN std_logic ;
         d_arr_relu_10_9 : IN std_logic ;
         d_arr_relu_10_8 : IN std_logic ;
         d_arr_relu_10_7 : IN std_logic ;
         d_arr_relu_10_6 : IN std_logic ;
         d_arr_relu_10_5 : IN std_logic ;
         d_arr_relu_10_4 : IN std_logic ;
         d_arr_relu_10_3 : IN std_logic ;
         d_arr_relu_10_2 : IN std_logic ;
         d_arr_relu_10_1 : IN std_logic ;
         d_arr_relu_10_0 : IN std_logic ;
         d_arr_relu_11_31 : IN std_logic ;
         d_arr_relu_11_30 : IN std_logic ;
         d_arr_relu_11_29 : IN std_logic ;
         d_arr_relu_11_28 : IN std_logic ;
         d_arr_relu_11_27 : IN std_logic ;
         d_arr_relu_11_26 : IN std_logic ;
         d_arr_relu_11_25 : IN std_logic ;
         d_arr_relu_11_24 : IN std_logic ;
         d_arr_relu_11_23 : IN std_logic ;
         d_arr_relu_11_22 : IN std_logic ;
         d_arr_relu_11_21 : IN std_logic ;
         d_arr_relu_11_20 : IN std_logic ;
         d_arr_relu_11_19 : IN std_logic ;
         d_arr_relu_11_18 : IN std_logic ;
         d_arr_relu_11_17 : IN std_logic ;
         d_arr_relu_11_16 : IN std_logic ;
         d_arr_relu_11_15 : IN std_logic ;
         d_arr_relu_11_14 : IN std_logic ;
         d_arr_relu_11_13 : IN std_logic ;
         d_arr_relu_11_12 : IN std_logic ;
         d_arr_relu_11_11 : IN std_logic ;
         d_arr_relu_11_10 : IN std_logic ;
         d_arr_relu_11_9 : IN std_logic ;
         d_arr_relu_11_8 : IN std_logic ;
         d_arr_relu_11_7 : IN std_logic ;
         d_arr_relu_11_6 : IN std_logic ;
         d_arr_relu_11_5 : IN std_logic ;
         d_arr_relu_11_4 : IN std_logic ;
         d_arr_relu_11_3 : IN std_logic ;
         d_arr_relu_11_2 : IN std_logic ;
         d_arr_relu_11_1 : IN std_logic ;
         d_arr_relu_11_0 : IN std_logic ;
         d_arr_relu_12_31 : IN std_logic ;
         d_arr_relu_12_30 : IN std_logic ;
         d_arr_relu_12_29 : IN std_logic ;
         d_arr_relu_12_28 : IN std_logic ;
         d_arr_relu_12_27 : IN std_logic ;
         d_arr_relu_12_26 : IN std_logic ;
         d_arr_relu_12_25 : IN std_logic ;
         d_arr_relu_12_24 : IN std_logic ;
         d_arr_relu_12_23 : IN std_logic ;
         d_arr_relu_12_22 : IN std_logic ;
         d_arr_relu_12_21 : IN std_logic ;
         d_arr_relu_12_20 : IN std_logic ;
         d_arr_relu_12_19 : IN std_logic ;
         d_arr_relu_12_18 : IN std_logic ;
         d_arr_relu_12_17 : IN std_logic ;
         d_arr_relu_12_16 : IN std_logic ;
         d_arr_relu_12_15 : IN std_logic ;
         d_arr_relu_12_14 : IN std_logic ;
         d_arr_relu_12_13 : IN std_logic ;
         d_arr_relu_12_12 : IN std_logic ;
         d_arr_relu_12_11 : IN std_logic ;
         d_arr_relu_12_10 : IN std_logic ;
         d_arr_relu_12_9 : IN std_logic ;
         d_arr_relu_12_8 : IN std_logic ;
         d_arr_relu_12_7 : IN std_logic ;
         d_arr_relu_12_6 : IN std_logic ;
         d_arr_relu_12_5 : IN std_logic ;
         d_arr_relu_12_4 : IN std_logic ;
         d_arr_relu_12_3 : IN std_logic ;
         d_arr_relu_12_2 : IN std_logic ;
         d_arr_relu_12_1 : IN std_logic ;
         d_arr_relu_12_0 : IN std_logic ;
         d_arr_relu_13_31 : IN std_logic ;
         d_arr_relu_13_30 : IN std_logic ;
         d_arr_relu_13_29 : IN std_logic ;
         d_arr_relu_13_28 : IN std_logic ;
         d_arr_relu_13_27 : IN std_logic ;
         d_arr_relu_13_26 : IN std_logic ;
         d_arr_relu_13_25 : IN std_logic ;
         d_arr_relu_13_24 : IN std_logic ;
         d_arr_relu_13_23 : IN std_logic ;
         d_arr_relu_13_22 : IN std_logic ;
         d_arr_relu_13_21 : IN std_logic ;
         d_arr_relu_13_20 : IN std_logic ;
         d_arr_relu_13_19 : IN std_logic ;
         d_arr_relu_13_18 : IN std_logic ;
         d_arr_relu_13_17 : IN std_logic ;
         d_arr_relu_13_16 : IN std_logic ;
         d_arr_relu_13_15 : IN std_logic ;
         d_arr_relu_13_14 : IN std_logic ;
         d_arr_relu_13_13 : IN std_logic ;
         d_arr_relu_13_12 : IN std_logic ;
         d_arr_relu_13_11 : IN std_logic ;
         d_arr_relu_13_10 : IN std_logic ;
         d_arr_relu_13_9 : IN std_logic ;
         d_arr_relu_13_8 : IN std_logic ;
         d_arr_relu_13_7 : IN std_logic ;
         d_arr_relu_13_6 : IN std_logic ;
         d_arr_relu_13_5 : IN std_logic ;
         d_arr_relu_13_4 : IN std_logic ;
         d_arr_relu_13_3 : IN std_logic ;
         d_arr_relu_13_2 : IN std_logic ;
         d_arr_relu_13_1 : IN std_logic ;
         d_arr_relu_13_0 : IN std_logic ;
         d_arr_relu_14_31 : IN std_logic ;
         d_arr_relu_14_30 : IN std_logic ;
         d_arr_relu_14_29 : IN std_logic ;
         d_arr_relu_14_28 : IN std_logic ;
         d_arr_relu_14_27 : IN std_logic ;
         d_arr_relu_14_26 : IN std_logic ;
         d_arr_relu_14_25 : IN std_logic ;
         d_arr_relu_14_24 : IN std_logic ;
         d_arr_relu_14_23 : IN std_logic ;
         d_arr_relu_14_22 : IN std_logic ;
         d_arr_relu_14_21 : IN std_logic ;
         d_arr_relu_14_20 : IN std_logic ;
         d_arr_relu_14_19 : IN std_logic ;
         d_arr_relu_14_18 : IN std_logic ;
         d_arr_relu_14_17 : IN std_logic ;
         d_arr_relu_14_16 : IN std_logic ;
         d_arr_relu_14_15 : IN std_logic ;
         d_arr_relu_14_14 : IN std_logic ;
         d_arr_relu_14_13 : IN std_logic ;
         d_arr_relu_14_12 : IN std_logic ;
         d_arr_relu_14_11 : IN std_logic ;
         d_arr_relu_14_10 : IN std_logic ;
         d_arr_relu_14_9 : IN std_logic ;
         d_arr_relu_14_8 : IN std_logic ;
         d_arr_relu_14_7 : IN std_logic ;
         d_arr_relu_14_6 : IN std_logic ;
         d_arr_relu_14_5 : IN std_logic ;
         d_arr_relu_14_4 : IN std_logic ;
         d_arr_relu_14_3 : IN std_logic ;
         d_arr_relu_14_2 : IN std_logic ;
         d_arr_relu_14_1 : IN std_logic ;
         d_arr_relu_14_0 : IN std_logic ;
         d_arr_relu_15_31 : IN std_logic ;
         d_arr_relu_15_30 : IN std_logic ;
         d_arr_relu_15_29 : IN std_logic ;
         d_arr_relu_15_28 : IN std_logic ;
         d_arr_relu_15_27 : IN std_logic ;
         d_arr_relu_15_26 : IN std_logic ;
         d_arr_relu_15_25 : IN std_logic ;
         d_arr_relu_15_24 : IN std_logic ;
         d_arr_relu_15_23 : IN std_logic ;
         d_arr_relu_15_22 : IN std_logic ;
         d_arr_relu_15_21 : IN std_logic ;
         d_arr_relu_15_20 : IN std_logic ;
         d_arr_relu_15_19 : IN std_logic ;
         d_arr_relu_15_18 : IN std_logic ;
         d_arr_relu_15_17 : IN std_logic ;
         d_arr_relu_15_16 : IN std_logic ;
         d_arr_relu_15_15 : IN std_logic ;
         d_arr_relu_15_14 : IN std_logic ;
         d_arr_relu_15_13 : IN std_logic ;
         d_arr_relu_15_12 : IN std_logic ;
         d_arr_relu_15_11 : IN std_logic ;
         d_arr_relu_15_10 : IN std_logic ;
         d_arr_relu_15_9 : IN std_logic ;
         d_arr_relu_15_8 : IN std_logic ;
         d_arr_relu_15_7 : IN std_logic ;
         d_arr_relu_15_6 : IN std_logic ;
         d_arr_relu_15_5 : IN std_logic ;
         d_arr_relu_15_4 : IN std_logic ;
         d_arr_relu_15_3 : IN std_logic ;
         d_arr_relu_15_2 : IN std_logic ;
         d_arr_relu_15_1 : IN std_logic ;
         d_arr_relu_15_0 : IN std_logic ;
         d_arr_relu_16_31 : IN std_logic ;
         d_arr_relu_16_30 : IN std_logic ;
         d_arr_relu_16_29 : IN std_logic ;
         d_arr_relu_16_28 : IN std_logic ;
         d_arr_relu_16_27 : IN std_logic ;
         d_arr_relu_16_26 : IN std_logic ;
         d_arr_relu_16_25 : IN std_logic ;
         d_arr_relu_16_24 : IN std_logic ;
         d_arr_relu_16_23 : IN std_logic ;
         d_arr_relu_16_22 : IN std_logic ;
         d_arr_relu_16_21 : IN std_logic ;
         d_arr_relu_16_20 : IN std_logic ;
         d_arr_relu_16_19 : IN std_logic ;
         d_arr_relu_16_18 : IN std_logic ;
         d_arr_relu_16_17 : IN std_logic ;
         d_arr_relu_16_16 : IN std_logic ;
         d_arr_relu_16_15 : IN std_logic ;
         d_arr_relu_16_14 : IN std_logic ;
         d_arr_relu_16_13 : IN std_logic ;
         d_arr_relu_16_12 : IN std_logic ;
         d_arr_relu_16_11 : IN std_logic ;
         d_arr_relu_16_10 : IN std_logic ;
         d_arr_relu_16_9 : IN std_logic ;
         d_arr_relu_16_8 : IN std_logic ;
         d_arr_relu_16_7 : IN std_logic ;
         d_arr_relu_16_6 : IN std_logic ;
         d_arr_relu_16_5 : IN std_logic ;
         d_arr_relu_16_4 : IN std_logic ;
         d_arr_relu_16_3 : IN std_logic ;
         d_arr_relu_16_2 : IN std_logic ;
         d_arr_relu_16_1 : IN std_logic ;
         d_arr_relu_16_0 : IN std_logic ;
         d_arr_relu_17_31 : IN std_logic ;
         d_arr_relu_17_30 : IN std_logic ;
         d_arr_relu_17_29 : IN std_logic ;
         d_arr_relu_17_28 : IN std_logic ;
         d_arr_relu_17_27 : IN std_logic ;
         d_arr_relu_17_26 : IN std_logic ;
         d_arr_relu_17_25 : IN std_logic ;
         d_arr_relu_17_24 : IN std_logic ;
         d_arr_relu_17_23 : IN std_logic ;
         d_arr_relu_17_22 : IN std_logic ;
         d_arr_relu_17_21 : IN std_logic ;
         d_arr_relu_17_20 : IN std_logic ;
         d_arr_relu_17_19 : IN std_logic ;
         d_arr_relu_17_18 : IN std_logic ;
         d_arr_relu_17_17 : IN std_logic ;
         d_arr_relu_17_16 : IN std_logic ;
         d_arr_relu_17_15 : IN std_logic ;
         d_arr_relu_17_14 : IN std_logic ;
         d_arr_relu_17_13 : IN std_logic ;
         d_arr_relu_17_12 : IN std_logic ;
         d_arr_relu_17_11 : IN std_logic ;
         d_arr_relu_17_10 : IN std_logic ;
         d_arr_relu_17_9 : IN std_logic ;
         d_arr_relu_17_8 : IN std_logic ;
         d_arr_relu_17_7 : IN std_logic ;
         d_arr_relu_17_6 : IN std_logic ;
         d_arr_relu_17_5 : IN std_logic ;
         d_arr_relu_17_4 : IN std_logic ;
         d_arr_relu_17_3 : IN std_logic ;
         d_arr_relu_17_2 : IN std_logic ;
         d_arr_relu_17_1 : IN std_logic ;
         d_arr_relu_17_0 : IN std_logic ;
         d_arr_relu_18_31 : IN std_logic ;
         d_arr_relu_18_30 : IN std_logic ;
         d_arr_relu_18_29 : IN std_logic ;
         d_arr_relu_18_28 : IN std_logic ;
         d_arr_relu_18_27 : IN std_logic ;
         d_arr_relu_18_26 : IN std_logic ;
         d_arr_relu_18_25 : IN std_logic ;
         d_arr_relu_18_24 : IN std_logic ;
         d_arr_relu_18_23 : IN std_logic ;
         d_arr_relu_18_22 : IN std_logic ;
         d_arr_relu_18_21 : IN std_logic ;
         d_arr_relu_18_20 : IN std_logic ;
         d_arr_relu_18_19 : IN std_logic ;
         d_arr_relu_18_18 : IN std_logic ;
         d_arr_relu_18_17 : IN std_logic ;
         d_arr_relu_18_16 : IN std_logic ;
         d_arr_relu_18_15 : IN std_logic ;
         d_arr_relu_18_14 : IN std_logic ;
         d_arr_relu_18_13 : IN std_logic ;
         d_arr_relu_18_12 : IN std_logic ;
         d_arr_relu_18_11 : IN std_logic ;
         d_arr_relu_18_10 : IN std_logic ;
         d_arr_relu_18_9 : IN std_logic ;
         d_arr_relu_18_8 : IN std_logic ;
         d_arr_relu_18_7 : IN std_logic ;
         d_arr_relu_18_6 : IN std_logic ;
         d_arr_relu_18_5 : IN std_logic ;
         d_arr_relu_18_4 : IN std_logic ;
         d_arr_relu_18_3 : IN std_logic ;
         d_arr_relu_18_2 : IN std_logic ;
         d_arr_relu_18_1 : IN std_logic ;
         d_arr_relu_18_0 : IN std_logic ;
         d_arr_relu_19_31 : IN std_logic ;
         d_arr_relu_19_30 : IN std_logic ;
         d_arr_relu_19_29 : IN std_logic ;
         d_arr_relu_19_28 : IN std_logic ;
         d_arr_relu_19_27 : IN std_logic ;
         d_arr_relu_19_26 : IN std_logic ;
         d_arr_relu_19_25 : IN std_logic ;
         d_arr_relu_19_24 : IN std_logic ;
         d_arr_relu_19_23 : IN std_logic ;
         d_arr_relu_19_22 : IN std_logic ;
         d_arr_relu_19_21 : IN std_logic ;
         d_arr_relu_19_20 : IN std_logic ;
         d_arr_relu_19_19 : IN std_logic ;
         d_arr_relu_19_18 : IN std_logic ;
         d_arr_relu_19_17 : IN std_logic ;
         d_arr_relu_19_16 : IN std_logic ;
         d_arr_relu_19_15 : IN std_logic ;
         d_arr_relu_19_14 : IN std_logic ;
         d_arr_relu_19_13 : IN std_logic ;
         d_arr_relu_19_12 : IN std_logic ;
         d_arr_relu_19_11 : IN std_logic ;
         d_arr_relu_19_10 : IN std_logic ;
         d_arr_relu_19_9 : IN std_logic ;
         d_arr_relu_19_8 : IN std_logic ;
         d_arr_relu_19_7 : IN std_logic ;
         d_arr_relu_19_6 : IN std_logic ;
         d_arr_relu_19_5 : IN std_logic ;
         d_arr_relu_19_4 : IN std_logic ;
         d_arr_relu_19_3 : IN std_logic ;
         d_arr_relu_19_2 : IN std_logic ;
         d_arr_relu_19_1 : IN std_logic ;
         d_arr_relu_19_0 : IN std_logic ;
         d_arr_relu_20_31 : IN std_logic ;
         d_arr_relu_20_30 : IN std_logic ;
         d_arr_relu_20_29 : IN std_logic ;
         d_arr_relu_20_28 : IN std_logic ;
         d_arr_relu_20_27 : IN std_logic ;
         d_arr_relu_20_26 : IN std_logic ;
         d_arr_relu_20_25 : IN std_logic ;
         d_arr_relu_20_24 : IN std_logic ;
         d_arr_relu_20_23 : IN std_logic ;
         d_arr_relu_20_22 : IN std_logic ;
         d_arr_relu_20_21 : IN std_logic ;
         d_arr_relu_20_20 : IN std_logic ;
         d_arr_relu_20_19 : IN std_logic ;
         d_arr_relu_20_18 : IN std_logic ;
         d_arr_relu_20_17 : IN std_logic ;
         d_arr_relu_20_16 : IN std_logic ;
         d_arr_relu_20_15 : IN std_logic ;
         d_arr_relu_20_14 : IN std_logic ;
         d_arr_relu_20_13 : IN std_logic ;
         d_arr_relu_20_12 : IN std_logic ;
         d_arr_relu_20_11 : IN std_logic ;
         d_arr_relu_20_10 : IN std_logic ;
         d_arr_relu_20_9 : IN std_logic ;
         d_arr_relu_20_8 : IN std_logic ;
         d_arr_relu_20_7 : IN std_logic ;
         d_arr_relu_20_6 : IN std_logic ;
         d_arr_relu_20_5 : IN std_logic ;
         d_arr_relu_20_4 : IN std_logic ;
         d_arr_relu_20_3 : IN std_logic ;
         d_arr_relu_20_2 : IN std_logic ;
         d_arr_relu_20_1 : IN std_logic ;
         d_arr_relu_20_0 : IN std_logic ;
         d_arr_relu_21_31 : IN std_logic ;
         d_arr_relu_21_30 : IN std_logic ;
         d_arr_relu_21_29 : IN std_logic ;
         d_arr_relu_21_28 : IN std_logic ;
         d_arr_relu_21_27 : IN std_logic ;
         d_arr_relu_21_26 : IN std_logic ;
         d_arr_relu_21_25 : IN std_logic ;
         d_arr_relu_21_24 : IN std_logic ;
         d_arr_relu_21_23 : IN std_logic ;
         d_arr_relu_21_22 : IN std_logic ;
         d_arr_relu_21_21 : IN std_logic ;
         d_arr_relu_21_20 : IN std_logic ;
         d_arr_relu_21_19 : IN std_logic ;
         d_arr_relu_21_18 : IN std_logic ;
         d_arr_relu_21_17 : IN std_logic ;
         d_arr_relu_21_16 : IN std_logic ;
         d_arr_relu_21_15 : IN std_logic ;
         d_arr_relu_21_14 : IN std_logic ;
         d_arr_relu_21_13 : IN std_logic ;
         d_arr_relu_21_12 : IN std_logic ;
         d_arr_relu_21_11 : IN std_logic ;
         d_arr_relu_21_10 : IN std_logic ;
         d_arr_relu_21_9 : IN std_logic ;
         d_arr_relu_21_8 : IN std_logic ;
         d_arr_relu_21_7 : IN std_logic ;
         d_arr_relu_21_6 : IN std_logic ;
         d_arr_relu_21_5 : IN std_logic ;
         d_arr_relu_21_4 : IN std_logic ;
         d_arr_relu_21_3 : IN std_logic ;
         d_arr_relu_21_2 : IN std_logic ;
         d_arr_relu_21_1 : IN std_logic ;
         d_arr_relu_21_0 : IN std_logic ;
         d_arr_relu_22_31 : IN std_logic ;
         d_arr_relu_22_30 : IN std_logic ;
         d_arr_relu_22_29 : IN std_logic ;
         d_arr_relu_22_28 : IN std_logic ;
         d_arr_relu_22_27 : IN std_logic ;
         d_arr_relu_22_26 : IN std_logic ;
         d_arr_relu_22_25 : IN std_logic ;
         d_arr_relu_22_24 : IN std_logic ;
         d_arr_relu_22_23 : IN std_logic ;
         d_arr_relu_22_22 : IN std_logic ;
         d_arr_relu_22_21 : IN std_logic ;
         d_arr_relu_22_20 : IN std_logic ;
         d_arr_relu_22_19 : IN std_logic ;
         d_arr_relu_22_18 : IN std_logic ;
         d_arr_relu_22_17 : IN std_logic ;
         d_arr_relu_22_16 : IN std_logic ;
         d_arr_relu_22_15 : IN std_logic ;
         d_arr_relu_22_14 : IN std_logic ;
         d_arr_relu_22_13 : IN std_logic ;
         d_arr_relu_22_12 : IN std_logic ;
         d_arr_relu_22_11 : IN std_logic ;
         d_arr_relu_22_10 : IN std_logic ;
         d_arr_relu_22_9 : IN std_logic ;
         d_arr_relu_22_8 : IN std_logic ;
         d_arr_relu_22_7 : IN std_logic ;
         d_arr_relu_22_6 : IN std_logic ;
         d_arr_relu_22_5 : IN std_logic ;
         d_arr_relu_22_4 : IN std_logic ;
         d_arr_relu_22_3 : IN std_logic ;
         d_arr_relu_22_2 : IN std_logic ;
         d_arr_relu_22_1 : IN std_logic ;
         d_arr_relu_22_0 : IN std_logic ;
         d_arr_relu_23_31 : IN std_logic ;
         d_arr_relu_23_30 : IN std_logic ;
         d_arr_relu_23_29 : IN std_logic ;
         d_arr_relu_23_28 : IN std_logic ;
         d_arr_relu_23_27 : IN std_logic ;
         d_arr_relu_23_26 : IN std_logic ;
         d_arr_relu_23_25 : IN std_logic ;
         d_arr_relu_23_24 : IN std_logic ;
         d_arr_relu_23_23 : IN std_logic ;
         d_arr_relu_23_22 : IN std_logic ;
         d_arr_relu_23_21 : IN std_logic ;
         d_arr_relu_23_20 : IN std_logic ;
         d_arr_relu_23_19 : IN std_logic ;
         d_arr_relu_23_18 : IN std_logic ;
         d_arr_relu_23_17 : IN std_logic ;
         d_arr_relu_23_16 : IN std_logic ;
         d_arr_relu_23_15 : IN std_logic ;
         d_arr_relu_23_14 : IN std_logic ;
         d_arr_relu_23_13 : IN std_logic ;
         d_arr_relu_23_12 : IN std_logic ;
         d_arr_relu_23_11 : IN std_logic ;
         d_arr_relu_23_10 : IN std_logic ;
         d_arr_relu_23_9 : IN std_logic ;
         d_arr_relu_23_8 : IN std_logic ;
         d_arr_relu_23_7 : IN std_logic ;
         d_arr_relu_23_6 : IN std_logic ;
         d_arr_relu_23_5 : IN std_logic ;
         d_arr_relu_23_4 : IN std_logic ;
         d_arr_relu_23_3 : IN std_logic ;
         d_arr_relu_23_2 : IN std_logic ;
         d_arr_relu_23_1 : IN std_logic ;
         d_arr_relu_23_0 : IN std_logic ;
         d_arr_relu_24_31 : IN std_logic ;
         d_arr_relu_24_30 : IN std_logic ;
         d_arr_relu_24_29 : IN std_logic ;
         d_arr_relu_24_28 : IN std_logic ;
         d_arr_relu_24_27 : IN std_logic ;
         d_arr_relu_24_26 : IN std_logic ;
         d_arr_relu_24_25 : IN std_logic ;
         d_arr_relu_24_24 : IN std_logic ;
         d_arr_relu_24_23 : IN std_logic ;
         d_arr_relu_24_22 : IN std_logic ;
         d_arr_relu_24_21 : IN std_logic ;
         d_arr_relu_24_20 : IN std_logic ;
         d_arr_relu_24_19 : IN std_logic ;
         d_arr_relu_24_18 : IN std_logic ;
         d_arr_relu_24_17 : IN std_logic ;
         d_arr_relu_24_16 : IN std_logic ;
         d_arr_relu_24_15 : IN std_logic ;
         d_arr_relu_24_14 : IN std_logic ;
         d_arr_relu_24_13 : IN std_logic ;
         d_arr_relu_24_12 : IN std_logic ;
         d_arr_relu_24_11 : IN std_logic ;
         d_arr_relu_24_10 : IN std_logic ;
         d_arr_relu_24_9 : IN std_logic ;
         d_arr_relu_24_8 : IN std_logic ;
         d_arr_relu_24_7 : IN std_logic ;
         d_arr_relu_24_6 : IN std_logic ;
         d_arr_relu_24_5 : IN std_logic ;
         d_arr_relu_24_4 : IN std_logic ;
         d_arr_relu_24_3 : IN std_logic ;
         d_arr_relu_24_2 : IN std_logic ;
         d_arr_relu_24_1 : IN std_logic ;
         d_arr_relu_24_0 : IN std_logic ;
         sel_mux : IN std_logic ;
         sel_mul : IN std_logic ;
         sel_add : IN std_logic ;
         sel_merge1 : IN std_logic ;
         sel_merge2 : IN std_logic ;
         sel_relu : IN std_logic ;
         d_arr_0_31 : OUT std_logic ;
         d_arr_0_30 : OUT std_logic ;
         d_arr_0_29 : OUT std_logic ;
         d_arr_0_28 : OUT std_logic ;
         d_arr_0_27 : OUT std_logic ;
         d_arr_0_26 : OUT std_logic ;
         d_arr_0_25 : OUT std_logic ;
         d_arr_0_24 : OUT std_logic ;
         d_arr_0_23 : OUT std_logic ;
         d_arr_0_22 : OUT std_logic ;
         d_arr_0_21 : OUT std_logic ;
         d_arr_0_20 : OUT std_logic ;
         d_arr_0_19 : OUT std_logic ;
         d_arr_0_18 : OUT std_logic ;
         d_arr_0_17 : OUT std_logic ;
         d_arr_0_16 : OUT std_logic ;
         d_arr_0_15 : OUT std_logic ;
         d_arr_0_14 : OUT std_logic ;
         d_arr_0_13 : OUT std_logic ;
         d_arr_0_12 : OUT std_logic ;
         d_arr_0_11 : OUT std_logic ;
         d_arr_0_10 : OUT std_logic ;
         d_arr_0_9 : OUT std_logic ;
         d_arr_0_8 : OUT std_logic ;
         d_arr_0_7 : OUT std_logic ;
         d_arr_0_6 : OUT std_logic ;
         d_arr_0_5 : OUT std_logic ;
         d_arr_0_4 : OUT std_logic ;
         d_arr_0_3 : OUT std_logic ;
         d_arr_0_2 : OUT std_logic ;
         d_arr_0_1 : OUT std_logic ;
         d_arr_0_0 : OUT std_logic ;
         d_arr_1_31 : OUT std_logic ;
         d_arr_1_30 : OUT std_logic ;
         d_arr_1_29 : OUT std_logic ;
         d_arr_1_28 : OUT std_logic ;
         d_arr_1_27 : OUT std_logic ;
         d_arr_1_26 : OUT std_logic ;
         d_arr_1_25 : OUT std_logic ;
         d_arr_1_24 : OUT std_logic ;
         d_arr_1_23 : OUT std_logic ;
         d_arr_1_22 : OUT std_logic ;
         d_arr_1_21 : OUT std_logic ;
         d_arr_1_20 : OUT std_logic ;
         d_arr_1_19 : OUT std_logic ;
         d_arr_1_18 : OUT std_logic ;
         d_arr_1_17 : OUT std_logic ;
         d_arr_1_16 : OUT std_logic ;
         d_arr_1_15 : OUT std_logic ;
         d_arr_1_14 : OUT std_logic ;
         d_arr_1_13 : OUT std_logic ;
         d_arr_1_12 : OUT std_logic ;
         d_arr_1_11 : OUT std_logic ;
         d_arr_1_10 : OUT std_logic ;
         d_arr_1_9 : OUT std_logic ;
         d_arr_1_8 : OUT std_logic ;
         d_arr_1_7 : OUT std_logic ;
         d_arr_1_6 : OUT std_logic ;
         d_arr_1_5 : OUT std_logic ;
         d_arr_1_4 : OUT std_logic ;
         d_arr_1_3 : OUT std_logic ;
         d_arr_1_2 : OUT std_logic ;
         d_arr_1_1 : OUT std_logic ;
         d_arr_1_0 : OUT std_logic ;
         d_arr_2_31 : OUT std_logic ;
         d_arr_2_30 : OUT std_logic ;
         d_arr_2_29 : OUT std_logic ;
         d_arr_2_28 : OUT std_logic ;
         d_arr_2_27 : OUT std_logic ;
         d_arr_2_26 : OUT std_logic ;
         d_arr_2_25 : OUT std_logic ;
         d_arr_2_24 : OUT std_logic ;
         d_arr_2_23 : OUT std_logic ;
         d_arr_2_22 : OUT std_logic ;
         d_arr_2_21 : OUT std_logic ;
         d_arr_2_20 : OUT std_logic ;
         d_arr_2_19 : OUT std_logic ;
         d_arr_2_18 : OUT std_logic ;
         d_arr_2_17 : OUT std_logic ;
         d_arr_2_16 : OUT std_logic ;
         d_arr_2_15 : OUT std_logic ;
         d_arr_2_14 : OUT std_logic ;
         d_arr_2_13 : OUT std_logic ;
         d_arr_2_12 : OUT std_logic ;
         d_arr_2_11 : OUT std_logic ;
         d_arr_2_10 : OUT std_logic ;
         d_arr_2_9 : OUT std_logic ;
         d_arr_2_8 : OUT std_logic ;
         d_arr_2_7 : OUT std_logic ;
         d_arr_2_6 : OUT std_logic ;
         d_arr_2_5 : OUT std_logic ;
         d_arr_2_4 : OUT std_logic ;
         d_arr_2_3 : OUT std_logic ;
         d_arr_2_2 : OUT std_logic ;
         d_arr_2_1 : OUT std_logic ;
         d_arr_2_0 : OUT std_logic ;
         d_arr_3_31 : OUT std_logic ;
         d_arr_3_30 : OUT std_logic ;
         d_arr_3_29 : OUT std_logic ;
         d_arr_3_28 : OUT std_logic ;
         d_arr_3_27 : OUT std_logic ;
         d_arr_3_26 : OUT std_logic ;
         d_arr_3_25 : OUT std_logic ;
         d_arr_3_24 : OUT std_logic ;
         d_arr_3_23 : OUT std_logic ;
         d_arr_3_22 : OUT std_logic ;
         d_arr_3_21 : OUT std_logic ;
         d_arr_3_20 : OUT std_logic ;
         d_arr_3_19 : OUT std_logic ;
         d_arr_3_18 : OUT std_logic ;
         d_arr_3_17 : OUT std_logic ;
         d_arr_3_16 : OUT std_logic ;
         d_arr_3_15 : OUT std_logic ;
         d_arr_3_14 : OUT std_logic ;
         d_arr_3_13 : OUT std_logic ;
         d_arr_3_12 : OUT std_logic ;
         d_arr_3_11 : OUT std_logic ;
         d_arr_3_10 : OUT std_logic ;
         d_arr_3_9 : OUT std_logic ;
         d_arr_3_8 : OUT std_logic ;
         d_arr_3_7 : OUT std_logic ;
         d_arr_3_6 : OUT std_logic ;
         d_arr_3_5 : OUT std_logic ;
         d_arr_3_4 : OUT std_logic ;
         d_arr_3_3 : OUT std_logic ;
         d_arr_3_2 : OUT std_logic ;
         d_arr_3_1 : OUT std_logic ;
         d_arr_3_0 : OUT std_logic ;
         d_arr_4_31 : OUT std_logic ;
         d_arr_4_30 : OUT std_logic ;
         d_arr_4_29 : OUT std_logic ;
         d_arr_4_28 : OUT std_logic ;
         d_arr_4_27 : OUT std_logic ;
         d_arr_4_26 : OUT std_logic ;
         d_arr_4_25 : OUT std_logic ;
         d_arr_4_24 : OUT std_logic ;
         d_arr_4_23 : OUT std_logic ;
         d_arr_4_22 : OUT std_logic ;
         d_arr_4_21 : OUT std_logic ;
         d_arr_4_20 : OUT std_logic ;
         d_arr_4_19 : OUT std_logic ;
         d_arr_4_18 : OUT std_logic ;
         d_arr_4_17 : OUT std_logic ;
         d_arr_4_16 : OUT std_logic ;
         d_arr_4_15 : OUT std_logic ;
         d_arr_4_14 : OUT std_logic ;
         d_arr_4_13 : OUT std_logic ;
         d_arr_4_12 : OUT std_logic ;
         d_arr_4_11 : OUT std_logic ;
         d_arr_4_10 : OUT std_logic ;
         d_arr_4_9 : OUT std_logic ;
         d_arr_4_8 : OUT std_logic ;
         d_arr_4_7 : OUT std_logic ;
         d_arr_4_6 : OUT std_logic ;
         d_arr_4_5 : OUT std_logic ;
         d_arr_4_4 : OUT std_logic ;
         d_arr_4_3 : OUT std_logic ;
         d_arr_4_2 : OUT std_logic ;
         d_arr_4_1 : OUT std_logic ;
         d_arr_4_0 : OUT std_logic ;
         d_arr_5_31 : OUT std_logic ;
         d_arr_5_30 : OUT std_logic ;
         d_arr_5_29 : OUT std_logic ;
         d_arr_5_28 : OUT std_logic ;
         d_arr_5_27 : OUT std_logic ;
         d_arr_5_26 : OUT std_logic ;
         d_arr_5_25 : OUT std_logic ;
         d_arr_5_24 : OUT std_logic ;
         d_arr_5_23 : OUT std_logic ;
         d_arr_5_22 : OUT std_logic ;
         d_arr_5_21 : OUT std_logic ;
         d_arr_5_20 : OUT std_logic ;
         d_arr_5_19 : OUT std_logic ;
         d_arr_5_18 : OUT std_logic ;
         d_arr_5_17 : OUT std_logic ;
         d_arr_5_16 : OUT std_logic ;
         d_arr_5_15 : OUT std_logic ;
         d_arr_5_14 : OUT std_logic ;
         d_arr_5_13 : OUT std_logic ;
         d_arr_5_12 : OUT std_logic ;
         d_arr_5_11 : OUT std_logic ;
         d_arr_5_10 : OUT std_logic ;
         d_arr_5_9 : OUT std_logic ;
         d_arr_5_8 : OUT std_logic ;
         d_arr_5_7 : OUT std_logic ;
         d_arr_5_6 : OUT std_logic ;
         d_arr_5_5 : OUT std_logic ;
         d_arr_5_4 : OUT std_logic ;
         d_arr_5_3 : OUT std_logic ;
         d_arr_5_2 : OUT std_logic ;
         d_arr_5_1 : OUT std_logic ;
         d_arr_5_0 : OUT std_logic ;
         d_arr_6_31 : OUT std_logic ;
         d_arr_6_30 : OUT std_logic ;
         d_arr_6_29 : OUT std_logic ;
         d_arr_6_28 : OUT std_logic ;
         d_arr_6_27 : OUT std_logic ;
         d_arr_6_26 : OUT std_logic ;
         d_arr_6_25 : OUT std_logic ;
         d_arr_6_24 : OUT std_logic ;
         d_arr_6_23 : OUT std_logic ;
         d_arr_6_22 : OUT std_logic ;
         d_arr_6_21 : OUT std_logic ;
         d_arr_6_20 : OUT std_logic ;
         d_arr_6_19 : OUT std_logic ;
         d_arr_6_18 : OUT std_logic ;
         d_arr_6_17 : OUT std_logic ;
         d_arr_6_16 : OUT std_logic ;
         d_arr_6_15 : OUT std_logic ;
         d_arr_6_14 : OUT std_logic ;
         d_arr_6_13 : OUT std_logic ;
         d_arr_6_12 : OUT std_logic ;
         d_arr_6_11 : OUT std_logic ;
         d_arr_6_10 : OUT std_logic ;
         d_arr_6_9 : OUT std_logic ;
         d_arr_6_8 : OUT std_logic ;
         d_arr_6_7 : OUT std_logic ;
         d_arr_6_6 : OUT std_logic ;
         d_arr_6_5 : OUT std_logic ;
         d_arr_6_4 : OUT std_logic ;
         d_arr_6_3 : OUT std_logic ;
         d_arr_6_2 : OUT std_logic ;
         d_arr_6_1 : OUT std_logic ;
         d_arr_6_0 : OUT std_logic ;
         d_arr_7_31 : OUT std_logic ;
         d_arr_7_30 : OUT std_logic ;
         d_arr_7_29 : OUT std_logic ;
         d_arr_7_28 : OUT std_logic ;
         d_arr_7_27 : OUT std_logic ;
         d_arr_7_26 : OUT std_logic ;
         d_arr_7_25 : OUT std_logic ;
         d_arr_7_24 : OUT std_logic ;
         d_arr_7_23 : OUT std_logic ;
         d_arr_7_22 : OUT std_logic ;
         d_arr_7_21 : OUT std_logic ;
         d_arr_7_20 : OUT std_logic ;
         d_arr_7_19 : OUT std_logic ;
         d_arr_7_18 : OUT std_logic ;
         d_arr_7_17 : OUT std_logic ;
         d_arr_7_16 : OUT std_logic ;
         d_arr_7_15 : OUT std_logic ;
         d_arr_7_14 : OUT std_logic ;
         d_arr_7_13 : OUT std_logic ;
         d_arr_7_12 : OUT std_logic ;
         d_arr_7_11 : OUT std_logic ;
         d_arr_7_10 : OUT std_logic ;
         d_arr_7_9 : OUT std_logic ;
         d_arr_7_8 : OUT std_logic ;
         d_arr_7_7 : OUT std_logic ;
         d_arr_7_6 : OUT std_logic ;
         d_arr_7_5 : OUT std_logic ;
         d_arr_7_4 : OUT std_logic ;
         d_arr_7_3 : OUT std_logic ;
         d_arr_7_2 : OUT std_logic ;
         d_arr_7_1 : OUT std_logic ;
         d_arr_7_0 : OUT std_logic ;
         d_arr_8_31 : OUT std_logic ;
         d_arr_8_30 : OUT std_logic ;
         d_arr_8_29 : OUT std_logic ;
         d_arr_8_28 : OUT std_logic ;
         d_arr_8_27 : OUT std_logic ;
         d_arr_8_26 : OUT std_logic ;
         d_arr_8_25 : OUT std_logic ;
         d_arr_8_24 : OUT std_logic ;
         d_arr_8_23 : OUT std_logic ;
         d_arr_8_22 : OUT std_logic ;
         d_arr_8_21 : OUT std_logic ;
         d_arr_8_20 : OUT std_logic ;
         d_arr_8_19 : OUT std_logic ;
         d_arr_8_18 : OUT std_logic ;
         d_arr_8_17 : OUT std_logic ;
         d_arr_8_16 : OUT std_logic ;
         d_arr_8_15 : OUT std_logic ;
         d_arr_8_14 : OUT std_logic ;
         d_arr_8_13 : OUT std_logic ;
         d_arr_8_12 : OUT std_logic ;
         d_arr_8_11 : OUT std_logic ;
         d_arr_8_10 : OUT std_logic ;
         d_arr_8_9 : OUT std_logic ;
         d_arr_8_8 : OUT std_logic ;
         d_arr_8_7 : OUT std_logic ;
         d_arr_8_6 : OUT std_logic ;
         d_arr_8_5 : OUT std_logic ;
         d_arr_8_4 : OUT std_logic ;
         d_arr_8_3 : OUT std_logic ;
         d_arr_8_2 : OUT std_logic ;
         d_arr_8_1 : OUT std_logic ;
         d_arr_8_0 : OUT std_logic ;
         d_arr_9_31 : OUT std_logic ;
         d_arr_9_30 : OUT std_logic ;
         d_arr_9_29 : OUT std_logic ;
         d_arr_9_28 : OUT std_logic ;
         d_arr_9_27 : OUT std_logic ;
         d_arr_9_26 : OUT std_logic ;
         d_arr_9_25 : OUT std_logic ;
         d_arr_9_24 : OUT std_logic ;
         d_arr_9_23 : OUT std_logic ;
         d_arr_9_22 : OUT std_logic ;
         d_arr_9_21 : OUT std_logic ;
         d_arr_9_20 : OUT std_logic ;
         d_arr_9_19 : OUT std_logic ;
         d_arr_9_18 : OUT std_logic ;
         d_arr_9_17 : OUT std_logic ;
         d_arr_9_16 : OUT std_logic ;
         d_arr_9_15 : OUT std_logic ;
         d_arr_9_14 : OUT std_logic ;
         d_arr_9_13 : OUT std_logic ;
         d_arr_9_12 : OUT std_logic ;
         d_arr_9_11 : OUT std_logic ;
         d_arr_9_10 : OUT std_logic ;
         d_arr_9_9 : OUT std_logic ;
         d_arr_9_8 : OUT std_logic ;
         d_arr_9_7 : OUT std_logic ;
         d_arr_9_6 : OUT std_logic ;
         d_arr_9_5 : OUT std_logic ;
         d_arr_9_4 : OUT std_logic ;
         d_arr_9_3 : OUT std_logic ;
         d_arr_9_2 : OUT std_logic ;
         d_arr_9_1 : OUT std_logic ;
         d_arr_9_0 : OUT std_logic ;
         d_arr_10_31 : OUT std_logic ;
         d_arr_10_30 : OUT std_logic ;
         d_arr_10_29 : OUT std_logic ;
         d_arr_10_28 : OUT std_logic ;
         d_arr_10_27 : OUT std_logic ;
         d_arr_10_26 : OUT std_logic ;
         d_arr_10_25 : OUT std_logic ;
         d_arr_10_24 : OUT std_logic ;
         d_arr_10_23 : OUT std_logic ;
         d_arr_10_22 : OUT std_logic ;
         d_arr_10_21 : OUT std_logic ;
         d_arr_10_20 : OUT std_logic ;
         d_arr_10_19 : OUT std_logic ;
         d_arr_10_18 : OUT std_logic ;
         d_arr_10_17 : OUT std_logic ;
         d_arr_10_16 : OUT std_logic ;
         d_arr_10_15 : OUT std_logic ;
         d_arr_10_14 : OUT std_logic ;
         d_arr_10_13 : OUT std_logic ;
         d_arr_10_12 : OUT std_logic ;
         d_arr_10_11 : OUT std_logic ;
         d_arr_10_10 : OUT std_logic ;
         d_arr_10_9 : OUT std_logic ;
         d_arr_10_8 : OUT std_logic ;
         d_arr_10_7 : OUT std_logic ;
         d_arr_10_6 : OUT std_logic ;
         d_arr_10_5 : OUT std_logic ;
         d_arr_10_4 : OUT std_logic ;
         d_arr_10_3 : OUT std_logic ;
         d_arr_10_2 : OUT std_logic ;
         d_arr_10_1 : OUT std_logic ;
         d_arr_10_0 : OUT std_logic ;
         d_arr_11_31 : OUT std_logic ;
         d_arr_11_30 : OUT std_logic ;
         d_arr_11_29 : OUT std_logic ;
         d_arr_11_28 : OUT std_logic ;
         d_arr_11_27 : OUT std_logic ;
         d_arr_11_26 : OUT std_logic ;
         d_arr_11_25 : OUT std_logic ;
         d_arr_11_24 : OUT std_logic ;
         d_arr_11_23 : OUT std_logic ;
         d_arr_11_22 : OUT std_logic ;
         d_arr_11_21 : OUT std_logic ;
         d_arr_11_20 : OUT std_logic ;
         d_arr_11_19 : OUT std_logic ;
         d_arr_11_18 : OUT std_logic ;
         d_arr_11_17 : OUT std_logic ;
         d_arr_11_16 : OUT std_logic ;
         d_arr_11_15 : OUT std_logic ;
         d_arr_11_14 : OUT std_logic ;
         d_arr_11_13 : OUT std_logic ;
         d_arr_11_12 : OUT std_logic ;
         d_arr_11_11 : OUT std_logic ;
         d_arr_11_10 : OUT std_logic ;
         d_arr_11_9 : OUT std_logic ;
         d_arr_11_8 : OUT std_logic ;
         d_arr_11_7 : OUT std_logic ;
         d_arr_11_6 : OUT std_logic ;
         d_arr_11_5 : OUT std_logic ;
         d_arr_11_4 : OUT std_logic ;
         d_arr_11_3 : OUT std_logic ;
         d_arr_11_2 : OUT std_logic ;
         d_arr_11_1 : OUT std_logic ;
         d_arr_11_0 : OUT std_logic ;
         d_arr_12_31 : OUT std_logic ;
         d_arr_12_30 : OUT std_logic ;
         d_arr_12_29 : OUT std_logic ;
         d_arr_12_28 : OUT std_logic ;
         d_arr_12_27 : OUT std_logic ;
         d_arr_12_26 : OUT std_logic ;
         d_arr_12_25 : OUT std_logic ;
         d_arr_12_24 : OUT std_logic ;
         d_arr_12_23 : OUT std_logic ;
         d_arr_12_22 : OUT std_logic ;
         d_arr_12_21 : OUT std_logic ;
         d_arr_12_20 : OUT std_logic ;
         d_arr_12_19 : OUT std_logic ;
         d_arr_12_18 : OUT std_logic ;
         d_arr_12_17 : OUT std_logic ;
         d_arr_12_16 : OUT std_logic ;
         d_arr_12_15 : OUT std_logic ;
         d_arr_12_14 : OUT std_logic ;
         d_arr_12_13 : OUT std_logic ;
         d_arr_12_12 : OUT std_logic ;
         d_arr_12_11 : OUT std_logic ;
         d_arr_12_10 : OUT std_logic ;
         d_arr_12_9 : OUT std_logic ;
         d_arr_12_8 : OUT std_logic ;
         d_arr_12_7 : OUT std_logic ;
         d_arr_12_6 : OUT std_logic ;
         d_arr_12_5 : OUT std_logic ;
         d_arr_12_4 : OUT std_logic ;
         d_arr_12_3 : OUT std_logic ;
         d_arr_12_2 : OUT std_logic ;
         d_arr_12_1 : OUT std_logic ;
         d_arr_12_0 : OUT std_logic ;
         d_arr_13_31 : OUT std_logic ;
         d_arr_13_30 : OUT std_logic ;
         d_arr_13_29 : OUT std_logic ;
         d_arr_13_28 : OUT std_logic ;
         d_arr_13_27 : OUT std_logic ;
         d_arr_13_26 : OUT std_logic ;
         d_arr_13_25 : OUT std_logic ;
         d_arr_13_24 : OUT std_logic ;
         d_arr_13_23 : OUT std_logic ;
         d_arr_13_22 : OUT std_logic ;
         d_arr_13_21 : OUT std_logic ;
         d_arr_13_20 : OUT std_logic ;
         d_arr_13_19 : OUT std_logic ;
         d_arr_13_18 : OUT std_logic ;
         d_arr_13_17 : OUT std_logic ;
         d_arr_13_16 : OUT std_logic ;
         d_arr_13_15 : OUT std_logic ;
         d_arr_13_14 : OUT std_logic ;
         d_arr_13_13 : OUT std_logic ;
         d_arr_13_12 : OUT std_logic ;
         d_arr_13_11 : OUT std_logic ;
         d_arr_13_10 : OUT std_logic ;
         d_arr_13_9 : OUT std_logic ;
         d_arr_13_8 : OUT std_logic ;
         d_arr_13_7 : OUT std_logic ;
         d_arr_13_6 : OUT std_logic ;
         d_arr_13_5 : OUT std_logic ;
         d_arr_13_4 : OUT std_logic ;
         d_arr_13_3 : OUT std_logic ;
         d_arr_13_2 : OUT std_logic ;
         d_arr_13_1 : OUT std_logic ;
         d_arr_13_0 : OUT std_logic ;
         d_arr_14_31 : OUT std_logic ;
         d_arr_14_30 : OUT std_logic ;
         d_arr_14_29 : OUT std_logic ;
         d_arr_14_28 : OUT std_logic ;
         d_arr_14_27 : OUT std_logic ;
         d_arr_14_26 : OUT std_logic ;
         d_arr_14_25 : OUT std_logic ;
         d_arr_14_24 : OUT std_logic ;
         d_arr_14_23 : OUT std_logic ;
         d_arr_14_22 : OUT std_logic ;
         d_arr_14_21 : OUT std_logic ;
         d_arr_14_20 : OUT std_logic ;
         d_arr_14_19 : OUT std_logic ;
         d_arr_14_18 : OUT std_logic ;
         d_arr_14_17 : OUT std_logic ;
         d_arr_14_16 : OUT std_logic ;
         d_arr_14_15 : OUT std_logic ;
         d_arr_14_14 : OUT std_logic ;
         d_arr_14_13 : OUT std_logic ;
         d_arr_14_12 : OUT std_logic ;
         d_arr_14_11 : OUT std_logic ;
         d_arr_14_10 : OUT std_logic ;
         d_arr_14_9 : OUT std_logic ;
         d_arr_14_8 : OUT std_logic ;
         d_arr_14_7 : OUT std_logic ;
         d_arr_14_6 : OUT std_logic ;
         d_arr_14_5 : OUT std_logic ;
         d_arr_14_4 : OUT std_logic ;
         d_arr_14_3 : OUT std_logic ;
         d_arr_14_2 : OUT std_logic ;
         d_arr_14_1 : OUT std_logic ;
         d_arr_14_0 : OUT std_logic ;
         d_arr_15_31 : OUT std_logic ;
         d_arr_15_30 : OUT std_logic ;
         d_arr_15_29 : OUT std_logic ;
         d_arr_15_28 : OUT std_logic ;
         d_arr_15_27 : OUT std_logic ;
         d_arr_15_26 : OUT std_logic ;
         d_arr_15_25 : OUT std_logic ;
         d_arr_15_24 : OUT std_logic ;
         d_arr_15_23 : OUT std_logic ;
         d_arr_15_22 : OUT std_logic ;
         d_arr_15_21 : OUT std_logic ;
         d_arr_15_20 : OUT std_logic ;
         d_arr_15_19 : OUT std_logic ;
         d_arr_15_18 : OUT std_logic ;
         d_arr_15_17 : OUT std_logic ;
         d_arr_15_16 : OUT std_logic ;
         d_arr_15_15 : OUT std_logic ;
         d_arr_15_14 : OUT std_logic ;
         d_arr_15_13 : OUT std_logic ;
         d_arr_15_12 : OUT std_logic ;
         d_arr_15_11 : OUT std_logic ;
         d_arr_15_10 : OUT std_logic ;
         d_arr_15_9 : OUT std_logic ;
         d_arr_15_8 : OUT std_logic ;
         d_arr_15_7 : OUT std_logic ;
         d_arr_15_6 : OUT std_logic ;
         d_arr_15_5 : OUT std_logic ;
         d_arr_15_4 : OUT std_logic ;
         d_arr_15_3 : OUT std_logic ;
         d_arr_15_2 : OUT std_logic ;
         d_arr_15_1 : OUT std_logic ;
         d_arr_15_0 : OUT std_logic ;
         d_arr_16_31 : OUT std_logic ;
         d_arr_16_30 : OUT std_logic ;
         d_arr_16_29 : OUT std_logic ;
         d_arr_16_28 : OUT std_logic ;
         d_arr_16_27 : OUT std_logic ;
         d_arr_16_26 : OUT std_logic ;
         d_arr_16_25 : OUT std_logic ;
         d_arr_16_24 : OUT std_logic ;
         d_arr_16_23 : OUT std_logic ;
         d_arr_16_22 : OUT std_logic ;
         d_arr_16_21 : OUT std_logic ;
         d_arr_16_20 : OUT std_logic ;
         d_arr_16_19 : OUT std_logic ;
         d_arr_16_18 : OUT std_logic ;
         d_arr_16_17 : OUT std_logic ;
         d_arr_16_16 : OUT std_logic ;
         d_arr_16_15 : OUT std_logic ;
         d_arr_16_14 : OUT std_logic ;
         d_arr_16_13 : OUT std_logic ;
         d_arr_16_12 : OUT std_logic ;
         d_arr_16_11 : OUT std_logic ;
         d_arr_16_10 : OUT std_logic ;
         d_arr_16_9 : OUT std_logic ;
         d_arr_16_8 : OUT std_logic ;
         d_arr_16_7 : OUT std_logic ;
         d_arr_16_6 : OUT std_logic ;
         d_arr_16_5 : OUT std_logic ;
         d_arr_16_4 : OUT std_logic ;
         d_arr_16_3 : OUT std_logic ;
         d_arr_16_2 : OUT std_logic ;
         d_arr_16_1 : OUT std_logic ;
         d_arr_16_0 : OUT std_logic ;
         d_arr_17_31 : OUT std_logic ;
         d_arr_17_30 : OUT std_logic ;
         d_arr_17_29 : OUT std_logic ;
         d_arr_17_28 : OUT std_logic ;
         d_arr_17_27 : OUT std_logic ;
         d_arr_17_26 : OUT std_logic ;
         d_arr_17_25 : OUT std_logic ;
         d_arr_17_24 : OUT std_logic ;
         d_arr_17_23 : OUT std_logic ;
         d_arr_17_22 : OUT std_logic ;
         d_arr_17_21 : OUT std_logic ;
         d_arr_17_20 : OUT std_logic ;
         d_arr_17_19 : OUT std_logic ;
         d_arr_17_18 : OUT std_logic ;
         d_arr_17_17 : OUT std_logic ;
         d_arr_17_16 : OUT std_logic ;
         d_arr_17_15 : OUT std_logic ;
         d_arr_17_14 : OUT std_logic ;
         d_arr_17_13 : OUT std_logic ;
         d_arr_17_12 : OUT std_logic ;
         d_arr_17_11 : OUT std_logic ;
         d_arr_17_10 : OUT std_logic ;
         d_arr_17_9 : OUT std_logic ;
         d_arr_17_8 : OUT std_logic ;
         d_arr_17_7 : OUT std_logic ;
         d_arr_17_6 : OUT std_logic ;
         d_arr_17_5 : OUT std_logic ;
         d_arr_17_4 : OUT std_logic ;
         d_arr_17_3 : OUT std_logic ;
         d_arr_17_2 : OUT std_logic ;
         d_arr_17_1 : OUT std_logic ;
         d_arr_17_0 : OUT std_logic ;
         d_arr_18_31 : OUT std_logic ;
         d_arr_18_30 : OUT std_logic ;
         d_arr_18_29 : OUT std_logic ;
         d_arr_18_28 : OUT std_logic ;
         d_arr_18_27 : OUT std_logic ;
         d_arr_18_26 : OUT std_logic ;
         d_arr_18_25 : OUT std_logic ;
         d_arr_18_24 : OUT std_logic ;
         d_arr_18_23 : OUT std_logic ;
         d_arr_18_22 : OUT std_logic ;
         d_arr_18_21 : OUT std_logic ;
         d_arr_18_20 : OUT std_logic ;
         d_arr_18_19 : OUT std_logic ;
         d_arr_18_18 : OUT std_logic ;
         d_arr_18_17 : OUT std_logic ;
         d_arr_18_16 : OUT std_logic ;
         d_arr_18_15 : OUT std_logic ;
         d_arr_18_14 : OUT std_logic ;
         d_arr_18_13 : OUT std_logic ;
         d_arr_18_12 : OUT std_logic ;
         d_arr_18_11 : OUT std_logic ;
         d_arr_18_10 : OUT std_logic ;
         d_arr_18_9 : OUT std_logic ;
         d_arr_18_8 : OUT std_logic ;
         d_arr_18_7 : OUT std_logic ;
         d_arr_18_6 : OUT std_logic ;
         d_arr_18_5 : OUT std_logic ;
         d_arr_18_4 : OUT std_logic ;
         d_arr_18_3 : OUT std_logic ;
         d_arr_18_2 : OUT std_logic ;
         d_arr_18_1 : OUT std_logic ;
         d_arr_18_0 : OUT std_logic ;
         d_arr_19_31 : OUT std_logic ;
         d_arr_19_30 : OUT std_logic ;
         d_arr_19_29 : OUT std_logic ;
         d_arr_19_28 : OUT std_logic ;
         d_arr_19_27 : OUT std_logic ;
         d_arr_19_26 : OUT std_logic ;
         d_arr_19_25 : OUT std_logic ;
         d_arr_19_24 : OUT std_logic ;
         d_arr_19_23 : OUT std_logic ;
         d_arr_19_22 : OUT std_logic ;
         d_arr_19_21 : OUT std_logic ;
         d_arr_19_20 : OUT std_logic ;
         d_arr_19_19 : OUT std_logic ;
         d_arr_19_18 : OUT std_logic ;
         d_arr_19_17 : OUT std_logic ;
         d_arr_19_16 : OUT std_logic ;
         d_arr_19_15 : OUT std_logic ;
         d_arr_19_14 : OUT std_logic ;
         d_arr_19_13 : OUT std_logic ;
         d_arr_19_12 : OUT std_logic ;
         d_arr_19_11 : OUT std_logic ;
         d_arr_19_10 : OUT std_logic ;
         d_arr_19_9 : OUT std_logic ;
         d_arr_19_8 : OUT std_logic ;
         d_arr_19_7 : OUT std_logic ;
         d_arr_19_6 : OUT std_logic ;
         d_arr_19_5 : OUT std_logic ;
         d_arr_19_4 : OUT std_logic ;
         d_arr_19_3 : OUT std_logic ;
         d_arr_19_2 : OUT std_logic ;
         d_arr_19_1 : OUT std_logic ;
         d_arr_19_0 : OUT std_logic ;
         d_arr_20_31 : OUT std_logic ;
         d_arr_20_30 : OUT std_logic ;
         d_arr_20_29 : OUT std_logic ;
         d_arr_20_28 : OUT std_logic ;
         d_arr_20_27 : OUT std_logic ;
         d_arr_20_26 : OUT std_logic ;
         d_arr_20_25 : OUT std_logic ;
         d_arr_20_24 : OUT std_logic ;
         d_arr_20_23 : OUT std_logic ;
         d_arr_20_22 : OUT std_logic ;
         d_arr_20_21 : OUT std_logic ;
         d_arr_20_20 : OUT std_logic ;
         d_arr_20_19 : OUT std_logic ;
         d_arr_20_18 : OUT std_logic ;
         d_arr_20_17 : OUT std_logic ;
         d_arr_20_16 : OUT std_logic ;
         d_arr_20_15 : OUT std_logic ;
         d_arr_20_14 : OUT std_logic ;
         d_arr_20_13 : OUT std_logic ;
         d_arr_20_12 : OUT std_logic ;
         d_arr_20_11 : OUT std_logic ;
         d_arr_20_10 : OUT std_logic ;
         d_arr_20_9 : OUT std_logic ;
         d_arr_20_8 : OUT std_logic ;
         d_arr_20_7 : OUT std_logic ;
         d_arr_20_6 : OUT std_logic ;
         d_arr_20_5 : OUT std_logic ;
         d_arr_20_4 : OUT std_logic ;
         d_arr_20_3 : OUT std_logic ;
         d_arr_20_2 : OUT std_logic ;
         d_arr_20_1 : OUT std_logic ;
         d_arr_20_0 : OUT std_logic ;
         d_arr_21_31 : OUT std_logic ;
         d_arr_21_30 : OUT std_logic ;
         d_arr_21_29 : OUT std_logic ;
         d_arr_21_28 : OUT std_logic ;
         d_arr_21_27 : OUT std_logic ;
         d_arr_21_26 : OUT std_logic ;
         d_arr_21_25 : OUT std_logic ;
         d_arr_21_24 : OUT std_logic ;
         d_arr_21_23 : OUT std_logic ;
         d_arr_21_22 : OUT std_logic ;
         d_arr_21_21 : OUT std_logic ;
         d_arr_21_20 : OUT std_logic ;
         d_arr_21_19 : OUT std_logic ;
         d_arr_21_18 : OUT std_logic ;
         d_arr_21_17 : OUT std_logic ;
         d_arr_21_16 : OUT std_logic ;
         d_arr_21_15 : OUT std_logic ;
         d_arr_21_14 : OUT std_logic ;
         d_arr_21_13 : OUT std_logic ;
         d_arr_21_12 : OUT std_logic ;
         d_arr_21_11 : OUT std_logic ;
         d_arr_21_10 : OUT std_logic ;
         d_arr_21_9 : OUT std_logic ;
         d_arr_21_8 : OUT std_logic ;
         d_arr_21_7 : OUT std_logic ;
         d_arr_21_6 : OUT std_logic ;
         d_arr_21_5 : OUT std_logic ;
         d_arr_21_4 : OUT std_logic ;
         d_arr_21_3 : OUT std_logic ;
         d_arr_21_2 : OUT std_logic ;
         d_arr_21_1 : OUT std_logic ;
         d_arr_21_0 : OUT std_logic ;
         d_arr_22_31 : OUT std_logic ;
         d_arr_22_30 : OUT std_logic ;
         d_arr_22_29 : OUT std_logic ;
         d_arr_22_28 : OUT std_logic ;
         d_arr_22_27 : OUT std_logic ;
         d_arr_22_26 : OUT std_logic ;
         d_arr_22_25 : OUT std_logic ;
         d_arr_22_24 : OUT std_logic ;
         d_arr_22_23 : OUT std_logic ;
         d_arr_22_22 : OUT std_logic ;
         d_arr_22_21 : OUT std_logic ;
         d_arr_22_20 : OUT std_logic ;
         d_arr_22_19 : OUT std_logic ;
         d_arr_22_18 : OUT std_logic ;
         d_arr_22_17 : OUT std_logic ;
         d_arr_22_16 : OUT std_logic ;
         d_arr_22_15 : OUT std_logic ;
         d_arr_22_14 : OUT std_logic ;
         d_arr_22_13 : OUT std_logic ;
         d_arr_22_12 : OUT std_logic ;
         d_arr_22_11 : OUT std_logic ;
         d_arr_22_10 : OUT std_logic ;
         d_arr_22_9 : OUT std_logic ;
         d_arr_22_8 : OUT std_logic ;
         d_arr_22_7 : OUT std_logic ;
         d_arr_22_6 : OUT std_logic ;
         d_arr_22_5 : OUT std_logic ;
         d_arr_22_4 : OUT std_logic ;
         d_arr_22_3 : OUT std_logic ;
         d_arr_22_2 : OUT std_logic ;
         d_arr_22_1 : OUT std_logic ;
         d_arr_22_0 : OUT std_logic ;
         d_arr_23_31 : OUT std_logic ;
         d_arr_23_30 : OUT std_logic ;
         d_arr_23_29 : OUT std_logic ;
         d_arr_23_28 : OUT std_logic ;
         d_arr_23_27 : OUT std_logic ;
         d_arr_23_26 : OUT std_logic ;
         d_arr_23_25 : OUT std_logic ;
         d_arr_23_24 : OUT std_logic ;
         d_arr_23_23 : OUT std_logic ;
         d_arr_23_22 : OUT std_logic ;
         d_arr_23_21 : OUT std_logic ;
         d_arr_23_20 : OUT std_logic ;
         d_arr_23_19 : OUT std_logic ;
         d_arr_23_18 : OUT std_logic ;
         d_arr_23_17 : OUT std_logic ;
         d_arr_23_16 : OUT std_logic ;
         d_arr_23_15 : OUT std_logic ;
         d_arr_23_14 : OUT std_logic ;
         d_arr_23_13 : OUT std_logic ;
         d_arr_23_12 : OUT std_logic ;
         d_arr_23_11 : OUT std_logic ;
         d_arr_23_10 : OUT std_logic ;
         d_arr_23_9 : OUT std_logic ;
         d_arr_23_8 : OUT std_logic ;
         d_arr_23_7 : OUT std_logic ;
         d_arr_23_6 : OUT std_logic ;
         d_arr_23_5 : OUT std_logic ;
         d_arr_23_4 : OUT std_logic ;
         d_arr_23_3 : OUT std_logic ;
         d_arr_23_2 : OUT std_logic ;
         d_arr_23_1 : OUT std_logic ;
         d_arr_23_0 : OUT std_logic ;
         d_arr_24_31 : OUT std_logic ;
         d_arr_24_30 : OUT std_logic ;
         d_arr_24_29 : OUT std_logic ;
         d_arr_24_28 : OUT std_logic ;
         d_arr_24_27 : OUT std_logic ;
         d_arr_24_26 : OUT std_logic ;
         d_arr_24_25 : OUT std_logic ;
         d_arr_24_24 : OUT std_logic ;
         d_arr_24_23 : OUT std_logic ;
         d_arr_24_22 : OUT std_logic ;
         d_arr_24_21 : OUT std_logic ;
         d_arr_24_20 : OUT std_logic ;
         d_arr_24_19 : OUT std_logic ;
         d_arr_24_18 : OUT std_logic ;
         d_arr_24_17 : OUT std_logic ;
         d_arr_24_16 : OUT std_logic ;
         d_arr_24_15 : OUT std_logic ;
         d_arr_24_14 : OUT std_logic ;
         d_arr_24_13 : OUT std_logic ;
         d_arr_24_12 : OUT std_logic ;
         d_arr_24_11 : OUT std_logic ;
         d_arr_24_10 : OUT std_logic ;
         d_arr_24_9 : OUT std_logic ;
         d_arr_24_8 : OUT std_logic ;
         d_arr_24_7 : OUT std_logic ;
         d_arr_24_6 : OUT std_logic ;
         d_arr_24_5 : OUT std_logic ;
         d_arr_24_4 : OUT std_logic ;
         d_arr_24_3 : OUT std_logic ;
         d_arr_24_2 : OUT std_logic ;
         d_arr_24_1 : OUT std_logic ;
         d_arr_24_0 : OUT std_logic) ;
   end component ;
   component MuxLayer
      port (
         img_data_0_31 : IN std_logic ;
         img_data_0_30 : IN std_logic ;
         img_data_0_29 : IN std_logic ;
         img_data_0_28 : IN std_logic ;
         img_data_0_27 : IN std_logic ;
         img_data_0_26 : IN std_logic ;
         img_data_0_25 : IN std_logic ;
         img_data_0_24 : IN std_logic ;
         img_data_0_23 : IN std_logic ;
         img_data_0_22 : IN std_logic ;
         img_data_0_21 : IN std_logic ;
         img_data_0_20 : IN std_logic ;
         img_data_0_19 : IN std_logic ;
         img_data_0_18 : IN std_logic ;
         img_data_0_17 : IN std_logic ;
         img_data_0_16 : IN std_logic ;
         img_data_0_15 : IN std_logic ;
         img_data_0_14 : IN std_logic ;
         img_data_0_13 : IN std_logic ;
         img_data_0_12 : IN std_logic ;
         img_data_0_11 : IN std_logic ;
         img_data_0_10 : IN std_logic ;
         img_data_0_9 : IN std_logic ;
         img_data_0_8 : IN std_logic ;
         img_data_0_7 : IN std_logic ;
         img_data_0_6 : IN std_logic ;
         img_data_0_5 : IN std_logic ;
         img_data_0_4 : IN std_logic ;
         img_data_0_3 : IN std_logic ;
         img_data_0_2 : IN std_logic ;
         img_data_0_1 : IN std_logic ;
         img_data_0_0 : IN std_logic ;
         img_data_1_31 : IN std_logic ;
         img_data_1_30 : IN std_logic ;
         img_data_1_29 : IN std_logic ;
         img_data_1_28 : IN std_logic ;
         img_data_1_27 : IN std_logic ;
         img_data_1_26 : IN std_logic ;
         img_data_1_25 : IN std_logic ;
         img_data_1_24 : IN std_logic ;
         img_data_1_23 : IN std_logic ;
         img_data_1_22 : IN std_logic ;
         img_data_1_21 : IN std_logic ;
         img_data_1_20 : IN std_logic ;
         img_data_1_19 : IN std_logic ;
         img_data_1_18 : IN std_logic ;
         img_data_1_17 : IN std_logic ;
         img_data_1_16 : IN std_logic ;
         img_data_1_15 : IN std_logic ;
         img_data_1_14 : IN std_logic ;
         img_data_1_13 : IN std_logic ;
         img_data_1_12 : IN std_logic ;
         img_data_1_11 : IN std_logic ;
         img_data_1_10 : IN std_logic ;
         img_data_1_9 : IN std_logic ;
         img_data_1_8 : IN std_logic ;
         img_data_1_7 : IN std_logic ;
         img_data_1_6 : IN std_logic ;
         img_data_1_5 : IN std_logic ;
         img_data_1_4 : IN std_logic ;
         img_data_1_3 : IN std_logic ;
         img_data_1_2 : IN std_logic ;
         img_data_1_1 : IN std_logic ;
         img_data_1_0 : IN std_logic ;
         img_data_2_31 : IN std_logic ;
         img_data_2_30 : IN std_logic ;
         img_data_2_29 : IN std_logic ;
         img_data_2_28 : IN std_logic ;
         img_data_2_27 : IN std_logic ;
         img_data_2_26 : IN std_logic ;
         img_data_2_25 : IN std_logic ;
         img_data_2_24 : IN std_logic ;
         img_data_2_23 : IN std_logic ;
         img_data_2_22 : IN std_logic ;
         img_data_2_21 : IN std_logic ;
         img_data_2_20 : IN std_logic ;
         img_data_2_19 : IN std_logic ;
         img_data_2_18 : IN std_logic ;
         img_data_2_17 : IN std_logic ;
         img_data_2_16 : IN std_logic ;
         img_data_2_15 : IN std_logic ;
         img_data_2_14 : IN std_logic ;
         img_data_2_13 : IN std_logic ;
         img_data_2_12 : IN std_logic ;
         img_data_2_11 : IN std_logic ;
         img_data_2_10 : IN std_logic ;
         img_data_2_9 : IN std_logic ;
         img_data_2_8 : IN std_logic ;
         img_data_2_7 : IN std_logic ;
         img_data_2_6 : IN std_logic ;
         img_data_2_5 : IN std_logic ;
         img_data_2_4 : IN std_logic ;
         img_data_2_3 : IN std_logic ;
         img_data_2_2 : IN std_logic ;
         img_data_2_1 : IN std_logic ;
         img_data_2_0 : IN std_logic ;
         img_data_3_31 : IN std_logic ;
         img_data_3_30 : IN std_logic ;
         img_data_3_29 : IN std_logic ;
         img_data_3_28 : IN std_logic ;
         img_data_3_27 : IN std_logic ;
         img_data_3_26 : IN std_logic ;
         img_data_3_25 : IN std_logic ;
         img_data_3_24 : IN std_logic ;
         img_data_3_23 : IN std_logic ;
         img_data_3_22 : IN std_logic ;
         img_data_3_21 : IN std_logic ;
         img_data_3_20 : IN std_logic ;
         img_data_3_19 : IN std_logic ;
         img_data_3_18 : IN std_logic ;
         img_data_3_17 : IN std_logic ;
         img_data_3_16 : IN std_logic ;
         img_data_3_15 : IN std_logic ;
         img_data_3_14 : IN std_logic ;
         img_data_3_13 : IN std_logic ;
         img_data_3_12 : IN std_logic ;
         img_data_3_11 : IN std_logic ;
         img_data_3_10 : IN std_logic ;
         img_data_3_9 : IN std_logic ;
         img_data_3_8 : IN std_logic ;
         img_data_3_7 : IN std_logic ;
         img_data_3_6 : IN std_logic ;
         img_data_3_5 : IN std_logic ;
         img_data_3_4 : IN std_logic ;
         img_data_3_3 : IN std_logic ;
         img_data_3_2 : IN std_logic ;
         img_data_3_1 : IN std_logic ;
         img_data_3_0 : IN std_logic ;
         img_data_4_31 : IN std_logic ;
         img_data_4_30 : IN std_logic ;
         img_data_4_29 : IN std_logic ;
         img_data_4_28 : IN std_logic ;
         img_data_4_27 : IN std_logic ;
         img_data_4_26 : IN std_logic ;
         img_data_4_25 : IN std_logic ;
         img_data_4_24 : IN std_logic ;
         img_data_4_23 : IN std_logic ;
         img_data_4_22 : IN std_logic ;
         img_data_4_21 : IN std_logic ;
         img_data_4_20 : IN std_logic ;
         img_data_4_19 : IN std_logic ;
         img_data_4_18 : IN std_logic ;
         img_data_4_17 : IN std_logic ;
         img_data_4_16 : IN std_logic ;
         img_data_4_15 : IN std_logic ;
         img_data_4_14 : IN std_logic ;
         img_data_4_13 : IN std_logic ;
         img_data_4_12 : IN std_logic ;
         img_data_4_11 : IN std_logic ;
         img_data_4_10 : IN std_logic ;
         img_data_4_9 : IN std_logic ;
         img_data_4_8 : IN std_logic ;
         img_data_4_7 : IN std_logic ;
         img_data_4_6 : IN std_logic ;
         img_data_4_5 : IN std_logic ;
         img_data_4_4 : IN std_logic ;
         img_data_4_3 : IN std_logic ;
         img_data_4_2 : IN std_logic ;
         img_data_4_1 : IN std_logic ;
         img_data_4_0 : IN std_logic ;
         img_data_5_31 : IN std_logic ;
         img_data_5_30 : IN std_logic ;
         img_data_5_29 : IN std_logic ;
         img_data_5_28 : IN std_logic ;
         img_data_5_27 : IN std_logic ;
         img_data_5_26 : IN std_logic ;
         img_data_5_25 : IN std_logic ;
         img_data_5_24 : IN std_logic ;
         img_data_5_23 : IN std_logic ;
         img_data_5_22 : IN std_logic ;
         img_data_5_21 : IN std_logic ;
         img_data_5_20 : IN std_logic ;
         img_data_5_19 : IN std_logic ;
         img_data_5_18 : IN std_logic ;
         img_data_5_17 : IN std_logic ;
         img_data_5_16 : IN std_logic ;
         img_data_5_15 : IN std_logic ;
         img_data_5_14 : IN std_logic ;
         img_data_5_13 : IN std_logic ;
         img_data_5_12 : IN std_logic ;
         img_data_5_11 : IN std_logic ;
         img_data_5_10 : IN std_logic ;
         img_data_5_9 : IN std_logic ;
         img_data_5_8 : IN std_logic ;
         img_data_5_7 : IN std_logic ;
         img_data_5_6 : IN std_logic ;
         img_data_5_5 : IN std_logic ;
         img_data_5_4 : IN std_logic ;
         img_data_5_3 : IN std_logic ;
         img_data_5_2 : IN std_logic ;
         img_data_5_1 : IN std_logic ;
         img_data_5_0 : IN std_logic ;
         img_data_6_31 : IN std_logic ;
         img_data_6_30 : IN std_logic ;
         img_data_6_29 : IN std_logic ;
         img_data_6_28 : IN std_logic ;
         img_data_6_27 : IN std_logic ;
         img_data_6_26 : IN std_logic ;
         img_data_6_25 : IN std_logic ;
         img_data_6_24 : IN std_logic ;
         img_data_6_23 : IN std_logic ;
         img_data_6_22 : IN std_logic ;
         img_data_6_21 : IN std_logic ;
         img_data_6_20 : IN std_logic ;
         img_data_6_19 : IN std_logic ;
         img_data_6_18 : IN std_logic ;
         img_data_6_17 : IN std_logic ;
         img_data_6_16 : IN std_logic ;
         img_data_6_15 : IN std_logic ;
         img_data_6_14 : IN std_logic ;
         img_data_6_13 : IN std_logic ;
         img_data_6_12 : IN std_logic ;
         img_data_6_11 : IN std_logic ;
         img_data_6_10 : IN std_logic ;
         img_data_6_9 : IN std_logic ;
         img_data_6_8 : IN std_logic ;
         img_data_6_7 : IN std_logic ;
         img_data_6_6 : IN std_logic ;
         img_data_6_5 : IN std_logic ;
         img_data_6_4 : IN std_logic ;
         img_data_6_3 : IN std_logic ;
         img_data_6_2 : IN std_logic ;
         img_data_6_1 : IN std_logic ;
         img_data_6_0 : IN std_logic ;
         img_data_7_31 : IN std_logic ;
         img_data_7_30 : IN std_logic ;
         img_data_7_29 : IN std_logic ;
         img_data_7_28 : IN std_logic ;
         img_data_7_27 : IN std_logic ;
         img_data_7_26 : IN std_logic ;
         img_data_7_25 : IN std_logic ;
         img_data_7_24 : IN std_logic ;
         img_data_7_23 : IN std_logic ;
         img_data_7_22 : IN std_logic ;
         img_data_7_21 : IN std_logic ;
         img_data_7_20 : IN std_logic ;
         img_data_7_19 : IN std_logic ;
         img_data_7_18 : IN std_logic ;
         img_data_7_17 : IN std_logic ;
         img_data_7_16 : IN std_logic ;
         img_data_7_15 : IN std_logic ;
         img_data_7_14 : IN std_logic ;
         img_data_7_13 : IN std_logic ;
         img_data_7_12 : IN std_logic ;
         img_data_7_11 : IN std_logic ;
         img_data_7_10 : IN std_logic ;
         img_data_7_9 : IN std_logic ;
         img_data_7_8 : IN std_logic ;
         img_data_7_7 : IN std_logic ;
         img_data_7_6 : IN std_logic ;
         img_data_7_5 : IN std_logic ;
         img_data_7_4 : IN std_logic ;
         img_data_7_3 : IN std_logic ;
         img_data_7_2 : IN std_logic ;
         img_data_7_1 : IN std_logic ;
         img_data_7_0 : IN std_logic ;
         img_data_8_31 : IN std_logic ;
         img_data_8_30 : IN std_logic ;
         img_data_8_29 : IN std_logic ;
         img_data_8_28 : IN std_logic ;
         img_data_8_27 : IN std_logic ;
         img_data_8_26 : IN std_logic ;
         img_data_8_25 : IN std_logic ;
         img_data_8_24 : IN std_logic ;
         img_data_8_23 : IN std_logic ;
         img_data_8_22 : IN std_logic ;
         img_data_8_21 : IN std_logic ;
         img_data_8_20 : IN std_logic ;
         img_data_8_19 : IN std_logic ;
         img_data_8_18 : IN std_logic ;
         img_data_8_17 : IN std_logic ;
         img_data_8_16 : IN std_logic ;
         img_data_8_15 : IN std_logic ;
         img_data_8_14 : IN std_logic ;
         img_data_8_13 : IN std_logic ;
         img_data_8_12 : IN std_logic ;
         img_data_8_11 : IN std_logic ;
         img_data_8_10 : IN std_logic ;
         img_data_8_9 : IN std_logic ;
         img_data_8_8 : IN std_logic ;
         img_data_8_7 : IN std_logic ;
         img_data_8_6 : IN std_logic ;
         img_data_8_5 : IN std_logic ;
         img_data_8_4 : IN std_logic ;
         img_data_8_3 : IN std_logic ;
         img_data_8_2 : IN std_logic ;
         img_data_8_1 : IN std_logic ;
         img_data_8_0 : IN std_logic ;
         img_data_9_31 : IN std_logic ;
         img_data_9_30 : IN std_logic ;
         img_data_9_29 : IN std_logic ;
         img_data_9_28 : IN std_logic ;
         img_data_9_27 : IN std_logic ;
         img_data_9_26 : IN std_logic ;
         img_data_9_25 : IN std_logic ;
         img_data_9_24 : IN std_logic ;
         img_data_9_23 : IN std_logic ;
         img_data_9_22 : IN std_logic ;
         img_data_9_21 : IN std_logic ;
         img_data_9_20 : IN std_logic ;
         img_data_9_19 : IN std_logic ;
         img_data_9_18 : IN std_logic ;
         img_data_9_17 : IN std_logic ;
         img_data_9_16 : IN std_logic ;
         img_data_9_15 : IN std_logic ;
         img_data_9_14 : IN std_logic ;
         img_data_9_13 : IN std_logic ;
         img_data_9_12 : IN std_logic ;
         img_data_9_11 : IN std_logic ;
         img_data_9_10 : IN std_logic ;
         img_data_9_9 : IN std_logic ;
         img_data_9_8 : IN std_logic ;
         img_data_9_7 : IN std_logic ;
         img_data_9_6 : IN std_logic ;
         img_data_9_5 : IN std_logic ;
         img_data_9_4 : IN std_logic ;
         img_data_9_3 : IN std_logic ;
         img_data_9_2 : IN std_logic ;
         img_data_9_1 : IN std_logic ;
         img_data_9_0 : IN std_logic ;
         img_data_10_31 : IN std_logic ;
         img_data_10_30 : IN std_logic ;
         img_data_10_29 : IN std_logic ;
         img_data_10_28 : IN std_logic ;
         img_data_10_27 : IN std_logic ;
         img_data_10_26 : IN std_logic ;
         img_data_10_25 : IN std_logic ;
         img_data_10_24 : IN std_logic ;
         img_data_10_23 : IN std_logic ;
         img_data_10_22 : IN std_logic ;
         img_data_10_21 : IN std_logic ;
         img_data_10_20 : IN std_logic ;
         img_data_10_19 : IN std_logic ;
         img_data_10_18 : IN std_logic ;
         img_data_10_17 : IN std_logic ;
         img_data_10_16 : IN std_logic ;
         img_data_10_15 : IN std_logic ;
         img_data_10_14 : IN std_logic ;
         img_data_10_13 : IN std_logic ;
         img_data_10_12 : IN std_logic ;
         img_data_10_11 : IN std_logic ;
         img_data_10_10 : IN std_logic ;
         img_data_10_9 : IN std_logic ;
         img_data_10_8 : IN std_logic ;
         img_data_10_7 : IN std_logic ;
         img_data_10_6 : IN std_logic ;
         img_data_10_5 : IN std_logic ;
         img_data_10_4 : IN std_logic ;
         img_data_10_3 : IN std_logic ;
         img_data_10_2 : IN std_logic ;
         img_data_10_1 : IN std_logic ;
         img_data_10_0 : IN std_logic ;
         img_data_11_31 : IN std_logic ;
         img_data_11_30 : IN std_logic ;
         img_data_11_29 : IN std_logic ;
         img_data_11_28 : IN std_logic ;
         img_data_11_27 : IN std_logic ;
         img_data_11_26 : IN std_logic ;
         img_data_11_25 : IN std_logic ;
         img_data_11_24 : IN std_logic ;
         img_data_11_23 : IN std_logic ;
         img_data_11_22 : IN std_logic ;
         img_data_11_21 : IN std_logic ;
         img_data_11_20 : IN std_logic ;
         img_data_11_19 : IN std_logic ;
         img_data_11_18 : IN std_logic ;
         img_data_11_17 : IN std_logic ;
         img_data_11_16 : IN std_logic ;
         img_data_11_15 : IN std_logic ;
         img_data_11_14 : IN std_logic ;
         img_data_11_13 : IN std_logic ;
         img_data_11_12 : IN std_logic ;
         img_data_11_11 : IN std_logic ;
         img_data_11_10 : IN std_logic ;
         img_data_11_9 : IN std_logic ;
         img_data_11_8 : IN std_logic ;
         img_data_11_7 : IN std_logic ;
         img_data_11_6 : IN std_logic ;
         img_data_11_5 : IN std_logic ;
         img_data_11_4 : IN std_logic ;
         img_data_11_3 : IN std_logic ;
         img_data_11_2 : IN std_logic ;
         img_data_11_1 : IN std_logic ;
         img_data_11_0 : IN std_logic ;
         img_data_12_31 : IN std_logic ;
         img_data_12_30 : IN std_logic ;
         img_data_12_29 : IN std_logic ;
         img_data_12_28 : IN std_logic ;
         img_data_12_27 : IN std_logic ;
         img_data_12_26 : IN std_logic ;
         img_data_12_25 : IN std_logic ;
         img_data_12_24 : IN std_logic ;
         img_data_12_23 : IN std_logic ;
         img_data_12_22 : IN std_logic ;
         img_data_12_21 : IN std_logic ;
         img_data_12_20 : IN std_logic ;
         img_data_12_19 : IN std_logic ;
         img_data_12_18 : IN std_logic ;
         img_data_12_17 : IN std_logic ;
         img_data_12_16 : IN std_logic ;
         img_data_12_15 : IN std_logic ;
         img_data_12_14 : IN std_logic ;
         img_data_12_13 : IN std_logic ;
         img_data_12_12 : IN std_logic ;
         img_data_12_11 : IN std_logic ;
         img_data_12_10 : IN std_logic ;
         img_data_12_9 : IN std_logic ;
         img_data_12_8 : IN std_logic ;
         img_data_12_7 : IN std_logic ;
         img_data_12_6 : IN std_logic ;
         img_data_12_5 : IN std_logic ;
         img_data_12_4 : IN std_logic ;
         img_data_12_3 : IN std_logic ;
         img_data_12_2 : IN std_logic ;
         img_data_12_1 : IN std_logic ;
         img_data_12_0 : IN std_logic ;
         img_data_13_31 : IN std_logic ;
         img_data_13_30 : IN std_logic ;
         img_data_13_29 : IN std_logic ;
         img_data_13_28 : IN std_logic ;
         img_data_13_27 : IN std_logic ;
         img_data_13_26 : IN std_logic ;
         img_data_13_25 : IN std_logic ;
         img_data_13_24 : IN std_logic ;
         img_data_13_23 : IN std_logic ;
         img_data_13_22 : IN std_logic ;
         img_data_13_21 : IN std_logic ;
         img_data_13_20 : IN std_logic ;
         img_data_13_19 : IN std_logic ;
         img_data_13_18 : IN std_logic ;
         img_data_13_17 : IN std_logic ;
         img_data_13_16 : IN std_logic ;
         img_data_13_15 : IN std_logic ;
         img_data_13_14 : IN std_logic ;
         img_data_13_13 : IN std_logic ;
         img_data_13_12 : IN std_logic ;
         img_data_13_11 : IN std_logic ;
         img_data_13_10 : IN std_logic ;
         img_data_13_9 : IN std_logic ;
         img_data_13_8 : IN std_logic ;
         img_data_13_7 : IN std_logic ;
         img_data_13_6 : IN std_logic ;
         img_data_13_5 : IN std_logic ;
         img_data_13_4 : IN std_logic ;
         img_data_13_3 : IN std_logic ;
         img_data_13_2 : IN std_logic ;
         img_data_13_1 : IN std_logic ;
         img_data_13_0 : IN std_logic ;
         img_data_14_31 : IN std_logic ;
         img_data_14_30 : IN std_logic ;
         img_data_14_29 : IN std_logic ;
         img_data_14_28 : IN std_logic ;
         img_data_14_27 : IN std_logic ;
         img_data_14_26 : IN std_logic ;
         img_data_14_25 : IN std_logic ;
         img_data_14_24 : IN std_logic ;
         img_data_14_23 : IN std_logic ;
         img_data_14_22 : IN std_logic ;
         img_data_14_21 : IN std_logic ;
         img_data_14_20 : IN std_logic ;
         img_data_14_19 : IN std_logic ;
         img_data_14_18 : IN std_logic ;
         img_data_14_17 : IN std_logic ;
         img_data_14_16 : IN std_logic ;
         img_data_14_15 : IN std_logic ;
         img_data_14_14 : IN std_logic ;
         img_data_14_13 : IN std_logic ;
         img_data_14_12 : IN std_logic ;
         img_data_14_11 : IN std_logic ;
         img_data_14_10 : IN std_logic ;
         img_data_14_9 : IN std_logic ;
         img_data_14_8 : IN std_logic ;
         img_data_14_7 : IN std_logic ;
         img_data_14_6 : IN std_logic ;
         img_data_14_5 : IN std_logic ;
         img_data_14_4 : IN std_logic ;
         img_data_14_3 : IN std_logic ;
         img_data_14_2 : IN std_logic ;
         img_data_14_1 : IN std_logic ;
         img_data_14_0 : IN std_logic ;
         img_data_15_31 : IN std_logic ;
         img_data_15_30 : IN std_logic ;
         img_data_15_29 : IN std_logic ;
         img_data_15_28 : IN std_logic ;
         img_data_15_27 : IN std_logic ;
         img_data_15_26 : IN std_logic ;
         img_data_15_25 : IN std_logic ;
         img_data_15_24 : IN std_logic ;
         img_data_15_23 : IN std_logic ;
         img_data_15_22 : IN std_logic ;
         img_data_15_21 : IN std_logic ;
         img_data_15_20 : IN std_logic ;
         img_data_15_19 : IN std_logic ;
         img_data_15_18 : IN std_logic ;
         img_data_15_17 : IN std_logic ;
         img_data_15_16 : IN std_logic ;
         img_data_15_15 : IN std_logic ;
         img_data_15_14 : IN std_logic ;
         img_data_15_13 : IN std_logic ;
         img_data_15_12 : IN std_logic ;
         img_data_15_11 : IN std_logic ;
         img_data_15_10 : IN std_logic ;
         img_data_15_9 : IN std_logic ;
         img_data_15_8 : IN std_logic ;
         img_data_15_7 : IN std_logic ;
         img_data_15_6 : IN std_logic ;
         img_data_15_5 : IN std_logic ;
         img_data_15_4 : IN std_logic ;
         img_data_15_3 : IN std_logic ;
         img_data_15_2 : IN std_logic ;
         img_data_15_1 : IN std_logic ;
         img_data_15_0 : IN std_logic ;
         img_data_16_31 : IN std_logic ;
         img_data_16_30 : IN std_logic ;
         img_data_16_29 : IN std_logic ;
         img_data_16_28 : IN std_logic ;
         img_data_16_27 : IN std_logic ;
         img_data_16_26 : IN std_logic ;
         img_data_16_25 : IN std_logic ;
         img_data_16_24 : IN std_logic ;
         img_data_16_23 : IN std_logic ;
         img_data_16_22 : IN std_logic ;
         img_data_16_21 : IN std_logic ;
         img_data_16_20 : IN std_logic ;
         img_data_16_19 : IN std_logic ;
         img_data_16_18 : IN std_logic ;
         img_data_16_17 : IN std_logic ;
         img_data_16_16 : IN std_logic ;
         img_data_16_15 : IN std_logic ;
         img_data_16_14 : IN std_logic ;
         img_data_16_13 : IN std_logic ;
         img_data_16_12 : IN std_logic ;
         img_data_16_11 : IN std_logic ;
         img_data_16_10 : IN std_logic ;
         img_data_16_9 : IN std_logic ;
         img_data_16_8 : IN std_logic ;
         img_data_16_7 : IN std_logic ;
         img_data_16_6 : IN std_logic ;
         img_data_16_5 : IN std_logic ;
         img_data_16_4 : IN std_logic ;
         img_data_16_3 : IN std_logic ;
         img_data_16_2 : IN std_logic ;
         img_data_16_1 : IN std_logic ;
         img_data_16_0 : IN std_logic ;
         img_data_17_31 : IN std_logic ;
         img_data_17_30 : IN std_logic ;
         img_data_17_29 : IN std_logic ;
         img_data_17_28 : IN std_logic ;
         img_data_17_27 : IN std_logic ;
         img_data_17_26 : IN std_logic ;
         img_data_17_25 : IN std_logic ;
         img_data_17_24 : IN std_logic ;
         img_data_17_23 : IN std_logic ;
         img_data_17_22 : IN std_logic ;
         img_data_17_21 : IN std_logic ;
         img_data_17_20 : IN std_logic ;
         img_data_17_19 : IN std_logic ;
         img_data_17_18 : IN std_logic ;
         img_data_17_17 : IN std_logic ;
         img_data_17_16 : IN std_logic ;
         img_data_17_15 : IN std_logic ;
         img_data_17_14 : IN std_logic ;
         img_data_17_13 : IN std_logic ;
         img_data_17_12 : IN std_logic ;
         img_data_17_11 : IN std_logic ;
         img_data_17_10 : IN std_logic ;
         img_data_17_9 : IN std_logic ;
         img_data_17_8 : IN std_logic ;
         img_data_17_7 : IN std_logic ;
         img_data_17_6 : IN std_logic ;
         img_data_17_5 : IN std_logic ;
         img_data_17_4 : IN std_logic ;
         img_data_17_3 : IN std_logic ;
         img_data_17_2 : IN std_logic ;
         img_data_17_1 : IN std_logic ;
         img_data_17_0 : IN std_logic ;
         img_data_18_31 : IN std_logic ;
         img_data_18_30 : IN std_logic ;
         img_data_18_29 : IN std_logic ;
         img_data_18_28 : IN std_logic ;
         img_data_18_27 : IN std_logic ;
         img_data_18_26 : IN std_logic ;
         img_data_18_25 : IN std_logic ;
         img_data_18_24 : IN std_logic ;
         img_data_18_23 : IN std_logic ;
         img_data_18_22 : IN std_logic ;
         img_data_18_21 : IN std_logic ;
         img_data_18_20 : IN std_logic ;
         img_data_18_19 : IN std_logic ;
         img_data_18_18 : IN std_logic ;
         img_data_18_17 : IN std_logic ;
         img_data_18_16 : IN std_logic ;
         img_data_18_15 : IN std_logic ;
         img_data_18_14 : IN std_logic ;
         img_data_18_13 : IN std_logic ;
         img_data_18_12 : IN std_logic ;
         img_data_18_11 : IN std_logic ;
         img_data_18_10 : IN std_logic ;
         img_data_18_9 : IN std_logic ;
         img_data_18_8 : IN std_logic ;
         img_data_18_7 : IN std_logic ;
         img_data_18_6 : IN std_logic ;
         img_data_18_5 : IN std_logic ;
         img_data_18_4 : IN std_logic ;
         img_data_18_3 : IN std_logic ;
         img_data_18_2 : IN std_logic ;
         img_data_18_1 : IN std_logic ;
         img_data_18_0 : IN std_logic ;
         img_data_19_31 : IN std_logic ;
         img_data_19_30 : IN std_logic ;
         img_data_19_29 : IN std_logic ;
         img_data_19_28 : IN std_logic ;
         img_data_19_27 : IN std_logic ;
         img_data_19_26 : IN std_logic ;
         img_data_19_25 : IN std_logic ;
         img_data_19_24 : IN std_logic ;
         img_data_19_23 : IN std_logic ;
         img_data_19_22 : IN std_logic ;
         img_data_19_21 : IN std_logic ;
         img_data_19_20 : IN std_logic ;
         img_data_19_19 : IN std_logic ;
         img_data_19_18 : IN std_logic ;
         img_data_19_17 : IN std_logic ;
         img_data_19_16 : IN std_logic ;
         img_data_19_15 : IN std_logic ;
         img_data_19_14 : IN std_logic ;
         img_data_19_13 : IN std_logic ;
         img_data_19_12 : IN std_logic ;
         img_data_19_11 : IN std_logic ;
         img_data_19_10 : IN std_logic ;
         img_data_19_9 : IN std_logic ;
         img_data_19_8 : IN std_logic ;
         img_data_19_7 : IN std_logic ;
         img_data_19_6 : IN std_logic ;
         img_data_19_5 : IN std_logic ;
         img_data_19_4 : IN std_logic ;
         img_data_19_3 : IN std_logic ;
         img_data_19_2 : IN std_logic ;
         img_data_19_1 : IN std_logic ;
         img_data_19_0 : IN std_logic ;
         img_data_20_31 : IN std_logic ;
         img_data_20_30 : IN std_logic ;
         img_data_20_29 : IN std_logic ;
         img_data_20_28 : IN std_logic ;
         img_data_20_27 : IN std_logic ;
         img_data_20_26 : IN std_logic ;
         img_data_20_25 : IN std_logic ;
         img_data_20_24 : IN std_logic ;
         img_data_20_23 : IN std_logic ;
         img_data_20_22 : IN std_logic ;
         img_data_20_21 : IN std_logic ;
         img_data_20_20 : IN std_logic ;
         img_data_20_19 : IN std_logic ;
         img_data_20_18 : IN std_logic ;
         img_data_20_17 : IN std_logic ;
         img_data_20_16 : IN std_logic ;
         img_data_20_15 : IN std_logic ;
         img_data_20_14 : IN std_logic ;
         img_data_20_13 : IN std_logic ;
         img_data_20_12 : IN std_logic ;
         img_data_20_11 : IN std_logic ;
         img_data_20_10 : IN std_logic ;
         img_data_20_9 : IN std_logic ;
         img_data_20_8 : IN std_logic ;
         img_data_20_7 : IN std_logic ;
         img_data_20_6 : IN std_logic ;
         img_data_20_5 : IN std_logic ;
         img_data_20_4 : IN std_logic ;
         img_data_20_3 : IN std_logic ;
         img_data_20_2 : IN std_logic ;
         img_data_20_1 : IN std_logic ;
         img_data_20_0 : IN std_logic ;
         img_data_21_31 : IN std_logic ;
         img_data_21_30 : IN std_logic ;
         img_data_21_29 : IN std_logic ;
         img_data_21_28 : IN std_logic ;
         img_data_21_27 : IN std_logic ;
         img_data_21_26 : IN std_logic ;
         img_data_21_25 : IN std_logic ;
         img_data_21_24 : IN std_logic ;
         img_data_21_23 : IN std_logic ;
         img_data_21_22 : IN std_logic ;
         img_data_21_21 : IN std_logic ;
         img_data_21_20 : IN std_logic ;
         img_data_21_19 : IN std_logic ;
         img_data_21_18 : IN std_logic ;
         img_data_21_17 : IN std_logic ;
         img_data_21_16 : IN std_logic ;
         img_data_21_15 : IN std_logic ;
         img_data_21_14 : IN std_logic ;
         img_data_21_13 : IN std_logic ;
         img_data_21_12 : IN std_logic ;
         img_data_21_11 : IN std_logic ;
         img_data_21_10 : IN std_logic ;
         img_data_21_9 : IN std_logic ;
         img_data_21_8 : IN std_logic ;
         img_data_21_7 : IN std_logic ;
         img_data_21_6 : IN std_logic ;
         img_data_21_5 : IN std_logic ;
         img_data_21_4 : IN std_logic ;
         img_data_21_3 : IN std_logic ;
         img_data_21_2 : IN std_logic ;
         img_data_21_1 : IN std_logic ;
         img_data_21_0 : IN std_logic ;
         img_data_22_31 : IN std_logic ;
         img_data_22_30 : IN std_logic ;
         img_data_22_29 : IN std_logic ;
         img_data_22_28 : IN std_logic ;
         img_data_22_27 : IN std_logic ;
         img_data_22_26 : IN std_logic ;
         img_data_22_25 : IN std_logic ;
         img_data_22_24 : IN std_logic ;
         img_data_22_23 : IN std_logic ;
         img_data_22_22 : IN std_logic ;
         img_data_22_21 : IN std_logic ;
         img_data_22_20 : IN std_logic ;
         img_data_22_19 : IN std_logic ;
         img_data_22_18 : IN std_logic ;
         img_data_22_17 : IN std_logic ;
         img_data_22_16 : IN std_logic ;
         img_data_22_15 : IN std_logic ;
         img_data_22_14 : IN std_logic ;
         img_data_22_13 : IN std_logic ;
         img_data_22_12 : IN std_logic ;
         img_data_22_11 : IN std_logic ;
         img_data_22_10 : IN std_logic ;
         img_data_22_9 : IN std_logic ;
         img_data_22_8 : IN std_logic ;
         img_data_22_7 : IN std_logic ;
         img_data_22_6 : IN std_logic ;
         img_data_22_5 : IN std_logic ;
         img_data_22_4 : IN std_logic ;
         img_data_22_3 : IN std_logic ;
         img_data_22_2 : IN std_logic ;
         img_data_22_1 : IN std_logic ;
         img_data_22_0 : IN std_logic ;
         img_data_23_31 : IN std_logic ;
         img_data_23_30 : IN std_logic ;
         img_data_23_29 : IN std_logic ;
         img_data_23_28 : IN std_logic ;
         img_data_23_27 : IN std_logic ;
         img_data_23_26 : IN std_logic ;
         img_data_23_25 : IN std_logic ;
         img_data_23_24 : IN std_logic ;
         img_data_23_23 : IN std_logic ;
         img_data_23_22 : IN std_logic ;
         img_data_23_21 : IN std_logic ;
         img_data_23_20 : IN std_logic ;
         img_data_23_19 : IN std_logic ;
         img_data_23_18 : IN std_logic ;
         img_data_23_17 : IN std_logic ;
         img_data_23_16 : IN std_logic ;
         img_data_23_15 : IN std_logic ;
         img_data_23_14 : IN std_logic ;
         img_data_23_13 : IN std_logic ;
         img_data_23_12 : IN std_logic ;
         img_data_23_11 : IN std_logic ;
         img_data_23_10 : IN std_logic ;
         img_data_23_9 : IN std_logic ;
         img_data_23_8 : IN std_logic ;
         img_data_23_7 : IN std_logic ;
         img_data_23_6 : IN std_logic ;
         img_data_23_5 : IN std_logic ;
         img_data_23_4 : IN std_logic ;
         img_data_23_3 : IN std_logic ;
         img_data_23_2 : IN std_logic ;
         img_data_23_1 : IN std_logic ;
         img_data_23_0 : IN std_logic ;
         img_data_24_31 : IN std_logic ;
         img_data_24_30 : IN std_logic ;
         img_data_24_29 : IN std_logic ;
         img_data_24_28 : IN std_logic ;
         img_data_24_27 : IN std_logic ;
         img_data_24_26 : IN std_logic ;
         img_data_24_25 : IN std_logic ;
         img_data_24_24 : IN std_logic ;
         img_data_24_23 : IN std_logic ;
         img_data_24_22 : IN std_logic ;
         img_data_24_21 : IN std_logic ;
         img_data_24_20 : IN std_logic ;
         img_data_24_19 : IN std_logic ;
         img_data_24_18 : IN std_logic ;
         img_data_24_17 : IN std_logic ;
         img_data_24_16 : IN std_logic ;
         img_data_24_15 : IN std_logic ;
         img_data_24_14 : IN std_logic ;
         img_data_24_13 : IN std_logic ;
         img_data_24_12 : IN std_logic ;
         img_data_24_11 : IN std_logic ;
         img_data_24_10 : IN std_logic ;
         img_data_24_9 : IN std_logic ;
         img_data_24_8 : IN std_logic ;
         img_data_24_7 : IN std_logic ;
         img_data_24_6 : IN std_logic ;
         img_data_24_5 : IN std_logic ;
         img_data_24_4 : IN std_logic ;
         img_data_24_3 : IN std_logic ;
         img_data_24_2 : IN std_logic ;
         img_data_24_1 : IN std_logic ;
         img_data_24_0 : IN std_logic ;
         filter_data_0_31 : IN std_logic ;
         filter_data_0_30 : IN std_logic ;
         filter_data_0_29 : IN std_logic ;
         filter_data_0_28 : IN std_logic ;
         filter_data_0_27 : IN std_logic ;
         filter_data_0_26 : IN std_logic ;
         filter_data_0_25 : IN std_logic ;
         filter_data_0_24 : IN std_logic ;
         filter_data_0_23 : IN std_logic ;
         filter_data_0_22 : IN std_logic ;
         filter_data_0_21 : IN std_logic ;
         filter_data_0_20 : IN std_logic ;
         filter_data_0_19 : IN std_logic ;
         filter_data_0_18 : IN std_logic ;
         filter_data_0_17 : IN std_logic ;
         filter_data_0_16 : IN std_logic ;
         filter_data_0_15 : IN std_logic ;
         filter_data_0_14 : IN std_logic ;
         filter_data_0_13 : IN std_logic ;
         filter_data_0_12 : IN std_logic ;
         filter_data_0_11 : IN std_logic ;
         filter_data_0_10 : IN std_logic ;
         filter_data_0_9 : IN std_logic ;
         filter_data_0_8 : IN std_logic ;
         filter_data_0_7 : IN std_logic ;
         filter_data_0_6 : IN std_logic ;
         filter_data_0_5 : IN std_logic ;
         filter_data_0_4 : IN std_logic ;
         filter_data_0_3 : IN std_logic ;
         filter_data_0_2 : IN std_logic ;
         filter_data_0_1 : IN std_logic ;
         filter_data_0_0 : IN std_logic ;
         filter_data_1_31 : IN std_logic ;
         filter_data_1_30 : IN std_logic ;
         filter_data_1_29 : IN std_logic ;
         filter_data_1_28 : IN std_logic ;
         filter_data_1_27 : IN std_logic ;
         filter_data_1_26 : IN std_logic ;
         filter_data_1_25 : IN std_logic ;
         filter_data_1_24 : IN std_logic ;
         filter_data_1_23 : IN std_logic ;
         filter_data_1_22 : IN std_logic ;
         filter_data_1_21 : IN std_logic ;
         filter_data_1_20 : IN std_logic ;
         filter_data_1_19 : IN std_logic ;
         filter_data_1_18 : IN std_logic ;
         filter_data_1_17 : IN std_logic ;
         filter_data_1_16 : IN std_logic ;
         filter_data_1_15 : IN std_logic ;
         filter_data_1_14 : IN std_logic ;
         filter_data_1_13 : IN std_logic ;
         filter_data_1_12 : IN std_logic ;
         filter_data_1_11 : IN std_logic ;
         filter_data_1_10 : IN std_logic ;
         filter_data_1_9 : IN std_logic ;
         filter_data_1_8 : IN std_logic ;
         filter_data_1_7 : IN std_logic ;
         filter_data_1_6 : IN std_logic ;
         filter_data_1_5 : IN std_logic ;
         filter_data_1_4 : IN std_logic ;
         filter_data_1_3 : IN std_logic ;
         filter_data_1_2 : IN std_logic ;
         filter_data_1_1 : IN std_logic ;
         filter_data_1_0 : IN std_logic ;
         filter_data_2_31 : IN std_logic ;
         filter_data_2_30 : IN std_logic ;
         filter_data_2_29 : IN std_logic ;
         filter_data_2_28 : IN std_logic ;
         filter_data_2_27 : IN std_logic ;
         filter_data_2_26 : IN std_logic ;
         filter_data_2_25 : IN std_logic ;
         filter_data_2_24 : IN std_logic ;
         filter_data_2_23 : IN std_logic ;
         filter_data_2_22 : IN std_logic ;
         filter_data_2_21 : IN std_logic ;
         filter_data_2_20 : IN std_logic ;
         filter_data_2_19 : IN std_logic ;
         filter_data_2_18 : IN std_logic ;
         filter_data_2_17 : IN std_logic ;
         filter_data_2_16 : IN std_logic ;
         filter_data_2_15 : IN std_logic ;
         filter_data_2_14 : IN std_logic ;
         filter_data_2_13 : IN std_logic ;
         filter_data_2_12 : IN std_logic ;
         filter_data_2_11 : IN std_logic ;
         filter_data_2_10 : IN std_logic ;
         filter_data_2_9 : IN std_logic ;
         filter_data_2_8 : IN std_logic ;
         filter_data_2_7 : IN std_logic ;
         filter_data_2_6 : IN std_logic ;
         filter_data_2_5 : IN std_logic ;
         filter_data_2_4 : IN std_logic ;
         filter_data_2_3 : IN std_logic ;
         filter_data_2_2 : IN std_logic ;
         filter_data_2_1 : IN std_logic ;
         filter_data_2_0 : IN std_logic ;
         filter_data_3_31 : IN std_logic ;
         filter_data_3_30 : IN std_logic ;
         filter_data_3_29 : IN std_logic ;
         filter_data_3_28 : IN std_logic ;
         filter_data_3_27 : IN std_logic ;
         filter_data_3_26 : IN std_logic ;
         filter_data_3_25 : IN std_logic ;
         filter_data_3_24 : IN std_logic ;
         filter_data_3_23 : IN std_logic ;
         filter_data_3_22 : IN std_logic ;
         filter_data_3_21 : IN std_logic ;
         filter_data_3_20 : IN std_logic ;
         filter_data_3_19 : IN std_logic ;
         filter_data_3_18 : IN std_logic ;
         filter_data_3_17 : IN std_logic ;
         filter_data_3_16 : IN std_logic ;
         filter_data_3_15 : IN std_logic ;
         filter_data_3_14 : IN std_logic ;
         filter_data_3_13 : IN std_logic ;
         filter_data_3_12 : IN std_logic ;
         filter_data_3_11 : IN std_logic ;
         filter_data_3_10 : IN std_logic ;
         filter_data_3_9 : IN std_logic ;
         filter_data_3_8 : IN std_logic ;
         filter_data_3_7 : IN std_logic ;
         filter_data_3_6 : IN std_logic ;
         filter_data_3_5 : IN std_logic ;
         filter_data_3_4 : IN std_logic ;
         filter_data_3_3 : IN std_logic ;
         filter_data_3_2 : IN std_logic ;
         filter_data_3_1 : IN std_logic ;
         filter_data_3_0 : IN std_logic ;
         filter_data_4_31 : IN std_logic ;
         filter_data_4_30 : IN std_logic ;
         filter_data_4_29 : IN std_logic ;
         filter_data_4_28 : IN std_logic ;
         filter_data_4_27 : IN std_logic ;
         filter_data_4_26 : IN std_logic ;
         filter_data_4_25 : IN std_logic ;
         filter_data_4_24 : IN std_logic ;
         filter_data_4_23 : IN std_logic ;
         filter_data_4_22 : IN std_logic ;
         filter_data_4_21 : IN std_logic ;
         filter_data_4_20 : IN std_logic ;
         filter_data_4_19 : IN std_logic ;
         filter_data_4_18 : IN std_logic ;
         filter_data_4_17 : IN std_logic ;
         filter_data_4_16 : IN std_logic ;
         filter_data_4_15 : IN std_logic ;
         filter_data_4_14 : IN std_logic ;
         filter_data_4_13 : IN std_logic ;
         filter_data_4_12 : IN std_logic ;
         filter_data_4_11 : IN std_logic ;
         filter_data_4_10 : IN std_logic ;
         filter_data_4_9 : IN std_logic ;
         filter_data_4_8 : IN std_logic ;
         filter_data_4_7 : IN std_logic ;
         filter_data_4_6 : IN std_logic ;
         filter_data_4_5 : IN std_logic ;
         filter_data_4_4 : IN std_logic ;
         filter_data_4_3 : IN std_logic ;
         filter_data_4_2 : IN std_logic ;
         filter_data_4_1 : IN std_logic ;
         filter_data_4_0 : IN std_logic ;
         filter_data_5_31 : IN std_logic ;
         filter_data_5_30 : IN std_logic ;
         filter_data_5_29 : IN std_logic ;
         filter_data_5_28 : IN std_logic ;
         filter_data_5_27 : IN std_logic ;
         filter_data_5_26 : IN std_logic ;
         filter_data_5_25 : IN std_logic ;
         filter_data_5_24 : IN std_logic ;
         filter_data_5_23 : IN std_logic ;
         filter_data_5_22 : IN std_logic ;
         filter_data_5_21 : IN std_logic ;
         filter_data_5_20 : IN std_logic ;
         filter_data_5_19 : IN std_logic ;
         filter_data_5_18 : IN std_logic ;
         filter_data_5_17 : IN std_logic ;
         filter_data_5_16 : IN std_logic ;
         filter_data_5_15 : IN std_logic ;
         filter_data_5_14 : IN std_logic ;
         filter_data_5_13 : IN std_logic ;
         filter_data_5_12 : IN std_logic ;
         filter_data_5_11 : IN std_logic ;
         filter_data_5_10 : IN std_logic ;
         filter_data_5_9 : IN std_logic ;
         filter_data_5_8 : IN std_logic ;
         filter_data_5_7 : IN std_logic ;
         filter_data_5_6 : IN std_logic ;
         filter_data_5_5 : IN std_logic ;
         filter_data_5_4 : IN std_logic ;
         filter_data_5_3 : IN std_logic ;
         filter_data_5_2 : IN std_logic ;
         filter_data_5_1 : IN std_logic ;
         filter_data_5_0 : IN std_logic ;
         filter_data_6_31 : IN std_logic ;
         filter_data_6_30 : IN std_logic ;
         filter_data_6_29 : IN std_logic ;
         filter_data_6_28 : IN std_logic ;
         filter_data_6_27 : IN std_logic ;
         filter_data_6_26 : IN std_logic ;
         filter_data_6_25 : IN std_logic ;
         filter_data_6_24 : IN std_logic ;
         filter_data_6_23 : IN std_logic ;
         filter_data_6_22 : IN std_logic ;
         filter_data_6_21 : IN std_logic ;
         filter_data_6_20 : IN std_logic ;
         filter_data_6_19 : IN std_logic ;
         filter_data_6_18 : IN std_logic ;
         filter_data_6_17 : IN std_logic ;
         filter_data_6_16 : IN std_logic ;
         filter_data_6_15 : IN std_logic ;
         filter_data_6_14 : IN std_logic ;
         filter_data_6_13 : IN std_logic ;
         filter_data_6_12 : IN std_logic ;
         filter_data_6_11 : IN std_logic ;
         filter_data_6_10 : IN std_logic ;
         filter_data_6_9 : IN std_logic ;
         filter_data_6_8 : IN std_logic ;
         filter_data_6_7 : IN std_logic ;
         filter_data_6_6 : IN std_logic ;
         filter_data_6_5 : IN std_logic ;
         filter_data_6_4 : IN std_logic ;
         filter_data_6_3 : IN std_logic ;
         filter_data_6_2 : IN std_logic ;
         filter_data_6_1 : IN std_logic ;
         filter_data_6_0 : IN std_logic ;
         filter_data_7_31 : IN std_logic ;
         filter_data_7_30 : IN std_logic ;
         filter_data_7_29 : IN std_logic ;
         filter_data_7_28 : IN std_logic ;
         filter_data_7_27 : IN std_logic ;
         filter_data_7_26 : IN std_logic ;
         filter_data_7_25 : IN std_logic ;
         filter_data_7_24 : IN std_logic ;
         filter_data_7_23 : IN std_logic ;
         filter_data_7_22 : IN std_logic ;
         filter_data_7_21 : IN std_logic ;
         filter_data_7_20 : IN std_logic ;
         filter_data_7_19 : IN std_logic ;
         filter_data_7_18 : IN std_logic ;
         filter_data_7_17 : IN std_logic ;
         filter_data_7_16 : IN std_logic ;
         filter_data_7_15 : IN std_logic ;
         filter_data_7_14 : IN std_logic ;
         filter_data_7_13 : IN std_logic ;
         filter_data_7_12 : IN std_logic ;
         filter_data_7_11 : IN std_logic ;
         filter_data_7_10 : IN std_logic ;
         filter_data_7_9 : IN std_logic ;
         filter_data_7_8 : IN std_logic ;
         filter_data_7_7 : IN std_logic ;
         filter_data_7_6 : IN std_logic ;
         filter_data_7_5 : IN std_logic ;
         filter_data_7_4 : IN std_logic ;
         filter_data_7_3 : IN std_logic ;
         filter_data_7_2 : IN std_logic ;
         filter_data_7_1 : IN std_logic ;
         filter_data_7_0 : IN std_logic ;
         filter_data_8_31 : IN std_logic ;
         filter_data_8_30 : IN std_logic ;
         filter_data_8_29 : IN std_logic ;
         filter_data_8_28 : IN std_logic ;
         filter_data_8_27 : IN std_logic ;
         filter_data_8_26 : IN std_logic ;
         filter_data_8_25 : IN std_logic ;
         filter_data_8_24 : IN std_logic ;
         filter_data_8_23 : IN std_logic ;
         filter_data_8_22 : IN std_logic ;
         filter_data_8_21 : IN std_logic ;
         filter_data_8_20 : IN std_logic ;
         filter_data_8_19 : IN std_logic ;
         filter_data_8_18 : IN std_logic ;
         filter_data_8_17 : IN std_logic ;
         filter_data_8_16 : IN std_logic ;
         filter_data_8_15 : IN std_logic ;
         filter_data_8_14 : IN std_logic ;
         filter_data_8_13 : IN std_logic ;
         filter_data_8_12 : IN std_logic ;
         filter_data_8_11 : IN std_logic ;
         filter_data_8_10 : IN std_logic ;
         filter_data_8_9 : IN std_logic ;
         filter_data_8_8 : IN std_logic ;
         filter_data_8_7 : IN std_logic ;
         filter_data_8_6 : IN std_logic ;
         filter_data_8_5 : IN std_logic ;
         filter_data_8_4 : IN std_logic ;
         filter_data_8_3 : IN std_logic ;
         filter_data_8_2 : IN std_logic ;
         filter_data_8_1 : IN std_logic ;
         filter_data_8_0 : IN std_logic ;
         filter_data_9_31 : IN std_logic ;
         filter_data_9_30 : IN std_logic ;
         filter_data_9_29 : IN std_logic ;
         filter_data_9_28 : IN std_logic ;
         filter_data_9_27 : IN std_logic ;
         filter_data_9_26 : IN std_logic ;
         filter_data_9_25 : IN std_logic ;
         filter_data_9_24 : IN std_logic ;
         filter_data_9_23 : IN std_logic ;
         filter_data_9_22 : IN std_logic ;
         filter_data_9_21 : IN std_logic ;
         filter_data_9_20 : IN std_logic ;
         filter_data_9_19 : IN std_logic ;
         filter_data_9_18 : IN std_logic ;
         filter_data_9_17 : IN std_logic ;
         filter_data_9_16 : IN std_logic ;
         filter_data_9_15 : IN std_logic ;
         filter_data_9_14 : IN std_logic ;
         filter_data_9_13 : IN std_logic ;
         filter_data_9_12 : IN std_logic ;
         filter_data_9_11 : IN std_logic ;
         filter_data_9_10 : IN std_logic ;
         filter_data_9_9 : IN std_logic ;
         filter_data_9_8 : IN std_logic ;
         filter_data_9_7 : IN std_logic ;
         filter_data_9_6 : IN std_logic ;
         filter_data_9_5 : IN std_logic ;
         filter_data_9_4 : IN std_logic ;
         filter_data_9_3 : IN std_logic ;
         filter_data_9_2 : IN std_logic ;
         filter_data_9_1 : IN std_logic ;
         filter_data_9_0 : IN std_logic ;
         filter_data_10_31 : IN std_logic ;
         filter_data_10_30 : IN std_logic ;
         filter_data_10_29 : IN std_logic ;
         filter_data_10_28 : IN std_logic ;
         filter_data_10_27 : IN std_logic ;
         filter_data_10_26 : IN std_logic ;
         filter_data_10_25 : IN std_logic ;
         filter_data_10_24 : IN std_logic ;
         filter_data_10_23 : IN std_logic ;
         filter_data_10_22 : IN std_logic ;
         filter_data_10_21 : IN std_logic ;
         filter_data_10_20 : IN std_logic ;
         filter_data_10_19 : IN std_logic ;
         filter_data_10_18 : IN std_logic ;
         filter_data_10_17 : IN std_logic ;
         filter_data_10_16 : IN std_logic ;
         filter_data_10_15 : IN std_logic ;
         filter_data_10_14 : IN std_logic ;
         filter_data_10_13 : IN std_logic ;
         filter_data_10_12 : IN std_logic ;
         filter_data_10_11 : IN std_logic ;
         filter_data_10_10 : IN std_logic ;
         filter_data_10_9 : IN std_logic ;
         filter_data_10_8 : IN std_logic ;
         filter_data_10_7 : IN std_logic ;
         filter_data_10_6 : IN std_logic ;
         filter_data_10_5 : IN std_logic ;
         filter_data_10_4 : IN std_logic ;
         filter_data_10_3 : IN std_logic ;
         filter_data_10_2 : IN std_logic ;
         filter_data_10_1 : IN std_logic ;
         filter_data_10_0 : IN std_logic ;
         filter_data_11_31 : IN std_logic ;
         filter_data_11_30 : IN std_logic ;
         filter_data_11_29 : IN std_logic ;
         filter_data_11_28 : IN std_logic ;
         filter_data_11_27 : IN std_logic ;
         filter_data_11_26 : IN std_logic ;
         filter_data_11_25 : IN std_logic ;
         filter_data_11_24 : IN std_logic ;
         filter_data_11_23 : IN std_logic ;
         filter_data_11_22 : IN std_logic ;
         filter_data_11_21 : IN std_logic ;
         filter_data_11_20 : IN std_logic ;
         filter_data_11_19 : IN std_logic ;
         filter_data_11_18 : IN std_logic ;
         filter_data_11_17 : IN std_logic ;
         filter_data_11_16 : IN std_logic ;
         filter_data_11_15 : IN std_logic ;
         filter_data_11_14 : IN std_logic ;
         filter_data_11_13 : IN std_logic ;
         filter_data_11_12 : IN std_logic ;
         filter_data_11_11 : IN std_logic ;
         filter_data_11_10 : IN std_logic ;
         filter_data_11_9 : IN std_logic ;
         filter_data_11_8 : IN std_logic ;
         filter_data_11_7 : IN std_logic ;
         filter_data_11_6 : IN std_logic ;
         filter_data_11_5 : IN std_logic ;
         filter_data_11_4 : IN std_logic ;
         filter_data_11_3 : IN std_logic ;
         filter_data_11_2 : IN std_logic ;
         filter_data_11_1 : IN std_logic ;
         filter_data_11_0 : IN std_logic ;
         filter_data_12_31 : IN std_logic ;
         filter_data_12_30 : IN std_logic ;
         filter_data_12_29 : IN std_logic ;
         filter_data_12_28 : IN std_logic ;
         filter_data_12_27 : IN std_logic ;
         filter_data_12_26 : IN std_logic ;
         filter_data_12_25 : IN std_logic ;
         filter_data_12_24 : IN std_logic ;
         filter_data_12_23 : IN std_logic ;
         filter_data_12_22 : IN std_logic ;
         filter_data_12_21 : IN std_logic ;
         filter_data_12_20 : IN std_logic ;
         filter_data_12_19 : IN std_logic ;
         filter_data_12_18 : IN std_logic ;
         filter_data_12_17 : IN std_logic ;
         filter_data_12_16 : IN std_logic ;
         filter_data_12_15 : IN std_logic ;
         filter_data_12_14 : IN std_logic ;
         filter_data_12_13 : IN std_logic ;
         filter_data_12_12 : IN std_logic ;
         filter_data_12_11 : IN std_logic ;
         filter_data_12_10 : IN std_logic ;
         filter_data_12_9 : IN std_logic ;
         filter_data_12_8 : IN std_logic ;
         filter_data_12_7 : IN std_logic ;
         filter_data_12_6 : IN std_logic ;
         filter_data_12_5 : IN std_logic ;
         filter_data_12_4 : IN std_logic ;
         filter_data_12_3 : IN std_logic ;
         filter_data_12_2 : IN std_logic ;
         filter_data_12_1 : IN std_logic ;
         filter_data_12_0 : IN std_logic ;
         filter_data_13_31 : IN std_logic ;
         filter_data_13_30 : IN std_logic ;
         filter_data_13_29 : IN std_logic ;
         filter_data_13_28 : IN std_logic ;
         filter_data_13_27 : IN std_logic ;
         filter_data_13_26 : IN std_logic ;
         filter_data_13_25 : IN std_logic ;
         filter_data_13_24 : IN std_logic ;
         filter_data_13_23 : IN std_logic ;
         filter_data_13_22 : IN std_logic ;
         filter_data_13_21 : IN std_logic ;
         filter_data_13_20 : IN std_logic ;
         filter_data_13_19 : IN std_logic ;
         filter_data_13_18 : IN std_logic ;
         filter_data_13_17 : IN std_logic ;
         filter_data_13_16 : IN std_logic ;
         filter_data_13_15 : IN std_logic ;
         filter_data_13_14 : IN std_logic ;
         filter_data_13_13 : IN std_logic ;
         filter_data_13_12 : IN std_logic ;
         filter_data_13_11 : IN std_logic ;
         filter_data_13_10 : IN std_logic ;
         filter_data_13_9 : IN std_logic ;
         filter_data_13_8 : IN std_logic ;
         filter_data_13_7 : IN std_logic ;
         filter_data_13_6 : IN std_logic ;
         filter_data_13_5 : IN std_logic ;
         filter_data_13_4 : IN std_logic ;
         filter_data_13_3 : IN std_logic ;
         filter_data_13_2 : IN std_logic ;
         filter_data_13_1 : IN std_logic ;
         filter_data_13_0 : IN std_logic ;
         filter_data_14_31 : IN std_logic ;
         filter_data_14_30 : IN std_logic ;
         filter_data_14_29 : IN std_logic ;
         filter_data_14_28 : IN std_logic ;
         filter_data_14_27 : IN std_logic ;
         filter_data_14_26 : IN std_logic ;
         filter_data_14_25 : IN std_logic ;
         filter_data_14_24 : IN std_logic ;
         filter_data_14_23 : IN std_logic ;
         filter_data_14_22 : IN std_logic ;
         filter_data_14_21 : IN std_logic ;
         filter_data_14_20 : IN std_logic ;
         filter_data_14_19 : IN std_logic ;
         filter_data_14_18 : IN std_logic ;
         filter_data_14_17 : IN std_logic ;
         filter_data_14_16 : IN std_logic ;
         filter_data_14_15 : IN std_logic ;
         filter_data_14_14 : IN std_logic ;
         filter_data_14_13 : IN std_logic ;
         filter_data_14_12 : IN std_logic ;
         filter_data_14_11 : IN std_logic ;
         filter_data_14_10 : IN std_logic ;
         filter_data_14_9 : IN std_logic ;
         filter_data_14_8 : IN std_logic ;
         filter_data_14_7 : IN std_logic ;
         filter_data_14_6 : IN std_logic ;
         filter_data_14_5 : IN std_logic ;
         filter_data_14_4 : IN std_logic ;
         filter_data_14_3 : IN std_logic ;
         filter_data_14_2 : IN std_logic ;
         filter_data_14_1 : IN std_logic ;
         filter_data_14_0 : IN std_logic ;
         filter_data_15_31 : IN std_logic ;
         filter_data_15_30 : IN std_logic ;
         filter_data_15_29 : IN std_logic ;
         filter_data_15_28 : IN std_logic ;
         filter_data_15_27 : IN std_logic ;
         filter_data_15_26 : IN std_logic ;
         filter_data_15_25 : IN std_logic ;
         filter_data_15_24 : IN std_logic ;
         filter_data_15_23 : IN std_logic ;
         filter_data_15_22 : IN std_logic ;
         filter_data_15_21 : IN std_logic ;
         filter_data_15_20 : IN std_logic ;
         filter_data_15_19 : IN std_logic ;
         filter_data_15_18 : IN std_logic ;
         filter_data_15_17 : IN std_logic ;
         filter_data_15_16 : IN std_logic ;
         filter_data_15_15 : IN std_logic ;
         filter_data_15_14 : IN std_logic ;
         filter_data_15_13 : IN std_logic ;
         filter_data_15_12 : IN std_logic ;
         filter_data_15_11 : IN std_logic ;
         filter_data_15_10 : IN std_logic ;
         filter_data_15_9 : IN std_logic ;
         filter_data_15_8 : IN std_logic ;
         filter_data_15_7 : IN std_logic ;
         filter_data_15_6 : IN std_logic ;
         filter_data_15_5 : IN std_logic ;
         filter_data_15_4 : IN std_logic ;
         filter_data_15_3 : IN std_logic ;
         filter_data_15_2 : IN std_logic ;
         filter_data_15_1 : IN std_logic ;
         filter_data_15_0 : IN std_logic ;
         filter_data_16_31 : IN std_logic ;
         filter_data_16_30 : IN std_logic ;
         filter_data_16_29 : IN std_logic ;
         filter_data_16_28 : IN std_logic ;
         filter_data_16_27 : IN std_logic ;
         filter_data_16_26 : IN std_logic ;
         filter_data_16_25 : IN std_logic ;
         filter_data_16_24 : IN std_logic ;
         filter_data_16_23 : IN std_logic ;
         filter_data_16_22 : IN std_logic ;
         filter_data_16_21 : IN std_logic ;
         filter_data_16_20 : IN std_logic ;
         filter_data_16_19 : IN std_logic ;
         filter_data_16_18 : IN std_logic ;
         filter_data_16_17 : IN std_logic ;
         filter_data_16_16 : IN std_logic ;
         filter_data_16_15 : IN std_logic ;
         filter_data_16_14 : IN std_logic ;
         filter_data_16_13 : IN std_logic ;
         filter_data_16_12 : IN std_logic ;
         filter_data_16_11 : IN std_logic ;
         filter_data_16_10 : IN std_logic ;
         filter_data_16_9 : IN std_logic ;
         filter_data_16_8 : IN std_logic ;
         filter_data_16_7 : IN std_logic ;
         filter_data_16_6 : IN std_logic ;
         filter_data_16_5 : IN std_logic ;
         filter_data_16_4 : IN std_logic ;
         filter_data_16_3 : IN std_logic ;
         filter_data_16_2 : IN std_logic ;
         filter_data_16_1 : IN std_logic ;
         filter_data_16_0 : IN std_logic ;
         filter_data_17_31 : IN std_logic ;
         filter_data_17_30 : IN std_logic ;
         filter_data_17_29 : IN std_logic ;
         filter_data_17_28 : IN std_logic ;
         filter_data_17_27 : IN std_logic ;
         filter_data_17_26 : IN std_logic ;
         filter_data_17_25 : IN std_logic ;
         filter_data_17_24 : IN std_logic ;
         filter_data_17_23 : IN std_logic ;
         filter_data_17_22 : IN std_logic ;
         filter_data_17_21 : IN std_logic ;
         filter_data_17_20 : IN std_logic ;
         filter_data_17_19 : IN std_logic ;
         filter_data_17_18 : IN std_logic ;
         filter_data_17_17 : IN std_logic ;
         filter_data_17_16 : IN std_logic ;
         filter_data_17_15 : IN std_logic ;
         filter_data_17_14 : IN std_logic ;
         filter_data_17_13 : IN std_logic ;
         filter_data_17_12 : IN std_logic ;
         filter_data_17_11 : IN std_logic ;
         filter_data_17_10 : IN std_logic ;
         filter_data_17_9 : IN std_logic ;
         filter_data_17_8 : IN std_logic ;
         filter_data_17_7 : IN std_logic ;
         filter_data_17_6 : IN std_logic ;
         filter_data_17_5 : IN std_logic ;
         filter_data_17_4 : IN std_logic ;
         filter_data_17_3 : IN std_logic ;
         filter_data_17_2 : IN std_logic ;
         filter_data_17_1 : IN std_logic ;
         filter_data_17_0 : IN std_logic ;
         filter_data_18_31 : IN std_logic ;
         filter_data_18_30 : IN std_logic ;
         filter_data_18_29 : IN std_logic ;
         filter_data_18_28 : IN std_logic ;
         filter_data_18_27 : IN std_logic ;
         filter_data_18_26 : IN std_logic ;
         filter_data_18_25 : IN std_logic ;
         filter_data_18_24 : IN std_logic ;
         filter_data_18_23 : IN std_logic ;
         filter_data_18_22 : IN std_logic ;
         filter_data_18_21 : IN std_logic ;
         filter_data_18_20 : IN std_logic ;
         filter_data_18_19 : IN std_logic ;
         filter_data_18_18 : IN std_logic ;
         filter_data_18_17 : IN std_logic ;
         filter_data_18_16 : IN std_logic ;
         filter_data_18_15 : IN std_logic ;
         filter_data_18_14 : IN std_logic ;
         filter_data_18_13 : IN std_logic ;
         filter_data_18_12 : IN std_logic ;
         filter_data_18_11 : IN std_logic ;
         filter_data_18_10 : IN std_logic ;
         filter_data_18_9 : IN std_logic ;
         filter_data_18_8 : IN std_logic ;
         filter_data_18_7 : IN std_logic ;
         filter_data_18_6 : IN std_logic ;
         filter_data_18_5 : IN std_logic ;
         filter_data_18_4 : IN std_logic ;
         filter_data_18_3 : IN std_logic ;
         filter_data_18_2 : IN std_logic ;
         filter_data_18_1 : IN std_logic ;
         filter_data_18_0 : IN std_logic ;
         filter_data_19_31 : IN std_logic ;
         filter_data_19_30 : IN std_logic ;
         filter_data_19_29 : IN std_logic ;
         filter_data_19_28 : IN std_logic ;
         filter_data_19_27 : IN std_logic ;
         filter_data_19_26 : IN std_logic ;
         filter_data_19_25 : IN std_logic ;
         filter_data_19_24 : IN std_logic ;
         filter_data_19_23 : IN std_logic ;
         filter_data_19_22 : IN std_logic ;
         filter_data_19_21 : IN std_logic ;
         filter_data_19_20 : IN std_logic ;
         filter_data_19_19 : IN std_logic ;
         filter_data_19_18 : IN std_logic ;
         filter_data_19_17 : IN std_logic ;
         filter_data_19_16 : IN std_logic ;
         filter_data_19_15 : IN std_logic ;
         filter_data_19_14 : IN std_logic ;
         filter_data_19_13 : IN std_logic ;
         filter_data_19_12 : IN std_logic ;
         filter_data_19_11 : IN std_logic ;
         filter_data_19_10 : IN std_logic ;
         filter_data_19_9 : IN std_logic ;
         filter_data_19_8 : IN std_logic ;
         filter_data_19_7 : IN std_logic ;
         filter_data_19_6 : IN std_logic ;
         filter_data_19_5 : IN std_logic ;
         filter_data_19_4 : IN std_logic ;
         filter_data_19_3 : IN std_logic ;
         filter_data_19_2 : IN std_logic ;
         filter_data_19_1 : IN std_logic ;
         filter_data_19_0 : IN std_logic ;
         filter_data_20_31 : IN std_logic ;
         filter_data_20_30 : IN std_logic ;
         filter_data_20_29 : IN std_logic ;
         filter_data_20_28 : IN std_logic ;
         filter_data_20_27 : IN std_logic ;
         filter_data_20_26 : IN std_logic ;
         filter_data_20_25 : IN std_logic ;
         filter_data_20_24 : IN std_logic ;
         filter_data_20_23 : IN std_logic ;
         filter_data_20_22 : IN std_logic ;
         filter_data_20_21 : IN std_logic ;
         filter_data_20_20 : IN std_logic ;
         filter_data_20_19 : IN std_logic ;
         filter_data_20_18 : IN std_logic ;
         filter_data_20_17 : IN std_logic ;
         filter_data_20_16 : IN std_logic ;
         filter_data_20_15 : IN std_logic ;
         filter_data_20_14 : IN std_logic ;
         filter_data_20_13 : IN std_logic ;
         filter_data_20_12 : IN std_logic ;
         filter_data_20_11 : IN std_logic ;
         filter_data_20_10 : IN std_logic ;
         filter_data_20_9 : IN std_logic ;
         filter_data_20_8 : IN std_logic ;
         filter_data_20_7 : IN std_logic ;
         filter_data_20_6 : IN std_logic ;
         filter_data_20_5 : IN std_logic ;
         filter_data_20_4 : IN std_logic ;
         filter_data_20_3 : IN std_logic ;
         filter_data_20_2 : IN std_logic ;
         filter_data_20_1 : IN std_logic ;
         filter_data_20_0 : IN std_logic ;
         filter_data_21_31 : IN std_logic ;
         filter_data_21_30 : IN std_logic ;
         filter_data_21_29 : IN std_logic ;
         filter_data_21_28 : IN std_logic ;
         filter_data_21_27 : IN std_logic ;
         filter_data_21_26 : IN std_logic ;
         filter_data_21_25 : IN std_logic ;
         filter_data_21_24 : IN std_logic ;
         filter_data_21_23 : IN std_logic ;
         filter_data_21_22 : IN std_logic ;
         filter_data_21_21 : IN std_logic ;
         filter_data_21_20 : IN std_logic ;
         filter_data_21_19 : IN std_logic ;
         filter_data_21_18 : IN std_logic ;
         filter_data_21_17 : IN std_logic ;
         filter_data_21_16 : IN std_logic ;
         filter_data_21_15 : IN std_logic ;
         filter_data_21_14 : IN std_logic ;
         filter_data_21_13 : IN std_logic ;
         filter_data_21_12 : IN std_logic ;
         filter_data_21_11 : IN std_logic ;
         filter_data_21_10 : IN std_logic ;
         filter_data_21_9 : IN std_logic ;
         filter_data_21_8 : IN std_logic ;
         filter_data_21_7 : IN std_logic ;
         filter_data_21_6 : IN std_logic ;
         filter_data_21_5 : IN std_logic ;
         filter_data_21_4 : IN std_logic ;
         filter_data_21_3 : IN std_logic ;
         filter_data_21_2 : IN std_logic ;
         filter_data_21_1 : IN std_logic ;
         filter_data_21_0 : IN std_logic ;
         filter_data_22_31 : IN std_logic ;
         filter_data_22_30 : IN std_logic ;
         filter_data_22_29 : IN std_logic ;
         filter_data_22_28 : IN std_logic ;
         filter_data_22_27 : IN std_logic ;
         filter_data_22_26 : IN std_logic ;
         filter_data_22_25 : IN std_logic ;
         filter_data_22_24 : IN std_logic ;
         filter_data_22_23 : IN std_logic ;
         filter_data_22_22 : IN std_logic ;
         filter_data_22_21 : IN std_logic ;
         filter_data_22_20 : IN std_logic ;
         filter_data_22_19 : IN std_logic ;
         filter_data_22_18 : IN std_logic ;
         filter_data_22_17 : IN std_logic ;
         filter_data_22_16 : IN std_logic ;
         filter_data_22_15 : IN std_logic ;
         filter_data_22_14 : IN std_logic ;
         filter_data_22_13 : IN std_logic ;
         filter_data_22_12 : IN std_logic ;
         filter_data_22_11 : IN std_logic ;
         filter_data_22_10 : IN std_logic ;
         filter_data_22_9 : IN std_logic ;
         filter_data_22_8 : IN std_logic ;
         filter_data_22_7 : IN std_logic ;
         filter_data_22_6 : IN std_logic ;
         filter_data_22_5 : IN std_logic ;
         filter_data_22_4 : IN std_logic ;
         filter_data_22_3 : IN std_logic ;
         filter_data_22_2 : IN std_logic ;
         filter_data_22_1 : IN std_logic ;
         filter_data_22_0 : IN std_logic ;
         filter_data_23_31 : IN std_logic ;
         filter_data_23_30 : IN std_logic ;
         filter_data_23_29 : IN std_logic ;
         filter_data_23_28 : IN std_logic ;
         filter_data_23_27 : IN std_logic ;
         filter_data_23_26 : IN std_logic ;
         filter_data_23_25 : IN std_logic ;
         filter_data_23_24 : IN std_logic ;
         filter_data_23_23 : IN std_logic ;
         filter_data_23_22 : IN std_logic ;
         filter_data_23_21 : IN std_logic ;
         filter_data_23_20 : IN std_logic ;
         filter_data_23_19 : IN std_logic ;
         filter_data_23_18 : IN std_logic ;
         filter_data_23_17 : IN std_logic ;
         filter_data_23_16 : IN std_logic ;
         filter_data_23_15 : IN std_logic ;
         filter_data_23_14 : IN std_logic ;
         filter_data_23_13 : IN std_logic ;
         filter_data_23_12 : IN std_logic ;
         filter_data_23_11 : IN std_logic ;
         filter_data_23_10 : IN std_logic ;
         filter_data_23_9 : IN std_logic ;
         filter_data_23_8 : IN std_logic ;
         filter_data_23_7 : IN std_logic ;
         filter_data_23_6 : IN std_logic ;
         filter_data_23_5 : IN std_logic ;
         filter_data_23_4 : IN std_logic ;
         filter_data_23_3 : IN std_logic ;
         filter_data_23_2 : IN std_logic ;
         filter_data_23_1 : IN std_logic ;
         filter_data_23_0 : IN std_logic ;
         filter_data_24_31 : IN std_logic ;
         filter_data_24_30 : IN std_logic ;
         filter_data_24_29 : IN std_logic ;
         filter_data_24_28 : IN std_logic ;
         filter_data_24_27 : IN std_logic ;
         filter_data_24_26 : IN std_logic ;
         filter_data_24_25 : IN std_logic ;
         filter_data_24_24 : IN std_logic ;
         filter_data_24_23 : IN std_logic ;
         filter_data_24_22 : IN std_logic ;
         filter_data_24_21 : IN std_logic ;
         filter_data_24_20 : IN std_logic ;
         filter_data_24_19 : IN std_logic ;
         filter_data_24_18 : IN std_logic ;
         filter_data_24_17 : IN std_logic ;
         filter_data_24_16 : IN std_logic ;
         filter_data_24_15 : IN std_logic ;
         filter_data_24_14 : IN std_logic ;
         filter_data_24_13 : IN std_logic ;
         filter_data_24_12 : IN std_logic ;
         filter_data_24_11 : IN std_logic ;
         filter_data_24_10 : IN std_logic ;
         filter_data_24_9 : IN std_logic ;
         filter_data_24_8 : IN std_logic ;
         filter_data_24_7 : IN std_logic ;
         filter_data_24_6 : IN std_logic ;
         filter_data_24_5 : IN std_logic ;
         filter_data_24_4 : IN std_logic ;
         filter_data_24_3 : IN std_logic ;
         filter_data_24_2 : IN std_logic ;
         filter_data_24_1 : IN std_logic ;
         filter_data_24_0 : IN std_logic ;
         filter_size : IN std_logic ;
         ordered_img_data_0_31 : OUT std_logic ;
         ordered_img_data_0_30 : OUT std_logic ;
         ordered_img_data_0_29 : OUT std_logic ;
         ordered_img_data_0_28 : OUT std_logic ;
         ordered_img_data_0_27 : OUT std_logic ;
         ordered_img_data_0_26 : OUT std_logic ;
         ordered_img_data_0_25 : OUT std_logic ;
         ordered_img_data_0_24 : OUT std_logic ;
         ordered_img_data_0_23 : OUT std_logic ;
         ordered_img_data_0_22 : OUT std_logic ;
         ordered_img_data_0_21 : OUT std_logic ;
         ordered_img_data_0_20 : OUT std_logic ;
         ordered_img_data_0_19 : OUT std_logic ;
         ordered_img_data_0_18 : OUT std_logic ;
         ordered_img_data_0_17 : OUT std_logic ;
         ordered_img_data_0_16 : OUT std_logic ;
         ordered_img_data_0_15 : OUT std_logic ;
         ordered_img_data_0_14 : OUT std_logic ;
         ordered_img_data_0_13 : OUT std_logic ;
         ordered_img_data_0_12 : OUT std_logic ;
         ordered_img_data_0_11 : OUT std_logic ;
         ordered_img_data_0_10 : OUT std_logic ;
         ordered_img_data_0_9 : OUT std_logic ;
         ordered_img_data_0_8 : OUT std_logic ;
         ordered_img_data_0_7 : OUT std_logic ;
         ordered_img_data_0_6 : OUT std_logic ;
         ordered_img_data_0_5 : OUT std_logic ;
         ordered_img_data_0_4 : OUT std_logic ;
         ordered_img_data_0_3 : OUT std_logic ;
         ordered_img_data_0_2 : OUT std_logic ;
         ordered_img_data_0_1 : OUT std_logic ;
         ordered_img_data_0_0 : OUT std_logic ;
         ordered_img_data_1_31 : OUT std_logic ;
         ordered_img_data_1_30 : OUT std_logic ;
         ordered_img_data_1_29 : OUT std_logic ;
         ordered_img_data_1_28 : OUT std_logic ;
         ordered_img_data_1_27 : OUT std_logic ;
         ordered_img_data_1_26 : OUT std_logic ;
         ordered_img_data_1_25 : OUT std_logic ;
         ordered_img_data_1_24 : OUT std_logic ;
         ordered_img_data_1_23 : OUT std_logic ;
         ordered_img_data_1_22 : OUT std_logic ;
         ordered_img_data_1_21 : OUT std_logic ;
         ordered_img_data_1_20 : OUT std_logic ;
         ordered_img_data_1_19 : OUT std_logic ;
         ordered_img_data_1_18 : OUT std_logic ;
         ordered_img_data_1_17 : OUT std_logic ;
         ordered_img_data_1_16 : OUT std_logic ;
         ordered_img_data_1_15 : OUT std_logic ;
         ordered_img_data_1_14 : OUT std_logic ;
         ordered_img_data_1_13 : OUT std_logic ;
         ordered_img_data_1_12 : OUT std_logic ;
         ordered_img_data_1_11 : OUT std_logic ;
         ordered_img_data_1_10 : OUT std_logic ;
         ordered_img_data_1_9 : OUT std_logic ;
         ordered_img_data_1_8 : OUT std_logic ;
         ordered_img_data_1_7 : OUT std_logic ;
         ordered_img_data_1_6 : OUT std_logic ;
         ordered_img_data_1_5 : OUT std_logic ;
         ordered_img_data_1_4 : OUT std_logic ;
         ordered_img_data_1_3 : OUT std_logic ;
         ordered_img_data_1_2 : OUT std_logic ;
         ordered_img_data_1_1 : OUT std_logic ;
         ordered_img_data_1_0 : OUT std_logic ;
         ordered_img_data_2_31 : OUT std_logic ;
         ordered_img_data_2_30 : OUT std_logic ;
         ordered_img_data_2_29 : OUT std_logic ;
         ordered_img_data_2_28 : OUT std_logic ;
         ordered_img_data_2_27 : OUT std_logic ;
         ordered_img_data_2_26 : OUT std_logic ;
         ordered_img_data_2_25 : OUT std_logic ;
         ordered_img_data_2_24 : OUT std_logic ;
         ordered_img_data_2_23 : OUT std_logic ;
         ordered_img_data_2_22 : OUT std_logic ;
         ordered_img_data_2_21 : OUT std_logic ;
         ordered_img_data_2_20 : OUT std_logic ;
         ordered_img_data_2_19 : OUT std_logic ;
         ordered_img_data_2_18 : OUT std_logic ;
         ordered_img_data_2_17 : OUT std_logic ;
         ordered_img_data_2_16 : OUT std_logic ;
         ordered_img_data_2_15 : OUT std_logic ;
         ordered_img_data_2_14 : OUT std_logic ;
         ordered_img_data_2_13 : OUT std_logic ;
         ordered_img_data_2_12 : OUT std_logic ;
         ordered_img_data_2_11 : OUT std_logic ;
         ordered_img_data_2_10 : OUT std_logic ;
         ordered_img_data_2_9 : OUT std_logic ;
         ordered_img_data_2_8 : OUT std_logic ;
         ordered_img_data_2_7 : OUT std_logic ;
         ordered_img_data_2_6 : OUT std_logic ;
         ordered_img_data_2_5 : OUT std_logic ;
         ordered_img_data_2_4 : OUT std_logic ;
         ordered_img_data_2_3 : OUT std_logic ;
         ordered_img_data_2_2 : OUT std_logic ;
         ordered_img_data_2_1 : OUT std_logic ;
         ordered_img_data_2_0 : OUT std_logic ;
         ordered_img_data_3_31 : OUT std_logic ;
         ordered_img_data_3_30 : OUT std_logic ;
         ordered_img_data_3_29 : OUT std_logic ;
         ordered_img_data_3_28 : OUT std_logic ;
         ordered_img_data_3_27 : OUT std_logic ;
         ordered_img_data_3_26 : OUT std_logic ;
         ordered_img_data_3_25 : OUT std_logic ;
         ordered_img_data_3_24 : OUT std_logic ;
         ordered_img_data_3_23 : OUT std_logic ;
         ordered_img_data_3_22 : OUT std_logic ;
         ordered_img_data_3_21 : OUT std_logic ;
         ordered_img_data_3_20 : OUT std_logic ;
         ordered_img_data_3_19 : OUT std_logic ;
         ordered_img_data_3_18 : OUT std_logic ;
         ordered_img_data_3_17 : OUT std_logic ;
         ordered_img_data_3_16 : OUT std_logic ;
         ordered_img_data_3_15 : OUT std_logic ;
         ordered_img_data_3_14 : OUT std_logic ;
         ordered_img_data_3_13 : OUT std_logic ;
         ordered_img_data_3_12 : OUT std_logic ;
         ordered_img_data_3_11 : OUT std_logic ;
         ordered_img_data_3_10 : OUT std_logic ;
         ordered_img_data_3_9 : OUT std_logic ;
         ordered_img_data_3_8 : OUT std_logic ;
         ordered_img_data_3_7 : OUT std_logic ;
         ordered_img_data_3_6 : OUT std_logic ;
         ordered_img_data_3_5 : OUT std_logic ;
         ordered_img_data_3_4 : OUT std_logic ;
         ordered_img_data_3_3 : OUT std_logic ;
         ordered_img_data_3_2 : OUT std_logic ;
         ordered_img_data_3_1 : OUT std_logic ;
         ordered_img_data_3_0 : OUT std_logic ;
         ordered_img_data_4_31 : OUT std_logic ;
         ordered_img_data_4_30 : OUT std_logic ;
         ordered_img_data_4_29 : OUT std_logic ;
         ordered_img_data_4_28 : OUT std_logic ;
         ordered_img_data_4_27 : OUT std_logic ;
         ordered_img_data_4_26 : OUT std_logic ;
         ordered_img_data_4_25 : OUT std_logic ;
         ordered_img_data_4_24 : OUT std_logic ;
         ordered_img_data_4_23 : OUT std_logic ;
         ordered_img_data_4_22 : OUT std_logic ;
         ordered_img_data_4_21 : OUT std_logic ;
         ordered_img_data_4_20 : OUT std_logic ;
         ordered_img_data_4_19 : OUT std_logic ;
         ordered_img_data_4_18 : OUT std_logic ;
         ordered_img_data_4_17 : OUT std_logic ;
         ordered_img_data_4_16 : OUT std_logic ;
         ordered_img_data_4_15 : OUT std_logic ;
         ordered_img_data_4_14 : OUT std_logic ;
         ordered_img_data_4_13 : OUT std_logic ;
         ordered_img_data_4_12 : OUT std_logic ;
         ordered_img_data_4_11 : OUT std_logic ;
         ordered_img_data_4_10 : OUT std_logic ;
         ordered_img_data_4_9 : OUT std_logic ;
         ordered_img_data_4_8 : OUT std_logic ;
         ordered_img_data_4_7 : OUT std_logic ;
         ordered_img_data_4_6 : OUT std_logic ;
         ordered_img_data_4_5 : OUT std_logic ;
         ordered_img_data_4_4 : OUT std_logic ;
         ordered_img_data_4_3 : OUT std_logic ;
         ordered_img_data_4_2 : OUT std_logic ;
         ordered_img_data_4_1 : OUT std_logic ;
         ordered_img_data_4_0 : OUT std_logic ;
         ordered_img_data_5_31 : OUT std_logic ;
         ordered_img_data_5_30 : OUT std_logic ;
         ordered_img_data_5_29 : OUT std_logic ;
         ordered_img_data_5_28 : OUT std_logic ;
         ordered_img_data_5_27 : OUT std_logic ;
         ordered_img_data_5_26 : OUT std_logic ;
         ordered_img_data_5_25 : OUT std_logic ;
         ordered_img_data_5_24 : OUT std_logic ;
         ordered_img_data_5_23 : OUT std_logic ;
         ordered_img_data_5_22 : OUT std_logic ;
         ordered_img_data_5_21 : OUT std_logic ;
         ordered_img_data_5_20 : OUT std_logic ;
         ordered_img_data_5_19 : OUT std_logic ;
         ordered_img_data_5_18 : OUT std_logic ;
         ordered_img_data_5_17 : OUT std_logic ;
         ordered_img_data_5_16 : OUT std_logic ;
         ordered_img_data_5_15 : OUT std_logic ;
         ordered_img_data_5_14 : OUT std_logic ;
         ordered_img_data_5_13 : OUT std_logic ;
         ordered_img_data_5_12 : OUT std_logic ;
         ordered_img_data_5_11 : OUT std_logic ;
         ordered_img_data_5_10 : OUT std_logic ;
         ordered_img_data_5_9 : OUT std_logic ;
         ordered_img_data_5_8 : OUT std_logic ;
         ordered_img_data_5_7 : OUT std_logic ;
         ordered_img_data_5_6 : OUT std_logic ;
         ordered_img_data_5_5 : OUT std_logic ;
         ordered_img_data_5_4 : OUT std_logic ;
         ordered_img_data_5_3 : OUT std_logic ;
         ordered_img_data_5_2 : OUT std_logic ;
         ordered_img_data_5_1 : OUT std_logic ;
         ordered_img_data_5_0 : OUT std_logic ;
         ordered_img_data_6_31 : OUT std_logic ;
         ordered_img_data_6_30 : OUT std_logic ;
         ordered_img_data_6_29 : OUT std_logic ;
         ordered_img_data_6_28 : OUT std_logic ;
         ordered_img_data_6_27 : OUT std_logic ;
         ordered_img_data_6_26 : OUT std_logic ;
         ordered_img_data_6_25 : OUT std_logic ;
         ordered_img_data_6_24 : OUT std_logic ;
         ordered_img_data_6_23 : OUT std_logic ;
         ordered_img_data_6_22 : OUT std_logic ;
         ordered_img_data_6_21 : OUT std_logic ;
         ordered_img_data_6_20 : OUT std_logic ;
         ordered_img_data_6_19 : OUT std_logic ;
         ordered_img_data_6_18 : OUT std_logic ;
         ordered_img_data_6_17 : OUT std_logic ;
         ordered_img_data_6_16 : OUT std_logic ;
         ordered_img_data_6_15 : OUT std_logic ;
         ordered_img_data_6_14 : OUT std_logic ;
         ordered_img_data_6_13 : OUT std_logic ;
         ordered_img_data_6_12 : OUT std_logic ;
         ordered_img_data_6_11 : OUT std_logic ;
         ordered_img_data_6_10 : OUT std_logic ;
         ordered_img_data_6_9 : OUT std_logic ;
         ordered_img_data_6_8 : OUT std_logic ;
         ordered_img_data_6_7 : OUT std_logic ;
         ordered_img_data_6_6 : OUT std_logic ;
         ordered_img_data_6_5 : OUT std_logic ;
         ordered_img_data_6_4 : OUT std_logic ;
         ordered_img_data_6_3 : OUT std_logic ;
         ordered_img_data_6_2 : OUT std_logic ;
         ordered_img_data_6_1 : OUT std_logic ;
         ordered_img_data_6_0 : OUT std_logic ;
         ordered_img_data_7_31 : OUT std_logic ;
         ordered_img_data_7_30 : OUT std_logic ;
         ordered_img_data_7_29 : OUT std_logic ;
         ordered_img_data_7_28 : OUT std_logic ;
         ordered_img_data_7_27 : OUT std_logic ;
         ordered_img_data_7_26 : OUT std_logic ;
         ordered_img_data_7_25 : OUT std_logic ;
         ordered_img_data_7_24 : OUT std_logic ;
         ordered_img_data_7_23 : OUT std_logic ;
         ordered_img_data_7_22 : OUT std_logic ;
         ordered_img_data_7_21 : OUT std_logic ;
         ordered_img_data_7_20 : OUT std_logic ;
         ordered_img_data_7_19 : OUT std_logic ;
         ordered_img_data_7_18 : OUT std_logic ;
         ordered_img_data_7_17 : OUT std_logic ;
         ordered_img_data_7_16 : OUT std_logic ;
         ordered_img_data_7_15 : OUT std_logic ;
         ordered_img_data_7_14 : OUT std_logic ;
         ordered_img_data_7_13 : OUT std_logic ;
         ordered_img_data_7_12 : OUT std_logic ;
         ordered_img_data_7_11 : OUT std_logic ;
         ordered_img_data_7_10 : OUT std_logic ;
         ordered_img_data_7_9 : OUT std_logic ;
         ordered_img_data_7_8 : OUT std_logic ;
         ordered_img_data_7_7 : OUT std_logic ;
         ordered_img_data_7_6 : OUT std_logic ;
         ordered_img_data_7_5 : OUT std_logic ;
         ordered_img_data_7_4 : OUT std_logic ;
         ordered_img_data_7_3 : OUT std_logic ;
         ordered_img_data_7_2 : OUT std_logic ;
         ordered_img_data_7_1 : OUT std_logic ;
         ordered_img_data_7_0 : OUT std_logic ;
         ordered_img_data_8_31 : OUT std_logic ;
         ordered_img_data_8_30 : OUT std_logic ;
         ordered_img_data_8_29 : OUT std_logic ;
         ordered_img_data_8_28 : OUT std_logic ;
         ordered_img_data_8_27 : OUT std_logic ;
         ordered_img_data_8_26 : OUT std_logic ;
         ordered_img_data_8_25 : OUT std_logic ;
         ordered_img_data_8_24 : OUT std_logic ;
         ordered_img_data_8_23 : OUT std_logic ;
         ordered_img_data_8_22 : OUT std_logic ;
         ordered_img_data_8_21 : OUT std_logic ;
         ordered_img_data_8_20 : OUT std_logic ;
         ordered_img_data_8_19 : OUT std_logic ;
         ordered_img_data_8_18 : OUT std_logic ;
         ordered_img_data_8_17 : OUT std_logic ;
         ordered_img_data_8_16 : OUT std_logic ;
         ordered_img_data_8_15 : OUT std_logic ;
         ordered_img_data_8_14 : OUT std_logic ;
         ordered_img_data_8_13 : OUT std_logic ;
         ordered_img_data_8_12 : OUT std_logic ;
         ordered_img_data_8_11 : OUT std_logic ;
         ordered_img_data_8_10 : OUT std_logic ;
         ordered_img_data_8_9 : OUT std_logic ;
         ordered_img_data_8_8 : OUT std_logic ;
         ordered_img_data_8_7 : OUT std_logic ;
         ordered_img_data_8_6 : OUT std_logic ;
         ordered_img_data_8_5 : OUT std_logic ;
         ordered_img_data_8_4 : OUT std_logic ;
         ordered_img_data_8_3 : OUT std_logic ;
         ordered_img_data_8_2 : OUT std_logic ;
         ordered_img_data_8_1 : OUT std_logic ;
         ordered_img_data_8_0 : OUT std_logic ;
         ordered_img_data_9_31 : OUT std_logic ;
         ordered_img_data_9_30 : OUT std_logic ;
         ordered_img_data_9_29 : OUT std_logic ;
         ordered_img_data_9_28 : OUT std_logic ;
         ordered_img_data_9_27 : OUT std_logic ;
         ordered_img_data_9_26 : OUT std_logic ;
         ordered_img_data_9_25 : OUT std_logic ;
         ordered_img_data_9_24 : OUT std_logic ;
         ordered_img_data_9_23 : OUT std_logic ;
         ordered_img_data_9_22 : OUT std_logic ;
         ordered_img_data_9_21 : OUT std_logic ;
         ordered_img_data_9_20 : OUT std_logic ;
         ordered_img_data_9_19 : OUT std_logic ;
         ordered_img_data_9_18 : OUT std_logic ;
         ordered_img_data_9_17 : OUT std_logic ;
         ordered_img_data_9_16 : OUT std_logic ;
         ordered_img_data_9_15 : OUT std_logic ;
         ordered_img_data_9_14 : OUT std_logic ;
         ordered_img_data_9_13 : OUT std_logic ;
         ordered_img_data_9_12 : OUT std_logic ;
         ordered_img_data_9_11 : OUT std_logic ;
         ordered_img_data_9_10 : OUT std_logic ;
         ordered_img_data_9_9 : OUT std_logic ;
         ordered_img_data_9_8 : OUT std_logic ;
         ordered_img_data_9_7 : OUT std_logic ;
         ordered_img_data_9_6 : OUT std_logic ;
         ordered_img_data_9_5 : OUT std_logic ;
         ordered_img_data_9_4 : OUT std_logic ;
         ordered_img_data_9_3 : OUT std_logic ;
         ordered_img_data_9_2 : OUT std_logic ;
         ordered_img_data_9_1 : OUT std_logic ;
         ordered_img_data_9_0 : OUT std_logic ;
         ordered_img_data_10_31 : OUT std_logic ;
         ordered_img_data_10_30 : OUT std_logic ;
         ordered_img_data_10_29 : OUT std_logic ;
         ordered_img_data_10_28 : OUT std_logic ;
         ordered_img_data_10_27 : OUT std_logic ;
         ordered_img_data_10_26 : OUT std_logic ;
         ordered_img_data_10_25 : OUT std_logic ;
         ordered_img_data_10_24 : OUT std_logic ;
         ordered_img_data_10_23 : OUT std_logic ;
         ordered_img_data_10_22 : OUT std_logic ;
         ordered_img_data_10_21 : OUT std_logic ;
         ordered_img_data_10_20 : OUT std_logic ;
         ordered_img_data_10_19 : OUT std_logic ;
         ordered_img_data_10_18 : OUT std_logic ;
         ordered_img_data_10_17 : OUT std_logic ;
         ordered_img_data_10_16 : OUT std_logic ;
         ordered_img_data_10_15 : OUT std_logic ;
         ordered_img_data_10_14 : OUT std_logic ;
         ordered_img_data_10_13 : OUT std_logic ;
         ordered_img_data_10_12 : OUT std_logic ;
         ordered_img_data_10_11 : OUT std_logic ;
         ordered_img_data_10_10 : OUT std_logic ;
         ordered_img_data_10_9 : OUT std_logic ;
         ordered_img_data_10_8 : OUT std_logic ;
         ordered_img_data_10_7 : OUT std_logic ;
         ordered_img_data_10_6 : OUT std_logic ;
         ordered_img_data_10_5 : OUT std_logic ;
         ordered_img_data_10_4 : OUT std_logic ;
         ordered_img_data_10_3 : OUT std_logic ;
         ordered_img_data_10_2 : OUT std_logic ;
         ordered_img_data_10_1 : OUT std_logic ;
         ordered_img_data_10_0 : OUT std_logic ;
         ordered_img_data_11_31 : OUT std_logic ;
         ordered_img_data_11_30 : OUT std_logic ;
         ordered_img_data_11_29 : OUT std_logic ;
         ordered_img_data_11_28 : OUT std_logic ;
         ordered_img_data_11_27 : OUT std_logic ;
         ordered_img_data_11_26 : OUT std_logic ;
         ordered_img_data_11_25 : OUT std_logic ;
         ordered_img_data_11_24 : OUT std_logic ;
         ordered_img_data_11_23 : OUT std_logic ;
         ordered_img_data_11_22 : OUT std_logic ;
         ordered_img_data_11_21 : OUT std_logic ;
         ordered_img_data_11_20 : OUT std_logic ;
         ordered_img_data_11_19 : OUT std_logic ;
         ordered_img_data_11_18 : OUT std_logic ;
         ordered_img_data_11_17 : OUT std_logic ;
         ordered_img_data_11_16 : OUT std_logic ;
         ordered_img_data_11_15 : OUT std_logic ;
         ordered_img_data_11_14 : OUT std_logic ;
         ordered_img_data_11_13 : OUT std_logic ;
         ordered_img_data_11_12 : OUT std_logic ;
         ordered_img_data_11_11 : OUT std_logic ;
         ordered_img_data_11_10 : OUT std_logic ;
         ordered_img_data_11_9 : OUT std_logic ;
         ordered_img_data_11_8 : OUT std_logic ;
         ordered_img_data_11_7 : OUT std_logic ;
         ordered_img_data_11_6 : OUT std_logic ;
         ordered_img_data_11_5 : OUT std_logic ;
         ordered_img_data_11_4 : OUT std_logic ;
         ordered_img_data_11_3 : OUT std_logic ;
         ordered_img_data_11_2 : OUT std_logic ;
         ordered_img_data_11_1 : OUT std_logic ;
         ordered_img_data_11_0 : OUT std_logic ;
         ordered_img_data_12_31 : OUT std_logic ;
         ordered_img_data_12_30 : OUT std_logic ;
         ordered_img_data_12_29 : OUT std_logic ;
         ordered_img_data_12_28 : OUT std_logic ;
         ordered_img_data_12_27 : OUT std_logic ;
         ordered_img_data_12_26 : OUT std_logic ;
         ordered_img_data_12_25 : OUT std_logic ;
         ordered_img_data_12_24 : OUT std_logic ;
         ordered_img_data_12_23 : OUT std_logic ;
         ordered_img_data_12_22 : OUT std_logic ;
         ordered_img_data_12_21 : OUT std_logic ;
         ordered_img_data_12_20 : OUT std_logic ;
         ordered_img_data_12_19 : OUT std_logic ;
         ordered_img_data_12_18 : OUT std_logic ;
         ordered_img_data_12_17 : OUT std_logic ;
         ordered_img_data_12_16 : OUT std_logic ;
         ordered_img_data_12_15 : OUT std_logic ;
         ordered_img_data_12_14 : OUT std_logic ;
         ordered_img_data_12_13 : OUT std_logic ;
         ordered_img_data_12_12 : OUT std_logic ;
         ordered_img_data_12_11 : OUT std_logic ;
         ordered_img_data_12_10 : OUT std_logic ;
         ordered_img_data_12_9 : OUT std_logic ;
         ordered_img_data_12_8 : OUT std_logic ;
         ordered_img_data_12_7 : OUT std_logic ;
         ordered_img_data_12_6 : OUT std_logic ;
         ordered_img_data_12_5 : OUT std_logic ;
         ordered_img_data_12_4 : OUT std_logic ;
         ordered_img_data_12_3 : OUT std_logic ;
         ordered_img_data_12_2 : OUT std_logic ;
         ordered_img_data_12_1 : OUT std_logic ;
         ordered_img_data_12_0 : OUT std_logic ;
         ordered_img_data_13_31 : OUT std_logic ;
         ordered_img_data_13_30 : OUT std_logic ;
         ordered_img_data_13_29 : OUT std_logic ;
         ordered_img_data_13_28 : OUT std_logic ;
         ordered_img_data_13_27 : OUT std_logic ;
         ordered_img_data_13_26 : OUT std_logic ;
         ordered_img_data_13_25 : OUT std_logic ;
         ordered_img_data_13_24 : OUT std_logic ;
         ordered_img_data_13_23 : OUT std_logic ;
         ordered_img_data_13_22 : OUT std_logic ;
         ordered_img_data_13_21 : OUT std_logic ;
         ordered_img_data_13_20 : OUT std_logic ;
         ordered_img_data_13_19 : OUT std_logic ;
         ordered_img_data_13_18 : OUT std_logic ;
         ordered_img_data_13_17 : OUT std_logic ;
         ordered_img_data_13_16 : OUT std_logic ;
         ordered_img_data_13_15 : OUT std_logic ;
         ordered_img_data_13_14 : OUT std_logic ;
         ordered_img_data_13_13 : OUT std_logic ;
         ordered_img_data_13_12 : OUT std_logic ;
         ordered_img_data_13_11 : OUT std_logic ;
         ordered_img_data_13_10 : OUT std_logic ;
         ordered_img_data_13_9 : OUT std_logic ;
         ordered_img_data_13_8 : OUT std_logic ;
         ordered_img_data_13_7 : OUT std_logic ;
         ordered_img_data_13_6 : OUT std_logic ;
         ordered_img_data_13_5 : OUT std_logic ;
         ordered_img_data_13_4 : OUT std_logic ;
         ordered_img_data_13_3 : OUT std_logic ;
         ordered_img_data_13_2 : OUT std_logic ;
         ordered_img_data_13_1 : OUT std_logic ;
         ordered_img_data_13_0 : OUT std_logic ;
         ordered_img_data_14_31 : OUT std_logic ;
         ordered_img_data_14_30 : OUT std_logic ;
         ordered_img_data_14_29 : OUT std_logic ;
         ordered_img_data_14_28 : OUT std_logic ;
         ordered_img_data_14_27 : OUT std_logic ;
         ordered_img_data_14_26 : OUT std_logic ;
         ordered_img_data_14_25 : OUT std_logic ;
         ordered_img_data_14_24 : OUT std_logic ;
         ordered_img_data_14_23 : OUT std_logic ;
         ordered_img_data_14_22 : OUT std_logic ;
         ordered_img_data_14_21 : OUT std_logic ;
         ordered_img_data_14_20 : OUT std_logic ;
         ordered_img_data_14_19 : OUT std_logic ;
         ordered_img_data_14_18 : OUT std_logic ;
         ordered_img_data_14_17 : OUT std_logic ;
         ordered_img_data_14_16 : OUT std_logic ;
         ordered_img_data_14_15 : OUT std_logic ;
         ordered_img_data_14_14 : OUT std_logic ;
         ordered_img_data_14_13 : OUT std_logic ;
         ordered_img_data_14_12 : OUT std_logic ;
         ordered_img_data_14_11 : OUT std_logic ;
         ordered_img_data_14_10 : OUT std_logic ;
         ordered_img_data_14_9 : OUT std_logic ;
         ordered_img_data_14_8 : OUT std_logic ;
         ordered_img_data_14_7 : OUT std_logic ;
         ordered_img_data_14_6 : OUT std_logic ;
         ordered_img_data_14_5 : OUT std_logic ;
         ordered_img_data_14_4 : OUT std_logic ;
         ordered_img_data_14_3 : OUT std_logic ;
         ordered_img_data_14_2 : OUT std_logic ;
         ordered_img_data_14_1 : OUT std_logic ;
         ordered_img_data_14_0 : OUT std_logic ;
         ordered_img_data_15_31 : OUT std_logic ;
         ordered_img_data_15_30 : OUT std_logic ;
         ordered_img_data_15_29 : OUT std_logic ;
         ordered_img_data_15_28 : OUT std_logic ;
         ordered_img_data_15_27 : OUT std_logic ;
         ordered_img_data_15_26 : OUT std_logic ;
         ordered_img_data_15_25 : OUT std_logic ;
         ordered_img_data_15_24 : OUT std_logic ;
         ordered_img_data_15_23 : OUT std_logic ;
         ordered_img_data_15_22 : OUT std_logic ;
         ordered_img_data_15_21 : OUT std_logic ;
         ordered_img_data_15_20 : OUT std_logic ;
         ordered_img_data_15_19 : OUT std_logic ;
         ordered_img_data_15_18 : OUT std_logic ;
         ordered_img_data_15_17 : OUT std_logic ;
         ordered_img_data_15_16 : OUT std_logic ;
         ordered_img_data_15_15 : OUT std_logic ;
         ordered_img_data_15_14 : OUT std_logic ;
         ordered_img_data_15_13 : OUT std_logic ;
         ordered_img_data_15_12 : OUT std_logic ;
         ordered_img_data_15_11 : OUT std_logic ;
         ordered_img_data_15_10 : OUT std_logic ;
         ordered_img_data_15_9 : OUT std_logic ;
         ordered_img_data_15_8 : OUT std_logic ;
         ordered_img_data_15_7 : OUT std_logic ;
         ordered_img_data_15_6 : OUT std_logic ;
         ordered_img_data_15_5 : OUT std_logic ;
         ordered_img_data_15_4 : OUT std_logic ;
         ordered_img_data_15_3 : OUT std_logic ;
         ordered_img_data_15_2 : OUT std_logic ;
         ordered_img_data_15_1 : OUT std_logic ;
         ordered_img_data_15_0 : OUT std_logic ;
         ordered_img_data_16_31 : OUT std_logic ;
         ordered_img_data_16_30 : OUT std_logic ;
         ordered_img_data_16_29 : OUT std_logic ;
         ordered_img_data_16_28 : OUT std_logic ;
         ordered_img_data_16_27 : OUT std_logic ;
         ordered_img_data_16_26 : OUT std_logic ;
         ordered_img_data_16_25 : OUT std_logic ;
         ordered_img_data_16_24 : OUT std_logic ;
         ordered_img_data_16_23 : OUT std_logic ;
         ordered_img_data_16_22 : OUT std_logic ;
         ordered_img_data_16_21 : OUT std_logic ;
         ordered_img_data_16_20 : OUT std_logic ;
         ordered_img_data_16_19 : OUT std_logic ;
         ordered_img_data_16_18 : OUT std_logic ;
         ordered_img_data_16_17 : OUT std_logic ;
         ordered_img_data_16_16 : OUT std_logic ;
         ordered_img_data_16_15 : OUT std_logic ;
         ordered_img_data_16_14 : OUT std_logic ;
         ordered_img_data_16_13 : OUT std_logic ;
         ordered_img_data_16_12 : OUT std_logic ;
         ordered_img_data_16_11 : OUT std_logic ;
         ordered_img_data_16_10 : OUT std_logic ;
         ordered_img_data_16_9 : OUT std_logic ;
         ordered_img_data_16_8 : OUT std_logic ;
         ordered_img_data_16_7 : OUT std_logic ;
         ordered_img_data_16_6 : OUT std_logic ;
         ordered_img_data_16_5 : OUT std_logic ;
         ordered_img_data_16_4 : OUT std_logic ;
         ordered_img_data_16_3 : OUT std_logic ;
         ordered_img_data_16_2 : OUT std_logic ;
         ordered_img_data_16_1 : OUT std_logic ;
         ordered_img_data_16_0 : OUT std_logic ;
         ordered_img_data_17_31 : OUT std_logic ;
         ordered_img_data_17_30 : OUT std_logic ;
         ordered_img_data_17_29 : OUT std_logic ;
         ordered_img_data_17_28 : OUT std_logic ;
         ordered_img_data_17_27 : OUT std_logic ;
         ordered_img_data_17_26 : OUT std_logic ;
         ordered_img_data_17_25 : OUT std_logic ;
         ordered_img_data_17_24 : OUT std_logic ;
         ordered_img_data_17_23 : OUT std_logic ;
         ordered_img_data_17_22 : OUT std_logic ;
         ordered_img_data_17_21 : OUT std_logic ;
         ordered_img_data_17_20 : OUT std_logic ;
         ordered_img_data_17_19 : OUT std_logic ;
         ordered_img_data_17_18 : OUT std_logic ;
         ordered_img_data_17_17 : OUT std_logic ;
         ordered_img_data_17_16 : OUT std_logic ;
         ordered_img_data_17_15 : OUT std_logic ;
         ordered_img_data_17_14 : OUT std_logic ;
         ordered_img_data_17_13 : OUT std_logic ;
         ordered_img_data_17_12 : OUT std_logic ;
         ordered_img_data_17_11 : OUT std_logic ;
         ordered_img_data_17_10 : OUT std_logic ;
         ordered_img_data_17_9 : OUT std_logic ;
         ordered_img_data_17_8 : OUT std_logic ;
         ordered_img_data_17_7 : OUT std_logic ;
         ordered_img_data_17_6 : OUT std_logic ;
         ordered_img_data_17_5 : OUT std_logic ;
         ordered_img_data_17_4 : OUT std_logic ;
         ordered_img_data_17_3 : OUT std_logic ;
         ordered_img_data_17_2 : OUT std_logic ;
         ordered_img_data_17_1 : OUT std_logic ;
         ordered_img_data_17_0 : OUT std_logic ;
         ordered_img_data_18_31 : OUT std_logic ;
         ordered_img_data_18_30 : OUT std_logic ;
         ordered_img_data_18_29 : OUT std_logic ;
         ordered_img_data_18_28 : OUT std_logic ;
         ordered_img_data_18_27 : OUT std_logic ;
         ordered_img_data_18_26 : OUT std_logic ;
         ordered_img_data_18_25 : OUT std_logic ;
         ordered_img_data_18_24 : OUT std_logic ;
         ordered_img_data_18_23 : OUT std_logic ;
         ordered_img_data_18_22 : OUT std_logic ;
         ordered_img_data_18_21 : OUT std_logic ;
         ordered_img_data_18_20 : OUT std_logic ;
         ordered_img_data_18_19 : OUT std_logic ;
         ordered_img_data_18_18 : OUT std_logic ;
         ordered_img_data_18_17 : OUT std_logic ;
         ordered_img_data_18_16 : OUT std_logic ;
         ordered_img_data_18_15 : OUT std_logic ;
         ordered_img_data_18_14 : OUT std_logic ;
         ordered_img_data_18_13 : OUT std_logic ;
         ordered_img_data_18_12 : OUT std_logic ;
         ordered_img_data_18_11 : OUT std_logic ;
         ordered_img_data_18_10 : OUT std_logic ;
         ordered_img_data_18_9 : OUT std_logic ;
         ordered_img_data_18_8 : OUT std_logic ;
         ordered_img_data_18_7 : OUT std_logic ;
         ordered_img_data_18_6 : OUT std_logic ;
         ordered_img_data_18_5 : OUT std_logic ;
         ordered_img_data_18_4 : OUT std_logic ;
         ordered_img_data_18_3 : OUT std_logic ;
         ordered_img_data_18_2 : OUT std_logic ;
         ordered_img_data_18_1 : OUT std_logic ;
         ordered_img_data_18_0 : OUT std_logic ;
         ordered_img_data_19_31 : OUT std_logic ;
         ordered_img_data_19_30 : OUT std_logic ;
         ordered_img_data_19_29 : OUT std_logic ;
         ordered_img_data_19_28 : OUT std_logic ;
         ordered_img_data_19_27 : OUT std_logic ;
         ordered_img_data_19_26 : OUT std_logic ;
         ordered_img_data_19_25 : OUT std_logic ;
         ordered_img_data_19_24 : OUT std_logic ;
         ordered_img_data_19_23 : OUT std_logic ;
         ordered_img_data_19_22 : OUT std_logic ;
         ordered_img_data_19_21 : OUT std_logic ;
         ordered_img_data_19_20 : OUT std_logic ;
         ordered_img_data_19_19 : OUT std_logic ;
         ordered_img_data_19_18 : OUT std_logic ;
         ordered_img_data_19_17 : OUT std_logic ;
         ordered_img_data_19_16 : OUT std_logic ;
         ordered_img_data_19_15 : OUT std_logic ;
         ordered_img_data_19_14 : OUT std_logic ;
         ordered_img_data_19_13 : OUT std_logic ;
         ordered_img_data_19_12 : OUT std_logic ;
         ordered_img_data_19_11 : OUT std_logic ;
         ordered_img_data_19_10 : OUT std_logic ;
         ordered_img_data_19_9 : OUT std_logic ;
         ordered_img_data_19_8 : OUT std_logic ;
         ordered_img_data_19_7 : OUT std_logic ;
         ordered_img_data_19_6 : OUT std_logic ;
         ordered_img_data_19_5 : OUT std_logic ;
         ordered_img_data_19_4 : OUT std_logic ;
         ordered_img_data_19_3 : OUT std_logic ;
         ordered_img_data_19_2 : OUT std_logic ;
         ordered_img_data_19_1 : OUT std_logic ;
         ordered_img_data_19_0 : OUT std_logic ;
         ordered_img_data_20_31 : OUT std_logic ;
         ordered_img_data_20_30 : OUT std_logic ;
         ordered_img_data_20_29 : OUT std_logic ;
         ordered_img_data_20_28 : OUT std_logic ;
         ordered_img_data_20_27 : OUT std_logic ;
         ordered_img_data_20_26 : OUT std_logic ;
         ordered_img_data_20_25 : OUT std_logic ;
         ordered_img_data_20_24 : OUT std_logic ;
         ordered_img_data_20_23 : OUT std_logic ;
         ordered_img_data_20_22 : OUT std_logic ;
         ordered_img_data_20_21 : OUT std_logic ;
         ordered_img_data_20_20 : OUT std_logic ;
         ordered_img_data_20_19 : OUT std_logic ;
         ordered_img_data_20_18 : OUT std_logic ;
         ordered_img_data_20_17 : OUT std_logic ;
         ordered_img_data_20_16 : OUT std_logic ;
         ordered_img_data_20_15 : OUT std_logic ;
         ordered_img_data_20_14 : OUT std_logic ;
         ordered_img_data_20_13 : OUT std_logic ;
         ordered_img_data_20_12 : OUT std_logic ;
         ordered_img_data_20_11 : OUT std_logic ;
         ordered_img_data_20_10 : OUT std_logic ;
         ordered_img_data_20_9 : OUT std_logic ;
         ordered_img_data_20_8 : OUT std_logic ;
         ordered_img_data_20_7 : OUT std_logic ;
         ordered_img_data_20_6 : OUT std_logic ;
         ordered_img_data_20_5 : OUT std_logic ;
         ordered_img_data_20_4 : OUT std_logic ;
         ordered_img_data_20_3 : OUT std_logic ;
         ordered_img_data_20_2 : OUT std_logic ;
         ordered_img_data_20_1 : OUT std_logic ;
         ordered_img_data_20_0 : OUT std_logic ;
         ordered_img_data_21_31 : OUT std_logic ;
         ordered_img_data_21_30 : OUT std_logic ;
         ordered_img_data_21_29 : OUT std_logic ;
         ordered_img_data_21_28 : OUT std_logic ;
         ordered_img_data_21_27 : OUT std_logic ;
         ordered_img_data_21_26 : OUT std_logic ;
         ordered_img_data_21_25 : OUT std_logic ;
         ordered_img_data_21_24 : OUT std_logic ;
         ordered_img_data_21_23 : OUT std_logic ;
         ordered_img_data_21_22 : OUT std_logic ;
         ordered_img_data_21_21 : OUT std_logic ;
         ordered_img_data_21_20 : OUT std_logic ;
         ordered_img_data_21_19 : OUT std_logic ;
         ordered_img_data_21_18 : OUT std_logic ;
         ordered_img_data_21_17 : OUT std_logic ;
         ordered_img_data_21_16 : OUT std_logic ;
         ordered_img_data_21_15 : OUT std_logic ;
         ordered_img_data_21_14 : OUT std_logic ;
         ordered_img_data_21_13 : OUT std_logic ;
         ordered_img_data_21_12 : OUT std_logic ;
         ordered_img_data_21_11 : OUT std_logic ;
         ordered_img_data_21_10 : OUT std_logic ;
         ordered_img_data_21_9 : OUT std_logic ;
         ordered_img_data_21_8 : OUT std_logic ;
         ordered_img_data_21_7 : OUT std_logic ;
         ordered_img_data_21_6 : OUT std_logic ;
         ordered_img_data_21_5 : OUT std_logic ;
         ordered_img_data_21_4 : OUT std_logic ;
         ordered_img_data_21_3 : OUT std_logic ;
         ordered_img_data_21_2 : OUT std_logic ;
         ordered_img_data_21_1 : OUT std_logic ;
         ordered_img_data_21_0 : OUT std_logic ;
         ordered_img_data_22_31 : OUT std_logic ;
         ordered_img_data_22_30 : OUT std_logic ;
         ordered_img_data_22_29 : OUT std_logic ;
         ordered_img_data_22_28 : OUT std_logic ;
         ordered_img_data_22_27 : OUT std_logic ;
         ordered_img_data_22_26 : OUT std_logic ;
         ordered_img_data_22_25 : OUT std_logic ;
         ordered_img_data_22_24 : OUT std_logic ;
         ordered_img_data_22_23 : OUT std_logic ;
         ordered_img_data_22_22 : OUT std_logic ;
         ordered_img_data_22_21 : OUT std_logic ;
         ordered_img_data_22_20 : OUT std_logic ;
         ordered_img_data_22_19 : OUT std_logic ;
         ordered_img_data_22_18 : OUT std_logic ;
         ordered_img_data_22_17 : OUT std_logic ;
         ordered_img_data_22_16 : OUT std_logic ;
         ordered_img_data_22_15 : OUT std_logic ;
         ordered_img_data_22_14 : OUT std_logic ;
         ordered_img_data_22_13 : OUT std_logic ;
         ordered_img_data_22_12 : OUT std_logic ;
         ordered_img_data_22_11 : OUT std_logic ;
         ordered_img_data_22_10 : OUT std_logic ;
         ordered_img_data_22_9 : OUT std_logic ;
         ordered_img_data_22_8 : OUT std_logic ;
         ordered_img_data_22_7 : OUT std_logic ;
         ordered_img_data_22_6 : OUT std_logic ;
         ordered_img_data_22_5 : OUT std_logic ;
         ordered_img_data_22_4 : OUT std_logic ;
         ordered_img_data_22_3 : OUT std_logic ;
         ordered_img_data_22_2 : OUT std_logic ;
         ordered_img_data_22_1 : OUT std_logic ;
         ordered_img_data_22_0 : OUT std_logic ;
         ordered_img_data_23_31 : OUT std_logic ;
         ordered_img_data_23_30 : OUT std_logic ;
         ordered_img_data_23_29 : OUT std_logic ;
         ordered_img_data_23_28 : OUT std_logic ;
         ordered_img_data_23_27 : OUT std_logic ;
         ordered_img_data_23_26 : OUT std_logic ;
         ordered_img_data_23_25 : OUT std_logic ;
         ordered_img_data_23_24 : OUT std_logic ;
         ordered_img_data_23_23 : OUT std_logic ;
         ordered_img_data_23_22 : OUT std_logic ;
         ordered_img_data_23_21 : OUT std_logic ;
         ordered_img_data_23_20 : OUT std_logic ;
         ordered_img_data_23_19 : OUT std_logic ;
         ordered_img_data_23_18 : OUT std_logic ;
         ordered_img_data_23_17 : OUT std_logic ;
         ordered_img_data_23_16 : OUT std_logic ;
         ordered_img_data_23_15 : OUT std_logic ;
         ordered_img_data_23_14 : OUT std_logic ;
         ordered_img_data_23_13 : OUT std_logic ;
         ordered_img_data_23_12 : OUT std_logic ;
         ordered_img_data_23_11 : OUT std_logic ;
         ordered_img_data_23_10 : OUT std_logic ;
         ordered_img_data_23_9 : OUT std_logic ;
         ordered_img_data_23_8 : OUT std_logic ;
         ordered_img_data_23_7 : OUT std_logic ;
         ordered_img_data_23_6 : OUT std_logic ;
         ordered_img_data_23_5 : OUT std_logic ;
         ordered_img_data_23_4 : OUT std_logic ;
         ordered_img_data_23_3 : OUT std_logic ;
         ordered_img_data_23_2 : OUT std_logic ;
         ordered_img_data_23_1 : OUT std_logic ;
         ordered_img_data_23_0 : OUT std_logic ;
         ordered_img_data_24_31 : OUT std_logic ;
         ordered_img_data_24_30 : OUT std_logic ;
         ordered_img_data_24_29 : OUT std_logic ;
         ordered_img_data_24_28 : OUT std_logic ;
         ordered_img_data_24_27 : OUT std_logic ;
         ordered_img_data_24_26 : OUT std_logic ;
         ordered_img_data_24_25 : OUT std_logic ;
         ordered_img_data_24_24 : OUT std_logic ;
         ordered_img_data_24_23 : OUT std_logic ;
         ordered_img_data_24_22 : OUT std_logic ;
         ordered_img_data_24_21 : OUT std_logic ;
         ordered_img_data_24_20 : OUT std_logic ;
         ordered_img_data_24_19 : OUT std_logic ;
         ordered_img_data_24_18 : OUT std_logic ;
         ordered_img_data_24_17 : OUT std_logic ;
         ordered_img_data_24_16 : OUT std_logic ;
         ordered_img_data_24_15 : OUT std_logic ;
         ordered_img_data_24_14 : OUT std_logic ;
         ordered_img_data_24_13 : OUT std_logic ;
         ordered_img_data_24_12 : OUT std_logic ;
         ordered_img_data_24_11 : OUT std_logic ;
         ordered_img_data_24_10 : OUT std_logic ;
         ordered_img_data_24_9 : OUT std_logic ;
         ordered_img_data_24_8 : OUT std_logic ;
         ordered_img_data_24_7 : OUT std_logic ;
         ordered_img_data_24_6 : OUT std_logic ;
         ordered_img_data_24_5 : OUT std_logic ;
         ordered_img_data_24_4 : OUT std_logic ;
         ordered_img_data_24_3 : OUT std_logic ;
         ordered_img_data_24_2 : OUT std_logic ;
         ordered_img_data_24_1 : OUT std_logic ;
         ordered_img_data_24_0 : OUT std_logic ;
         ordered_filter_data_0_31 : OUT std_logic ;
         ordered_filter_data_0_30 : OUT std_logic ;
         ordered_filter_data_0_29 : OUT std_logic ;
         ordered_filter_data_0_28 : OUT std_logic ;
         ordered_filter_data_0_27 : OUT std_logic ;
         ordered_filter_data_0_26 : OUT std_logic ;
         ordered_filter_data_0_25 : OUT std_logic ;
         ordered_filter_data_0_24 : OUT std_logic ;
         ordered_filter_data_0_23 : OUT std_logic ;
         ordered_filter_data_0_22 : OUT std_logic ;
         ordered_filter_data_0_21 : OUT std_logic ;
         ordered_filter_data_0_20 : OUT std_logic ;
         ordered_filter_data_0_19 : OUT std_logic ;
         ordered_filter_data_0_18 : OUT std_logic ;
         ordered_filter_data_0_17 : OUT std_logic ;
         ordered_filter_data_0_16 : OUT std_logic ;
         ordered_filter_data_0_15 : OUT std_logic ;
         ordered_filter_data_0_14 : OUT std_logic ;
         ordered_filter_data_0_13 : OUT std_logic ;
         ordered_filter_data_0_12 : OUT std_logic ;
         ordered_filter_data_0_11 : OUT std_logic ;
         ordered_filter_data_0_10 : OUT std_logic ;
         ordered_filter_data_0_9 : OUT std_logic ;
         ordered_filter_data_0_8 : OUT std_logic ;
         ordered_filter_data_0_7 : OUT std_logic ;
         ordered_filter_data_0_6 : OUT std_logic ;
         ordered_filter_data_0_5 : OUT std_logic ;
         ordered_filter_data_0_4 : OUT std_logic ;
         ordered_filter_data_0_3 : OUT std_logic ;
         ordered_filter_data_0_2 : OUT std_logic ;
         ordered_filter_data_0_1 : OUT std_logic ;
         ordered_filter_data_0_0 : OUT std_logic ;
         ordered_filter_data_1_31 : OUT std_logic ;
         ordered_filter_data_1_30 : OUT std_logic ;
         ordered_filter_data_1_29 : OUT std_logic ;
         ordered_filter_data_1_28 : OUT std_logic ;
         ordered_filter_data_1_27 : OUT std_logic ;
         ordered_filter_data_1_26 : OUT std_logic ;
         ordered_filter_data_1_25 : OUT std_logic ;
         ordered_filter_data_1_24 : OUT std_logic ;
         ordered_filter_data_1_23 : OUT std_logic ;
         ordered_filter_data_1_22 : OUT std_logic ;
         ordered_filter_data_1_21 : OUT std_logic ;
         ordered_filter_data_1_20 : OUT std_logic ;
         ordered_filter_data_1_19 : OUT std_logic ;
         ordered_filter_data_1_18 : OUT std_logic ;
         ordered_filter_data_1_17 : OUT std_logic ;
         ordered_filter_data_1_16 : OUT std_logic ;
         ordered_filter_data_1_15 : OUT std_logic ;
         ordered_filter_data_1_14 : OUT std_logic ;
         ordered_filter_data_1_13 : OUT std_logic ;
         ordered_filter_data_1_12 : OUT std_logic ;
         ordered_filter_data_1_11 : OUT std_logic ;
         ordered_filter_data_1_10 : OUT std_logic ;
         ordered_filter_data_1_9 : OUT std_logic ;
         ordered_filter_data_1_8 : OUT std_logic ;
         ordered_filter_data_1_7 : OUT std_logic ;
         ordered_filter_data_1_6 : OUT std_logic ;
         ordered_filter_data_1_5 : OUT std_logic ;
         ordered_filter_data_1_4 : OUT std_logic ;
         ordered_filter_data_1_3 : OUT std_logic ;
         ordered_filter_data_1_2 : OUT std_logic ;
         ordered_filter_data_1_1 : OUT std_logic ;
         ordered_filter_data_1_0 : OUT std_logic ;
         ordered_filter_data_2_31 : OUT std_logic ;
         ordered_filter_data_2_30 : OUT std_logic ;
         ordered_filter_data_2_29 : OUT std_logic ;
         ordered_filter_data_2_28 : OUT std_logic ;
         ordered_filter_data_2_27 : OUT std_logic ;
         ordered_filter_data_2_26 : OUT std_logic ;
         ordered_filter_data_2_25 : OUT std_logic ;
         ordered_filter_data_2_24 : OUT std_logic ;
         ordered_filter_data_2_23 : OUT std_logic ;
         ordered_filter_data_2_22 : OUT std_logic ;
         ordered_filter_data_2_21 : OUT std_logic ;
         ordered_filter_data_2_20 : OUT std_logic ;
         ordered_filter_data_2_19 : OUT std_logic ;
         ordered_filter_data_2_18 : OUT std_logic ;
         ordered_filter_data_2_17 : OUT std_logic ;
         ordered_filter_data_2_16 : OUT std_logic ;
         ordered_filter_data_2_15 : OUT std_logic ;
         ordered_filter_data_2_14 : OUT std_logic ;
         ordered_filter_data_2_13 : OUT std_logic ;
         ordered_filter_data_2_12 : OUT std_logic ;
         ordered_filter_data_2_11 : OUT std_logic ;
         ordered_filter_data_2_10 : OUT std_logic ;
         ordered_filter_data_2_9 : OUT std_logic ;
         ordered_filter_data_2_8 : OUT std_logic ;
         ordered_filter_data_2_7 : OUT std_logic ;
         ordered_filter_data_2_6 : OUT std_logic ;
         ordered_filter_data_2_5 : OUT std_logic ;
         ordered_filter_data_2_4 : OUT std_logic ;
         ordered_filter_data_2_3 : OUT std_logic ;
         ordered_filter_data_2_2 : OUT std_logic ;
         ordered_filter_data_2_1 : OUT std_logic ;
         ordered_filter_data_2_0 : OUT std_logic ;
         ordered_filter_data_3_31 : OUT std_logic ;
         ordered_filter_data_3_30 : OUT std_logic ;
         ordered_filter_data_3_29 : OUT std_logic ;
         ordered_filter_data_3_28 : OUT std_logic ;
         ordered_filter_data_3_27 : OUT std_logic ;
         ordered_filter_data_3_26 : OUT std_logic ;
         ordered_filter_data_3_25 : OUT std_logic ;
         ordered_filter_data_3_24 : OUT std_logic ;
         ordered_filter_data_3_23 : OUT std_logic ;
         ordered_filter_data_3_22 : OUT std_logic ;
         ordered_filter_data_3_21 : OUT std_logic ;
         ordered_filter_data_3_20 : OUT std_logic ;
         ordered_filter_data_3_19 : OUT std_logic ;
         ordered_filter_data_3_18 : OUT std_logic ;
         ordered_filter_data_3_17 : OUT std_logic ;
         ordered_filter_data_3_16 : OUT std_logic ;
         ordered_filter_data_3_15 : OUT std_logic ;
         ordered_filter_data_3_14 : OUT std_logic ;
         ordered_filter_data_3_13 : OUT std_logic ;
         ordered_filter_data_3_12 : OUT std_logic ;
         ordered_filter_data_3_11 : OUT std_logic ;
         ordered_filter_data_3_10 : OUT std_logic ;
         ordered_filter_data_3_9 : OUT std_logic ;
         ordered_filter_data_3_8 : OUT std_logic ;
         ordered_filter_data_3_7 : OUT std_logic ;
         ordered_filter_data_3_6 : OUT std_logic ;
         ordered_filter_data_3_5 : OUT std_logic ;
         ordered_filter_data_3_4 : OUT std_logic ;
         ordered_filter_data_3_3 : OUT std_logic ;
         ordered_filter_data_3_2 : OUT std_logic ;
         ordered_filter_data_3_1 : OUT std_logic ;
         ordered_filter_data_3_0 : OUT std_logic ;
         ordered_filter_data_4_31 : OUT std_logic ;
         ordered_filter_data_4_30 : OUT std_logic ;
         ordered_filter_data_4_29 : OUT std_logic ;
         ordered_filter_data_4_28 : OUT std_logic ;
         ordered_filter_data_4_27 : OUT std_logic ;
         ordered_filter_data_4_26 : OUT std_logic ;
         ordered_filter_data_4_25 : OUT std_logic ;
         ordered_filter_data_4_24 : OUT std_logic ;
         ordered_filter_data_4_23 : OUT std_logic ;
         ordered_filter_data_4_22 : OUT std_logic ;
         ordered_filter_data_4_21 : OUT std_logic ;
         ordered_filter_data_4_20 : OUT std_logic ;
         ordered_filter_data_4_19 : OUT std_logic ;
         ordered_filter_data_4_18 : OUT std_logic ;
         ordered_filter_data_4_17 : OUT std_logic ;
         ordered_filter_data_4_16 : OUT std_logic ;
         ordered_filter_data_4_15 : OUT std_logic ;
         ordered_filter_data_4_14 : OUT std_logic ;
         ordered_filter_data_4_13 : OUT std_logic ;
         ordered_filter_data_4_12 : OUT std_logic ;
         ordered_filter_data_4_11 : OUT std_logic ;
         ordered_filter_data_4_10 : OUT std_logic ;
         ordered_filter_data_4_9 : OUT std_logic ;
         ordered_filter_data_4_8 : OUT std_logic ;
         ordered_filter_data_4_7 : OUT std_logic ;
         ordered_filter_data_4_6 : OUT std_logic ;
         ordered_filter_data_4_5 : OUT std_logic ;
         ordered_filter_data_4_4 : OUT std_logic ;
         ordered_filter_data_4_3 : OUT std_logic ;
         ordered_filter_data_4_2 : OUT std_logic ;
         ordered_filter_data_4_1 : OUT std_logic ;
         ordered_filter_data_4_0 : OUT std_logic ;
         ordered_filter_data_5_31 : OUT std_logic ;
         ordered_filter_data_5_30 : OUT std_logic ;
         ordered_filter_data_5_29 : OUT std_logic ;
         ordered_filter_data_5_28 : OUT std_logic ;
         ordered_filter_data_5_27 : OUT std_logic ;
         ordered_filter_data_5_26 : OUT std_logic ;
         ordered_filter_data_5_25 : OUT std_logic ;
         ordered_filter_data_5_24 : OUT std_logic ;
         ordered_filter_data_5_23 : OUT std_logic ;
         ordered_filter_data_5_22 : OUT std_logic ;
         ordered_filter_data_5_21 : OUT std_logic ;
         ordered_filter_data_5_20 : OUT std_logic ;
         ordered_filter_data_5_19 : OUT std_logic ;
         ordered_filter_data_5_18 : OUT std_logic ;
         ordered_filter_data_5_17 : OUT std_logic ;
         ordered_filter_data_5_16 : OUT std_logic ;
         ordered_filter_data_5_15 : OUT std_logic ;
         ordered_filter_data_5_14 : OUT std_logic ;
         ordered_filter_data_5_13 : OUT std_logic ;
         ordered_filter_data_5_12 : OUT std_logic ;
         ordered_filter_data_5_11 : OUT std_logic ;
         ordered_filter_data_5_10 : OUT std_logic ;
         ordered_filter_data_5_9 : OUT std_logic ;
         ordered_filter_data_5_8 : OUT std_logic ;
         ordered_filter_data_5_7 : OUT std_logic ;
         ordered_filter_data_5_6 : OUT std_logic ;
         ordered_filter_data_5_5 : OUT std_logic ;
         ordered_filter_data_5_4 : OUT std_logic ;
         ordered_filter_data_5_3 : OUT std_logic ;
         ordered_filter_data_5_2 : OUT std_logic ;
         ordered_filter_data_5_1 : OUT std_logic ;
         ordered_filter_data_5_0 : OUT std_logic ;
         ordered_filter_data_6_31 : OUT std_logic ;
         ordered_filter_data_6_30 : OUT std_logic ;
         ordered_filter_data_6_29 : OUT std_logic ;
         ordered_filter_data_6_28 : OUT std_logic ;
         ordered_filter_data_6_27 : OUT std_logic ;
         ordered_filter_data_6_26 : OUT std_logic ;
         ordered_filter_data_6_25 : OUT std_logic ;
         ordered_filter_data_6_24 : OUT std_logic ;
         ordered_filter_data_6_23 : OUT std_logic ;
         ordered_filter_data_6_22 : OUT std_logic ;
         ordered_filter_data_6_21 : OUT std_logic ;
         ordered_filter_data_6_20 : OUT std_logic ;
         ordered_filter_data_6_19 : OUT std_logic ;
         ordered_filter_data_6_18 : OUT std_logic ;
         ordered_filter_data_6_17 : OUT std_logic ;
         ordered_filter_data_6_16 : OUT std_logic ;
         ordered_filter_data_6_15 : OUT std_logic ;
         ordered_filter_data_6_14 : OUT std_logic ;
         ordered_filter_data_6_13 : OUT std_logic ;
         ordered_filter_data_6_12 : OUT std_logic ;
         ordered_filter_data_6_11 : OUT std_logic ;
         ordered_filter_data_6_10 : OUT std_logic ;
         ordered_filter_data_6_9 : OUT std_logic ;
         ordered_filter_data_6_8 : OUT std_logic ;
         ordered_filter_data_6_7 : OUT std_logic ;
         ordered_filter_data_6_6 : OUT std_logic ;
         ordered_filter_data_6_5 : OUT std_logic ;
         ordered_filter_data_6_4 : OUT std_logic ;
         ordered_filter_data_6_3 : OUT std_logic ;
         ordered_filter_data_6_2 : OUT std_logic ;
         ordered_filter_data_6_1 : OUT std_logic ;
         ordered_filter_data_6_0 : OUT std_logic ;
         ordered_filter_data_7_31 : OUT std_logic ;
         ordered_filter_data_7_30 : OUT std_logic ;
         ordered_filter_data_7_29 : OUT std_logic ;
         ordered_filter_data_7_28 : OUT std_logic ;
         ordered_filter_data_7_27 : OUT std_logic ;
         ordered_filter_data_7_26 : OUT std_logic ;
         ordered_filter_data_7_25 : OUT std_logic ;
         ordered_filter_data_7_24 : OUT std_logic ;
         ordered_filter_data_7_23 : OUT std_logic ;
         ordered_filter_data_7_22 : OUT std_logic ;
         ordered_filter_data_7_21 : OUT std_logic ;
         ordered_filter_data_7_20 : OUT std_logic ;
         ordered_filter_data_7_19 : OUT std_logic ;
         ordered_filter_data_7_18 : OUT std_logic ;
         ordered_filter_data_7_17 : OUT std_logic ;
         ordered_filter_data_7_16 : OUT std_logic ;
         ordered_filter_data_7_15 : OUT std_logic ;
         ordered_filter_data_7_14 : OUT std_logic ;
         ordered_filter_data_7_13 : OUT std_logic ;
         ordered_filter_data_7_12 : OUT std_logic ;
         ordered_filter_data_7_11 : OUT std_logic ;
         ordered_filter_data_7_10 : OUT std_logic ;
         ordered_filter_data_7_9 : OUT std_logic ;
         ordered_filter_data_7_8 : OUT std_logic ;
         ordered_filter_data_7_7 : OUT std_logic ;
         ordered_filter_data_7_6 : OUT std_logic ;
         ordered_filter_data_7_5 : OUT std_logic ;
         ordered_filter_data_7_4 : OUT std_logic ;
         ordered_filter_data_7_3 : OUT std_logic ;
         ordered_filter_data_7_2 : OUT std_logic ;
         ordered_filter_data_7_1 : OUT std_logic ;
         ordered_filter_data_7_0 : OUT std_logic ;
         ordered_filter_data_8_31 : OUT std_logic ;
         ordered_filter_data_8_30 : OUT std_logic ;
         ordered_filter_data_8_29 : OUT std_logic ;
         ordered_filter_data_8_28 : OUT std_logic ;
         ordered_filter_data_8_27 : OUT std_logic ;
         ordered_filter_data_8_26 : OUT std_logic ;
         ordered_filter_data_8_25 : OUT std_logic ;
         ordered_filter_data_8_24 : OUT std_logic ;
         ordered_filter_data_8_23 : OUT std_logic ;
         ordered_filter_data_8_22 : OUT std_logic ;
         ordered_filter_data_8_21 : OUT std_logic ;
         ordered_filter_data_8_20 : OUT std_logic ;
         ordered_filter_data_8_19 : OUT std_logic ;
         ordered_filter_data_8_18 : OUT std_logic ;
         ordered_filter_data_8_17 : OUT std_logic ;
         ordered_filter_data_8_16 : OUT std_logic ;
         ordered_filter_data_8_15 : OUT std_logic ;
         ordered_filter_data_8_14 : OUT std_logic ;
         ordered_filter_data_8_13 : OUT std_logic ;
         ordered_filter_data_8_12 : OUT std_logic ;
         ordered_filter_data_8_11 : OUT std_logic ;
         ordered_filter_data_8_10 : OUT std_logic ;
         ordered_filter_data_8_9 : OUT std_logic ;
         ordered_filter_data_8_8 : OUT std_logic ;
         ordered_filter_data_8_7 : OUT std_logic ;
         ordered_filter_data_8_6 : OUT std_logic ;
         ordered_filter_data_8_5 : OUT std_logic ;
         ordered_filter_data_8_4 : OUT std_logic ;
         ordered_filter_data_8_3 : OUT std_logic ;
         ordered_filter_data_8_2 : OUT std_logic ;
         ordered_filter_data_8_1 : OUT std_logic ;
         ordered_filter_data_8_0 : OUT std_logic ;
         ordered_filter_data_9_31 : OUT std_logic ;
         ordered_filter_data_9_30 : OUT std_logic ;
         ordered_filter_data_9_29 : OUT std_logic ;
         ordered_filter_data_9_28 : OUT std_logic ;
         ordered_filter_data_9_27 : OUT std_logic ;
         ordered_filter_data_9_26 : OUT std_logic ;
         ordered_filter_data_9_25 : OUT std_logic ;
         ordered_filter_data_9_24 : OUT std_logic ;
         ordered_filter_data_9_23 : OUT std_logic ;
         ordered_filter_data_9_22 : OUT std_logic ;
         ordered_filter_data_9_21 : OUT std_logic ;
         ordered_filter_data_9_20 : OUT std_logic ;
         ordered_filter_data_9_19 : OUT std_logic ;
         ordered_filter_data_9_18 : OUT std_logic ;
         ordered_filter_data_9_17 : OUT std_logic ;
         ordered_filter_data_9_16 : OUT std_logic ;
         ordered_filter_data_9_15 : OUT std_logic ;
         ordered_filter_data_9_14 : OUT std_logic ;
         ordered_filter_data_9_13 : OUT std_logic ;
         ordered_filter_data_9_12 : OUT std_logic ;
         ordered_filter_data_9_11 : OUT std_logic ;
         ordered_filter_data_9_10 : OUT std_logic ;
         ordered_filter_data_9_9 : OUT std_logic ;
         ordered_filter_data_9_8 : OUT std_logic ;
         ordered_filter_data_9_7 : OUT std_logic ;
         ordered_filter_data_9_6 : OUT std_logic ;
         ordered_filter_data_9_5 : OUT std_logic ;
         ordered_filter_data_9_4 : OUT std_logic ;
         ordered_filter_data_9_3 : OUT std_logic ;
         ordered_filter_data_9_2 : OUT std_logic ;
         ordered_filter_data_9_1 : OUT std_logic ;
         ordered_filter_data_9_0 : OUT std_logic ;
         ordered_filter_data_10_31 : OUT std_logic ;
         ordered_filter_data_10_30 : OUT std_logic ;
         ordered_filter_data_10_29 : OUT std_logic ;
         ordered_filter_data_10_28 : OUT std_logic ;
         ordered_filter_data_10_27 : OUT std_logic ;
         ordered_filter_data_10_26 : OUT std_logic ;
         ordered_filter_data_10_25 : OUT std_logic ;
         ordered_filter_data_10_24 : OUT std_logic ;
         ordered_filter_data_10_23 : OUT std_logic ;
         ordered_filter_data_10_22 : OUT std_logic ;
         ordered_filter_data_10_21 : OUT std_logic ;
         ordered_filter_data_10_20 : OUT std_logic ;
         ordered_filter_data_10_19 : OUT std_logic ;
         ordered_filter_data_10_18 : OUT std_logic ;
         ordered_filter_data_10_17 : OUT std_logic ;
         ordered_filter_data_10_16 : OUT std_logic ;
         ordered_filter_data_10_15 : OUT std_logic ;
         ordered_filter_data_10_14 : OUT std_logic ;
         ordered_filter_data_10_13 : OUT std_logic ;
         ordered_filter_data_10_12 : OUT std_logic ;
         ordered_filter_data_10_11 : OUT std_logic ;
         ordered_filter_data_10_10 : OUT std_logic ;
         ordered_filter_data_10_9 : OUT std_logic ;
         ordered_filter_data_10_8 : OUT std_logic ;
         ordered_filter_data_10_7 : OUT std_logic ;
         ordered_filter_data_10_6 : OUT std_logic ;
         ordered_filter_data_10_5 : OUT std_logic ;
         ordered_filter_data_10_4 : OUT std_logic ;
         ordered_filter_data_10_3 : OUT std_logic ;
         ordered_filter_data_10_2 : OUT std_logic ;
         ordered_filter_data_10_1 : OUT std_logic ;
         ordered_filter_data_10_0 : OUT std_logic ;
         ordered_filter_data_11_31 : OUT std_logic ;
         ordered_filter_data_11_30 : OUT std_logic ;
         ordered_filter_data_11_29 : OUT std_logic ;
         ordered_filter_data_11_28 : OUT std_logic ;
         ordered_filter_data_11_27 : OUT std_logic ;
         ordered_filter_data_11_26 : OUT std_logic ;
         ordered_filter_data_11_25 : OUT std_logic ;
         ordered_filter_data_11_24 : OUT std_logic ;
         ordered_filter_data_11_23 : OUT std_logic ;
         ordered_filter_data_11_22 : OUT std_logic ;
         ordered_filter_data_11_21 : OUT std_logic ;
         ordered_filter_data_11_20 : OUT std_logic ;
         ordered_filter_data_11_19 : OUT std_logic ;
         ordered_filter_data_11_18 : OUT std_logic ;
         ordered_filter_data_11_17 : OUT std_logic ;
         ordered_filter_data_11_16 : OUT std_logic ;
         ordered_filter_data_11_15 : OUT std_logic ;
         ordered_filter_data_11_14 : OUT std_logic ;
         ordered_filter_data_11_13 : OUT std_logic ;
         ordered_filter_data_11_12 : OUT std_logic ;
         ordered_filter_data_11_11 : OUT std_logic ;
         ordered_filter_data_11_10 : OUT std_logic ;
         ordered_filter_data_11_9 : OUT std_logic ;
         ordered_filter_data_11_8 : OUT std_logic ;
         ordered_filter_data_11_7 : OUT std_logic ;
         ordered_filter_data_11_6 : OUT std_logic ;
         ordered_filter_data_11_5 : OUT std_logic ;
         ordered_filter_data_11_4 : OUT std_logic ;
         ordered_filter_data_11_3 : OUT std_logic ;
         ordered_filter_data_11_2 : OUT std_logic ;
         ordered_filter_data_11_1 : OUT std_logic ;
         ordered_filter_data_11_0 : OUT std_logic ;
         ordered_filter_data_12_31 : OUT std_logic ;
         ordered_filter_data_12_30 : OUT std_logic ;
         ordered_filter_data_12_29 : OUT std_logic ;
         ordered_filter_data_12_28 : OUT std_logic ;
         ordered_filter_data_12_27 : OUT std_logic ;
         ordered_filter_data_12_26 : OUT std_logic ;
         ordered_filter_data_12_25 : OUT std_logic ;
         ordered_filter_data_12_24 : OUT std_logic ;
         ordered_filter_data_12_23 : OUT std_logic ;
         ordered_filter_data_12_22 : OUT std_logic ;
         ordered_filter_data_12_21 : OUT std_logic ;
         ordered_filter_data_12_20 : OUT std_logic ;
         ordered_filter_data_12_19 : OUT std_logic ;
         ordered_filter_data_12_18 : OUT std_logic ;
         ordered_filter_data_12_17 : OUT std_logic ;
         ordered_filter_data_12_16 : OUT std_logic ;
         ordered_filter_data_12_15 : OUT std_logic ;
         ordered_filter_data_12_14 : OUT std_logic ;
         ordered_filter_data_12_13 : OUT std_logic ;
         ordered_filter_data_12_12 : OUT std_logic ;
         ordered_filter_data_12_11 : OUT std_logic ;
         ordered_filter_data_12_10 : OUT std_logic ;
         ordered_filter_data_12_9 : OUT std_logic ;
         ordered_filter_data_12_8 : OUT std_logic ;
         ordered_filter_data_12_7 : OUT std_logic ;
         ordered_filter_data_12_6 : OUT std_logic ;
         ordered_filter_data_12_5 : OUT std_logic ;
         ordered_filter_data_12_4 : OUT std_logic ;
         ordered_filter_data_12_3 : OUT std_logic ;
         ordered_filter_data_12_2 : OUT std_logic ;
         ordered_filter_data_12_1 : OUT std_logic ;
         ordered_filter_data_12_0 : OUT std_logic ;
         ordered_filter_data_13_31 : OUT std_logic ;
         ordered_filter_data_13_30 : OUT std_logic ;
         ordered_filter_data_13_29 : OUT std_logic ;
         ordered_filter_data_13_28 : OUT std_logic ;
         ordered_filter_data_13_27 : OUT std_logic ;
         ordered_filter_data_13_26 : OUT std_logic ;
         ordered_filter_data_13_25 : OUT std_logic ;
         ordered_filter_data_13_24 : OUT std_logic ;
         ordered_filter_data_13_23 : OUT std_logic ;
         ordered_filter_data_13_22 : OUT std_logic ;
         ordered_filter_data_13_21 : OUT std_logic ;
         ordered_filter_data_13_20 : OUT std_logic ;
         ordered_filter_data_13_19 : OUT std_logic ;
         ordered_filter_data_13_18 : OUT std_logic ;
         ordered_filter_data_13_17 : OUT std_logic ;
         ordered_filter_data_13_16 : OUT std_logic ;
         ordered_filter_data_13_15 : OUT std_logic ;
         ordered_filter_data_13_14 : OUT std_logic ;
         ordered_filter_data_13_13 : OUT std_logic ;
         ordered_filter_data_13_12 : OUT std_logic ;
         ordered_filter_data_13_11 : OUT std_logic ;
         ordered_filter_data_13_10 : OUT std_logic ;
         ordered_filter_data_13_9 : OUT std_logic ;
         ordered_filter_data_13_8 : OUT std_logic ;
         ordered_filter_data_13_7 : OUT std_logic ;
         ordered_filter_data_13_6 : OUT std_logic ;
         ordered_filter_data_13_5 : OUT std_logic ;
         ordered_filter_data_13_4 : OUT std_logic ;
         ordered_filter_data_13_3 : OUT std_logic ;
         ordered_filter_data_13_2 : OUT std_logic ;
         ordered_filter_data_13_1 : OUT std_logic ;
         ordered_filter_data_13_0 : OUT std_logic ;
         ordered_filter_data_14_31 : OUT std_logic ;
         ordered_filter_data_14_30 : OUT std_logic ;
         ordered_filter_data_14_29 : OUT std_logic ;
         ordered_filter_data_14_28 : OUT std_logic ;
         ordered_filter_data_14_27 : OUT std_logic ;
         ordered_filter_data_14_26 : OUT std_logic ;
         ordered_filter_data_14_25 : OUT std_logic ;
         ordered_filter_data_14_24 : OUT std_logic ;
         ordered_filter_data_14_23 : OUT std_logic ;
         ordered_filter_data_14_22 : OUT std_logic ;
         ordered_filter_data_14_21 : OUT std_logic ;
         ordered_filter_data_14_20 : OUT std_logic ;
         ordered_filter_data_14_19 : OUT std_logic ;
         ordered_filter_data_14_18 : OUT std_logic ;
         ordered_filter_data_14_17 : OUT std_logic ;
         ordered_filter_data_14_16 : OUT std_logic ;
         ordered_filter_data_14_15 : OUT std_logic ;
         ordered_filter_data_14_14 : OUT std_logic ;
         ordered_filter_data_14_13 : OUT std_logic ;
         ordered_filter_data_14_12 : OUT std_logic ;
         ordered_filter_data_14_11 : OUT std_logic ;
         ordered_filter_data_14_10 : OUT std_logic ;
         ordered_filter_data_14_9 : OUT std_logic ;
         ordered_filter_data_14_8 : OUT std_logic ;
         ordered_filter_data_14_7 : OUT std_logic ;
         ordered_filter_data_14_6 : OUT std_logic ;
         ordered_filter_data_14_5 : OUT std_logic ;
         ordered_filter_data_14_4 : OUT std_logic ;
         ordered_filter_data_14_3 : OUT std_logic ;
         ordered_filter_data_14_2 : OUT std_logic ;
         ordered_filter_data_14_1 : OUT std_logic ;
         ordered_filter_data_14_0 : OUT std_logic ;
         ordered_filter_data_15_31 : OUT std_logic ;
         ordered_filter_data_15_30 : OUT std_logic ;
         ordered_filter_data_15_29 : OUT std_logic ;
         ordered_filter_data_15_28 : OUT std_logic ;
         ordered_filter_data_15_27 : OUT std_logic ;
         ordered_filter_data_15_26 : OUT std_logic ;
         ordered_filter_data_15_25 : OUT std_logic ;
         ordered_filter_data_15_24 : OUT std_logic ;
         ordered_filter_data_15_23 : OUT std_logic ;
         ordered_filter_data_15_22 : OUT std_logic ;
         ordered_filter_data_15_21 : OUT std_logic ;
         ordered_filter_data_15_20 : OUT std_logic ;
         ordered_filter_data_15_19 : OUT std_logic ;
         ordered_filter_data_15_18 : OUT std_logic ;
         ordered_filter_data_15_17 : OUT std_logic ;
         ordered_filter_data_15_16 : OUT std_logic ;
         ordered_filter_data_15_15 : OUT std_logic ;
         ordered_filter_data_15_14 : OUT std_logic ;
         ordered_filter_data_15_13 : OUT std_logic ;
         ordered_filter_data_15_12 : OUT std_logic ;
         ordered_filter_data_15_11 : OUT std_logic ;
         ordered_filter_data_15_10 : OUT std_logic ;
         ordered_filter_data_15_9 : OUT std_logic ;
         ordered_filter_data_15_8 : OUT std_logic ;
         ordered_filter_data_15_7 : OUT std_logic ;
         ordered_filter_data_15_6 : OUT std_logic ;
         ordered_filter_data_15_5 : OUT std_logic ;
         ordered_filter_data_15_4 : OUT std_logic ;
         ordered_filter_data_15_3 : OUT std_logic ;
         ordered_filter_data_15_2 : OUT std_logic ;
         ordered_filter_data_15_1 : OUT std_logic ;
         ordered_filter_data_15_0 : OUT std_logic ;
         ordered_filter_data_16_31 : OUT std_logic ;
         ordered_filter_data_16_30 : OUT std_logic ;
         ordered_filter_data_16_29 : OUT std_logic ;
         ordered_filter_data_16_28 : OUT std_logic ;
         ordered_filter_data_16_27 : OUT std_logic ;
         ordered_filter_data_16_26 : OUT std_logic ;
         ordered_filter_data_16_25 : OUT std_logic ;
         ordered_filter_data_16_24 : OUT std_logic ;
         ordered_filter_data_16_23 : OUT std_logic ;
         ordered_filter_data_16_22 : OUT std_logic ;
         ordered_filter_data_16_21 : OUT std_logic ;
         ordered_filter_data_16_20 : OUT std_logic ;
         ordered_filter_data_16_19 : OUT std_logic ;
         ordered_filter_data_16_18 : OUT std_logic ;
         ordered_filter_data_16_17 : OUT std_logic ;
         ordered_filter_data_16_16 : OUT std_logic ;
         ordered_filter_data_16_15 : OUT std_logic ;
         ordered_filter_data_16_14 : OUT std_logic ;
         ordered_filter_data_16_13 : OUT std_logic ;
         ordered_filter_data_16_12 : OUT std_logic ;
         ordered_filter_data_16_11 : OUT std_logic ;
         ordered_filter_data_16_10 : OUT std_logic ;
         ordered_filter_data_16_9 : OUT std_logic ;
         ordered_filter_data_16_8 : OUT std_logic ;
         ordered_filter_data_16_7 : OUT std_logic ;
         ordered_filter_data_16_6 : OUT std_logic ;
         ordered_filter_data_16_5 : OUT std_logic ;
         ordered_filter_data_16_4 : OUT std_logic ;
         ordered_filter_data_16_3 : OUT std_logic ;
         ordered_filter_data_16_2 : OUT std_logic ;
         ordered_filter_data_16_1 : OUT std_logic ;
         ordered_filter_data_16_0 : OUT std_logic ;
         ordered_filter_data_17_31 : OUT std_logic ;
         ordered_filter_data_17_30 : OUT std_logic ;
         ordered_filter_data_17_29 : OUT std_logic ;
         ordered_filter_data_17_28 : OUT std_logic ;
         ordered_filter_data_17_27 : OUT std_logic ;
         ordered_filter_data_17_26 : OUT std_logic ;
         ordered_filter_data_17_25 : OUT std_logic ;
         ordered_filter_data_17_24 : OUT std_logic ;
         ordered_filter_data_17_23 : OUT std_logic ;
         ordered_filter_data_17_22 : OUT std_logic ;
         ordered_filter_data_17_21 : OUT std_logic ;
         ordered_filter_data_17_20 : OUT std_logic ;
         ordered_filter_data_17_19 : OUT std_logic ;
         ordered_filter_data_17_18 : OUT std_logic ;
         ordered_filter_data_17_17 : OUT std_logic ;
         ordered_filter_data_17_16 : OUT std_logic ;
         ordered_filter_data_17_15 : OUT std_logic ;
         ordered_filter_data_17_14 : OUT std_logic ;
         ordered_filter_data_17_13 : OUT std_logic ;
         ordered_filter_data_17_12 : OUT std_logic ;
         ordered_filter_data_17_11 : OUT std_logic ;
         ordered_filter_data_17_10 : OUT std_logic ;
         ordered_filter_data_17_9 : OUT std_logic ;
         ordered_filter_data_17_8 : OUT std_logic ;
         ordered_filter_data_17_7 : OUT std_logic ;
         ordered_filter_data_17_6 : OUT std_logic ;
         ordered_filter_data_17_5 : OUT std_logic ;
         ordered_filter_data_17_4 : OUT std_logic ;
         ordered_filter_data_17_3 : OUT std_logic ;
         ordered_filter_data_17_2 : OUT std_logic ;
         ordered_filter_data_17_1 : OUT std_logic ;
         ordered_filter_data_17_0 : OUT std_logic ;
         ordered_filter_data_18_31 : OUT std_logic ;
         ordered_filter_data_18_30 : OUT std_logic ;
         ordered_filter_data_18_29 : OUT std_logic ;
         ordered_filter_data_18_28 : OUT std_logic ;
         ordered_filter_data_18_27 : OUT std_logic ;
         ordered_filter_data_18_26 : OUT std_logic ;
         ordered_filter_data_18_25 : OUT std_logic ;
         ordered_filter_data_18_24 : OUT std_logic ;
         ordered_filter_data_18_23 : OUT std_logic ;
         ordered_filter_data_18_22 : OUT std_logic ;
         ordered_filter_data_18_21 : OUT std_logic ;
         ordered_filter_data_18_20 : OUT std_logic ;
         ordered_filter_data_18_19 : OUT std_logic ;
         ordered_filter_data_18_18 : OUT std_logic ;
         ordered_filter_data_18_17 : OUT std_logic ;
         ordered_filter_data_18_16 : OUT std_logic ;
         ordered_filter_data_18_15 : OUT std_logic ;
         ordered_filter_data_18_14 : OUT std_logic ;
         ordered_filter_data_18_13 : OUT std_logic ;
         ordered_filter_data_18_12 : OUT std_logic ;
         ordered_filter_data_18_11 : OUT std_logic ;
         ordered_filter_data_18_10 : OUT std_logic ;
         ordered_filter_data_18_9 : OUT std_logic ;
         ordered_filter_data_18_8 : OUT std_logic ;
         ordered_filter_data_18_7 : OUT std_logic ;
         ordered_filter_data_18_6 : OUT std_logic ;
         ordered_filter_data_18_5 : OUT std_logic ;
         ordered_filter_data_18_4 : OUT std_logic ;
         ordered_filter_data_18_3 : OUT std_logic ;
         ordered_filter_data_18_2 : OUT std_logic ;
         ordered_filter_data_18_1 : OUT std_logic ;
         ordered_filter_data_18_0 : OUT std_logic ;
         ordered_filter_data_19_31 : OUT std_logic ;
         ordered_filter_data_19_30 : OUT std_logic ;
         ordered_filter_data_19_29 : OUT std_logic ;
         ordered_filter_data_19_28 : OUT std_logic ;
         ordered_filter_data_19_27 : OUT std_logic ;
         ordered_filter_data_19_26 : OUT std_logic ;
         ordered_filter_data_19_25 : OUT std_logic ;
         ordered_filter_data_19_24 : OUT std_logic ;
         ordered_filter_data_19_23 : OUT std_logic ;
         ordered_filter_data_19_22 : OUT std_logic ;
         ordered_filter_data_19_21 : OUT std_logic ;
         ordered_filter_data_19_20 : OUT std_logic ;
         ordered_filter_data_19_19 : OUT std_logic ;
         ordered_filter_data_19_18 : OUT std_logic ;
         ordered_filter_data_19_17 : OUT std_logic ;
         ordered_filter_data_19_16 : OUT std_logic ;
         ordered_filter_data_19_15 : OUT std_logic ;
         ordered_filter_data_19_14 : OUT std_logic ;
         ordered_filter_data_19_13 : OUT std_logic ;
         ordered_filter_data_19_12 : OUT std_logic ;
         ordered_filter_data_19_11 : OUT std_logic ;
         ordered_filter_data_19_10 : OUT std_logic ;
         ordered_filter_data_19_9 : OUT std_logic ;
         ordered_filter_data_19_8 : OUT std_logic ;
         ordered_filter_data_19_7 : OUT std_logic ;
         ordered_filter_data_19_6 : OUT std_logic ;
         ordered_filter_data_19_5 : OUT std_logic ;
         ordered_filter_data_19_4 : OUT std_logic ;
         ordered_filter_data_19_3 : OUT std_logic ;
         ordered_filter_data_19_2 : OUT std_logic ;
         ordered_filter_data_19_1 : OUT std_logic ;
         ordered_filter_data_19_0 : OUT std_logic ;
         ordered_filter_data_20_31 : OUT std_logic ;
         ordered_filter_data_20_30 : OUT std_logic ;
         ordered_filter_data_20_29 : OUT std_logic ;
         ordered_filter_data_20_28 : OUT std_logic ;
         ordered_filter_data_20_27 : OUT std_logic ;
         ordered_filter_data_20_26 : OUT std_logic ;
         ordered_filter_data_20_25 : OUT std_logic ;
         ordered_filter_data_20_24 : OUT std_logic ;
         ordered_filter_data_20_23 : OUT std_logic ;
         ordered_filter_data_20_22 : OUT std_logic ;
         ordered_filter_data_20_21 : OUT std_logic ;
         ordered_filter_data_20_20 : OUT std_logic ;
         ordered_filter_data_20_19 : OUT std_logic ;
         ordered_filter_data_20_18 : OUT std_logic ;
         ordered_filter_data_20_17 : OUT std_logic ;
         ordered_filter_data_20_16 : OUT std_logic ;
         ordered_filter_data_20_15 : OUT std_logic ;
         ordered_filter_data_20_14 : OUT std_logic ;
         ordered_filter_data_20_13 : OUT std_logic ;
         ordered_filter_data_20_12 : OUT std_logic ;
         ordered_filter_data_20_11 : OUT std_logic ;
         ordered_filter_data_20_10 : OUT std_logic ;
         ordered_filter_data_20_9 : OUT std_logic ;
         ordered_filter_data_20_8 : OUT std_logic ;
         ordered_filter_data_20_7 : OUT std_logic ;
         ordered_filter_data_20_6 : OUT std_logic ;
         ordered_filter_data_20_5 : OUT std_logic ;
         ordered_filter_data_20_4 : OUT std_logic ;
         ordered_filter_data_20_3 : OUT std_logic ;
         ordered_filter_data_20_2 : OUT std_logic ;
         ordered_filter_data_20_1 : OUT std_logic ;
         ordered_filter_data_20_0 : OUT std_logic ;
         ordered_filter_data_21_31 : OUT std_logic ;
         ordered_filter_data_21_30 : OUT std_logic ;
         ordered_filter_data_21_29 : OUT std_logic ;
         ordered_filter_data_21_28 : OUT std_logic ;
         ordered_filter_data_21_27 : OUT std_logic ;
         ordered_filter_data_21_26 : OUT std_logic ;
         ordered_filter_data_21_25 : OUT std_logic ;
         ordered_filter_data_21_24 : OUT std_logic ;
         ordered_filter_data_21_23 : OUT std_logic ;
         ordered_filter_data_21_22 : OUT std_logic ;
         ordered_filter_data_21_21 : OUT std_logic ;
         ordered_filter_data_21_20 : OUT std_logic ;
         ordered_filter_data_21_19 : OUT std_logic ;
         ordered_filter_data_21_18 : OUT std_logic ;
         ordered_filter_data_21_17 : OUT std_logic ;
         ordered_filter_data_21_16 : OUT std_logic ;
         ordered_filter_data_21_15 : OUT std_logic ;
         ordered_filter_data_21_14 : OUT std_logic ;
         ordered_filter_data_21_13 : OUT std_logic ;
         ordered_filter_data_21_12 : OUT std_logic ;
         ordered_filter_data_21_11 : OUT std_logic ;
         ordered_filter_data_21_10 : OUT std_logic ;
         ordered_filter_data_21_9 : OUT std_logic ;
         ordered_filter_data_21_8 : OUT std_logic ;
         ordered_filter_data_21_7 : OUT std_logic ;
         ordered_filter_data_21_6 : OUT std_logic ;
         ordered_filter_data_21_5 : OUT std_logic ;
         ordered_filter_data_21_4 : OUT std_logic ;
         ordered_filter_data_21_3 : OUT std_logic ;
         ordered_filter_data_21_2 : OUT std_logic ;
         ordered_filter_data_21_1 : OUT std_logic ;
         ordered_filter_data_21_0 : OUT std_logic ;
         ordered_filter_data_22_31 : OUT std_logic ;
         ordered_filter_data_22_30 : OUT std_logic ;
         ordered_filter_data_22_29 : OUT std_logic ;
         ordered_filter_data_22_28 : OUT std_logic ;
         ordered_filter_data_22_27 : OUT std_logic ;
         ordered_filter_data_22_26 : OUT std_logic ;
         ordered_filter_data_22_25 : OUT std_logic ;
         ordered_filter_data_22_24 : OUT std_logic ;
         ordered_filter_data_22_23 : OUT std_logic ;
         ordered_filter_data_22_22 : OUT std_logic ;
         ordered_filter_data_22_21 : OUT std_logic ;
         ordered_filter_data_22_20 : OUT std_logic ;
         ordered_filter_data_22_19 : OUT std_logic ;
         ordered_filter_data_22_18 : OUT std_logic ;
         ordered_filter_data_22_17 : OUT std_logic ;
         ordered_filter_data_22_16 : OUT std_logic ;
         ordered_filter_data_22_15 : OUT std_logic ;
         ordered_filter_data_22_14 : OUT std_logic ;
         ordered_filter_data_22_13 : OUT std_logic ;
         ordered_filter_data_22_12 : OUT std_logic ;
         ordered_filter_data_22_11 : OUT std_logic ;
         ordered_filter_data_22_10 : OUT std_logic ;
         ordered_filter_data_22_9 : OUT std_logic ;
         ordered_filter_data_22_8 : OUT std_logic ;
         ordered_filter_data_22_7 : OUT std_logic ;
         ordered_filter_data_22_6 : OUT std_logic ;
         ordered_filter_data_22_5 : OUT std_logic ;
         ordered_filter_data_22_4 : OUT std_logic ;
         ordered_filter_data_22_3 : OUT std_logic ;
         ordered_filter_data_22_2 : OUT std_logic ;
         ordered_filter_data_22_1 : OUT std_logic ;
         ordered_filter_data_22_0 : OUT std_logic ;
         ordered_filter_data_23_31 : OUT std_logic ;
         ordered_filter_data_23_30 : OUT std_logic ;
         ordered_filter_data_23_29 : OUT std_logic ;
         ordered_filter_data_23_28 : OUT std_logic ;
         ordered_filter_data_23_27 : OUT std_logic ;
         ordered_filter_data_23_26 : OUT std_logic ;
         ordered_filter_data_23_25 : OUT std_logic ;
         ordered_filter_data_23_24 : OUT std_logic ;
         ordered_filter_data_23_23 : OUT std_logic ;
         ordered_filter_data_23_22 : OUT std_logic ;
         ordered_filter_data_23_21 : OUT std_logic ;
         ordered_filter_data_23_20 : OUT std_logic ;
         ordered_filter_data_23_19 : OUT std_logic ;
         ordered_filter_data_23_18 : OUT std_logic ;
         ordered_filter_data_23_17 : OUT std_logic ;
         ordered_filter_data_23_16 : OUT std_logic ;
         ordered_filter_data_23_15 : OUT std_logic ;
         ordered_filter_data_23_14 : OUT std_logic ;
         ordered_filter_data_23_13 : OUT std_logic ;
         ordered_filter_data_23_12 : OUT std_logic ;
         ordered_filter_data_23_11 : OUT std_logic ;
         ordered_filter_data_23_10 : OUT std_logic ;
         ordered_filter_data_23_9 : OUT std_logic ;
         ordered_filter_data_23_8 : OUT std_logic ;
         ordered_filter_data_23_7 : OUT std_logic ;
         ordered_filter_data_23_6 : OUT std_logic ;
         ordered_filter_data_23_5 : OUT std_logic ;
         ordered_filter_data_23_4 : OUT std_logic ;
         ordered_filter_data_23_3 : OUT std_logic ;
         ordered_filter_data_23_2 : OUT std_logic ;
         ordered_filter_data_23_1 : OUT std_logic ;
         ordered_filter_data_23_0 : OUT std_logic ;
         ordered_filter_data_24_31 : OUT std_logic ;
         ordered_filter_data_24_30 : OUT std_logic ;
         ordered_filter_data_24_29 : OUT std_logic ;
         ordered_filter_data_24_28 : OUT std_logic ;
         ordered_filter_data_24_27 : OUT std_logic ;
         ordered_filter_data_24_26 : OUT std_logic ;
         ordered_filter_data_24_25 : OUT std_logic ;
         ordered_filter_data_24_24 : OUT std_logic ;
         ordered_filter_data_24_23 : OUT std_logic ;
         ordered_filter_data_24_22 : OUT std_logic ;
         ordered_filter_data_24_21 : OUT std_logic ;
         ordered_filter_data_24_20 : OUT std_logic ;
         ordered_filter_data_24_19 : OUT std_logic ;
         ordered_filter_data_24_18 : OUT std_logic ;
         ordered_filter_data_24_17 : OUT std_logic ;
         ordered_filter_data_24_16 : OUT std_logic ;
         ordered_filter_data_24_15 : OUT std_logic ;
         ordered_filter_data_24_14 : OUT std_logic ;
         ordered_filter_data_24_13 : OUT std_logic ;
         ordered_filter_data_24_12 : OUT std_logic ;
         ordered_filter_data_24_11 : OUT std_logic ;
         ordered_filter_data_24_10 : OUT std_logic ;
         ordered_filter_data_24_9 : OUT std_logic ;
         ordered_filter_data_24_8 : OUT std_logic ;
         ordered_filter_data_24_7 : OUT std_logic ;
         ordered_filter_data_24_6 : OUT std_logic ;
         ordered_filter_data_24_5 : OUT std_logic ;
         ordered_filter_data_24_4 : OUT std_logic ;
         ordered_filter_data_24_3 : OUT std_logic ;
         ordered_filter_data_24_2 : OUT std_logic ;
         ordered_filter_data_24_1 : OUT std_logic ;
         ordered_filter_data_24_0 : OUT std_logic) ;
   end component ;
   component MergeLayer
      port (
         d_arr_0_31 : OUT std_logic ;
         d_arr_0_30 : OUT std_logic ;
         d_arr_0_29 : OUT std_logic ;
         d_arr_0_28 : OUT std_logic ;
         d_arr_0_27 : OUT std_logic ;
         d_arr_0_26 : OUT std_logic ;
         d_arr_0_25 : OUT std_logic ;
         d_arr_0_24 : OUT std_logic ;
         d_arr_0_23 : OUT std_logic ;
         d_arr_0_22 : OUT std_logic ;
         d_arr_0_21 : OUT std_logic ;
         d_arr_0_20 : OUT std_logic ;
         d_arr_0_19 : OUT std_logic ;
         d_arr_0_18 : OUT std_logic ;
         d_arr_0_17 : OUT std_logic ;
         d_arr_0_16 : OUT std_logic ;
         d_arr_0_15 : OUT std_logic ;
         d_arr_0_14 : OUT std_logic ;
         d_arr_0_13 : OUT std_logic ;
         d_arr_0_12 : OUT std_logic ;
         d_arr_0_11 : OUT std_logic ;
         d_arr_0_10 : OUT std_logic ;
         d_arr_0_9 : OUT std_logic ;
         d_arr_0_8 : OUT std_logic ;
         d_arr_0_7 : OUT std_logic ;
         d_arr_0_6 : OUT std_logic ;
         d_arr_0_5 : OUT std_logic ;
         d_arr_0_4 : OUT std_logic ;
         d_arr_0_3 : OUT std_logic ;
         d_arr_0_2 : OUT std_logic ;
         d_arr_0_1 : OUT std_logic ;
         d_arr_0_0 : OUT std_logic ;
         d_arr_1_31 : OUT std_logic ;
         d_arr_1_30 : OUT std_logic ;
         d_arr_1_29 : OUT std_logic ;
         d_arr_1_28 : OUT std_logic ;
         d_arr_1_27 : OUT std_logic ;
         d_arr_1_26 : OUT std_logic ;
         d_arr_1_25 : OUT std_logic ;
         d_arr_1_24 : OUT std_logic ;
         d_arr_1_23 : OUT std_logic ;
         d_arr_1_22 : OUT std_logic ;
         d_arr_1_21 : OUT std_logic ;
         d_arr_1_20 : OUT std_logic ;
         d_arr_1_19 : OUT std_logic ;
         d_arr_1_18 : OUT std_logic ;
         d_arr_1_17 : OUT std_logic ;
         d_arr_1_16 : OUT std_logic ;
         d_arr_1_15 : OUT std_logic ;
         d_arr_1_14 : OUT std_logic ;
         d_arr_1_13 : OUT std_logic ;
         d_arr_1_12 : OUT std_logic ;
         d_arr_1_11 : OUT std_logic ;
         d_arr_1_10 : OUT std_logic ;
         d_arr_1_9 : OUT std_logic ;
         d_arr_1_8 : OUT std_logic ;
         d_arr_1_7 : OUT std_logic ;
         d_arr_1_6 : OUT std_logic ;
         d_arr_1_5 : OUT std_logic ;
         d_arr_1_4 : OUT std_logic ;
         d_arr_1_3 : OUT std_logic ;
         d_arr_1_2 : OUT std_logic ;
         d_arr_1_1 : OUT std_logic ;
         d_arr_1_0 : OUT std_logic ;
         d_arr_2_31 : OUT std_logic ;
         d_arr_2_30 : OUT std_logic ;
         d_arr_2_29 : OUT std_logic ;
         d_arr_2_28 : OUT std_logic ;
         d_arr_2_27 : OUT std_logic ;
         d_arr_2_26 : OUT std_logic ;
         d_arr_2_25 : OUT std_logic ;
         d_arr_2_24 : OUT std_logic ;
         d_arr_2_23 : OUT std_logic ;
         d_arr_2_22 : OUT std_logic ;
         d_arr_2_21 : OUT std_logic ;
         d_arr_2_20 : OUT std_logic ;
         d_arr_2_19 : OUT std_logic ;
         d_arr_2_18 : OUT std_logic ;
         d_arr_2_17 : OUT std_logic ;
         d_arr_2_16 : OUT std_logic ;
         d_arr_2_15 : OUT std_logic ;
         d_arr_2_14 : OUT std_logic ;
         d_arr_2_13 : OUT std_logic ;
         d_arr_2_12 : OUT std_logic ;
         d_arr_2_11 : OUT std_logic ;
         d_arr_2_10 : OUT std_logic ;
         d_arr_2_9 : OUT std_logic ;
         d_arr_2_8 : OUT std_logic ;
         d_arr_2_7 : OUT std_logic ;
         d_arr_2_6 : OUT std_logic ;
         d_arr_2_5 : OUT std_logic ;
         d_arr_2_4 : OUT std_logic ;
         d_arr_2_3 : OUT std_logic ;
         d_arr_2_2 : OUT std_logic ;
         d_arr_2_1 : OUT std_logic ;
         d_arr_2_0 : OUT std_logic ;
         d_arr_3_31 : OUT std_logic ;
         d_arr_3_30 : OUT std_logic ;
         d_arr_3_29 : OUT std_logic ;
         d_arr_3_28 : OUT std_logic ;
         d_arr_3_27 : OUT std_logic ;
         d_arr_3_26 : OUT std_logic ;
         d_arr_3_25 : OUT std_logic ;
         d_arr_3_24 : OUT std_logic ;
         d_arr_3_23 : OUT std_logic ;
         d_arr_3_22 : OUT std_logic ;
         d_arr_3_21 : OUT std_logic ;
         d_arr_3_20 : OUT std_logic ;
         d_arr_3_19 : OUT std_logic ;
         d_arr_3_18 : OUT std_logic ;
         d_arr_3_17 : OUT std_logic ;
         d_arr_3_16 : OUT std_logic ;
         d_arr_3_15 : OUT std_logic ;
         d_arr_3_14 : OUT std_logic ;
         d_arr_3_13 : OUT std_logic ;
         d_arr_3_12 : OUT std_logic ;
         d_arr_3_11 : OUT std_logic ;
         d_arr_3_10 : OUT std_logic ;
         d_arr_3_9 : OUT std_logic ;
         d_arr_3_8 : OUT std_logic ;
         d_arr_3_7 : OUT std_logic ;
         d_arr_3_6 : OUT std_logic ;
         d_arr_3_5 : OUT std_logic ;
         d_arr_3_4 : OUT std_logic ;
         d_arr_3_3 : OUT std_logic ;
         d_arr_3_2 : OUT std_logic ;
         d_arr_3_1 : OUT std_logic ;
         d_arr_3_0 : OUT std_logic ;
         d_arr_4_31 : OUT std_logic ;
         d_arr_4_30 : OUT std_logic ;
         d_arr_4_29 : OUT std_logic ;
         d_arr_4_28 : OUT std_logic ;
         d_arr_4_27 : OUT std_logic ;
         d_arr_4_26 : OUT std_logic ;
         d_arr_4_25 : OUT std_logic ;
         d_arr_4_24 : OUT std_logic ;
         d_arr_4_23 : OUT std_logic ;
         d_arr_4_22 : OUT std_logic ;
         d_arr_4_21 : OUT std_logic ;
         d_arr_4_20 : OUT std_logic ;
         d_arr_4_19 : OUT std_logic ;
         d_arr_4_18 : OUT std_logic ;
         d_arr_4_17 : OUT std_logic ;
         d_arr_4_16 : OUT std_logic ;
         d_arr_4_15 : OUT std_logic ;
         d_arr_4_14 : OUT std_logic ;
         d_arr_4_13 : OUT std_logic ;
         d_arr_4_12 : OUT std_logic ;
         d_arr_4_11 : OUT std_logic ;
         d_arr_4_10 : OUT std_logic ;
         d_arr_4_9 : OUT std_logic ;
         d_arr_4_8 : OUT std_logic ;
         d_arr_4_7 : OUT std_logic ;
         d_arr_4_6 : OUT std_logic ;
         d_arr_4_5 : OUT std_logic ;
         d_arr_4_4 : OUT std_logic ;
         d_arr_4_3 : OUT std_logic ;
         d_arr_4_2 : OUT std_logic ;
         d_arr_4_1 : OUT std_logic ;
         d_arr_4_0 : OUT std_logic ;
         d_arr_5_31 : OUT std_logic ;
         d_arr_5_30 : OUT std_logic ;
         d_arr_5_29 : OUT std_logic ;
         d_arr_5_28 : OUT std_logic ;
         d_arr_5_27 : OUT std_logic ;
         d_arr_5_26 : OUT std_logic ;
         d_arr_5_25 : OUT std_logic ;
         d_arr_5_24 : OUT std_logic ;
         d_arr_5_23 : OUT std_logic ;
         d_arr_5_22 : OUT std_logic ;
         d_arr_5_21 : OUT std_logic ;
         d_arr_5_20 : OUT std_logic ;
         d_arr_5_19 : OUT std_logic ;
         d_arr_5_18 : OUT std_logic ;
         d_arr_5_17 : OUT std_logic ;
         d_arr_5_16 : OUT std_logic ;
         d_arr_5_15 : OUT std_logic ;
         d_arr_5_14 : OUT std_logic ;
         d_arr_5_13 : OUT std_logic ;
         d_arr_5_12 : OUT std_logic ;
         d_arr_5_11 : OUT std_logic ;
         d_arr_5_10 : OUT std_logic ;
         d_arr_5_9 : OUT std_logic ;
         d_arr_5_8 : OUT std_logic ;
         d_arr_5_7 : OUT std_logic ;
         d_arr_5_6 : OUT std_logic ;
         d_arr_5_5 : OUT std_logic ;
         d_arr_5_4 : OUT std_logic ;
         d_arr_5_3 : OUT std_logic ;
         d_arr_5_2 : OUT std_logic ;
         d_arr_5_1 : OUT std_logic ;
         d_arr_5_0 : OUT std_logic ;
         d_arr_6_31 : OUT std_logic ;
         d_arr_6_30 : OUT std_logic ;
         d_arr_6_29 : OUT std_logic ;
         d_arr_6_28 : OUT std_logic ;
         d_arr_6_27 : OUT std_logic ;
         d_arr_6_26 : OUT std_logic ;
         d_arr_6_25 : OUT std_logic ;
         d_arr_6_24 : OUT std_logic ;
         d_arr_6_23 : OUT std_logic ;
         d_arr_6_22 : OUT std_logic ;
         d_arr_6_21 : OUT std_logic ;
         d_arr_6_20 : OUT std_logic ;
         d_arr_6_19 : OUT std_logic ;
         d_arr_6_18 : OUT std_logic ;
         d_arr_6_17 : OUT std_logic ;
         d_arr_6_16 : OUT std_logic ;
         d_arr_6_15 : OUT std_logic ;
         d_arr_6_14 : OUT std_logic ;
         d_arr_6_13 : OUT std_logic ;
         d_arr_6_12 : OUT std_logic ;
         d_arr_6_11 : OUT std_logic ;
         d_arr_6_10 : OUT std_logic ;
         d_arr_6_9 : OUT std_logic ;
         d_arr_6_8 : OUT std_logic ;
         d_arr_6_7 : OUT std_logic ;
         d_arr_6_6 : OUT std_logic ;
         d_arr_6_5 : OUT std_logic ;
         d_arr_6_4 : OUT std_logic ;
         d_arr_6_3 : OUT std_logic ;
         d_arr_6_2 : OUT std_logic ;
         d_arr_6_1 : OUT std_logic ;
         d_arr_6_0 : OUT std_logic ;
         d_arr_7_31 : OUT std_logic ;
         d_arr_7_30 : OUT std_logic ;
         d_arr_7_29 : OUT std_logic ;
         d_arr_7_28 : OUT std_logic ;
         d_arr_7_27 : OUT std_logic ;
         d_arr_7_26 : OUT std_logic ;
         d_arr_7_25 : OUT std_logic ;
         d_arr_7_24 : OUT std_logic ;
         d_arr_7_23 : OUT std_logic ;
         d_arr_7_22 : OUT std_logic ;
         d_arr_7_21 : OUT std_logic ;
         d_arr_7_20 : OUT std_logic ;
         d_arr_7_19 : OUT std_logic ;
         d_arr_7_18 : OUT std_logic ;
         d_arr_7_17 : OUT std_logic ;
         d_arr_7_16 : OUT std_logic ;
         d_arr_7_15 : OUT std_logic ;
         d_arr_7_14 : OUT std_logic ;
         d_arr_7_13 : OUT std_logic ;
         d_arr_7_12 : OUT std_logic ;
         d_arr_7_11 : OUT std_logic ;
         d_arr_7_10 : OUT std_logic ;
         d_arr_7_9 : OUT std_logic ;
         d_arr_7_8 : OUT std_logic ;
         d_arr_7_7 : OUT std_logic ;
         d_arr_7_6 : OUT std_logic ;
         d_arr_7_5 : OUT std_logic ;
         d_arr_7_4 : OUT std_logic ;
         d_arr_7_3 : OUT std_logic ;
         d_arr_7_2 : OUT std_logic ;
         d_arr_7_1 : OUT std_logic ;
         d_arr_7_0 : OUT std_logic ;
         d_arr_8_31 : OUT std_logic ;
         d_arr_8_30 : OUT std_logic ;
         d_arr_8_29 : OUT std_logic ;
         d_arr_8_28 : OUT std_logic ;
         d_arr_8_27 : OUT std_logic ;
         d_arr_8_26 : OUT std_logic ;
         d_arr_8_25 : OUT std_logic ;
         d_arr_8_24 : OUT std_logic ;
         d_arr_8_23 : OUT std_logic ;
         d_arr_8_22 : OUT std_logic ;
         d_arr_8_21 : OUT std_logic ;
         d_arr_8_20 : OUT std_logic ;
         d_arr_8_19 : OUT std_logic ;
         d_arr_8_18 : OUT std_logic ;
         d_arr_8_17 : OUT std_logic ;
         d_arr_8_16 : OUT std_logic ;
         d_arr_8_15 : OUT std_logic ;
         d_arr_8_14 : OUT std_logic ;
         d_arr_8_13 : OUT std_logic ;
         d_arr_8_12 : OUT std_logic ;
         d_arr_8_11 : OUT std_logic ;
         d_arr_8_10 : OUT std_logic ;
         d_arr_8_9 : OUT std_logic ;
         d_arr_8_8 : OUT std_logic ;
         d_arr_8_7 : OUT std_logic ;
         d_arr_8_6 : OUT std_logic ;
         d_arr_8_5 : OUT std_logic ;
         d_arr_8_4 : OUT std_logic ;
         d_arr_8_3 : OUT std_logic ;
         d_arr_8_2 : OUT std_logic ;
         d_arr_8_1 : OUT std_logic ;
         d_arr_8_0 : OUT std_logic ;
         d_arr_9_31 : OUT std_logic ;
         d_arr_9_30 : OUT std_logic ;
         d_arr_9_29 : OUT std_logic ;
         d_arr_9_28 : OUT std_logic ;
         d_arr_9_27 : OUT std_logic ;
         d_arr_9_26 : OUT std_logic ;
         d_arr_9_25 : OUT std_logic ;
         d_arr_9_24 : OUT std_logic ;
         d_arr_9_23 : OUT std_logic ;
         d_arr_9_22 : OUT std_logic ;
         d_arr_9_21 : OUT std_logic ;
         d_arr_9_20 : OUT std_logic ;
         d_arr_9_19 : OUT std_logic ;
         d_arr_9_18 : OUT std_logic ;
         d_arr_9_17 : OUT std_logic ;
         d_arr_9_16 : OUT std_logic ;
         d_arr_9_15 : OUT std_logic ;
         d_arr_9_14 : OUT std_logic ;
         d_arr_9_13 : OUT std_logic ;
         d_arr_9_12 : OUT std_logic ;
         d_arr_9_11 : OUT std_logic ;
         d_arr_9_10 : OUT std_logic ;
         d_arr_9_9 : OUT std_logic ;
         d_arr_9_8 : OUT std_logic ;
         d_arr_9_7 : OUT std_logic ;
         d_arr_9_6 : OUT std_logic ;
         d_arr_9_5 : OUT std_logic ;
         d_arr_9_4 : OUT std_logic ;
         d_arr_9_3 : OUT std_logic ;
         d_arr_9_2 : OUT std_logic ;
         d_arr_9_1 : OUT std_logic ;
         d_arr_9_0 : OUT std_logic ;
         d_arr_10_31 : OUT std_logic ;
         d_arr_10_30 : OUT std_logic ;
         d_arr_10_29 : OUT std_logic ;
         d_arr_10_28 : OUT std_logic ;
         d_arr_10_27 : OUT std_logic ;
         d_arr_10_26 : OUT std_logic ;
         d_arr_10_25 : OUT std_logic ;
         d_arr_10_24 : OUT std_logic ;
         d_arr_10_23 : OUT std_logic ;
         d_arr_10_22 : OUT std_logic ;
         d_arr_10_21 : OUT std_logic ;
         d_arr_10_20 : OUT std_logic ;
         d_arr_10_19 : OUT std_logic ;
         d_arr_10_18 : OUT std_logic ;
         d_arr_10_17 : OUT std_logic ;
         d_arr_10_16 : OUT std_logic ;
         d_arr_10_15 : OUT std_logic ;
         d_arr_10_14 : OUT std_logic ;
         d_arr_10_13 : OUT std_logic ;
         d_arr_10_12 : OUT std_logic ;
         d_arr_10_11 : OUT std_logic ;
         d_arr_10_10 : OUT std_logic ;
         d_arr_10_9 : OUT std_logic ;
         d_arr_10_8 : OUT std_logic ;
         d_arr_10_7 : OUT std_logic ;
         d_arr_10_6 : OUT std_logic ;
         d_arr_10_5 : OUT std_logic ;
         d_arr_10_4 : OUT std_logic ;
         d_arr_10_3 : OUT std_logic ;
         d_arr_10_2 : OUT std_logic ;
         d_arr_10_1 : OUT std_logic ;
         d_arr_10_0 : OUT std_logic ;
         d_arr_11_31 : OUT std_logic ;
         d_arr_11_30 : OUT std_logic ;
         d_arr_11_29 : OUT std_logic ;
         d_arr_11_28 : OUT std_logic ;
         d_arr_11_27 : OUT std_logic ;
         d_arr_11_26 : OUT std_logic ;
         d_arr_11_25 : OUT std_logic ;
         d_arr_11_24 : OUT std_logic ;
         d_arr_11_23 : OUT std_logic ;
         d_arr_11_22 : OUT std_logic ;
         d_arr_11_21 : OUT std_logic ;
         d_arr_11_20 : OUT std_logic ;
         d_arr_11_19 : OUT std_logic ;
         d_arr_11_18 : OUT std_logic ;
         d_arr_11_17 : OUT std_logic ;
         d_arr_11_16 : OUT std_logic ;
         d_arr_11_15 : OUT std_logic ;
         d_arr_11_14 : OUT std_logic ;
         d_arr_11_13 : OUT std_logic ;
         d_arr_11_12 : OUT std_logic ;
         d_arr_11_11 : OUT std_logic ;
         d_arr_11_10 : OUT std_logic ;
         d_arr_11_9 : OUT std_logic ;
         d_arr_11_8 : OUT std_logic ;
         d_arr_11_7 : OUT std_logic ;
         d_arr_11_6 : OUT std_logic ;
         d_arr_11_5 : OUT std_logic ;
         d_arr_11_4 : OUT std_logic ;
         d_arr_11_3 : OUT std_logic ;
         d_arr_11_2 : OUT std_logic ;
         d_arr_11_1 : OUT std_logic ;
         d_arr_11_0 : OUT std_logic ;
         d_arr_12_31 : OUT std_logic ;
         d_arr_12_30 : OUT std_logic ;
         d_arr_12_29 : OUT std_logic ;
         d_arr_12_28 : OUT std_logic ;
         d_arr_12_27 : OUT std_logic ;
         d_arr_12_26 : OUT std_logic ;
         d_arr_12_25 : OUT std_logic ;
         d_arr_12_24 : OUT std_logic ;
         d_arr_12_23 : OUT std_logic ;
         d_arr_12_22 : OUT std_logic ;
         d_arr_12_21 : OUT std_logic ;
         d_arr_12_20 : OUT std_logic ;
         d_arr_12_19 : OUT std_logic ;
         d_arr_12_18 : OUT std_logic ;
         d_arr_12_17 : OUT std_logic ;
         d_arr_12_16 : OUT std_logic ;
         d_arr_12_15 : OUT std_logic ;
         d_arr_12_14 : OUT std_logic ;
         d_arr_12_13 : OUT std_logic ;
         d_arr_12_12 : OUT std_logic ;
         d_arr_12_11 : OUT std_logic ;
         d_arr_12_10 : OUT std_logic ;
         d_arr_12_9 : OUT std_logic ;
         d_arr_12_8 : OUT std_logic ;
         d_arr_12_7 : OUT std_logic ;
         d_arr_12_6 : OUT std_logic ;
         d_arr_12_5 : OUT std_logic ;
         d_arr_12_4 : OUT std_logic ;
         d_arr_12_3 : OUT std_logic ;
         d_arr_12_2 : OUT std_logic ;
         d_arr_12_1 : OUT std_logic ;
         d_arr_12_0 : OUT std_logic ;
         d_arr_13_31 : OUT std_logic ;
         d_arr_13_30 : OUT std_logic ;
         d_arr_13_29 : OUT std_logic ;
         d_arr_13_28 : OUT std_logic ;
         d_arr_13_27 : OUT std_logic ;
         d_arr_13_26 : OUT std_logic ;
         d_arr_13_25 : OUT std_logic ;
         d_arr_13_24 : OUT std_logic ;
         d_arr_13_23 : OUT std_logic ;
         d_arr_13_22 : OUT std_logic ;
         d_arr_13_21 : OUT std_logic ;
         d_arr_13_20 : OUT std_logic ;
         d_arr_13_19 : OUT std_logic ;
         d_arr_13_18 : OUT std_logic ;
         d_arr_13_17 : OUT std_logic ;
         d_arr_13_16 : OUT std_logic ;
         d_arr_13_15 : OUT std_logic ;
         d_arr_13_14 : OUT std_logic ;
         d_arr_13_13 : OUT std_logic ;
         d_arr_13_12 : OUT std_logic ;
         d_arr_13_11 : OUT std_logic ;
         d_arr_13_10 : OUT std_logic ;
         d_arr_13_9 : OUT std_logic ;
         d_arr_13_8 : OUT std_logic ;
         d_arr_13_7 : OUT std_logic ;
         d_arr_13_6 : OUT std_logic ;
         d_arr_13_5 : OUT std_logic ;
         d_arr_13_4 : OUT std_logic ;
         d_arr_13_3 : OUT std_logic ;
         d_arr_13_2 : OUT std_logic ;
         d_arr_13_1 : OUT std_logic ;
         d_arr_13_0 : OUT std_logic ;
         d_arr_14_31 : OUT std_logic ;
         d_arr_14_30 : OUT std_logic ;
         d_arr_14_29 : OUT std_logic ;
         d_arr_14_28 : OUT std_logic ;
         d_arr_14_27 : OUT std_logic ;
         d_arr_14_26 : OUT std_logic ;
         d_arr_14_25 : OUT std_logic ;
         d_arr_14_24 : OUT std_logic ;
         d_arr_14_23 : OUT std_logic ;
         d_arr_14_22 : OUT std_logic ;
         d_arr_14_21 : OUT std_logic ;
         d_arr_14_20 : OUT std_logic ;
         d_arr_14_19 : OUT std_logic ;
         d_arr_14_18 : OUT std_logic ;
         d_arr_14_17 : OUT std_logic ;
         d_arr_14_16 : OUT std_logic ;
         d_arr_14_15 : OUT std_logic ;
         d_arr_14_14 : OUT std_logic ;
         d_arr_14_13 : OUT std_logic ;
         d_arr_14_12 : OUT std_logic ;
         d_arr_14_11 : OUT std_logic ;
         d_arr_14_10 : OUT std_logic ;
         d_arr_14_9 : OUT std_logic ;
         d_arr_14_8 : OUT std_logic ;
         d_arr_14_7 : OUT std_logic ;
         d_arr_14_6 : OUT std_logic ;
         d_arr_14_5 : OUT std_logic ;
         d_arr_14_4 : OUT std_logic ;
         d_arr_14_3 : OUT std_logic ;
         d_arr_14_2 : OUT std_logic ;
         d_arr_14_1 : OUT std_logic ;
         d_arr_14_0 : OUT std_logic ;
         d_arr_15_31 : OUT std_logic ;
         d_arr_15_30 : OUT std_logic ;
         d_arr_15_29 : OUT std_logic ;
         d_arr_15_28 : OUT std_logic ;
         d_arr_15_27 : OUT std_logic ;
         d_arr_15_26 : OUT std_logic ;
         d_arr_15_25 : OUT std_logic ;
         d_arr_15_24 : OUT std_logic ;
         d_arr_15_23 : OUT std_logic ;
         d_arr_15_22 : OUT std_logic ;
         d_arr_15_21 : OUT std_logic ;
         d_arr_15_20 : OUT std_logic ;
         d_arr_15_19 : OUT std_logic ;
         d_arr_15_18 : OUT std_logic ;
         d_arr_15_17 : OUT std_logic ;
         d_arr_15_16 : OUT std_logic ;
         d_arr_15_15 : OUT std_logic ;
         d_arr_15_14 : OUT std_logic ;
         d_arr_15_13 : OUT std_logic ;
         d_arr_15_12 : OUT std_logic ;
         d_arr_15_11 : OUT std_logic ;
         d_arr_15_10 : OUT std_logic ;
         d_arr_15_9 : OUT std_logic ;
         d_arr_15_8 : OUT std_logic ;
         d_arr_15_7 : OUT std_logic ;
         d_arr_15_6 : OUT std_logic ;
         d_arr_15_5 : OUT std_logic ;
         d_arr_15_4 : OUT std_logic ;
         d_arr_15_3 : OUT std_logic ;
         d_arr_15_2 : OUT std_logic ;
         d_arr_15_1 : OUT std_logic ;
         d_arr_15_0 : OUT std_logic ;
         d_arr_16_31 : OUT std_logic ;
         d_arr_16_30 : OUT std_logic ;
         d_arr_16_29 : OUT std_logic ;
         d_arr_16_28 : OUT std_logic ;
         d_arr_16_27 : OUT std_logic ;
         d_arr_16_26 : OUT std_logic ;
         d_arr_16_25 : OUT std_logic ;
         d_arr_16_24 : OUT std_logic ;
         d_arr_16_23 : OUT std_logic ;
         d_arr_16_22 : OUT std_logic ;
         d_arr_16_21 : OUT std_logic ;
         d_arr_16_20 : OUT std_logic ;
         d_arr_16_19 : OUT std_logic ;
         d_arr_16_18 : OUT std_logic ;
         d_arr_16_17 : OUT std_logic ;
         d_arr_16_16 : OUT std_logic ;
         d_arr_16_15 : OUT std_logic ;
         d_arr_16_14 : OUT std_logic ;
         d_arr_16_13 : OUT std_logic ;
         d_arr_16_12 : OUT std_logic ;
         d_arr_16_11 : OUT std_logic ;
         d_arr_16_10 : OUT std_logic ;
         d_arr_16_9 : OUT std_logic ;
         d_arr_16_8 : OUT std_logic ;
         d_arr_16_7 : OUT std_logic ;
         d_arr_16_6 : OUT std_logic ;
         d_arr_16_5 : OUT std_logic ;
         d_arr_16_4 : OUT std_logic ;
         d_arr_16_3 : OUT std_logic ;
         d_arr_16_2 : OUT std_logic ;
         d_arr_16_1 : OUT std_logic ;
         d_arr_16_0 : OUT std_logic ;
         d_arr_17_31 : OUT std_logic ;
         d_arr_17_30 : OUT std_logic ;
         d_arr_17_29 : OUT std_logic ;
         d_arr_17_28 : OUT std_logic ;
         d_arr_17_27 : OUT std_logic ;
         d_arr_17_26 : OUT std_logic ;
         d_arr_17_25 : OUT std_logic ;
         d_arr_17_24 : OUT std_logic ;
         d_arr_17_23 : OUT std_logic ;
         d_arr_17_22 : OUT std_logic ;
         d_arr_17_21 : OUT std_logic ;
         d_arr_17_20 : OUT std_logic ;
         d_arr_17_19 : OUT std_logic ;
         d_arr_17_18 : OUT std_logic ;
         d_arr_17_17 : OUT std_logic ;
         d_arr_17_16 : OUT std_logic ;
         d_arr_17_15 : OUT std_logic ;
         d_arr_17_14 : OUT std_logic ;
         d_arr_17_13 : OUT std_logic ;
         d_arr_17_12 : OUT std_logic ;
         d_arr_17_11 : OUT std_logic ;
         d_arr_17_10 : OUT std_logic ;
         d_arr_17_9 : OUT std_logic ;
         d_arr_17_8 : OUT std_logic ;
         d_arr_17_7 : OUT std_logic ;
         d_arr_17_6 : OUT std_logic ;
         d_arr_17_5 : OUT std_logic ;
         d_arr_17_4 : OUT std_logic ;
         d_arr_17_3 : OUT std_logic ;
         d_arr_17_2 : OUT std_logic ;
         d_arr_17_1 : OUT std_logic ;
         d_arr_17_0 : OUT std_logic ;
         d_arr_18_31 : OUT std_logic ;
         d_arr_18_30 : OUT std_logic ;
         d_arr_18_29 : OUT std_logic ;
         d_arr_18_28 : OUT std_logic ;
         d_arr_18_27 : OUT std_logic ;
         d_arr_18_26 : OUT std_logic ;
         d_arr_18_25 : OUT std_logic ;
         d_arr_18_24 : OUT std_logic ;
         d_arr_18_23 : OUT std_logic ;
         d_arr_18_22 : OUT std_logic ;
         d_arr_18_21 : OUT std_logic ;
         d_arr_18_20 : OUT std_logic ;
         d_arr_18_19 : OUT std_logic ;
         d_arr_18_18 : OUT std_logic ;
         d_arr_18_17 : OUT std_logic ;
         d_arr_18_16 : OUT std_logic ;
         d_arr_18_15 : OUT std_logic ;
         d_arr_18_14 : OUT std_logic ;
         d_arr_18_13 : OUT std_logic ;
         d_arr_18_12 : OUT std_logic ;
         d_arr_18_11 : OUT std_logic ;
         d_arr_18_10 : OUT std_logic ;
         d_arr_18_9 : OUT std_logic ;
         d_arr_18_8 : OUT std_logic ;
         d_arr_18_7 : OUT std_logic ;
         d_arr_18_6 : OUT std_logic ;
         d_arr_18_5 : OUT std_logic ;
         d_arr_18_4 : OUT std_logic ;
         d_arr_18_3 : OUT std_logic ;
         d_arr_18_2 : OUT std_logic ;
         d_arr_18_1 : OUT std_logic ;
         d_arr_18_0 : OUT std_logic ;
         d_arr_19_31 : OUT std_logic ;
         d_arr_19_30 : OUT std_logic ;
         d_arr_19_29 : OUT std_logic ;
         d_arr_19_28 : OUT std_logic ;
         d_arr_19_27 : OUT std_logic ;
         d_arr_19_26 : OUT std_logic ;
         d_arr_19_25 : OUT std_logic ;
         d_arr_19_24 : OUT std_logic ;
         d_arr_19_23 : OUT std_logic ;
         d_arr_19_22 : OUT std_logic ;
         d_arr_19_21 : OUT std_logic ;
         d_arr_19_20 : OUT std_logic ;
         d_arr_19_19 : OUT std_logic ;
         d_arr_19_18 : OUT std_logic ;
         d_arr_19_17 : OUT std_logic ;
         d_arr_19_16 : OUT std_logic ;
         d_arr_19_15 : OUT std_logic ;
         d_arr_19_14 : OUT std_logic ;
         d_arr_19_13 : OUT std_logic ;
         d_arr_19_12 : OUT std_logic ;
         d_arr_19_11 : OUT std_logic ;
         d_arr_19_10 : OUT std_logic ;
         d_arr_19_9 : OUT std_logic ;
         d_arr_19_8 : OUT std_logic ;
         d_arr_19_7 : OUT std_logic ;
         d_arr_19_6 : OUT std_logic ;
         d_arr_19_5 : OUT std_logic ;
         d_arr_19_4 : OUT std_logic ;
         d_arr_19_3 : OUT std_logic ;
         d_arr_19_2 : OUT std_logic ;
         d_arr_19_1 : OUT std_logic ;
         d_arr_19_0 : OUT std_logic ;
         d_arr_20_31 : OUT std_logic ;
         d_arr_20_30 : OUT std_logic ;
         d_arr_20_29 : OUT std_logic ;
         d_arr_20_28 : OUT std_logic ;
         d_arr_20_27 : OUT std_logic ;
         d_arr_20_26 : OUT std_logic ;
         d_arr_20_25 : OUT std_logic ;
         d_arr_20_24 : OUT std_logic ;
         d_arr_20_23 : OUT std_logic ;
         d_arr_20_22 : OUT std_logic ;
         d_arr_20_21 : OUT std_logic ;
         d_arr_20_20 : OUT std_logic ;
         d_arr_20_19 : OUT std_logic ;
         d_arr_20_18 : OUT std_logic ;
         d_arr_20_17 : OUT std_logic ;
         d_arr_20_16 : OUT std_logic ;
         d_arr_20_15 : OUT std_logic ;
         d_arr_20_14 : OUT std_logic ;
         d_arr_20_13 : OUT std_logic ;
         d_arr_20_12 : OUT std_logic ;
         d_arr_20_11 : OUT std_logic ;
         d_arr_20_10 : OUT std_logic ;
         d_arr_20_9 : OUT std_logic ;
         d_arr_20_8 : OUT std_logic ;
         d_arr_20_7 : OUT std_logic ;
         d_arr_20_6 : OUT std_logic ;
         d_arr_20_5 : OUT std_logic ;
         d_arr_20_4 : OUT std_logic ;
         d_arr_20_3 : OUT std_logic ;
         d_arr_20_2 : OUT std_logic ;
         d_arr_20_1 : OUT std_logic ;
         d_arr_20_0 : OUT std_logic ;
         d_arr_21_31 : OUT std_logic ;
         d_arr_21_30 : OUT std_logic ;
         d_arr_21_29 : OUT std_logic ;
         d_arr_21_28 : OUT std_logic ;
         d_arr_21_27 : OUT std_logic ;
         d_arr_21_26 : OUT std_logic ;
         d_arr_21_25 : OUT std_logic ;
         d_arr_21_24 : OUT std_logic ;
         d_arr_21_23 : OUT std_logic ;
         d_arr_21_22 : OUT std_logic ;
         d_arr_21_21 : OUT std_logic ;
         d_arr_21_20 : OUT std_logic ;
         d_arr_21_19 : OUT std_logic ;
         d_arr_21_18 : OUT std_logic ;
         d_arr_21_17 : OUT std_logic ;
         d_arr_21_16 : OUT std_logic ;
         d_arr_21_15 : OUT std_logic ;
         d_arr_21_14 : OUT std_logic ;
         d_arr_21_13 : OUT std_logic ;
         d_arr_21_12 : OUT std_logic ;
         d_arr_21_11 : OUT std_logic ;
         d_arr_21_10 : OUT std_logic ;
         d_arr_21_9 : OUT std_logic ;
         d_arr_21_8 : OUT std_logic ;
         d_arr_21_7 : OUT std_logic ;
         d_arr_21_6 : OUT std_logic ;
         d_arr_21_5 : OUT std_logic ;
         d_arr_21_4 : OUT std_logic ;
         d_arr_21_3 : OUT std_logic ;
         d_arr_21_2 : OUT std_logic ;
         d_arr_21_1 : OUT std_logic ;
         d_arr_21_0 : OUT std_logic ;
         d_arr_22_31 : OUT std_logic ;
         d_arr_22_30 : OUT std_logic ;
         d_arr_22_29 : OUT std_logic ;
         d_arr_22_28 : OUT std_logic ;
         d_arr_22_27 : OUT std_logic ;
         d_arr_22_26 : OUT std_logic ;
         d_arr_22_25 : OUT std_logic ;
         d_arr_22_24 : OUT std_logic ;
         d_arr_22_23 : OUT std_logic ;
         d_arr_22_22 : OUT std_logic ;
         d_arr_22_21 : OUT std_logic ;
         d_arr_22_20 : OUT std_logic ;
         d_arr_22_19 : OUT std_logic ;
         d_arr_22_18 : OUT std_logic ;
         d_arr_22_17 : OUT std_logic ;
         d_arr_22_16 : OUT std_logic ;
         d_arr_22_15 : OUT std_logic ;
         d_arr_22_14 : OUT std_logic ;
         d_arr_22_13 : OUT std_logic ;
         d_arr_22_12 : OUT std_logic ;
         d_arr_22_11 : OUT std_logic ;
         d_arr_22_10 : OUT std_logic ;
         d_arr_22_9 : OUT std_logic ;
         d_arr_22_8 : OUT std_logic ;
         d_arr_22_7 : OUT std_logic ;
         d_arr_22_6 : OUT std_logic ;
         d_arr_22_5 : OUT std_logic ;
         d_arr_22_4 : OUT std_logic ;
         d_arr_22_3 : OUT std_logic ;
         d_arr_22_2 : OUT std_logic ;
         d_arr_22_1 : OUT std_logic ;
         d_arr_22_0 : OUT std_logic ;
         d_arr_23_31 : OUT std_logic ;
         d_arr_23_30 : OUT std_logic ;
         d_arr_23_29 : OUT std_logic ;
         d_arr_23_28 : OUT std_logic ;
         d_arr_23_27 : OUT std_logic ;
         d_arr_23_26 : OUT std_logic ;
         d_arr_23_25 : OUT std_logic ;
         d_arr_23_24 : OUT std_logic ;
         d_arr_23_23 : OUT std_logic ;
         d_arr_23_22 : OUT std_logic ;
         d_arr_23_21 : OUT std_logic ;
         d_arr_23_20 : OUT std_logic ;
         d_arr_23_19 : OUT std_logic ;
         d_arr_23_18 : OUT std_logic ;
         d_arr_23_17 : OUT std_logic ;
         d_arr_23_16 : OUT std_logic ;
         d_arr_23_15 : OUT std_logic ;
         d_arr_23_14 : OUT std_logic ;
         d_arr_23_13 : OUT std_logic ;
         d_arr_23_12 : OUT std_logic ;
         d_arr_23_11 : OUT std_logic ;
         d_arr_23_10 : OUT std_logic ;
         d_arr_23_9 : OUT std_logic ;
         d_arr_23_8 : OUT std_logic ;
         d_arr_23_7 : OUT std_logic ;
         d_arr_23_6 : OUT std_logic ;
         d_arr_23_5 : OUT std_logic ;
         d_arr_23_4 : OUT std_logic ;
         d_arr_23_3 : OUT std_logic ;
         d_arr_23_2 : OUT std_logic ;
         d_arr_23_1 : OUT std_logic ;
         d_arr_23_0 : OUT std_logic ;
         d_arr_24_31 : OUT std_logic ;
         d_arr_24_30 : OUT std_logic ;
         d_arr_24_29 : OUT std_logic ;
         d_arr_24_28 : OUT std_logic ;
         d_arr_24_27 : OUT std_logic ;
         d_arr_24_26 : OUT std_logic ;
         d_arr_24_25 : OUT std_logic ;
         d_arr_24_24 : OUT std_logic ;
         d_arr_24_23 : OUT std_logic ;
         d_arr_24_22 : OUT std_logic ;
         d_arr_24_21 : OUT std_logic ;
         d_arr_24_20 : OUT std_logic ;
         d_arr_24_19 : OUT std_logic ;
         d_arr_24_18 : OUT std_logic ;
         d_arr_24_17 : OUT std_logic ;
         d_arr_24_16 : OUT std_logic ;
         d_arr_24_15 : OUT std_logic ;
         d_arr_24_14 : OUT std_logic ;
         d_arr_24_13 : OUT std_logic ;
         d_arr_24_12 : OUT std_logic ;
         d_arr_24_11 : OUT std_logic ;
         d_arr_24_10 : OUT std_logic ;
         d_arr_24_9 : OUT std_logic ;
         d_arr_24_8 : OUT std_logic ;
         d_arr_24_7 : OUT std_logic ;
         d_arr_24_6 : OUT std_logic ;
         d_arr_24_5 : OUT std_logic ;
         d_arr_24_4 : OUT std_logic ;
         d_arr_24_3 : OUT std_logic ;
         d_arr_24_2 : OUT std_logic ;
         d_arr_24_1 : OUT std_logic ;
         d_arr_24_0 : OUT std_logic ;
         q_arr_0_31 : IN std_logic ;
         q_arr_0_30 : IN std_logic ;
         q_arr_0_29 : IN std_logic ;
         q_arr_0_28 : IN std_logic ;
         q_arr_0_27 : IN std_logic ;
         q_arr_0_26 : IN std_logic ;
         q_arr_0_25 : IN std_logic ;
         q_arr_0_24 : IN std_logic ;
         q_arr_0_23 : IN std_logic ;
         q_arr_0_22 : IN std_logic ;
         q_arr_0_21 : IN std_logic ;
         q_arr_0_20 : IN std_logic ;
         q_arr_0_19 : IN std_logic ;
         q_arr_0_18 : IN std_logic ;
         q_arr_0_17 : IN std_logic ;
         q_arr_0_16 : IN std_logic ;
         q_arr_0_15 : IN std_logic ;
         q_arr_0_14 : IN std_logic ;
         q_arr_0_13 : IN std_logic ;
         q_arr_0_12 : IN std_logic ;
         q_arr_0_11 : IN std_logic ;
         q_arr_0_10 : IN std_logic ;
         q_arr_0_9 : IN std_logic ;
         q_arr_0_8 : IN std_logic ;
         q_arr_0_7 : IN std_logic ;
         q_arr_0_6 : IN std_logic ;
         q_arr_0_5 : IN std_logic ;
         q_arr_0_4 : IN std_logic ;
         q_arr_0_3 : IN std_logic ;
         q_arr_0_2 : IN std_logic ;
         q_arr_0_1 : IN std_logic ;
         q_arr_0_0 : IN std_logic ;
         q_arr_1_31 : IN std_logic ;
         q_arr_1_30 : IN std_logic ;
         q_arr_1_29 : IN std_logic ;
         q_arr_1_28 : IN std_logic ;
         q_arr_1_27 : IN std_logic ;
         q_arr_1_26 : IN std_logic ;
         q_arr_1_25 : IN std_logic ;
         q_arr_1_24 : IN std_logic ;
         q_arr_1_23 : IN std_logic ;
         q_arr_1_22 : IN std_logic ;
         q_arr_1_21 : IN std_logic ;
         q_arr_1_20 : IN std_logic ;
         q_arr_1_19 : IN std_logic ;
         q_arr_1_18 : IN std_logic ;
         q_arr_1_17 : IN std_logic ;
         q_arr_1_16 : IN std_logic ;
         q_arr_1_15 : IN std_logic ;
         q_arr_1_14 : IN std_logic ;
         q_arr_1_13 : IN std_logic ;
         q_arr_1_12 : IN std_logic ;
         q_arr_1_11 : IN std_logic ;
         q_arr_1_10 : IN std_logic ;
         q_arr_1_9 : IN std_logic ;
         q_arr_1_8 : IN std_logic ;
         q_arr_1_7 : IN std_logic ;
         q_arr_1_6 : IN std_logic ;
         q_arr_1_5 : IN std_logic ;
         q_arr_1_4 : IN std_logic ;
         q_arr_1_3 : IN std_logic ;
         q_arr_1_2 : IN std_logic ;
         q_arr_1_1 : IN std_logic ;
         q_arr_1_0 : IN std_logic ;
         q_arr_2_31 : IN std_logic ;
         q_arr_2_30 : IN std_logic ;
         q_arr_2_29 : IN std_logic ;
         q_arr_2_28 : IN std_logic ;
         q_arr_2_27 : IN std_logic ;
         q_arr_2_26 : IN std_logic ;
         q_arr_2_25 : IN std_logic ;
         q_arr_2_24 : IN std_logic ;
         q_arr_2_23 : IN std_logic ;
         q_arr_2_22 : IN std_logic ;
         q_arr_2_21 : IN std_logic ;
         q_arr_2_20 : IN std_logic ;
         q_arr_2_19 : IN std_logic ;
         q_arr_2_18 : IN std_logic ;
         q_arr_2_17 : IN std_logic ;
         q_arr_2_16 : IN std_logic ;
         q_arr_2_15 : IN std_logic ;
         q_arr_2_14 : IN std_logic ;
         q_arr_2_13 : IN std_logic ;
         q_arr_2_12 : IN std_logic ;
         q_arr_2_11 : IN std_logic ;
         q_arr_2_10 : IN std_logic ;
         q_arr_2_9 : IN std_logic ;
         q_arr_2_8 : IN std_logic ;
         q_arr_2_7 : IN std_logic ;
         q_arr_2_6 : IN std_logic ;
         q_arr_2_5 : IN std_logic ;
         q_arr_2_4 : IN std_logic ;
         q_arr_2_3 : IN std_logic ;
         q_arr_2_2 : IN std_logic ;
         q_arr_2_1 : IN std_logic ;
         q_arr_2_0 : IN std_logic ;
         q_arr_3_31 : IN std_logic ;
         q_arr_3_30 : IN std_logic ;
         q_arr_3_29 : IN std_logic ;
         q_arr_3_28 : IN std_logic ;
         q_arr_3_27 : IN std_logic ;
         q_arr_3_26 : IN std_logic ;
         q_arr_3_25 : IN std_logic ;
         q_arr_3_24 : IN std_logic ;
         q_arr_3_23 : IN std_logic ;
         q_arr_3_22 : IN std_logic ;
         q_arr_3_21 : IN std_logic ;
         q_arr_3_20 : IN std_logic ;
         q_arr_3_19 : IN std_logic ;
         q_arr_3_18 : IN std_logic ;
         q_arr_3_17 : IN std_logic ;
         q_arr_3_16 : IN std_logic ;
         q_arr_3_15 : IN std_logic ;
         q_arr_3_14 : IN std_logic ;
         q_arr_3_13 : IN std_logic ;
         q_arr_3_12 : IN std_logic ;
         q_arr_3_11 : IN std_logic ;
         q_arr_3_10 : IN std_logic ;
         q_arr_3_9 : IN std_logic ;
         q_arr_3_8 : IN std_logic ;
         q_arr_3_7 : IN std_logic ;
         q_arr_3_6 : IN std_logic ;
         q_arr_3_5 : IN std_logic ;
         q_arr_3_4 : IN std_logic ;
         q_arr_3_3 : IN std_logic ;
         q_arr_3_2 : IN std_logic ;
         q_arr_3_1 : IN std_logic ;
         q_arr_3_0 : IN std_logic ;
         q_arr_4_31 : IN std_logic ;
         q_arr_4_30 : IN std_logic ;
         q_arr_4_29 : IN std_logic ;
         q_arr_4_28 : IN std_logic ;
         q_arr_4_27 : IN std_logic ;
         q_arr_4_26 : IN std_logic ;
         q_arr_4_25 : IN std_logic ;
         q_arr_4_24 : IN std_logic ;
         q_arr_4_23 : IN std_logic ;
         q_arr_4_22 : IN std_logic ;
         q_arr_4_21 : IN std_logic ;
         q_arr_4_20 : IN std_logic ;
         q_arr_4_19 : IN std_logic ;
         q_arr_4_18 : IN std_logic ;
         q_arr_4_17 : IN std_logic ;
         q_arr_4_16 : IN std_logic ;
         q_arr_4_15 : IN std_logic ;
         q_arr_4_14 : IN std_logic ;
         q_arr_4_13 : IN std_logic ;
         q_arr_4_12 : IN std_logic ;
         q_arr_4_11 : IN std_logic ;
         q_arr_4_10 : IN std_logic ;
         q_arr_4_9 : IN std_logic ;
         q_arr_4_8 : IN std_logic ;
         q_arr_4_7 : IN std_logic ;
         q_arr_4_6 : IN std_logic ;
         q_arr_4_5 : IN std_logic ;
         q_arr_4_4 : IN std_logic ;
         q_arr_4_3 : IN std_logic ;
         q_arr_4_2 : IN std_logic ;
         q_arr_4_1 : IN std_logic ;
         q_arr_4_0 : IN std_logic ;
         q_arr_5_31 : IN std_logic ;
         q_arr_5_30 : IN std_logic ;
         q_arr_5_29 : IN std_logic ;
         q_arr_5_28 : IN std_logic ;
         q_arr_5_27 : IN std_logic ;
         q_arr_5_26 : IN std_logic ;
         q_arr_5_25 : IN std_logic ;
         q_arr_5_24 : IN std_logic ;
         q_arr_5_23 : IN std_logic ;
         q_arr_5_22 : IN std_logic ;
         q_arr_5_21 : IN std_logic ;
         q_arr_5_20 : IN std_logic ;
         q_arr_5_19 : IN std_logic ;
         q_arr_5_18 : IN std_logic ;
         q_arr_5_17 : IN std_logic ;
         q_arr_5_16 : IN std_logic ;
         q_arr_5_15 : IN std_logic ;
         q_arr_5_14 : IN std_logic ;
         q_arr_5_13 : IN std_logic ;
         q_arr_5_12 : IN std_logic ;
         q_arr_5_11 : IN std_logic ;
         q_arr_5_10 : IN std_logic ;
         q_arr_5_9 : IN std_logic ;
         q_arr_5_8 : IN std_logic ;
         q_arr_5_7 : IN std_logic ;
         q_arr_5_6 : IN std_logic ;
         q_arr_5_5 : IN std_logic ;
         q_arr_5_4 : IN std_logic ;
         q_arr_5_3 : IN std_logic ;
         q_arr_5_2 : IN std_logic ;
         q_arr_5_1 : IN std_logic ;
         q_arr_5_0 : IN std_logic ;
         q_arr_6_31 : IN std_logic ;
         q_arr_6_30 : IN std_logic ;
         q_arr_6_29 : IN std_logic ;
         q_arr_6_28 : IN std_logic ;
         q_arr_6_27 : IN std_logic ;
         q_arr_6_26 : IN std_logic ;
         q_arr_6_25 : IN std_logic ;
         q_arr_6_24 : IN std_logic ;
         q_arr_6_23 : IN std_logic ;
         q_arr_6_22 : IN std_logic ;
         q_arr_6_21 : IN std_logic ;
         q_arr_6_20 : IN std_logic ;
         q_arr_6_19 : IN std_logic ;
         q_arr_6_18 : IN std_logic ;
         q_arr_6_17 : IN std_logic ;
         q_arr_6_16 : IN std_logic ;
         q_arr_6_15 : IN std_logic ;
         q_arr_6_14 : IN std_logic ;
         q_arr_6_13 : IN std_logic ;
         q_arr_6_12 : IN std_logic ;
         q_arr_6_11 : IN std_logic ;
         q_arr_6_10 : IN std_logic ;
         q_arr_6_9 : IN std_logic ;
         q_arr_6_8 : IN std_logic ;
         q_arr_6_7 : IN std_logic ;
         q_arr_6_6 : IN std_logic ;
         q_arr_6_5 : IN std_logic ;
         q_arr_6_4 : IN std_logic ;
         q_arr_6_3 : IN std_logic ;
         q_arr_6_2 : IN std_logic ;
         q_arr_6_1 : IN std_logic ;
         q_arr_6_0 : IN std_logic ;
         q_arr_7_31 : IN std_logic ;
         q_arr_7_30 : IN std_logic ;
         q_arr_7_29 : IN std_logic ;
         q_arr_7_28 : IN std_logic ;
         q_arr_7_27 : IN std_logic ;
         q_arr_7_26 : IN std_logic ;
         q_arr_7_25 : IN std_logic ;
         q_arr_7_24 : IN std_logic ;
         q_arr_7_23 : IN std_logic ;
         q_arr_7_22 : IN std_logic ;
         q_arr_7_21 : IN std_logic ;
         q_arr_7_20 : IN std_logic ;
         q_arr_7_19 : IN std_logic ;
         q_arr_7_18 : IN std_logic ;
         q_arr_7_17 : IN std_logic ;
         q_arr_7_16 : IN std_logic ;
         q_arr_7_15 : IN std_logic ;
         q_arr_7_14 : IN std_logic ;
         q_arr_7_13 : IN std_logic ;
         q_arr_7_12 : IN std_logic ;
         q_arr_7_11 : IN std_logic ;
         q_arr_7_10 : IN std_logic ;
         q_arr_7_9 : IN std_logic ;
         q_arr_7_8 : IN std_logic ;
         q_arr_7_7 : IN std_logic ;
         q_arr_7_6 : IN std_logic ;
         q_arr_7_5 : IN std_logic ;
         q_arr_7_4 : IN std_logic ;
         q_arr_7_3 : IN std_logic ;
         q_arr_7_2 : IN std_logic ;
         q_arr_7_1 : IN std_logic ;
         q_arr_7_0 : IN std_logic ;
         q_arr_8_31 : IN std_logic ;
         q_arr_8_30 : IN std_logic ;
         q_arr_8_29 : IN std_logic ;
         q_arr_8_28 : IN std_logic ;
         q_arr_8_27 : IN std_logic ;
         q_arr_8_26 : IN std_logic ;
         q_arr_8_25 : IN std_logic ;
         q_arr_8_24 : IN std_logic ;
         q_arr_8_23 : IN std_logic ;
         q_arr_8_22 : IN std_logic ;
         q_arr_8_21 : IN std_logic ;
         q_arr_8_20 : IN std_logic ;
         q_arr_8_19 : IN std_logic ;
         q_arr_8_18 : IN std_logic ;
         q_arr_8_17 : IN std_logic ;
         q_arr_8_16 : IN std_logic ;
         q_arr_8_15 : IN std_logic ;
         q_arr_8_14 : IN std_logic ;
         q_arr_8_13 : IN std_logic ;
         q_arr_8_12 : IN std_logic ;
         q_arr_8_11 : IN std_logic ;
         q_arr_8_10 : IN std_logic ;
         q_arr_8_9 : IN std_logic ;
         q_arr_8_8 : IN std_logic ;
         q_arr_8_7 : IN std_logic ;
         q_arr_8_6 : IN std_logic ;
         q_arr_8_5 : IN std_logic ;
         q_arr_8_4 : IN std_logic ;
         q_arr_8_3 : IN std_logic ;
         q_arr_8_2 : IN std_logic ;
         q_arr_8_1 : IN std_logic ;
         q_arr_8_0 : IN std_logic ;
         q_arr_9_31 : IN std_logic ;
         q_arr_9_30 : IN std_logic ;
         q_arr_9_29 : IN std_logic ;
         q_arr_9_28 : IN std_logic ;
         q_arr_9_27 : IN std_logic ;
         q_arr_9_26 : IN std_logic ;
         q_arr_9_25 : IN std_logic ;
         q_arr_9_24 : IN std_logic ;
         q_arr_9_23 : IN std_logic ;
         q_arr_9_22 : IN std_logic ;
         q_arr_9_21 : IN std_logic ;
         q_arr_9_20 : IN std_logic ;
         q_arr_9_19 : IN std_logic ;
         q_arr_9_18 : IN std_logic ;
         q_arr_9_17 : IN std_logic ;
         q_arr_9_16 : IN std_logic ;
         q_arr_9_15 : IN std_logic ;
         q_arr_9_14 : IN std_logic ;
         q_arr_9_13 : IN std_logic ;
         q_arr_9_12 : IN std_logic ;
         q_arr_9_11 : IN std_logic ;
         q_arr_9_10 : IN std_logic ;
         q_arr_9_9 : IN std_logic ;
         q_arr_9_8 : IN std_logic ;
         q_arr_9_7 : IN std_logic ;
         q_arr_9_6 : IN std_logic ;
         q_arr_9_5 : IN std_logic ;
         q_arr_9_4 : IN std_logic ;
         q_arr_9_3 : IN std_logic ;
         q_arr_9_2 : IN std_logic ;
         q_arr_9_1 : IN std_logic ;
         q_arr_9_0 : IN std_logic ;
         q_arr_10_31 : IN std_logic ;
         q_arr_10_30 : IN std_logic ;
         q_arr_10_29 : IN std_logic ;
         q_arr_10_28 : IN std_logic ;
         q_arr_10_27 : IN std_logic ;
         q_arr_10_26 : IN std_logic ;
         q_arr_10_25 : IN std_logic ;
         q_arr_10_24 : IN std_logic ;
         q_arr_10_23 : IN std_logic ;
         q_arr_10_22 : IN std_logic ;
         q_arr_10_21 : IN std_logic ;
         q_arr_10_20 : IN std_logic ;
         q_arr_10_19 : IN std_logic ;
         q_arr_10_18 : IN std_logic ;
         q_arr_10_17 : IN std_logic ;
         q_arr_10_16 : IN std_logic ;
         q_arr_10_15 : IN std_logic ;
         q_arr_10_14 : IN std_logic ;
         q_arr_10_13 : IN std_logic ;
         q_arr_10_12 : IN std_logic ;
         q_arr_10_11 : IN std_logic ;
         q_arr_10_10 : IN std_logic ;
         q_arr_10_9 : IN std_logic ;
         q_arr_10_8 : IN std_logic ;
         q_arr_10_7 : IN std_logic ;
         q_arr_10_6 : IN std_logic ;
         q_arr_10_5 : IN std_logic ;
         q_arr_10_4 : IN std_logic ;
         q_arr_10_3 : IN std_logic ;
         q_arr_10_2 : IN std_logic ;
         q_arr_10_1 : IN std_logic ;
         q_arr_10_0 : IN std_logic ;
         q_arr_11_31 : IN std_logic ;
         q_arr_11_30 : IN std_logic ;
         q_arr_11_29 : IN std_logic ;
         q_arr_11_28 : IN std_logic ;
         q_arr_11_27 : IN std_logic ;
         q_arr_11_26 : IN std_logic ;
         q_arr_11_25 : IN std_logic ;
         q_arr_11_24 : IN std_logic ;
         q_arr_11_23 : IN std_logic ;
         q_arr_11_22 : IN std_logic ;
         q_arr_11_21 : IN std_logic ;
         q_arr_11_20 : IN std_logic ;
         q_arr_11_19 : IN std_logic ;
         q_arr_11_18 : IN std_logic ;
         q_arr_11_17 : IN std_logic ;
         q_arr_11_16 : IN std_logic ;
         q_arr_11_15 : IN std_logic ;
         q_arr_11_14 : IN std_logic ;
         q_arr_11_13 : IN std_logic ;
         q_arr_11_12 : IN std_logic ;
         q_arr_11_11 : IN std_logic ;
         q_arr_11_10 : IN std_logic ;
         q_arr_11_9 : IN std_logic ;
         q_arr_11_8 : IN std_logic ;
         q_arr_11_7 : IN std_logic ;
         q_arr_11_6 : IN std_logic ;
         q_arr_11_5 : IN std_logic ;
         q_arr_11_4 : IN std_logic ;
         q_arr_11_3 : IN std_logic ;
         q_arr_11_2 : IN std_logic ;
         q_arr_11_1 : IN std_logic ;
         q_arr_11_0 : IN std_logic ;
         q_arr_12_31 : IN std_logic ;
         q_arr_12_30 : IN std_logic ;
         q_arr_12_29 : IN std_logic ;
         q_arr_12_28 : IN std_logic ;
         q_arr_12_27 : IN std_logic ;
         q_arr_12_26 : IN std_logic ;
         q_arr_12_25 : IN std_logic ;
         q_arr_12_24 : IN std_logic ;
         q_arr_12_23 : IN std_logic ;
         q_arr_12_22 : IN std_logic ;
         q_arr_12_21 : IN std_logic ;
         q_arr_12_20 : IN std_logic ;
         q_arr_12_19 : IN std_logic ;
         q_arr_12_18 : IN std_logic ;
         q_arr_12_17 : IN std_logic ;
         q_arr_12_16 : IN std_logic ;
         q_arr_12_15 : IN std_logic ;
         q_arr_12_14 : IN std_logic ;
         q_arr_12_13 : IN std_logic ;
         q_arr_12_12 : IN std_logic ;
         q_arr_12_11 : IN std_logic ;
         q_arr_12_10 : IN std_logic ;
         q_arr_12_9 : IN std_logic ;
         q_arr_12_8 : IN std_logic ;
         q_arr_12_7 : IN std_logic ;
         q_arr_12_6 : IN std_logic ;
         q_arr_12_5 : IN std_logic ;
         q_arr_12_4 : IN std_logic ;
         q_arr_12_3 : IN std_logic ;
         q_arr_12_2 : IN std_logic ;
         q_arr_12_1 : IN std_logic ;
         q_arr_12_0 : IN std_logic ;
         q_arr_13_31 : IN std_logic ;
         q_arr_13_30 : IN std_logic ;
         q_arr_13_29 : IN std_logic ;
         q_arr_13_28 : IN std_logic ;
         q_arr_13_27 : IN std_logic ;
         q_arr_13_26 : IN std_logic ;
         q_arr_13_25 : IN std_logic ;
         q_arr_13_24 : IN std_logic ;
         q_arr_13_23 : IN std_logic ;
         q_arr_13_22 : IN std_logic ;
         q_arr_13_21 : IN std_logic ;
         q_arr_13_20 : IN std_logic ;
         q_arr_13_19 : IN std_logic ;
         q_arr_13_18 : IN std_logic ;
         q_arr_13_17 : IN std_logic ;
         q_arr_13_16 : IN std_logic ;
         q_arr_13_15 : IN std_logic ;
         q_arr_13_14 : IN std_logic ;
         q_arr_13_13 : IN std_logic ;
         q_arr_13_12 : IN std_logic ;
         q_arr_13_11 : IN std_logic ;
         q_arr_13_10 : IN std_logic ;
         q_arr_13_9 : IN std_logic ;
         q_arr_13_8 : IN std_logic ;
         q_arr_13_7 : IN std_logic ;
         q_arr_13_6 : IN std_logic ;
         q_arr_13_5 : IN std_logic ;
         q_arr_13_4 : IN std_logic ;
         q_arr_13_3 : IN std_logic ;
         q_arr_13_2 : IN std_logic ;
         q_arr_13_1 : IN std_logic ;
         q_arr_13_0 : IN std_logic ;
         q_arr_14_31 : IN std_logic ;
         q_arr_14_30 : IN std_logic ;
         q_arr_14_29 : IN std_logic ;
         q_arr_14_28 : IN std_logic ;
         q_arr_14_27 : IN std_logic ;
         q_arr_14_26 : IN std_logic ;
         q_arr_14_25 : IN std_logic ;
         q_arr_14_24 : IN std_logic ;
         q_arr_14_23 : IN std_logic ;
         q_arr_14_22 : IN std_logic ;
         q_arr_14_21 : IN std_logic ;
         q_arr_14_20 : IN std_logic ;
         q_arr_14_19 : IN std_logic ;
         q_arr_14_18 : IN std_logic ;
         q_arr_14_17 : IN std_logic ;
         q_arr_14_16 : IN std_logic ;
         q_arr_14_15 : IN std_logic ;
         q_arr_14_14 : IN std_logic ;
         q_arr_14_13 : IN std_logic ;
         q_arr_14_12 : IN std_logic ;
         q_arr_14_11 : IN std_logic ;
         q_arr_14_10 : IN std_logic ;
         q_arr_14_9 : IN std_logic ;
         q_arr_14_8 : IN std_logic ;
         q_arr_14_7 : IN std_logic ;
         q_arr_14_6 : IN std_logic ;
         q_arr_14_5 : IN std_logic ;
         q_arr_14_4 : IN std_logic ;
         q_arr_14_3 : IN std_logic ;
         q_arr_14_2 : IN std_logic ;
         q_arr_14_1 : IN std_logic ;
         q_arr_14_0 : IN std_logic ;
         q_arr_15_31 : IN std_logic ;
         q_arr_15_30 : IN std_logic ;
         q_arr_15_29 : IN std_logic ;
         q_arr_15_28 : IN std_logic ;
         q_arr_15_27 : IN std_logic ;
         q_arr_15_26 : IN std_logic ;
         q_arr_15_25 : IN std_logic ;
         q_arr_15_24 : IN std_logic ;
         q_arr_15_23 : IN std_logic ;
         q_arr_15_22 : IN std_logic ;
         q_arr_15_21 : IN std_logic ;
         q_arr_15_20 : IN std_logic ;
         q_arr_15_19 : IN std_logic ;
         q_arr_15_18 : IN std_logic ;
         q_arr_15_17 : IN std_logic ;
         q_arr_15_16 : IN std_logic ;
         q_arr_15_15 : IN std_logic ;
         q_arr_15_14 : IN std_logic ;
         q_arr_15_13 : IN std_logic ;
         q_arr_15_12 : IN std_logic ;
         q_arr_15_11 : IN std_logic ;
         q_arr_15_10 : IN std_logic ;
         q_arr_15_9 : IN std_logic ;
         q_arr_15_8 : IN std_logic ;
         q_arr_15_7 : IN std_logic ;
         q_arr_15_6 : IN std_logic ;
         q_arr_15_5 : IN std_logic ;
         q_arr_15_4 : IN std_logic ;
         q_arr_15_3 : IN std_logic ;
         q_arr_15_2 : IN std_logic ;
         q_arr_15_1 : IN std_logic ;
         q_arr_15_0 : IN std_logic ;
         q_arr_16_31 : IN std_logic ;
         q_arr_16_30 : IN std_logic ;
         q_arr_16_29 : IN std_logic ;
         q_arr_16_28 : IN std_logic ;
         q_arr_16_27 : IN std_logic ;
         q_arr_16_26 : IN std_logic ;
         q_arr_16_25 : IN std_logic ;
         q_arr_16_24 : IN std_logic ;
         q_arr_16_23 : IN std_logic ;
         q_arr_16_22 : IN std_logic ;
         q_arr_16_21 : IN std_logic ;
         q_arr_16_20 : IN std_logic ;
         q_arr_16_19 : IN std_logic ;
         q_arr_16_18 : IN std_logic ;
         q_arr_16_17 : IN std_logic ;
         q_arr_16_16 : IN std_logic ;
         q_arr_16_15 : IN std_logic ;
         q_arr_16_14 : IN std_logic ;
         q_arr_16_13 : IN std_logic ;
         q_arr_16_12 : IN std_logic ;
         q_arr_16_11 : IN std_logic ;
         q_arr_16_10 : IN std_logic ;
         q_arr_16_9 : IN std_logic ;
         q_arr_16_8 : IN std_logic ;
         q_arr_16_7 : IN std_logic ;
         q_arr_16_6 : IN std_logic ;
         q_arr_16_5 : IN std_logic ;
         q_arr_16_4 : IN std_logic ;
         q_arr_16_3 : IN std_logic ;
         q_arr_16_2 : IN std_logic ;
         q_arr_16_1 : IN std_logic ;
         q_arr_16_0 : IN std_logic ;
         q_arr_17_31 : IN std_logic ;
         q_arr_17_30 : IN std_logic ;
         q_arr_17_29 : IN std_logic ;
         q_arr_17_28 : IN std_logic ;
         q_arr_17_27 : IN std_logic ;
         q_arr_17_26 : IN std_logic ;
         q_arr_17_25 : IN std_logic ;
         q_arr_17_24 : IN std_logic ;
         q_arr_17_23 : IN std_logic ;
         q_arr_17_22 : IN std_logic ;
         q_arr_17_21 : IN std_logic ;
         q_arr_17_20 : IN std_logic ;
         q_arr_17_19 : IN std_logic ;
         q_arr_17_18 : IN std_logic ;
         q_arr_17_17 : IN std_logic ;
         q_arr_17_16 : IN std_logic ;
         q_arr_17_15 : IN std_logic ;
         q_arr_17_14 : IN std_logic ;
         q_arr_17_13 : IN std_logic ;
         q_arr_17_12 : IN std_logic ;
         q_arr_17_11 : IN std_logic ;
         q_arr_17_10 : IN std_logic ;
         q_arr_17_9 : IN std_logic ;
         q_arr_17_8 : IN std_logic ;
         q_arr_17_7 : IN std_logic ;
         q_arr_17_6 : IN std_logic ;
         q_arr_17_5 : IN std_logic ;
         q_arr_17_4 : IN std_logic ;
         q_arr_17_3 : IN std_logic ;
         q_arr_17_2 : IN std_logic ;
         q_arr_17_1 : IN std_logic ;
         q_arr_17_0 : IN std_logic ;
         q_arr_18_31 : IN std_logic ;
         q_arr_18_30 : IN std_logic ;
         q_arr_18_29 : IN std_logic ;
         q_arr_18_28 : IN std_logic ;
         q_arr_18_27 : IN std_logic ;
         q_arr_18_26 : IN std_logic ;
         q_arr_18_25 : IN std_logic ;
         q_arr_18_24 : IN std_logic ;
         q_arr_18_23 : IN std_logic ;
         q_arr_18_22 : IN std_logic ;
         q_arr_18_21 : IN std_logic ;
         q_arr_18_20 : IN std_logic ;
         q_arr_18_19 : IN std_logic ;
         q_arr_18_18 : IN std_logic ;
         q_arr_18_17 : IN std_logic ;
         q_arr_18_16 : IN std_logic ;
         q_arr_18_15 : IN std_logic ;
         q_arr_18_14 : IN std_logic ;
         q_arr_18_13 : IN std_logic ;
         q_arr_18_12 : IN std_logic ;
         q_arr_18_11 : IN std_logic ;
         q_arr_18_10 : IN std_logic ;
         q_arr_18_9 : IN std_logic ;
         q_arr_18_8 : IN std_logic ;
         q_arr_18_7 : IN std_logic ;
         q_arr_18_6 : IN std_logic ;
         q_arr_18_5 : IN std_logic ;
         q_arr_18_4 : IN std_logic ;
         q_arr_18_3 : IN std_logic ;
         q_arr_18_2 : IN std_logic ;
         q_arr_18_1 : IN std_logic ;
         q_arr_18_0 : IN std_logic ;
         q_arr_19_31 : IN std_logic ;
         q_arr_19_30 : IN std_logic ;
         q_arr_19_29 : IN std_logic ;
         q_arr_19_28 : IN std_logic ;
         q_arr_19_27 : IN std_logic ;
         q_arr_19_26 : IN std_logic ;
         q_arr_19_25 : IN std_logic ;
         q_arr_19_24 : IN std_logic ;
         q_arr_19_23 : IN std_logic ;
         q_arr_19_22 : IN std_logic ;
         q_arr_19_21 : IN std_logic ;
         q_arr_19_20 : IN std_logic ;
         q_arr_19_19 : IN std_logic ;
         q_arr_19_18 : IN std_logic ;
         q_arr_19_17 : IN std_logic ;
         q_arr_19_16 : IN std_logic ;
         q_arr_19_15 : IN std_logic ;
         q_arr_19_14 : IN std_logic ;
         q_arr_19_13 : IN std_logic ;
         q_arr_19_12 : IN std_logic ;
         q_arr_19_11 : IN std_logic ;
         q_arr_19_10 : IN std_logic ;
         q_arr_19_9 : IN std_logic ;
         q_arr_19_8 : IN std_logic ;
         q_arr_19_7 : IN std_logic ;
         q_arr_19_6 : IN std_logic ;
         q_arr_19_5 : IN std_logic ;
         q_arr_19_4 : IN std_logic ;
         q_arr_19_3 : IN std_logic ;
         q_arr_19_2 : IN std_logic ;
         q_arr_19_1 : IN std_logic ;
         q_arr_19_0 : IN std_logic ;
         q_arr_20_31 : IN std_logic ;
         q_arr_20_30 : IN std_logic ;
         q_arr_20_29 : IN std_logic ;
         q_arr_20_28 : IN std_logic ;
         q_arr_20_27 : IN std_logic ;
         q_arr_20_26 : IN std_logic ;
         q_arr_20_25 : IN std_logic ;
         q_arr_20_24 : IN std_logic ;
         q_arr_20_23 : IN std_logic ;
         q_arr_20_22 : IN std_logic ;
         q_arr_20_21 : IN std_logic ;
         q_arr_20_20 : IN std_logic ;
         q_arr_20_19 : IN std_logic ;
         q_arr_20_18 : IN std_logic ;
         q_arr_20_17 : IN std_logic ;
         q_arr_20_16 : IN std_logic ;
         q_arr_20_15 : IN std_logic ;
         q_arr_20_14 : IN std_logic ;
         q_arr_20_13 : IN std_logic ;
         q_arr_20_12 : IN std_logic ;
         q_arr_20_11 : IN std_logic ;
         q_arr_20_10 : IN std_logic ;
         q_arr_20_9 : IN std_logic ;
         q_arr_20_8 : IN std_logic ;
         q_arr_20_7 : IN std_logic ;
         q_arr_20_6 : IN std_logic ;
         q_arr_20_5 : IN std_logic ;
         q_arr_20_4 : IN std_logic ;
         q_arr_20_3 : IN std_logic ;
         q_arr_20_2 : IN std_logic ;
         q_arr_20_1 : IN std_logic ;
         q_arr_20_0 : IN std_logic ;
         q_arr_21_31 : IN std_logic ;
         q_arr_21_30 : IN std_logic ;
         q_arr_21_29 : IN std_logic ;
         q_arr_21_28 : IN std_logic ;
         q_arr_21_27 : IN std_logic ;
         q_arr_21_26 : IN std_logic ;
         q_arr_21_25 : IN std_logic ;
         q_arr_21_24 : IN std_logic ;
         q_arr_21_23 : IN std_logic ;
         q_arr_21_22 : IN std_logic ;
         q_arr_21_21 : IN std_logic ;
         q_arr_21_20 : IN std_logic ;
         q_arr_21_19 : IN std_logic ;
         q_arr_21_18 : IN std_logic ;
         q_arr_21_17 : IN std_logic ;
         q_arr_21_16 : IN std_logic ;
         q_arr_21_15 : IN std_logic ;
         q_arr_21_14 : IN std_logic ;
         q_arr_21_13 : IN std_logic ;
         q_arr_21_12 : IN std_logic ;
         q_arr_21_11 : IN std_logic ;
         q_arr_21_10 : IN std_logic ;
         q_arr_21_9 : IN std_logic ;
         q_arr_21_8 : IN std_logic ;
         q_arr_21_7 : IN std_logic ;
         q_arr_21_6 : IN std_logic ;
         q_arr_21_5 : IN std_logic ;
         q_arr_21_4 : IN std_logic ;
         q_arr_21_3 : IN std_logic ;
         q_arr_21_2 : IN std_logic ;
         q_arr_21_1 : IN std_logic ;
         q_arr_21_0 : IN std_logic ;
         q_arr_22_31 : IN std_logic ;
         q_arr_22_30 : IN std_logic ;
         q_arr_22_29 : IN std_logic ;
         q_arr_22_28 : IN std_logic ;
         q_arr_22_27 : IN std_logic ;
         q_arr_22_26 : IN std_logic ;
         q_arr_22_25 : IN std_logic ;
         q_arr_22_24 : IN std_logic ;
         q_arr_22_23 : IN std_logic ;
         q_arr_22_22 : IN std_logic ;
         q_arr_22_21 : IN std_logic ;
         q_arr_22_20 : IN std_logic ;
         q_arr_22_19 : IN std_logic ;
         q_arr_22_18 : IN std_logic ;
         q_arr_22_17 : IN std_logic ;
         q_arr_22_16 : IN std_logic ;
         q_arr_22_15 : IN std_logic ;
         q_arr_22_14 : IN std_logic ;
         q_arr_22_13 : IN std_logic ;
         q_arr_22_12 : IN std_logic ;
         q_arr_22_11 : IN std_logic ;
         q_arr_22_10 : IN std_logic ;
         q_arr_22_9 : IN std_logic ;
         q_arr_22_8 : IN std_logic ;
         q_arr_22_7 : IN std_logic ;
         q_arr_22_6 : IN std_logic ;
         q_arr_22_5 : IN std_logic ;
         q_arr_22_4 : IN std_logic ;
         q_arr_22_3 : IN std_logic ;
         q_arr_22_2 : IN std_logic ;
         q_arr_22_1 : IN std_logic ;
         q_arr_22_0 : IN std_logic ;
         q_arr_23_31 : IN std_logic ;
         q_arr_23_30 : IN std_logic ;
         q_arr_23_29 : IN std_logic ;
         q_arr_23_28 : IN std_logic ;
         q_arr_23_27 : IN std_logic ;
         q_arr_23_26 : IN std_logic ;
         q_arr_23_25 : IN std_logic ;
         q_arr_23_24 : IN std_logic ;
         q_arr_23_23 : IN std_logic ;
         q_arr_23_22 : IN std_logic ;
         q_arr_23_21 : IN std_logic ;
         q_arr_23_20 : IN std_logic ;
         q_arr_23_19 : IN std_logic ;
         q_arr_23_18 : IN std_logic ;
         q_arr_23_17 : IN std_logic ;
         q_arr_23_16 : IN std_logic ;
         q_arr_23_15 : IN std_logic ;
         q_arr_23_14 : IN std_logic ;
         q_arr_23_13 : IN std_logic ;
         q_arr_23_12 : IN std_logic ;
         q_arr_23_11 : IN std_logic ;
         q_arr_23_10 : IN std_logic ;
         q_arr_23_9 : IN std_logic ;
         q_arr_23_8 : IN std_logic ;
         q_arr_23_7 : IN std_logic ;
         q_arr_23_6 : IN std_logic ;
         q_arr_23_5 : IN std_logic ;
         q_arr_23_4 : IN std_logic ;
         q_arr_23_3 : IN std_logic ;
         q_arr_23_2 : IN std_logic ;
         q_arr_23_1 : IN std_logic ;
         q_arr_23_0 : IN std_logic ;
         q_arr_24_31 : IN std_logic ;
         q_arr_24_30 : IN std_logic ;
         q_arr_24_29 : IN std_logic ;
         q_arr_24_28 : IN std_logic ;
         q_arr_24_27 : IN std_logic ;
         q_arr_24_26 : IN std_logic ;
         q_arr_24_25 : IN std_logic ;
         q_arr_24_24 : IN std_logic ;
         q_arr_24_23 : IN std_logic ;
         q_arr_24_22 : IN std_logic ;
         q_arr_24_21 : IN std_logic ;
         q_arr_24_20 : IN std_logic ;
         q_arr_24_19 : IN std_logic ;
         q_arr_24_18 : IN std_logic ;
         q_arr_24_17 : IN std_logic ;
         q_arr_24_16 : IN std_logic ;
         q_arr_24_15 : IN std_logic ;
         q_arr_24_14 : IN std_logic ;
         q_arr_24_13 : IN std_logic ;
         q_arr_24_12 : IN std_logic ;
         q_arr_24_11 : IN std_logic ;
         q_arr_24_10 : IN std_logic ;
         q_arr_24_9 : IN std_logic ;
         q_arr_24_8 : IN std_logic ;
         q_arr_24_7 : IN std_logic ;
         q_arr_24_6 : IN std_logic ;
         q_arr_24_5 : IN std_logic ;
         q_arr_24_4 : IN std_logic ;
         q_arr_24_3 : IN std_logic ;
         q_arr_24_2 : IN std_logic ;
         q_arr_24_1 : IN std_logic ;
         q_arr_24_0 : IN std_logic ;
         operation : IN std_logic ;
         filter_size : IN std_logic) ;
   end component ;
   component ReluLayer
      port (
         d_arr_0_31 : OUT std_logic ;
         d_arr_0_30 : OUT std_logic ;
         d_arr_0_29 : OUT std_logic ;
         d_arr_0_28 : OUT std_logic ;
         d_arr_0_27 : OUT std_logic ;
         d_arr_0_26 : OUT std_logic ;
         d_arr_0_25 : OUT std_logic ;
         d_arr_0_24 : OUT std_logic ;
         d_arr_0_23 : OUT std_logic ;
         d_arr_0_22 : OUT std_logic ;
         d_arr_0_21 : OUT std_logic ;
         d_arr_0_20 : OUT std_logic ;
         d_arr_0_19 : OUT std_logic ;
         d_arr_0_18 : OUT std_logic ;
         d_arr_0_17 : OUT std_logic ;
         d_arr_0_16 : OUT std_logic ;
         d_arr_0_15 : OUT std_logic ;
         d_arr_0_14 : OUT std_logic ;
         d_arr_0_13 : OUT std_logic ;
         d_arr_0_12 : OUT std_logic ;
         d_arr_0_11 : OUT std_logic ;
         d_arr_0_10 : OUT std_logic ;
         d_arr_0_9 : OUT std_logic ;
         d_arr_0_8 : OUT std_logic ;
         d_arr_0_7 : OUT std_logic ;
         d_arr_0_6 : OUT std_logic ;
         d_arr_0_5 : OUT std_logic ;
         d_arr_0_4 : OUT std_logic ;
         d_arr_0_3 : OUT std_logic ;
         d_arr_0_2 : OUT std_logic ;
         d_arr_0_1 : OUT std_logic ;
         d_arr_0_0 : OUT std_logic ;
         d_arr_1_31 : OUT std_logic ;
         d_arr_1_30 : OUT std_logic ;
         d_arr_1_29 : OUT std_logic ;
         d_arr_1_28 : OUT std_logic ;
         d_arr_1_27 : OUT std_logic ;
         d_arr_1_26 : OUT std_logic ;
         d_arr_1_25 : OUT std_logic ;
         d_arr_1_24 : OUT std_logic ;
         d_arr_1_23 : OUT std_logic ;
         d_arr_1_22 : OUT std_logic ;
         d_arr_1_21 : OUT std_logic ;
         d_arr_1_20 : OUT std_logic ;
         d_arr_1_19 : OUT std_logic ;
         d_arr_1_18 : OUT std_logic ;
         d_arr_1_17 : OUT std_logic ;
         d_arr_1_16 : OUT std_logic ;
         d_arr_1_15 : OUT std_logic ;
         d_arr_1_14 : OUT std_logic ;
         d_arr_1_13 : OUT std_logic ;
         d_arr_1_12 : OUT std_logic ;
         d_arr_1_11 : OUT std_logic ;
         d_arr_1_10 : OUT std_logic ;
         d_arr_1_9 : OUT std_logic ;
         d_arr_1_8 : OUT std_logic ;
         d_arr_1_7 : OUT std_logic ;
         d_arr_1_6 : OUT std_logic ;
         d_arr_1_5 : OUT std_logic ;
         d_arr_1_4 : OUT std_logic ;
         d_arr_1_3 : OUT std_logic ;
         d_arr_1_2 : OUT std_logic ;
         d_arr_1_1 : OUT std_logic ;
         d_arr_1_0 : OUT std_logic ;
         d_arr_2_31 : OUT std_logic ;
         d_arr_2_30 : OUT std_logic ;
         d_arr_2_29 : OUT std_logic ;
         d_arr_2_28 : OUT std_logic ;
         d_arr_2_27 : OUT std_logic ;
         d_arr_2_26 : OUT std_logic ;
         d_arr_2_25 : OUT std_logic ;
         d_arr_2_24 : OUT std_logic ;
         d_arr_2_23 : OUT std_logic ;
         d_arr_2_22 : OUT std_logic ;
         d_arr_2_21 : OUT std_logic ;
         d_arr_2_20 : OUT std_logic ;
         d_arr_2_19 : OUT std_logic ;
         d_arr_2_18 : OUT std_logic ;
         d_arr_2_17 : OUT std_logic ;
         d_arr_2_16 : OUT std_logic ;
         d_arr_2_15 : OUT std_logic ;
         d_arr_2_14 : OUT std_logic ;
         d_arr_2_13 : OUT std_logic ;
         d_arr_2_12 : OUT std_logic ;
         d_arr_2_11 : OUT std_logic ;
         d_arr_2_10 : OUT std_logic ;
         d_arr_2_9 : OUT std_logic ;
         d_arr_2_8 : OUT std_logic ;
         d_arr_2_7 : OUT std_logic ;
         d_arr_2_6 : OUT std_logic ;
         d_arr_2_5 : OUT std_logic ;
         d_arr_2_4 : OUT std_logic ;
         d_arr_2_3 : OUT std_logic ;
         d_arr_2_2 : OUT std_logic ;
         d_arr_2_1 : OUT std_logic ;
         d_arr_2_0 : OUT std_logic ;
         d_arr_3_31 : OUT std_logic ;
         d_arr_3_30 : OUT std_logic ;
         d_arr_3_29 : OUT std_logic ;
         d_arr_3_28 : OUT std_logic ;
         d_arr_3_27 : OUT std_logic ;
         d_arr_3_26 : OUT std_logic ;
         d_arr_3_25 : OUT std_logic ;
         d_arr_3_24 : OUT std_logic ;
         d_arr_3_23 : OUT std_logic ;
         d_arr_3_22 : OUT std_logic ;
         d_arr_3_21 : OUT std_logic ;
         d_arr_3_20 : OUT std_logic ;
         d_arr_3_19 : OUT std_logic ;
         d_arr_3_18 : OUT std_logic ;
         d_arr_3_17 : OUT std_logic ;
         d_arr_3_16 : OUT std_logic ;
         d_arr_3_15 : OUT std_logic ;
         d_arr_3_14 : OUT std_logic ;
         d_arr_3_13 : OUT std_logic ;
         d_arr_3_12 : OUT std_logic ;
         d_arr_3_11 : OUT std_logic ;
         d_arr_3_10 : OUT std_logic ;
         d_arr_3_9 : OUT std_logic ;
         d_arr_3_8 : OUT std_logic ;
         d_arr_3_7 : OUT std_logic ;
         d_arr_3_6 : OUT std_logic ;
         d_arr_3_5 : OUT std_logic ;
         d_arr_3_4 : OUT std_logic ;
         d_arr_3_3 : OUT std_logic ;
         d_arr_3_2 : OUT std_logic ;
         d_arr_3_1 : OUT std_logic ;
         d_arr_3_0 : OUT std_logic ;
         d_arr_4_31 : OUT std_logic ;
         d_arr_4_30 : OUT std_logic ;
         d_arr_4_29 : OUT std_logic ;
         d_arr_4_28 : OUT std_logic ;
         d_arr_4_27 : OUT std_logic ;
         d_arr_4_26 : OUT std_logic ;
         d_arr_4_25 : OUT std_logic ;
         d_arr_4_24 : OUT std_logic ;
         d_arr_4_23 : OUT std_logic ;
         d_arr_4_22 : OUT std_logic ;
         d_arr_4_21 : OUT std_logic ;
         d_arr_4_20 : OUT std_logic ;
         d_arr_4_19 : OUT std_logic ;
         d_arr_4_18 : OUT std_logic ;
         d_arr_4_17 : OUT std_logic ;
         d_arr_4_16 : OUT std_logic ;
         d_arr_4_15 : OUT std_logic ;
         d_arr_4_14 : OUT std_logic ;
         d_arr_4_13 : OUT std_logic ;
         d_arr_4_12 : OUT std_logic ;
         d_arr_4_11 : OUT std_logic ;
         d_arr_4_10 : OUT std_logic ;
         d_arr_4_9 : OUT std_logic ;
         d_arr_4_8 : OUT std_logic ;
         d_arr_4_7 : OUT std_logic ;
         d_arr_4_6 : OUT std_logic ;
         d_arr_4_5 : OUT std_logic ;
         d_arr_4_4 : OUT std_logic ;
         d_arr_4_3 : OUT std_logic ;
         d_arr_4_2 : OUT std_logic ;
         d_arr_4_1 : OUT std_logic ;
         d_arr_4_0 : OUT std_logic ;
         d_arr_5_31 : OUT std_logic ;
         d_arr_5_30 : OUT std_logic ;
         d_arr_5_29 : OUT std_logic ;
         d_arr_5_28 : OUT std_logic ;
         d_arr_5_27 : OUT std_logic ;
         d_arr_5_26 : OUT std_logic ;
         d_arr_5_25 : OUT std_logic ;
         d_arr_5_24 : OUT std_logic ;
         d_arr_5_23 : OUT std_logic ;
         d_arr_5_22 : OUT std_logic ;
         d_arr_5_21 : OUT std_logic ;
         d_arr_5_20 : OUT std_logic ;
         d_arr_5_19 : OUT std_logic ;
         d_arr_5_18 : OUT std_logic ;
         d_arr_5_17 : OUT std_logic ;
         d_arr_5_16 : OUT std_logic ;
         d_arr_5_15 : OUT std_logic ;
         d_arr_5_14 : OUT std_logic ;
         d_arr_5_13 : OUT std_logic ;
         d_arr_5_12 : OUT std_logic ;
         d_arr_5_11 : OUT std_logic ;
         d_arr_5_10 : OUT std_logic ;
         d_arr_5_9 : OUT std_logic ;
         d_arr_5_8 : OUT std_logic ;
         d_arr_5_7 : OUT std_logic ;
         d_arr_5_6 : OUT std_logic ;
         d_arr_5_5 : OUT std_logic ;
         d_arr_5_4 : OUT std_logic ;
         d_arr_5_3 : OUT std_logic ;
         d_arr_5_2 : OUT std_logic ;
         d_arr_5_1 : OUT std_logic ;
         d_arr_5_0 : OUT std_logic ;
         d_arr_6_31 : OUT std_logic ;
         d_arr_6_30 : OUT std_logic ;
         d_arr_6_29 : OUT std_logic ;
         d_arr_6_28 : OUT std_logic ;
         d_arr_6_27 : OUT std_logic ;
         d_arr_6_26 : OUT std_logic ;
         d_arr_6_25 : OUT std_logic ;
         d_arr_6_24 : OUT std_logic ;
         d_arr_6_23 : OUT std_logic ;
         d_arr_6_22 : OUT std_logic ;
         d_arr_6_21 : OUT std_logic ;
         d_arr_6_20 : OUT std_logic ;
         d_arr_6_19 : OUT std_logic ;
         d_arr_6_18 : OUT std_logic ;
         d_arr_6_17 : OUT std_logic ;
         d_arr_6_16 : OUT std_logic ;
         d_arr_6_15 : OUT std_logic ;
         d_arr_6_14 : OUT std_logic ;
         d_arr_6_13 : OUT std_logic ;
         d_arr_6_12 : OUT std_logic ;
         d_arr_6_11 : OUT std_logic ;
         d_arr_6_10 : OUT std_logic ;
         d_arr_6_9 : OUT std_logic ;
         d_arr_6_8 : OUT std_logic ;
         d_arr_6_7 : OUT std_logic ;
         d_arr_6_6 : OUT std_logic ;
         d_arr_6_5 : OUT std_logic ;
         d_arr_6_4 : OUT std_logic ;
         d_arr_6_3 : OUT std_logic ;
         d_arr_6_2 : OUT std_logic ;
         d_arr_6_1 : OUT std_logic ;
         d_arr_6_0 : OUT std_logic ;
         d_arr_7_31 : OUT std_logic ;
         d_arr_7_30 : OUT std_logic ;
         d_arr_7_29 : OUT std_logic ;
         d_arr_7_28 : OUT std_logic ;
         d_arr_7_27 : OUT std_logic ;
         d_arr_7_26 : OUT std_logic ;
         d_arr_7_25 : OUT std_logic ;
         d_arr_7_24 : OUT std_logic ;
         d_arr_7_23 : OUT std_logic ;
         d_arr_7_22 : OUT std_logic ;
         d_arr_7_21 : OUT std_logic ;
         d_arr_7_20 : OUT std_logic ;
         d_arr_7_19 : OUT std_logic ;
         d_arr_7_18 : OUT std_logic ;
         d_arr_7_17 : OUT std_logic ;
         d_arr_7_16 : OUT std_logic ;
         d_arr_7_15 : OUT std_logic ;
         d_arr_7_14 : OUT std_logic ;
         d_arr_7_13 : OUT std_logic ;
         d_arr_7_12 : OUT std_logic ;
         d_arr_7_11 : OUT std_logic ;
         d_arr_7_10 : OUT std_logic ;
         d_arr_7_9 : OUT std_logic ;
         d_arr_7_8 : OUT std_logic ;
         d_arr_7_7 : OUT std_logic ;
         d_arr_7_6 : OUT std_logic ;
         d_arr_7_5 : OUT std_logic ;
         d_arr_7_4 : OUT std_logic ;
         d_arr_7_3 : OUT std_logic ;
         d_arr_7_2 : OUT std_logic ;
         d_arr_7_1 : OUT std_logic ;
         d_arr_7_0 : OUT std_logic ;
         d_arr_8_31 : OUT std_logic ;
         d_arr_8_30 : OUT std_logic ;
         d_arr_8_29 : OUT std_logic ;
         d_arr_8_28 : OUT std_logic ;
         d_arr_8_27 : OUT std_logic ;
         d_arr_8_26 : OUT std_logic ;
         d_arr_8_25 : OUT std_logic ;
         d_arr_8_24 : OUT std_logic ;
         d_arr_8_23 : OUT std_logic ;
         d_arr_8_22 : OUT std_logic ;
         d_arr_8_21 : OUT std_logic ;
         d_arr_8_20 : OUT std_logic ;
         d_arr_8_19 : OUT std_logic ;
         d_arr_8_18 : OUT std_logic ;
         d_arr_8_17 : OUT std_logic ;
         d_arr_8_16 : OUT std_logic ;
         d_arr_8_15 : OUT std_logic ;
         d_arr_8_14 : OUT std_logic ;
         d_arr_8_13 : OUT std_logic ;
         d_arr_8_12 : OUT std_logic ;
         d_arr_8_11 : OUT std_logic ;
         d_arr_8_10 : OUT std_logic ;
         d_arr_8_9 : OUT std_logic ;
         d_arr_8_8 : OUT std_logic ;
         d_arr_8_7 : OUT std_logic ;
         d_arr_8_6 : OUT std_logic ;
         d_arr_8_5 : OUT std_logic ;
         d_arr_8_4 : OUT std_logic ;
         d_arr_8_3 : OUT std_logic ;
         d_arr_8_2 : OUT std_logic ;
         d_arr_8_1 : OUT std_logic ;
         d_arr_8_0 : OUT std_logic ;
         d_arr_9_31 : OUT std_logic ;
         d_arr_9_30 : OUT std_logic ;
         d_arr_9_29 : OUT std_logic ;
         d_arr_9_28 : OUT std_logic ;
         d_arr_9_27 : OUT std_logic ;
         d_arr_9_26 : OUT std_logic ;
         d_arr_9_25 : OUT std_logic ;
         d_arr_9_24 : OUT std_logic ;
         d_arr_9_23 : OUT std_logic ;
         d_arr_9_22 : OUT std_logic ;
         d_arr_9_21 : OUT std_logic ;
         d_arr_9_20 : OUT std_logic ;
         d_arr_9_19 : OUT std_logic ;
         d_arr_9_18 : OUT std_logic ;
         d_arr_9_17 : OUT std_logic ;
         d_arr_9_16 : OUT std_logic ;
         d_arr_9_15 : OUT std_logic ;
         d_arr_9_14 : OUT std_logic ;
         d_arr_9_13 : OUT std_logic ;
         d_arr_9_12 : OUT std_logic ;
         d_arr_9_11 : OUT std_logic ;
         d_arr_9_10 : OUT std_logic ;
         d_arr_9_9 : OUT std_logic ;
         d_arr_9_8 : OUT std_logic ;
         d_arr_9_7 : OUT std_logic ;
         d_arr_9_6 : OUT std_logic ;
         d_arr_9_5 : OUT std_logic ;
         d_arr_9_4 : OUT std_logic ;
         d_arr_9_3 : OUT std_logic ;
         d_arr_9_2 : OUT std_logic ;
         d_arr_9_1 : OUT std_logic ;
         d_arr_9_0 : OUT std_logic ;
         d_arr_10_31 : OUT std_logic ;
         d_arr_10_30 : OUT std_logic ;
         d_arr_10_29 : OUT std_logic ;
         d_arr_10_28 : OUT std_logic ;
         d_arr_10_27 : OUT std_logic ;
         d_arr_10_26 : OUT std_logic ;
         d_arr_10_25 : OUT std_logic ;
         d_arr_10_24 : OUT std_logic ;
         d_arr_10_23 : OUT std_logic ;
         d_arr_10_22 : OUT std_logic ;
         d_arr_10_21 : OUT std_logic ;
         d_arr_10_20 : OUT std_logic ;
         d_arr_10_19 : OUT std_logic ;
         d_arr_10_18 : OUT std_logic ;
         d_arr_10_17 : OUT std_logic ;
         d_arr_10_16 : OUT std_logic ;
         d_arr_10_15 : OUT std_logic ;
         d_arr_10_14 : OUT std_logic ;
         d_arr_10_13 : OUT std_logic ;
         d_arr_10_12 : OUT std_logic ;
         d_arr_10_11 : OUT std_logic ;
         d_arr_10_10 : OUT std_logic ;
         d_arr_10_9 : OUT std_logic ;
         d_arr_10_8 : OUT std_logic ;
         d_arr_10_7 : OUT std_logic ;
         d_arr_10_6 : OUT std_logic ;
         d_arr_10_5 : OUT std_logic ;
         d_arr_10_4 : OUT std_logic ;
         d_arr_10_3 : OUT std_logic ;
         d_arr_10_2 : OUT std_logic ;
         d_arr_10_1 : OUT std_logic ;
         d_arr_10_0 : OUT std_logic ;
         d_arr_11_31 : OUT std_logic ;
         d_arr_11_30 : OUT std_logic ;
         d_arr_11_29 : OUT std_logic ;
         d_arr_11_28 : OUT std_logic ;
         d_arr_11_27 : OUT std_logic ;
         d_arr_11_26 : OUT std_logic ;
         d_arr_11_25 : OUT std_logic ;
         d_arr_11_24 : OUT std_logic ;
         d_arr_11_23 : OUT std_logic ;
         d_arr_11_22 : OUT std_logic ;
         d_arr_11_21 : OUT std_logic ;
         d_arr_11_20 : OUT std_logic ;
         d_arr_11_19 : OUT std_logic ;
         d_arr_11_18 : OUT std_logic ;
         d_arr_11_17 : OUT std_logic ;
         d_arr_11_16 : OUT std_logic ;
         d_arr_11_15 : OUT std_logic ;
         d_arr_11_14 : OUT std_logic ;
         d_arr_11_13 : OUT std_logic ;
         d_arr_11_12 : OUT std_logic ;
         d_arr_11_11 : OUT std_logic ;
         d_arr_11_10 : OUT std_logic ;
         d_arr_11_9 : OUT std_logic ;
         d_arr_11_8 : OUT std_logic ;
         d_arr_11_7 : OUT std_logic ;
         d_arr_11_6 : OUT std_logic ;
         d_arr_11_5 : OUT std_logic ;
         d_arr_11_4 : OUT std_logic ;
         d_arr_11_3 : OUT std_logic ;
         d_arr_11_2 : OUT std_logic ;
         d_arr_11_1 : OUT std_logic ;
         d_arr_11_0 : OUT std_logic ;
         d_arr_12_31 : OUT std_logic ;
         d_arr_12_30 : OUT std_logic ;
         d_arr_12_29 : OUT std_logic ;
         d_arr_12_28 : OUT std_logic ;
         d_arr_12_27 : OUT std_logic ;
         d_arr_12_26 : OUT std_logic ;
         d_arr_12_25 : OUT std_logic ;
         d_arr_12_24 : OUT std_logic ;
         d_arr_12_23 : OUT std_logic ;
         d_arr_12_22 : OUT std_logic ;
         d_arr_12_21 : OUT std_logic ;
         d_arr_12_20 : OUT std_logic ;
         d_arr_12_19 : OUT std_logic ;
         d_arr_12_18 : OUT std_logic ;
         d_arr_12_17 : OUT std_logic ;
         d_arr_12_16 : OUT std_logic ;
         d_arr_12_15 : OUT std_logic ;
         d_arr_12_14 : OUT std_logic ;
         d_arr_12_13 : OUT std_logic ;
         d_arr_12_12 : OUT std_logic ;
         d_arr_12_11 : OUT std_logic ;
         d_arr_12_10 : OUT std_logic ;
         d_arr_12_9 : OUT std_logic ;
         d_arr_12_8 : OUT std_logic ;
         d_arr_12_7 : OUT std_logic ;
         d_arr_12_6 : OUT std_logic ;
         d_arr_12_5 : OUT std_logic ;
         d_arr_12_4 : OUT std_logic ;
         d_arr_12_3 : OUT std_logic ;
         d_arr_12_2 : OUT std_logic ;
         d_arr_12_1 : OUT std_logic ;
         d_arr_12_0 : OUT std_logic ;
         d_arr_13_31 : OUT std_logic ;
         d_arr_13_30 : OUT std_logic ;
         d_arr_13_29 : OUT std_logic ;
         d_arr_13_28 : OUT std_logic ;
         d_arr_13_27 : OUT std_logic ;
         d_arr_13_26 : OUT std_logic ;
         d_arr_13_25 : OUT std_logic ;
         d_arr_13_24 : OUT std_logic ;
         d_arr_13_23 : OUT std_logic ;
         d_arr_13_22 : OUT std_logic ;
         d_arr_13_21 : OUT std_logic ;
         d_arr_13_20 : OUT std_logic ;
         d_arr_13_19 : OUT std_logic ;
         d_arr_13_18 : OUT std_logic ;
         d_arr_13_17 : OUT std_logic ;
         d_arr_13_16 : OUT std_logic ;
         d_arr_13_15 : OUT std_logic ;
         d_arr_13_14 : OUT std_logic ;
         d_arr_13_13 : OUT std_logic ;
         d_arr_13_12 : OUT std_logic ;
         d_arr_13_11 : OUT std_logic ;
         d_arr_13_10 : OUT std_logic ;
         d_arr_13_9 : OUT std_logic ;
         d_arr_13_8 : OUT std_logic ;
         d_arr_13_7 : OUT std_logic ;
         d_arr_13_6 : OUT std_logic ;
         d_arr_13_5 : OUT std_logic ;
         d_arr_13_4 : OUT std_logic ;
         d_arr_13_3 : OUT std_logic ;
         d_arr_13_2 : OUT std_logic ;
         d_arr_13_1 : OUT std_logic ;
         d_arr_13_0 : OUT std_logic ;
         d_arr_14_31 : OUT std_logic ;
         d_arr_14_30 : OUT std_logic ;
         d_arr_14_29 : OUT std_logic ;
         d_arr_14_28 : OUT std_logic ;
         d_arr_14_27 : OUT std_logic ;
         d_arr_14_26 : OUT std_logic ;
         d_arr_14_25 : OUT std_logic ;
         d_arr_14_24 : OUT std_logic ;
         d_arr_14_23 : OUT std_logic ;
         d_arr_14_22 : OUT std_logic ;
         d_arr_14_21 : OUT std_logic ;
         d_arr_14_20 : OUT std_logic ;
         d_arr_14_19 : OUT std_logic ;
         d_arr_14_18 : OUT std_logic ;
         d_arr_14_17 : OUT std_logic ;
         d_arr_14_16 : OUT std_logic ;
         d_arr_14_15 : OUT std_logic ;
         d_arr_14_14 : OUT std_logic ;
         d_arr_14_13 : OUT std_logic ;
         d_arr_14_12 : OUT std_logic ;
         d_arr_14_11 : OUT std_logic ;
         d_arr_14_10 : OUT std_logic ;
         d_arr_14_9 : OUT std_logic ;
         d_arr_14_8 : OUT std_logic ;
         d_arr_14_7 : OUT std_logic ;
         d_arr_14_6 : OUT std_logic ;
         d_arr_14_5 : OUT std_logic ;
         d_arr_14_4 : OUT std_logic ;
         d_arr_14_3 : OUT std_logic ;
         d_arr_14_2 : OUT std_logic ;
         d_arr_14_1 : OUT std_logic ;
         d_arr_14_0 : OUT std_logic ;
         d_arr_15_31 : OUT std_logic ;
         d_arr_15_30 : OUT std_logic ;
         d_arr_15_29 : OUT std_logic ;
         d_arr_15_28 : OUT std_logic ;
         d_arr_15_27 : OUT std_logic ;
         d_arr_15_26 : OUT std_logic ;
         d_arr_15_25 : OUT std_logic ;
         d_arr_15_24 : OUT std_logic ;
         d_arr_15_23 : OUT std_logic ;
         d_arr_15_22 : OUT std_logic ;
         d_arr_15_21 : OUT std_logic ;
         d_arr_15_20 : OUT std_logic ;
         d_arr_15_19 : OUT std_logic ;
         d_arr_15_18 : OUT std_logic ;
         d_arr_15_17 : OUT std_logic ;
         d_arr_15_16 : OUT std_logic ;
         d_arr_15_15 : OUT std_logic ;
         d_arr_15_14 : OUT std_logic ;
         d_arr_15_13 : OUT std_logic ;
         d_arr_15_12 : OUT std_logic ;
         d_arr_15_11 : OUT std_logic ;
         d_arr_15_10 : OUT std_logic ;
         d_arr_15_9 : OUT std_logic ;
         d_arr_15_8 : OUT std_logic ;
         d_arr_15_7 : OUT std_logic ;
         d_arr_15_6 : OUT std_logic ;
         d_arr_15_5 : OUT std_logic ;
         d_arr_15_4 : OUT std_logic ;
         d_arr_15_3 : OUT std_logic ;
         d_arr_15_2 : OUT std_logic ;
         d_arr_15_1 : OUT std_logic ;
         d_arr_15_0 : OUT std_logic ;
         d_arr_16_31 : OUT std_logic ;
         d_arr_16_30 : OUT std_logic ;
         d_arr_16_29 : OUT std_logic ;
         d_arr_16_28 : OUT std_logic ;
         d_arr_16_27 : OUT std_logic ;
         d_arr_16_26 : OUT std_logic ;
         d_arr_16_25 : OUT std_logic ;
         d_arr_16_24 : OUT std_logic ;
         d_arr_16_23 : OUT std_logic ;
         d_arr_16_22 : OUT std_logic ;
         d_arr_16_21 : OUT std_logic ;
         d_arr_16_20 : OUT std_logic ;
         d_arr_16_19 : OUT std_logic ;
         d_arr_16_18 : OUT std_logic ;
         d_arr_16_17 : OUT std_logic ;
         d_arr_16_16 : OUT std_logic ;
         d_arr_16_15 : OUT std_logic ;
         d_arr_16_14 : OUT std_logic ;
         d_arr_16_13 : OUT std_logic ;
         d_arr_16_12 : OUT std_logic ;
         d_arr_16_11 : OUT std_logic ;
         d_arr_16_10 : OUT std_logic ;
         d_arr_16_9 : OUT std_logic ;
         d_arr_16_8 : OUT std_logic ;
         d_arr_16_7 : OUT std_logic ;
         d_arr_16_6 : OUT std_logic ;
         d_arr_16_5 : OUT std_logic ;
         d_arr_16_4 : OUT std_logic ;
         d_arr_16_3 : OUT std_logic ;
         d_arr_16_2 : OUT std_logic ;
         d_arr_16_1 : OUT std_logic ;
         d_arr_16_0 : OUT std_logic ;
         d_arr_17_31 : OUT std_logic ;
         d_arr_17_30 : OUT std_logic ;
         d_arr_17_29 : OUT std_logic ;
         d_arr_17_28 : OUT std_logic ;
         d_arr_17_27 : OUT std_logic ;
         d_arr_17_26 : OUT std_logic ;
         d_arr_17_25 : OUT std_logic ;
         d_arr_17_24 : OUT std_logic ;
         d_arr_17_23 : OUT std_logic ;
         d_arr_17_22 : OUT std_logic ;
         d_arr_17_21 : OUT std_logic ;
         d_arr_17_20 : OUT std_logic ;
         d_arr_17_19 : OUT std_logic ;
         d_arr_17_18 : OUT std_logic ;
         d_arr_17_17 : OUT std_logic ;
         d_arr_17_16 : OUT std_logic ;
         d_arr_17_15 : OUT std_logic ;
         d_arr_17_14 : OUT std_logic ;
         d_arr_17_13 : OUT std_logic ;
         d_arr_17_12 : OUT std_logic ;
         d_arr_17_11 : OUT std_logic ;
         d_arr_17_10 : OUT std_logic ;
         d_arr_17_9 : OUT std_logic ;
         d_arr_17_8 : OUT std_logic ;
         d_arr_17_7 : OUT std_logic ;
         d_arr_17_6 : OUT std_logic ;
         d_arr_17_5 : OUT std_logic ;
         d_arr_17_4 : OUT std_logic ;
         d_arr_17_3 : OUT std_logic ;
         d_arr_17_2 : OUT std_logic ;
         d_arr_17_1 : OUT std_logic ;
         d_arr_17_0 : OUT std_logic ;
         d_arr_18_31 : OUT std_logic ;
         d_arr_18_30 : OUT std_logic ;
         d_arr_18_29 : OUT std_logic ;
         d_arr_18_28 : OUT std_logic ;
         d_arr_18_27 : OUT std_logic ;
         d_arr_18_26 : OUT std_logic ;
         d_arr_18_25 : OUT std_logic ;
         d_arr_18_24 : OUT std_logic ;
         d_arr_18_23 : OUT std_logic ;
         d_arr_18_22 : OUT std_logic ;
         d_arr_18_21 : OUT std_logic ;
         d_arr_18_20 : OUT std_logic ;
         d_arr_18_19 : OUT std_logic ;
         d_arr_18_18 : OUT std_logic ;
         d_arr_18_17 : OUT std_logic ;
         d_arr_18_16 : OUT std_logic ;
         d_arr_18_15 : OUT std_logic ;
         d_arr_18_14 : OUT std_logic ;
         d_arr_18_13 : OUT std_logic ;
         d_arr_18_12 : OUT std_logic ;
         d_arr_18_11 : OUT std_logic ;
         d_arr_18_10 : OUT std_logic ;
         d_arr_18_9 : OUT std_logic ;
         d_arr_18_8 : OUT std_logic ;
         d_arr_18_7 : OUT std_logic ;
         d_arr_18_6 : OUT std_logic ;
         d_arr_18_5 : OUT std_logic ;
         d_arr_18_4 : OUT std_logic ;
         d_arr_18_3 : OUT std_logic ;
         d_arr_18_2 : OUT std_logic ;
         d_arr_18_1 : OUT std_logic ;
         d_arr_18_0 : OUT std_logic ;
         d_arr_19_31 : OUT std_logic ;
         d_arr_19_30 : OUT std_logic ;
         d_arr_19_29 : OUT std_logic ;
         d_arr_19_28 : OUT std_logic ;
         d_arr_19_27 : OUT std_logic ;
         d_arr_19_26 : OUT std_logic ;
         d_arr_19_25 : OUT std_logic ;
         d_arr_19_24 : OUT std_logic ;
         d_arr_19_23 : OUT std_logic ;
         d_arr_19_22 : OUT std_logic ;
         d_arr_19_21 : OUT std_logic ;
         d_arr_19_20 : OUT std_logic ;
         d_arr_19_19 : OUT std_logic ;
         d_arr_19_18 : OUT std_logic ;
         d_arr_19_17 : OUT std_logic ;
         d_arr_19_16 : OUT std_logic ;
         d_arr_19_15 : OUT std_logic ;
         d_arr_19_14 : OUT std_logic ;
         d_arr_19_13 : OUT std_logic ;
         d_arr_19_12 : OUT std_logic ;
         d_arr_19_11 : OUT std_logic ;
         d_arr_19_10 : OUT std_logic ;
         d_arr_19_9 : OUT std_logic ;
         d_arr_19_8 : OUT std_logic ;
         d_arr_19_7 : OUT std_logic ;
         d_arr_19_6 : OUT std_logic ;
         d_arr_19_5 : OUT std_logic ;
         d_arr_19_4 : OUT std_logic ;
         d_arr_19_3 : OUT std_logic ;
         d_arr_19_2 : OUT std_logic ;
         d_arr_19_1 : OUT std_logic ;
         d_arr_19_0 : OUT std_logic ;
         d_arr_20_31 : OUT std_logic ;
         d_arr_20_30 : OUT std_logic ;
         d_arr_20_29 : OUT std_logic ;
         d_arr_20_28 : OUT std_logic ;
         d_arr_20_27 : OUT std_logic ;
         d_arr_20_26 : OUT std_logic ;
         d_arr_20_25 : OUT std_logic ;
         d_arr_20_24 : OUT std_logic ;
         d_arr_20_23 : OUT std_logic ;
         d_arr_20_22 : OUT std_logic ;
         d_arr_20_21 : OUT std_logic ;
         d_arr_20_20 : OUT std_logic ;
         d_arr_20_19 : OUT std_logic ;
         d_arr_20_18 : OUT std_logic ;
         d_arr_20_17 : OUT std_logic ;
         d_arr_20_16 : OUT std_logic ;
         d_arr_20_15 : OUT std_logic ;
         d_arr_20_14 : OUT std_logic ;
         d_arr_20_13 : OUT std_logic ;
         d_arr_20_12 : OUT std_logic ;
         d_arr_20_11 : OUT std_logic ;
         d_arr_20_10 : OUT std_logic ;
         d_arr_20_9 : OUT std_logic ;
         d_arr_20_8 : OUT std_logic ;
         d_arr_20_7 : OUT std_logic ;
         d_arr_20_6 : OUT std_logic ;
         d_arr_20_5 : OUT std_logic ;
         d_arr_20_4 : OUT std_logic ;
         d_arr_20_3 : OUT std_logic ;
         d_arr_20_2 : OUT std_logic ;
         d_arr_20_1 : OUT std_logic ;
         d_arr_20_0 : OUT std_logic ;
         d_arr_21_31 : OUT std_logic ;
         d_arr_21_30 : OUT std_logic ;
         d_arr_21_29 : OUT std_logic ;
         d_arr_21_28 : OUT std_logic ;
         d_arr_21_27 : OUT std_logic ;
         d_arr_21_26 : OUT std_logic ;
         d_arr_21_25 : OUT std_logic ;
         d_arr_21_24 : OUT std_logic ;
         d_arr_21_23 : OUT std_logic ;
         d_arr_21_22 : OUT std_logic ;
         d_arr_21_21 : OUT std_logic ;
         d_arr_21_20 : OUT std_logic ;
         d_arr_21_19 : OUT std_logic ;
         d_arr_21_18 : OUT std_logic ;
         d_arr_21_17 : OUT std_logic ;
         d_arr_21_16 : OUT std_logic ;
         d_arr_21_15 : OUT std_logic ;
         d_arr_21_14 : OUT std_logic ;
         d_arr_21_13 : OUT std_logic ;
         d_arr_21_12 : OUT std_logic ;
         d_arr_21_11 : OUT std_logic ;
         d_arr_21_10 : OUT std_logic ;
         d_arr_21_9 : OUT std_logic ;
         d_arr_21_8 : OUT std_logic ;
         d_arr_21_7 : OUT std_logic ;
         d_arr_21_6 : OUT std_logic ;
         d_arr_21_5 : OUT std_logic ;
         d_arr_21_4 : OUT std_logic ;
         d_arr_21_3 : OUT std_logic ;
         d_arr_21_2 : OUT std_logic ;
         d_arr_21_1 : OUT std_logic ;
         d_arr_21_0 : OUT std_logic ;
         d_arr_22_31 : OUT std_logic ;
         d_arr_22_30 : OUT std_logic ;
         d_arr_22_29 : OUT std_logic ;
         d_arr_22_28 : OUT std_logic ;
         d_arr_22_27 : OUT std_logic ;
         d_arr_22_26 : OUT std_logic ;
         d_arr_22_25 : OUT std_logic ;
         d_arr_22_24 : OUT std_logic ;
         d_arr_22_23 : OUT std_logic ;
         d_arr_22_22 : OUT std_logic ;
         d_arr_22_21 : OUT std_logic ;
         d_arr_22_20 : OUT std_logic ;
         d_arr_22_19 : OUT std_logic ;
         d_arr_22_18 : OUT std_logic ;
         d_arr_22_17 : OUT std_logic ;
         d_arr_22_16 : OUT std_logic ;
         d_arr_22_15 : OUT std_logic ;
         d_arr_22_14 : OUT std_logic ;
         d_arr_22_13 : OUT std_logic ;
         d_arr_22_12 : OUT std_logic ;
         d_arr_22_11 : OUT std_logic ;
         d_arr_22_10 : OUT std_logic ;
         d_arr_22_9 : OUT std_logic ;
         d_arr_22_8 : OUT std_logic ;
         d_arr_22_7 : OUT std_logic ;
         d_arr_22_6 : OUT std_logic ;
         d_arr_22_5 : OUT std_logic ;
         d_arr_22_4 : OUT std_logic ;
         d_arr_22_3 : OUT std_logic ;
         d_arr_22_2 : OUT std_logic ;
         d_arr_22_1 : OUT std_logic ;
         d_arr_22_0 : OUT std_logic ;
         d_arr_23_31 : OUT std_logic ;
         d_arr_23_30 : OUT std_logic ;
         d_arr_23_29 : OUT std_logic ;
         d_arr_23_28 : OUT std_logic ;
         d_arr_23_27 : OUT std_logic ;
         d_arr_23_26 : OUT std_logic ;
         d_arr_23_25 : OUT std_logic ;
         d_arr_23_24 : OUT std_logic ;
         d_arr_23_23 : OUT std_logic ;
         d_arr_23_22 : OUT std_logic ;
         d_arr_23_21 : OUT std_logic ;
         d_arr_23_20 : OUT std_logic ;
         d_arr_23_19 : OUT std_logic ;
         d_arr_23_18 : OUT std_logic ;
         d_arr_23_17 : OUT std_logic ;
         d_arr_23_16 : OUT std_logic ;
         d_arr_23_15 : OUT std_logic ;
         d_arr_23_14 : OUT std_logic ;
         d_arr_23_13 : OUT std_logic ;
         d_arr_23_12 : OUT std_logic ;
         d_arr_23_11 : OUT std_logic ;
         d_arr_23_10 : OUT std_logic ;
         d_arr_23_9 : OUT std_logic ;
         d_arr_23_8 : OUT std_logic ;
         d_arr_23_7 : OUT std_logic ;
         d_arr_23_6 : OUT std_logic ;
         d_arr_23_5 : OUT std_logic ;
         d_arr_23_4 : OUT std_logic ;
         d_arr_23_3 : OUT std_logic ;
         d_arr_23_2 : OUT std_logic ;
         d_arr_23_1 : OUT std_logic ;
         d_arr_23_0 : OUT std_logic ;
         d_arr_24_31 : OUT std_logic ;
         d_arr_24_30 : OUT std_logic ;
         d_arr_24_29 : OUT std_logic ;
         d_arr_24_28 : OUT std_logic ;
         d_arr_24_27 : OUT std_logic ;
         d_arr_24_26 : OUT std_logic ;
         d_arr_24_25 : OUT std_logic ;
         d_arr_24_24 : OUT std_logic ;
         d_arr_24_23 : OUT std_logic ;
         d_arr_24_22 : OUT std_logic ;
         d_arr_24_21 : OUT std_logic ;
         d_arr_24_20 : OUT std_logic ;
         d_arr_24_19 : OUT std_logic ;
         d_arr_24_18 : OUT std_logic ;
         d_arr_24_17 : OUT std_logic ;
         d_arr_24_16 : OUT std_logic ;
         d_arr_24_15 : OUT std_logic ;
         d_arr_24_14 : OUT std_logic ;
         d_arr_24_13 : OUT std_logic ;
         d_arr_24_12 : OUT std_logic ;
         d_arr_24_11 : OUT std_logic ;
         d_arr_24_10 : OUT std_logic ;
         d_arr_24_9 : OUT std_logic ;
         d_arr_24_8 : OUT std_logic ;
         d_arr_24_7 : OUT std_logic ;
         d_arr_24_6 : OUT std_logic ;
         d_arr_24_5 : OUT std_logic ;
         d_arr_24_4 : OUT std_logic ;
         d_arr_24_3 : OUT std_logic ;
         d_arr_24_2 : OUT std_logic ;
         d_arr_24_1 : OUT std_logic ;
         d_arr_24_0 : OUT std_logic ;
         q_arr_0_31 : IN std_logic ;
         q_arr_0_30 : IN std_logic ;
         q_arr_0_29 : IN std_logic ;
         q_arr_0_28 : IN std_logic ;
         q_arr_0_27 : IN std_logic ;
         q_arr_0_26 : IN std_logic ;
         q_arr_0_25 : IN std_logic ;
         q_arr_0_24 : IN std_logic ;
         q_arr_0_23 : IN std_logic ;
         q_arr_0_22 : IN std_logic ;
         q_arr_0_21 : IN std_logic ;
         q_arr_0_20 : IN std_logic ;
         q_arr_0_19 : IN std_logic ;
         q_arr_0_18 : IN std_logic ;
         q_arr_0_17 : IN std_logic ;
         q_arr_0_16 : IN std_logic ;
         q_arr_0_15 : IN std_logic ;
         q_arr_0_14 : IN std_logic ;
         q_arr_0_13 : IN std_logic ;
         q_arr_0_12 : IN std_logic ;
         q_arr_0_11 : IN std_logic ;
         q_arr_0_10 : IN std_logic ;
         q_arr_0_9 : IN std_logic ;
         q_arr_0_8 : IN std_logic ;
         q_arr_0_7 : IN std_logic ;
         q_arr_0_6 : IN std_logic ;
         q_arr_0_5 : IN std_logic ;
         q_arr_0_4 : IN std_logic ;
         q_arr_0_3 : IN std_logic ;
         q_arr_0_2 : IN std_logic ;
         q_arr_0_1 : IN std_logic ;
         q_arr_0_0 : IN std_logic ;
         q_arr_1_31 : IN std_logic ;
         q_arr_1_30 : IN std_logic ;
         q_arr_1_29 : IN std_logic ;
         q_arr_1_28 : IN std_logic ;
         q_arr_1_27 : IN std_logic ;
         q_arr_1_26 : IN std_logic ;
         q_arr_1_25 : IN std_logic ;
         q_arr_1_24 : IN std_logic ;
         q_arr_1_23 : IN std_logic ;
         q_arr_1_22 : IN std_logic ;
         q_arr_1_21 : IN std_logic ;
         q_arr_1_20 : IN std_logic ;
         q_arr_1_19 : IN std_logic ;
         q_arr_1_18 : IN std_logic ;
         q_arr_1_17 : IN std_logic ;
         q_arr_1_16 : IN std_logic ;
         q_arr_1_15 : IN std_logic ;
         q_arr_1_14 : IN std_logic ;
         q_arr_1_13 : IN std_logic ;
         q_arr_1_12 : IN std_logic ;
         q_arr_1_11 : IN std_logic ;
         q_arr_1_10 : IN std_logic ;
         q_arr_1_9 : IN std_logic ;
         q_arr_1_8 : IN std_logic ;
         q_arr_1_7 : IN std_logic ;
         q_arr_1_6 : IN std_logic ;
         q_arr_1_5 : IN std_logic ;
         q_arr_1_4 : IN std_logic ;
         q_arr_1_3 : IN std_logic ;
         q_arr_1_2 : IN std_logic ;
         q_arr_1_1 : IN std_logic ;
         q_arr_1_0 : IN std_logic ;
         q_arr_2_31 : IN std_logic ;
         q_arr_2_30 : IN std_logic ;
         q_arr_2_29 : IN std_logic ;
         q_arr_2_28 : IN std_logic ;
         q_arr_2_27 : IN std_logic ;
         q_arr_2_26 : IN std_logic ;
         q_arr_2_25 : IN std_logic ;
         q_arr_2_24 : IN std_logic ;
         q_arr_2_23 : IN std_logic ;
         q_arr_2_22 : IN std_logic ;
         q_arr_2_21 : IN std_logic ;
         q_arr_2_20 : IN std_logic ;
         q_arr_2_19 : IN std_logic ;
         q_arr_2_18 : IN std_logic ;
         q_arr_2_17 : IN std_logic ;
         q_arr_2_16 : IN std_logic ;
         q_arr_2_15 : IN std_logic ;
         q_arr_2_14 : IN std_logic ;
         q_arr_2_13 : IN std_logic ;
         q_arr_2_12 : IN std_logic ;
         q_arr_2_11 : IN std_logic ;
         q_arr_2_10 : IN std_logic ;
         q_arr_2_9 : IN std_logic ;
         q_arr_2_8 : IN std_logic ;
         q_arr_2_7 : IN std_logic ;
         q_arr_2_6 : IN std_logic ;
         q_arr_2_5 : IN std_logic ;
         q_arr_2_4 : IN std_logic ;
         q_arr_2_3 : IN std_logic ;
         q_arr_2_2 : IN std_logic ;
         q_arr_2_1 : IN std_logic ;
         q_arr_2_0 : IN std_logic ;
         q_arr_3_31 : IN std_logic ;
         q_arr_3_30 : IN std_logic ;
         q_arr_3_29 : IN std_logic ;
         q_arr_3_28 : IN std_logic ;
         q_arr_3_27 : IN std_logic ;
         q_arr_3_26 : IN std_logic ;
         q_arr_3_25 : IN std_logic ;
         q_arr_3_24 : IN std_logic ;
         q_arr_3_23 : IN std_logic ;
         q_arr_3_22 : IN std_logic ;
         q_arr_3_21 : IN std_logic ;
         q_arr_3_20 : IN std_logic ;
         q_arr_3_19 : IN std_logic ;
         q_arr_3_18 : IN std_logic ;
         q_arr_3_17 : IN std_logic ;
         q_arr_3_16 : IN std_logic ;
         q_arr_3_15 : IN std_logic ;
         q_arr_3_14 : IN std_logic ;
         q_arr_3_13 : IN std_logic ;
         q_arr_3_12 : IN std_logic ;
         q_arr_3_11 : IN std_logic ;
         q_arr_3_10 : IN std_logic ;
         q_arr_3_9 : IN std_logic ;
         q_arr_3_8 : IN std_logic ;
         q_arr_3_7 : IN std_logic ;
         q_arr_3_6 : IN std_logic ;
         q_arr_3_5 : IN std_logic ;
         q_arr_3_4 : IN std_logic ;
         q_arr_3_3 : IN std_logic ;
         q_arr_3_2 : IN std_logic ;
         q_arr_3_1 : IN std_logic ;
         q_arr_3_0 : IN std_logic ;
         q_arr_4_31 : IN std_logic ;
         q_arr_4_30 : IN std_logic ;
         q_arr_4_29 : IN std_logic ;
         q_arr_4_28 : IN std_logic ;
         q_arr_4_27 : IN std_logic ;
         q_arr_4_26 : IN std_logic ;
         q_arr_4_25 : IN std_logic ;
         q_arr_4_24 : IN std_logic ;
         q_arr_4_23 : IN std_logic ;
         q_arr_4_22 : IN std_logic ;
         q_arr_4_21 : IN std_logic ;
         q_arr_4_20 : IN std_logic ;
         q_arr_4_19 : IN std_logic ;
         q_arr_4_18 : IN std_logic ;
         q_arr_4_17 : IN std_logic ;
         q_arr_4_16 : IN std_logic ;
         q_arr_4_15 : IN std_logic ;
         q_arr_4_14 : IN std_logic ;
         q_arr_4_13 : IN std_logic ;
         q_arr_4_12 : IN std_logic ;
         q_arr_4_11 : IN std_logic ;
         q_arr_4_10 : IN std_logic ;
         q_arr_4_9 : IN std_logic ;
         q_arr_4_8 : IN std_logic ;
         q_arr_4_7 : IN std_logic ;
         q_arr_4_6 : IN std_logic ;
         q_arr_4_5 : IN std_logic ;
         q_arr_4_4 : IN std_logic ;
         q_arr_4_3 : IN std_logic ;
         q_arr_4_2 : IN std_logic ;
         q_arr_4_1 : IN std_logic ;
         q_arr_4_0 : IN std_logic ;
         q_arr_5_31 : IN std_logic ;
         q_arr_5_30 : IN std_logic ;
         q_arr_5_29 : IN std_logic ;
         q_arr_5_28 : IN std_logic ;
         q_arr_5_27 : IN std_logic ;
         q_arr_5_26 : IN std_logic ;
         q_arr_5_25 : IN std_logic ;
         q_arr_5_24 : IN std_logic ;
         q_arr_5_23 : IN std_logic ;
         q_arr_5_22 : IN std_logic ;
         q_arr_5_21 : IN std_logic ;
         q_arr_5_20 : IN std_logic ;
         q_arr_5_19 : IN std_logic ;
         q_arr_5_18 : IN std_logic ;
         q_arr_5_17 : IN std_logic ;
         q_arr_5_16 : IN std_logic ;
         q_arr_5_15 : IN std_logic ;
         q_arr_5_14 : IN std_logic ;
         q_arr_5_13 : IN std_logic ;
         q_arr_5_12 : IN std_logic ;
         q_arr_5_11 : IN std_logic ;
         q_arr_5_10 : IN std_logic ;
         q_arr_5_9 : IN std_logic ;
         q_arr_5_8 : IN std_logic ;
         q_arr_5_7 : IN std_logic ;
         q_arr_5_6 : IN std_logic ;
         q_arr_5_5 : IN std_logic ;
         q_arr_5_4 : IN std_logic ;
         q_arr_5_3 : IN std_logic ;
         q_arr_5_2 : IN std_logic ;
         q_arr_5_1 : IN std_logic ;
         q_arr_5_0 : IN std_logic ;
         q_arr_6_31 : IN std_logic ;
         q_arr_6_30 : IN std_logic ;
         q_arr_6_29 : IN std_logic ;
         q_arr_6_28 : IN std_logic ;
         q_arr_6_27 : IN std_logic ;
         q_arr_6_26 : IN std_logic ;
         q_arr_6_25 : IN std_logic ;
         q_arr_6_24 : IN std_logic ;
         q_arr_6_23 : IN std_logic ;
         q_arr_6_22 : IN std_logic ;
         q_arr_6_21 : IN std_logic ;
         q_arr_6_20 : IN std_logic ;
         q_arr_6_19 : IN std_logic ;
         q_arr_6_18 : IN std_logic ;
         q_arr_6_17 : IN std_logic ;
         q_arr_6_16 : IN std_logic ;
         q_arr_6_15 : IN std_logic ;
         q_arr_6_14 : IN std_logic ;
         q_arr_6_13 : IN std_logic ;
         q_arr_6_12 : IN std_logic ;
         q_arr_6_11 : IN std_logic ;
         q_arr_6_10 : IN std_logic ;
         q_arr_6_9 : IN std_logic ;
         q_arr_6_8 : IN std_logic ;
         q_arr_6_7 : IN std_logic ;
         q_arr_6_6 : IN std_logic ;
         q_arr_6_5 : IN std_logic ;
         q_arr_6_4 : IN std_logic ;
         q_arr_6_3 : IN std_logic ;
         q_arr_6_2 : IN std_logic ;
         q_arr_6_1 : IN std_logic ;
         q_arr_6_0 : IN std_logic ;
         q_arr_7_31 : IN std_logic ;
         q_arr_7_30 : IN std_logic ;
         q_arr_7_29 : IN std_logic ;
         q_arr_7_28 : IN std_logic ;
         q_arr_7_27 : IN std_logic ;
         q_arr_7_26 : IN std_logic ;
         q_arr_7_25 : IN std_logic ;
         q_arr_7_24 : IN std_logic ;
         q_arr_7_23 : IN std_logic ;
         q_arr_7_22 : IN std_logic ;
         q_arr_7_21 : IN std_logic ;
         q_arr_7_20 : IN std_logic ;
         q_arr_7_19 : IN std_logic ;
         q_arr_7_18 : IN std_logic ;
         q_arr_7_17 : IN std_logic ;
         q_arr_7_16 : IN std_logic ;
         q_arr_7_15 : IN std_logic ;
         q_arr_7_14 : IN std_logic ;
         q_arr_7_13 : IN std_logic ;
         q_arr_7_12 : IN std_logic ;
         q_arr_7_11 : IN std_logic ;
         q_arr_7_10 : IN std_logic ;
         q_arr_7_9 : IN std_logic ;
         q_arr_7_8 : IN std_logic ;
         q_arr_7_7 : IN std_logic ;
         q_arr_7_6 : IN std_logic ;
         q_arr_7_5 : IN std_logic ;
         q_arr_7_4 : IN std_logic ;
         q_arr_7_3 : IN std_logic ;
         q_arr_7_2 : IN std_logic ;
         q_arr_7_1 : IN std_logic ;
         q_arr_7_0 : IN std_logic ;
         q_arr_8_31 : IN std_logic ;
         q_arr_8_30 : IN std_logic ;
         q_arr_8_29 : IN std_logic ;
         q_arr_8_28 : IN std_logic ;
         q_arr_8_27 : IN std_logic ;
         q_arr_8_26 : IN std_logic ;
         q_arr_8_25 : IN std_logic ;
         q_arr_8_24 : IN std_logic ;
         q_arr_8_23 : IN std_logic ;
         q_arr_8_22 : IN std_logic ;
         q_arr_8_21 : IN std_logic ;
         q_arr_8_20 : IN std_logic ;
         q_arr_8_19 : IN std_logic ;
         q_arr_8_18 : IN std_logic ;
         q_arr_8_17 : IN std_logic ;
         q_arr_8_16 : IN std_logic ;
         q_arr_8_15 : IN std_logic ;
         q_arr_8_14 : IN std_logic ;
         q_arr_8_13 : IN std_logic ;
         q_arr_8_12 : IN std_logic ;
         q_arr_8_11 : IN std_logic ;
         q_arr_8_10 : IN std_logic ;
         q_arr_8_9 : IN std_logic ;
         q_arr_8_8 : IN std_logic ;
         q_arr_8_7 : IN std_logic ;
         q_arr_8_6 : IN std_logic ;
         q_arr_8_5 : IN std_logic ;
         q_arr_8_4 : IN std_logic ;
         q_arr_8_3 : IN std_logic ;
         q_arr_8_2 : IN std_logic ;
         q_arr_8_1 : IN std_logic ;
         q_arr_8_0 : IN std_logic ;
         q_arr_9_31 : IN std_logic ;
         q_arr_9_30 : IN std_logic ;
         q_arr_9_29 : IN std_logic ;
         q_arr_9_28 : IN std_logic ;
         q_arr_9_27 : IN std_logic ;
         q_arr_9_26 : IN std_logic ;
         q_arr_9_25 : IN std_logic ;
         q_arr_9_24 : IN std_logic ;
         q_arr_9_23 : IN std_logic ;
         q_arr_9_22 : IN std_logic ;
         q_arr_9_21 : IN std_logic ;
         q_arr_9_20 : IN std_logic ;
         q_arr_9_19 : IN std_logic ;
         q_arr_9_18 : IN std_logic ;
         q_arr_9_17 : IN std_logic ;
         q_arr_9_16 : IN std_logic ;
         q_arr_9_15 : IN std_logic ;
         q_arr_9_14 : IN std_logic ;
         q_arr_9_13 : IN std_logic ;
         q_arr_9_12 : IN std_logic ;
         q_arr_9_11 : IN std_logic ;
         q_arr_9_10 : IN std_logic ;
         q_arr_9_9 : IN std_logic ;
         q_arr_9_8 : IN std_logic ;
         q_arr_9_7 : IN std_logic ;
         q_arr_9_6 : IN std_logic ;
         q_arr_9_5 : IN std_logic ;
         q_arr_9_4 : IN std_logic ;
         q_arr_9_3 : IN std_logic ;
         q_arr_9_2 : IN std_logic ;
         q_arr_9_1 : IN std_logic ;
         q_arr_9_0 : IN std_logic ;
         q_arr_10_31 : IN std_logic ;
         q_arr_10_30 : IN std_logic ;
         q_arr_10_29 : IN std_logic ;
         q_arr_10_28 : IN std_logic ;
         q_arr_10_27 : IN std_logic ;
         q_arr_10_26 : IN std_logic ;
         q_arr_10_25 : IN std_logic ;
         q_arr_10_24 : IN std_logic ;
         q_arr_10_23 : IN std_logic ;
         q_arr_10_22 : IN std_logic ;
         q_arr_10_21 : IN std_logic ;
         q_arr_10_20 : IN std_logic ;
         q_arr_10_19 : IN std_logic ;
         q_arr_10_18 : IN std_logic ;
         q_arr_10_17 : IN std_logic ;
         q_arr_10_16 : IN std_logic ;
         q_arr_10_15 : IN std_logic ;
         q_arr_10_14 : IN std_logic ;
         q_arr_10_13 : IN std_logic ;
         q_arr_10_12 : IN std_logic ;
         q_arr_10_11 : IN std_logic ;
         q_arr_10_10 : IN std_logic ;
         q_arr_10_9 : IN std_logic ;
         q_arr_10_8 : IN std_logic ;
         q_arr_10_7 : IN std_logic ;
         q_arr_10_6 : IN std_logic ;
         q_arr_10_5 : IN std_logic ;
         q_arr_10_4 : IN std_logic ;
         q_arr_10_3 : IN std_logic ;
         q_arr_10_2 : IN std_logic ;
         q_arr_10_1 : IN std_logic ;
         q_arr_10_0 : IN std_logic ;
         q_arr_11_31 : IN std_logic ;
         q_arr_11_30 : IN std_logic ;
         q_arr_11_29 : IN std_logic ;
         q_arr_11_28 : IN std_logic ;
         q_arr_11_27 : IN std_logic ;
         q_arr_11_26 : IN std_logic ;
         q_arr_11_25 : IN std_logic ;
         q_arr_11_24 : IN std_logic ;
         q_arr_11_23 : IN std_logic ;
         q_arr_11_22 : IN std_logic ;
         q_arr_11_21 : IN std_logic ;
         q_arr_11_20 : IN std_logic ;
         q_arr_11_19 : IN std_logic ;
         q_arr_11_18 : IN std_logic ;
         q_arr_11_17 : IN std_logic ;
         q_arr_11_16 : IN std_logic ;
         q_arr_11_15 : IN std_logic ;
         q_arr_11_14 : IN std_logic ;
         q_arr_11_13 : IN std_logic ;
         q_arr_11_12 : IN std_logic ;
         q_arr_11_11 : IN std_logic ;
         q_arr_11_10 : IN std_logic ;
         q_arr_11_9 : IN std_logic ;
         q_arr_11_8 : IN std_logic ;
         q_arr_11_7 : IN std_logic ;
         q_arr_11_6 : IN std_logic ;
         q_arr_11_5 : IN std_logic ;
         q_arr_11_4 : IN std_logic ;
         q_arr_11_3 : IN std_logic ;
         q_arr_11_2 : IN std_logic ;
         q_arr_11_1 : IN std_logic ;
         q_arr_11_0 : IN std_logic ;
         q_arr_12_31 : IN std_logic ;
         q_arr_12_30 : IN std_logic ;
         q_arr_12_29 : IN std_logic ;
         q_arr_12_28 : IN std_logic ;
         q_arr_12_27 : IN std_logic ;
         q_arr_12_26 : IN std_logic ;
         q_arr_12_25 : IN std_logic ;
         q_arr_12_24 : IN std_logic ;
         q_arr_12_23 : IN std_logic ;
         q_arr_12_22 : IN std_logic ;
         q_arr_12_21 : IN std_logic ;
         q_arr_12_20 : IN std_logic ;
         q_arr_12_19 : IN std_logic ;
         q_arr_12_18 : IN std_logic ;
         q_arr_12_17 : IN std_logic ;
         q_arr_12_16 : IN std_logic ;
         q_arr_12_15 : IN std_logic ;
         q_arr_12_14 : IN std_logic ;
         q_arr_12_13 : IN std_logic ;
         q_arr_12_12 : IN std_logic ;
         q_arr_12_11 : IN std_logic ;
         q_arr_12_10 : IN std_logic ;
         q_arr_12_9 : IN std_logic ;
         q_arr_12_8 : IN std_logic ;
         q_arr_12_7 : IN std_logic ;
         q_arr_12_6 : IN std_logic ;
         q_arr_12_5 : IN std_logic ;
         q_arr_12_4 : IN std_logic ;
         q_arr_12_3 : IN std_logic ;
         q_arr_12_2 : IN std_logic ;
         q_arr_12_1 : IN std_logic ;
         q_arr_12_0 : IN std_logic ;
         q_arr_13_31 : IN std_logic ;
         q_arr_13_30 : IN std_logic ;
         q_arr_13_29 : IN std_logic ;
         q_arr_13_28 : IN std_logic ;
         q_arr_13_27 : IN std_logic ;
         q_arr_13_26 : IN std_logic ;
         q_arr_13_25 : IN std_logic ;
         q_arr_13_24 : IN std_logic ;
         q_arr_13_23 : IN std_logic ;
         q_arr_13_22 : IN std_logic ;
         q_arr_13_21 : IN std_logic ;
         q_arr_13_20 : IN std_logic ;
         q_arr_13_19 : IN std_logic ;
         q_arr_13_18 : IN std_logic ;
         q_arr_13_17 : IN std_logic ;
         q_arr_13_16 : IN std_logic ;
         q_arr_13_15 : IN std_logic ;
         q_arr_13_14 : IN std_logic ;
         q_arr_13_13 : IN std_logic ;
         q_arr_13_12 : IN std_logic ;
         q_arr_13_11 : IN std_logic ;
         q_arr_13_10 : IN std_logic ;
         q_arr_13_9 : IN std_logic ;
         q_arr_13_8 : IN std_logic ;
         q_arr_13_7 : IN std_logic ;
         q_arr_13_6 : IN std_logic ;
         q_arr_13_5 : IN std_logic ;
         q_arr_13_4 : IN std_logic ;
         q_arr_13_3 : IN std_logic ;
         q_arr_13_2 : IN std_logic ;
         q_arr_13_1 : IN std_logic ;
         q_arr_13_0 : IN std_logic ;
         q_arr_14_31 : IN std_logic ;
         q_arr_14_30 : IN std_logic ;
         q_arr_14_29 : IN std_logic ;
         q_arr_14_28 : IN std_logic ;
         q_arr_14_27 : IN std_logic ;
         q_arr_14_26 : IN std_logic ;
         q_arr_14_25 : IN std_logic ;
         q_arr_14_24 : IN std_logic ;
         q_arr_14_23 : IN std_logic ;
         q_arr_14_22 : IN std_logic ;
         q_arr_14_21 : IN std_logic ;
         q_arr_14_20 : IN std_logic ;
         q_arr_14_19 : IN std_logic ;
         q_arr_14_18 : IN std_logic ;
         q_arr_14_17 : IN std_logic ;
         q_arr_14_16 : IN std_logic ;
         q_arr_14_15 : IN std_logic ;
         q_arr_14_14 : IN std_logic ;
         q_arr_14_13 : IN std_logic ;
         q_arr_14_12 : IN std_logic ;
         q_arr_14_11 : IN std_logic ;
         q_arr_14_10 : IN std_logic ;
         q_arr_14_9 : IN std_logic ;
         q_arr_14_8 : IN std_logic ;
         q_arr_14_7 : IN std_logic ;
         q_arr_14_6 : IN std_logic ;
         q_arr_14_5 : IN std_logic ;
         q_arr_14_4 : IN std_logic ;
         q_arr_14_3 : IN std_logic ;
         q_arr_14_2 : IN std_logic ;
         q_arr_14_1 : IN std_logic ;
         q_arr_14_0 : IN std_logic ;
         q_arr_15_31 : IN std_logic ;
         q_arr_15_30 : IN std_logic ;
         q_arr_15_29 : IN std_logic ;
         q_arr_15_28 : IN std_logic ;
         q_arr_15_27 : IN std_logic ;
         q_arr_15_26 : IN std_logic ;
         q_arr_15_25 : IN std_logic ;
         q_arr_15_24 : IN std_logic ;
         q_arr_15_23 : IN std_logic ;
         q_arr_15_22 : IN std_logic ;
         q_arr_15_21 : IN std_logic ;
         q_arr_15_20 : IN std_logic ;
         q_arr_15_19 : IN std_logic ;
         q_arr_15_18 : IN std_logic ;
         q_arr_15_17 : IN std_logic ;
         q_arr_15_16 : IN std_logic ;
         q_arr_15_15 : IN std_logic ;
         q_arr_15_14 : IN std_logic ;
         q_arr_15_13 : IN std_logic ;
         q_arr_15_12 : IN std_logic ;
         q_arr_15_11 : IN std_logic ;
         q_arr_15_10 : IN std_logic ;
         q_arr_15_9 : IN std_logic ;
         q_arr_15_8 : IN std_logic ;
         q_arr_15_7 : IN std_logic ;
         q_arr_15_6 : IN std_logic ;
         q_arr_15_5 : IN std_logic ;
         q_arr_15_4 : IN std_logic ;
         q_arr_15_3 : IN std_logic ;
         q_arr_15_2 : IN std_logic ;
         q_arr_15_1 : IN std_logic ;
         q_arr_15_0 : IN std_logic ;
         q_arr_16_31 : IN std_logic ;
         q_arr_16_30 : IN std_logic ;
         q_arr_16_29 : IN std_logic ;
         q_arr_16_28 : IN std_logic ;
         q_arr_16_27 : IN std_logic ;
         q_arr_16_26 : IN std_logic ;
         q_arr_16_25 : IN std_logic ;
         q_arr_16_24 : IN std_logic ;
         q_arr_16_23 : IN std_logic ;
         q_arr_16_22 : IN std_logic ;
         q_arr_16_21 : IN std_logic ;
         q_arr_16_20 : IN std_logic ;
         q_arr_16_19 : IN std_logic ;
         q_arr_16_18 : IN std_logic ;
         q_arr_16_17 : IN std_logic ;
         q_arr_16_16 : IN std_logic ;
         q_arr_16_15 : IN std_logic ;
         q_arr_16_14 : IN std_logic ;
         q_arr_16_13 : IN std_logic ;
         q_arr_16_12 : IN std_logic ;
         q_arr_16_11 : IN std_logic ;
         q_arr_16_10 : IN std_logic ;
         q_arr_16_9 : IN std_logic ;
         q_arr_16_8 : IN std_logic ;
         q_arr_16_7 : IN std_logic ;
         q_arr_16_6 : IN std_logic ;
         q_arr_16_5 : IN std_logic ;
         q_arr_16_4 : IN std_logic ;
         q_arr_16_3 : IN std_logic ;
         q_arr_16_2 : IN std_logic ;
         q_arr_16_1 : IN std_logic ;
         q_arr_16_0 : IN std_logic ;
         q_arr_17_31 : IN std_logic ;
         q_arr_17_30 : IN std_logic ;
         q_arr_17_29 : IN std_logic ;
         q_arr_17_28 : IN std_logic ;
         q_arr_17_27 : IN std_logic ;
         q_arr_17_26 : IN std_logic ;
         q_arr_17_25 : IN std_logic ;
         q_arr_17_24 : IN std_logic ;
         q_arr_17_23 : IN std_logic ;
         q_arr_17_22 : IN std_logic ;
         q_arr_17_21 : IN std_logic ;
         q_arr_17_20 : IN std_logic ;
         q_arr_17_19 : IN std_logic ;
         q_arr_17_18 : IN std_logic ;
         q_arr_17_17 : IN std_logic ;
         q_arr_17_16 : IN std_logic ;
         q_arr_17_15 : IN std_logic ;
         q_arr_17_14 : IN std_logic ;
         q_arr_17_13 : IN std_logic ;
         q_arr_17_12 : IN std_logic ;
         q_arr_17_11 : IN std_logic ;
         q_arr_17_10 : IN std_logic ;
         q_arr_17_9 : IN std_logic ;
         q_arr_17_8 : IN std_logic ;
         q_arr_17_7 : IN std_logic ;
         q_arr_17_6 : IN std_logic ;
         q_arr_17_5 : IN std_logic ;
         q_arr_17_4 : IN std_logic ;
         q_arr_17_3 : IN std_logic ;
         q_arr_17_2 : IN std_logic ;
         q_arr_17_1 : IN std_logic ;
         q_arr_17_0 : IN std_logic ;
         q_arr_18_31 : IN std_logic ;
         q_arr_18_30 : IN std_logic ;
         q_arr_18_29 : IN std_logic ;
         q_arr_18_28 : IN std_logic ;
         q_arr_18_27 : IN std_logic ;
         q_arr_18_26 : IN std_logic ;
         q_arr_18_25 : IN std_logic ;
         q_arr_18_24 : IN std_logic ;
         q_arr_18_23 : IN std_logic ;
         q_arr_18_22 : IN std_logic ;
         q_arr_18_21 : IN std_logic ;
         q_arr_18_20 : IN std_logic ;
         q_arr_18_19 : IN std_logic ;
         q_arr_18_18 : IN std_logic ;
         q_arr_18_17 : IN std_logic ;
         q_arr_18_16 : IN std_logic ;
         q_arr_18_15 : IN std_logic ;
         q_arr_18_14 : IN std_logic ;
         q_arr_18_13 : IN std_logic ;
         q_arr_18_12 : IN std_logic ;
         q_arr_18_11 : IN std_logic ;
         q_arr_18_10 : IN std_logic ;
         q_arr_18_9 : IN std_logic ;
         q_arr_18_8 : IN std_logic ;
         q_arr_18_7 : IN std_logic ;
         q_arr_18_6 : IN std_logic ;
         q_arr_18_5 : IN std_logic ;
         q_arr_18_4 : IN std_logic ;
         q_arr_18_3 : IN std_logic ;
         q_arr_18_2 : IN std_logic ;
         q_arr_18_1 : IN std_logic ;
         q_arr_18_0 : IN std_logic ;
         q_arr_19_31 : IN std_logic ;
         q_arr_19_30 : IN std_logic ;
         q_arr_19_29 : IN std_logic ;
         q_arr_19_28 : IN std_logic ;
         q_arr_19_27 : IN std_logic ;
         q_arr_19_26 : IN std_logic ;
         q_arr_19_25 : IN std_logic ;
         q_arr_19_24 : IN std_logic ;
         q_arr_19_23 : IN std_logic ;
         q_arr_19_22 : IN std_logic ;
         q_arr_19_21 : IN std_logic ;
         q_arr_19_20 : IN std_logic ;
         q_arr_19_19 : IN std_logic ;
         q_arr_19_18 : IN std_logic ;
         q_arr_19_17 : IN std_logic ;
         q_arr_19_16 : IN std_logic ;
         q_arr_19_15 : IN std_logic ;
         q_arr_19_14 : IN std_logic ;
         q_arr_19_13 : IN std_logic ;
         q_arr_19_12 : IN std_logic ;
         q_arr_19_11 : IN std_logic ;
         q_arr_19_10 : IN std_logic ;
         q_arr_19_9 : IN std_logic ;
         q_arr_19_8 : IN std_logic ;
         q_arr_19_7 : IN std_logic ;
         q_arr_19_6 : IN std_logic ;
         q_arr_19_5 : IN std_logic ;
         q_arr_19_4 : IN std_logic ;
         q_arr_19_3 : IN std_logic ;
         q_arr_19_2 : IN std_logic ;
         q_arr_19_1 : IN std_logic ;
         q_arr_19_0 : IN std_logic ;
         q_arr_20_31 : IN std_logic ;
         q_arr_20_30 : IN std_logic ;
         q_arr_20_29 : IN std_logic ;
         q_arr_20_28 : IN std_logic ;
         q_arr_20_27 : IN std_logic ;
         q_arr_20_26 : IN std_logic ;
         q_arr_20_25 : IN std_logic ;
         q_arr_20_24 : IN std_logic ;
         q_arr_20_23 : IN std_logic ;
         q_arr_20_22 : IN std_logic ;
         q_arr_20_21 : IN std_logic ;
         q_arr_20_20 : IN std_logic ;
         q_arr_20_19 : IN std_logic ;
         q_arr_20_18 : IN std_logic ;
         q_arr_20_17 : IN std_logic ;
         q_arr_20_16 : IN std_logic ;
         q_arr_20_15 : IN std_logic ;
         q_arr_20_14 : IN std_logic ;
         q_arr_20_13 : IN std_logic ;
         q_arr_20_12 : IN std_logic ;
         q_arr_20_11 : IN std_logic ;
         q_arr_20_10 : IN std_logic ;
         q_arr_20_9 : IN std_logic ;
         q_arr_20_8 : IN std_logic ;
         q_arr_20_7 : IN std_logic ;
         q_arr_20_6 : IN std_logic ;
         q_arr_20_5 : IN std_logic ;
         q_arr_20_4 : IN std_logic ;
         q_arr_20_3 : IN std_logic ;
         q_arr_20_2 : IN std_logic ;
         q_arr_20_1 : IN std_logic ;
         q_arr_20_0 : IN std_logic ;
         q_arr_21_31 : IN std_logic ;
         q_arr_21_30 : IN std_logic ;
         q_arr_21_29 : IN std_logic ;
         q_arr_21_28 : IN std_logic ;
         q_arr_21_27 : IN std_logic ;
         q_arr_21_26 : IN std_logic ;
         q_arr_21_25 : IN std_logic ;
         q_arr_21_24 : IN std_logic ;
         q_arr_21_23 : IN std_logic ;
         q_arr_21_22 : IN std_logic ;
         q_arr_21_21 : IN std_logic ;
         q_arr_21_20 : IN std_logic ;
         q_arr_21_19 : IN std_logic ;
         q_arr_21_18 : IN std_logic ;
         q_arr_21_17 : IN std_logic ;
         q_arr_21_16 : IN std_logic ;
         q_arr_21_15 : IN std_logic ;
         q_arr_21_14 : IN std_logic ;
         q_arr_21_13 : IN std_logic ;
         q_arr_21_12 : IN std_logic ;
         q_arr_21_11 : IN std_logic ;
         q_arr_21_10 : IN std_logic ;
         q_arr_21_9 : IN std_logic ;
         q_arr_21_8 : IN std_logic ;
         q_arr_21_7 : IN std_logic ;
         q_arr_21_6 : IN std_logic ;
         q_arr_21_5 : IN std_logic ;
         q_arr_21_4 : IN std_logic ;
         q_arr_21_3 : IN std_logic ;
         q_arr_21_2 : IN std_logic ;
         q_arr_21_1 : IN std_logic ;
         q_arr_21_0 : IN std_logic ;
         q_arr_22_31 : IN std_logic ;
         q_arr_22_30 : IN std_logic ;
         q_arr_22_29 : IN std_logic ;
         q_arr_22_28 : IN std_logic ;
         q_arr_22_27 : IN std_logic ;
         q_arr_22_26 : IN std_logic ;
         q_arr_22_25 : IN std_logic ;
         q_arr_22_24 : IN std_logic ;
         q_arr_22_23 : IN std_logic ;
         q_arr_22_22 : IN std_logic ;
         q_arr_22_21 : IN std_logic ;
         q_arr_22_20 : IN std_logic ;
         q_arr_22_19 : IN std_logic ;
         q_arr_22_18 : IN std_logic ;
         q_arr_22_17 : IN std_logic ;
         q_arr_22_16 : IN std_logic ;
         q_arr_22_15 : IN std_logic ;
         q_arr_22_14 : IN std_logic ;
         q_arr_22_13 : IN std_logic ;
         q_arr_22_12 : IN std_logic ;
         q_arr_22_11 : IN std_logic ;
         q_arr_22_10 : IN std_logic ;
         q_arr_22_9 : IN std_logic ;
         q_arr_22_8 : IN std_logic ;
         q_arr_22_7 : IN std_logic ;
         q_arr_22_6 : IN std_logic ;
         q_arr_22_5 : IN std_logic ;
         q_arr_22_4 : IN std_logic ;
         q_arr_22_3 : IN std_logic ;
         q_arr_22_2 : IN std_logic ;
         q_arr_22_1 : IN std_logic ;
         q_arr_22_0 : IN std_logic ;
         q_arr_23_31 : IN std_logic ;
         q_arr_23_30 : IN std_logic ;
         q_arr_23_29 : IN std_logic ;
         q_arr_23_28 : IN std_logic ;
         q_arr_23_27 : IN std_logic ;
         q_arr_23_26 : IN std_logic ;
         q_arr_23_25 : IN std_logic ;
         q_arr_23_24 : IN std_logic ;
         q_arr_23_23 : IN std_logic ;
         q_arr_23_22 : IN std_logic ;
         q_arr_23_21 : IN std_logic ;
         q_arr_23_20 : IN std_logic ;
         q_arr_23_19 : IN std_logic ;
         q_arr_23_18 : IN std_logic ;
         q_arr_23_17 : IN std_logic ;
         q_arr_23_16 : IN std_logic ;
         q_arr_23_15 : IN std_logic ;
         q_arr_23_14 : IN std_logic ;
         q_arr_23_13 : IN std_logic ;
         q_arr_23_12 : IN std_logic ;
         q_arr_23_11 : IN std_logic ;
         q_arr_23_10 : IN std_logic ;
         q_arr_23_9 : IN std_logic ;
         q_arr_23_8 : IN std_logic ;
         q_arr_23_7 : IN std_logic ;
         q_arr_23_6 : IN std_logic ;
         q_arr_23_5 : IN std_logic ;
         q_arr_23_4 : IN std_logic ;
         q_arr_23_3 : IN std_logic ;
         q_arr_23_2 : IN std_logic ;
         q_arr_23_1 : IN std_logic ;
         q_arr_23_0 : IN std_logic ;
         q_arr_24_31 : IN std_logic ;
         q_arr_24_30 : IN std_logic ;
         q_arr_24_29 : IN std_logic ;
         q_arr_24_28 : IN std_logic ;
         q_arr_24_27 : IN std_logic ;
         q_arr_24_26 : IN std_logic ;
         q_arr_24_25 : IN std_logic ;
         q_arr_24_24 : IN std_logic ;
         q_arr_24_23 : IN std_logic ;
         q_arr_24_22 : IN std_logic ;
         q_arr_24_21 : IN std_logic ;
         q_arr_24_20 : IN std_logic ;
         q_arr_24_19 : IN std_logic ;
         q_arr_24_18 : IN std_logic ;
         q_arr_24_17 : IN std_logic ;
         q_arr_24_16 : IN std_logic ;
         q_arr_24_15 : IN std_logic ;
         q_arr_24_14 : IN std_logic ;
         q_arr_24_13 : IN std_logic ;
         q_arr_24_12 : IN std_logic ;
         q_arr_24_11 : IN std_logic ;
         q_arr_24_10 : IN std_logic ;
         q_arr_24_9 : IN std_logic ;
         q_arr_24_8 : IN std_logic ;
         q_arr_24_7 : IN std_logic ;
         q_arr_24_6 : IN std_logic ;
         q_arr_24_5 : IN std_logic ;
         q_arr_24_4 : IN std_logic ;
         q_arr_24_3 : IN std_logic ;
         q_arr_24_2 : IN std_logic ;
         q_arr_24_1 : IN std_logic ;
         q_arr_24_0 : IN std_logic) ;
   end component ;
   component ModifiedBoothMultiplier
      port (
         M : IN std_logic_vector (15 DOWNTO 0) ;
         R : IN std_logic_vector (15 DOWNTO 0) ;
         cnt_enable : IN std_logic ;
         product : OUT std_logic_vector (31 DOWNTO 0) ;
         clk : IN std_logic) ;
   end component ;
   component NAdder_32
      port (
         a : IN std_logic_vector (31 DOWNTO 0) ;
         b : IN std_logic_vector (31 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (31 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   component NAdder_32_unfolded0
      port (
         a : IN std_logic_vector (31 DOWNTO 0) ;
         b : IN std_logic_vector (31 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (31 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal buffer_ready_EXMPLR, semi_ready_EXMPLR, counter_15, counter_14, 
      counter_13, counter_0, ordered_filter_data_3_15, 
      ordered_filter_data_3_14, ordered_filter_data_3_13, 
      ordered_filter_data_3_12, ordered_filter_data_3_11, 
      ordered_filter_data_3_10, ordered_filter_data_3_9, 
      ordered_filter_data_3_8, ordered_filter_data_3_7, 
      ordered_filter_data_3_6, ordered_filter_data_3_5, 
      ordered_filter_data_3_4, ordered_filter_data_3_3, 
      ordered_filter_data_3_2, ordered_filter_data_3_1, 
      ordered_filter_data_3_0, ordered_filter_data_4_15, 
      ordered_filter_data_4_14, ordered_filter_data_4_13, 
      ordered_filter_data_4_12, ordered_filter_data_4_11, 
      ordered_filter_data_4_10, ordered_filter_data_4_9, 
      ordered_filter_data_4_8, ordered_filter_data_4_7, 
      ordered_filter_data_4_6, ordered_filter_data_4_5, 
      ordered_filter_data_4_4, ordered_filter_data_4_3, 
      ordered_filter_data_4_2, ordered_filter_data_4_1, 
      ordered_filter_data_4_0, ordered_filter_data_5_15, 
      ordered_filter_data_5_14, ordered_filter_data_5_13, 
      ordered_filter_data_5_12, ordered_filter_data_5_11, 
      ordered_filter_data_5_10, ordered_filter_data_5_9, 
      ordered_filter_data_5_8, ordered_filter_data_5_7, 
      ordered_filter_data_5_6, ordered_filter_data_5_5, 
      ordered_filter_data_5_4, ordered_filter_data_5_3, 
      ordered_filter_data_5_2, ordered_filter_data_5_1, 
      ordered_filter_data_5_0, ordered_filter_data_6_15, 
      ordered_filter_data_6_14, ordered_filter_data_6_13, 
      ordered_filter_data_6_12, ordered_filter_data_6_11, 
      ordered_filter_data_6_10, ordered_filter_data_6_9, 
      ordered_filter_data_6_8, ordered_filter_data_6_7, 
      ordered_filter_data_6_6, ordered_filter_data_6_5, 
      ordered_filter_data_6_4, ordered_filter_data_6_3, 
      ordered_filter_data_6_2, ordered_filter_data_6_1, 
      ordered_filter_data_6_0, ordered_filter_data_7_15, 
      ordered_filter_data_7_14, ordered_filter_data_7_13, 
      ordered_filter_data_7_12, ordered_filter_data_7_11, 
      ordered_filter_data_7_10, ordered_filter_data_7_9, 
      ordered_filter_data_7_8, ordered_filter_data_7_7, 
      ordered_filter_data_7_6, ordered_filter_data_7_5, 
      ordered_filter_data_7_4, ordered_filter_data_7_3, 
      ordered_filter_data_7_2, ordered_filter_data_7_1, 
      ordered_filter_data_7_0, ordered_filter_data_8_15, 
      ordered_filter_data_8_14, ordered_filter_data_8_13, 
      ordered_filter_data_8_12, ordered_filter_data_8_11, 
      ordered_filter_data_8_10, ordered_filter_data_8_9, 
      ordered_filter_data_8_8, ordered_filter_data_8_7, 
      ordered_filter_data_8_6, ordered_filter_data_8_5, 
      ordered_filter_data_8_4, ordered_filter_data_8_3, 
      ordered_filter_data_8_2, ordered_filter_data_8_1, 
      ordered_filter_data_8_0, ordered_filter_data_9_15, 
      ordered_filter_data_9_14, ordered_filter_data_9_13, 
      ordered_filter_data_9_12, ordered_filter_data_9_11, 
      ordered_filter_data_9_10, ordered_filter_data_9_9, 
      ordered_filter_data_9_8, ordered_filter_data_9_7, 
      ordered_filter_data_9_6, ordered_filter_data_9_5, 
      ordered_filter_data_9_4, ordered_filter_data_9_3, 
      ordered_filter_data_9_2, ordered_filter_data_9_1, 
      ordered_filter_data_9_0, ordered_filter_data_10_15, 
      ordered_filter_data_10_14, ordered_filter_data_10_13, 
      ordered_filter_data_10_12, ordered_filter_data_10_11, 
      ordered_filter_data_10_10, ordered_filter_data_10_9, 
      ordered_filter_data_10_8, ordered_filter_data_10_7, 
      ordered_filter_data_10_6, ordered_filter_data_10_5, 
      ordered_filter_data_10_4, ordered_filter_data_10_3, 
      ordered_filter_data_10_2, ordered_filter_data_10_1, 
      ordered_filter_data_10_0, ordered_filter_data_11_15, 
      ordered_filter_data_11_14, ordered_filter_data_11_13, 
      ordered_filter_data_11_12, ordered_filter_data_11_11, 
      ordered_filter_data_11_10, ordered_filter_data_11_9, 
      ordered_filter_data_11_8, ordered_filter_data_11_7, 
      ordered_filter_data_11_6, ordered_filter_data_11_5, 
      ordered_filter_data_11_4, ordered_filter_data_11_3, 
      ordered_filter_data_11_2, ordered_filter_data_11_1, 
      ordered_filter_data_11_0, ordered_filter_data_12_15, 
      ordered_filter_data_12_14, ordered_filter_data_12_13, 
      ordered_filter_data_12_12, ordered_filter_data_12_11, 
      ordered_filter_data_12_10, ordered_filter_data_12_9, 
      ordered_filter_data_12_8, ordered_filter_data_12_7, 
      ordered_filter_data_12_6, ordered_filter_data_12_5, 
      ordered_filter_data_12_4, ordered_filter_data_12_3, 
      ordered_filter_data_12_2, ordered_filter_data_12_1, 
      ordered_filter_data_12_0, ordered_filter_data_13_15, 
      ordered_filter_data_13_14, ordered_filter_data_13_13, 
      ordered_filter_data_13_12, ordered_filter_data_13_11, 
      ordered_filter_data_13_10, ordered_filter_data_13_9, 
      ordered_filter_data_13_8, ordered_filter_data_13_7, 
      ordered_filter_data_13_6, ordered_filter_data_13_5, 
      ordered_filter_data_13_4, ordered_filter_data_13_3, 
      ordered_filter_data_13_2, ordered_filter_data_13_1, 
      ordered_filter_data_13_0, ordered_filter_data_14_15, 
      ordered_filter_data_14_14, ordered_filter_data_14_13, 
      ordered_filter_data_14_12, ordered_filter_data_14_11, 
      ordered_filter_data_14_10, ordered_filter_data_14_9, 
      ordered_filter_data_14_8, ordered_filter_data_14_7, 
      ordered_filter_data_14_6, ordered_filter_data_14_5, 
      ordered_filter_data_14_4, ordered_filter_data_14_3, 
      ordered_filter_data_14_2, ordered_filter_data_14_1, 
      ordered_filter_data_14_0, ordered_filter_data_15_15, 
      ordered_filter_data_15_14, ordered_filter_data_15_13, 
      ordered_filter_data_15_12, ordered_filter_data_15_11, 
      ordered_filter_data_15_10, ordered_filter_data_15_9, 
      ordered_filter_data_15_8, ordered_filter_data_15_7, 
      ordered_filter_data_15_6, ordered_filter_data_15_5, 
      ordered_filter_data_15_4, ordered_filter_data_15_3, 
      ordered_filter_data_15_2, ordered_filter_data_15_1, 
      ordered_filter_data_15_0, ordered_filter_data_16_15, 
      ordered_filter_data_16_14, ordered_filter_data_16_13, 
      ordered_filter_data_16_12, ordered_filter_data_16_11, 
      ordered_filter_data_16_10, ordered_filter_data_16_9, 
      ordered_filter_data_16_8, ordered_filter_data_16_7, 
      ordered_filter_data_16_6, ordered_filter_data_16_5, 
      ordered_filter_data_16_4, ordered_filter_data_16_3, 
      ordered_filter_data_16_2, ordered_filter_data_16_1, 
      ordered_filter_data_16_0, ordered_filter_data_17_15, 
      ordered_filter_data_17_14, ordered_filter_data_17_13, 
      ordered_filter_data_17_12, ordered_filter_data_17_11, 
      ordered_filter_data_17_10, ordered_filter_data_17_9, 
      ordered_filter_data_17_8, ordered_filter_data_17_7, 
      ordered_filter_data_17_6, ordered_filter_data_17_5, 
      ordered_filter_data_17_4, ordered_filter_data_17_3, 
      ordered_filter_data_17_2, ordered_filter_data_17_1, 
      ordered_filter_data_17_0, ordered_img_data_9_31, ordered_img_data_9_14, 
      ordered_img_data_9_13, ordered_img_data_9_12, ordered_img_data_9_11, 
      ordered_img_data_9_10, ordered_img_data_9_9, ordered_img_data_9_8, 
      ordered_img_data_9_7, ordered_img_data_9_6, ordered_img_data_9_5, 
      ordered_img_data_9_4, ordered_img_data_9_3, ordered_img_data_9_2, 
      ordered_img_data_9_1, ordered_img_data_9_0, ordered_img_data_10_31, 
      ordered_img_data_10_14, ordered_img_data_10_13, ordered_img_data_10_12, 
      ordered_img_data_10_11, ordered_img_data_10_10, ordered_img_data_10_9, 
      ordered_img_data_10_8, ordered_img_data_10_7, ordered_img_data_10_6, 
      ordered_img_data_10_5, ordered_img_data_10_4, ordered_img_data_10_3, 
      ordered_img_data_10_2, ordered_img_data_10_1, ordered_img_data_10_0, 
      ordered_img_data_11_31, ordered_img_data_11_14, ordered_img_data_11_13, 
      ordered_img_data_11_12, ordered_img_data_11_11, ordered_img_data_11_10, 
      ordered_img_data_11_9, ordered_img_data_11_8, ordered_img_data_11_7, 
      ordered_img_data_11_6, ordered_img_data_11_5, ordered_img_data_11_4, 
      ordered_img_data_11_3, ordered_img_data_11_2, ordered_img_data_11_1, 
      ordered_img_data_11_0, ordered_img_data_12_31, ordered_img_data_12_14, 
      ordered_img_data_12_13, ordered_img_data_12_12, ordered_img_data_12_11, 
      ordered_img_data_12_10, ordered_img_data_12_9, ordered_img_data_12_8, 
      ordered_img_data_12_7, ordered_img_data_12_6, ordered_img_data_12_5, 
      ordered_img_data_12_4, ordered_img_data_12_3, ordered_img_data_12_2, 
      ordered_img_data_12_1, ordered_img_data_12_0, ordered_img_data_13_31, 
      ordered_img_data_13_14, ordered_img_data_13_13, ordered_img_data_13_12, 
      ordered_img_data_13_11, ordered_img_data_13_10, ordered_img_data_13_9, 
      ordered_img_data_13_8, ordered_img_data_13_7, ordered_img_data_13_6, 
      ordered_img_data_13_5, ordered_img_data_13_4, ordered_img_data_13_3, 
      ordered_img_data_13_2, ordered_img_data_13_1, ordered_img_data_13_0, 
      ordered_img_data_14_31, ordered_img_data_14_14, ordered_img_data_14_13, 
      ordered_img_data_14_12, ordered_img_data_14_11, ordered_img_data_14_10, 
      ordered_img_data_14_9, ordered_img_data_14_8, ordered_img_data_14_7, 
      ordered_img_data_14_6, ordered_img_data_14_5, ordered_img_data_14_4, 
      ordered_img_data_14_3, ordered_img_data_14_2, ordered_img_data_14_1, 
      ordered_img_data_14_0, ordered_img_data_15_31, ordered_img_data_15_14, 
      ordered_img_data_15_13, ordered_img_data_15_12, ordered_img_data_15_11, 
      ordered_img_data_15_10, ordered_img_data_15_9, ordered_img_data_15_8, 
      ordered_img_data_15_7, ordered_img_data_15_6, ordered_img_data_15_5, 
      ordered_img_data_15_4, ordered_img_data_15_3, ordered_img_data_15_2, 
      ordered_img_data_15_1, ordered_img_data_15_0, ordered_img_data_16_31, 
      ordered_img_data_16_14, ordered_img_data_16_13, ordered_img_data_16_12, 
      ordered_img_data_16_11, ordered_img_data_16_10, ordered_img_data_16_9, 
      ordered_img_data_16_8, ordered_img_data_16_7, ordered_img_data_16_6, 
      ordered_img_data_16_5, ordered_img_data_16_4, ordered_img_data_16_3, 
      ordered_img_data_16_2, ordered_img_data_16_1, ordered_img_data_16_0, 
      ordered_img_data_17_31, ordered_img_data_17_14, ordered_img_data_17_13, 
      ordered_img_data_17_12, ordered_img_data_17_11, ordered_img_data_17_10, 
      ordered_img_data_17_9, ordered_img_data_17_8, ordered_img_data_17_7, 
      ordered_img_data_17_6, ordered_img_data_17_5, ordered_img_data_17_4, 
      ordered_img_data_17_3, ordered_img_data_17_2, ordered_img_data_17_1, 
      ordered_img_data_17_0, d_arr_mul_0_31, d_arr_mul_0_30, d_arr_mul_0_29, 
      d_arr_mul_0_28, d_arr_mul_0_27, d_arr_mul_0_26, d_arr_mul_0_25, 
      d_arr_mul_0_24, d_arr_mul_0_23, d_arr_mul_0_22, d_arr_mul_0_21, 
      d_arr_mul_0_20, d_arr_mul_0_19, d_arr_mul_0_18, d_arr_mul_0_17, 
      d_arr_mul_0_16, d_arr_mul_0_15, d_arr_mul_0_14, d_arr_mul_0_13, 
      d_arr_mul_0_12, d_arr_mul_0_11, d_arr_mul_0_10, d_arr_mul_0_9, 
      d_arr_mul_0_8, d_arr_mul_0_7, d_arr_mul_0_6, d_arr_mul_0_5, 
      d_arr_mul_0_4, d_arr_mul_0_3, d_arr_mul_0_2, d_arr_mul_0_1, 
      d_arr_mul_0_0, d_arr_mul_1_31, d_arr_mul_1_30, d_arr_mul_1_29, 
      d_arr_mul_1_28, d_arr_mul_1_27, d_arr_mul_1_26, d_arr_mul_1_25, 
      d_arr_mul_1_24, d_arr_mul_1_23, d_arr_mul_1_22, d_arr_mul_1_21, 
      d_arr_mul_1_20, d_arr_mul_1_19, d_arr_mul_1_18, d_arr_mul_1_17, 
      d_arr_mul_1_16, d_arr_mul_1_15, d_arr_mul_1_14, d_arr_mul_1_13, 
      d_arr_mul_1_12, d_arr_mul_1_11, d_arr_mul_1_10, d_arr_mul_1_9, 
      d_arr_mul_1_8, d_arr_mul_1_7, d_arr_mul_1_6, d_arr_mul_1_5, 
      d_arr_mul_1_4, d_arr_mul_1_3, d_arr_mul_1_2, d_arr_mul_1_1, 
      d_arr_mul_1_0, d_arr_mul_2_31, d_arr_mul_2_30, d_arr_mul_2_29, 
      d_arr_mul_2_28, d_arr_mul_2_27, d_arr_mul_2_26, d_arr_mul_2_25, 
      d_arr_mul_2_24, d_arr_mul_2_23, d_arr_mul_2_22, d_arr_mul_2_21, 
      d_arr_mul_2_20, d_arr_mul_2_19, d_arr_mul_2_18, d_arr_mul_2_17, 
      d_arr_mul_2_16, d_arr_mul_2_15, d_arr_mul_2_14, d_arr_mul_2_13, 
      d_arr_mul_2_12, d_arr_mul_2_11, d_arr_mul_2_10, d_arr_mul_2_9, 
      d_arr_mul_2_8, d_arr_mul_2_7, d_arr_mul_2_6, d_arr_mul_2_5, 
      d_arr_mul_2_4, d_arr_mul_2_3, d_arr_mul_2_2, d_arr_mul_2_1, 
      d_arr_mul_2_0, d_arr_mul_3_31, d_arr_mul_3_30, d_arr_mul_3_29, 
      d_arr_mul_3_28, d_arr_mul_3_27, d_arr_mul_3_26, d_arr_mul_3_25, 
      d_arr_mul_3_24, d_arr_mul_3_23, d_arr_mul_3_22, d_arr_mul_3_21, 
      d_arr_mul_3_20, d_arr_mul_3_19, d_arr_mul_3_18, d_arr_mul_3_17, 
      d_arr_mul_3_16, d_arr_mul_3_15, d_arr_mul_3_14, d_arr_mul_3_13, 
      d_arr_mul_3_12, d_arr_mul_3_11, d_arr_mul_3_10, d_arr_mul_3_9, 
      d_arr_mul_3_8, d_arr_mul_3_7, d_arr_mul_3_6, d_arr_mul_3_5, 
      d_arr_mul_3_4, d_arr_mul_3_3, d_arr_mul_3_2, d_arr_mul_3_1, 
      d_arr_mul_3_0, d_arr_mul_4_31, d_arr_mul_4_30, d_arr_mul_4_29, 
      d_arr_mul_4_28, d_arr_mul_4_27, d_arr_mul_4_26, d_arr_mul_4_25, 
      d_arr_mul_4_24, d_arr_mul_4_23, d_arr_mul_4_22, d_arr_mul_4_21, 
      d_arr_mul_4_20, d_arr_mul_4_19, d_arr_mul_4_18, d_arr_mul_4_17, 
      d_arr_mul_4_16, d_arr_mul_4_15, d_arr_mul_4_14, d_arr_mul_4_13, 
      d_arr_mul_4_12, d_arr_mul_4_11, d_arr_mul_4_10, d_arr_mul_4_9, 
      d_arr_mul_4_8, d_arr_mul_4_7, d_arr_mul_4_6, d_arr_mul_4_5, 
      d_arr_mul_4_4, d_arr_mul_4_3, d_arr_mul_4_2, d_arr_mul_4_1, 
      d_arr_mul_4_0, d_arr_mul_5_31, d_arr_mul_5_30, d_arr_mul_5_29, 
      d_arr_mul_5_28, d_arr_mul_5_27, d_arr_mul_5_26, d_arr_mul_5_25, 
      d_arr_mul_5_24, d_arr_mul_5_23, d_arr_mul_5_22, d_arr_mul_5_21, 
      d_arr_mul_5_20, d_arr_mul_5_19, d_arr_mul_5_18, d_arr_mul_5_17, 
      d_arr_mul_5_16, d_arr_mul_5_15, d_arr_mul_5_14, d_arr_mul_5_13, 
      d_arr_mul_5_12, d_arr_mul_5_11, d_arr_mul_5_10, d_arr_mul_5_9, 
      d_arr_mul_5_8, d_arr_mul_5_7, d_arr_mul_5_6, d_arr_mul_5_5, 
      d_arr_mul_5_4, d_arr_mul_5_3, d_arr_mul_5_2, d_arr_mul_5_1, 
      d_arr_mul_5_0, d_arr_mul_6_31, d_arr_mul_6_30, d_arr_mul_6_29, 
      d_arr_mul_6_28, d_arr_mul_6_27, d_arr_mul_6_26, d_arr_mul_6_25, 
      d_arr_mul_6_24, d_arr_mul_6_23, d_arr_mul_6_22, d_arr_mul_6_21, 
      d_arr_mul_6_20, d_arr_mul_6_19, d_arr_mul_6_18, d_arr_mul_6_17, 
      d_arr_mul_6_16, d_arr_mul_6_15, d_arr_mul_6_14, d_arr_mul_6_13, 
      d_arr_mul_6_12, d_arr_mul_6_11, d_arr_mul_6_10, d_arr_mul_6_9, 
      d_arr_mul_6_8, d_arr_mul_6_7, d_arr_mul_6_6, d_arr_mul_6_5, 
      d_arr_mul_6_4, d_arr_mul_6_3, d_arr_mul_6_2, d_arr_mul_6_1, 
      d_arr_mul_6_0, d_arr_mul_7_31, d_arr_mul_7_30, d_arr_mul_7_29, 
      d_arr_mul_7_28, d_arr_mul_7_27, d_arr_mul_7_26, d_arr_mul_7_25, 
      d_arr_mul_7_24, d_arr_mul_7_23, d_arr_mul_7_22, d_arr_mul_7_21, 
      d_arr_mul_7_20, d_arr_mul_7_19, d_arr_mul_7_18, d_arr_mul_7_17, 
      d_arr_mul_7_16, d_arr_mul_7_15, d_arr_mul_7_14, d_arr_mul_7_13, 
      d_arr_mul_7_12, d_arr_mul_7_11, d_arr_mul_7_10, d_arr_mul_7_9, 
      d_arr_mul_7_8, d_arr_mul_7_7, d_arr_mul_7_6, d_arr_mul_7_5, 
      d_arr_mul_7_4, d_arr_mul_7_3, d_arr_mul_7_2, d_arr_mul_7_1, 
      d_arr_mul_7_0, d_arr_mul_8_31, d_arr_mul_8_30, d_arr_mul_8_29, 
      d_arr_mul_8_28, d_arr_mul_8_27, d_arr_mul_8_26, d_arr_mul_8_25, 
      d_arr_mul_8_24, d_arr_mul_8_23, d_arr_mul_8_22, d_arr_mul_8_21, 
      d_arr_mul_8_20, d_arr_mul_8_19, d_arr_mul_8_18, d_arr_mul_8_17, 
      d_arr_mul_8_16, d_arr_mul_8_15, d_arr_mul_8_14, d_arr_mul_8_13, 
      d_arr_mul_8_12, d_arr_mul_8_11, d_arr_mul_8_10, d_arr_mul_8_9, 
      d_arr_mul_8_8, d_arr_mul_8_7, d_arr_mul_8_6, d_arr_mul_8_5, 
      d_arr_mul_8_4, d_arr_mul_8_3, d_arr_mul_8_2, d_arr_mul_8_1, 
      d_arr_mul_8_0, d_arr_mul_9_31, d_arr_mul_9_30, d_arr_mul_9_29, 
      d_arr_mul_9_28, d_arr_mul_9_27, d_arr_mul_9_26, d_arr_mul_9_25, 
      d_arr_mul_9_24, d_arr_mul_9_23, d_arr_mul_9_22, d_arr_mul_9_21, 
      d_arr_mul_9_20, d_arr_mul_9_19, d_arr_mul_9_18, d_arr_mul_9_17, 
      d_arr_mul_9_16, d_arr_mul_9_15, d_arr_mul_9_14, d_arr_mul_9_13, 
      d_arr_mul_9_12, d_arr_mul_9_11, d_arr_mul_9_10, d_arr_mul_9_9, 
      d_arr_mul_9_8, d_arr_mul_9_7, d_arr_mul_9_6, d_arr_mul_9_5, 
      d_arr_mul_9_4, d_arr_mul_9_3, d_arr_mul_9_2, d_arr_mul_9_1, 
      d_arr_mul_9_0, d_arr_mul_10_31, d_arr_mul_10_30, d_arr_mul_10_29, 
      d_arr_mul_10_28, d_arr_mul_10_27, d_arr_mul_10_26, d_arr_mul_10_25, 
      d_arr_mul_10_24, d_arr_mul_10_23, d_arr_mul_10_22, d_arr_mul_10_21, 
      d_arr_mul_10_20, d_arr_mul_10_19, d_arr_mul_10_18, d_arr_mul_10_17, 
      d_arr_mul_10_16, d_arr_mul_10_15, d_arr_mul_10_14, d_arr_mul_10_13, 
      d_arr_mul_10_12, d_arr_mul_10_11, d_arr_mul_10_10, d_arr_mul_10_9, 
      d_arr_mul_10_8, d_arr_mul_10_7, d_arr_mul_10_6, d_arr_mul_10_5, 
      d_arr_mul_10_4, d_arr_mul_10_3, d_arr_mul_10_2, d_arr_mul_10_1, 
      d_arr_mul_10_0, d_arr_mul_11_31, d_arr_mul_11_30, d_arr_mul_11_29, 
      d_arr_mul_11_28, d_arr_mul_11_27, d_arr_mul_11_26, d_arr_mul_11_25, 
      d_arr_mul_11_24, d_arr_mul_11_23, d_arr_mul_11_22, d_arr_mul_11_21, 
      d_arr_mul_11_20, d_arr_mul_11_19, d_arr_mul_11_18, d_arr_mul_11_17, 
      d_arr_mul_11_16, d_arr_mul_11_15, d_arr_mul_11_14, d_arr_mul_11_13, 
      d_arr_mul_11_12, d_arr_mul_11_11, d_arr_mul_11_10, d_arr_mul_11_9, 
      d_arr_mul_11_8, d_arr_mul_11_7, d_arr_mul_11_6, d_arr_mul_11_5, 
      d_arr_mul_11_4, d_arr_mul_11_3, d_arr_mul_11_2, d_arr_mul_11_1, 
      d_arr_mul_11_0, d_arr_mul_12_31, d_arr_mul_12_30, d_arr_mul_12_29, 
      d_arr_mul_12_28, d_arr_mul_12_27, d_arr_mul_12_26, d_arr_mul_12_25, 
      d_arr_mul_12_24, d_arr_mul_12_23, d_arr_mul_12_22, d_arr_mul_12_21, 
      d_arr_mul_12_20, d_arr_mul_12_19, d_arr_mul_12_18, d_arr_mul_12_17, 
      d_arr_mul_12_16, d_arr_mul_12_15, d_arr_mul_12_14, d_arr_mul_12_13, 
      d_arr_mul_12_12, d_arr_mul_12_11, d_arr_mul_12_10, d_arr_mul_12_9, 
      d_arr_mul_12_8, d_arr_mul_12_7, d_arr_mul_12_6, d_arr_mul_12_5, 
      d_arr_mul_12_4, d_arr_mul_12_3, d_arr_mul_12_2, d_arr_mul_12_1, 
      d_arr_mul_12_0, d_arr_mul_13_31, d_arr_mul_13_30, d_arr_mul_13_29, 
      d_arr_mul_13_28, d_arr_mul_13_27, d_arr_mul_13_26, d_arr_mul_13_25, 
      d_arr_mul_13_24, d_arr_mul_13_23, d_arr_mul_13_22, d_arr_mul_13_21, 
      d_arr_mul_13_20, d_arr_mul_13_19, d_arr_mul_13_18, d_arr_mul_13_17, 
      d_arr_mul_13_16, d_arr_mul_13_15, d_arr_mul_13_14, d_arr_mul_13_13, 
      d_arr_mul_13_12, d_arr_mul_13_11, d_arr_mul_13_10, d_arr_mul_13_9, 
      d_arr_mul_13_8, d_arr_mul_13_7, d_arr_mul_13_6, d_arr_mul_13_5, 
      d_arr_mul_13_4, d_arr_mul_13_3, d_arr_mul_13_2, d_arr_mul_13_1, 
      d_arr_mul_13_0, d_arr_mul_14_31, d_arr_mul_14_30, d_arr_mul_14_29, 
      d_arr_mul_14_28, d_arr_mul_14_27, d_arr_mul_14_26, d_arr_mul_14_25, 
      d_arr_mul_14_24, d_arr_mul_14_23, d_arr_mul_14_22, d_arr_mul_14_21, 
      d_arr_mul_14_20, d_arr_mul_14_19, d_arr_mul_14_18, d_arr_mul_14_17, 
      d_arr_mul_14_16, d_arr_mul_14_15, d_arr_mul_14_14, d_arr_mul_14_13, 
      d_arr_mul_14_12, d_arr_mul_14_11, d_arr_mul_14_10, d_arr_mul_14_9, 
      d_arr_mul_14_8, d_arr_mul_14_7, d_arr_mul_14_6, d_arr_mul_14_5, 
      d_arr_mul_14_4, d_arr_mul_14_3, d_arr_mul_14_2, d_arr_mul_14_1, 
      d_arr_mul_14_0, d_arr_mul_15_31, d_arr_mul_15_30, d_arr_mul_15_29, 
      d_arr_mul_15_28, d_arr_mul_15_27, d_arr_mul_15_26, d_arr_mul_15_25, 
      d_arr_mul_15_24, d_arr_mul_15_23, d_arr_mul_15_22, d_arr_mul_15_21, 
      d_arr_mul_15_20, d_arr_mul_15_19, d_arr_mul_15_18, d_arr_mul_15_17, 
      d_arr_mul_15_16, d_arr_mul_15_15, d_arr_mul_15_14, d_arr_mul_15_13, 
      d_arr_mul_15_12, d_arr_mul_15_11, d_arr_mul_15_10, d_arr_mul_15_9, 
      d_arr_mul_15_8, d_arr_mul_15_7, d_arr_mul_15_6, d_arr_mul_15_5, 
      d_arr_mul_15_4, d_arr_mul_15_3, d_arr_mul_15_2, d_arr_mul_15_1, 
      d_arr_mul_15_0, d_arr_mul_16_31, d_arr_mul_16_30, d_arr_mul_16_29, 
      d_arr_mul_16_28, d_arr_mul_16_27, d_arr_mul_16_26, d_arr_mul_16_25, 
      d_arr_mul_16_24, d_arr_mul_16_23, d_arr_mul_16_22, d_arr_mul_16_21, 
      d_arr_mul_16_20, d_arr_mul_16_19, d_arr_mul_16_18, d_arr_mul_16_17, 
      d_arr_mul_16_16, d_arr_mul_16_15, d_arr_mul_16_14, d_arr_mul_16_13, 
      d_arr_mul_16_12, d_arr_mul_16_11, d_arr_mul_16_10, d_arr_mul_16_9, 
      d_arr_mul_16_8, d_arr_mul_16_7, d_arr_mul_16_6, d_arr_mul_16_5, 
      d_arr_mul_16_4, d_arr_mul_16_3, d_arr_mul_16_2, d_arr_mul_16_1, 
      d_arr_mul_16_0, d_arr_mul_17_31, d_arr_mul_17_30, d_arr_mul_17_29, 
      d_arr_mul_17_28, d_arr_mul_17_27, d_arr_mul_17_26, d_arr_mul_17_25, 
      d_arr_mul_17_24, d_arr_mul_17_23, d_arr_mul_17_22, d_arr_mul_17_21, 
      d_arr_mul_17_20, d_arr_mul_17_19, d_arr_mul_17_18, d_arr_mul_17_17, 
      d_arr_mul_17_16, d_arr_mul_17_15, d_arr_mul_17_14, d_arr_mul_17_13, 
      d_arr_mul_17_12, d_arr_mul_17_11, d_arr_mul_17_10, d_arr_mul_17_9, 
      d_arr_mul_17_8, d_arr_mul_17_7, d_arr_mul_17_6, d_arr_mul_17_5, 
      d_arr_mul_17_4, d_arr_mul_17_3, d_arr_mul_17_2, d_arr_mul_17_1, 
      d_arr_mul_17_0, d_arr_mul_18_31, d_arr_mul_18_30, d_arr_mul_18_29, 
      d_arr_mul_18_28, d_arr_mul_18_27, d_arr_mul_18_26, d_arr_mul_18_25, 
      d_arr_mul_18_24, d_arr_mul_18_23, d_arr_mul_18_22, d_arr_mul_18_21, 
      d_arr_mul_18_20, d_arr_mul_18_19, d_arr_mul_18_18, d_arr_mul_18_17, 
      d_arr_mul_18_16, d_arr_mul_18_15, d_arr_mul_18_14, d_arr_mul_18_13, 
      d_arr_mul_18_12, d_arr_mul_18_11, d_arr_mul_18_10, d_arr_mul_18_9, 
      d_arr_mul_18_8, d_arr_mul_18_7, d_arr_mul_18_6, d_arr_mul_18_5, 
      d_arr_mul_18_4, d_arr_mul_18_3, d_arr_mul_18_2, d_arr_mul_18_1, 
      d_arr_mul_18_0, d_arr_mul_19_31, d_arr_mul_19_30, d_arr_mul_19_29, 
      d_arr_mul_19_28, d_arr_mul_19_27, d_arr_mul_19_26, d_arr_mul_19_25, 
      d_arr_mul_19_24, d_arr_mul_19_23, d_arr_mul_19_22, d_arr_mul_19_21, 
      d_arr_mul_19_20, d_arr_mul_19_19, d_arr_mul_19_18, d_arr_mul_19_17, 
      d_arr_mul_19_16, d_arr_mul_19_15, d_arr_mul_19_14, d_arr_mul_19_13, 
      d_arr_mul_19_12, d_arr_mul_19_11, d_arr_mul_19_10, d_arr_mul_19_9, 
      d_arr_mul_19_8, d_arr_mul_19_7, d_arr_mul_19_6, d_arr_mul_19_5, 
      d_arr_mul_19_4, d_arr_mul_19_3, d_arr_mul_19_2, d_arr_mul_19_1, 
      d_arr_mul_19_0, d_arr_mul_20_31, d_arr_mul_20_30, d_arr_mul_20_29, 
      d_arr_mul_20_28, d_arr_mul_20_27, d_arr_mul_20_26, d_arr_mul_20_25, 
      d_arr_mul_20_24, d_arr_mul_20_23, d_arr_mul_20_22, d_arr_mul_20_21, 
      d_arr_mul_20_20, d_arr_mul_20_19, d_arr_mul_20_18, d_arr_mul_20_17, 
      d_arr_mul_20_16, d_arr_mul_20_15, d_arr_mul_20_14, d_arr_mul_20_13, 
      d_arr_mul_20_12, d_arr_mul_20_11, d_arr_mul_20_10, d_arr_mul_20_9, 
      d_arr_mul_20_8, d_arr_mul_20_7, d_arr_mul_20_6, d_arr_mul_20_5, 
      d_arr_mul_20_4, d_arr_mul_20_3, d_arr_mul_20_2, d_arr_mul_20_1, 
      d_arr_mul_20_0, d_arr_mul_21_31, d_arr_mul_21_30, d_arr_mul_21_29, 
      d_arr_mul_21_28, d_arr_mul_21_27, d_arr_mul_21_26, d_arr_mul_21_25, 
      d_arr_mul_21_24, d_arr_mul_21_23, d_arr_mul_21_22, d_arr_mul_21_21, 
      d_arr_mul_21_20, d_arr_mul_21_19, d_arr_mul_21_18, d_arr_mul_21_17, 
      d_arr_mul_21_16, d_arr_mul_21_15, d_arr_mul_21_14, d_arr_mul_21_13, 
      d_arr_mul_21_12, d_arr_mul_21_11, d_arr_mul_21_10, d_arr_mul_21_9, 
      d_arr_mul_21_8, d_arr_mul_21_7, d_arr_mul_21_6, d_arr_mul_21_5, 
      d_arr_mul_21_4, d_arr_mul_21_3, d_arr_mul_21_2, d_arr_mul_21_1, 
      d_arr_mul_21_0, d_arr_mul_22_31, d_arr_mul_22_30, d_arr_mul_22_29, 
      d_arr_mul_22_28, d_arr_mul_22_27, d_arr_mul_22_26, d_arr_mul_22_25, 
      d_arr_mul_22_24, d_arr_mul_22_23, d_arr_mul_22_22, d_arr_mul_22_21, 
      d_arr_mul_22_20, d_arr_mul_22_19, d_arr_mul_22_18, d_arr_mul_22_17, 
      d_arr_mul_22_16, d_arr_mul_22_15, d_arr_mul_22_14, d_arr_mul_22_13, 
      d_arr_mul_22_12, d_arr_mul_22_11, d_arr_mul_22_10, d_arr_mul_22_9, 
      d_arr_mul_22_8, d_arr_mul_22_7, d_arr_mul_22_6, d_arr_mul_22_5, 
      d_arr_mul_22_4, d_arr_mul_22_3, d_arr_mul_22_2, d_arr_mul_22_1, 
      d_arr_mul_22_0, d_arr_mul_23_31, d_arr_mul_23_30, d_arr_mul_23_29, 
      d_arr_mul_23_28, d_arr_mul_23_27, d_arr_mul_23_26, d_arr_mul_23_25, 
      d_arr_mul_23_24, d_arr_mul_23_23, d_arr_mul_23_22, d_arr_mul_23_21, 
      d_arr_mul_23_20, d_arr_mul_23_19, d_arr_mul_23_18, d_arr_mul_23_17, 
      d_arr_mul_23_16, d_arr_mul_23_15, d_arr_mul_23_14, d_arr_mul_23_13, 
      d_arr_mul_23_12, d_arr_mul_23_11, d_arr_mul_23_10, d_arr_mul_23_9, 
      d_arr_mul_23_8, d_arr_mul_23_7, d_arr_mul_23_6, d_arr_mul_23_5, 
      d_arr_mul_23_4, d_arr_mul_23_3, d_arr_mul_23_2, d_arr_mul_23_1, 
      d_arr_mul_23_0, d_arr_mul_24_31, d_arr_mul_24_30, d_arr_mul_24_29, 
      d_arr_mul_24_28, d_arr_mul_24_27, d_arr_mul_24_26, d_arr_mul_24_25, 
      d_arr_mul_24_24, d_arr_mul_24_23, d_arr_mul_24_22, d_arr_mul_24_21, 
      d_arr_mul_24_20, d_arr_mul_24_19, d_arr_mul_24_18, d_arr_mul_24_17, 
      d_arr_mul_24_16, d_arr_mul_24_15, d_arr_mul_24_14, d_arr_mul_24_13, 
      d_arr_mul_24_12, d_arr_mul_24_11, d_arr_mul_24_10, d_arr_mul_24_9, 
      d_arr_mul_24_8, d_arr_mul_24_7, d_arr_mul_24_6, d_arr_mul_24_5, 
      d_arr_mul_24_4, d_arr_mul_24_3, d_arr_mul_24_2, d_arr_mul_24_1, 
      d_arr_mul_24_0, d_arr_add_0_31, d_arr_add_0_30, d_arr_add_0_29, 
      d_arr_add_0_28, d_arr_add_0_27, d_arr_add_0_26, d_arr_add_0_25, 
      d_arr_add_0_24, d_arr_add_0_23, d_arr_add_0_22, d_arr_add_0_21, 
      d_arr_add_0_20, d_arr_add_0_19, d_arr_add_0_18, d_arr_add_0_17, 
      d_arr_add_0_16, d_arr_add_0_15, d_arr_add_0_14, d_arr_add_0_13, 
      d_arr_add_0_12, d_arr_add_0_11, d_arr_add_0_10, d_arr_add_0_9, 
      d_arr_add_0_8, d_arr_add_0_7, d_arr_add_0_6, d_arr_add_0_5, 
      d_arr_add_0_4, d_arr_add_0_3, d_arr_add_0_2, d_arr_add_0_1, 
      d_arr_add_0_0, d_arr_add_1_31, d_arr_add_1_30, d_arr_add_1_29, 
      d_arr_add_1_28, d_arr_add_1_27, d_arr_add_1_26, d_arr_add_1_25, 
      d_arr_add_1_24, d_arr_add_1_23, d_arr_add_1_22, d_arr_add_1_21, 
      d_arr_add_1_20, d_arr_add_1_19, d_arr_add_1_18, d_arr_add_1_17, 
      d_arr_add_1_16, d_arr_add_1_15, d_arr_add_1_14, d_arr_add_1_13, 
      d_arr_add_1_12, d_arr_add_1_11, d_arr_add_1_10, d_arr_add_1_9, 
      d_arr_add_1_8, d_arr_add_1_7, d_arr_add_1_6, d_arr_add_1_5, 
      d_arr_add_1_4, d_arr_add_1_3, d_arr_add_1_2, d_arr_add_1_1, 
      d_arr_add_1_0, d_arr_add_2_31, d_arr_add_2_30, d_arr_add_2_29, 
      d_arr_add_2_28, d_arr_add_2_27, d_arr_add_2_26, d_arr_add_2_25, 
      d_arr_add_2_24, d_arr_add_2_23, d_arr_add_2_22, d_arr_add_2_21, 
      d_arr_add_2_20, d_arr_add_2_19, d_arr_add_2_18, d_arr_add_2_17, 
      d_arr_add_2_16, d_arr_add_2_15, d_arr_add_2_14, d_arr_add_2_13, 
      d_arr_add_2_12, d_arr_add_2_11, d_arr_add_2_10, d_arr_add_2_9, 
      d_arr_add_2_8, d_arr_add_2_7, d_arr_add_2_6, d_arr_add_2_5, 
      d_arr_add_2_4, d_arr_add_2_3, d_arr_add_2_2, d_arr_add_2_1, 
      d_arr_add_2_0, d_arr_add_3_31, d_arr_add_3_30, d_arr_add_3_29, 
      d_arr_add_3_28, d_arr_add_3_27, d_arr_add_3_26, d_arr_add_3_25, 
      d_arr_add_3_24, d_arr_add_3_23, d_arr_add_3_22, d_arr_add_3_21, 
      d_arr_add_3_20, d_arr_add_3_19, d_arr_add_3_18, d_arr_add_3_17, 
      d_arr_add_3_16, d_arr_add_3_15, d_arr_add_3_14, d_arr_add_3_13, 
      d_arr_add_3_12, d_arr_add_3_11, d_arr_add_3_10, d_arr_add_3_9, 
      d_arr_add_3_8, d_arr_add_3_7, d_arr_add_3_6, d_arr_add_3_5, 
      d_arr_add_3_4, d_arr_add_3_3, d_arr_add_3_2, d_arr_add_3_1, 
      d_arr_add_3_0, d_arr_add_9_31, d_arr_add_9_30, d_arr_add_9_29, 
      d_arr_add_9_28, d_arr_add_9_27, d_arr_add_9_26, d_arr_add_9_25, 
      d_arr_add_9_24, d_arr_add_9_23, d_arr_add_9_22, d_arr_add_9_21, 
      d_arr_add_9_20, d_arr_add_9_19, d_arr_add_9_18, d_arr_add_9_17, 
      d_arr_add_9_16, d_arr_add_9_15, d_arr_add_9_14, d_arr_add_9_13, 
      d_arr_add_9_12, d_arr_add_9_11, d_arr_add_9_10, d_arr_add_9_9, 
      d_arr_add_9_8, d_arr_add_9_7, d_arr_add_9_6, d_arr_add_9_5, 
      d_arr_add_9_4, d_arr_add_9_3, d_arr_add_9_2, d_arr_add_9_1, 
      d_arr_add_9_0, d_arr_add_10_31, d_arr_add_10_30, d_arr_add_10_29, 
      d_arr_add_10_28, d_arr_add_10_27, d_arr_add_10_26, d_arr_add_10_25, 
      d_arr_add_10_24, d_arr_add_10_23, d_arr_add_10_22, d_arr_add_10_21, 
      d_arr_add_10_20, d_arr_add_10_19, d_arr_add_10_18, d_arr_add_10_17, 
      d_arr_add_10_16, d_arr_add_10_15, d_arr_add_10_14, d_arr_add_10_13, 
      d_arr_add_10_12, d_arr_add_10_11, d_arr_add_10_10, d_arr_add_10_9, 
      d_arr_add_10_8, d_arr_add_10_7, d_arr_add_10_6, d_arr_add_10_5, 
      d_arr_add_10_4, d_arr_add_10_3, d_arr_add_10_2, d_arr_add_10_1, 
      d_arr_add_10_0, d_arr_add_11_31, d_arr_add_11_30, d_arr_add_11_29, 
      d_arr_add_11_28, d_arr_add_11_27, d_arr_add_11_26, d_arr_add_11_25, 
      d_arr_add_11_24, d_arr_add_11_23, d_arr_add_11_22, d_arr_add_11_21, 
      d_arr_add_11_20, d_arr_add_11_19, d_arr_add_11_18, d_arr_add_11_17, 
      d_arr_add_11_16, d_arr_add_11_15, d_arr_add_11_14, d_arr_add_11_13, 
      d_arr_add_11_12, d_arr_add_11_11, d_arr_add_11_10, d_arr_add_11_9, 
      d_arr_add_11_8, d_arr_add_11_7, d_arr_add_11_6, d_arr_add_11_5, 
      d_arr_add_11_4, d_arr_add_11_3, d_arr_add_11_2, d_arr_add_11_1, 
      d_arr_add_11_0, d_arr_add_12_31, d_arr_add_12_30, d_arr_add_12_29, 
      d_arr_add_12_28, d_arr_add_12_27, d_arr_add_12_26, d_arr_add_12_25, 
      d_arr_add_12_24, d_arr_add_12_23, d_arr_add_12_22, d_arr_add_12_21, 
      d_arr_add_12_20, d_arr_add_12_19, d_arr_add_12_18, d_arr_add_12_17, 
      d_arr_add_12_16, d_arr_add_12_15, d_arr_add_12_14, d_arr_add_12_13, 
      d_arr_add_12_12, d_arr_add_12_11, d_arr_add_12_10, d_arr_add_12_9, 
      d_arr_add_12_8, d_arr_add_12_7, d_arr_add_12_6, d_arr_add_12_5, 
      d_arr_add_12_4, d_arr_add_12_3, d_arr_add_12_2, d_arr_add_12_1, 
      d_arr_add_12_0, d_arr_add_18_31, d_arr_add_18_30, d_arr_add_18_29, 
      d_arr_add_18_28, d_arr_add_18_27, d_arr_add_18_26, d_arr_add_18_25, 
      d_arr_add_18_24, d_arr_add_18_23, d_arr_add_18_22, d_arr_add_18_21, 
      d_arr_add_18_20, d_arr_add_18_19, d_arr_add_18_18, d_arr_add_18_17, 
      d_arr_add_18_16, d_arr_add_18_15, d_arr_add_18_14, d_arr_add_18_13, 
      d_arr_add_18_12, d_arr_add_18_11, d_arr_add_18_10, d_arr_add_18_9, 
      d_arr_add_18_8, d_arr_add_18_7, d_arr_add_18_6, d_arr_add_18_5, 
      d_arr_add_18_4, d_arr_add_18_3, d_arr_add_18_2, d_arr_add_18_1, 
      d_arr_add_18_0, d_arr_add_19_31, d_arr_add_19_30, d_arr_add_19_29, 
      d_arr_add_19_28, d_arr_add_19_27, d_arr_add_19_26, d_arr_add_19_25, 
      d_arr_add_19_24, d_arr_add_19_23, d_arr_add_19_22, d_arr_add_19_21, 
      d_arr_add_19_20, d_arr_add_19_19, d_arr_add_19_18, d_arr_add_19_17, 
      d_arr_add_19_16, d_arr_add_19_15, d_arr_add_19_14, d_arr_add_19_13, 
      d_arr_add_19_12, d_arr_add_19_11, d_arr_add_19_10, d_arr_add_19_9, 
      d_arr_add_19_8, d_arr_add_19_7, d_arr_add_19_6, d_arr_add_19_5, 
      d_arr_add_19_4, d_arr_add_19_3, d_arr_add_19_2, d_arr_add_19_1, 
      d_arr_add_19_0, d_arr_add_20_31, d_arr_add_20_30, d_arr_add_20_29, 
      d_arr_add_20_28, d_arr_add_20_27, d_arr_add_20_26, d_arr_add_20_25, 
      d_arr_add_20_24, d_arr_add_20_23, d_arr_add_20_22, d_arr_add_20_21, 
      d_arr_add_20_20, d_arr_add_20_19, d_arr_add_20_18, d_arr_add_20_17, 
      d_arr_add_20_16, d_arr_add_20_15, d_arr_add_20_14, d_arr_add_20_13, 
      d_arr_add_20_12, d_arr_add_20_11, d_arr_add_20_10, d_arr_add_20_9, 
      d_arr_add_20_8, d_arr_add_20_7, d_arr_add_20_6, d_arr_add_20_5, 
      d_arr_add_20_4, d_arr_add_20_3, d_arr_add_20_2, d_arr_add_20_1, 
      d_arr_add_20_0, d_arr_merge1_0_31, d_arr_merge1_0_30, 
      d_arr_merge1_0_29, d_arr_merge1_0_28, d_arr_merge1_0_27, 
      d_arr_merge1_0_26, d_arr_merge1_0_25, d_arr_merge1_0_24, 
      d_arr_merge1_0_23, d_arr_merge1_0_22, d_arr_merge1_0_21, 
      d_arr_merge1_0_20, d_arr_merge1_0_19, d_arr_merge1_0_18, 
      d_arr_merge1_0_17, d_arr_merge1_0_16, d_arr_merge1_0_15, 
      d_arr_merge1_0_14, d_arr_merge1_0_13, d_arr_merge1_0_12, 
      d_arr_merge1_0_11, d_arr_merge1_0_10, d_arr_merge1_0_9, 
      d_arr_merge1_0_8, d_arr_merge1_0_7, d_arr_merge1_0_6, d_arr_merge1_0_5, 
      d_arr_merge1_0_4, d_arr_merge1_0_3, d_arr_merge1_0_2, d_arr_merge1_0_1, 
      d_arr_merge1_0_0, d_arr_merge1_1_31, d_arr_merge1_1_30, 
      d_arr_merge1_1_29, d_arr_merge1_1_28, d_arr_merge1_1_27, 
      d_arr_merge1_1_26, d_arr_merge1_1_25, d_arr_merge1_1_24, 
      d_arr_merge1_1_23, d_arr_merge1_1_22, d_arr_merge1_1_21, 
      d_arr_merge1_1_20, d_arr_merge1_1_19, d_arr_merge1_1_18, 
      d_arr_merge1_1_17, d_arr_merge1_1_16, d_arr_merge1_1_15, 
      d_arr_merge1_1_14, d_arr_merge1_1_13, d_arr_merge1_1_12, 
      d_arr_merge1_1_11, d_arr_merge1_1_10, d_arr_merge1_1_9, 
      d_arr_merge1_1_8, d_arr_merge1_1_7, d_arr_merge1_1_6, d_arr_merge1_1_5, 
      d_arr_merge1_1_4, d_arr_merge1_1_3, d_arr_merge1_1_2, d_arr_merge1_1_1, 
      d_arr_merge1_1_0, d_arr_merge2_0_31, d_arr_merge2_0_26, 
      d_arr_merge2_0_25, d_arr_merge2_0_24, d_arr_merge2_0_23, 
      d_arr_merge2_0_22, d_arr_merge2_0_21, d_arr_merge2_0_20, 
      d_arr_merge2_0_19, d_arr_merge2_0_18, d_arr_merge2_0_17, 
      d_arr_merge2_0_16, d_arr_merge2_0_15, d_arr_merge2_0_14, 
      d_arr_merge2_0_13, d_arr_merge2_0_12, d_arr_merge2_0_11, 
      d_arr_merge2_0_10, d_arr_merge2_0_9, d_arr_merge2_0_8, 
      d_arr_merge2_0_7, d_arr_merge2_0_6, d_arr_merge2_0_5, d_arr_merge2_0_4, 
      d_arr_merge2_0_3, d_arr_merge2_0_2, d_arr_merge2_0_1, d_arr_merge2_0_0, 
      d_arr_merge2_1_31, d_arr_merge2_1_26, d_arr_merge2_1_25, 
      d_arr_merge2_1_24, d_arr_merge2_1_23, d_arr_merge2_1_22, 
      d_arr_merge2_1_21, d_arr_merge2_1_20, d_arr_merge2_1_19, 
      d_arr_merge2_1_18, d_arr_merge2_1_17, d_arr_merge2_1_16, 
      d_arr_merge2_1_15, d_arr_merge2_1_14, d_arr_merge2_1_13, 
      d_arr_merge2_1_12, d_arr_merge2_1_11, d_arr_merge2_1_10, 
      d_arr_merge2_1_9, d_arr_merge2_1_8, d_arr_merge2_1_7, d_arr_merge2_1_6, 
      d_arr_merge2_1_5, d_arr_merge2_1_4, d_arr_merge2_1_3, d_arr_merge2_1_2, 
      d_arr_merge2_1_1, d_arr_merge2_1_0, d_arr_relu_0_31, d_arr_relu_0_30, 
      d_arr_relu_0_29, d_arr_relu_0_28, d_arr_relu_0_27, d_arr_relu_0_26, 
      d_arr_relu_0_25, d_arr_relu_0_24, d_arr_relu_0_23, d_arr_relu_0_22, 
      d_arr_relu_0_21, d_arr_relu_0_20, d_arr_relu_0_19, d_arr_relu_0_18, 
      d_arr_relu_0_17, d_arr_relu_0_16, d_arr_relu_0_14, d_arr_relu_0_13, 
      d_arr_relu_0_12, d_arr_relu_0_11, d_arr_relu_0_10, d_arr_relu_0_9, 
      d_arr_relu_0_8, d_arr_relu_0_7, d_arr_relu_0_6, d_arr_relu_0_5, 
      d_arr_relu_0_4, d_arr_relu_0_3, d_arr_relu_0_2, d_arr_relu_0_1, 
      d_arr_relu_0_0, d_arr_relu_1_31, d_arr_relu_1_30, d_arr_relu_1_29, 
      d_arr_relu_1_28, d_arr_relu_1_27, d_arr_relu_1_26, d_arr_relu_1_25, 
      d_arr_relu_1_24, d_arr_relu_1_23, d_arr_relu_1_22, d_arr_relu_1_21, 
      d_arr_relu_1_20, d_arr_relu_1_19, d_arr_relu_1_18, d_arr_relu_1_17, 
      d_arr_relu_1_16, d_arr_relu_1_14, d_arr_relu_1_13, d_arr_relu_1_12, 
      d_arr_relu_1_11, d_arr_relu_1_10, d_arr_relu_1_9, d_arr_relu_1_8, 
      d_arr_relu_1_7, d_arr_relu_1_6, d_arr_relu_1_5, d_arr_relu_1_4, 
      d_arr_relu_1_3, d_arr_relu_1_2, d_arr_relu_1_1, d_arr_relu_1_0, 
      sel_mul, sel_add, GND0, counter_12, counter_11, counter_10, counter_9, 
      counter_7, counter_6, counter_5, counter_4, counter_3, counter_2, 
      counter_1, nx20, nx92, nx194, nx16101, nx16115, nx16125, nx16135, 
      nx16145, nx16155, nx16165, nx16175, nx16185, nx16195, nx16205, nx16215, 
      nx16225, nx16235, nx16245, nx16255, nx16265, nx16276, nx16278, nx16281, 
      nx16285, nx16289, nx16293, nx16295, nx16299, nx16301, nx16306, nx16309, 
      nx16313, nx16315, nx16319, nx16321, nx16325, nx16327, nx16331, nx16333, 
      nx16337, nx16339, nx16343, nx16345, nx16349, nx16351, nx16353, nx16361, 
      nx16363, nx16366, nx16371, nx16373, nx16375, nx16380, nx16382, nx16386, 
      nx16388, nx16390, nx16399, nx16401, nx16403, nx16405, nx16407, nx16409, 
      nx16411, nx16413, nx16415, nx16417, nx16419, nx16421, nx16423, nx16425, 
      nx16427, nx16429, nx16431, nx16433, nx16435, nx16437, nx16439, nx16441, 
      nx16443, nx16445, nx16447, nx16449, nx16451, nx16453, nx16455, nx16457, 
      nx16459, nx16461, nx16463, nx16465, nx16467, nx16469, nx16471, nx16473, 
      nx16475, nx16477, nx16479, nx16481, nx16483, nx16485, nx16487, nx16489, 
      nx16491, nx16497, nx16499, nx16501, nx16503, nx16505, nx16507, nx16509, 
      nx16511, nx16513, nx16515, nx16517, nx16519, nx16521, nx16523, nx16525, 
      nx16527, nx16529, nx16531, nx16533, nx16535, nx16537, nx16539, nx16541, 
      nx16543, nx16545, nx16547, nx16549, nx16551, nx16553, nx16555, nx16557, 
      nx16559, nx16561, nx16563, nx16565, nx16567, nx16569, nx16571, nx16573, 
      nx16575, nx16577, nx16579, nx16581, nx16583, nx16585, nx16587, nx16589, 
      nx16591, nx16593, nx16595, nx16597, nx16599, nx16601, nx16603, nx16605, 
      nx16607, nx16609, nx16611, nx16613, nx16615, nx16617, nx16619, nx16621, 
      nx16623, nx16625, nx16627, nx16629, nx16631, nx16633, nx16635, nx16637, 
      nx16639, nx16641, nx16643, nx16645, nx16651, nx16653, nx16659, nx16661, 
      nx16663, nx16665, nx16667, nx19388, nx19390, nx19396, nx19398, nx19400, 
      nx19402, nx19404, nx19406, nx19408, nx19410, nx19412, nx19414, nx19416, 
      nx19418, nx19420, nx19422, nx19424, nx19426, nx19428, nx19430, nx19432, 
      nx19434, nx19436, nx19438, nx19440, nx19442, nx19444, nx19446, nx19448, 
      nx19450, nx19452, nx19454, nx19456, nx19458, nx19460, nx19462, nx19464, 
      nx19466, nx19468, nx19470, nx19472, nx19474, nx19476, nx19478, nx19480, 
      nx19482, nx19484, nx19486, nx19488, nx19490, nx19492, nx19494: 
   std_logic ;
   
   signal DANGLING : std_logic_vector (2710 downto 0 );

begin
   buffer_ready <= buffer_ready_EXMPLR ;
   semi_ready <= semi_ready_EXMPLR ;
   cache_muxer_gen : CacheMuxer port map ( d_arr_mux_0_31=>img_data_0_15, 
      d_arr_mux_0_30=>GND0, d_arr_mux_0_29=>GND0, d_arr_mux_0_28=>GND0, 
      d_arr_mux_0_27=>GND0, d_arr_mux_0_26=>GND0, d_arr_mux_0_25=>GND0, 
      d_arr_mux_0_24=>GND0, d_arr_mux_0_23=>GND0, d_arr_mux_0_22=>GND0, 
      d_arr_mux_0_21=>GND0, d_arr_mux_0_20=>GND0, d_arr_mux_0_19=>GND0, 
      d_arr_mux_0_18=>GND0, d_arr_mux_0_17=>GND0, d_arr_mux_0_16=>GND0, 
      d_arr_mux_0_15=>GND0, d_arr_mux_0_14=>nx19396, d_arr_mux_0_13=>
      img_data_0_13, d_arr_mux_0_12=>img_data_0_12, d_arr_mux_0_11=>
      img_data_0_11, d_arr_mux_0_10=>img_data_0_10, d_arr_mux_0_9=>
      img_data_0_9, d_arr_mux_0_8=>img_data_0_8, d_arr_mux_0_7=>img_data_0_7, 
      d_arr_mux_0_6=>img_data_0_6, d_arr_mux_0_5=>img_data_0_5, 
      d_arr_mux_0_4=>img_data_0_4, d_arr_mux_0_3=>img_data_0_3, 
      d_arr_mux_0_2=>img_data_0_2, d_arr_mux_0_1=>img_data_0_1, 
      d_arr_mux_0_0=>img_data_0_0, d_arr_mux_1_31=>img_data_1_15, 
      d_arr_mux_1_30=>GND0, d_arr_mux_1_29=>GND0, d_arr_mux_1_28=>GND0, 
      d_arr_mux_1_27=>GND0, d_arr_mux_1_26=>GND0, d_arr_mux_1_25=>GND0, 
      d_arr_mux_1_24=>GND0, d_arr_mux_1_23=>GND0, d_arr_mux_1_22=>GND0, 
      d_arr_mux_1_21=>GND0, d_arr_mux_1_20=>GND0, d_arr_mux_1_19=>GND0, 
      d_arr_mux_1_18=>GND0, d_arr_mux_1_17=>GND0, d_arr_mux_1_16=>GND0, 
      d_arr_mux_1_15=>GND0, d_arr_mux_1_14=>nx19398, d_arr_mux_1_13=>
      img_data_1_13, d_arr_mux_1_12=>img_data_1_12, d_arr_mux_1_11=>
      img_data_1_11, d_arr_mux_1_10=>nx19402, d_arr_mux_1_9=>img_data_1_9, 
      d_arr_mux_1_8=>img_data_1_8, d_arr_mux_1_7=>img_data_1_7, 
      d_arr_mux_1_6=>img_data_1_6, d_arr_mux_1_5=>img_data_1_5, 
      d_arr_mux_1_4=>img_data_1_4, d_arr_mux_1_3=>img_data_1_3, 
      d_arr_mux_1_2=>img_data_1_2, d_arr_mux_1_1=>img_data_1_1, 
      d_arr_mux_1_0=>img_data_1_0, d_arr_mux_2_31=>img_data_2_15, 
      d_arr_mux_2_30=>GND0, d_arr_mux_2_29=>GND0, d_arr_mux_2_28=>GND0, 
      d_arr_mux_2_27=>GND0, d_arr_mux_2_26=>GND0, d_arr_mux_2_25=>GND0, 
      d_arr_mux_2_24=>GND0, d_arr_mux_2_23=>GND0, d_arr_mux_2_22=>GND0, 
      d_arr_mux_2_21=>GND0, d_arr_mux_2_20=>GND0, d_arr_mux_2_19=>GND0, 
      d_arr_mux_2_18=>GND0, d_arr_mux_2_17=>GND0, d_arr_mux_2_16=>GND0, 
      d_arr_mux_2_15=>GND0, d_arr_mux_2_14=>nx19404, d_arr_mux_2_13=>
      img_data_2_13, d_arr_mux_2_12=>img_data_2_12, d_arr_mux_2_11=>
      img_data_2_11, d_arr_mux_2_10=>nx19408, d_arr_mux_2_9=>img_data_2_9, 
      d_arr_mux_2_8=>img_data_2_8, d_arr_mux_2_7=>img_data_2_7, 
      d_arr_mux_2_6=>img_data_2_6, d_arr_mux_2_5=>img_data_2_5, 
      d_arr_mux_2_4=>img_data_2_4, d_arr_mux_2_3=>img_data_2_3, 
      d_arr_mux_2_2=>img_data_2_2, d_arr_mux_2_1=>img_data_2_1, 
      d_arr_mux_2_0=>img_data_2_0, d_arr_mux_3_31=>img_data_5_15, 
      d_arr_mux_3_30=>GND0, d_arr_mux_3_29=>GND0, d_arr_mux_3_28=>GND0, 
      d_arr_mux_3_27=>GND0, d_arr_mux_3_26=>GND0, d_arr_mux_3_25=>GND0, 
      d_arr_mux_3_24=>GND0, d_arr_mux_3_23=>GND0, d_arr_mux_3_22=>GND0, 
      d_arr_mux_3_21=>GND0, d_arr_mux_3_20=>GND0, d_arr_mux_3_19=>GND0, 
      d_arr_mux_3_18=>GND0, d_arr_mux_3_17=>GND0, d_arr_mux_3_16=>GND0, 
      d_arr_mux_3_15=>GND0, d_arr_mux_3_14=>nx19410, d_arr_mux_3_13=>
      img_data_5_13, d_arr_mux_3_12=>img_data_5_12, d_arr_mux_3_11=>
      img_data_5_11, d_arr_mux_3_10=>img_data_5_10, d_arr_mux_3_9=>
      img_data_5_9, d_arr_mux_3_8=>img_data_5_8, d_arr_mux_3_7=>img_data_5_7, 
      d_arr_mux_3_6=>img_data_5_6, d_arr_mux_3_5=>img_data_5_5, 
      d_arr_mux_3_4=>img_data_5_4, d_arr_mux_3_3=>img_data_5_3, 
      d_arr_mux_3_2=>img_data_5_2, d_arr_mux_3_1=>img_data_5_1, 
      d_arr_mux_3_0=>img_data_5_0, d_arr_mux_4_31=>img_data_6_15, 
      d_arr_mux_4_30=>GND0, d_arr_mux_4_29=>GND0, d_arr_mux_4_28=>GND0, 
      d_arr_mux_4_27=>GND0, d_arr_mux_4_26=>GND0, d_arr_mux_4_25=>GND0, 
      d_arr_mux_4_24=>GND0, d_arr_mux_4_23=>GND0, d_arr_mux_4_22=>GND0, 
      d_arr_mux_4_21=>GND0, d_arr_mux_4_20=>GND0, d_arr_mux_4_19=>GND0, 
      d_arr_mux_4_18=>GND0, d_arr_mux_4_17=>GND0, d_arr_mux_4_16=>GND0, 
      d_arr_mux_4_15=>GND0, d_arr_mux_4_14=>nx19412, d_arr_mux_4_13=>
      img_data_6_13, d_arr_mux_4_12=>img_data_6_12, d_arr_mux_4_11=>
      img_data_6_11, d_arr_mux_4_10=>nx19416, d_arr_mux_4_9=>img_data_6_9, 
      d_arr_mux_4_8=>img_data_6_8, d_arr_mux_4_7=>img_data_6_7, 
      d_arr_mux_4_6=>img_data_6_6, d_arr_mux_4_5=>img_data_6_5, 
      d_arr_mux_4_4=>img_data_6_4, d_arr_mux_4_3=>img_data_6_3, 
      d_arr_mux_4_2=>img_data_6_2, d_arr_mux_4_1=>img_data_6_1, 
      d_arr_mux_4_0=>img_data_6_0, d_arr_mux_5_31=>nx16659, d_arr_mux_5_30=>
      GND0, d_arr_mux_5_29=>GND0, d_arr_mux_5_28=>GND0, d_arr_mux_5_27=>GND0, 
      d_arr_mux_5_26=>GND0, d_arr_mux_5_25=>GND0, d_arr_mux_5_24=>GND0, 
      d_arr_mux_5_23=>GND0, d_arr_mux_5_22=>GND0, d_arr_mux_5_21=>GND0, 
      d_arr_mux_5_20=>GND0, d_arr_mux_5_19=>GND0, d_arr_mux_5_18=>GND0, 
      d_arr_mux_5_17=>GND0, d_arr_mux_5_16=>GND0, d_arr_mux_5_15=>GND0, 
      d_arr_mux_5_14=>nx19418, d_arr_mux_5_13=>img_data_7_13, d_arr_mux_5_12
      =>img_data_7_12, d_arr_mux_5_11=>img_data_7_11, d_arr_mux_5_10=>
      nx19422, d_arr_mux_5_9=>img_data_7_9, d_arr_mux_5_8=>img_data_7_8, 
      d_arr_mux_5_7=>img_data_7_7, d_arr_mux_5_6=>img_data_7_6, 
      d_arr_mux_5_5=>img_data_7_5, d_arr_mux_5_4=>img_data_7_4, 
      d_arr_mux_5_3=>img_data_7_3, d_arr_mux_5_2=>img_data_7_2, 
      d_arr_mux_5_1=>img_data_7_1, d_arr_mux_5_0=>img_data_7_0, 
      d_arr_mux_6_31=>img_data_10_15, d_arr_mux_6_30=>GND0, d_arr_mux_6_29=>
      GND0, d_arr_mux_6_28=>GND0, d_arr_mux_6_27=>GND0, d_arr_mux_6_26=>GND0, 
      d_arr_mux_6_25=>GND0, d_arr_mux_6_24=>GND0, d_arr_mux_6_23=>GND0, 
      d_arr_mux_6_22=>GND0, d_arr_mux_6_21=>GND0, d_arr_mux_6_20=>GND0, 
      d_arr_mux_6_19=>GND0, d_arr_mux_6_18=>GND0, d_arr_mux_6_17=>GND0, 
      d_arr_mux_6_16=>GND0, d_arr_mux_6_15=>GND0, d_arr_mux_6_14=>nx19424, 
      d_arr_mux_6_13=>img_data_10_13, d_arr_mux_6_12=>img_data_10_12, 
      d_arr_mux_6_11=>img_data_10_11, d_arr_mux_6_10=>img_data_10_10, 
      d_arr_mux_6_9=>img_data_10_9, d_arr_mux_6_8=>img_data_10_8, 
      d_arr_mux_6_7=>img_data_10_7, d_arr_mux_6_6=>img_data_10_6, 
      d_arr_mux_6_5=>img_data_10_5, d_arr_mux_6_4=>img_data_10_4, 
      d_arr_mux_6_3=>img_data_10_3, d_arr_mux_6_2=>img_data_10_2, 
      d_arr_mux_6_1=>img_data_10_1, d_arr_mux_6_0=>img_data_10_0, 
      d_arr_mux_7_31=>nx16661, d_arr_mux_7_30=>GND0, d_arr_mux_7_29=>GND0, 
      d_arr_mux_7_28=>GND0, d_arr_mux_7_27=>GND0, d_arr_mux_7_26=>GND0, 
      d_arr_mux_7_25=>GND0, d_arr_mux_7_24=>GND0, d_arr_mux_7_23=>GND0, 
      d_arr_mux_7_22=>GND0, d_arr_mux_7_21=>GND0, d_arr_mux_7_20=>GND0, 
      d_arr_mux_7_19=>GND0, d_arr_mux_7_18=>GND0, d_arr_mux_7_17=>GND0, 
      d_arr_mux_7_16=>GND0, d_arr_mux_7_15=>GND0, d_arr_mux_7_14=>nx19426, 
      d_arr_mux_7_13=>img_data_11_13, d_arr_mux_7_12=>img_data_11_12, 
      d_arr_mux_7_11=>img_data_11_11, d_arr_mux_7_10=>nx19430, d_arr_mux_7_9
      =>img_data_11_9, d_arr_mux_7_8=>img_data_11_8, d_arr_mux_7_7=>
      img_data_11_7, d_arr_mux_7_6=>img_data_11_6, d_arr_mux_7_5=>
      img_data_11_5, d_arr_mux_7_4=>img_data_11_4, d_arr_mux_7_3=>
      img_data_11_3, d_arr_mux_7_2=>img_data_11_2, d_arr_mux_7_1=>
      img_data_11_1, d_arr_mux_7_0=>img_data_11_0, d_arr_mux_8_31=>nx16663, 
      d_arr_mux_8_30=>GND0, d_arr_mux_8_29=>GND0, d_arr_mux_8_28=>GND0, 
      d_arr_mux_8_27=>GND0, d_arr_mux_8_26=>GND0, d_arr_mux_8_25=>GND0, 
      d_arr_mux_8_24=>GND0, d_arr_mux_8_23=>GND0, d_arr_mux_8_22=>GND0, 
      d_arr_mux_8_21=>GND0, d_arr_mux_8_20=>GND0, d_arr_mux_8_19=>GND0, 
      d_arr_mux_8_18=>GND0, d_arr_mux_8_17=>GND0, d_arr_mux_8_16=>GND0, 
      d_arr_mux_8_15=>GND0, d_arr_mux_8_14=>nx19432, d_arr_mux_8_13=>
      img_data_12_13, d_arr_mux_8_12=>img_data_12_12, d_arr_mux_8_11=>
      img_data_12_11, d_arr_mux_8_10=>nx19436, d_arr_mux_8_9=>img_data_12_9, 
      d_arr_mux_8_8=>img_data_12_8, d_arr_mux_8_7=>img_data_12_7, 
      d_arr_mux_8_6=>img_data_12_6, d_arr_mux_8_5=>img_data_12_5, 
      d_arr_mux_8_4=>img_data_12_4, d_arr_mux_8_3=>img_data_12_3, 
      d_arr_mux_8_2=>img_data_12_2, d_arr_mux_8_1=>img_data_12_1, 
      d_arr_mux_8_0=>img_data_12_0, d_arr_mux_9_31=>nx16401, d_arr_mux_9_30
      =>nx16401, d_arr_mux_9_29=>nx16401, d_arr_mux_9_28=>nx16401, 
      d_arr_mux_9_27=>nx16401, d_arr_mux_9_26=>nx16401, d_arr_mux_9_25=>
      nx16401, d_arr_mux_9_24=>nx16403, d_arr_mux_9_23=>nx16403, 
      d_arr_mux_9_22=>nx16403, d_arr_mux_9_21=>nx16403, d_arr_mux_9_20=>
      nx16403, d_arr_mux_9_19=>nx16403, d_arr_mux_9_18=>nx16403, 
      d_arr_mux_9_17=>nx16405, d_arr_mux_9_16=>nx16405, d_arr_mux_9_15=>
      nx16405, d_arr_mux_9_14=>ordered_img_data_9_14, d_arr_mux_9_13=>
      ordered_img_data_9_13, d_arr_mux_9_12=>ordered_img_data_9_12, 
      d_arr_mux_9_11=>ordered_img_data_9_11, d_arr_mux_9_10=>
      ordered_img_data_9_10, d_arr_mux_9_9=>ordered_img_data_9_9, 
      d_arr_mux_9_8=>ordered_img_data_9_8, d_arr_mux_9_7=>
      ordered_img_data_9_7, d_arr_mux_9_6=>ordered_img_data_9_6, 
      d_arr_mux_9_5=>ordered_img_data_9_5, d_arr_mux_9_4=>
      ordered_img_data_9_4, d_arr_mux_9_3=>ordered_img_data_9_3, 
      d_arr_mux_9_2=>ordered_img_data_9_2, d_arr_mux_9_1=>
      ordered_img_data_9_1, d_arr_mux_9_0=>ordered_img_data_9_0, 
      d_arr_mux_10_31=>nx16409, d_arr_mux_10_30=>nx16409, d_arr_mux_10_29=>
      nx16409, d_arr_mux_10_28=>nx16409, d_arr_mux_10_27=>nx16409, 
      d_arr_mux_10_26=>nx16409, d_arr_mux_10_25=>nx16409, d_arr_mux_10_24=>
      nx16411, d_arr_mux_10_23=>nx16411, d_arr_mux_10_22=>nx16411, 
      d_arr_mux_10_21=>nx16411, d_arr_mux_10_20=>nx16411, d_arr_mux_10_19=>
      nx16411, d_arr_mux_10_18=>nx16411, d_arr_mux_10_17=>nx16413, 
      d_arr_mux_10_16=>nx16413, d_arr_mux_10_15=>nx16413, d_arr_mux_10_14=>
      ordered_img_data_10_14, d_arr_mux_10_13=>ordered_img_data_10_13, 
      d_arr_mux_10_12=>ordered_img_data_10_12, d_arr_mux_10_11=>
      ordered_img_data_10_11, d_arr_mux_10_10=>ordered_img_data_10_10, 
      d_arr_mux_10_9=>ordered_img_data_10_9, d_arr_mux_10_8=>
      ordered_img_data_10_8, d_arr_mux_10_7=>ordered_img_data_10_7, 
      d_arr_mux_10_6=>ordered_img_data_10_6, d_arr_mux_10_5=>
      ordered_img_data_10_5, d_arr_mux_10_4=>ordered_img_data_10_4, 
      d_arr_mux_10_3=>ordered_img_data_10_3, d_arr_mux_10_2=>
      ordered_img_data_10_2, d_arr_mux_10_1=>ordered_img_data_10_1, 
      d_arr_mux_10_0=>ordered_img_data_10_0, d_arr_mux_11_31=>nx16417, 
      d_arr_mux_11_30=>nx16417, d_arr_mux_11_29=>nx16417, d_arr_mux_11_28=>
      nx16417, d_arr_mux_11_27=>nx16417, d_arr_mux_11_26=>nx16417, 
      d_arr_mux_11_25=>nx16417, d_arr_mux_11_24=>nx16419, d_arr_mux_11_23=>
      nx16419, d_arr_mux_11_22=>nx16419, d_arr_mux_11_21=>nx16419, 
      d_arr_mux_11_20=>nx16419, d_arr_mux_11_19=>nx16419, d_arr_mux_11_18=>
      nx16419, d_arr_mux_11_17=>nx16421, d_arr_mux_11_16=>nx16421, 
      d_arr_mux_11_15=>nx16421, d_arr_mux_11_14=>ordered_img_data_11_14, 
      d_arr_mux_11_13=>ordered_img_data_11_13, d_arr_mux_11_12=>
      ordered_img_data_11_12, d_arr_mux_11_11=>ordered_img_data_11_11, 
      d_arr_mux_11_10=>ordered_img_data_11_10, d_arr_mux_11_9=>
      ordered_img_data_11_9, d_arr_mux_11_8=>ordered_img_data_11_8, 
      d_arr_mux_11_7=>ordered_img_data_11_7, d_arr_mux_11_6=>
      ordered_img_data_11_6, d_arr_mux_11_5=>ordered_img_data_11_5, 
      d_arr_mux_11_4=>ordered_img_data_11_4, d_arr_mux_11_3=>
      ordered_img_data_11_3, d_arr_mux_11_2=>ordered_img_data_11_2, 
      d_arr_mux_11_1=>ordered_img_data_11_1, d_arr_mux_11_0=>
      ordered_img_data_11_0, d_arr_mux_12_31=>nx16425, d_arr_mux_12_30=>
      nx16425, d_arr_mux_12_29=>nx16425, d_arr_mux_12_28=>nx16425, 
      d_arr_mux_12_27=>nx16425, d_arr_mux_12_26=>nx16425, d_arr_mux_12_25=>
      nx16425, d_arr_mux_12_24=>nx16427, d_arr_mux_12_23=>nx16427, 
      d_arr_mux_12_22=>nx16427, d_arr_mux_12_21=>nx16427, d_arr_mux_12_20=>
      nx16427, d_arr_mux_12_19=>nx16427, d_arr_mux_12_18=>nx16427, 
      d_arr_mux_12_17=>nx16429, d_arr_mux_12_16=>nx16429, d_arr_mux_12_15=>
      nx16429, d_arr_mux_12_14=>ordered_img_data_12_14, d_arr_mux_12_13=>
      ordered_img_data_12_13, d_arr_mux_12_12=>ordered_img_data_12_12, 
      d_arr_mux_12_11=>ordered_img_data_12_11, d_arr_mux_12_10=>
      ordered_img_data_12_10, d_arr_mux_12_9=>ordered_img_data_12_9, 
      d_arr_mux_12_8=>ordered_img_data_12_8, d_arr_mux_12_7=>
      ordered_img_data_12_7, d_arr_mux_12_6=>ordered_img_data_12_6, 
      d_arr_mux_12_5=>ordered_img_data_12_5, d_arr_mux_12_4=>
      ordered_img_data_12_4, d_arr_mux_12_3=>ordered_img_data_12_3, 
      d_arr_mux_12_2=>ordered_img_data_12_2, d_arr_mux_12_1=>
      ordered_img_data_12_1, d_arr_mux_12_0=>ordered_img_data_12_0, 
      d_arr_mux_13_31=>nx16433, d_arr_mux_13_30=>nx16433, d_arr_mux_13_29=>
      nx16433, d_arr_mux_13_28=>nx16433, d_arr_mux_13_27=>nx16433, 
      d_arr_mux_13_26=>nx16433, d_arr_mux_13_25=>nx16433, d_arr_mux_13_24=>
      nx16435, d_arr_mux_13_23=>nx16435, d_arr_mux_13_22=>nx16435, 
      d_arr_mux_13_21=>nx16435, d_arr_mux_13_20=>nx16435, d_arr_mux_13_19=>
      nx16435, d_arr_mux_13_18=>nx16435, d_arr_mux_13_17=>nx16437, 
      d_arr_mux_13_16=>nx16437, d_arr_mux_13_15=>nx16437, d_arr_mux_13_14=>
      ordered_img_data_13_14, d_arr_mux_13_13=>ordered_img_data_13_13, 
      d_arr_mux_13_12=>ordered_img_data_13_12, d_arr_mux_13_11=>
      ordered_img_data_13_11, d_arr_mux_13_10=>ordered_img_data_13_10, 
      d_arr_mux_13_9=>ordered_img_data_13_9, d_arr_mux_13_8=>
      ordered_img_data_13_8, d_arr_mux_13_7=>ordered_img_data_13_7, 
      d_arr_mux_13_6=>ordered_img_data_13_6, d_arr_mux_13_5=>
      ordered_img_data_13_5, d_arr_mux_13_4=>ordered_img_data_13_4, 
      d_arr_mux_13_3=>ordered_img_data_13_3, d_arr_mux_13_2=>
      ordered_img_data_13_2, d_arr_mux_13_1=>ordered_img_data_13_1, 
      d_arr_mux_13_0=>ordered_img_data_13_0, d_arr_mux_14_31=>nx16441, 
      d_arr_mux_14_30=>nx16441, d_arr_mux_14_29=>nx16441, d_arr_mux_14_28=>
      nx16441, d_arr_mux_14_27=>nx16441, d_arr_mux_14_26=>nx16441, 
      d_arr_mux_14_25=>nx16441, d_arr_mux_14_24=>nx16443, d_arr_mux_14_23=>
      nx16443, d_arr_mux_14_22=>nx16443, d_arr_mux_14_21=>nx16443, 
      d_arr_mux_14_20=>nx16443, d_arr_mux_14_19=>nx16443, d_arr_mux_14_18=>
      nx16443, d_arr_mux_14_17=>nx16445, d_arr_mux_14_16=>nx16445, 
      d_arr_mux_14_15=>nx16445, d_arr_mux_14_14=>ordered_img_data_14_14, 
      d_arr_mux_14_13=>ordered_img_data_14_13, d_arr_mux_14_12=>
      ordered_img_data_14_12, d_arr_mux_14_11=>ordered_img_data_14_11, 
      d_arr_mux_14_10=>ordered_img_data_14_10, d_arr_mux_14_9=>
      ordered_img_data_14_9, d_arr_mux_14_8=>ordered_img_data_14_8, 
      d_arr_mux_14_7=>ordered_img_data_14_7, d_arr_mux_14_6=>
      ordered_img_data_14_6, d_arr_mux_14_5=>ordered_img_data_14_5, 
      d_arr_mux_14_4=>ordered_img_data_14_4, d_arr_mux_14_3=>
      ordered_img_data_14_3, d_arr_mux_14_2=>ordered_img_data_14_2, 
      d_arr_mux_14_1=>ordered_img_data_14_1, d_arr_mux_14_0=>
      ordered_img_data_14_0, d_arr_mux_15_31=>nx16449, d_arr_mux_15_30=>
      nx16449, d_arr_mux_15_29=>nx16449, d_arr_mux_15_28=>nx16449, 
      d_arr_mux_15_27=>nx16449, d_arr_mux_15_26=>nx16449, d_arr_mux_15_25=>
      nx16449, d_arr_mux_15_24=>nx16451, d_arr_mux_15_23=>nx16451, 
      d_arr_mux_15_22=>nx16451, d_arr_mux_15_21=>nx16451, d_arr_mux_15_20=>
      nx16451, d_arr_mux_15_19=>nx16451, d_arr_mux_15_18=>nx16451, 
      d_arr_mux_15_17=>nx16453, d_arr_mux_15_16=>nx16453, d_arr_mux_15_15=>
      nx16453, d_arr_mux_15_14=>ordered_img_data_15_14, d_arr_mux_15_13=>
      ordered_img_data_15_13, d_arr_mux_15_12=>ordered_img_data_15_12, 
      d_arr_mux_15_11=>ordered_img_data_15_11, d_arr_mux_15_10=>
      ordered_img_data_15_10, d_arr_mux_15_9=>ordered_img_data_15_9, 
      d_arr_mux_15_8=>ordered_img_data_15_8, d_arr_mux_15_7=>
      ordered_img_data_15_7, d_arr_mux_15_6=>ordered_img_data_15_6, 
      d_arr_mux_15_5=>ordered_img_data_15_5, d_arr_mux_15_4=>
      ordered_img_data_15_4, d_arr_mux_15_3=>ordered_img_data_15_3, 
      d_arr_mux_15_2=>ordered_img_data_15_2, d_arr_mux_15_1=>
      ordered_img_data_15_1, d_arr_mux_15_0=>ordered_img_data_15_0, 
      d_arr_mux_16_31=>nx16457, d_arr_mux_16_30=>nx16457, d_arr_mux_16_29=>
      nx16457, d_arr_mux_16_28=>nx16457, d_arr_mux_16_27=>nx16457, 
      d_arr_mux_16_26=>nx16457, d_arr_mux_16_25=>nx16457, d_arr_mux_16_24=>
      nx16459, d_arr_mux_16_23=>nx16459, d_arr_mux_16_22=>nx16459, 
      d_arr_mux_16_21=>nx16459, d_arr_mux_16_20=>nx16459, d_arr_mux_16_19=>
      nx16459, d_arr_mux_16_18=>nx16459, d_arr_mux_16_17=>nx16461, 
      d_arr_mux_16_16=>nx16461, d_arr_mux_16_15=>nx16461, d_arr_mux_16_14=>
      ordered_img_data_16_14, d_arr_mux_16_13=>ordered_img_data_16_13, 
      d_arr_mux_16_12=>ordered_img_data_16_12, d_arr_mux_16_11=>
      ordered_img_data_16_11, d_arr_mux_16_10=>ordered_img_data_16_10, 
      d_arr_mux_16_9=>ordered_img_data_16_9, d_arr_mux_16_8=>
      ordered_img_data_16_8, d_arr_mux_16_7=>ordered_img_data_16_7, 
      d_arr_mux_16_6=>ordered_img_data_16_6, d_arr_mux_16_5=>
      ordered_img_data_16_5, d_arr_mux_16_4=>ordered_img_data_16_4, 
      d_arr_mux_16_3=>ordered_img_data_16_3, d_arr_mux_16_2=>
      ordered_img_data_16_2, d_arr_mux_16_1=>ordered_img_data_16_1, 
      d_arr_mux_16_0=>ordered_img_data_16_0, d_arr_mux_17_31=>nx16465, 
      d_arr_mux_17_30=>nx16465, d_arr_mux_17_29=>nx16465, d_arr_mux_17_28=>
      nx16465, d_arr_mux_17_27=>nx16465, d_arr_mux_17_26=>nx16465, 
      d_arr_mux_17_25=>nx16465, d_arr_mux_17_24=>nx16467, d_arr_mux_17_23=>
      nx16467, d_arr_mux_17_22=>nx16467, d_arr_mux_17_21=>nx16467, 
      d_arr_mux_17_20=>nx16467, d_arr_mux_17_19=>nx16467, d_arr_mux_17_18=>
      nx16467, d_arr_mux_17_17=>nx16469, d_arr_mux_17_16=>nx16469, 
      d_arr_mux_17_15=>nx16469, d_arr_mux_17_14=>ordered_img_data_17_14, 
      d_arr_mux_17_13=>ordered_img_data_17_13, d_arr_mux_17_12=>
      ordered_img_data_17_12, d_arr_mux_17_11=>ordered_img_data_17_11, 
      d_arr_mux_17_10=>ordered_img_data_17_10, d_arr_mux_17_9=>
      ordered_img_data_17_9, d_arr_mux_17_8=>ordered_img_data_17_8, 
      d_arr_mux_17_7=>ordered_img_data_17_7, d_arr_mux_17_6=>
      ordered_img_data_17_6, d_arr_mux_17_5=>ordered_img_data_17_5, 
      d_arr_mux_17_4=>ordered_img_data_17_4, d_arr_mux_17_3=>
      ordered_img_data_17_3, d_arr_mux_17_2=>ordered_img_data_17_2, 
      d_arr_mux_17_1=>ordered_img_data_17_1, d_arr_mux_17_0=>
      ordered_img_data_17_0, d_arr_mux_18_31=>img_data_18_15, 
      d_arr_mux_18_30=>GND0, d_arr_mux_18_29=>GND0, d_arr_mux_18_28=>GND0, 
      d_arr_mux_18_27=>GND0, d_arr_mux_18_26=>GND0, d_arr_mux_18_25=>GND0, 
      d_arr_mux_18_24=>GND0, d_arr_mux_18_23=>GND0, d_arr_mux_18_22=>GND0, 
      d_arr_mux_18_21=>GND0, d_arr_mux_18_20=>GND0, d_arr_mux_18_19=>GND0, 
      d_arr_mux_18_18=>GND0, d_arr_mux_18_17=>GND0, d_arr_mux_18_16=>GND0, 
      d_arr_mux_18_15=>GND0, d_arr_mux_18_14=>nx19438, d_arr_mux_18_13=>
      img_data_18_13, d_arr_mux_18_12=>img_data_18_12, d_arr_mux_18_11=>
      img_data_18_11, d_arr_mux_18_10=>img_data_18_10, d_arr_mux_18_9=>
      img_data_18_9, d_arr_mux_18_8=>img_data_18_8, d_arr_mux_18_7=>
      img_data_18_7, d_arr_mux_18_6=>img_data_18_6, d_arr_mux_18_5=>
      img_data_18_5, d_arr_mux_18_4=>img_data_18_4, d_arr_mux_18_3=>
      img_data_18_3, d_arr_mux_18_2=>img_data_18_2, d_arr_mux_18_1=>
      img_data_18_1, d_arr_mux_18_0=>img_data_18_0, d_arr_mux_19_31=>
      img_data_19_15, d_arr_mux_19_30=>GND0, d_arr_mux_19_29=>GND0, 
      d_arr_mux_19_28=>GND0, d_arr_mux_19_27=>GND0, d_arr_mux_19_26=>GND0, 
      d_arr_mux_19_25=>GND0, d_arr_mux_19_24=>GND0, d_arr_mux_19_23=>GND0, 
      d_arr_mux_19_22=>GND0, d_arr_mux_19_21=>GND0, d_arr_mux_19_20=>GND0, 
      d_arr_mux_19_19=>GND0, d_arr_mux_19_18=>GND0, d_arr_mux_19_17=>GND0, 
      d_arr_mux_19_16=>GND0, d_arr_mux_19_15=>GND0, d_arr_mux_19_14=>
      img_data_19_14, d_arr_mux_19_13=>img_data_19_13, d_arr_mux_19_12=>
      img_data_19_12, d_arr_mux_19_11=>img_data_19_11, d_arr_mux_19_10=>
      img_data_19_10, d_arr_mux_19_9=>img_data_19_9, d_arr_mux_19_8=>
      img_data_19_8, d_arr_mux_19_7=>img_data_19_7, d_arr_mux_19_6=>
      img_data_19_6, d_arr_mux_19_5=>img_data_19_5, d_arr_mux_19_4=>
      img_data_19_4, d_arr_mux_19_3=>img_data_19_3, d_arr_mux_19_2=>
      img_data_19_2, d_arr_mux_19_1=>img_data_19_1, d_arr_mux_19_0=>
      img_data_19_0, d_arr_mux_20_31=>img_data_20_15, d_arr_mux_20_30=>GND0, 
      d_arr_mux_20_29=>GND0, d_arr_mux_20_28=>GND0, d_arr_mux_20_27=>GND0, 
      d_arr_mux_20_26=>GND0, d_arr_mux_20_25=>GND0, d_arr_mux_20_24=>GND0, 
      d_arr_mux_20_23=>GND0, d_arr_mux_20_22=>GND0, d_arr_mux_20_21=>GND0, 
      d_arr_mux_20_20=>GND0, d_arr_mux_20_19=>GND0, d_arr_mux_20_18=>GND0, 
      d_arr_mux_20_17=>GND0, d_arr_mux_20_16=>GND0, d_arr_mux_20_15=>GND0, 
      d_arr_mux_20_14=>nx19440, d_arr_mux_20_13=>img_data_20_13, 
      d_arr_mux_20_12=>img_data_20_12, d_arr_mux_20_11=>img_data_20_11, 
      d_arr_mux_20_10=>img_data_20_10, d_arr_mux_20_9=>img_data_20_9, 
      d_arr_mux_20_8=>img_data_20_8, d_arr_mux_20_7=>img_data_20_7, 
      d_arr_mux_20_6=>img_data_20_6, d_arr_mux_20_5=>img_data_20_5, 
      d_arr_mux_20_4=>img_data_20_4, d_arr_mux_20_3=>img_data_20_3, 
      d_arr_mux_20_2=>img_data_20_2, d_arr_mux_20_1=>img_data_20_1, 
      d_arr_mux_20_0=>img_data_20_0, d_arr_mux_21_31=>img_data_21_15, 
      d_arr_mux_21_30=>GND0, d_arr_mux_21_29=>GND0, d_arr_mux_21_28=>GND0, 
      d_arr_mux_21_27=>GND0, d_arr_mux_21_26=>GND0, d_arr_mux_21_25=>GND0, 
      d_arr_mux_21_24=>GND0, d_arr_mux_21_23=>GND0, d_arr_mux_21_22=>GND0, 
      d_arr_mux_21_21=>GND0, d_arr_mux_21_20=>GND0, d_arr_mux_21_19=>GND0, 
      d_arr_mux_21_18=>GND0, d_arr_mux_21_17=>GND0, d_arr_mux_21_16=>GND0, 
      d_arr_mux_21_15=>GND0, d_arr_mux_21_14=>nx19442, d_arr_mux_21_13=>
      img_data_21_13, d_arr_mux_21_12=>img_data_21_12, d_arr_mux_21_11=>
      img_data_21_11, d_arr_mux_21_10=>img_data_21_10, d_arr_mux_21_9=>
      img_data_21_9, d_arr_mux_21_8=>img_data_21_8, d_arr_mux_21_7=>
      img_data_21_7, d_arr_mux_21_6=>img_data_21_6, d_arr_mux_21_5=>
      img_data_21_5, d_arr_mux_21_4=>img_data_21_4, d_arr_mux_21_3=>
      img_data_21_3, d_arr_mux_21_2=>img_data_21_2, d_arr_mux_21_1=>
      img_data_21_1, d_arr_mux_21_0=>img_data_21_0, d_arr_mux_22_31=>
      img_data_22_15, d_arr_mux_22_30=>GND0, d_arr_mux_22_29=>GND0, 
      d_arr_mux_22_28=>GND0, d_arr_mux_22_27=>GND0, d_arr_mux_22_26=>GND0, 
      d_arr_mux_22_25=>GND0, d_arr_mux_22_24=>GND0, d_arr_mux_22_23=>GND0, 
      d_arr_mux_22_22=>GND0, d_arr_mux_22_21=>GND0, d_arr_mux_22_20=>GND0, 
      d_arr_mux_22_19=>GND0, d_arr_mux_22_18=>GND0, d_arr_mux_22_17=>GND0, 
      d_arr_mux_22_16=>GND0, d_arr_mux_22_15=>GND0, d_arr_mux_22_14=>nx19444, 
      d_arr_mux_22_13=>img_data_22_13, d_arr_mux_22_12=>img_data_22_12, 
      d_arr_mux_22_11=>img_data_22_11, d_arr_mux_22_10=>img_data_22_10, 
      d_arr_mux_22_9=>img_data_22_9, d_arr_mux_22_8=>img_data_22_8, 
      d_arr_mux_22_7=>img_data_22_7, d_arr_mux_22_6=>img_data_22_6, 
      d_arr_mux_22_5=>img_data_22_5, d_arr_mux_22_4=>img_data_22_4, 
      d_arr_mux_22_3=>img_data_22_3, d_arr_mux_22_2=>img_data_22_2, 
      d_arr_mux_22_1=>img_data_22_1, d_arr_mux_22_0=>img_data_22_0, 
      d_arr_mux_23_31=>img_data_23_15, d_arr_mux_23_30=>GND0, 
      d_arr_mux_23_29=>GND0, d_arr_mux_23_28=>GND0, d_arr_mux_23_27=>GND0, 
      d_arr_mux_23_26=>GND0, d_arr_mux_23_25=>GND0, d_arr_mux_23_24=>GND0, 
      d_arr_mux_23_23=>GND0, d_arr_mux_23_22=>GND0, d_arr_mux_23_21=>GND0, 
      d_arr_mux_23_20=>GND0, d_arr_mux_23_19=>GND0, d_arr_mux_23_18=>GND0, 
      d_arr_mux_23_17=>GND0, d_arr_mux_23_16=>GND0, d_arr_mux_23_15=>GND0, 
      d_arr_mux_23_14=>nx19446, d_arr_mux_23_13=>img_data_23_13, 
      d_arr_mux_23_12=>img_data_23_12, d_arr_mux_23_11=>img_data_23_11, 
      d_arr_mux_23_10=>img_data_23_10, d_arr_mux_23_9=>img_data_23_9, 
      d_arr_mux_23_8=>img_data_23_8, d_arr_mux_23_7=>img_data_23_7, 
      d_arr_mux_23_6=>img_data_23_6, d_arr_mux_23_5=>img_data_23_5, 
      d_arr_mux_23_4=>img_data_23_4, d_arr_mux_23_3=>img_data_23_3, 
      d_arr_mux_23_2=>img_data_23_2, d_arr_mux_23_1=>img_data_23_1, 
      d_arr_mux_23_0=>img_data_23_0, d_arr_mux_24_31=>img_data_24_15, 
      d_arr_mux_24_30=>GND0, d_arr_mux_24_29=>GND0, d_arr_mux_24_28=>GND0, 
      d_arr_mux_24_27=>GND0, d_arr_mux_24_26=>GND0, d_arr_mux_24_25=>GND0, 
      d_arr_mux_24_24=>GND0, d_arr_mux_24_23=>GND0, d_arr_mux_24_22=>GND0, 
      d_arr_mux_24_21=>GND0, d_arr_mux_24_20=>GND0, d_arr_mux_24_19=>GND0, 
      d_arr_mux_24_18=>GND0, d_arr_mux_24_17=>GND0, d_arr_mux_24_16=>GND0, 
      d_arr_mux_24_15=>GND0, d_arr_mux_24_14=>img_data_24_14, 
      d_arr_mux_24_13=>img_data_24_13, d_arr_mux_24_12=>img_data_24_12, 
      d_arr_mux_24_11=>img_data_24_11, d_arr_mux_24_10=>img_data_24_10, 
      d_arr_mux_24_9=>img_data_24_9, d_arr_mux_24_8=>img_data_24_8, 
      d_arr_mux_24_7=>img_data_24_7, d_arr_mux_24_6=>img_data_24_6, 
      d_arr_mux_24_5=>img_data_24_5, d_arr_mux_24_4=>img_data_24_4, 
      d_arr_mux_24_3=>img_data_24_3, d_arr_mux_24_2=>img_data_24_2, 
      d_arr_mux_24_1=>img_data_24_1, d_arr_mux_24_0=>img_data_24_0, 
      d_arr_mul_0_31=>d_arr_mul_0_31, d_arr_mul_0_30=>d_arr_mul_0_30, 
      d_arr_mul_0_29=>d_arr_mul_0_29, d_arr_mul_0_28=>d_arr_mul_0_28, 
      d_arr_mul_0_27=>d_arr_mul_0_27, d_arr_mul_0_26=>d_arr_mul_0_26, 
      d_arr_mul_0_25=>d_arr_mul_0_25, d_arr_mul_0_24=>d_arr_mul_0_24, 
      d_arr_mul_0_23=>d_arr_mul_0_23, d_arr_mul_0_22=>d_arr_mul_0_22, 
      d_arr_mul_0_21=>d_arr_mul_0_21, d_arr_mul_0_20=>d_arr_mul_0_20, 
      d_arr_mul_0_19=>d_arr_mul_0_19, d_arr_mul_0_18=>d_arr_mul_0_18, 
      d_arr_mul_0_17=>d_arr_mul_0_17, d_arr_mul_0_16=>d_arr_mul_0_16, 
      d_arr_mul_0_15=>d_arr_mul_0_15, d_arr_mul_0_14=>d_arr_mul_0_14, 
      d_arr_mul_0_13=>d_arr_mul_0_13, d_arr_mul_0_12=>d_arr_mul_0_12, 
      d_arr_mul_0_11=>d_arr_mul_0_11, d_arr_mul_0_10=>d_arr_mul_0_10, 
      d_arr_mul_0_9=>d_arr_mul_0_9, d_arr_mul_0_8=>d_arr_mul_0_8, 
      d_arr_mul_0_7=>d_arr_mul_0_7, d_arr_mul_0_6=>d_arr_mul_0_6, 
      d_arr_mul_0_5=>d_arr_mul_0_5, d_arr_mul_0_4=>d_arr_mul_0_4, 
      d_arr_mul_0_3=>d_arr_mul_0_3, d_arr_mul_0_2=>d_arr_mul_0_2, 
      d_arr_mul_0_1=>d_arr_mul_0_1, d_arr_mul_0_0=>d_arr_mul_0_0, 
      d_arr_mul_1_31=>d_arr_mul_1_31, d_arr_mul_1_30=>d_arr_mul_1_30, 
      d_arr_mul_1_29=>d_arr_mul_1_29, d_arr_mul_1_28=>d_arr_mul_1_28, 
      d_arr_mul_1_27=>d_arr_mul_1_27, d_arr_mul_1_26=>d_arr_mul_1_26, 
      d_arr_mul_1_25=>d_arr_mul_1_25, d_arr_mul_1_24=>d_arr_mul_1_24, 
      d_arr_mul_1_23=>d_arr_mul_1_23, d_arr_mul_1_22=>d_arr_mul_1_22, 
      d_arr_mul_1_21=>d_arr_mul_1_21, d_arr_mul_1_20=>d_arr_mul_1_20, 
      d_arr_mul_1_19=>d_arr_mul_1_19, d_arr_mul_1_18=>d_arr_mul_1_18, 
      d_arr_mul_1_17=>d_arr_mul_1_17, d_arr_mul_1_16=>d_arr_mul_1_16, 
      d_arr_mul_1_15=>d_arr_mul_1_15, d_arr_mul_1_14=>d_arr_mul_1_14, 
      d_arr_mul_1_13=>d_arr_mul_1_13, d_arr_mul_1_12=>d_arr_mul_1_12, 
      d_arr_mul_1_11=>d_arr_mul_1_11, d_arr_mul_1_10=>d_arr_mul_1_10, 
      d_arr_mul_1_9=>d_arr_mul_1_9, d_arr_mul_1_8=>d_arr_mul_1_8, 
      d_arr_mul_1_7=>d_arr_mul_1_7, d_arr_mul_1_6=>d_arr_mul_1_6, 
      d_arr_mul_1_5=>d_arr_mul_1_5, d_arr_mul_1_4=>d_arr_mul_1_4, 
      d_arr_mul_1_3=>d_arr_mul_1_3, d_arr_mul_1_2=>d_arr_mul_1_2, 
      d_arr_mul_1_1=>d_arr_mul_1_1, d_arr_mul_1_0=>d_arr_mul_1_0, 
      d_arr_mul_2_31=>d_arr_mul_2_31, d_arr_mul_2_30=>d_arr_mul_2_30, 
      d_arr_mul_2_29=>d_arr_mul_2_29, d_arr_mul_2_28=>d_arr_mul_2_28, 
      d_arr_mul_2_27=>d_arr_mul_2_27, d_arr_mul_2_26=>d_arr_mul_2_26, 
      d_arr_mul_2_25=>d_arr_mul_2_25, d_arr_mul_2_24=>d_arr_mul_2_24, 
      d_arr_mul_2_23=>d_arr_mul_2_23, d_arr_mul_2_22=>d_arr_mul_2_22, 
      d_arr_mul_2_21=>d_arr_mul_2_21, d_arr_mul_2_20=>d_arr_mul_2_20, 
      d_arr_mul_2_19=>d_arr_mul_2_19, d_arr_mul_2_18=>d_arr_mul_2_18, 
      d_arr_mul_2_17=>d_arr_mul_2_17, d_arr_mul_2_16=>d_arr_mul_2_16, 
      d_arr_mul_2_15=>d_arr_mul_2_15, d_arr_mul_2_14=>d_arr_mul_2_14, 
      d_arr_mul_2_13=>d_arr_mul_2_13, d_arr_mul_2_12=>d_arr_mul_2_12, 
      d_arr_mul_2_11=>d_arr_mul_2_11, d_arr_mul_2_10=>d_arr_mul_2_10, 
      d_arr_mul_2_9=>d_arr_mul_2_9, d_arr_mul_2_8=>d_arr_mul_2_8, 
      d_arr_mul_2_7=>d_arr_mul_2_7, d_arr_mul_2_6=>d_arr_mul_2_6, 
      d_arr_mul_2_5=>d_arr_mul_2_5, d_arr_mul_2_4=>d_arr_mul_2_4, 
      d_arr_mul_2_3=>d_arr_mul_2_3, d_arr_mul_2_2=>d_arr_mul_2_2, 
      d_arr_mul_2_1=>d_arr_mul_2_1, d_arr_mul_2_0=>d_arr_mul_2_0, 
      d_arr_mul_3_31=>d_arr_mul_3_31, d_arr_mul_3_30=>d_arr_mul_3_30, 
      d_arr_mul_3_29=>d_arr_mul_3_29, d_arr_mul_3_28=>d_arr_mul_3_28, 
      d_arr_mul_3_27=>d_arr_mul_3_27, d_arr_mul_3_26=>d_arr_mul_3_26, 
      d_arr_mul_3_25=>d_arr_mul_3_25, d_arr_mul_3_24=>d_arr_mul_3_24, 
      d_arr_mul_3_23=>d_arr_mul_3_23, d_arr_mul_3_22=>d_arr_mul_3_22, 
      d_arr_mul_3_21=>d_arr_mul_3_21, d_arr_mul_3_20=>d_arr_mul_3_20, 
      d_arr_mul_3_19=>d_arr_mul_3_19, d_arr_mul_3_18=>d_arr_mul_3_18, 
      d_arr_mul_3_17=>d_arr_mul_3_17, d_arr_mul_3_16=>d_arr_mul_3_16, 
      d_arr_mul_3_15=>d_arr_mul_3_15, d_arr_mul_3_14=>d_arr_mul_3_14, 
      d_arr_mul_3_13=>d_arr_mul_3_13, d_arr_mul_3_12=>d_arr_mul_3_12, 
      d_arr_mul_3_11=>d_arr_mul_3_11, d_arr_mul_3_10=>d_arr_mul_3_10, 
      d_arr_mul_3_9=>d_arr_mul_3_9, d_arr_mul_3_8=>d_arr_mul_3_8, 
      d_arr_mul_3_7=>d_arr_mul_3_7, d_arr_mul_3_6=>d_arr_mul_3_6, 
      d_arr_mul_3_5=>d_arr_mul_3_5, d_arr_mul_3_4=>d_arr_mul_3_4, 
      d_arr_mul_3_3=>d_arr_mul_3_3, d_arr_mul_3_2=>d_arr_mul_3_2, 
      d_arr_mul_3_1=>d_arr_mul_3_1, d_arr_mul_3_0=>d_arr_mul_3_0, 
      d_arr_mul_4_31=>d_arr_mul_4_31, d_arr_mul_4_30=>d_arr_mul_4_30, 
      d_arr_mul_4_29=>d_arr_mul_4_29, d_arr_mul_4_28=>d_arr_mul_4_28, 
      d_arr_mul_4_27=>d_arr_mul_4_27, d_arr_mul_4_26=>d_arr_mul_4_26, 
      d_arr_mul_4_25=>d_arr_mul_4_25, d_arr_mul_4_24=>d_arr_mul_4_24, 
      d_arr_mul_4_23=>d_arr_mul_4_23, d_arr_mul_4_22=>d_arr_mul_4_22, 
      d_arr_mul_4_21=>d_arr_mul_4_21, d_arr_mul_4_20=>d_arr_mul_4_20, 
      d_arr_mul_4_19=>d_arr_mul_4_19, d_arr_mul_4_18=>d_arr_mul_4_18, 
      d_arr_mul_4_17=>d_arr_mul_4_17, d_arr_mul_4_16=>d_arr_mul_4_16, 
      d_arr_mul_4_15=>d_arr_mul_4_15, d_arr_mul_4_14=>d_arr_mul_4_14, 
      d_arr_mul_4_13=>d_arr_mul_4_13, d_arr_mul_4_12=>d_arr_mul_4_12, 
      d_arr_mul_4_11=>d_arr_mul_4_11, d_arr_mul_4_10=>d_arr_mul_4_10, 
      d_arr_mul_4_9=>d_arr_mul_4_9, d_arr_mul_4_8=>d_arr_mul_4_8, 
      d_arr_mul_4_7=>d_arr_mul_4_7, d_arr_mul_4_6=>d_arr_mul_4_6, 
      d_arr_mul_4_5=>d_arr_mul_4_5, d_arr_mul_4_4=>d_arr_mul_4_4, 
      d_arr_mul_4_3=>d_arr_mul_4_3, d_arr_mul_4_2=>d_arr_mul_4_2, 
      d_arr_mul_4_1=>d_arr_mul_4_1, d_arr_mul_4_0=>d_arr_mul_4_0, 
      d_arr_mul_5_31=>d_arr_mul_5_31, d_arr_mul_5_30=>d_arr_mul_5_30, 
      d_arr_mul_5_29=>d_arr_mul_5_29, d_arr_mul_5_28=>d_arr_mul_5_28, 
      d_arr_mul_5_27=>d_arr_mul_5_27, d_arr_mul_5_26=>d_arr_mul_5_26, 
      d_arr_mul_5_25=>d_arr_mul_5_25, d_arr_mul_5_24=>d_arr_mul_5_24, 
      d_arr_mul_5_23=>d_arr_mul_5_23, d_arr_mul_5_22=>d_arr_mul_5_22, 
      d_arr_mul_5_21=>d_arr_mul_5_21, d_arr_mul_5_20=>d_arr_mul_5_20, 
      d_arr_mul_5_19=>d_arr_mul_5_19, d_arr_mul_5_18=>d_arr_mul_5_18, 
      d_arr_mul_5_17=>d_arr_mul_5_17, d_arr_mul_5_16=>d_arr_mul_5_16, 
      d_arr_mul_5_15=>d_arr_mul_5_15, d_arr_mul_5_14=>d_arr_mul_5_14, 
      d_arr_mul_5_13=>d_arr_mul_5_13, d_arr_mul_5_12=>d_arr_mul_5_12, 
      d_arr_mul_5_11=>d_arr_mul_5_11, d_arr_mul_5_10=>d_arr_mul_5_10, 
      d_arr_mul_5_9=>d_arr_mul_5_9, d_arr_mul_5_8=>d_arr_mul_5_8, 
      d_arr_mul_5_7=>d_arr_mul_5_7, d_arr_mul_5_6=>d_arr_mul_5_6, 
      d_arr_mul_5_5=>d_arr_mul_5_5, d_arr_mul_5_4=>d_arr_mul_5_4, 
      d_arr_mul_5_3=>d_arr_mul_5_3, d_arr_mul_5_2=>d_arr_mul_5_2, 
      d_arr_mul_5_1=>d_arr_mul_5_1, d_arr_mul_5_0=>d_arr_mul_5_0, 
      d_arr_mul_6_31=>d_arr_mul_6_31, d_arr_mul_6_30=>d_arr_mul_6_30, 
      d_arr_mul_6_29=>d_arr_mul_6_29, d_arr_mul_6_28=>d_arr_mul_6_28, 
      d_arr_mul_6_27=>d_arr_mul_6_27, d_arr_mul_6_26=>d_arr_mul_6_26, 
      d_arr_mul_6_25=>d_arr_mul_6_25, d_arr_mul_6_24=>d_arr_mul_6_24, 
      d_arr_mul_6_23=>d_arr_mul_6_23, d_arr_mul_6_22=>d_arr_mul_6_22, 
      d_arr_mul_6_21=>d_arr_mul_6_21, d_arr_mul_6_20=>d_arr_mul_6_20, 
      d_arr_mul_6_19=>d_arr_mul_6_19, d_arr_mul_6_18=>d_arr_mul_6_18, 
      d_arr_mul_6_17=>d_arr_mul_6_17, d_arr_mul_6_16=>d_arr_mul_6_16, 
      d_arr_mul_6_15=>d_arr_mul_6_15, d_arr_mul_6_14=>d_arr_mul_6_14, 
      d_arr_mul_6_13=>d_arr_mul_6_13, d_arr_mul_6_12=>d_arr_mul_6_12, 
      d_arr_mul_6_11=>d_arr_mul_6_11, d_arr_mul_6_10=>d_arr_mul_6_10, 
      d_arr_mul_6_9=>d_arr_mul_6_9, d_arr_mul_6_8=>d_arr_mul_6_8, 
      d_arr_mul_6_7=>d_arr_mul_6_7, d_arr_mul_6_6=>d_arr_mul_6_6, 
      d_arr_mul_6_5=>d_arr_mul_6_5, d_arr_mul_6_4=>d_arr_mul_6_4, 
      d_arr_mul_6_3=>d_arr_mul_6_3, d_arr_mul_6_2=>d_arr_mul_6_2, 
      d_arr_mul_6_1=>d_arr_mul_6_1, d_arr_mul_6_0=>d_arr_mul_6_0, 
      d_arr_mul_7_31=>d_arr_mul_7_31, d_arr_mul_7_30=>d_arr_mul_7_30, 
      d_arr_mul_7_29=>d_arr_mul_7_29, d_arr_mul_7_28=>d_arr_mul_7_28, 
      d_arr_mul_7_27=>d_arr_mul_7_27, d_arr_mul_7_26=>d_arr_mul_7_26, 
      d_arr_mul_7_25=>d_arr_mul_7_25, d_arr_mul_7_24=>d_arr_mul_7_24, 
      d_arr_mul_7_23=>d_arr_mul_7_23, d_arr_mul_7_22=>d_arr_mul_7_22, 
      d_arr_mul_7_21=>d_arr_mul_7_21, d_arr_mul_7_20=>d_arr_mul_7_20, 
      d_arr_mul_7_19=>d_arr_mul_7_19, d_arr_mul_7_18=>d_arr_mul_7_18, 
      d_arr_mul_7_17=>d_arr_mul_7_17, d_arr_mul_7_16=>d_arr_mul_7_16, 
      d_arr_mul_7_15=>d_arr_mul_7_15, d_arr_mul_7_14=>d_arr_mul_7_14, 
      d_arr_mul_7_13=>d_arr_mul_7_13, d_arr_mul_7_12=>d_arr_mul_7_12, 
      d_arr_mul_7_11=>d_arr_mul_7_11, d_arr_mul_7_10=>d_arr_mul_7_10, 
      d_arr_mul_7_9=>d_arr_mul_7_9, d_arr_mul_7_8=>d_arr_mul_7_8, 
      d_arr_mul_7_7=>d_arr_mul_7_7, d_arr_mul_7_6=>d_arr_mul_7_6, 
      d_arr_mul_7_5=>d_arr_mul_7_5, d_arr_mul_7_4=>d_arr_mul_7_4, 
      d_arr_mul_7_3=>d_arr_mul_7_3, d_arr_mul_7_2=>d_arr_mul_7_2, 
      d_arr_mul_7_1=>d_arr_mul_7_1, d_arr_mul_7_0=>d_arr_mul_7_0, 
      d_arr_mul_8_31=>d_arr_mul_8_31, d_arr_mul_8_30=>d_arr_mul_8_30, 
      d_arr_mul_8_29=>d_arr_mul_8_29, d_arr_mul_8_28=>d_arr_mul_8_28, 
      d_arr_mul_8_27=>d_arr_mul_8_27, d_arr_mul_8_26=>d_arr_mul_8_26, 
      d_arr_mul_8_25=>d_arr_mul_8_25, d_arr_mul_8_24=>d_arr_mul_8_24, 
      d_arr_mul_8_23=>d_arr_mul_8_23, d_arr_mul_8_22=>d_arr_mul_8_22, 
      d_arr_mul_8_21=>d_arr_mul_8_21, d_arr_mul_8_20=>d_arr_mul_8_20, 
      d_arr_mul_8_19=>d_arr_mul_8_19, d_arr_mul_8_18=>d_arr_mul_8_18, 
      d_arr_mul_8_17=>d_arr_mul_8_17, d_arr_mul_8_16=>d_arr_mul_8_16, 
      d_arr_mul_8_15=>d_arr_mul_8_15, d_arr_mul_8_14=>d_arr_mul_8_14, 
      d_arr_mul_8_13=>d_arr_mul_8_13, d_arr_mul_8_12=>d_arr_mul_8_12, 
      d_arr_mul_8_11=>d_arr_mul_8_11, d_arr_mul_8_10=>d_arr_mul_8_10, 
      d_arr_mul_8_9=>d_arr_mul_8_9, d_arr_mul_8_8=>d_arr_mul_8_8, 
      d_arr_mul_8_7=>d_arr_mul_8_7, d_arr_mul_8_6=>d_arr_mul_8_6, 
      d_arr_mul_8_5=>d_arr_mul_8_5, d_arr_mul_8_4=>d_arr_mul_8_4, 
      d_arr_mul_8_3=>d_arr_mul_8_3, d_arr_mul_8_2=>d_arr_mul_8_2, 
      d_arr_mul_8_1=>d_arr_mul_8_1, d_arr_mul_8_0=>d_arr_mul_8_0, 
      d_arr_mul_9_31=>d_arr_mul_9_31, d_arr_mul_9_30=>d_arr_mul_9_30, 
      d_arr_mul_9_29=>d_arr_mul_9_29, d_arr_mul_9_28=>d_arr_mul_9_28, 
      d_arr_mul_9_27=>d_arr_mul_9_27, d_arr_mul_9_26=>d_arr_mul_9_26, 
      d_arr_mul_9_25=>d_arr_mul_9_25, d_arr_mul_9_24=>d_arr_mul_9_24, 
      d_arr_mul_9_23=>d_arr_mul_9_23, d_arr_mul_9_22=>d_arr_mul_9_22, 
      d_arr_mul_9_21=>d_arr_mul_9_21, d_arr_mul_9_20=>d_arr_mul_9_20, 
      d_arr_mul_9_19=>d_arr_mul_9_19, d_arr_mul_9_18=>d_arr_mul_9_18, 
      d_arr_mul_9_17=>d_arr_mul_9_17, d_arr_mul_9_16=>d_arr_mul_9_16, 
      d_arr_mul_9_15=>d_arr_mul_9_15, d_arr_mul_9_14=>d_arr_mul_9_14, 
      d_arr_mul_9_13=>d_arr_mul_9_13, d_arr_mul_9_12=>d_arr_mul_9_12, 
      d_arr_mul_9_11=>d_arr_mul_9_11, d_arr_mul_9_10=>d_arr_mul_9_10, 
      d_arr_mul_9_9=>d_arr_mul_9_9, d_arr_mul_9_8=>d_arr_mul_9_8, 
      d_arr_mul_9_7=>d_arr_mul_9_7, d_arr_mul_9_6=>d_arr_mul_9_6, 
      d_arr_mul_9_5=>d_arr_mul_9_5, d_arr_mul_9_4=>d_arr_mul_9_4, 
      d_arr_mul_9_3=>d_arr_mul_9_3, d_arr_mul_9_2=>d_arr_mul_9_2, 
      d_arr_mul_9_1=>d_arr_mul_9_1, d_arr_mul_9_0=>d_arr_mul_9_0, 
      d_arr_mul_10_31=>d_arr_mul_10_31, d_arr_mul_10_30=>d_arr_mul_10_30, 
      d_arr_mul_10_29=>d_arr_mul_10_29, d_arr_mul_10_28=>d_arr_mul_10_28, 
      d_arr_mul_10_27=>d_arr_mul_10_27, d_arr_mul_10_26=>d_arr_mul_10_26, 
      d_arr_mul_10_25=>d_arr_mul_10_25, d_arr_mul_10_24=>d_arr_mul_10_24, 
      d_arr_mul_10_23=>d_arr_mul_10_23, d_arr_mul_10_22=>d_arr_mul_10_22, 
      d_arr_mul_10_21=>d_arr_mul_10_21, d_arr_mul_10_20=>d_arr_mul_10_20, 
      d_arr_mul_10_19=>d_arr_mul_10_19, d_arr_mul_10_18=>d_arr_mul_10_18, 
      d_arr_mul_10_17=>d_arr_mul_10_17, d_arr_mul_10_16=>d_arr_mul_10_16, 
      d_arr_mul_10_15=>d_arr_mul_10_15, d_arr_mul_10_14=>d_arr_mul_10_14, 
      d_arr_mul_10_13=>d_arr_mul_10_13, d_arr_mul_10_12=>d_arr_mul_10_12, 
      d_arr_mul_10_11=>d_arr_mul_10_11, d_arr_mul_10_10=>d_arr_mul_10_10, 
      d_arr_mul_10_9=>d_arr_mul_10_9, d_arr_mul_10_8=>d_arr_mul_10_8, 
      d_arr_mul_10_7=>d_arr_mul_10_7, d_arr_mul_10_6=>d_arr_mul_10_6, 
      d_arr_mul_10_5=>d_arr_mul_10_5, d_arr_mul_10_4=>d_arr_mul_10_4, 
      d_arr_mul_10_3=>d_arr_mul_10_3, d_arr_mul_10_2=>d_arr_mul_10_2, 
      d_arr_mul_10_1=>d_arr_mul_10_1, d_arr_mul_10_0=>d_arr_mul_10_0, 
      d_arr_mul_11_31=>d_arr_mul_11_31, d_arr_mul_11_30=>d_arr_mul_11_30, 
      d_arr_mul_11_29=>d_arr_mul_11_29, d_arr_mul_11_28=>d_arr_mul_11_28, 
      d_arr_mul_11_27=>d_arr_mul_11_27, d_arr_mul_11_26=>d_arr_mul_11_26, 
      d_arr_mul_11_25=>d_arr_mul_11_25, d_arr_mul_11_24=>d_arr_mul_11_24, 
      d_arr_mul_11_23=>d_arr_mul_11_23, d_arr_mul_11_22=>d_arr_mul_11_22, 
      d_arr_mul_11_21=>d_arr_mul_11_21, d_arr_mul_11_20=>d_arr_mul_11_20, 
      d_arr_mul_11_19=>d_arr_mul_11_19, d_arr_mul_11_18=>d_arr_mul_11_18, 
      d_arr_mul_11_17=>d_arr_mul_11_17, d_arr_mul_11_16=>d_arr_mul_11_16, 
      d_arr_mul_11_15=>d_arr_mul_11_15, d_arr_mul_11_14=>d_arr_mul_11_14, 
      d_arr_mul_11_13=>d_arr_mul_11_13, d_arr_mul_11_12=>d_arr_mul_11_12, 
      d_arr_mul_11_11=>d_arr_mul_11_11, d_arr_mul_11_10=>d_arr_mul_11_10, 
      d_arr_mul_11_9=>d_arr_mul_11_9, d_arr_mul_11_8=>d_arr_mul_11_8, 
      d_arr_mul_11_7=>d_arr_mul_11_7, d_arr_mul_11_6=>d_arr_mul_11_6, 
      d_arr_mul_11_5=>d_arr_mul_11_5, d_arr_mul_11_4=>d_arr_mul_11_4, 
      d_arr_mul_11_3=>d_arr_mul_11_3, d_arr_mul_11_2=>d_arr_mul_11_2, 
      d_arr_mul_11_1=>d_arr_mul_11_1, d_arr_mul_11_0=>d_arr_mul_11_0, 
      d_arr_mul_12_31=>d_arr_mul_12_31, d_arr_mul_12_30=>d_arr_mul_12_30, 
      d_arr_mul_12_29=>d_arr_mul_12_29, d_arr_mul_12_28=>d_arr_mul_12_28, 
      d_arr_mul_12_27=>d_arr_mul_12_27, d_arr_mul_12_26=>d_arr_mul_12_26, 
      d_arr_mul_12_25=>d_arr_mul_12_25, d_arr_mul_12_24=>d_arr_mul_12_24, 
      d_arr_mul_12_23=>d_arr_mul_12_23, d_arr_mul_12_22=>d_arr_mul_12_22, 
      d_arr_mul_12_21=>d_arr_mul_12_21, d_arr_mul_12_20=>d_arr_mul_12_20, 
      d_arr_mul_12_19=>d_arr_mul_12_19, d_arr_mul_12_18=>d_arr_mul_12_18, 
      d_arr_mul_12_17=>d_arr_mul_12_17, d_arr_mul_12_16=>d_arr_mul_12_16, 
      d_arr_mul_12_15=>d_arr_mul_12_15, d_arr_mul_12_14=>d_arr_mul_12_14, 
      d_arr_mul_12_13=>d_arr_mul_12_13, d_arr_mul_12_12=>d_arr_mul_12_12, 
      d_arr_mul_12_11=>d_arr_mul_12_11, d_arr_mul_12_10=>d_arr_mul_12_10, 
      d_arr_mul_12_9=>d_arr_mul_12_9, d_arr_mul_12_8=>d_arr_mul_12_8, 
      d_arr_mul_12_7=>d_arr_mul_12_7, d_arr_mul_12_6=>d_arr_mul_12_6, 
      d_arr_mul_12_5=>d_arr_mul_12_5, d_arr_mul_12_4=>d_arr_mul_12_4, 
      d_arr_mul_12_3=>d_arr_mul_12_3, d_arr_mul_12_2=>d_arr_mul_12_2, 
      d_arr_mul_12_1=>d_arr_mul_12_1, d_arr_mul_12_0=>d_arr_mul_12_0, 
      d_arr_mul_13_31=>d_arr_mul_13_31, d_arr_mul_13_30=>d_arr_mul_13_30, 
      d_arr_mul_13_29=>d_arr_mul_13_29, d_arr_mul_13_28=>d_arr_mul_13_28, 
      d_arr_mul_13_27=>d_arr_mul_13_27, d_arr_mul_13_26=>d_arr_mul_13_26, 
      d_arr_mul_13_25=>d_arr_mul_13_25, d_arr_mul_13_24=>d_arr_mul_13_24, 
      d_arr_mul_13_23=>d_arr_mul_13_23, d_arr_mul_13_22=>d_arr_mul_13_22, 
      d_arr_mul_13_21=>d_arr_mul_13_21, d_arr_mul_13_20=>d_arr_mul_13_20, 
      d_arr_mul_13_19=>d_arr_mul_13_19, d_arr_mul_13_18=>d_arr_mul_13_18, 
      d_arr_mul_13_17=>d_arr_mul_13_17, d_arr_mul_13_16=>d_arr_mul_13_16, 
      d_arr_mul_13_15=>d_arr_mul_13_15, d_arr_mul_13_14=>d_arr_mul_13_14, 
      d_arr_mul_13_13=>d_arr_mul_13_13, d_arr_mul_13_12=>d_arr_mul_13_12, 
      d_arr_mul_13_11=>d_arr_mul_13_11, d_arr_mul_13_10=>d_arr_mul_13_10, 
      d_arr_mul_13_9=>d_arr_mul_13_9, d_arr_mul_13_8=>d_arr_mul_13_8, 
      d_arr_mul_13_7=>d_arr_mul_13_7, d_arr_mul_13_6=>d_arr_mul_13_6, 
      d_arr_mul_13_5=>d_arr_mul_13_5, d_arr_mul_13_4=>d_arr_mul_13_4, 
      d_arr_mul_13_3=>d_arr_mul_13_3, d_arr_mul_13_2=>d_arr_mul_13_2, 
      d_arr_mul_13_1=>d_arr_mul_13_1, d_arr_mul_13_0=>d_arr_mul_13_0, 
      d_arr_mul_14_31=>d_arr_mul_14_31, d_arr_mul_14_30=>d_arr_mul_14_30, 
      d_arr_mul_14_29=>d_arr_mul_14_29, d_arr_mul_14_28=>d_arr_mul_14_28, 
      d_arr_mul_14_27=>d_arr_mul_14_27, d_arr_mul_14_26=>d_arr_mul_14_26, 
      d_arr_mul_14_25=>d_arr_mul_14_25, d_arr_mul_14_24=>d_arr_mul_14_24, 
      d_arr_mul_14_23=>d_arr_mul_14_23, d_arr_mul_14_22=>d_arr_mul_14_22, 
      d_arr_mul_14_21=>d_arr_mul_14_21, d_arr_mul_14_20=>d_arr_mul_14_20, 
      d_arr_mul_14_19=>d_arr_mul_14_19, d_arr_mul_14_18=>d_arr_mul_14_18, 
      d_arr_mul_14_17=>d_arr_mul_14_17, d_arr_mul_14_16=>d_arr_mul_14_16, 
      d_arr_mul_14_15=>d_arr_mul_14_15, d_arr_mul_14_14=>d_arr_mul_14_14, 
      d_arr_mul_14_13=>d_arr_mul_14_13, d_arr_mul_14_12=>d_arr_mul_14_12, 
      d_arr_mul_14_11=>d_arr_mul_14_11, d_arr_mul_14_10=>d_arr_mul_14_10, 
      d_arr_mul_14_9=>d_arr_mul_14_9, d_arr_mul_14_8=>d_arr_mul_14_8, 
      d_arr_mul_14_7=>d_arr_mul_14_7, d_arr_mul_14_6=>d_arr_mul_14_6, 
      d_arr_mul_14_5=>d_arr_mul_14_5, d_arr_mul_14_4=>d_arr_mul_14_4, 
      d_arr_mul_14_3=>d_arr_mul_14_3, d_arr_mul_14_2=>d_arr_mul_14_2, 
      d_arr_mul_14_1=>d_arr_mul_14_1, d_arr_mul_14_0=>d_arr_mul_14_0, 
      d_arr_mul_15_31=>d_arr_mul_15_31, d_arr_mul_15_30=>d_arr_mul_15_30, 
      d_arr_mul_15_29=>d_arr_mul_15_29, d_arr_mul_15_28=>d_arr_mul_15_28, 
      d_arr_mul_15_27=>d_arr_mul_15_27, d_arr_mul_15_26=>d_arr_mul_15_26, 
      d_arr_mul_15_25=>d_arr_mul_15_25, d_arr_mul_15_24=>d_arr_mul_15_24, 
      d_arr_mul_15_23=>d_arr_mul_15_23, d_arr_mul_15_22=>d_arr_mul_15_22, 
      d_arr_mul_15_21=>d_arr_mul_15_21, d_arr_mul_15_20=>d_arr_mul_15_20, 
      d_arr_mul_15_19=>d_arr_mul_15_19, d_arr_mul_15_18=>d_arr_mul_15_18, 
      d_arr_mul_15_17=>d_arr_mul_15_17, d_arr_mul_15_16=>d_arr_mul_15_16, 
      d_arr_mul_15_15=>d_arr_mul_15_15, d_arr_mul_15_14=>d_arr_mul_15_14, 
      d_arr_mul_15_13=>d_arr_mul_15_13, d_arr_mul_15_12=>d_arr_mul_15_12, 
      d_arr_mul_15_11=>d_arr_mul_15_11, d_arr_mul_15_10=>d_arr_mul_15_10, 
      d_arr_mul_15_9=>d_arr_mul_15_9, d_arr_mul_15_8=>d_arr_mul_15_8, 
      d_arr_mul_15_7=>d_arr_mul_15_7, d_arr_mul_15_6=>d_arr_mul_15_6, 
      d_arr_mul_15_5=>d_arr_mul_15_5, d_arr_mul_15_4=>d_arr_mul_15_4, 
      d_arr_mul_15_3=>d_arr_mul_15_3, d_arr_mul_15_2=>d_arr_mul_15_2, 
      d_arr_mul_15_1=>d_arr_mul_15_1, d_arr_mul_15_0=>d_arr_mul_15_0, 
      d_arr_mul_16_31=>d_arr_mul_16_31, d_arr_mul_16_30=>d_arr_mul_16_30, 
      d_arr_mul_16_29=>d_arr_mul_16_29, d_arr_mul_16_28=>d_arr_mul_16_28, 
      d_arr_mul_16_27=>d_arr_mul_16_27, d_arr_mul_16_26=>d_arr_mul_16_26, 
      d_arr_mul_16_25=>d_arr_mul_16_25, d_arr_mul_16_24=>d_arr_mul_16_24, 
      d_arr_mul_16_23=>d_arr_mul_16_23, d_arr_mul_16_22=>d_arr_mul_16_22, 
      d_arr_mul_16_21=>d_arr_mul_16_21, d_arr_mul_16_20=>d_arr_mul_16_20, 
      d_arr_mul_16_19=>d_arr_mul_16_19, d_arr_mul_16_18=>d_arr_mul_16_18, 
      d_arr_mul_16_17=>d_arr_mul_16_17, d_arr_mul_16_16=>d_arr_mul_16_16, 
      d_arr_mul_16_15=>d_arr_mul_16_15, d_arr_mul_16_14=>d_arr_mul_16_14, 
      d_arr_mul_16_13=>d_arr_mul_16_13, d_arr_mul_16_12=>d_arr_mul_16_12, 
      d_arr_mul_16_11=>d_arr_mul_16_11, d_arr_mul_16_10=>d_arr_mul_16_10, 
      d_arr_mul_16_9=>d_arr_mul_16_9, d_arr_mul_16_8=>d_arr_mul_16_8, 
      d_arr_mul_16_7=>d_arr_mul_16_7, d_arr_mul_16_6=>d_arr_mul_16_6, 
      d_arr_mul_16_5=>d_arr_mul_16_5, d_arr_mul_16_4=>d_arr_mul_16_4, 
      d_arr_mul_16_3=>d_arr_mul_16_3, d_arr_mul_16_2=>d_arr_mul_16_2, 
      d_arr_mul_16_1=>d_arr_mul_16_1, d_arr_mul_16_0=>d_arr_mul_16_0, 
      d_arr_mul_17_31=>d_arr_mul_17_31, d_arr_mul_17_30=>d_arr_mul_17_30, 
      d_arr_mul_17_29=>d_arr_mul_17_29, d_arr_mul_17_28=>d_arr_mul_17_28, 
      d_arr_mul_17_27=>d_arr_mul_17_27, d_arr_mul_17_26=>d_arr_mul_17_26, 
      d_arr_mul_17_25=>d_arr_mul_17_25, d_arr_mul_17_24=>d_arr_mul_17_24, 
      d_arr_mul_17_23=>d_arr_mul_17_23, d_arr_mul_17_22=>d_arr_mul_17_22, 
      d_arr_mul_17_21=>d_arr_mul_17_21, d_arr_mul_17_20=>d_arr_mul_17_20, 
      d_arr_mul_17_19=>d_arr_mul_17_19, d_arr_mul_17_18=>d_arr_mul_17_18, 
      d_arr_mul_17_17=>d_arr_mul_17_17, d_arr_mul_17_16=>d_arr_mul_17_16, 
      d_arr_mul_17_15=>d_arr_mul_17_15, d_arr_mul_17_14=>d_arr_mul_17_14, 
      d_arr_mul_17_13=>d_arr_mul_17_13, d_arr_mul_17_12=>d_arr_mul_17_12, 
      d_arr_mul_17_11=>d_arr_mul_17_11, d_arr_mul_17_10=>d_arr_mul_17_10, 
      d_arr_mul_17_9=>d_arr_mul_17_9, d_arr_mul_17_8=>d_arr_mul_17_8, 
      d_arr_mul_17_7=>d_arr_mul_17_7, d_arr_mul_17_6=>d_arr_mul_17_6, 
      d_arr_mul_17_5=>d_arr_mul_17_5, d_arr_mul_17_4=>d_arr_mul_17_4, 
      d_arr_mul_17_3=>d_arr_mul_17_3, d_arr_mul_17_2=>d_arr_mul_17_2, 
      d_arr_mul_17_1=>d_arr_mul_17_1, d_arr_mul_17_0=>d_arr_mul_17_0, 
      d_arr_mul_18_31=>d_arr_mul_18_31, d_arr_mul_18_30=>d_arr_mul_18_30, 
      d_arr_mul_18_29=>d_arr_mul_18_29, d_arr_mul_18_28=>d_arr_mul_18_28, 
      d_arr_mul_18_27=>d_arr_mul_18_27, d_arr_mul_18_26=>d_arr_mul_18_26, 
      d_arr_mul_18_25=>d_arr_mul_18_25, d_arr_mul_18_24=>d_arr_mul_18_24, 
      d_arr_mul_18_23=>d_arr_mul_18_23, d_arr_mul_18_22=>d_arr_mul_18_22, 
      d_arr_mul_18_21=>d_arr_mul_18_21, d_arr_mul_18_20=>d_arr_mul_18_20, 
      d_arr_mul_18_19=>d_arr_mul_18_19, d_arr_mul_18_18=>d_arr_mul_18_18, 
      d_arr_mul_18_17=>d_arr_mul_18_17, d_arr_mul_18_16=>d_arr_mul_18_16, 
      d_arr_mul_18_15=>d_arr_mul_18_15, d_arr_mul_18_14=>d_arr_mul_18_14, 
      d_arr_mul_18_13=>d_arr_mul_18_13, d_arr_mul_18_12=>d_arr_mul_18_12, 
      d_arr_mul_18_11=>d_arr_mul_18_11, d_arr_mul_18_10=>d_arr_mul_18_10, 
      d_arr_mul_18_9=>d_arr_mul_18_9, d_arr_mul_18_8=>d_arr_mul_18_8, 
      d_arr_mul_18_7=>d_arr_mul_18_7, d_arr_mul_18_6=>d_arr_mul_18_6, 
      d_arr_mul_18_5=>d_arr_mul_18_5, d_arr_mul_18_4=>d_arr_mul_18_4, 
      d_arr_mul_18_3=>d_arr_mul_18_3, d_arr_mul_18_2=>d_arr_mul_18_2, 
      d_arr_mul_18_1=>d_arr_mul_18_1, d_arr_mul_18_0=>d_arr_mul_18_0, 
      d_arr_mul_19_31=>d_arr_mul_19_31, d_arr_mul_19_30=>d_arr_mul_19_30, 
      d_arr_mul_19_29=>d_arr_mul_19_29, d_arr_mul_19_28=>d_arr_mul_19_28, 
      d_arr_mul_19_27=>d_arr_mul_19_27, d_arr_mul_19_26=>d_arr_mul_19_26, 
      d_arr_mul_19_25=>d_arr_mul_19_25, d_arr_mul_19_24=>d_arr_mul_19_24, 
      d_arr_mul_19_23=>d_arr_mul_19_23, d_arr_mul_19_22=>d_arr_mul_19_22, 
      d_arr_mul_19_21=>d_arr_mul_19_21, d_arr_mul_19_20=>d_arr_mul_19_20, 
      d_arr_mul_19_19=>d_arr_mul_19_19, d_arr_mul_19_18=>d_arr_mul_19_18, 
      d_arr_mul_19_17=>d_arr_mul_19_17, d_arr_mul_19_16=>d_arr_mul_19_16, 
      d_arr_mul_19_15=>d_arr_mul_19_15, d_arr_mul_19_14=>d_arr_mul_19_14, 
      d_arr_mul_19_13=>d_arr_mul_19_13, d_arr_mul_19_12=>d_arr_mul_19_12, 
      d_arr_mul_19_11=>d_arr_mul_19_11, d_arr_mul_19_10=>d_arr_mul_19_10, 
      d_arr_mul_19_9=>d_arr_mul_19_9, d_arr_mul_19_8=>d_arr_mul_19_8, 
      d_arr_mul_19_7=>d_arr_mul_19_7, d_arr_mul_19_6=>d_arr_mul_19_6, 
      d_arr_mul_19_5=>d_arr_mul_19_5, d_arr_mul_19_4=>d_arr_mul_19_4, 
      d_arr_mul_19_3=>d_arr_mul_19_3, d_arr_mul_19_2=>d_arr_mul_19_2, 
      d_arr_mul_19_1=>d_arr_mul_19_1, d_arr_mul_19_0=>d_arr_mul_19_0, 
      d_arr_mul_20_31=>d_arr_mul_20_31, d_arr_mul_20_30=>d_arr_mul_20_30, 
      d_arr_mul_20_29=>d_arr_mul_20_29, d_arr_mul_20_28=>d_arr_mul_20_28, 
      d_arr_mul_20_27=>d_arr_mul_20_27, d_arr_mul_20_26=>d_arr_mul_20_26, 
      d_arr_mul_20_25=>d_arr_mul_20_25, d_arr_mul_20_24=>d_arr_mul_20_24, 
      d_arr_mul_20_23=>d_arr_mul_20_23, d_arr_mul_20_22=>d_arr_mul_20_22, 
      d_arr_mul_20_21=>d_arr_mul_20_21, d_arr_mul_20_20=>d_arr_mul_20_20, 
      d_arr_mul_20_19=>d_arr_mul_20_19, d_arr_mul_20_18=>d_arr_mul_20_18, 
      d_arr_mul_20_17=>d_arr_mul_20_17, d_arr_mul_20_16=>d_arr_mul_20_16, 
      d_arr_mul_20_15=>d_arr_mul_20_15, d_arr_mul_20_14=>d_arr_mul_20_14, 
      d_arr_mul_20_13=>d_arr_mul_20_13, d_arr_mul_20_12=>d_arr_mul_20_12, 
      d_arr_mul_20_11=>d_arr_mul_20_11, d_arr_mul_20_10=>d_arr_mul_20_10, 
      d_arr_mul_20_9=>d_arr_mul_20_9, d_arr_mul_20_8=>d_arr_mul_20_8, 
      d_arr_mul_20_7=>d_arr_mul_20_7, d_arr_mul_20_6=>d_arr_mul_20_6, 
      d_arr_mul_20_5=>d_arr_mul_20_5, d_arr_mul_20_4=>d_arr_mul_20_4, 
      d_arr_mul_20_3=>d_arr_mul_20_3, d_arr_mul_20_2=>d_arr_mul_20_2, 
      d_arr_mul_20_1=>d_arr_mul_20_1, d_arr_mul_20_0=>d_arr_mul_20_0, 
      d_arr_mul_21_31=>d_arr_mul_21_31, d_arr_mul_21_30=>d_arr_mul_21_30, 
      d_arr_mul_21_29=>d_arr_mul_21_29, d_arr_mul_21_28=>d_arr_mul_21_28, 
      d_arr_mul_21_27=>d_arr_mul_21_27, d_arr_mul_21_26=>d_arr_mul_21_26, 
      d_arr_mul_21_25=>d_arr_mul_21_25, d_arr_mul_21_24=>d_arr_mul_21_24, 
      d_arr_mul_21_23=>d_arr_mul_21_23, d_arr_mul_21_22=>d_arr_mul_21_22, 
      d_arr_mul_21_21=>d_arr_mul_21_21, d_arr_mul_21_20=>d_arr_mul_21_20, 
      d_arr_mul_21_19=>d_arr_mul_21_19, d_arr_mul_21_18=>d_arr_mul_21_18, 
      d_arr_mul_21_17=>d_arr_mul_21_17, d_arr_mul_21_16=>d_arr_mul_21_16, 
      d_arr_mul_21_15=>d_arr_mul_21_15, d_arr_mul_21_14=>d_arr_mul_21_14, 
      d_arr_mul_21_13=>d_arr_mul_21_13, d_arr_mul_21_12=>d_arr_mul_21_12, 
      d_arr_mul_21_11=>d_arr_mul_21_11, d_arr_mul_21_10=>d_arr_mul_21_10, 
      d_arr_mul_21_9=>d_arr_mul_21_9, d_arr_mul_21_8=>d_arr_mul_21_8, 
      d_arr_mul_21_7=>d_arr_mul_21_7, d_arr_mul_21_6=>d_arr_mul_21_6, 
      d_arr_mul_21_5=>d_arr_mul_21_5, d_arr_mul_21_4=>d_arr_mul_21_4, 
      d_arr_mul_21_3=>d_arr_mul_21_3, d_arr_mul_21_2=>d_arr_mul_21_2, 
      d_arr_mul_21_1=>d_arr_mul_21_1, d_arr_mul_21_0=>d_arr_mul_21_0, 
      d_arr_mul_22_31=>d_arr_mul_22_31, d_arr_mul_22_30=>d_arr_mul_22_30, 
      d_arr_mul_22_29=>d_arr_mul_22_29, d_arr_mul_22_28=>d_arr_mul_22_28, 
      d_arr_mul_22_27=>d_arr_mul_22_27, d_arr_mul_22_26=>d_arr_mul_22_26, 
      d_arr_mul_22_25=>d_arr_mul_22_25, d_arr_mul_22_24=>d_arr_mul_22_24, 
      d_arr_mul_22_23=>d_arr_mul_22_23, d_arr_mul_22_22=>d_arr_mul_22_22, 
      d_arr_mul_22_21=>d_arr_mul_22_21, d_arr_mul_22_20=>d_arr_mul_22_20, 
      d_arr_mul_22_19=>d_arr_mul_22_19, d_arr_mul_22_18=>d_arr_mul_22_18, 
      d_arr_mul_22_17=>d_arr_mul_22_17, d_arr_mul_22_16=>d_arr_mul_22_16, 
      d_arr_mul_22_15=>d_arr_mul_22_15, d_arr_mul_22_14=>d_arr_mul_22_14, 
      d_arr_mul_22_13=>d_arr_mul_22_13, d_arr_mul_22_12=>d_arr_mul_22_12, 
      d_arr_mul_22_11=>d_arr_mul_22_11, d_arr_mul_22_10=>d_arr_mul_22_10, 
      d_arr_mul_22_9=>d_arr_mul_22_9, d_arr_mul_22_8=>d_arr_mul_22_8, 
      d_arr_mul_22_7=>d_arr_mul_22_7, d_arr_mul_22_6=>d_arr_mul_22_6, 
      d_arr_mul_22_5=>d_arr_mul_22_5, d_arr_mul_22_4=>d_arr_mul_22_4, 
      d_arr_mul_22_3=>d_arr_mul_22_3, d_arr_mul_22_2=>d_arr_mul_22_2, 
      d_arr_mul_22_1=>d_arr_mul_22_1, d_arr_mul_22_0=>d_arr_mul_22_0, 
      d_arr_mul_23_31=>d_arr_mul_23_31, d_arr_mul_23_30=>d_arr_mul_23_30, 
      d_arr_mul_23_29=>d_arr_mul_23_29, d_arr_mul_23_28=>d_arr_mul_23_28, 
      d_arr_mul_23_27=>d_arr_mul_23_27, d_arr_mul_23_26=>d_arr_mul_23_26, 
      d_arr_mul_23_25=>d_arr_mul_23_25, d_arr_mul_23_24=>d_arr_mul_23_24, 
      d_arr_mul_23_23=>d_arr_mul_23_23, d_arr_mul_23_22=>d_arr_mul_23_22, 
      d_arr_mul_23_21=>d_arr_mul_23_21, d_arr_mul_23_20=>d_arr_mul_23_20, 
      d_arr_mul_23_19=>d_arr_mul_23_19, d_arr_mul_23_18=>d_arr_mul_23_18, 
      d_arr_mul_23_17=>d_arr_mul_23_17, d_arr_mul_23_16=>d_arr_mul_23_16, 
      d_arr_mul_23_15=>d_arr_mul_23_15, d_arr_mul_23_14=>d_arr_mul_23_14, 
      d_arr_mul_23_13=>d_arr_mul_23_13, d_arr_mul_23_12=>d_arr_mul_23_12, 
      d_arr_mul_23_11=>d_arr_mul_23_11, d_arr_mul_23_10=>d_arr_mul_23_10, 
      d_arr_mul_23_9=>d_arr_mul_23_9, d_arr_mul_23_8=>d_arr_mul_23_8, 
      d_arr_mul_23_7=>d_arr_mul_23_7, d_arr_mul_23_6=>d_arr_mul_23_6, 
      d_arr_mul_23_5=>d_arr_mul_23_5, d_arr_mul_23_4=>d_arr_mul_23_4, 
      d_arr_mul_23_3=>d_arr_mul_23_3, d_arr_mul_23_2=>d_arr_mul_23_2, 
      d_arr_mul_23_1=>d_arr_mul_23_1, d_arr_mul_23_0=>d_arr_mul_23_0, 
      d_arr_mul_24_31=>d_arr_mul_24_31, d_arr_mul_24_30=>d_arr_mul_24_30, 
      d_arr_mul_24_29=>d_arr_mul_24_29, d_arr_mul_24_28=>d_arr_mul_24_28, 
      d_arr_mul_24_27=>d_arr_mul_24_27, d_arr_mul_24_26=>d_arr_mul_24_26, 
      d_arr_mul_24_25=>d_arr_mul_24_25, d_arr_mul_24_24=>d_arr_mul_24_24, 
      d_arr_mul_24_23=>d_arr_mul_24_23, d_arr_mul_24_22=>d_arr_mul_24_22, 
      d_arr_mul_24_21=>d_arr_mul_24_21, d_arr_mul_24_20=>d_arr_mul_24_20, 
      d_arr_mul_24_19=>d_arr_mul_24_19, d_arr_mul_24_18=>d_arr_mul_24_18, 
      d_arr_mul_24_17=>d_arr_mul_24_17, d_arr_mul_24_16=>d_arr_mul_24_16, 
      d_arr_mul_24_15=>d_arr_mul_24_15, d_arr_mul_24_14=>d_arr_mul_24_14, 
      d_arr_mul_24_13=>d_arr_mul_24_13, d_arr_mul_24_12=>d_arr_mul_24_12, 
      d_arr_mul_24_11=>d_arr_mul_24_11, d_arr_mul_24_10=>d_arr_mul_24_10, 
      d_arr_mul_24_9=>d_arr_mul_24_9, d_arr_mul_24_8=>d_arr_mul_24_8, 
      d_arr_mul_24_7=>d_arr_mul_24_7, d_arr_mul_24_6=>d_arr_mul_24_6, 
      d_arr_mul_24_5=>d_arr_mul_24_5, d_arr_mul_24_4=>d_arr_mul_24_4, 
      d_arr_mul_24_3=>d_arr_mul_24_3, d_arr_mul_24_2=>d_arr_mul_24_2, 
      d_arr_mul_24_1=>d_arr_mul_24_1, d_arr_mul_24_0=>d_arr_mul_24_0, 
      d_arr_add_0_31=>d_arr_add_0_31, d_arr_add_0_30=>d_arr_add_0_30, 
      d_arr_add_0_29=>d_arr_add_0_29, d_arr_add_0_28=>d_arr_add_0_28, 
      d_arr_add_0_27=>d_arr_add_0_27, d_arr_add_0_26=>d_arr_add_0_26, 
      d_arr_add_0_25=>d_arr_add_0_25, d_arr_add_0_24=>d_arr_add_0_24, 
      d_arr_add_0_23=>d_arr_add_0_23, d_arr_add_0_22=>d_arr_add_0_22, 
      d_arr_add_0_21=>d_arr_add_0_21, d_arr_add_0_20=>d_arr_add_0_20, 
      d_arr_add_0_19=>d_arr_add_0_19, d_arr_add_0_18=>d_arr_add_0_18, 
      d_arr_add_0_17=>d_arr_add_0_17, d_arr_add_0_16=>d_arr_add_0_16, 
      d_arr_add_0_15=>d_arr_add_0_15, d_arr_add_0_14=>d_arr_add_0_14, 
      d_arr_add_0_13=>d_arr_add_0_13, d_arr_add_0_12=>d_arr_add_0_12, 
      d_arr_add_0_11=>d_arr_add_0_11, d_arr_add_0_10=>d_arr_add_0_10, 
      d_arr_add_0_9=>d_arr_add_0_9, d_arr_add_0_8=>d_arr_add_0_8, 
      d_arr_add_0_7=>d_arr_add_0_7, d_arr_add_0_6=>d_arr_add_0_6, 
      d_arr_add_0_5=>d_arr_add_0_5, d_arr_add_0_4=>d_arr_add_0_4, 
      d_arr_add_0_3=>d_arr_add_0_3, d_arr_add_0_2=>d_arr_add_0_2, 
      d_arr_add_0_1=>d_arr_add_0_1, d_arr_add_0_0=>d_arr_add_0_0, 
      d_arr_add_1_31=>d_arr_add_1_31, d_arr_add_1_30=>d_arr_add_1_30, 
      d_arr_add_1_29=>d_arr_add_1_29, d_arr_add_1_28=>d_arr_add_1_28, 
      d_arr_add_1_27=>d_arr_add_1_27, d_arr_add_1_26=>d_arr_add_1_26, 
      d_arr_add_1_25=>d_arr_add_1_25, d_arr_add_1_24=>d_arr_add_1_24, 
      d_arr_add_1_23=>d_arr_add_1_23, d_arr_add_1_22=>d_arr_add_1_22, 
      d_arr_add_1_21=>d_arr_add_1_21, d_arr_add_1_20=>d_arr_add_1_20, 
      d_arr_add_1_19=>d_arr_add_1_19, d_arr_add_1_18=>d_arr_add_1_18, 
      d_arr_add_1_17=>d_arr_add_1_17, d_arr_add_1_16=>d_arr_add_1_16, 
      d_arr_add_1_15=>d_arr_add_1_15, d_arr_add_1_14=>d_arr_add_1_14, 
      d_arr_add_1_13=>d_arr_add_1_13, d_arr_add_1_12=>d_arr_add_1_12, 
      d_arr_add_1_11=>d_arr_add_1_11, d_arr_add_1_10=>d_arr_add_1_10, 
      d_arr_add_1_9=>d_arr_add_1_9, d_arr_add_1_8=>d_arr_add_1_8, 
      d_arr_add_1_7=>d_arr_add_1_7, d_arr_add_1_6=>d_arr_add_1_6, 
      d_arr_add_1_5=>d_arr_add_1_5, d_arr_add_1_4=>d_arr_add_1_4, 
      d_arr_add_1_3=>d_arr_add_1_3, d_arr_add_1_2=>d_arr_add_1_2, 
      d_arr_add_1_1=>d_arr_add_1_1, d_arr_add_1_0=>d_arr_add_1_0, 
      d_arr_add_2_31=>d_arr_add_2_31, d_arr_add_2_30=>d_arr_add_2_30, 
      d_arr_add_2_29=>d_arr_add_2_29, d_arr_add_2_28=>d_arr_add_2_28, 
      d_arr_add_2_27=>d_arr_add_2_27, d_arr_add_2_26=>d_arr_add_2_26, 
      d_arr_add_2_25=>d_arr_add_2_25, d_arr_add_2_24=>d_arr_add_2_24, 
      d_arr_add_2_23=>d_arr_add_2_23, d_arr_add_2_22=>d_arr_add_2_22, 
      d_arr_add_2_21=>d_arr_add_2_21, d_arr_add_2_20=>d_arr_add_2_20, 
      d_arr_add_2_19=>d_arr_add_2_19, d_arr_add_2_18=>d_arr_add_2_18, 
      d_arr_add_2_17=>d_arr_add_2_17, d_arr_add_2_16=>d_arr_add_2_16, 
      d_arr_add_2_15=>d_arr_add_2_15, d_arr_add_2_14=>d_arr_add_2_14, 
      d_arr_add_2_13=>d_arr_add_2_13, d_arr_add_2_12=>d_arr_add_2_12, 
      d_arr_add_2_11=>d_arr_add_2_11, d_arr_add_2_10=>d_arr_add_2_10, 
      d_arr_add_2_9=>d_arr_add_2_9, d_arr_add_2_8=>d_arr_add_2_8, 
      d_arr_add_2_7=>d_arr_add_2_7, d_arr_add_2_6=>d_arr_add_2_6, 
      d_arr_add_2_5=>d_arr_add_2_5, d_arr_add_2_4=>d_arr_add_2_4, 
      d_arr_add_2_3=>d_arr_add_2_3, d_arr_add_2_2=>d_arr_add_2_2, 
      d_arr_add_2_1=>d_arr_add_2_1, d_arr_add_2_0=>d_arr_add_2_0, 
      d_arr_add_3_31=>d_arr_add_3_31, d_arr_add_3_30=>d_arr_add_3_30, 
      d_arr_add_3_29=>d_arr_add_3_29, d_arr_add_3_28=>d_arr_add_3_28, 
      d_arr_add_3_27=>d_arr_add_3_27, d_arr_add_3_26=>d_arr_add_3_26, 
      d_arr_add_3_25=>d_arr_add_3_25, d_arr_add_3_24=>d_arr_add_3_24, 
      d_arr_add_3_23=>d_arr_add_3_23, d_arr_add_3_22=>d_arr_add_3_22, 
      d_arr_add_3_21=>d_arr_add_3_21, d_arr_add_3_20=>d_arr_add_3_20, 
      d_arr_add_3_19=>d_arr_add_3_19, d_arr_add_3_18=>d_arr_add_3_18, 
      d_arr_add_3_17=>d_arr_add_3_17, d_arr_add_3_16=>d_arr_add_3_16, 
      d_arr_add_3_15=>d_arr_add_3_15, d_arr_add_3_14=>d_arr_add_3_14, 
      d_arr_add_3_13=>d_arr_add_3_13, d_arr_add_3_12=>d_arr_add_3_12, 
      d_arr_add_3_11=>d_arr_add_3_11, d_arr_add_3_10=>d_arr_add_3_10, 
      d_arr_add_3_9=>d_arr_add_3_9, d_arr_add_3_8=>d_arr_add_3_8, 
      d_arr_add_3_7=>d_arr_add_3_7, d_arr_add_3_6=>d_arr_add_3_6, 
      d_arr_add_3_5=>d_arr_add_3_5, d_arr_add_3_4=>d_arr_add_3_4, 
      d_arr_add_3_3=>d_arr_add_3_3, d_arr_add_3_2=>d_arr_add_3_2, 
      d_arr_add_3_1=>d_arr_add_3_1, d_arr_add_3_0=>d_arr_add_3_0, 
      d_arr_add_4_31=>q_arr_8_31, d_arr_add_4_30=>q_arr_8_30, d_arr_add_4_29
      =>q_arr_8_29, d_arr_add_4_28=>q_arr_8_28, d_arr_add_4_27=>q_arr_8_27, 
      d_arr_add_4_26=>q_arr_8_26, d_arr_add_4_25=>q_arr_8_25, d_arr_add_4_24
      =>q_arr_8_24, d_arr_add_4_23=>q_arr_8_23, d_arr_add_4_22=>q_arr_8_22, 
      d_arr_add_4_21=>q_arr_8_21, d_arr_add_4_20=>q_arr_8_20, d_arr_add_4_19
      =>q_arr_8_19, d_arr_add_4_18=>q_arr_8_18, d_arr_add_4_17=>q_arr_8_17, 
      d_arr_add_4_16=>q_arr_8_16, d_arr_add_4_15=>q_arr_8_15, d_arr_add_4_14
      =>q_arr_8_14, d_arr_add_4_13=>q_arr_8_13, d_arr_add_4_12=>q_arr_8_12, 
      d_arr_add_4_11=>q_arr_8_11, d_arr_add_4_10=>q_arr_8_10, d_arr_add_4_9
      =>q_arr_8_9, d_arr_add_4_8=>q_arr_8_8, d_arr_add_4_7=>q_arr_8_7, 
      d_arr_add_4_6=>q_arr_8_6, d_arr_add_4_5=>q_arr_8_5, d_arr_add_4_4=>
      q_arr_8_4, d_arr_add_4_3=>q_arr_8_3, d_arr_add_4_2=>q_arr_8_2, 
      d_arr_add_4_1=>q_arr_8_1, d_arr_add_4_0=>q_arr_8_0, d_arr_add_5_31=>
      GND0, d_arr_add_5_30=>GND0, d_arr_add_5_29=>GND0, d_arr_add_5_28=>GND0, 
      d_arr_add_5_27=>GND0, d_arr_add_5_26=>GND0, d_arr_add_5_25=>GND0, 
      d_arr_add_5_24=>GND0, d_arr_add_5_23=>GND0, d_arr_add_5_22=>GND0, 
      d_arr_add_5_21=>GND0, d_arr_add_5_20=>GND0, d_arr_add_5_19=>GND0, 
      d_arr_add_5_18=>GND0, d_arr_add_5_17=>GND0, d_arr_add_5_16=>GND0, 
      d_arr_add_5_15=>GND0, d_arr_add_5_14=>GND0, d_arr_add_5_13=>GND0, 
      d_arr_add_5_12=>GND0, d_arr_add_5_11=>GND0, d_arr_add_5_10=>GND0, 
      d_arr_add_5_9=>GND0, d_arr_add_5_8=>GND0, d_arr_add_5_7=>GND0, 
      d_arr_add_5_6=>GND0, d_arr_add_5_5=>GND0, d_arr_add_5_4=>GND0, 
      d_arr_add_5_3=>GND0, d_arr_add_5_2=>GND0, d_arr_add_5_1=>GND0, 
      d_arr_add_5_0=>GND0, d_arr_add_6_31=>GND0, d_arr_add_6_30=>GND0, 
      d_arr_add_6_29=>GND0, d_arr_add_6_28=>GND0, d_arr_add_6_27=>GND0, 
      d_arr_add_6_26=>GND0, d_arr_add_6_25=>GND0, d_arr_add_6_24=>GND0, 
      d_arr_add_6_23=>GND0, d_arr_add_6_22=>GND0, d_arr_add_6_21=>GND0, 
      d_arr_add_6_20=>GND0, d_arr_add_6_19=>GND0, d_arr_add_6_18=>GND0, 
      d_arr_add_6_17=>GND0, d_arr_add_6_16=>GND0, d_arr_add_6_15=>GND0, 
      d_arr_add_6_14=>GND0, d_arr_add_6_13=>GND0, d_arr_add_6_12=>GND0, 
      d_arr_add_6_11=>GND0, d_arr_add_6_10=>GND0, d_arr_add_6_9=>GND0, 
      d_arr_add_6_8=>GND0, d_arr_add_6_7=>GND0, d_arr_add_6_6=>GND0, 
      d_arr_add_6_5=>GND0, d_arr_add_6_4=>GND0, d_arr_add_6_3=>GND0, 
      d_arr_add_6_2=>GND0, d_arr_add_6_1=>GND0, d_arr_add_6_0=>GND0, 
      d_arr_add_7_31=>GND0, d_arr_add_7_30=>GND0, d_arr_add_7_29=>GND0, 
      d_arr_add_7_28=>GND0, d_arr_add_7_27=>GND0, d_arr_add_7_26=>GND0, 
      d_arr_add_7_25=>GND0, d_arr_add_7_24=>GND0, d_arr_add_7_23=>GND0, 
      d_arr_add_7_22=>GND0, d_arr_add_7_21=>GND0, d_arr_add_7_20=>GND0, 
      d_arr_add_7_19=>GND0, d_arr_add_7_18=>GND0, d_arr_add_7_17=>GND0, 
      d_arr_add_7_16=>GND0, d_arr_add_7_15=>GND0, d_arr_add_7_14=>GND0, 
      d_arr_add_7_13=>GND0, d_arr_add_7_12=>GND0, d_arr_add_7_11=>GND0, 
      d_arr_add_7_10=>GND0, d_arr_add_7_9=>GND0, d_arr_add_7_8=>GND0, 
      d_arr_add_7_7=>GND0, d_arr_add_7_6=>GND0, d_arr_add_7_5=>GND0, 
      d_arr_add_7_4=>GND0, d_arr_add_7_3=>GND0, d_arr_add_7_2=>GND0, 
      d_arr_add_7_1=>GND0, d_arr_add_7_0=>GND0, d_arr_add_8_31=>GND0, 
      d_arr_add_8_30=>GND0, d_arr_add_8_29=>GND0, d_arr_add_8_28=>GND0, 
      d_arr_add_8_27=>GND0, d_arr_add_8_26=>GND0, d_arr_add_8_25=>GND0, 
      d_arr_add_8_24=>GND0, d_arr_add_8_23=>GND0, d_arr_add_8_22=>GND0, 
      d_arr_add_8_21=>GND0, d_arr_add_8_20=>GND0, d_arr_add_8_19=>GND0, 
      d_arr_add_8_18=>GND0, d_arr_add_8_17=>GND0, d_arr_add_8_16=>GND0, 
      d_arr_add_8_15=>GND0, d_arr_add_8_14=>GND0, d_arr_add_8_13=>GND0, 
      d_arr_add_8_12=>GND0, d_arr_add_8_11=>GND0, d_arr_add_8_10=>GND0, 
      d_arr_add_8_9=>GND0, d_arr_add_8_8=>GND0, d_arr_add_8_7=>GND0, 
      d_arr_add_8_6=>GND0, d_arr_add_8_5=>GND0, d_arr_add_8_4=>GND0, 
      d_arr_add_8_3=>GND0, d_arr_add_8_2=>GND0, d_arr_add_8_1=>GND0, 
      d_arr_add_8_0=>GND0, d_arr_add_9_31=>d_arr_add_9_31, d_arr_add_9_30=>
      d_arr_add_9_30, d_arr_add_9_29=>d_arr_add_9_29, d_arr_add_9_28=>
      d_arr_add_9_28, d_arr_add_9_27=>d_arr_add_9_27, d_arr_add_9_26=>
      d_arr_add_9_26, d_arr_add_9_25=>d_arr_add_9_25, d_arr_add_9_24=>
      d_arr_add_9_24, d_arr_add_9_23=>d_arr_add_9_23, d_arr_add_9_22=>
      d_arr_add_9_22, d_arr_add_9_21=>d_arr_add_9_21, d_arr_add_9_20=>
      d_arr_add_9_20, d_arr_add_9_19=>d_arr_add_9_19, d_arr_add_9_18=>
      d_arr_add_9_18, d_arr_add_9_17=>d_arr_add_9_17, d_arr_add_9_16=>
      d_arr_add_9_16, d_arr_add_9_15=>d_arr_add_9_15, d_arr_add_9_14=>
      d_arr_add_9_14, d_arr_add_9_13=>d_arr_add_9_13, d_arr_add_9_12=>
      d_arr_add_9_12, d_arr_add_9_11=>d_arr_add_9_11, d_arr_add_9_10=>
      d_arr_add_9_10, d_arr_add_9_9=>d_arr_add_9_9, d_arr_add_9_8=>
      d_arr_add_9_8, d_arr_add_9_7=>d_arr_add_9_7, d_arr_add_9_6=>
      d_arr_add_9_6, d_arr_add_9_5=>d_arr_add_9_5, d_arr_add_9_4=>
      d_arr_add_9_4, d_arr_add_9_3=>d_arr_add_9_3, d_arr_add_9_2=>
      d_arr_add_9_2, d_arr_add_9_1=>d_arr_add_9_1, d_arr_add_9_0=>
      d_arr_add_9_0, d_arr_add_10_31=>d_arr_add_10_31, d_arr_add_10_30=>
      d_arr_add_10_30, d_arr_add_10_29=>d_arr_add_10_29, d_arr_add_10_28=>
      d_arr_add_10_28, d_arr_add_10_27=>d_arr_add_10_27, d_arr_add_10_26=>
      d_arr_add_10_26, d_arr_add_10_25=>d_arr_add_10_25, d_arr_add_10_24=>
      d_arr_add_10_24, d_arr_add_10_23=>d_arr_add_10_23, d_arr_add_10_22=>
      d_arr_add_10_22, d_arr_add_10_21=>d_arr_add_10_21, d_arr_add_10_20=>
      d_arr_add_10_20, d_arr_add_10_19=>d_arr_add_10_19, d_arr_add_10_18=>
      d_arr_add_10_18, d_arr_add_10_17=>d_arr_add_10_17, d_arr_add_10_16=>
      d_arr_add_10_16, d_arr_add_10_15=>d_arr_add_10_15, d_arr_add_10_14=>
      d_arr_add_10_14, d_arr_add_10_13=>d_arr_add_10_13, d_arr_add_10_12=>
      d_arr_add_10_12, d_arr_add_10_11=>d_arr_add_10_11, d_arr_add_10_10=>
      d_arr_add_10_10, d_arr_add_10_9=>d_arr_add_10_9, d_arr_add_10_8=>
      d_arr_add_10_8, d_arr_add_10_7=>d_arr_add_10_7, d_arr_add_10_6=>
      d_arr_add_10_6, d_arr_add_10_5=>d_arr_add_10_5, d_arr_add_10_4=>
      d_arr_add_10_4, d_arr_add_10_3=>d_arr_add_10_3, d_arr_add_10_2=>
      d_arr_add_10_2, d_arr_add_10_1=>d_arr_add_10_1, d_arr_add_10_0=>
      d_arr_add_10_0, d_arr_add_11_31=>d_arr_add_11_31, d_arr_add_11_30=>
      d_arr_add_11_30, d_arr_add_11_29=>d_arr_add_11_29, d_arr_add_11_28=>
      d_arr_add_11_28, d_arr_add_11_27=>d_arr_add_11_27, d_arr_add_11_26=>
      d_arr_add_11_26, d_arr_add_11_25=>d_arr_add_11_25, d_arr_add_11_24=>
      d_arr_add_11_24, d_arr_add_11_23=>d_arr_add_11_23, d_arr_add_11_22=>
      d_arr_add_11_22, d_arr_add_11_21=>d_arr_add_11_21, d_arr_add_11_20=>
      d_arr_add_11_20, d_arr_add_11_19=>d_arr_add_11_19, d_arr_add_11_18=>
      d_arr_add_11_18, d_arr_add_11_17=>d_arr_add_11_17, d_arr_add_11_16=>
      d_arr_add_11_16, d_arr_add_11_15=>d_arr_add_11_15, d_arr_add_11_14=>
      d_arr_add_11_14, d_arr_add_11_13=>d_arr_add_11_13, d_arr_add_11_12=>
      d_arr_add_11_12, d_arr_add_11_11=>d_arr_add_11_11, d_arr_add_11_10=>
      d_arr_add_11_10, d_arr_add_11_9=>d_arr_add_11_9, d_arr_add_11_8=>
      d_arr_add_11_8, d_arr_add_11_7=>d_arr_add_11_7, d_arr_add_11_6=>
      d_arr_add_11_6, d_arr_add_11_5=>d_arr_add_11_5, d_arr_add_11_4=>
      d_arr_add_11_4, d_arr_add_11_3=>d_arr_add_11_3, d_arr_add_11_2=>
      d_arr_add_11_2, d_arr_add_11_1=>d_arr_add_11_1, d_arr_add_11_0=>
      d_arr_add_11_0, d_arr_add_12_31=>d_arr_add_12_31, d_arr_add_12_30=>
      d_arr_add_12_30, d_arr_add_12_29=>d_arr_add_12_29, d_arr_add_12_28=>
      d_arr_add_12_28, d_arr_add_12_27=>d_arr_add_12_27, d_arr_add_12_26=>
      d_arr_add_12_26, d_arr_add_12_25=>d_arr_add_12_25, d_arr_add_12_24=>
      d_arr_add_12_24, d_arr_add_12_23=>d_arr_add_12_23, d_arr_add_12_22=>
      d_arr_add_12_22, d_arr_add_12_21=>d_arr_add_12_21, d_arr_add_12_20=>
      d_arr_add_12_20, d_arr_add_12_19=>d_arr_add_12_19, d_arr_add_12_18=>
      d_arr_add_12_18, d_arr_add_12_17=>d_arr_add_12_17, d_arr_add_12_16=>
      d_arr_add_12_16, d_arr_add_12_15=>d_arr_add_12_15, d_arr_add_12_14=>
      d_arr_add_12_14, d_arr_add_12_13=>d_arr_add_12_13, d_arr_add_12_12=>
      d_arr_add_12_12, d_arr_add_12_11=>d_arr_add_12_11, d_arr_add_12_10=>
      d_arr_add_12_10, d_arr_add_12_9=>d_arr_add_12_9, d_arr_add_12_8=>
      d_arr_add_12_8, d_arr_add_12_7=>d_arr_add_12_7, d_arr_add_12_6=>
      d_arr_add_12_6, d_arr_add_12_5=>d_arr_add_12_5, d_arr_add_12_4=>
      d_arr_add_12_4, d_arr_add_12_3=>d_arr_add_12_3, d_arr_add_12_2=>
      d_arr_add_12_2, d_arr_add_12_1=>d_arr_add_12_1, d_arr_add_12_0=>
      d_arr_add_12_0, d_arr_add_13_31=>q_arr_17_31, d_arr_add_13_30=>
      q_arr_17_30, d_arr_add_13_29=>q_arr_17_29, d_arr_add_13_28=>
      q_arr_17_28, d_arr_add_13_27=>q_arr_17_27, d_arr_add_13_26=>
      q_arr_17_26, d_arr_add_13_25=>q_arr_17_25, d_arr_add_13_24=>
      q_arr_17_24, d_arr_add_13_23=>q_arr_17_23, d_arr_add_13_22=>
      q_arr_17_22, d_arr_add_13_21=>q_arr_17_21, d_arr_add_13_20=>
      q_arr_17_20, d_arr_add_13_19=>q_arr_17_19, d_arr_add_13_18=>
      q_arr_17_18, d_arr_add_13_17=>q_arr_17_17, d_arr_add_13_16=>
      q_arr_17_16, d_arr_add_13_15=>q_arr_17_15, d_arr_add_13_14=>
      q_arr_17_14, d_arr_add_13_13=>q_arr_17_13, d_arr_add_13_12=>
      q_arr_17_12, d_arr_add_13_11=>q_arr_17_11, d_arr_add_13_10=>
      q_arr_17_10, d_arr_add_13_9=>q_arr_17_9, d_arr_add_13_8=>q_arr_17_8, 
      d_arr_add_13_7=>q_arr_17_7, d_arr_add_13_6=>q_arr_17_6, d_arr_add_13_5
      =>q_arr_17_5, d_arr_add_13_4=>q_arr_17_4, d_arr_add_13_3=>q_arr_17_3, 
      d_arr_add_13_2=>q_arr_17_2, d_arr_add_13_1=>q_arr_17_1, d_arr_add_13_0
      =>q_arr_17_0, d_arr_add_14_31=>GND0, d_arr_add_14_30=>GND0, 
      d_arr_add_14_29=>GND0, d_arr_add_14_28=>GND0, d_arr_add_14_27=>GND0, 
      d_arr_add_14_26=>GND0, d_arr_add_14_25=>GND0, d_arr_add_14_24=>GND0, 
      d_arr_add_14_23=>GND0, d_arr_add_14_22=>GND0, d_arr_add_14_21=>GND0, 
      d_arr_add_14_20=>GND0, d_arr_add_14_19=>GND0, d_arr_add_14_18=>GND0, 
      d_arr_add_14_17=>GND0, d_arr_add_14_16=>GND0, d_arr_add_14_15=>GND0, 
      d_arr_add_14_14=>GND0, d_arr_add_14_13=>GND0, d_arr_add_14_12=>GND0, 
      d_arr_add_14_11=>GND0, d_arr_add_14_10=>GND0, d_arr_add_14_9=>GND0, 
      d_arr_add_14_8=>GND0, d_arr_add_14_7=>GND0, d_arr_add_14_6=>GND0, 
      d_arr_add_14_5=>GND0, d_arr_add_14_4=>GND0, d_arr_add_14_3=>GND0, 
      d_arr_add_14_2=>GND0, d_arr_add_14_1=>GND0, d_arr_add_14_0=>GND0, 
      d_arr_add_15_31=>GND0, d_arr_add_15_30=>GND0, d_arr_add_15_29=>GND0, 
      d_arr_add_15_28=>GND0, d_arr_add_15_27=>GND0, d_arr_add_15_26=>GND0, 
      d_arr_add_15_25=>GND0, d_arr_add_15_24=>GND0, d_arr_add_15_23=>GND0, 
      d_arr_add_15_22=>GND0, d_arr_add_15_21=>GND0, d_arr_add_15_20=>GND0, 
      d_arr_add_15_19=>GND0, d_arr_add_15_18=>GND0, d_arr_add_15_17=>GND0, 
      d_arr_add_15_16=>GND0, d_arr_add_15_15=>GND0, d_arr_add_15_14=>GND0, 
      d_arr_add_15_13=>GND0, d_arr_add_15_12=>GND0, d_arr_add_15_11=>GND0, 
      d_arr_add_15_10=>GND0, d_arr_add_15_9=>GND0, d_arr_add_15_8=>GND0, 
      d_arr_add_15_7=>GND0, d_arr_add_15_6=>GND0, d_arr_add_15_5=>GND0, 
      d_arr_add_15_4=>GND0, d_arr_add_15_3=>GND0, d_arr_add_15_2=>GND0, 
      d_arr_add_15_1=>GND0, d_arr_add_15_0=>GND0, d_arr_add_16_31=>GND0, 
      d_arr_add_16_30=>GND0, d_arr_add_16_29=>GND0, d_arr_add_16_28=>GND0, 
      d_arr_add_16_27=>GND0, d_arr_add_16_26=>GND0, d_arr_add_16_25=>GND0, 
      d_arr_add_16_24=>GND0, d_arr_add_16_23=>GND0, d_arr_add_16_22=>GND0, 
      d_arr_add_16_21=>GND0, d_arr_add_16_20=>GND0, d_arr_add_16_19=>GND0, 
      d_arr_add_16_18=>GND0, d_arr_add_16_17=>GND0, d_arr_add_16_16=>GND0, 
      d_arr_add_16_15=>GND0, d_arr_add_16_14=>GND0, d_arr_add_16_13=>GND0, 
      d_arr_add_16_12=>GND0, d_arr_add_16_11=>GND0, d_arr_add_16_10=>GND0, 
      d_arr_add_16_9=>GND0, d_arr_add_16_8=>GND0, d_arr_add_16_7=>GND0, 
      d_arr_add_16_6=>GND0, d_arr_add_16_5=>GND0, d_arr_add_16_4=>GND0, 
      d_arr_add_16_3=>GND0, d_arr_add_16_2=>GND0, d_arr_add_16_1=>GND0, 
      d_arr_add_16_0=>GND0, d_arr_add_17_31=>GND0, d_arr_add_17_30=>GND0, 
      d_arr_add_17_29=>GND0, d_arr_add_17_28=>GND0, d_arr_add_17_27=>GND0, 
      d_arr_add_17_26=>GND0, d_arr_add_17_25=>GND0, d_arr_add_17_24=>GND0, 
      d_arr_add_17_23=>GND0, d_arr_add_17_22=>GND0, d_arr_add_17_21=>GND0, 
      d_arr_add_17_20=>GND0, d_arr_add_17_19=>GND0, d_arr_add_17_18=>GND0, 
      d_arr_add_17_17=>GND0, d_arr_add_17_16=>GND0, d_arr_add_17_15=>GND0, 
      d_arr_add_17_14=>GND0, d_arr_add_17_13=>GND0, d_arr_add_17_12=>GND0, 
      d_arr_add_17_11=>GND0, d_arr_add_17_10=>GND0, d_arr_add_17_9=>GND0, 
      d_arr_add_17_8=>GND0, d_arr_add_17_7=>GND0, d_arr_add_17_6=>GND0, 
      d_arr_add_17_5=>GND0, d_arr_add_17_4=>GND0, d_arr_add_17_3=>GND0, 
      d_arr_add_17_2=>GND0, d_arr_add_17_1=>GND0, d_arr_add_17_0=>GND0, 
      d_arr_add_18_31=>d_arr_add_18_31, d_arr_add_18_30=>d_arr_add_18_30, 
      d_arr_add_18_29=>d_arr_add_18_29, d_arr_add_18_28=>d_arr_add_18_28, 
      d_arr_add_18_27=>d_arr_add_18_27, d_arr_add_18_26=>d_arr_add_18_26, 
      d_arr_add_18_25=>d_arr_add_18_25, d_arr_add_18_24=>d_arr_add_18_24, 
      d_arr_add_18_23=>d_arr_add_18_23, d_arr_add_18_22=>d_arr_add_18_22, 
      d_arr_add_18_21=>d_arr_add_18_21, d_arr_add_18_20=>d_arr_add_18_20, 
      d_arr_add_18_19=>d_arr_add_18_19, d_arr_add_18_18=>d_arr_add_18_18, 
      d_arr_add_18_17=>d_arr_add_18_17, d_arr_add_18_16=>d_arr_add_18_16, 
      d_arr_add_18_15=>d_arr_add_18_15, d_arr_add_18_14=>d_arr_add_18_14, 
      d_arr_add_18_13=>d_arr_add_18_13, d_arr_add_18_12=>d_arr_add_18_12, 
      d_arr_add_18_11=>d_arr_add_18_11, d_arr_add_18_10=>d_arr_add_18_10, 
      d_arr_add_18_9=>d_arr_add_18_9, d_arr_add_18_8=>d_arr_add_18_8, 
      d_arr_add_18_7=>d_arr_add_18_7, d_arr_add_18_6=>d_arr_add_18_6, 
      d_arr_add_18_5=>d_arr_add_18_5, d_arr_add_18_4=>d_arr_add_18_4, 
      d_arr_add_18_3=>d_arr_add_18_3, d_arr_add_18_2=>d_arr_add_18_2, 
      d_arr_add_18_1=>d_arr_add_18_1, d_arr_add_18_0=>d_arr_add_18_0, 
      d_arr_add_19_31=>d_arr_add_19_31, d_arr_add_19_30=>d_arr_add_19_30, 
      d_arr_add_19_29=>d_arr_add_19_29, d_arr_add_19_28=>d_arr_add_19_28, 
      d_arr_add_19_27=>d_arr_add_19_27, d_arr_add_19_26=>d_arr_add_19_26, 
      d_arr_add_19_25=>d_arr_add_19_25, d_arr_add_19_24=>d_arr_add_19_24, 
      d_arr_add_19_23=>d_arr_add_19_23, d_arr_add_19_22=>d_arr_add_19_22, 
      d_arr_add_19_21=>d_arr_add_19_21, d_arr_add_19_20=>d_arr_add_19_20, 
      d_arr_add_19_19=>d_arr_add_19_19, d_arr_add_19_18=>d_arr_add_19_18, 
      d_arr_add_19_17=>d_arr_add_19_17, d_arr_add_19_16=>d_arr_add_19_16, 
      d_arr_add_19_15=>d_arr_add_19_15, d_arr_add_19_14=>d_arr_add_19_14, 
      d_arr_add_19_13=>d_arr_add_19_13, d_arr_add_19_12=>d_arr_add_19_12, 
      d_arr_add_19_11=>d_arr_add_19_11, d_arr_add_19_10=>d_arr_add_19_10, 
      d_arr_add_19_9=>d_arr_add_19_9, d_arr_add_19_8=>d_arr_add_19_8, 
      d_arr_add_19_7=>d_arr_add_19_7, d_arr_add_19_6=>d_arr_add_19_6, 
      d_arr_add_19_5=>d_arr_add_19_5, d_arr_add_19_4=>d_arr_add_19_4, 
      d_arr_add_19_3=>d_arr_add_19_3, d_arr_add_19_2=>d_arr_add_19_2, 
      d_arr_add_19_1=>d_arr_add_19_1, d_arr_add_19_0=>d_arr_add_19_0, 
      d_arr_add_20_31=>d_arr_add_20_31, d_arr_add_20_30=>d_arr_add_20_30, 
      d_arr_add_20_29=>d_arr_add_20_29, d_arr_add_20_28=>d_arr_add_20_28, 
      d_arr_add_20_27=>d_arr_add_20_27, d_arr_add_20_26=>d_arr_add_20_26, 
      d_arr_add_20_25=>d_arr_add_20_25, d_arr_add_20_24=>d_arr_add_20_24, 
      d_arr_add_20_23=>d_arr_add_20_23, d_arr_add_20_22=>d_arr_add_20_22, 
      d_arr_add_20_21=>d_arr_add_20_21, d_arr_add_20_20=>d_arr_add_20_20, 
      d_arr_add_20_19=>d_arr_add_20_19, d_arr_add_20_18=>d_arr_add_20_18, 
      d_arr_add_20_17=>d_arr_add_20_17, d_arr_add_20_16=>d_arr_add_20_16, 
      d_arr_add_20_15=>d_arr_add_20_15, d_arr_add_20_14=>d_arr_add_20_14, 
      d_arr_add_20_13=>d_arr_add_20_13, d_arr_add_20_12=>d_arr_add_20_12, 
      d_arr_add_20_11=>d_arr_add_20_11, d_arr_add_20_10=>d_arr_add_20_10, 
      d_arr_add_20_9=>d_arr_add_20_9, d_arr_add_20_8=>d_arr_add_20_8, 
      d_arr_add_20_7=>d_arr_add_20_7, d_arr_add_20_6=>d_arr_add_20_6, 
      d_arr_add_20_5=>d_arr_add_20_5, d_arr_add_20_4=>d_arr_add_20_4, 
      d_arr_add_20_3=>d_arr_add_20_3, d_arr_add_20_2=>d_arr_add_20_2, 
      d_arr_add_20_1=>d_arr_add_20_1, d_arr_add_20_0=>d_arr_add_20_0, 
      d_arr_add_21_31=>q_arr_24_31, d_arr_add_21_30=>q_arr_24_30, 
      d_arr_add_21_29=>q_arr_24_29, d_arr_add_21_28=>q_arr_24_28, 
      d_arr_add_21_27=>q_arr_24_27, d_arr_add_21_26=>q_arr_24_26, 
      d_arr_add_21_25=>q_arr_24_25, d_arr_add_21_24=>q_arr_24_24, 
      d_arr_add_21_23=>q_arr_24_23, d_arr_add_21_22=>q_arr_24_22, 
      d_arr_add_21_21=>q_arr_24_21, d_arr_add_21_20=>q_arr_24_20, 
      d_arr_add_21_19=>q_arr_24_19, d_arr_add_21_18=>q_arr_24_18, 
      d_arr_add_21_17=>q_arr_24_17, d_arr_add_21_16=>q_arr_24_16, 
      d_arr_add_21_15=>q_arr_24_15, d_arr_add_21_14=>q_arr_24_14, 
      d_arr_add_21_13=>q_arr_24_13, d_arr_add_21_12=>q_arr_24_12, 
      d_arr_add_21_11=>q_arr_24_11, d_arr_add_21_10=>q_arr_24_10, 
      d_arr_add_21_9=>q_arr_24_9, d_arr_add_21_8=>q_arr_24_8, d_arr_add_21_7
      =>q_arr_24_7, d_arr_add_21_6=>q_arr_24_6, d_arr_add_21_5=>q_arr_24_5, 
      d_arr_add_21_4=>q_arr_24_4, d_arr_add_21_3=>q_arr_24_3, d_arr_add_21_2
      =>q_arr_24_2, d_arr_add_21_1=>q_arr_24_1, d_arr_add_21_0=>q_arr_24_0, 
      d_arr_add_22_31=>GND0, d_arr_add_22_30=>GND0, d_arr_add_22_29=>GND0, 
      d_arr_add_22_28=>GND0, d_arr_add_22_27=>GND0, d_arr_add_22_26=>GND0, 
      d_arr_add_22_25=>GND0, d_arr_add_22_24=>GND0, d_arr_add_22_23=>GND0, 
      d_arr_add_22_22=>GND0, d_arr_add_22_21=>GND0, d_arr_add_22_20=>GND0, 
      d_arr_add_22_19=>GND0, d_arr_add_22_18=>GND0, d_arr_add_22_17=>GND0, 
      d_arr_add_22_16=>GND0, d_arr_add_22_15=>GND0, d_arr_add_22_14=>GND0, 
      d_arr_add_22_13=>GND0, d_arr_add_22_12=>GND0, d_arr_add_22_11=>GND0, 
      d_arr_add_22_10=>GND0, d_arr_add_22_9=>GND0, d_arr_add_22_8=>GND0, 
      d_arr_add_22_7=>GND0, d_arr_add_22_6=>GND0, d_arr_add_22_5=>GND0, 
      d_arr_add_22_4=>GND0, d_arr_add_22_3=>GND0, d_arr_add_22_2=>GND0, 
      d_arr_add_22_1=>GND0, d_arr_add_22_0=>GND0, d_arr_add_23_31=>GND0, 
      d_arr_add_23_30=>GND0, d_arr_add_23_29=>GND0, d_arr_add_23_28=>GND0, 
      d_arr_add_23_27=>GND0, d_arr_add_23_26=>GND0, d_arr_add_23_25=>GND0, 
      d_arr_add_23_24=>GND0, d_arr_add_23_23=>GND0, d_arr_add_23_22=>GND0, 
      d_arr_add_23_21=>GND0, d_arr_add_23_20=>GND0, d_arr_add_23_19=>GND0, 
      d_arr_add_23_18=>GND0, d_arr_add_23_17=>GND0, d_arr_add_23_16=>GND0, 
      d_arr_add_23_15=>GND0, d_arr_add_23_14=>GND0, d_arr_add_23_13=>GND0, 
      d_arr_add_23_12=>GND0, d_arr_add_23_11=>GND0, d_arr_add_23_10=>GND0, 
      d_arr_add_23_9=>GND0, d_arr_add_23_8=>GND0, d_arr_add_23_7=>GND0, 
      d_arr_add_23_6=>GND0, d_arr_add_23_5=>GND0, d_arr_add_23_4=>GND0, 
      d_arr_add_23_3=>GND0, d_arr_add_23_2=>GND0, d_arr_add_23_1=>GND0, 
      d_arr_add_23_0=>GND0, d_arr_add_24_31=>GND0, d_arr_add_24_30=>GND0, 
      d_arr_add_24_29=>GND0, d_arr_add_24_28=>GND0, d_arr_add_24_27=>GND0, 
      d_arr_add_24_26=>GND0, d_arr_add_24_25=>GND0, d_arr_add_24_24=>GND0, 
      d_arr_add_24_23=>GND0, d_arr_add_24_22=>GND0, d_arr_add_24_21=>GND0, 
      d_arr_add_24_20=>GND0, d_arr_add_24_19=>GND0, d_arr_add_24_18=>GND0, 
      d_arr_add_24_17=>GND0, d_arr_add_24_16=>GND0, d_arr_add_24_15=>GND0, 
      d_arr_add_24_14=>GND0, d_arr_add_24_13=>GND0, d_arr_add_24_12=>GND0, 
      d_arr_add_24_11=>GND0, d_arr_add_24_10=>GND0, d_arr_add_24_9=>GND0, 
      d_arr_add_24_8=>GND0, d_arr_add_24_7=>GND0, d_arr_add_24_6=>GND0, 
      d_arr_add_24_5=>GND0, d_arr_add_24_4=>GND0, d_arr_add_24_3=>GND0, 
      d_arr_add_24_2=>GND0, d_arr_add_24_1=>GND0, d_arr_add_24_0=>GND0, 
      d_arr_merge1_0_31=>d_arr_merge1_0_31, d_arr_merge1_0_30=>
      d_arr_merge1_0_30, d_arr_merge1_0_29=>d_arr_merge1_0_29, 
      d_arr_merge1_0_28=>d_arr_merge1_0_28, d_arr_merge1_0_27=>
      d_arr_merge1_0_27, d_arr_merge1_0_26=>d_arr_merge1_0_26, 
      d_arr_merge1_0_25=>d_arr_merge1_0_25, d_arr_merge1_0_24=>
      d_arr_merge1_0_24, d_arr_merge1_0_23=>d_arr_merge1_0_23, 
      d_arr_merge1_0_22=>d_arr_merge1_0_22, d_arr_merge1_0_21=>
      d_arr_merge1_0_21, d_arr_merge1_0_20=>d_arr_merge1_0_20, 
      d_arr_merge1_0_19=>d_arr_merge1_0_19, d_arr_merge1_0_18=>
      d_arr_merge1_0_18, d_arr_merge1_0_17=>d_arr_merge1_0_17, 
      d_arr_merge1_0_16=>d_arr_merge1_0_16, d_arr_merge1_0_15=>
      d_arr_merge1_0_15, d_arr_merge1_0_14=>d_arr_merge1_0_14, 
      d_arr_merge1_0_13=>d_arr_merge1_0_13, d_arr_merge1_0_12=>
      d_arr_merge1_0_12, d_arr_merge1_0_11=>d_arr_merge1_0_11, 
      d_arr_merge1_0_10=>d_arr_merge1_0_10, d_arr_merge1_0_9=>
      d_arr_merge1_0_9, d_arr_merge1_0_8=>d_arr_merge1_0_8, d_arr_merge1_0_7
      =>d_arr_merge1_0_7, d_arr_merge1_0_6=>d_arr_merge1_0_6, 
      d_arr_merge1_0_5=>d_arr_merge1_0_5, d_arr_merge1_0_4=>d_arr_merge1_0_4, 
      d_arr_merge1_0_3=>d_arr_merge1_0_3, d_arr_merge1_0_2=>d_arr_merge1_0_2, 
      d_arr_merge1_0_1=>d_arr_merge1_0_1, d_arr_merge1_0_0=>d_arr_merge1_0_0, 
      d_arr_merge1_1_31=>d_arr_merge1_1_31, d_arr_merge1_1_30=>
      d_arr_merge1_1_30, d_arr_merge1_1_29=>d_arr_merge1_1_29, 
      d_arr_merge1_1_28=>d_arr_merge1_1_28, d_arr_merge1_1_27=>
      d_arr_merge1_1_27, d_arr_merge1_1_26=>d_arr_merge1_1_26, 
      d_arr_merge1_1_25=>d_arr_merge1_1_25, d_arr_merge1_1_24=>
      d_arr_merge1_1_24, d_arr_merge1_1_23=>d_arr_merge1_1_23, 
      d_arr_merge1_1_22=>d_arr_merge1_1_22, d_arr_merge1_1_21=>
      d_arr_merge1_1_21, d_arr_merge1_1_20=>d_arr_merge1_1_20, 
      d_arr_merge1_1_19=>d_arr_merge1_1_19, d_arr_merge1_1_18=>
      d_arr_merge1_1_18, d_arr_merge1_1_17=>d_arr_merge1_1_17, 
      d_arr_merge1_1_16=>d_arr_merge1_1_16, d_arr_merge1_1_15=>
      d_arr_merge1_1_15, d_arr_merge1_1_14=>d_arr_merge1_1_14, 
      d_arr_merge1_1_13=>d_arr_merge1_1_13, d_arr_merge1_1_12=>
      d_arr_merge1_1_12, d_arr_merge1_1_11=>d_arr_merge1_1_11, 
      d_arr_merge1_1_10=>d_arr_merge1_1_10, d_arr_merge1_1_9=>
      d_arr_merge1_1_9, d_arr_merge1_1_8=>d_arr_merge1_1_8, d_arr_merge1_1_7
      =>d_arr_merge1_1_7, d_arr_merge1_1_6=>d_arr_merge1_1_6, 
      d_arr_merge1_1_5=>d_arr_merge1_1_5, d_arr_merge1_1_4=>d_arr_merge1_1_4, 
      d_arr_merge1_1_3=>d_arr_merge1_1_3, d_arr_merge1_1_2=>d_arr_merge1_1_2, 
      d_arr_merge1_1_1=>d_arr_merge1_1_1, d_arr_merge1_1_0=>d_arr_merge1_1_0, 
      d_arr_merge1_2_31=>GND0, d_arr_merge1_2_30=>GND0, d_arr_merge1_2_29=>
      GND0, d_arr_merge1_2_28=>GND0, d_arr_merge1_2_27=>GND0, 
      d_arr_merge1_2_26=>GND0, d_arr_merge1_2_25=>GND0, d_arr_merge1_2_24=>
      GND0, d_arr_merge1_2_23=>GND0, d_arr_merge1_2_22=>GND0, 
      d_arr_merge1_2_21=>GND0, d_arr_merge1_2_20=>GND0, d_arr_merge1_2_19=>
      GND0, d_arr_merge1_2_18=>GND0, d_arr_merge1_2_17=>GND0, 
      d_arr_merge1_2_16=>GND0, d_arr_merge1_2_15=>GND0, d_arr_merge1_2_14=>
      GND0, d_arr_merge1_2_13=>GND0, d_arr_merge1_2_12=>GND0, 
      d_arr_merge1_2_11=>GND0, d_arr_merge1_2_10=>GND0, d_arr_merge1_2_9=>
      GND0, d_arr_merge1_2_8=>GND0, d_arr_merge1_2_7=>GND0, d_arr_merge1_2_6
      =>GND0, d_arr_merge1_2_5=>GND0, d_arr_merge1_2_4=>GND0, 
      d_arr_merge1_2_3=>GND0, d_arr_merge1_2_2=>GND0, d_arr_merge1_2_1=>GND0, 
      d_arr_merge1_2_0=>GND0, d_arr_merge1_3_31=>GND0, d_arr_merge1_3_30=>
      GND0, d_arr_merge1_3_29=>GND0, d_arr_merge1_3_28=>GND0, 
      d_arr_merge1_3_27=>GND0, d_arr_merge1_3_26=>GND0, d_arr_merge1_3_25=>
      GND0, d_arr_merge1_3_24=>GND0, d_arr_merge1_3_23=>GND0, 
      d_arr_merge1_3_22=>GND0, d_arr_merge1_3_21=>GND0, d_arr_merge1_3_20=>
      GND0, d_arr_merge1_3_19=>GND0, d_arr_merge1_3_18=>GND0, 
      d_arr_merge1_3_17=>GND0, d_arr_merge1_3_16=>GND0, d_arr_merge1_3_15=>
      GND0, d_arr_merge1_3_14=>GND0, d_arr_merge1_3_13=>GND0, 
      d_arr_merge1_3_12=>GND0, d_arr_merge1_3_11=>GND0, d_arr_merge1_3_10=>
      GND0, d_arr_merge1_3_9=>GND0, d_arr_merge1_3_8=>GND0, d_arr_merge1_3_7
      =>GND0, d_arr_merge1_3_6=>GND0, d_arr_merge1_3_5=>GND0, 
      d_arr_merge1_3_4=>GND0, d_arr_merge1_3_3=>GND0, d_arr_merge1_3_2=>GND0, 
      d_arr_merge1_3_1=>GND0, d_arr_merge1_3_0=>GND0, d_arr_merge1_4_31=>
      GND0, d_arr_merge1_4_30=>GND0, d_arr_merge1_4_29=>GND0, 
      d_arr_merge1_4_28=>GND0, d_arr_merge1_4_27=>GND0, d_arr_merge1_4_26=>
      GND0, d_arr_merge1_4_25=>GND0, d_arr_merge1_4_24=>GND0, 
      d_arr_merge1_4_23=>GND0, d_arr_merge1_4_22=>GND0, d_arr_merge1_4_21=>
      GND0, d_arr_merge1_4_20=>GND0, d_arr_merge1_4_19=>GND0, 
      d_arr_merge1_4_18=>GND0, d_arr_merge1_4_17=>GND0, d_arr_merge1_4_16=>
      GND0, d_arr_merge1_4_15=>GND0, d_arr_merge1_4_14=>GND0, 
      d_arr_merge1_4_13=>GND0, d_arr_merge1_4_12=>GND0, d_arr_merge1_4_11=>
      GND0, d_arr_merge1_4_10=>GND0, d_arr_merge1_4_9=>GND0, 
      d_arr_merge1_4_8=>GND0, d_arr_merge1_4_7=>GND0, d_arr_merge1_4_6=>GND0, 
      d_arr_merge1_4_5=>GND0, d_arr_merge1_4_4=>GND0, d_arr_merge1_4_3=>GND0, 
      d_arr_merge1_4_2=>GND0, d_arr_merge1_4_1=>GND0, d_arr_merge1_4_0=>GND0, 
      d_arr_merge1_5_31=>GND0, d_arr_merge1_5_30=>GND0, d_arr_merge1_5_29=>
      GND0, d_arr_merge1_5_28=>GND0, d_arr_merge1_5_27=>GND0, 
      d_arr_merge1_5_26=>GND0, d_arr_merge1_5_25=>GND0, d_arr_merge1_5_24=>
      GND0, d_arr_merge1_5_23=>GND0, d_arr_merge1_5_22=>GND0, 
      d_arr_merge1_5_21=>GND0, d_arr_merge1_5_20=>GND0, d_arr_merge1_5_19=>
      GND0, d_arr_merge1_5_18=>GND0, d_arr_merge1_5_17=>GND0, 
      d_arr_merge1_5_16=>GND0, d_arr_merge1_5_15=>GND0, d_arr_merge1_5_14=>
      GND0, d_arr_merge1_5_13=>GND0, d_arr_merge1_5_12=>GND0, 
      d_arr_merge1_5_11=>GND0, d_arr_merge1_5_10=>GND0, d_arr_merge1_5_9=>
      GND0, d_arr_merge1_5_8=>GND0, d_arr_merge1_5_7=>GND0, d_arr_merge1_5_6
      =>GND0, d_arr_merge1_5_5=>GND0, d_arr_merge1_5_4=>GND0, 
      d_arr_merge1_5_3=>GND0, d_arr_merge1_5_2=>GND0, d_arr_merge1_5_1=>GND0, 
      d_arr_merge1_5_0=>GND0, d_arr_merge1_6_31=>GND0, d_arr_merge1_6_30=>
      GND0, d_arr_merge1_6_29=>GND0, d_arr_merge1_6_28=>GND0, 
      d_arr_merge1_6_27=>GND0, d_arr_merge1_6_26=>GND0, d_arr_merge1_6_25=>
      GND0, d_arr_merge1_6_24=>GND0, d_arr_merge1_6_23=>GND0, 
      d_arr_merge1_6_22=>GND0, d_arr_merge1_6_21=>GND0, d_arr_merge1_6_20=>
      GND0, d_arr_merge1_6_19=>GND0, d_arr_merge1_6_18=>GND0, 
      d_arr_merge1_6_17=>GND0, d_arr_merge1_6_16=>GND0, d_arr_merge1_6_15=>
      GND0, d_arr_merge1_6_14=>GND0, d_arr_merge1_6_13=>GND0, 
      d_arr_merge1_6_12=>GND0, d_arr_merge1_6_11=>GND0, d_arr_merge1_6_10=>
      GND0, d_arr_merge1_6_9=>GND0, d_arr_merge1_6_8=>GND0, d_arr_merge1_6_7
      =>GND0, d_arr_merge1_6_6=>GND0, d_arr_merge1_6_5=>GND0, 
      d_arr_merge1_6_4=>GND0, d_arr_merge1_6_3=>GND0, d_arr_merge1_6_2=>GND0, 
      d_arr_merge1_6_1=>GND0, d_arr_merge1_6_0=>GND0, d_arr_merge1_7_31=>
      GND0, d_arr_merge1_7_30=>GND0, d_arr_merge1_7_29=>GND0, 
      d_arr_merge1_7_28=>GND0, d_arr_merge1_7_27=>GND0, d_arr_merge1_7_26=>
      GND0, d_arr_merge1_7_25=>GND0, d_arr_merge1_7_24=>GND0, 
      d_arr_merge1_7_23=>GND0, d_arr_merge1_7_22=>GND0, d_arr_merge1_7_21=>
      GND0, d_arr_merge1_7_20=>GND0, d_arr_merge1_7_19=>GND0, 
      d_arr_merge1_7_18=>GND0, d_arr_merge1_7_17=>GND0, d_arr_merge1_7_16=>
      GND0, d_arr_merge1_7_15=>GND0, d_arr_merge1_7_14=>GND0, 
      d_arr_merge1_7_13=>GND0, d_arr_merge1_7_12=>GND0, d_arr_merge1_7_11=>
      GND0, d_arr_merge1_7_10=>GND0, d_arr_merge1_7_9=>GND0, 
      d_arr_merge1_7_8=>GND0, d_arr_merge1_7_7=>GND0, d_arr_merge1_7_6=>GND0, 
      d_arr_merge1_7_5=>GND0, d_arr_merge1_7_4=>GND0, d_arr_merge1_7_3=>GND0, 
      d_arr_merge1_7_2=>GND0, d_arr_merge1_7_1=>GND0, d_arr_merge1_7_0=>GND0, 
      d_arr_merge1_8_31=>GND0, d_arr_merge1_8_30=>GND0, d_arr_merge1_8_29=>
      GND0, d_arr_merge1_8_28=>GND0, d_arr_merge1_8_27=>GND0, 
      d_arr_merge1_8_26=>GND0, d_arr_merge1_8_25=>GND0, d_arr_merge1_8_24=>
      GND0, d_arr_merge1_8_23=>GND0, d_arr_merge1_8_22=>GND0, 
      d_arr_merge1_8_21=>GND0, d_arr_merge1_8_20=>GND0, d_arr_merge1_8_19=>
      GND0, d_arr_merge1_8_18=>GND0, d_arr_merge1_8_17=>GND0, 
      d_arr_merge1_8_16=>GND0, d_arr_merge1_8_15=>GND0, d_arr_merge1_8_14=>
      GND0, d_arr_merge1_8_13=>GND0, d_arr_merge1_8_12=>GND0, 
      d_arr_merge1_8_11=>GND0, d_arr_merge1_8_10=>GND0, d_arr_merge1_8_9=>
      GND0, d_arr_merge1_8_8=>GND0, d_arr_merge1_8_7=>GND0, d_arr_merge1_8_6
      =>GND0, d_arr_merge1_8_5=>GND0, d_arr_merge1_8_4=>GND0, 
      d_arr_merge1_8_3=>GND0, d_arr_merge1_8_2=>GND0, d_arr_merge1_8_1=>GND0, 
      d_arr_merge1_8_0=>GND0, d_arr_merge1_9_31=>GND0, d_arr_merge1_9_30=>
      GND0, d_arr_merge1_9_29=>GND0, d_arr_merge1_9_28=>GND0, 
      d_arr_merge1_9_27=>GND0, d_arr_merge1_9_26=>GND0, d_arr_merge1_9_25=>
      GND0, d_arr_merge1_9_24=>GND0, d_arr_merge1_9_23=>GND0, 
      d_arr_merge1_9_22=>GND0, d_arr_merge1_9_21=>GND0, d_arr_merge1_9_20=>
      GND0, d_arr_merge1_9_19=>GND0, d_arr_merge1_9_18=>GND0, 
      d_arr_merge1_9_17=>GND0, d_arr_merge1_9_16=>GND0, d_arr_merge1_9_15=>
      GND0, d_arr_merge1_9_14=>GND0, d_arr_merge1_9_13=>GND0, 
      d_arr_merge1_9_12=>GND0, d_arr_merge1_9_11=>GND0, d_arr_merge1_9_10=>
      GND0, d_arr_merge1_9_9=>GND0, d_arr_merge1_9_8=>GND0, d_arr_merge1_9_7
      =>GND0, d_arr_merge1_9_6=>GND0, d_arr_merge1_9_5=>GND0, 
      d_arr_merge1_9_4=>GND0, d_arr_merge1_9_3=>GND0, d_arr_merge1_9_2=>GND0, 
      d_arr_merge1_9_1=>GND0, d_arr_merge1_9_0=>GND0, d_arr_merge1_10_31=>
      GND0, d_arr_merge1_10_30=>GND0, d_arr_merge1_10_29=>GND0, 
      d_arr_merge1_10_28=>GND0, d_arr_merge1_10_27=>GND0, d_arr_merge1_10_26
      =>GND0, d_arr_merge1_10_25=>GND0, d_arr_merge1_10_24=>GND0, 
      d_arr_merge1_10_23=>GND0, d_arr_merge1_10_22=>GND0, d_arr_merge1_10_21
      =>GND0, d_arr_merge1_10_20=>GND0, d_arr_merge1_10_19=>GND0, 
      d_arr_merge1_10_18=>GND0, d_arr_merge1_10_17=>GND0, d_arr_merge1_10_16
      =>GND0, d_arr_merge1_10_15=>GND0, d_arr_merge1_10_14=>GND0, 
      d_arr_merge1_10_13=>GND0, d_arr_merge1_10_12=>GND0, d_arr_merge1_10_11
      =>GND0, d_arr_merge1_10_10=>GND0, d_arr_merge1_10_9=>GND0, 
      d_arr_merge1_10_8=>GND0, d_arr_merge1_10_7=>GND0, d_arr_merge1_10_6=>
      GND0, d_arr_merge1_10_5=>GND0, d_arr_merge1_10_4=>GND0, 
      d_arr_merge1_10_3=>GND0, d_arr_merge1_10_2=>GND0, d_arr_merge1_10_1=>
      GND0, d_arr_merge1_10_0=>GND0, d_arr_merge1_11_31=>GND0, 
      d_arr_merge1_11_30=>GND0, d_arr_merge1_11_29=>GND0, d_arr_merge1_11_28
      =>GND0, d_arr_merge1_11_27=>GND0, d_arr_merge1_11_26=>GND0, 
      d_arr_merge1_11_25=>GND0, d_arr_merge1_11_24=>GND0, d_arr_merge1_11_23
      =>GND0, d_arr_merge1_11_22=>GND0, d_arr_merge1_11_21=>GND0, 
      d_arr_merge1_11_20=>GND0, d_arr_merge1_11_19=>GND0, d_arr_merge1_11_18
      =>GND0, d_arr_merge1_11_17=>GND0, d_arr_merge1_11_16=>GND0, 
      d_arr_merge1_11_15=>GND0, d_arr_merge1_11_14=>GND0, d_arr_merge1_11_13
      =>GND0, d_arr_merge1_11_12=>GND0, d_arr_merge1_11_11=>GND0, 
      d_arr_merge1_11_10=>GND0, d_arr_merge1_11_9=>GND0, d_arr_merge1_11_8=>
      GND0, d_arr_merge1_11_7=>GND0, d_arr_merge1_11_6=>GND0, 
      d_arr_merge1_11_5=>GND0, d_arr_merge1_11_4=>GND0, d_arr_merge1_11_3=>
      GND0, d_arr_merge1_11_2=>GND0, d_arr_merge1_11_1=>GND0, 
      d_arr_merge1_11_0=>GND0, d_arr_merge1_12_31=>GND0, d_arr_merge1_12_30
      =>GND0, d_arr_merge1_12_29=>GND0, d_arr_merge1_12_28=>GND0, 
      d_arr_merge1_12_27=>GND0, d_arr_merge1_12_26=>GND0, d_arr_merge1_12_25
      =>GND0, d_arr_merge1_12_24=>GND0, d_arr_merge1_12_23=>GND0, 
      d_arr_merge1_12_22=>GND0, d_arr_merge1_12_21=>GND0, d_arr_merge1_12_20
      =>GND0, d_arr_merge1_12_19=>GND0, d_arr_merge1_12_18=>GND0, 
      d_arr_merge1_12_17=>GND0, d_arr_merge1_12_16=>GND0, d_arr_merge1_12_15
      =>GND0, d_arr_merge1_12_14=>GND0, d_arr_merge1_12_13=>GND0, 
      d_arr_merge1_12_12=>GND0, d_arr_merge1_12_11=>GND0, d_arr_merge1_12_10
      =>GND0, d_arr_merge1_12_9=>GND0, d_arr_merge1_12_8=>GND0, 
      d_arr_merge1_12_7=>GND0, d_arr_merge1_12_6=>GND0, d_arr_merge1_12_5=>
      GND0, d_arr_merge1_12_4=>GND0, d_arr_merge1_12_3=>GND0, 
      d_arr_merge1_12_2=>GND0, d_arr_merge1_12_1=>GND0, d_arr_merge1_12_0=>
      GND0, d_arr_merge1_13_31=>GND0, d_arr_merge1_13_30=>GND0, 
      d_arr_merge1_13_29=>GND0, d_arr_merge1_13_28=>GND0, d_arr_merge1_13_27
      =>GND0, d_arr_merge1_13_26=>GND0, d_arr_merge1_13_25=>GND0, 
      d_arr_merge1_13_24=>GND0, d_arr_merge1_13_23=>GND0, d_arr_merge1_13_22
      =>GND0, d_arr_merge1_13_21=>GND0, d_arr_merge1_13_20=>GND0, 
      d_arr_merge1_13_19=>GND0, d_arr_merge1_13_18=>GND0, d_arr_merge1_13_17
      =>GND0, d_arr_merge1_13_16=>GND0, d_arr_merge1_13_15=>GND0, 
      d_arr_merge1_13_14=>GND0, d_arr_merge1_13_13=>GND0, d_arr_merge1_13_12
      =>GND0, d_arr_merge1_13_11=>GND0, d_arr_merge1_13_10=>GND0, 
      d_arr_merge1_13_9=>GND0, d_arr_merge1_13_8=>GND0, d_arr_merge1_13_7=>
      GND0, d_arr_merge1_13_6=>GND0, d_arr_merge1_13_5=>GND0, 
      d_arr_merge1_13_4=>GND0, d_arr_merge1_13_3=>GND0, d_arr_merge1_13_2=>
      GND0, d_arr_merge1_13_1=>GND0, d_arr_merge1_13_0=>GND0, 
      d_arr_merge1_14_31=>GND0, d_arr_merge1_14_30=>GND0, d_arr_merge1_14_29
      =>GND0, d_arr_merge1_14_28=>GND0, d_arr_merge1_14_27=>GND0, 
      d_arr_merge1_14_26=>GND0, d_arr_merge1_14_25=>GND0, d_arr_merge1_14_24
      =>GND0, d_arr_merge1_14_23=>GND0, d_arr_merge1_14_22=>GND0, 
      d_arr_merge1_14_21=>GND0, d_arr_merge1_14_20=>GND0, d_arr_merge1_14_19
      =>GND0, d_arr_merge1_14_18=>GND0, d_arr_merge1_14_17=>GND0, 
      d_arr_merge1_14_16=>GND0, d_arr_merge1_14_15=>GND0, d_arr_merge1_14_14
      =>GND0, d_arr_merge1_14_13=>GND0, d_arr_merge1_14_12=>GND0, 
      d_arr_merge1_14_11=>GND0, d_arr_merge1_14_10=>GND0, d_arr_merge1_14_9
      =>GND0, d_arr_merge1_14_8=>GND0, d_arr_merge1_14_7=>GND0, 
      d_arr_merge1_14_6=>GND0, d_arr_merge1_14_5=>GND0, d_arr_merge1_14_4=>
      GND0, d_arr_merge1_14_3=>GND0, d_arr_merge1_14_2=>GND0, 
      d_arr_merge1_14_1=>GND0, d_arr_merge1_14_0=>GND0, d_arr_merge1_15_31=>
      GND0, d_arr_merge1_15_30=>GND0, d_arr_merge1_15_29=>GND0, 
      d_arr_merge1_15_28=>GND0, d_arr_merge1_15_27=>GND0, d_arr_merge1_15_26
      =>GND0, d_arr_merge1_15_25=>GND0, d_arr_merge1_15_24=>GND0, 
      d_arr_merge1_15_23=>GND0, d_arr_merge1_15_22=>GND0, d_arr_merge1_15_21
      =>GND0, d_arr_merge1_15_20=>GND0, d_arr_merge1_15_19=>GND0, 
      d_arr_merge1_15_18=>GND0, d_arr_merge1_15_17=>GND0, d_arr_merge1_15_16
      =>GND0, d_arr_merge1_15_15=>GND0, d_arr_merge1_15_14=>GND0, 
      d_arr_merge1_15_13=>GND0, d_arr_merge1_15_12=>GND0, d_arr_merge1_15_11
      =>GND0, d_arr_merge1_15_10=>GND0, d_arr_merge1_15_9=>GND0, 
      d_arr_merge1_15_8=>GND0, d_arr_merge1_15_7=>GND0, d_arr_merge1_15_6=>
      GND0, d_arr_merge1_15_5=>GND0, d_arr_merge1_15_4=>GND0, 
      d_arr_merge1_15_3=>GND0, d_arr_merge1_15_2=>GND0, d_arr_merge1_15_1=>
      GND0, d_arr_merge1_15_0=>GND0, d_arr_merge1_16_31=>GND0, 
      d_arr_merge1_16_30=>GND0, d_arr_merge1_16_29=>GND0, d_arr_merge1_16_28
      =>GND0, d_arr_merge1_16_27=>GND0, d_arr_merge1_16_26=>GND0, 
      d_arr_merge1_16_25=>GND0, d_arr_merge1_16_24=>GND0, d_arr_merge1_16_23
      =>GND0, d_arr_merge1_16_22=>GND0, d_arr_merge1_16_21=>GND0, 
      d_arr_merge1_16_20=>GND0, d_arr_merge1_16_19=>GND0, d_arr_merge1_16_18
      =>GND0, d_arr_merge1_16_17=>GND0, d_arr_merge1_16_16=>GND0, 
      d_arr_merge1_16_15=>GND0, d_arr_merge1_16_14=>GND0, d_arr_merge1_16_13
      =>GND0, d_arr_merge1_16_12=>GND0, d_arr_merge1_16_11=>GND0, 
      d_arr_merge1_16_10=>GND0, d_arr_merge1_16_9=>GND0, d_arr_merge1_16_8=>
      GND0, d_arr_merge1_16_7=>GND0, d_arr_merge1_16_6=>GND0, 
      d_arr_merge1_16_5=>GND0, d_arr_merge1_16_4=>GND0, d_arr_merge1_16_3=>
      GND0, d_arr_merge1_16_2=>GND0, d_arr_merge1_16_1=>GND0, 
      d_arr_merge1_16_0=>GND0, d_arr_merge1_17_31=>GND0, d_arr_merge1_17_30
      =>GND0, d_arr_merge1_17_29=>GND0, d_arr_merge1_17_28=>GND0, 
      d_arr_merge1_17_27=>GND0, d_arr_merge1_17_26=>GND0, d_arr_merge1_17_25
      =>GND0, d_arr_merge1_17_24=>GND0, d_arr_merge1_17_23=>GND0, 
      d_arr_merge1_17_22=>GND0, d_arr_merge1_17_21=>GND0, d_arr_merge1_17_20
      =>GND0, d_arr_merge1_17_19=>GND0, d_arr_merge1_17_18=>GND0, 
      d_arr_merge1_17_17=>GND0, d_arr_merge1_17_16=>GND0, d_arr_merge1_17_15
      =>GND0, d_arr_merge1_17_14=>GND0, d_arr_merge1_17_13=>GND0, 
      d_arr_merge1_17_12=>GND0, d_arr_merge1_17_11=>GND0, d_arr_merge1_17_10
      =>GND0, d_arr_merge1_17_9=>GND0, d_arr_merge1_17_8=>GND0, 
      d_arr_merge1_17_7=>GND0, d_arr_merge1_17_6=>GND0, d_arr_merge1_17_5=>
      GND0, d_arr_merge1_17_4=>GND0, d_arr_merge1_17_3=>GND0, 
      d_arr_merge1_17_2=>GND0, d_arr_merge1_17_1=>GND0, d_arr_merge1_17_0=>
      GND0, d_arr_merge1_18_31=>GND0, d_arr_merge1_18_30=>GND0, 
      d_arr_merge1_18_29=>GND0, d_arr_merge1_18_28=>GND0, d_arr_merge1_18_27
      =>GND0, d_arr_merge1_18_26=>GND0, d_arr_merge1_18_25=>GND0, 
      d_arr_merge1_18_24=>GND0, d_arr_merge1_18_23=>GND0, d_arr_merge1_18_22
      =>GND0, d_arr_merge1_18_21=>GND0, d_arr_merge1_18_20=>GND0, 
      d_arr_merge1_18_19=>GND0, d_arr_merge1_18_18=>GND0, d_arr_merge1_18_17
      =>GND0, d_arr_merge1_18_16=>GND0, d_arr_merge1_18_15=>GND0, 
      d_arr_merge1_18_14=>GND0, d_arr_merge1_18_13=>GND0, d_arr_merge1_18_12
      =>GND0, d_arr_merge1_18_11=>GND0, d_arr_merge1_18_10=>GND0, 
      d_arr_merge1_18_9=>GND0, d_arr_merge1_18_8=>GND0, d_arr_merge1_18_7=>
      GND0, d_arr_merge1_18_6=>GND0, d_arr_merge1_18_5=>GND0, 
      d_arr_merge1_18_4=>GND0, d_arr_merge1_18_3=>GND0, d_arr_merge1_18_2=>
      GND0, d_arr_merge1_18_1=>GND0, d_arr_merge1_18_0=>GND0, 
      d_arr_merge1_19_31=>GND0, d_arr_merge1_19_30=>GND0, d_arr_merge1_19_29
      =>GND0, d_arr_merge1_19_28=>GND0, d_arr_merge1_19_27=>GND0, 
      d_arr_merge1_19_26=>GND0, d_arr_merge1_19_25=>GND0, d_arr_merge1_19_24
      =>GND0, d_arr_merge1_19_23=>GND0, d_arr_merge1_19_22=>GND0, 
      d_arr_merge1_19_21=>GND0, d_arr_merge1_19_20=>GND0, d_arr_merge1_19_19
      =>GND0, d_arr_merge1_19_18=>GND0, d_arr_merge1_19_17=>GND0, 
      d_arr_merge1_19_16=>GND0, d_arr_merge1_19_15=>GND0, d_arr_merge1_19_14
      =>GND0, d_arr_merge1_19_13=>GND0, d_arr_merge1_19_12=>GND0, 
      d_arr_merge1_19_11=>GND0, d_arr_merge1_19_10=>GND0, d_arr_merge1_19_9
      =>GND0, d_arr_merge1_19_8=>GND0, d_arr_merge1_19_7=>GND0, 
      d_arr_merge1_19_6=>GND0, d_arr_merge1_19_5=>GND0, d_arr_merge1_19_4=>
      GND0, d_arr_merge1_19_3=>GND0, d_arr_merge1_19_2=>GND0, 
      d_arr_merge1_19_1=>GND0, d_arr_merge1_19_0=>GND0, d_arr_merge1_20_31=>
      GND0, d_arr_merge1_20_30=>GND0, d_arr_merge1_20_29=>GND0, 
      d_arr_merge1_20_28=>GND0, d_arr_merge1_20_27=>GND0, d_arr_merge1_20_26
      =>GND0, d_arr_merge1_20_25=>GND0, d_arr_merge1_20_24=>GND0, 
      d_arr_merge1_20_23=>GND0, d_arr_merge1_20_22=>GND0, d_arr_merge1_20_21
      =>GND0, d_arr_merge1_20_20=>GND0, d_arr_merge1_20_19=>GND0, 
      d_arr_merge1_20_18=>GND0, d_arr_merge1_20_17=>GND0, d_arr_merge1_20_16
      =>GND0, d_arr_merge1_20_15=>GND0, d_arr_merge1_20_14=>GND0, 
      d_arr_merge1_20_13=>GND0, d_arr_merge1_20_12=>GND0, d_arr_merge1_20_11
      =>GND0, d_arr_merge1_20_10=>GND0, d_arr_merge1_20_9=>GND0, 
      d_arr_merge1_20_8=>GND0, d_arr_merge1_20_7=>GND0, d_arr_merge1_20_6=>
      GND0, d_arr_merge1_20_5=>GND0, d_arr_merge1_20_4=>GND0, 
      d_arr_merge1_20_3=>GND0, d_arr_merge1_20_2=>GND0, d_arr_merge1_20_1=>
      GND0, d_arr_merge1_20_0=>GND0, d_arr_merge1_21_31=>GND0, 
      d_arr_merge1_21_30=>GND0, d_arr_merge1_21_29=>GND0, d_arr_merge1_21_28
      =>GND0, d_arr_merge1_21_27=>GND0, d_arr_merge1_21_26=>GND0, 
      d_arr_merge1_21_25=>GND0, d_arr_merge1_21_24=>GND0, d_arr_merge1_21_23
      =>GND0, d_arr_merge1_21_22=>GND0, d_arr_merge1_21_21=>GND0, 
      d_arr_merge1_21_20=>GND0, d_arr_merge1_21_19=>GND0, d_arr_merge1_21_18
      =>GND0, d_arr_merge1_21_17=>GND0, d_arr_merge1_21_16=>GND0, 
      d_arr_merge1_21_15=>GND0, d_arr_merge1_21_14=>GND0, d_arr_merge1_21_13
      =>GND0, d_arr_merge1_21_12=>GND0, d_arr_merge1_21_11=>GND0, 
      d_arr_merge1_21_10=>GND0, d_arr_merge1_21_9=>GND0, d_arr_merge1_21_8=>
      GND0, d_arr_merge1_21_7=>GND0, d_arr_merge1_21_6=>GND0, 
      d_arr_merge1_21_5=>GND0, d_arr_merge1_21_4=>GND0, d_arr_merge1_21_3=>
      GND0, d_arr_merge1_21_2=>GND0, d_arr_merge1_21_1=>GND0, 
      d_arr_merge1_21_0=>GND0, d_arr_merge1_22_31=>GND0, d_arr_merge1_22_30
      =>GND0, d_arr_merge1_22_29=>GND0, d_arr_merge1_22_28=>GND0, 
      d_arr_merge1_22_27=>GND0, d_arr_merge1_22_26=>GND0, d_arr_merge1_22_25
      =>GND0, d_arr_merge1_22_24=>GND0, d_arr_merge1_22_23=>GND0, 
      d_arr_merge1_22_22=>GND0, d_arr_merge1_22_21=>GND0, d_arr_merge1_22_20
      =>GND0, d_arr_merge1_22_19=>GND0, d_arr_merge1_22_18=>GND0, 
      d_arr_merge1_22_17=>GND0, d_arr_merge1_22_16=>GND0, d_arr_merge1_22_15
      =>GND0, d_arr_merge1_22_14=>GND0, d_arr_merge1_22_13=>GND0, 
      d_arr_merge1_22_12=>GND0, d_arr_merge1_22_11=>GND0, d_arr_merge1_22_10
      =>GND0, d_arr_merge1_22_9=>GND0, d_arr_merge1_22_8=>GND0, 
      d_arr_merge1_22_7=>GND0, d_arr_merge1_22_6=>GND0, d_arr_merge1_22_5=>
      GND0, d_arr_merge1_22_4=>GND0, d_arr_merge1_22_3=>GND0, 
      d_arr_merge1_22_2=>GND0, d_arr_merge1_22_1=>GND0, d_arr_merge1_22_0=>
      GND0, d_arr_merge1_23_31=>GND0, d_arr_merge1_23_30=>GND0, 
      d_arr_merge1_23_29=>GND0, d_arr_merge1_23_28=>GND0, d_arr_merge1_23_27
      =>GND0, d_arr_merge1_23_26=>GND0, d_arr_merge1_23_25=>GND0, 
      d_arr_merge1_23_24=>GND0, d_arr_merge1_23_23=>GND0, d_arr_merge1_23_22
      =>GND0, d_arr_merge1_23_21=>GND0, d_arr_merge1_23_20=>GND0, 
      d_arr_merge1_23_19=>GND0, d_arr_merge1_23_18=>GND0, d_arr_merge1_23_17
      =>GND0, d_arr_merge1_23_16=>GND0, d_arr_merge1_23_15=>GND0, 
      d_arr_merge1_23_14=>GND0, d_arr_merge1_23_13=>GND0, d_arr_merge1_23_12
      =>GND0, d_arr_merge1_23_11=>GND0, d_arr_merge1_23_10=>GND0, 
      d_arr_merge1_23_9=>GND0, d_arr_merge1_23_8=>GND0, d_arr_merge1_23_7=>
      GND0, d_arr_merge1_23_6=>GND0, d_arr_merge1_23_5=>GND0, 
      d_arr_merge1_23_4=>GND0, d_arr_merge1_23_3=>GND0, d_arr_merge1_23_2=>
      GND0, d_arr_merge1_23_1=>GND0, d_arr_merge1_23_0=>GND0, 
      d_arr_merge1_24_31=>GND0, d_arr_merge1_24_30=>GND0, d_arr_merge1_24_29
      =>GND0, d_arr_merge1_24_28=>GND0, d_arr_merge1_24_27=>GND0, 
      d_arr_merge1_24_26=>GND0, d_arr_merge1_24_25=>GND0, d_arr_merge1_24_24
      =>GND0, d_arr_merge1_24_23=>GND0, d_arr_merge1_24_22=>GND0, 
      d_arr_merge1_24_21=>GND0, d_arr_merge1_24_20=>GND0, d_arr_merge1_24_19
      =>GND0, d_arr_merge1_24_18=>GND0, d_arr_merge1_24_17=>GND0, 
      d_arr_merge1_24_16=>GND0, d_arr_merge1_24_15=>GND0, d_arr_merge1_24_14
      =>GND0, d_arr_merge1_24_13=>GND0, d_arr_merge1_24_12=>GND0, 
      d_arr_merge1_24_11=>GND0, d_arr_merge1_24_10=>GND0, d_arr_merge1_24_9
      =>GND0, d_arr_merge1_24_8=>GND0, d_arr_merge1_24_7=>GND0, 
      d_arr_merge1_24_6=>GND0, d_arr_merge1_24_5=>GND0, d_arr_merge1_24_4=>
      GND0, d_arr_merge1_24_3=>GND0, d_arr_merge1_24_2=>GND0, 
      d_arr_merge1_24_1=>GND0, d_arr_merge1_24_0=>GND0, d_arr_merge2_0_31=>
      d_arr_merge2_0_31, d_arr_merge2_0_30=>d_arr_merge2_0_31, 
      d_arr_merge2_0_29=>d_arr_merge2_0_31, d_arr_merge2_0_28=>
      d_arr_merge2_0_31, d_arr_merge2_0_27=>d_arr_merge2_0_31, 
      d_arr_merge2_0_26=>d_arr_merge2_0_26, d_arr_merge2_0_25=>
      d_arr_merge2_0_25, d_arr_merge2_0_24=>d_arr_merge2_0_24, 
      d_arr_merge2_0_23=>d_arr_merge2_0_23, d_arr_merge2_0_22=>
      d_arr_merge2_0_22, d_arr_merge2_0_21=>d_arr_merge2_0_21, 
      d_arr_merge2_0_20=>d_arr_merge2_0_20, d_arr_merge2_0_19=>
      d_arr_merge2_0_19, d_arr_merge2_0_18=>d_arr_merge2_0_18, 
      d_arr_merge2_0_17=>d_arr_merge2_0_17, d_arr_merge2_0_16=>
      d_arr_merge2_0_16, d_arr_merge2_0_15=>d_arr_merge2_0_15, 
      d_arr_merge2_0_14=>d_arr_merge2_0_14, d_arr_merge2_0_13=>
      d_arr_merge2_0_13, d_arr_merge2_0_12=>d_arr_merge2_0_12, 
      d_arr_merge2_0_11=>d_arr_merge2_0_11, d_arr_merge2_0_10=>
      d_arr_merge2_0_10, d_arr_merge2_0_9=>d_arr_merge2_0_9, 
      d_arr_merge2_0_8=>d_arr_merge2_0_8, d_arr_merge2_0_7=>d_arr_merge2_0_7, 
      d_arr_merge2_0_6=>d_arr_merge2_0_6, d_arr_merge2_0_5=>d_arr_merge2_0_5, 
      d_arr_merge2_0_4=>d_arr_merge2_0_4, d_arr_merge2_0_3=>d_arr_merge2_0_3, 
      d_arr_merge2_0_2=>d_arr_merge2_0_2, d_arr_merge2_0_1=>d_arr_merge2_0_1, 
      d_arr_merge2_0_0=>d_arr_merge2_0_0, d_arr_merge2_1_31=>
      d_arr_merge2_1_31, d_arr_merge2_1_30=>d_arr_merge2_1_31, 
      d_arr_merge2_1_29=>d_arr_merge2_1_31, d_arr_merge2_1_28=>
      d_arr_merge2_1_31, d_arr_merge2_1_27=>d_arr_merge2_1_31, 
      d_arr_merge2_1_26=>d_arr_merge2_1_26, d_arr_merge2_1_25=>
      d_arr_merge2_1_25, d_arr_merge2_1_24=>d_arr_merge2_1_24, 
      d_arr_merge2_1_23=>d_arr_merge2_1_23, d_arr_merge2_1_22=>
      d_arr_merge2_1_22, d_arr_merge2_1_21=>d_arr_merge2_1_21, 
      d_arr_merge2_1_20=>d_arr_merge2_1_20, d_arr_merge2_1_19=>
      d_arr_merge2_1_19, d_arr_merge2_1_18=>d_arr_merge2_1_18, 
      d_arr_merge2_1_17=>d_arr_merge2_1_17, d_arr_merge2_1_16=>
      d_arr_merge2_1_16, d_arr_merge2_1_15=>d_arr_merge2_1_15, 
      d_arr_merge2_1_14=>d_arr_merge2_1_14, d_arr_merge2_1_13=>
      d_arr_merge2_1_13, d_arr_merge2_1_12=>d_arr_merge2_1_12, 
      d_arr_merge2_1_11=>d_arr_merge2_1_11, d_arr_merge2_1_10=>
      d_arr_merge2_1_10, d_arr_merge2_1_9=>d_arr_merge2_1_9, 
      d_arr_merge2_1_8=>d_arr_merge2_1_8, d_arr_merge2_1_7=>d_arr_merge2_1_7, 
      d_arr_merge2_1_6=>d_arr_merge2_1_6, d_arr_merge2_1_5=>d_arr_merge2_1_5, 
      d_arr_merge2_1_4=>d_arr_merge2_1_4, d_arr_merge2_1_3=>d_arr_merge2_1_3, 
      d_arr_merge2_1_2=>d_arr_merge2_1_2, d_arr_merge2_1_1=>d_arr_merge2_1_1, 
      d_arr_merge2_1_0=>d_arr_merge2_1_0, d_arr_merge2_2_31=>GND0, 
      d_arr_merge2_2_30=>GND0, d_arr_merge2_2_29=>GND0, d_arr_merge2_2_28=>
      GND0, d_arr_merge2_2_27=>GND0, d_arr_merge2_2_26=>GND0, 
      d_arr_merge2_2_25=>GND0, d_arr_merge2_2_24=>GND0, d_arr_merge2_2_23=>
      GND0, d_arr_merge2_2_22=>GND0, d_arr_merge2_2_21=>GND0, 
      d_arr_merge2_2_20=>GND0, d_arr_merge2_2_19=>GND0, d_arr_merge2_2_18=>
      GND0, d_arr_merge2_2_17=>GND0, d_arr_merge2_2_16=>GND0, 
      d_arr_merge2_2_15=>GND0, d_arr_merge2_2_14=>GND0, d_arr_merge2_2_13=>
      GND0, d_arr_merge2_2_12=>GND0, d_arr_merge2_2_11=>GND0, 
      d_arr_merge2_2_10=>GND0, d_arr_merge2_2_9=>GND0, d_arr_merge2_2_8=>
      GND0, d_arr_merge2_2_7=>GND0, d_arr_merge2_2_6=>GND0, d_arr_merge2_2_5
      =>GND0, d_arr_merge2_2_4=>GND0, d_arr_merge2_2_3=>GND0, 
      d_arr_merge2_2_2=>GND0, d_arr_merge2_2_1=>GND0, d_arr_merge2_2_0=>GND0, 
      d_arr_merge2_3_31=>GND0, d_arr_merge2_3_30=>GND0, d_arr_merge2_3_29=>
      GND0, d_arr_merge2_3_28=>GND0, d_arr_merge2_3_27=>GND0, 
      d_arr_merge2_3_26=>GND0, d_arr_merge2_3_25=>GND0, d_arr_merge2_3_24=>
      GND0, d_arr_merge2_3_23=>GND0, d_arr_merge2_3_22=>GND0, 
      d_arr_merge2_3_21=>GND0, d_arr_merge2_3_20=>GND0, d_arr_merge2_3_19=>
      GND0, d_arr_merge2_3_18=>GND0, d_arr_merge2_3_17=>GND0, 
      d_arr_merge2_3_16=>GND0, d_arr_merge2_3_15=>GND0, d_arr_merge2_3_14=>
      GND0, d_arr_merge2_3_13=>GND0, d_arr_merge2_3_12=>GND0, 
      d_arr_merge2_3_11=>GND0, d_arr_merge2_3_10=>GND0, d_arr_merge2_3_9=>
      GND0, d_arr_merge2_3_8=>GND0, d_arr_merge2_3_7=>GND0, d_arr_merge2_3_6
      =>GND0, d_arr_merge2_3_5=>GND0, d_arr_merge2_3_4=>GND0, 
      d_arr_merge2_3_3=>GND0, d_arr_merge2_3_2=>GND0, d_arr_merge2_3_1=>GND0, 
      d_arr_merge2_3_0=>GND0, d_arr_merge2_4_31=>GND0, d_arr_merge2_4_30=>
      GND0, d_arr_merge2_4_29=>GND0, d_arr_merge2_4_28=>GND0, 
      d_arr_merge2_4_27=>GND0, d_arr_merge2_4_26=>GND0, d_arr_merge2_4_25=>
      GND0, d_arr_merge2_4_24=>GND0, d_arr_merge2_4_23=>GND0, 
      d_arr_merge2_4_22=>GND0, d_arr_merge2_4_21=>GND0, d_arr_merge2_4_20=>
      GND0, d_arr_merge2_4_19=>GND0, d_arr_merge2_4_18=>GND0, 
      d_arr_merge2_4_17=>GND0, d_arr_merge2_4_16=>GND0, d_arr_merge2_4_15=>
      GND0, d_arr_merge2_4_14=>GND0, d_arr_merge2_4_13=>GND0, 
      d_arr_merge2_4_12=>GND0, d_arr_merge2_4_11=>GND0, d_arr_merge2_4_10=>
      GND0, d_arr_merge2_4_9=>GND0, d_arr_merge2_4_8=>GND0, d_arr_merge2_4_7
      =>GND0, d_arr_merge2_4_6=>GND0, d_arr_merge2_4_5=>GND0, 
      d_arr_merge2_4_4=>GND0, d_arr_merge2_4_3=>GND0, d_arr_merge2_4_2=>GND0, 
      d_arr_merge2_4_1=>GND0, d_arr_merge2_4_0=>GND0, d_arr_merge2_5_31=>
      GND0, d_arr_merge2_5_30=>GND0, d_arr_merge2_5_29=>GND0, 
      d_arr_merge2_5_28=>GND0, d_arr_merge2_5_27=>GND0, d_arr_merge2_5_26=>
      GND0, d_arr_merge2_5_25=>GND0, d_arr_merge2_5_24=>GND0, 
      d_arr_merge2_5_23=>GND0, d_arr_merge2_5_22=>GND0, d_arr_merge2_5_21=>
      GND0, d_arr_merge2_5_20=>GND0, d_arr_merge2_5_19=>GND0, 
      d_arr_merge2_5_18=>GND0, d_arr_merge2_5_17=>GND0, d_arr_merge2_5_16=>
      GND0, d_arr_merge2_5_15=>GND0, d_arr_merge2_5_14=>GND0, 
      d_arr_merge2_5_13=>GND0, d_arr_merge2_5_12=>GND0, d_arr_merge2_5_11=>
      GND0, d_arr_merge2_5_10=>GND0, d_arr_merge2_5_9=>GND0, 
      d_arr_merge2_5_8=>GND0, d_arr_merge2_5_7=>GND0, d_arr_merge2_5_6=>GND0, 
      d_arr_merge2_5_5=>GND0, d_arr_merge2_5_4=>GND0, d_arr_merge2_5_3=>GND0, 
      d_arr_merge2_5_2=>GND0, d_arr_merge2_5_1=>GND0, d_arr_merge2_5_0=>GND0, 
      d_arr_merge2_6_31=>GND0, d_arr_merge2_6_30=>GND0, d_arr_merge2_6_29=>
      GND0, d_arr_merge2_6_28=>GND0, d_arr_merge2_6_27=>GND0, 
      d_arr_merge2_6_26=>GND0, d_arr_merge2_6_25=>GND0, d_arr_merge2_6_24=>
      GND0, d_arr_merge2_6_23=>GND0, d_arr_merge2_6_22=>GND0, 
      d_arr_merge2_6_21=>GND0, d_arr_merge2_6_20=>GND0, d_arr_merge2_6_19=>
      GND0, d_arr_merge2_6_18=>GND0, d_arr_merge2_6_17=>GND0, 
      d_arr_merge2_6_16=>GND0, d_arr_merge2_6_15=>GND0, d_arr_merge2_6_14=>
      GND0, d_arr_merge2_6_13=>GND0, d_arr_merge2_6_12=>GND0, 
      d_arr_merge2_6_11=>GND0, d_arr_merge2_6_10=>GND0, d_arr_merge2_6_9=>
      GND0, d_arr_merge2_6_8=>GND0, d_arr_merge2_6_7=>GND0, d_arr_merge2_6_6
      =>GND0, d_arr_merge2_6_5=>GND0, d_arr_merge2_6_4=>GND0, 
      d_arr_merge2_6_3=>GND0, d_arr_merge2_6_2=>GND0, d_arr_merge2_6_1=>GND0, 
      d_arr_merge2_6_0=>GND0, d_arr_merge2_7_31=>GND0, d_arr_merge2_7_30=>
      GND0, d_arr_merge2_7_29=>GND0, d_arr_merge2_7_28=>GND0, 
      d_arr_merge2_7_27=>GND0, d_arr_merge2_7_26=>GND0, d_arr_merge2_7_25=>
      GND0, d_arr_merge2_7_24=>GND0, d_arr_merge2_7_23=>GND0, 
      d_arr_merge2_7_22=>GND0, d_arr_merge2_7_21=>GND0, d_arr_merge2_7_20=>
      GND0, d_arr_merge2_7_19=>GND0, d_arr_merge2_7_18=>GND0, 
      d_arr_merge2_7_17=>GND0, d_arr_merge2_7_16=>GND0, d_arr_merge2_7_15=>
      GND0, d_arr_merge2_7_14=>GND0, d_arr_merge2_7_13=>GND0, 
      d_arr_merge2_7_12=>GND0, d_arr_merge2_7_11=>GND0, d_arr_merge2_7_10=>
      GND0, d_arr_merge2_7_9=>GND0, d_arr_merge2_7_8=>GND0, d_arr_merge2_7_7
      =>GND0, d_arr_merge2_7_6=>GND0, d_arr_merge2_7_5=>GND0, 
      d_arr_merge2_7_4=>GND0, d_arr_merge2_7_3=>GND0, d_arr_merge2_7_2=>GND0, 
      d_arr_merge2_7_1=>GND0, d_arr_merge2_7_0=>GND0, d_arr_merge2_8_31=>
      GND0, d_arr_merge2_8_30=>GND0, d_arr_merge2_8_29=>GND0, 
      d_arr_merge2_8_28=>GND0, d_arr_merge2_8_27=>GND0, d_arr_merge2_8_26=>
      GND0, d_arr_merge2_8_25=>GND0, d_arr_merge2_8_24=>GND0, 
      d_arr_merge2_8_23=>GND0, d_arr_merge2_8_22=>GND0, d_arr_merge2_8_21=>
      GND0, d_arr_merge2_8_20=>GND0, d_arr_merge2_8_19=>GND0, 
      d_arr_merge2_8_18=>GND0, d_arr_merge2_8_17=>GND0, d_arr_merge2_8_16=>
      GND0, d_arr_merge2_8_15=>GND0, d_arr_merge2_8_14=>GND0, 
      d_arr_merge2_8_13=>GND0, d_arr_merge2_8_12=>GND0, d_arr_merge2_8_11=>
      GND0, d_arr_merge2_8_10=>GND0, d_arr_merge2_8_9=>GND0, 
      d_arr_merge2_8_8=>GND0, d_arr_merge2_8_7=>GND0, d_arr_merge2_8_6=>GND0, 
      d_arr_merge2_8_5=>GND0, d_arr_merge2_8_4=>GND0, d_arr_merge2_8_3=>GND0, 
      d_arr_merge2_8_2=>GND0, d_arr_merge2_8_1=>GND0, d_arr_merge2_8_0=>GND0, 
      d_arr_merge2_9_31=>GND0, d_arr_merge2_9_30=>GND0, d_arr_merge2_9_29=>
      GND0, d_arr_merge2_9_28=>GND0, d_arr_merge2_9_27=>GND0, 
      d_arr_merge2_9_26=>GND0, d_arr_merge2_9_25=>GND0, d_arr_merge2_9_24=>
      GND0, d_arr_merge2_9_23=>GND0, d_arr_merge2_9_22=>GND0, 
      d_arr_merge2_9_21=>GND0, d_arr_merge2_9_20=>GND0, d_arr_merge2_9_19=>
      GND0, d_arr_merge2_9_18=>GND0, d_arr_merge2_9_17=>GND0, 
      d_arr_merge2_9_16=>GND0, d_arr_merge2_9_15=>GND0, d_arr_merge2_9_14=>
      GND0, d_arr_merge2_9_13=>GND0, d_arr_merge2_9_12=>GND0, 
      d_arr_merge2_9_11=>GND0, d_arr_merge2_9_10=>GND0, d_arr_merge2_9_9=>
      GND0, d_arr_merge2_9_8=>GND0, d_arr_merge2_9_7=>GND0, d_arr_merge2_9_6
      =>GND0, d_arr_merge2_9_5=>GND0, d_arr_merge2_9_4=>GND0, 
      d_arr_merge2_9_3=>GND0, d_arr_merge2_9_2=>GND0, d_arr_merge2_9_1=>GND0, 
      d_arr_merge2_9_0=>GND0, d_arr_merge2_10_31=>GND0, d_arr_merge2_10_30=>
      GND0, d_arr_merge2_10_29=>GND0, d_arr_merge2_10_28=>GND0, 
      d_arr_merge2_10_27=>GND0, d_arr_merge2_10_26=>GND0, d_arr_merge2_10_25
      =>GND0, d_arr_merge2_10_24=>GND0, d_arr_merge2_10_23=>GND0, 
      d_arr_merge2_10_22=>GND0, d_arr_merge2_10_21=>GND0, d_arr_merge2_10_20
      =>GND0, d_arr_merge2_10_19=>GND0, d_arr_merge2_10_18=>GND0, 
      d_arr_merge2_10_17=>GND0, d_arr_merge2_10_16=>GND0, d_arr_merge2_10_15
      =>GND0, d_arr_merge2_10_14=>GND0, d_arr_merge2_10_13=>GND0, 
      d_arr_merge2_10_12=>GND0, d_arr_merge2_10_11=>GND0, d_arr_merge2_10_10
      =>GND0, d_arr_merge2_10_9=>GND0, d_arr_merge2_10_8=>GND0, 
      d_arr_merge2_10_7=>GND0, d_arr_merge2_10_6=>GND0, d_arr_merge2_10_5=>
      GND0, d_arr_merge2_10_4=>GND0, d_arr_merge2_10_3=>GND0, 
      d_arr_merge2_10_2=>GND0, d_arr_merge2_10_1=>GND0, d_arr_merge2_10_0=>
      GND0, d_arr_merge2_11_31=>GND0, d_arr_merge2_11_30=>GND0, 
      d_arr_merge2_11_29=>GND0, d_arr_merge2_11_28=>GND0, d_arr_merge2_11_27
      =>GND0, d_arr_merge2_11_26=>GND0, d_arr_merge2_11_25=>GND0, 
      d_arr_merge2_11_24=>GND0, d_arr_merge2_11_23=>GND0, d_arr_merge2_11_22
      =>GND0, d_arr_merge2_11_21=>GND0, d_arr_merge2_11_20=>GND0, 
      d_arr_merge2_11_19=>GND0, d_arr_merge2_11_18=>GND0, d_arr_merge2_11_17
      =>GND0, d_arr_merge2_11_16=>GND0, d_arr_merge2_11_15=>GND0, 
      d_arr_merge2_11_14=>GND0, d_arr_merge2_11_13=>GND0, d_arr_merge2_11_12
      =>GND0, d_arr_merge2_11_11=>GND0, d_arr_merge2_11_10=>GND0, 
      d_arr_merge2_11_9=>GND0, d_arr_merge2_11_8=>GND0, d_arr_merge2_11_7=>
      GND0, d_arr_merge2_11_6=>GND0, d_arr_merge2_11_5=>GND0, 
      d_arr_merge2_11_4=>GND0, d_arr_merge2_11_3=>GND0, d_arr_merge2_11_2=>
      GND0, d_arr_merge2_11_1=>GND0, d_arr_merge2_11_0=>GND0, 
      d_arr_merge2_12_31=>GND0, d_arr_merge2_12_30=>GND0, d_arr_merge2_12_29
      =>GND0, d_arr_merge2_12_28=>GND0, d_arr_merge2_12_27=>GND0, 
      d_arr_merge2_12_26=>GND0, d_arr_merge2_12_25=>GND0, d_arr_merge2_12_24
      =>GND0, d_arr_merge2_12_23=>GND0, d_arr_merge2_12_22=>GND0, 
      d_arr_merge2_12_21=>GND0, d_arr_merge2_12_20=>GND0, d_arr_merge2_12_19
      =>GND0, d_arr_merge2_12_18=>GND0, d_arr_merge2_12_17=>GND0, 
      d_arr_merge2_12_16=>GND0, d_arr_merge2_12_15=>GND0, d_arr_merge2_12_14
      =>GND0, d_arr_merge2_12_13=>GND0, d_arr_merge2_12_12=>GND0, 
      d_arr_merge2_12_11=>GND0, d_arr_merge2_12_10=>GND0, d_arr_merge2_12_9
      =>GND0, d_arr_merge2_12_8=>GND0, d_arr_merge2_12_7=>GND0, 
      d_arr_merge2_12_6=>GND0, d_arr_merge2_12_5=>GND0, d_arr_merge2_12_4=>
      GND0, d_arr_merge2_12_3=>GND0, d_arr_merge2_12_2=>GND0, 
      d_arr_merge2_12_1=>GND0, d_arr_merge2_12_0=>GND0, d_arr_merge2_13_31=>
      GND0, d_arr_merge2_13_30=>GND0, d_arr_merge2_13_29=>GND0, 
      d_arr_merge2_13_28=>GND0, d_arr_merge2_13_27=>GND0, d_arr_merge2_13_26
      =>GND0, d_arr_merge2_13_25=>GND0, d_arr_merge2_13_24=>GND0, 
      d_arr_merge2_13_23=>GND0, d_arr_merge2_13_22=>GND0, d_arr_merge2_13_21
      =>GND0, d_arr_merge2_13_20=>GND0, d_arr_merge2_13_19=>GND0, 
      d_arr_merge2_13_18=>GND0, d_arr_merge2_13_17=>GND0, d_arr_merge2_13_16
      =>GND0, d_arr_merge2_13_15=>GND0, d_arr_merge2_13_14=>GND0, 
      d_arr_merge2_13_13=>GND0, d_arr_merge2_13_12=>GND0, d_arr_merge2_13_11
      =>GND0, d_arr_merge2_13_10=>GND0, d_arr_merge2_13_9=>GND0, 
      d_arr_merge2_13_8=>GND0, d_arr_merge2_13_7=>GND0, d_arr_merge2_13_6=>
      GND0, d_arr_merge2_13_5=>GND0, d_arr_merge2_13_4=>GND0, 
      d_arr_merge2_13_3=>GND0, d_arr_merge2_13_2=>GND0, d_arr_merge2_13_1=>
      GND0, d_arr_merge2_13_0=>GND0, d_arr_merge2_14_31=>GND0, 
      d_arr_merge2_14_30=>GND0, d_arr_merge2_14_29=>GND0, d_arr_merge2_14_28
      =>GND0, d_arr_merge2_14_27=>GND0, d_arr_merge2_14_26=>GND0, 
      d_arr_merge2_14_25=>GND0, d_arr_merge2_14_24=>GND0, d_arr_merge2_14_23
      =>GND0, d_arr_merge2_14_22=>GND0, d_arr_merge2_14_21=>GND0, 
      d_arr_merge2_14_20=>GND0, d_arr_merge2_14_19=>GND0, d_arr_merge2_14_18
      =>GND0, d_arr_merge2_14_17=>GND0, d_arr_merge2_14_16=>GND0, 
      d_arr_merge2_14_15=>GND0, d_arr_merge2_14_14=>GND0, d_arr_merge2_14_13
      =>GND0, d_arr_merge2_14_12=>GND0, d_arr_merge2_14_11=>GND0, 
      d_arr_merge2_14_10=>GND0, d_arr_merge2_14_9=>GND0, d_arr_merge2_14_8=>
      GND0, d_arr_merge2_14_7=>GND0, d_arr_merge2_14_6=>GND0, 
      d_arr_merge2_14_5=>GND0, d_arr_merge2_14_4=>GND0, d_arr_merge2_14_3=>
      GND0, d_arr_merge2_14_2=>GND0, d_arr_merge2_14_1=>GND0, 
      d_arr_merge2_14_0=>GND0, d_arr_merge2_15_31=>GND0, d_arr_merge2_15_30
      =>GND0, d_arr_merge2_15_29=>GND0, d_arr_merge2_15_28=>GND0, 
      d_arr_merge2_15_27=>GND0, d_arr_merge2_15_26=>GND0, d_arr_merge2_15_25
      =>GND0, d_arr_merge2_15_24=>GND0, d_arr_merge2_15_23=>GND0, 
      d_arr_merge2_15_22=>GND0, d_arr_merge2_15_21=>GND0, d_arr_merge2_15_20
      =>GND0, d_arr_merge2_15_19=>GND0, d_arr_merge2_15_18=>GND0, 
      d_arr_merge2_15_17=>GND0, d_arr_merge2_15_16=>GND0, d_arr_merge2_15_15
      =>GND0, d_arr_merge2_15_14=>GND0, d_arr_merge2_15_13=>GND0, 
      d_arr_merge2_15_12=>GND0, d_arr_merge2_15_11=>GND0, d_arr_merge2_15_10
      =>GND0, d_arr_merge2_15_9=>GND0, d_arr_merge2_15_8=>GND0, 
      d_arr_merge2_15_7=>GND0, d_arr_merge2_15_6=>GND0, d_arr_merge2_15_5=>
      GND0, d_arr_merge2_15_4=>GND0, d_arr_merge2_15_3=>GND0, 
      d_arr_merge2_15_2=>GND0, d_arr_merge2_15_1=>GND0, d_arr_merge2_15_0=>
      GND0, d_arr_merge2_16_31=>GND0, d_arr_merge2_16_30=>GND0, 
      d_arr_merge2_16_29=>GND0, d_arr_merge2_16_28=>GND0, d_arr_merge2_16_27
      =>GND0, d_arr_merge2_16_26=>GND0, d_arr_merge2_16_25=>GND0, 
      d_arr_merge2_16_24=>GND0, d_arr_merge2_16_23=>GND0, d_arr_merge2_16_22
      =>GND0, d_arr_merge2_16_21=>GND0, d_arr_merge2_16_20=>GND0, 
      d_arr_merge2_16_19=>GND0, d_arr_merge2_16_18=>GND0, d_arr_merge2_16_17
      =>GND0, d_arr_merge2_16_16=>GND0, d_arr_merge2_16_15=>GND0, 
      d_arr_merge2_16_14=>GND0, d_arr_merge2_16_13=>GND0, d_arr_merge2_16_12
      =>GND0, d_arr_merge2_16_11=>GND0, d_arr_merge2_16_10=>GND0, 
      d_arr_merge2_16_9=>GND0, d_arr_merge2_16_8=>GND0, d_arr_merge2_16_7=>
      GND0, d_arr_merge2_16_6=>GND0, d_arr_merge2_16_5=>GND0, 
      d_arr_merge2_16_4=>GND0, d_arr_merge2_16_3=>GND0, d_arr_merge2_16_2=>
      GND0, d_arr_merge2_16_1=>GND0, d_arr_merge2_16_0=>GND0, 
      d_arr_merge2_17_31=>GND0, d_arr_merge2_17_30=>GND0, d_arr_merge2_17_29
      =>GND0, d_arr_merge2_17_28=>GND0, d_arr_merge2_17_27=>GND0, 
      d_arr_merge2_17_26=>GND0, d_arr_merge2_17_25=>GND0, d_arr_merge2_17_24
      =>GND0, d_arr_merge2_17_23=>GND0, d_arr_merge2_17_22=>GND0, 
      d_arr_merge2_17_21=>GND0, d_arr_merge2_17_20=>GND0, d_arr_merge2_17_19
      =>GND0, d_arr_merge2_17_18=>GND0, d_arr_merge2_17_17=>GND0, 
      d_arr_merge2_17_16=>GND0, d_arr_merge2_17_15=>GND0, d_arr_merge2_17_14
      =>GND0, d_arr_merge2_17_13=>GND0, d_arr_merge2_17_12=>GND0, 
      d_arr_merge2_17_11=>GND0, d_arr_merge2_17_10=>GND0, d_arr_merge2_17_9
      =>GND0, d_arr_merge2_17_8=>GND0, d_arr_merge2_17_7=>GND0, 
      d_arr_merge2_17_6=>GND0, d_arr_merge2_17_5=>GND0, d_arr_merge2_17_4=>
      GND0, d_arr_merge2_17_3=>GND0, d_arr_merge2_17_2=>GND0, 
      d_arr_merge2_17_1=>GND0, d_arr_merge2_17_0=>GND0, d_arr_merge2_18_31=>
      GND0, d_arr_merge2_18_30=>GND0, d_arr_merge2_18_29=>GND0, 
      d_arr_merge2_18_28=>GND0, d_arr_merge2_18_27=>GND0, d_arr_merge2_18_26
      =>GND0, d_arr_merge2_18_25=>GND0, d_arr_merge2_18_24=>GND0, 
      d_arr_merge2_18_23=>GND0, d_arr_merge2_18_22=>GND0, d_arr_merge2_18_21
      =>GND0, d_arr_merge2_18_20=>GND0, d_arr_merge2_18_19=>GND0, 
      d_arr_merge2_18_18=>GND0, d_arr_merge2_18_17=>GND0, d_arr_merge2_18_16
      =>GND0, d_arr_merge2_18_15=>GND0, d_arr_merge2_18_14=>GND0, 
      d_arr_merge2_18_13=>GND0, d_arr_merge2_18_12=>GND0, d_arr_merge2_18_11
      =>GND0, d_arr_merge2_18_10=>GND0, d_arr_merge2_18_9=>GND0, 
      d_arr_merge2_18_8=>GND0, d_arr_merge2_18_7=>GND0, d_arr_merge2_18_6=>
      GND0, d_arr_merge2_18_5=>GND0, d_arr_merge2_18_4=>GND0, 
      d_arr_merge2_18_3=>GND0, d_arr_merge2_18_2=>GND0, d_arr_merge2_18_1=>
      GND0, d_arr_merge2_18_0=>GND0, d_arr_merge2_19_31=>GND0, 
      d_arr_merge2_19_30=>GND0, d_arr_merge2_19_29=>GND0, d_arr_merge2_19_28
      =>GND0, d_arr_merge2_19_27=>GND0, d_arr_merge2_19_26=>GND0, 
      d_arr_merge2_19_25=>GND0, d_arr_merge2_19_24=>GND0, d_arr_merge2_19_23
      =>GND0, d_arr_merge2_19_22=>GND0, d_arr_merge2_19_21=>GND0, 
      d_arr_merge2_19_20=>GND0, d_arr_merge2_19_19=>GND0, d_arr_merge2_19_18
      =>GND0, d_arr_merge2_19_17=>GND0, d_arr_merge2_19_16=>GND0, 
      d_arr_merge2_19_15=>GND0, d_arr_merge2_19_14=>GND0, d_arr_merge2_19_13
      =>GND0, d_arr_merge2_19_12=>GND0, d_arr_merge2_19_11=>GND0, 
      d_arr_merge2_19_10=>GND0, d_arr_merge2_19_9=>GND0, d_arr_merge2_19_8=>
      GND0, d_arr_merge2_19_7=>GND0, d_arr_merge2_19_6=>GND0, 
      d_arr_merge2_19_5=>GND0, d_arr_merge2_19_4=>GND0, d_arr_merge2_19_3=>
      GND0, d_arr_merge2_19_2=>GND0, d_arr_merge2_19_1=>GND0, 
      d_arr_merge2_19_0=>GND0, d_arr_merge2_20_31=>GND0, d_arr_merge2_20_30
      =>GND0, d_arr_merge2_20_29=>GND0, d_arr_merge2_20_28=>GND0, 
      d_arr_merge2_20_27=>GND0, d_arr_merge2_20_26=>GND0, d_arr_merge2_20_25
      =>GND0, d_arr_merge2_20_24=>GND0, d_arr_merge2_20_23=>GND0, 
      d_arr_merge2_20_22=>GND0, d_arr_merge2_20_21=>GND0, d_arr_merge2_20_20
      =>GND0, d_arr_merge2_20_19=>GND0, d_arr_merge2_20_18=>GND0, 
      d_arr_merge2_20_17=>GND0, d_arr_merge2_20_16=>GND0, d_arr_merge2_20_15
      =>GND0, d_arr_merge2_20_14=>GND0, d_arr_merge2_20_13=>GND0, 
      d_arr_merge2_20_12=>GND0, d_arr_merge2_20_11=>GND0, d_arr_merge2_20_10
      =>GND0, d_arr_merge2_20_9=>GND0, d_arr_merge2_20_8=>GND0, 
      d_arr_merge2_20_7=>GND0, d_arr_merge2_20_6=>GND0, d_arr_merge2_20_5=>
      GND0, d_arr_merge2_20_4=>GND0, d_arr_merge2_20_3=>GND0, 
      d_arr_merge2_20_2=>GND0, d_arr_merge2_20_1=>GND0, d_arr_merge2_20_0=>
      GND0, d_arr_merge2_21_31=>GND0, d_arr_merge2_21_30=>GND0, 
      d_arr_merge2_21_29=>GND0, d_arr_merge2_21_28=>GND0, d_arr_merge2_21_27
      =>GND0, d_arr_merge2_21_26=>GND0, d_arr_merge2_21_25=>GND0, 
      d_arr_merge2_21_24=>GND0, d_arr_merge2_21_23=>GND0, d_arr_merge2_21_22
      =>GND0, d_arr_merge2_21_21=>GND0, d_arr_merge2_21_20=>GND0, 
      d_arr_merge2_21_19=>GND0, d_arr_merge2_21_18=>GND0, d_arr_merge2_21_17
      =>GND0, d_arr_merge2_21_16=>GND0, d_arr_merge2_21_15=>GND0, 
      d_arr_merge2_21_14=>GND0, d_arr_merge2_21_13=>GND0, d_arr_merge2_21_12
      =>GND0, d_arr_merge2_21_11=>GND0, d_arr_merge2_21_10=>GND0, 
      d_arr_merge2_21_9=>GND0, d_arr_merge2_21_8=>GND0, d_arr_merge2_21_7=>
      GND0, d_arr_merge2_21_6=>GND0, d_arr_merge2_21_5=>GND0, 
      d_arr_merge2_21_4=>GND0, d_arr_merge2_21_3=>GND0, d_arr_merge2_21_2=>
      GND0, d_arr_merge2_21_1=>GND0, d_arr_merge2_21_0=>GND0, 
      d_arr_merge2_22_31=>GND0, d_arr_merge2_22_30=>GND0, d_arr_merge2_22_29
      =>GND0, d_arr_merge2_22_28=>GND0, d_arr_merge2_22_27=>GND0, 
      d_arr_merge2_22_26=>GND0, d_arr_merge2_22_25=>GND0, d_arr_merge2_22_24
      =>GND0, d_arr_merge2_22_23=>GND0, d_arr_merge2_22_22=>GND0, 
      d_arr_merge2_22_21=>GND0, d_arr_merge2_22_20=>GND0, d_arr_merge2_22_19
      =>GND0, d_arr_merge2_22_18=>GND0, d_arr_merge2_22_17=>GND0, 
      d_arr_merge2_22_16=>GND0, d_arr_merge2_22_15=>GND0, d_arr_merge2_22_14
      =>GND0, d_arr_merge2_22_13=>GND0, d_arr_merge2_22_12=>GND0, 
      d_arr_merge2_22_11=>GND0, d_arr_merge2_22_10=>GND0, d_arr_merge2_22_9
      =>GND0, d_arr_merge2_22_8=>GND0, d_arr_merge2_22_7=>GND0, 
      d_arr_merge2_22_6=>GND0, d_arr_merge2_22_5=>GND0, d_arr_merge2_22_4=>
      GND0, d_arr_merge2_22_3=>GND0, d_arr_merge2_22_2=>GND0, 
      d_arr_merge2_22_1=>GND0, d_arr_merge2_22_0=>GND0, d_arr_merge2_23_31=>
      GND0, d_arr_merge2_23_30=>GND0, d_arr_merge2_23_29=>GND0, 
      d_arr_merge2_23_28=>GND0, d_arr_merge2_23_27=>GND0, d_arr_merge2_23_26
      =>GND0, d_arr_merge2_23_25=>GND0, d_arr_merge2_23_24=>GND0, 
      d_arr_merge2_23_23=>GND0, d_arr_merge2_23_22=>GND0, d_arr_merge2_23_21
      =>GND0, d_arr_merge2_23_20=>GND0, d_arr_merge2_23_19=>GND0, 
      d_arr_merge2_23_18=>GND0, d_arr_merge2_23_17=>GND0, d_arr_merge2_23_16
      =>GND0, d_arr_merge2_23_15=>GND0, d_arr_merge2_23_14=>GND0, 
      d_arr_merge2_23_13=>GND0, d_arr_merge2_23_12=>GND0, d_arr_merge2_23_11
      =>GND0, d_arr_merge2_23_10=>GND0, d_arr_merge2_23_9=>GND0, 
      d_arr_merge2_23_8=>GND0, d_arr_merge2_23_7=>GND0, d_arr_merge2_23_6=>
      GND0, d_arr_merge2_23_5=>GND0, d_arr_merge2_23_4=>GND0, 
      d_arr_merge2_23_3=>GND0, d_arr_merge2_23_2=>GND0, d_arr_merge2_23_1=>
      GND0, d_arr_merge2_23_0=>GND0, d_arr_merge2_24_31=>GND0, 
      d_arr_merge2_24_30=>GND0, d_arr_merge2_24_29=>GND0, d_arr_merge2_24_28
      =>GND0, d_arr_merge2_24_27=>GND0, d_arr_merge2_24_26=>GND0, 
      d_arr_merge2_24_25=>GND0, d_arr_merge2_24_24=>GND0, d_arr_merge2_24_23
      =>GND0, d_arr_merge2_24_22=>GND0, d_arr_merge2_24_21=>GND0, 
      d_arr_merge2_24_20=>GND0, d_arr_merge2_24_19=>GND0, d_arr_merge2_24_18
      =>GND0, d_arr_merge2_24_17=>GND0, d_arr_merge2_24_16=>GND0, 
      d_arr_merge2_24_15=>GND0, d_arr_merge2_24_14=>GND0, d_arr_merge2_24_13
      =>GND0, d_arr_merge2_24_12=>GND0, d_arr_merge2_24_11=>GND0, 
      d_arr_merge2_24_10=>GND0, d_arr_merge2_24_9=>GND0, d_arr_merge2_24_8=>
      GND0, d_arr_merge2_24_7=>GND0, d_arr_merge2_24_6=>GND0, 
      d_arr_merge2_24_5=>GND0, d_arr_merge2_24_4=>GND0, d_arr_merge2_24_3=>
      GND0, d_arr_merge2_24_2=>GND0, d_arr_merge2_24_1=>GND0, 
      d_arr_merge2_24_0=>GND0, d_arr_relu_0_31=>d_arr_relu_0_31, 
      d_arr_relu_0_30=>d_arr_relu_0_30, d_arr_relu_0_29=>d_arr_relu_0_29, 
      d_arr_relu_0_28=>d_arr_relu_0_28, d_arr_relu_0_27=>d_arr_relu_0_27, 
      d_arr_relu_0_26=>d_arr_relu_0_26, d_arr_relu_0_25=>d_arr_relu_0_25, 
      d_arr_relu_0_24=>d_arr_relu_0_24, d_arr_relu_0_23=>d_arr_relu_0_23, 
      d_arr_relu_0_22=>d_arr_relu_0_22, d_arr_relu_0_21=>d_arr_relu_0_21, 
      d_arr_relu_0_20=>d_arr_relu_0_20, d_arr_relu_0_19=>d_arr_relu_0_19, 
      d_arr_relu_0_18=>d_arr_relu_0_18, d_arr_relu_0_17=>d_arr_relu_0_17, 
      d_arr_relu_0_16=>d_arr_relu_0_16, d_arr_relu_0_15=>GND0, 
      d_arr_relu_0_14=>d_arr_relu_0_14, d_arr_relu_0_13=>d_arr_relu_0_13, 
      d_arr_relu_0_12=>d_arr_relu_0_12, d_arr_relu_0_11=>d_arr_relu_0_11, 
      d_arr_relu_0_10=>d_arr_relu_0_10, d_arr_relu_0_9=>d_arr_relu_0_9, 
      d_arr_relu_0_8=>d_arr_relu_0_8, d_arr_relu_0_7=>d_arr_relu_0_7, 
      d_arr_relu_0_6=>d_arr_relu_0_6, d_arr_relu_0_5=>d_arr_relu_0_5, 
      d_arr_relu_0_4=>d_arr_relu_0_4, d_arr_relu_0_3=>d_arr_relu_0_3, 
      d_arr_relu_0_2=>d_arr_relu_0_2, d_arr_relu_0_1=>d_arr_relu_0_1, 
      d_arr_relu_0_0=>d_arr_relu_0_0, d_arr_relu_1_31=>d_arr_relu_1_31, 
      d_arr_relu_1_30=>d_arr_relu_1_30, d_arr_relu_1_29=>d_arr_relu_1_29, 
      d_arr_relu_1_28=>d_arr_relu_1_28, d_arr_relu_1_27=>d_arr_relu_1_27, 
      d_arr_relu_1_26=>d_arr_relu_1_26, d_arr_relu_1_25=>d_arr_relu_1_25, 
      d_arr_relu_1_24=>d_arr_relu_1_24, d_arr_relu_1_23=>d_arr_relu_1_23, 
      d_arr_relu_1_22=>d_arr_relu_1_22, d_arr_relu_1_21=>d_arr_relu_1_21, 
      d_arr_relu_1_20=>d_arr_relu_1_20, d_arr_relu_1_19=>d_arr_relu_1_19, 
      d_arr_relu_1_18=>d_arr_relu_1_18, d_arr_relu_1_17=>d_arr_relu_1_17, 
      d_arr_relu_1_16=>d_arr_relu_1_16, d_arr_relu_1_15=>GND0, 
      d_arr_relu_1_14=>d_arr_relu_1_14, d_arr_relu_1_13=>d_arr_relu_1_13, 
      d_arr_relu_1_12=>d_arr_relu_1_12, d_arr_relu_1_11=>d_arr_relu_1_11, 
      d_arr_relu_1_10=>d_arr_relu_1_10, d_arr_relu_1_9=>d_arr_relu_1_9, 
      d_arr_relu_1_8=>d_arr_relu_1_8, d_arr_relu_1_7=>d_arr_relu_1_7, 
      d_arr_relu_1_6=>d_arr_relu_1_6, d_arr_relu_1_5=>d_arr_relu_1_5, 
      d_arr_relu_1_4=>d_arr_relu_1_4, d_arr_relu_1_3=>d_arr_relu_1_3, 
      d_arr_relu_1_2=>d_arr_relu_1_2, d_arr_relu_1_1=>d_arr_relu_1_1, 
      d_arr_relu_1_0=>d_arr_relu_1_0, d_arr_relu_2_31=>GND0, d_arr_relu_2_30
      =>GND0, d_arr_relu_2_29=>GND0, d_arr_relu_2_28=>GND0, d_arr_relu_2_27
      =>GND0, d_arr_relu_2_26=>GND0, d_arr_relu_2_25=>GND0, d_arr_relu_2_24
      =>GND0, d_arr_relu_2_23=>GND0, d_arr_relu_2_22=>GND0, d_arr_relu_2_21
      =>GND0, d_arr_relu_2_20=>GND0, d_arr_relu_2_19=>GND0, d_arr_relu_2_18
      =>GND0, d_arr_relu_2_17=>GND0, d_arr_relu_2_16=>GND0, d_arr_relu_2_15
      =>GND0, d_arr_relu_2_14=>GND0, d_arr_relu_2_13=>GND0, d_arr_relu_2_12
      =>GND0, d_arr_relu_2_11=>GND0, d_arr_relu_2_10=>GND0, d_arr_relu_2_9=>
      GND0, d_arr_relu_2_8=>GND0, d_arr_relu_2_7=>GND0, d_arr_relu_2_6=>GND0, 
      d_arr_relu_2_5=>GND0, d_arr_relu_2_4=>GND0, d_arr_relu_2_3=>GND0, 
      d_arr_relu_2_2=>GND0, d_arr_relu_2_1=>GND0, d_arr_relu_2_0=>GND0, 
      d_arr_relu_3_31=>GND0, d_arr_relu_3_30=>GND0, d_arr_relu_3_29=>GND0, 
      d_arr_relu_3_28=>GND0, d_arr_relu_3_27=>GND0, d_arr_relu_3_26=>GND0, 
      d_arr_relu_3_25=>GND0, d_arr_relu_3_24=>GND0, d_arr_relu_3_23=>GND0, 
      d_arr_relu_3_22=>GND0, d_arr_relu_3_21=>GND0, d_arr_relu_3_20=>GND0, 
      d_arr_relu_3_19=>GND0, d_arr_relu_3_18=>GND0, d_arr_relu_3_17=>GND0, 
      d_arr_relu_3_16=>GND0, d_arr_relu_3_15=>GND0, d_arr_relu_3_14=>GND0, 
      d_arr_relu_3_13=>GND0, d_arr_relu_3_12=>GND0, d_arr_relu_3_11=>GND0, 
      d_arr_relu_3_10=>GND0, d_arr_relu_3_9=>GND0, d_arr_relu_3_8=>GND0, 
      d_arr_relu_3_7=>GND0, d_arr_relu_3_6=>GND0, d_arr_relu_3_5=>GND0, 
      d_arr_relu_3_4=>GND0, d_arr_relu_3_3=>GND0, d_arr_relu_3_2=>GND0, 
      d_arr_relu_3_1=>GND0, d_arr_relu_3_0=>GND0, d_arr_relu_4_31=>GND0, 
      d_arr_relu_4_30=>GND0, d_arr_relu_4_29=>GND0, d_arr_relu_4_28=>GND0, 
      d_arr_relu_4_27=>GND0, d_arr_relu_4_26=>GND0, d_arr_relu_4_25=>GND0, 
      d_arr_relu_4_24=>GND0, d_arr_relu_4_23=>GND0, d_arr_relu_4_22=>GND0, 
      d_arr_relu_4_21=>GND0, d_arr_relu_4_20=>GND0, d_arr_relu_4_19=>GND0, 
      d_arr_relu_4_18=>GND0, d_arr_relu_4_17=>GND0, d_arr_relu_4_16=>GND0, 
      d_arr_relu_4_15=>GND0, d_arr_relu_4_14=>GND0, d_arr_relu_4_13=>GND0, 
      d_arr_relu_4_12=>GND0, d_arr_relu_4_11=>GND0, d_arr_relu_4_10=>GND0, 
      d_arr_relu_4_9=>GND0, d_arr_relu_4_8=>GND0, d_arr_relu_4_7=>GND0, 
      d_arr_relu_4_6=>GND0, d_arr_relu_4_5=>GND0, d_arr_relu_4_4=>GND0, 
      d_arr_relu_4_3=>GND0, d_arr_relu_4_2=>GND0, d_arr_relu_4_1=>GND0, 
      d_arr_relu_4_0=>GND0, d_arr_relu_5_31=>GND0, d_arr_relu_5_30=>GND0, 
      d_arr_relu_5_29=>GND0, d_arr_relu_5_28=>GND0, d_arr_relu_5_27=>GND0, 
      d_arr_relu_5_26=>GND0, d_arr_relu_5_25=>GND0, d_arr_relu_5_24=>GND0, 
      d_arr_relu_5_23=>GND0, d_arr_relu_5_22=>GND0, d_arr_relu_5_21=>GND0, 
      d_arr_relu_5_20=>GND0, d_arr_relu_5_19=>GND0, d_arr_relu_5_18=>GND0, 
      d_arr_relu_5_17=>GND0, d_arr_relu_5_16=>GND0, d_arr_relu_5_15=>GND0, 
      d_arr_relu_5_14=>GND0, d_arr_relu_5_13=>GND0, d_arr_relu_5_12=>GND0, 
      d_arr_relu_5_11=>GND0, d_arr_relu_5_10=>GND0, d_arr_relu_5_9=>GND0, 
      d_arr_relu_5_8=>GND0, d_arr_relu_5_7=>GND0, d_arr_relu_5_6=>GND0, 
      d_arr_relu_5_5=>GND0, d_arr_relu_5_4=>GND0, d_arr_relu_5_3=>GND0, 
      d_arr_relu_5_2=>GND0, d_arr_relu_5_1=>GND0, d_arr_relu_5_0=>GND0, 
      d_arr_relu_6_31=>GND0, d_arr_relu_6_30=>GND0, d_arr_relu_6_29=>GND0, 
      d_arr_relu_6_28=>GND0, d_arr_relu_6_27=>GND0, d_arr_relu_6_26=>GND0, 
      d_arr_relu_6_25=>GND0, d_arr_relu_6_24=>GND0, d_arr_relu_6_23=>GND0, 
      d_arr_relu_6_22=>GND0, d_arr_relu_6_21=>GND0, d_arr_relu_6_20=>GND0, 
      d_arr_relu_6_19=>GND0, d_arr_relu_6_18=>GND0, d_arr_relu_6_17=>GND0, 
      d_arr_relu_6_16=>GND0, d_arr_relu_6_15=>GND0, d_arr_relu_6_14=>GND0, 
      d_arr_relu_6_13=>GND0, d_arr_relu_6_12=>GND0, d_arr_relu_6_11=>GND0, 
      d_arr_relu_6_10=>GND0, d_arr_relu_6_9=>GND0, d_arr_relu_6_8=>GND0, 
      d_arr_relu_6_7=>GND0, d_arr_relu_6_6=>GND0, d_arr_relu_6_5=>GND0, 
      d_arr_relu_6_4=>GND0, d_arr_relu_6_3=>GND0, d_arr_relu_6_2=>GND0, 
      d_arr_relu_6_1=>GND0, d_arr_relu_6_0=>GND0, d_arr_relu_7_31=>GND0, 
      d_arr_relu_7_30=>GND0, d_arr_relu_7_29=>GND0, d_arr_relu_7_28=>GND0, 
      d_arr_relu_7_27=>GND0, d_arr_relu_7_26=>GND0, d_arr_relu_7_25=>GND0, 
      d_arr_relu_7_24=>GND0, d_arr_relu_7_23=>GND0, d_arr_relu_7_22=>GND0, 
      d_arr_relu_7_21=>GND0, d_arr_relu_7_20=>GND0, d_arr_relu_7_19=>GND0, 
      d_arr_relu_7_18=>GND0, d_arr_relu_7_17=>GND0, d_arr_relu_7_16=>GND0, 
      d_arr_relu_7_15=>GND0, d_arr_relu_7_14=>GND0, d_arr_relu_7_13=>GND0, 
      d_arr_relu_7_12=>GND0, d_arr_relu_7_11=>GND0, d_arr_relu_7_10=>GND0, 
      d_arr_relu_7_9=>GND0, d_arr_relu_7_8=>GND0, d_arr_relu_7_7=>GND0, 
      d_arr_relu_7_6=>GND0, d_arr_relu_7_5=>GND0, d_arr_relu_7_4=>GND0, 
      d_arr_relu_7_3=>GND0, d_arr_relu_7_2=>GND0, d_arr_relu_7_1=>GND0, 
      d_arr_relu_7_0=>GND0, d_arr_relu_8_31=>GND0, d_arr_relu_8_30=>GND0, 
      d_arr_relu_8_29=>GND0, d_arr_relu_8_28=>GND0, d_arr_relu_8_27=>GND0, 
      d_arr_relu_8_26=>GND0, d_arr_relu_8_25=>GND0, d_arr_relu_8_24=>GND0, 
      d_arr_relu_8_23=>GND0, d_arr_relu_8_22=>GND0, d_arr_relu_8_21=>GND0, 
      d_arr_relu_8_20=>GND0, d_arr_relu_8_19=>GND0, d_arr_relu_8_18=>GND0, 
      d_arr_relu_8_17=>GND0, d_arr_relu_8_16=>GND0, d_arr_relu_8_15=>GND0, 
      d_arr_relu_8_14=>GND0, d_arr_relu_8_13=>GND0, d_arr_relu_8_12=>GND0, 
      d_arr_relu_8_11=>GND0, d_arr_relu_8_10=>GND0, d_arr_relu_8_9=>GND0, 
      d_arr_relu_8_8=>GND0, d_arr_relu_8_7=>GND0, d_arr_relu_8_6=>GND0, 
      d_arr_relu_8_5=>GND0, d_arr_relu_8_4=>GND0, d_arr_relu_8_3=>GND0, 
      d_arr_relu_8_2=>GND0, d_arr_relu_8_1=>GND0, d_arr_relu_8_0=>GND0, 
      d_arr_relu_9_31=>GND0, d_arr_relu_9_30=>GND0, d_arr_relu_9_29=>GND0, 
      d_arr_relu_9_28=>GND0, d_arr_relu_9_27=>GND0, d_arr_relu_9_26=>GND0, 
      d_arr_relu_9_25=>GND0, d_arr_relu_9_24=>GND0, d_arr_relu_9_23=>GND0, 
      d_arr_relu_9_22=>GND0, d_arr_relu_9_21=>GND0, d_arr_relu_9_20=>GND0, 
      d_arr_relu_9_19=>GND0, d_arr_relu_9_18=>GND0, d_arr_relu_9_17=>GND0, 
      d_arr_relu_9_16=>GND0, d_arr_relu_9_15=>GND0, d_arr_relu_9_14=>GND0, 
      d_arr_relu_9_13=>GND0, d_arr_relu_9_12=>GND0, d_arr_relu_9_11=>GND0, 
      d_arr_relu_9_10=>GND0, d_arr_relu_9_9=>GND0, d_arr_relu_9_8=>GND0, 
      d_arr_relu_9_7=>GND0, d_arr_relu_9_6=>GND0, d_arr_relu_9_5=>GND0, 
      d_arr_relu_9_4=>GND0, d_arr_relu_9_3=>GND0, d_arr_relu_9_2=>GND0, 
      d_arr_relu_9_1=>GND0, d_arr_relu_9_0=>GND0, d_arr_relu_10_31=>GND0, 
      d_arr_relu_10_30=>GND0, d_arr_relu_10_29=>GND0, d_arr_relu_10_28=>GND0, 
      d_arr_relu_10_27=>GND0, d_arr_relu_10_26=>GND0, d_arr_relu_10_25=>GND0, 
      d_arr_relu_10_24=>GND0, d_arr_relu_10_23=>GND0, d_arr_relu_10_22=>GND0, 
      d_arr_relu_10_21=>GND0, d_arr_relu_10_20=>GND0, d_arr_relu_10_19=>GND0, 
      d_arr_relu_10_18=>GND0, d_arr_relu_10_17=>GND0, d_arr_relu_10_16=>GND0, 
      d_arr_relu_10_15=>GND0, d_arr_relu_10_14=>GND0, d_arr_relu_10_13=>GND0, 
      d_arr_relu_10_12=>GND0, d_arr_relu_10_11=>GND0, d_arr_relu_10_10=>GND0, 
      d_arr_relu_10_9=>GND0, d_arr_relu_10_8=>GND0, d_arr_relu_10_7=>GND0, 
      d_arr_relu_10_6=>GND0, d_arr_relu_10_5=>GND0, d_arr_relu_10_4=>GND0, 
      d_arr_relu_10_3=>GND0, d_arr_relu_10_2=>GND0, d_arr_relu_10_1=>GND0, 
      d_arr_relu_10_0=>GND0, d_arr_relu_11_31=>GND0, d_arr_relu_11_30=>GND0, 
      d_arr_relu_11_29=>GND0, d_arr_relu_11_28=>GND0, d_arr_relu_11_27=>GND0, 
      d_arr_relu_11_26=>GND0, d_arr_relu_11_25=>GND0, d_arr_relu_11_24=>GND0, 
      d_arr_relu_11_23=>GND0, d_arr_relu_11_22=>GND0, d_arr_relu_11_21=>GND0, 
      d_arr_relu_11_20=>GND0, d_arr_relu_11_19=>GND0, d_arr_relu_11_18=>GND0, 
      d_arr_relu_11_17=>GND0, d_arr_relu_11_16=>GND0, d_arr_relu_11_15=>GND0, 
      d_arr_relu_11_14=>GND0, d_arr_relu_11_13=>GND0, d_arr_relu_11_12=>GND0, 
      d_arr_relu_11_11=>GND0, d_arr_relu_11_10=>GND0, d_arr_relu_11_9=>GND0, 
      d_arr_relu_11_8=>GND0, d_arr_relu_11_7=>GND0, d_arr_relu_11_6=>GND0, 
      d_arr_relu_11_5=>GND0, d_arr_relu_11_4=>GND0, d_arr_relu_11_3=>GND0, 
      d_arr_relu_11_2=>GND0, d_arr_relu_11_1=>GND0, d_arr_relu_11_0=>GND0, 
      d_arr_relu_12_31=>GND0, d_arr_relu_12_30=>GND0, d_arr_relu_12_29=>GND0, 
      d_arr_relu_12_28=>GND0, d_arr_relu_12_27=>GND0, d_arr_relu_12_26=>GND0, 
      d_arr_relu_12_25=>GND0, d_arr_relu_12_24=>GND0, d_arr_relu_12_23=>GND0, 
      d_arr_relu_12_22=>GND0, d_arr_relu_12_21=>GND0, d_arr_relu_12_20=>GND0, 
      d_arr_relu_12_19=>GND0, d_arr_relu_12_18=>GND0, d_arr_relu_12_17=>GND0, 
      d_arr_relu_12_16=>GND0, d_arr_relu_12_15=>GND0, d_arr_relu_12_14=>GND0, 
      d_arr_relu_12_13=>GND0, d_arr_relu_12_12=>GND0, d_arr_relu_12_11=>GND0, 
      d_arr_relu_12_10=>GND0, d_arr_relu_12_9=>GND0, d_arr_relu_12_8=>GND0, 
      d_arr_relu_12_7=>GND0, d_arr_relu_12_6=>GND0, d_arr_relu_12_5=>GND0, 
      d_arr_relu_12_4=>GND0, d_arr_relu_12_3=>GND0, d_arr_relu_12_2=>GND0, 
      d_arr_relu_12_1=>GND0, d_arr_relu_12_0=>GND0, d_arr_relu_13_31=>GND0, 
      d_arr_relu_13_30=>GND0, d_arr_relu_13_29=>GND0, d_arr_relu_13_28=>GND0, 
      d_arr_relu_13_27=>GND0, d_arr_relu_13_26=>GND0, d_arr_relu_13_25=>GND0, 
      d_arr_relu_13_24=>GND0, d_arr_relu_13_23=>GND0, d_arr_relu_13_22=>GND0, 
      d_arr_relu_13_21=>GND0, d_arr_relu_13_20=>GND0, d_arr_relu_13_19=>GND0, 
      d_arr_relu_13_18=>GND0, d_arr_relu_13_17=>GND0, d_arr_relu_13_16=>GND0, 
      d_arr_relu_13_15=>GND0, d_arr_relu_13_14=>GND0, d_arr_relu_13_13=>GND0, 
      d_arr_relu_13_12=>GND0, d_arr_relu_13_11=>GND0, d_arr_relu_13_10=>GND0, 
      d_arr_relu_13_9=>GND0, d_arr_relu_13_8=>GND0, d_arr_relu_13_7=>GND0, 
      d_arr_relu_13_6=>GND0, d_arr_relu_13_5=>GND0, d_arr_relu_13_4=>GND0, 
      d_arr_relu_13_3=>GND0, d_arr_relu_13_2=>GND0, d_arr_relu_13_1=>GND0, 
      d_arr_relu_13_0=>GND0, d_arr_relu_14_31=>GND0, d_arr_relu_14_30=>GND0, 
      d_arr_relu_14_29=>GND0, d_arr_relu_14_28=>GND0, d_arr_relu_14_27=>GND0, 
      d_arr_relu_14_26=>GND0, d_arr_relu_14_25=>GND0, d_arr_relu_14_24=>GND0, 
      d_arr_relu_14_23=>GND0, d_arr_relu_14_22=>GND0, d_arr_relu_14_21=>GND0, 
      d_arr_relu_14_20=>GND0, d_arr_relu_14_19=>GND0, d_arr_relu_14_18=>GND0, 
      d_arr_relu_14_17=>GND0, d_arr_relu_14_16=>GND0, d_arr_relu_14_15=>GND0, 
      d_arr_relu_14_14=>GND0, d_arr_relu_14_13=>GND0, d_arr_relu_14_12=>GND0, 
      d_arr_relu_14_11=>GND0, d_arr_relu_14_10=>GND0, d_arr_relu_14_9=>GND0, 
      d_arr_relu_14_8=>GND0, d_arr_relu_14_7=>GND0, d_arr_relu_14_6=>GND0, 
      d_arr_relu_14_5=>GND0, d_arr_relu_14_4=>GND0, d_arr_relu_14_3=>GND0, 
      d_arr_relu_14_2=>GND0, d_arr_relu_14_1=>GND0, d_arr_relu_14_0=>GND0, 
      d_arr_relu_15_31=>GND0, d_arr_relu_15_30=>GND0, d_arr_relu_15_29=>GND0, 
      d_arr_relu_15_28=>GND0, d_arr_relu_15_27=>GND0, d_arr_relu_15_26=>GND0, 
      d_arr_relu_15_25=>GND0, d_arr_relu_15_24=>GND0, d_arr_relu_15_23=>GND0, 
      d_arr_relu_15_22=>GND0, d_arr_relu_15_21=>GND0, d_arr_relu_15_20=>GND0, 
      d_arr_relu_15_19=>GND0, d_arr_relu_15_18=>GND0, d_arr_relu_15_17=>GND0, 
      d_arr_relu_15_16=>GND0, d_arr_relu_15_15=>GND0, d_arr_relu_15_14=>GND0, 
      d_arr_relu_15_13=>GND0, d_arr_relu_15_12=>GND0, d_arr_relu_15_11=>GND0, 
      d_arr_relu_15_10=>GND0, d_arr_relu_15_9=>GND0, d_arr_relu_15_8=>GND0, 
      d_arr_relu_15_7=>GND0, d_arr_relu_15_6=>GND0, d_arr_relu_15_5=>GND0, 
      d_arr_relu_15_4=>GND0, d_arr_relu_15_3=>GND0, d_arr_relu_15_2=>GND0, 
      d_arr_relu_15_1=>GND0, d_arr_relu_15_0=>GND0, d_arr_relu_16_31=>GND0, 
      d_arr_relu_16_30=>GND0, d_arr_relu_16_29=>GND0, d_arr_relu_16_28=>GND0, 
      d_arr_relu_16_27=>GND0, d_arr_relu_16_26=>GND0, d_arr_relu_16_25=>GND0, 
      d_arr_relu_16_24=>GND0, d_arr_relu_16_23=>GND0, d_arr_relu_16_22=>GND0, 
      d_arr_relu_16_21=>GND0, d_arr_relu_16_20=>GND0, d_arr_relu_16_19=>GND0, 
      d_arr_relu_16_18=>GND0, d_arr_relu_16_17=>GND0, d_arr_relu_16_16=>GND0, 
      d_arr_relu_16_15=>GND0, d_arr_relu_16_14=>GND0, d_arr_relu_16_13=>GND0, 
      d_arr_relu_16_12=>GND0, d_arr_relu_16_11=>GND0, d_arr_relu_16_10=>GND0, 
      d_arr_relu_16_9=>GND0, d_arr_relu_16_8=>GND0, d_arr_relu_16_7=>GND0, 
      d_arr_relu_16_6=>GND0, d_arr_relu_16_5=>GND0, d_arr_relu_16_4=>GND0, 
      d_arr_relu_16_3=>GND0, d_arr_relu_16_2=>GND0, d_arr_relu_16_1=>GND0, 
      d_arr_relu_16_0=>GND0, d_arr_relu_17_31=>GND0, d_arr_relu_17_30=>GND0, 
      d_arr_relu_17_29=>GND0, d_arr_relu_17_28=>GND0, d_arr_relu_17_27=>GND0, 
      d_arr_relu_17_26=>GND0, d_arr_relu_17_25=>GND0, d_arr_relu_17_24=>GND0, 
      d_arr_relu_17_23=>GND0, d_arr_relu_17_22=>GND0, d_arr_relu_17_21=>GND0, 
      d_arr_relu_17_20=>GND0, d_arr_relu_17_19=>GND0, d_arr_relu_17_18=>GND0, 
      d_arr_relu_17_17=>GND0, d_arr_relu_17_16=>GND0, d_arr_relu_17_15=>GND0, 
      d_arr_relu_17_14=>GND0, d_arr_relu_17_13=>GND0, d_arr_relu_17_12=>GND0, 
      d_arr_relu_17_11=>GND0, d_arr_relu_17_10=>GND0, d_arr_relu_17_9=>GND0, 
      d_arr_relu_17_8=>GND0, d_arr_relu_17_7=>GND0, d_arr_relu_17_6=>GND0, 
      d_arr_relu_17_5=>GND0, d_arr_relu_17_4=>GND0, d_arr_relu_17_3=>GND0, 
      d_arr_relu_17_2=>GND0, d_arr_relu_17_1=>GND0, d_arr_relu_17_0=>GND0, 
      d_arr_relu_18_31=>GND0, d_arr_relu_18_30=>GND0, d_arr_relu_18_29=>GND0, 
      d_arr_relu_18_28=>GND0, d_arr_relu_18_27=>GND0, d_arr_relu_18_26=>GND0, 
      d_arr_relu_18_25=>GND0, d_arr_relu_18_24=>GND0, d_arr_relu_18_23=>GND0, 
      d_arr_relu_18_22=>GND0, d_arr_relu_18_21=>GND0, d_arr_relu_18_20=>GND0, 
      d_arr_relu_18_19=>GND0, d_arr_relu_18_18=>GND0, d_arr_relu_18_17=>GND0, 
      d_arr_relu_18_16=>GND0, d_arr_relu_18_15=>GND0, d_arr_relu_18_14=>GND0, 
      d_arr_relu_18_13=>GND0, d_arr_relu_18_12=>GND0, d_arr_relu_18_11=>GND0, 
      d_arr_relu_18_10=>GND0, d_arr_relu_18_9=>GND0, d_arr_relu_18_8=>GND0, 
      d_arr_relu_18_7=>GND0, d_arr_relu_18_6=>GND0, d_arr_relu_18_5=>GND0, 
      d_arr_relu_18_4=>GND0, d_arr_relu_18_3=>GND0, d_arr_relu_18_2=>GND0, 
      d_arr_relu_18_1=>GND0, d_arr_relu_18_0=>GND0, d_arr_relu_19_31=>GND0, 
      d_arr_relu_19_30=>GND0, d_arr_relu_19_29=>GND0, d_arr_relu_19_28=>GND0, 
      d_arr_relu_19_27=>GND0, d_arr_relu_19_26=>GND0, d_arr_relu_19_25=>GND0, 
      d_arr_relu_19_24=>GND0, d_arr_relu_19_23=>GND0, d_arr_relu_19_22=>GND0, 
      d_arr_relu_19_21=>GND0, d_arr_relu_19_20=>GND0, d_arr_relu_19_19=>GND0, 
      d_arr_relu_19_18=>GND0, d_arr_relu_19_17=>GND0, d_arr_relu_19_16=>GND0, 
      d_arr_relu_19_15=>GND0, d_arr_relu_19_14=>GND0, d_arr_relu_19_13=>GND0, 
      d_arr_relu_19_12=>GND0, d_arr_relu_19_11=>GND0, d_arr_relu_19_10=>GND0, 
      d_arr_relu_19_9=>GND0, d_arr_relu_19_8=>GND0, d_arr_relu_19_7=>GND0, 
      d_arr_relu_19_6=>GND0, d_arr_relu_19_5=>GND0, d_arr_relu_19_4=>GND0, 
      d_arr_relu_19_3=>GND0, d_arr_relu_19_2=>GND0, d_arr_relu_19_1=>GND0, 
      d_arr_relu_19_0=>GND0, d_arr_relu_20_31=>GND0, d_arr_relu_20_30=>GND0, 
      d_arr_relu_20_29=>GND0, d_arr_relu_20_28=>GND0, d_arr_relu_20_27=>GND0, 
      d_arr_relu_20_26=>GND0, d_arr_relu_20_25=>GND0, d_arr_relu_20_24=>GND0, 
      d_arr_relu_20_23=>GND0, d_arr_relu_20_22=>GND0, d_arr_relu_20_21=>GND0, 
      d_arr_relu_20_20=>GND0, d_arr_relu_20_19=>GND0, d_arr_relu_20_18=>GND0, 
      d_arr_relu_20_17=>GND0, d_arr_relu_20_16=>GND0, d_arr_relu_20_15=>GND0, 
      d_arr_relu_20_14=>GND0, d_arr_relu_20_13=>GND0, d_arr_relu_20_12=>GND0, 
      d_arr_relu_20_11=>GND0, d_arr_relu_20_10=>GND0, d_arr_relu_20_9=>GND0, 
      d_arr_relu_20_8=>GND0, d_arr_relu_20_7=>GND0, d_arr_relu_20_6=>GND0, 
      d_arr_relu_20_5=>GND0, d_arr_relu_20_4=>GND0, d_arr_relu_20_3=>GND0, 
      d_arr_relu_20_2=>GND0, d_arr_relu_20_1=>GND0, d_arr_relu_20_0=>GND0, 
      d_arr_relu_21_31=>GND0, d_arr_relu_21_30=>GND0, d_arr_relu_21_29=>GND0, 
      d_arr_relu_21_28=>GND0, d_arr_relu_21_27=>GND0, d_arr_relu_21_26=>GND0, 
      d_arr_relu_21_25=>GND0, d_arr_relu_21_24=>GND0, d_arr_relu_21_23=>GND0, 
      d_arr_relu_21_22=>GND0, d_arr_relu_21_21=>GND0, d_arr_relu_21_20=>GND0, 
      d_arr_relu_21_19=>GND0, d_arr_relu_21_18=>GND0, d_arr_relu_21_17=>GND0, 
      d_arr_relu_21_16=>GND0, d_arr_relu_21_15=>GND0, d_arr_relu_21_14=>GND0, 
      d_arr_relu_21_13=>GND0, d_arr_relu_21_12=>GND0, d_arr_relu_21_11=>GND0, 
      d_arr_relu_21_10=>GND0, d_arr_relu_21_9=>GND0, d_arr_relu_21_8=>GND0, 
      d_arr_relu_21_7=>GND0, d_arr_relu_21_6=>GND0, d_arr_relu_21_5=>GND0, 
      d_arr_relu_21_4=>GND0, d_arr_relu_21_3=>GND0, d_arr_relu_21_2=>GND0, 
      d_arr_relu_21_1=>GND0, d_arr_relu_21_0=>GND0, d_arr_relu_22_31=>GND0, 
      d_arr_relu_22_30=>GND0, d_arr_relu_22_29=>GND0, d_arr_relu_22_28=>GND0, 
      d_arr_relu_22_27=>GND0, d_arr_relu_22_26=>GND0, d_arr_relu_22_25=>GND0, 
      d_arr_relu_22_24=>GND0, d_arr_relu_22_23=>GND0, d_arr_relu_22_22=>GND0, 
      d_arr_relu_22_21=>GND0, d_arr_relu_22_20=>GND0, d_arr_relu_22_19=>GND0, 
      d_arr_relu_22_18=>GND0, d_arr_relu_22_17=>GND0, d_arr_relu_22_16=>GND0, 
      d_arr_relu_22_15=>GND0, d_arr_relu_22_14=>GND0, d_arr_relu_22_13=>GND0, 
      d_arr_relu_22_12=>GND0, d_arr_relu_22_11=>GND0, d_arr_relu_22_10=>GND0, 
      d_arr_relu_22_9=>GND0, d_arr_relu_22_8=>GND0, d_arr_relu_22_7=>GND0, 
      d_arr_relu_22_6=>GND0, d_arr_relu_22_5=>GND0, d_arr_relu_22_4=>GND0, 
      d_arr_relu_22_3=>GND0, d_arr_relu_22_2=>GND0, d_arr_relu_22_1=>GND0, 
      d_arr_relu_22_0=>GND0, d_arr_relu_23_31=>GND0, d_arr_relu_23_30=>GND0, 
      d_arr_relu_23_29=>GND0, d_arr_relu_23_28=>GND0, d_arr_relu_23_27=>GND0, 
      d_arr_relu_23_26=>GND0, d_arr_relu_23_25=>GND0, d_arr_relu_23_24=>GND0, 
      d_arr_relu_23_23=>GND0, d_arr_relu_23_22=>GND0, d_arr_relu_23_21=>GND0, 
      d_arr_relu_23_20=>GND0, d_arr_relu_23_19=>GND0, d_arr_relu_23_18=>GND0, 
      d_arr_relu_23_17=>GND0, d_arr_relu_23_16=>GND0, d_arr_relu_23_15=>GND0, 
      d_arr_relu_23_14=>GND0, d_arr_relu_23_13=>GND0, d_arr_relu_23_12=>GND0, 
      d_arr_relu_23_11=>GND0, d_arr_relu_23_10=>GND0, d_arr_relu_23_9=>GND0, 
      d_arr_relu_23_8=>GND0, d_arr_relu_23_7=>GND0, d_arr_relu_23_6=>GND0, 
      d_arr_relu_23_5=>GND0, d_arr_relu_23_4=>GND0, d_arr_relu_23_3=>GND0, 
      d_arr_relu_23_2=>GND0, d_arr_relu_23_1=>GND0, d_arr_relu_23_0=>GND0, 
      d_arr_relu_24_31=>GND0, d_arr_relu_24_30=>GND0, d_arr_relu_24_29=>GND0, 
      d_arr_relu_24_28=>GND0, d_arr_relu_24_27=>GND0, d_arr_relu_24_26=>GND0, 
      d_arr_relu_24_25=>GND0, d_arr_relu_24_24=>GND0, d_arr_relu_24_23=>GND0, 
      d_arr_relu_24_22=>GND0, d_arr_relu_24_21=>GND0, d_arr_relu_24_20=>GND0, 
      d_arr_relu_24_19=>GND0, d_arr_relu_24_18=>GND0, d_arr_relu_24_17=>GND0, 
      d_arr_relu_24_16=>GND0, d_arr_relu_24_15=>GND0, d_arr_relu_24_14=>GND0, 
      d_arr_relu_24_13=>GND0, d_arr_relu_24_12=>GND0, d_arr_relu_24_11=>GND0, 
      d_arr_relu_24_10=>GND0, d_arr_relu_24_9=>GND0, d_arr_relu_24_8=>GND0, 
      d_arr_relu_24_7=>GND0, d_arr_relu_24_6=>GND0, d_arr_relu_24_5=>GND0, 
      d_arr_relu_24_4=>GND0, d_arr_relu_24_3=>GND0, d_arr_relu_24_2=>GND0, 
      d_arr_relu_24_1=>GND0, d_arr_relu_24_0=>GND0, sel_mux=>counter_0, 
      sel_mul=>nx16627, sel_add=>sel_add, sel_merge1=>counter_13, sel_merge2
      =>counter_14, sel_relu=>counter_15, d_arr_0_31=>d_arr_0_31, d_arr_0_30
      =>d_arr_0_30, d_arr_0_29=>d_arr_0_29, d_arr_0_28=>d_arr_0_28, 
      d_arr_0_27=>d_arr_0_27, d_arr_0_26=>d_arr_0_26, d_arr_0_25=>d_arr_0_25, 
      d_arr_0_24=>d_arr_0_24, d_arr_0_23=>d_arr_0_23, d_arr_0_22=>d_arr_0_22, 
      d_arr_0_21=>d_arr_0_21, d_arr_0_20=>d_arr_0_20, d_arr_0_19=>d_arr_0_19, 
      d_arr_0_18=>d_arr_0_18, d_arr_0_17=>d_arr_0_17, d_arr_0_16=>d_arr_0_16, 
      d_arr_0_15=>d_arr_0_15, d_arr_0_14=>d_arr_0_14, d_arr_0_13=>d_arr_0_13, 
      d_arr_0_12=>d_arr_0_12, d_arr_0_11=>d_arr_0_11, d_arr_0_10=>d_arr_0_10, 
      d_arr_0_9=>d_arr_0_9, d_arr_0_8=>d_arr_0_8, d_arr_0_7=>d_arr_0_7, 
      d_arr_0_6=>d_arr_0_6, d_arr_0_5=>d_arr_0_5, d_arr_0_4=>d_arr_0_4, 
      d_arr_0_3=>d_arr_0_3, d_arr_0_2=>d_arr_0_2, d_arr_0_1=>d_arr_0_1, 
      d_arr_0_0=>d_arr_0_0, d_arr_1_31=>d_arr_1_31, d_arr_1_30=>d_arr_1_30, 
      d_arr_1_29=>d_arr_1_29, d_arr_1_28=>d_arr_1_28, d_arr_1_27=>d_arr_1_27, 
      d_arr_1_26=>d_arr_1_26, d_arr_1_25=>d_arr_1_25, d_arr_1_24=>d_arr_1_24, 
      d_arr_1_23=>d_arr_1_23, d_arr_1_22=>d_arr_1_22, d_arr_1_21=>d_arr_1_21, 
      d_arr_1_20=>d_arr_1_20, d_arr_1_19=>d_arr_1_19, d_arr_1_18=>d_arr_1_18, 
      d_arr_1_17=>d_arr_1_17, d_arr_1_16=>d_arr_1_16, d_arr_1_15=>d_arr_1_15, 
      d_arr_1_14=>d_arr_1_14, d_arr_1_13=>d_arr_1_13, d_arr_1_12=>d_arr_1_12, 
      d_arr_1_11=>d_arr_1_11, d_arr_1_10=>d_arr_1_10, d_arr_1_9=>d_arr_1_9, 
      d_arr_1_8=>d_arr_1_8, d_arr_1_7=>d_arr_1_7, d_arr_1_6=>d_arr_1_6, 
      d_arr_1_5=>d_arr_1_5, d_arr_1_4=>d_arr_1_4, d_arr_1_3=>d_arr_1_3, 
      d_arr_1_2=>d_arr_1_2, d_arr_1_1=>d_arr_1_1, d_arr_1_0=>d_arr_1_0, 
      d_arr_2_31=>d_arr_2_31, d_arr_2_30=>d_arr_2_30, d_arr_2_29=>d_arr_2_29, 
      d_arr_2_28=>d_arr_2_28, d_arr_2_27=>d_arr_2_27, d_arr_2_26=>d_arr_2_26, 
      d_arr_2_25=>d_arr_2_25, d_arr_2_24=>d_arr_2_24, d_arr_2_23=>d_arr_2_23, 
      d_arr_2_22=>d_arr_2_22, d_arr_2_21=>d_arr_2_21, d_arr_2_20=>d_arr_2_20, 
      d_arr_2_19=>d_arr_2_19, d_arr_2_18=>d_arr_2_18, d_arr_2_17=>d_arr_2_17, 
      d_arr_2_16=>d_arr_2_16, d_arr_2_15=>d_arr_2_15, d_arr_2_14=>d_arr_2_14, 
      d_arr_2_13=>d_arr_2_13, d_arr_2_12=>d_arr_2_12, d_arr_2_11=>d_arr_2_11, 
      d_arr_2_10=>d_arr_2_10, d_arr_2_9=>d_arr_2_9, d_arr_2_8=>d_arr_2_8, 
      d_arr_2_7=>d_arr_2_7, d_arr_2_6=>d_arr_2_6, d_arr_2_5=>d_arr_2_5, 
      d_arr_2_4=>d_arr_2_4, d_arr_2_3=>d_arr_2_3, d_arr_2_2=>d_arr_2_2, 
      d_arr_2_1=>d_arr_2_1, d_arr_2_0=>d_arr_2_0, d_arr_3_31=>d_arr_3_31, 
      d_arr_3_30=>d_arr_3_30, d_arr_3_29=>d_arr_3_29, d_arr_3_28=>d_arr_3_28, 
      d_arr_3_27=>d_arr_3_27, d_arr_3_26=>d_arr_3_26, d_arr_3_25=>d_arr_3_25, 
      d_arr_3_24=>d_arr_3_24, d_arr_3_23=>d_arr_3_23, d_arr_3_22=>d_arr_3_22, 
      d_arr_3_21=>d_arr_3_21, d_arr_3_20=>d_arr_3_20, d_arr_3_19=>d_arr_3_19, 
      d_arr_3_18=>d_arr_3_18, d_arr_3_17=>d_arr_3_17, d_arr_3_16=>d_arr_3_16, 
      d_arr_3_15=>d_arr_3_15, d_arr_3_14=>d_arr_3_14, d_arr_3_13=>d_arr_3_13, 
      d_arr_3_12=>d_arr_3_12, d_arr_3_11=>d_arr_3_11, d_arr_3_10=>d_arr_3_10, 
      d_arr_3_9=>d_arr_3_9, d_arr_3_8=>d_arr_3_8, d_arr_3_7=>d_arr_3_7, 
      d_arr_3_6=>d_arr_3_6, d_arr_3_5=>d_arr_3_5, d_arr_3_4=>d_arr_3_4, 
      d_arr_3_3=>d_arr_3_3, d_arr_3_2=>d_arr_3_2, d_arr_3_1=>d_arr_3_1, 
      d_arr_3_0=>d_arr_3_0, d_arr_4_31=>d_arr_4_31, d_arr_4_30=>d_arr_4_30, 
      d_arr_4_29=>d_arr_4_29, d_arr_4_28=>d_arr_4_28, d_arr_4_27=>d_arr_4_27, 
      d_arr_4_26=>d_arr_4_26, d_arr_4_25=>d_arr_4_25, d_arr_4_24=>d_arr_4_24, 
      d_arr_4_23=>d_arr_4_23, d_arr_4_22=>d_arr_4_22, d_arr_4_21=>d_arr_4_21, 
      d_arr_4_20=>d_arr_4_20, d_arr_4_19=>d_arr_4_19, d_arr_4_18=>d_arr_4_18, 
      d_arr_4_17=>d_arr_4_17, d_arr_4_16=>d_arr_4_16, d_arr_4_15=>d_arr_4_15, 
      d_arr_4_14=>d_arr_4_14, d_arr_4_13=>d_arr_4_13, d_arr_4_12=>d_arr_4_12, 
      d_arr_4_11=>d_arr_4_11, d_arr_4_10=>d_arr_4_10, d_arr_4_9=>d_arr_4_9, 
      d_arr_4_8=>d_arr_4_8, d_arr_4_7=>d_arr_4_7, d_arr_4_6=>d_arr_4_6, 
      d_arr_4_5=>d_arr_4_5, d_arr_4_4=>d_arr_4_4, d_arr_4_3=>d_arr_4_3, 
      d_arr_4_2=>d_arr_4_2, d_arr_4_1=>d_arr_4_1, d_arr_4_0=>d_arr_4_0, 
      d_arr_5_31=>d_arr_5_31, d_arr_5_30=>d_arr_5_30, d_arr_5_29=>d_arr_5_29, 
      d_arr_5_28=>d_arr_5_28, d_arr_5_27=>d_arr_5_27, d_arr_5_26=>d_arr_5_26, 
      d_arr_5_25=>d_arr_5_25, d_arr_5_24=>d_arr_5_24, d_arr_5_23=>d_arr_5_23, 
      d_arr_5_22=>d_arr_5_22, d_arr_5_21=>d_arr_5_21, d_arr_5_20=>d_arr_5_20, 
      d_arr_5_19=>d_arr_5_19, d_arr_5_18=>d_arr_5_18, d_arr_5_17=>d_arr_5_17, 
      d_arr_5_16=>d_arr_5_16, d_arr_5_15=>d_arr_5_15, d_arr_5_14=>d_arr_5_14, 
      d_arr_5_13=>d_arr_5_13, d_arr_5_12=>d_arr_5_12, d_arr_5_11=>d_arr_5_11, 
      d_arr_5_10=>d_arr_5_10, d_arr_5_9=>d_arr_5_9, d_arr_5_8=>d_arr_5_8, 
      d_arr_5_7=>d_arr_5_7, d_arr_5_6=>d_arr_5_6, d_arr_5_5=>d_arr_5_5, 
      d_arr_5_4=>d_arr_5_4, d_arr_5_3=>d_arr_5_3, d_arr_5_2=>d_arr_5_2, 
      d_arr_5_1=>d_arr_5_1, d_arr_5_0=>d_arr_5_0, d_arr_6_31=>d_arr_6_31, 
      d_arr_6_30=>d_arr_6_30, d_arr_6_29=>d_arr_6_29, d_arr_6_28=>d_arr_6_28, 
      d_arr_6_27=>d_arr_6_27, d_arr_6_26=>d_arr_6_26, d_arr_6_25=>d_arr_6_25, 
      d_arr_6_24=>d_arr_6_24, d_arr_6_23=>d_arr_6_23, d_arr_6_22=>d_arr_6_22, 
      d_arr_6_21=>d_arr_6_21, d_arr_6_20=>d_arr_6_20, d_arr_6_19=>d_arr_6_19, 
      d_arr_6_18=>d_arr_6_18, d_arr_6_17=>d_arr_6_17, d_arr_6_16=>d_arr_6_16, 
      d_arr_6_15=>d_arr_6_15, d_arr_6_14=>d_arr_6_14, d_arr_6_13=>d_arr_6_13, 
      d_arr_6_12=>d_arr_6_12, d_arr_6_11=>d_arr_6_11, d_arr_6_10=>d_arr_6_10, 
      d_arr_6_9=>d_arr_6_9, d_arr_6_8=>d_arr_6_8, d_arr_6_7=>d_arr_6_7, 
      d_arr_6_6=>d_arr_6_6, d_arr_6_5=>d_arr_6_5, d_arr_6_4=>d_arr_6_4, 
      d_arr_6_3=>d_arr_6_3, d_arr_6_2=>d_arr_6_2, d_arr_6_1=>d_arr_6_1, 
      d_arr_6_0=>d_arr_6_0, d_arr_7_31=>d_arr_7_31, d_arr_7_30=>d_arr_7_30, 
      d_arr_7_29=>d_arr_7_29, d_arr_7_28=>d_arr_7_28, d_arr_7_27=>d_arr_7_27, 
      d_arr_7_26=>d_arr_7_26, d_arr_7_25=>d_arr_7_25, d_arr_7_24=>d_arr_7_24, 
      d_arr_7_23=>d_arr_7_23, d_arr_7_22=>d_arr_7_22, d_arr_7_21=>d_arr_7_21, 
      d_arr_7_20=>d_arr_7_20, d_arr_7_19=>d_arr_7_19, d_arr_7_18=>d_arr_7_18, 
      d_arr_7_17=>d_arr_7_17, d_arr_7_16=>d_arr_7_16, d_arr_7_15=>d_arr_7_15, 
      d_arr_7_14=>d_arr_7_14, d_arr_7_13=>d_arr_7_13, d_arr_7_12=>d_arr_7_12, 
      d_arr_7_11=>d_arr_7_11, d_arr_7_10=>d_arr_7_10, d_arr_7_9=>d_arr_7_9, 
      d_arr_7_8=>d_arr_7_8, d_arr_7_7=>d_arr_7_7, d_arr_7_6=>d_arr_7_6, 
      d_arr_7_5=>d_arr_7_5, d_arr_7_4=>d_arr_7_4, d_arr_7_3=>d_arr_7_3, 
      d_arr_7_2=>d_arr_7_2, d_arr_7_1=>d_arr_7_1, d_arr_7_0=>d_arr_7_0, 
      d_arr_8_31=>d_arr_8_31, d_arr_8_30=>d_arr_8_30, d_arr_8_29=>d_arr_8_29, 
      d_arr_8_28=>d_arr_8_28, d_arr_8_27=>d_arr_8_27, d_arr_8_26=>d_arr_8_26, 
      d_arr_8_25=>d_arr_8_25, d_arr_8_24=>d_arr_8_24, d_arr_8_23=>d_arr_8_23, 
      d_arr_8_22=>d_arr_8_22, d_arr_8_21=>d_arr_8_21, d_arr_8_20=>d_arr_8_20, 
      d_arr_8_19=>d_arr_8_19, d_arr_8_18=>d_arr_8_18, d_arr_8_17=>d_arr_8_17, 
      d_arr_8_16=>d_arr_8_16, d_arr_8_15=>d_arr_8_15, d_arr_8_14=>d_arr_8_14, 
      d_arr_8_13=>d_arr_8_13, d_arr_8_12=>d_arr_8_12, d_arr_8_11=>d_arr_8_11, 
      d_arr_8_10=>d_arr_8_10, d_arr_8_9=>d_arr_8_9, d_arr_8_8=>d_arr_8_8, 
      d_arr_8_7=>d_arr_8_7, d_arr_8_6=>d_arr_8_6, d_arr_8_5=>d_arr_8_5, 
      d_arr_8_4=>d_arr_8_4, d_arr_8_3=>d_arr_8_3, d_arr_8_2=>d_arr_8_2, 
      d_arr_8_1=>d_arr_8_1, d_arr_8_0=>d_arr_8_0, d_arr_9_31=>d_arr_9_31, 
      d_arr_9_30=>d_arr_9_30, d_arr_9_29=>d_arr_9_29, d_arr_9_28=>d_arr_9_28, 
      d_arr_9_27=>d_arr_9_27, d_arr_9_26=>d_arr_9_26, d_arr_9_25=>d_arr_9_25, 
      d_arr_9_24=>d_arr_9_24, d_arr_9_23=>d_arr_9_23, d_arr_9_22=>d_arr_9_22, 
      d_arr_9_21=>d_arr_9_21, d_arr_9_20=>d_arr_9_20, d_arr_9_19=>d_arr_9_19, 
      d_arr_9_18=>d_arr_9_18, d_arr_9_17=>d_arr_9_17, d_arr_9_16=>d_arr_9_16, 
      d_arr_9_15=>d_arr_9_15, d_arr_9_14=>d_arr_9_14, d_arr_9_13=>d_arr_9_13, 
      d_arr_9_12=>d_arr_9_12, d_arr_9_11=>d_arr_9_11, d_arr_9_10=>d_arr_9_10, 
      d_arr_9_9=>d_arr_9_9, d_arr_9_8=>d_arr_9_8, d_arr_9_7=>d_arr_9_7, 
      d_arr_9_6=>d_arr_9_6, d_arr_9_5=>d_arr_9_5, d_arr_9_4=>d_arr_9_4, 
      d_arr_9_3=>d_arr_9_3, d_arr_9_2=>d_arr_9_2, d_arr_9_1=>d_arr_9_1, 
      d_arr_9_0=>d_arr_9_0, d_arr_10_31=>d_arr_10_31, d_arr_10_30=>
      d_arr_10_30, d_arr_10_29=>d_arr_10_29, d_arr_10_28=>d_arr_10_28, 
      d_arr_10_27=>d_arr_10_27, d_arr_10_26=>d_arr_10_26, d_arr_10_25=>
      d_arr_10_25, d_arr_10_24=>d_arr_10_24, d_arr_10_23=>d_arr_10_23, 
      d_arr_10_22=>d_arr_10_22, d_arr_10_21=>d_arr_10_21, d_arr_10_20=>
      d_arr_10_20, d_arr_10_19=>d_arr_10_19, d_arr_10_18=>d_arr_10_18, 
      d_arr_10_17=>d_arr_10_17, d_arr_10_16=>d_arr_10_16, d_arr_10_15=>
      d_arr_10_15, d_arr_10_14=>d_arr_10_14, d_arr_10_13=>d_arr_10_13, 
      d_arr_10_12=>d_arr_10_12, d_arr_10_11=>d_arr_10_11, d_arr_10_10=>
      d_arr_10_10, d_arr_10_9=>d_arr_10_9, d_arr_10_8=>d_arr_10_8, 
      d_arr_10_7=>d_arr_10_7, d_arr_10_6=>d_arr_10_6, d_arr_10_5=>d_arr_10_5, 
      d_arr_10_4=>d_arr_10_4, d_arr_10_3=>d_arr_10_3, d_arr_10_2=>d_arr_10_2, 
      d_arr_10_1=>d_arr_10_1, d_arr_10_0=>d_arr_10_0, d_arr_11_31=>
      d_arr_11_31, d_arr_11_30=>d_arr_11_30, d_arr_11_29=>d_arr_11_29, 
      d_arr_11_28=>d_arr_11_28, d_arr_11_27=>d_arr_11_27, d_arr_11_26=>
      d_arr_11_26, d_arr_11_25=>d_arr_11_25, d_arr_11_24=>d_arr_11_24, 
      d_arr_11_23=>d_arr_11_23, d_arr_11_22=>d_arr_11_22, d_arr_11_21=>
      d_arr_11_21, d_arr_11_20=>d_arr_11_20, d_arr_11_19=>d_arr_11_19, 
      d_arr_11_18=>d_arr_11_18, d_arr_11_17=>d_arr_11_17, d_arr_11_16=>
      d_arr_11_16, d_arr_11_15=>d_arr_11_15, d_arr_11_14=>d_arr_11_14, 
      d_arr_11_13=>d_arr_11_13, d_arr_11_12=>d_arr_11_12, d_arr_11_11=>
      d_arr_11_11, d_arr_11_10=>d_arr_11_10, d_arr_11_9=>d_arr_11_9, 
      d_arr_11_8=>d_arr_11_8, d_arr_11_7=>d_arr_11_7, d_arr_11_6=>d_arr_11_6, 
      d_arr_11_5=>d_arr_11_5, d_arr_11_4=>d_arr_11_4, d_arr_11_3=>d_arr_11_3, 
      d_arr_11_2=>d_arr_11_2, d_arr_11_1=>d_arr_11_1, d_arr_11_0=>d_arr_11_0, 
      d_arr_12_31=>d_arr_12_31, d_arr_12_30=>d_arr_12_30, d_arr_12_29=>
      d_arr_12_29, d_arr_12_28=>d_arr_12_28, d_arr_12_27=>d_arr_12_27, 
      d_arr_12_26=>d_arr_12_26, d_arr_12_25=>d_arr_12_25, d_arr_12_24=>
      d_arr_12_24, d_arr_12_23=>d_arr_12_23, d_arr_12_22=>d_arr_12_22, 
      d_arr_12_21=>d_arr_12_21, d_arr_12_20=>d_arr_12_20, d_arr_12_19=>
      d_arr_12_19, d_arr_12_18=>d_arr_12_18, d_arr_12_17=>d_arr_12_17, 
      d_arr_12_16=>d_arr_12_16, d_arr_12_15=>d_arr_12_15, d_arr_12_14=>
      d_arr_12_14, d_arr_12_13=>d_arr_12_13, d_arr_12_12=>d_arr_12_12, 
      d_arr_12_11=>d_arr_12_11, d_arr_12_10=>d_arr_12_10, d_arr_12_9=>
      d_arr_12_9, d_arr_12_8=>d_arr_12_8, d_arr_12_7=>d_arr_12_7, d_arr_12_6
      =>d_arr_12_6, d_arr_12_5=>d_arr_12_5, d_arr_12_4=>d_arr_12_4, 
      d_arr_12_3=>d_arr_12_3, d_arr_12_2=>d_arr_12_2, d_arr_12_1=>d_arr_12_1, 
      d_arr_12_0=>d_arr_12_0, d_arr_13_31=>d_arr_13_31, d_arr_13_30=>
      d_arr_13_30, d_arr_13_29=>d_arr_13_29, d_arr_13_28=>d_arr_13_28, 
      d_arr_13_27=>d_arr_13_27, d_arr_13_26=>d_arr_13_26, d_arr_13_25=>
      d_arr_13_25, d_arr_13_24=>d_arr_13_24, d_arr_13_23=>d_arr_13_23, 
      d_arr_13_22=>d_arr_13_22, d_arr_13_21=>d_arr_13_21, d_arr_13_20=>
      d_arr_13_20, d_arr_13_19=>d_arr_13_19, d_arr_13_18=>d_arr_13_18, 
      d_arr_13_17=>d_arr_13_17, d_arr_13_16=>d_arr_13_16, d_arr_13_15=>
      d_arr_13_15, d_arr_13_14=>d_arr_13_14, d_arr_13_13=>d_arr_13_13, 
      d_arr_13_12=>d_arr_13_12, d_arr_13_11=>d_arr_13_11, d_arr_13_10=>
      d_arr_13_10, d_arr_13_9=>d_arr_13_9, d_arr_13_8=>d_arr_13_8, 
      d_arr_13_7=>d_arr_13_7, d_arr_13_6=>d_arr_13_6, d_arr_13_5=>d_arr_13_5, 
      d_arr_13_4=>d_arr_13_4, d_arr_13_3=>d_arr_13_3, d_arr_13_2=>d_arr_13_2, 
      d_arr_13_1=>d_arr_13_1, d_arr_13_0=>d_arr_13_0, d_arr_14_31=>
      d_arr_14_31, d_arr_14_30=>d_arr_14_30, d_arr_14_29=>d_arr_14_29, 
      d_arr_14_28=>d_arr_14_28, d_arr_14_27=>d_arr_14_27, d_arr_14_26=>
      d_arr_14_26, d_arr_14_25=>d_arr_14_25, d_arr_14_24=>d_arr_14_24, 
      d_arr_14_23=>d_arr_14_23, d_arr_14_22=>d_arr_14_22, d_arr_14_21=>
      d_arr_14_21, d_arr_14_20=>d_arr_14_20, d_arr_14_19=>d_arr_14_19, 
      d_arr_14_18=>d_arr_14_18, d_arr_14_17=>d_arr_14_17, d_arr_14_16=>
      d_arr_14_16, d_arr_14_15=>d_arr_14_15, d_arr_14_14=>d_arr_14_14, 
      d_arr_14_13=>d_arr_14_13, d_arr_14_12=>d_arr_14_12, d_arr_14_11=>
      d_arr_14_11, d_arr_14_10=>d_arr_14_10, d_arr_14_9=>d_arr_14_9, 
      d_arr_14_8=>d_arr_14_8, d_arr_14_7=>d_arr_14_7, d_arr_14_6=>d_arr_14_6, 
      d_arr_14_5=>d_arr_14_5, d_arr_14_4=>d_arr_14_4, d_arr_14_3=>d_arr_14_3, 
      d_arr_14_2=>d_arr_14_2, d_arr_14_1=>d_arr_14_1, d_arr_14_0=>d_arr_14_0, 
      d_arr_15_31=>d_arr_15_31, d_arr_15_30=>d_arr_15_30, d_arr_15_29=>
      d_arr_15_29, d_arr_15_28=>d_arr_15_28, d_arr_15_27=>d_arr_15_27, 
      d_arr_15_26=>d_arr_15_26, d_arr_15_25=>d_arr_15_25, d_arr_15_24=>
      d_arr_15_24, d_arr_15_23=>d_arr_15_23, d_arr_15_22=>d_arr_15_22, 
      d_arr_15_21=>d_arr_15_21, d_arr_15_20=>d_arr_15_20, d_arr_15_19=>
      d_arr_15_19, d_arr_15_18=>d_arr_15_18, d_arr_15_17=>d_arr_15_17, 
      d_arr_15_16=>d_arr_15_16, d_arr_15_15=>d_arr_15_15, d_arr_15_14=>
      d_arr_15_14, d_arr_15_13=>d_arr_15_13, d_arr_15_12=>d_arr_15_12, 
      d_arr_15_11=>d_arr_15_11, d_arr_15_10=>d_arr_15_10, d_arr_15_9=>
      d_arr_15_9, d_arr_15_8=>d_arr_15_8, d_arr_15_7=>d_arr_15_7, d_arr_15_6
      =>d_arr_15_6, d_arr_15_5=>d_arr_15_5, d_arr_15_4=>d_arr_15_4, 
      d_arr_15_3=>d_arr_15_3, d_arr_15_2=>d_arr_15_2, d_arr_15_1=>d_arr_15_1, 
      d_arr_15_0=>d_arr_15_0, d_arr_16_31=>d_arr_16_31, d_arr_16_30=>
      d_arr_16_30, d_arr_16_29=>d_arr_16_29, d_arr_16_28=>d_arr_16_28, 
      d_arr_16_27=>d_arr_16_27, d_arr_16_26=>d_arr_16_26, d_arr_16_25=>
      d_arr_16_25, d_arr_16_24=>d_arr_16_24, d_arr_16_23=>d_arr_16_23, 
      d_arr_16_22=>d_arr_16_22, d_arr_16_21=>d_arr_16_21, d_arr_16_20=>
      d_arr_16_20, d_arr_16_19=>d_arr_16_19, d_arr_16_18=>d_arr_16_18, 
      d_arr_16_17=>d_arr_16_17, d_arr_16_16=>d_arr_16_16, d_arr_16_15=>
      d_arr_16_15, d_arr_16_14=>d_arr_16_14, d_arr_16_13=>d_arr_16_13, 
      d_arr_16_12=>d_arr_16_12, d_arr_16_11=>d_arr_16_11, d_arr_16_10=>
      d_arr_16_10, d_arr_16_9=>d_arr_16_9, d_arr_16_8=>d_arr_16_8, 
      d_arr_16_7=>d_arr_16_7, d_arr_16_6=>d_arr_16_6, d_arr_16_5=>d_arr_16_5, 
      d_arr_16_4=>d_arr_16_4, d_arr_16_3=>d_arr_16_3, d_arr_16_2=>d_arr_16_2, 
      d_arr_16_1=>d_arr_16_1, d_arr_16_0=>d_arr_16_0, d_arr_17_31=>
      d_arr_17_31, d_arr_17_30=>d_arr_17_30, d_arr_17_29=>d_arr_17_29, 
      d_arr_17_28=>d_arr_17_28, d_arr_17_27=>d_arr_17_27, d_arr_17_26=>
      d_arr_17_26, d_arr_17_25=>d_arr_17_25, d_arr_17_24=>d_arr_17_24, 
      d_arr_17_23=>d_arr_17_23, d_arr_17_22=>d_arr_17_22, d_arr_17_21=>
      d_arr_17_21, d_arr_17_20=>d_arr_17_20, d_arr_17_19=>d_arr_17_19, 
      d_arr_17_18=>d_arr_17_18, d_arr_17_17=>d_arr_17_17, d_arr_17_16=>
      d_arr_17_16, d_arr_17_15=>d_arr_17_15, d_arr_17_14=>d_arr_17_14, 
      d_arr_17_13=>d_arr_17_13, d_arr_17_12=>d_arr_17_12, d_arr_17_11=>
      d_arr_17_11, d_arr_17_10=>d_arr_17_10, d_arr_17_9=>d_arr_17_9, 
      d_arr_17_8=>d_arr_17_8, d_arr_17_7=>d_arr_17_7, d_arr_17_6=>d_arr_17_6, 
      d_arr_17_5=>d_arr_17_5, d_arr_17_4=>d_arr_17_4, d_arr_17_3=>d_arr_17_3, 
      d_arr_17_2=>d_arr_17_2, d_arr_17_1=>d_arr_17_1, d_arr_17_0=>d_arr_17_0, 
      d_arr_18_31=>d_arr_18_31, d_arr_18_30=>d_arr_18_30, d_arr_18_29=>
      d_arr_18_29, d_arr_18_28=>d_arr_18_28, d_arr_18_27=>d_arr_18_27, 
      d_arr_18_26=>d_arr_18_26, d_arr_18_25=>d_arr_18_25, d_arr_18_24=>
      d_arr_18_24, d_arr_18_23=>d_arr_18_23, d_arr_18_22=>d_arr_18_22, 
      d_arr_18_21=>d_arr_18_21, d_arr_18_20=>d_arr_18_20, d_arr_18_19=>
      d_arr_18_19, d_arr_18_18=>d_arr_18_18, d_arr_18_17=>d_arr_18_17, 
      d_arr_18_16=>d_arr_18_16, d_arr_18_15=>d_arr_18_15, d_arr_18_14=>
      d_arr_18_14, d_arr_18_13=>d_arr_18_13, d_arr_18_12=>d_arr_18_12, 
      d_arr_18_11=>d_arr_18_11, d_arr_18_10=>d_arr_18_10, d_arr_18_9=>
      d_arr_18_9, d_arr_18_8=>d_arr_18_8, d_arr_18_7=>d_arr_18_7, d_arr_18_6
      =>d_arr_18_6, d_arr_18_5=>d_arr_18_5, d_arr_18_4=>d_arr_18_4, 
      d_arr_18_3=>d_arr_18_3, d_arr_18_2=>d_arr_18_2, d_arr_18_1=>d_arr_18_1, 
      d_arr_18_0=>d_arr_18_0, d_arr_19_31=>d_arr_19_31, d_arr_19_30=>
      d_arr_19_30, d_arr_19_29=>d_arr_19_29, d_arr_19_28=>d_arr_19_28, 
      d_arr_19_27=>d_arr_19_27, d_arr_19_26=>d_arr_19_26, d_arr_19_25=>
      d_arr_19_25, d_arr_19_24=>d_arr_19_24, d_arr_19_23=>d_arr_19_23, 
      d_arr_19_22=>d_arr_19_22, d_arr_19_21=>d_arr_19_21, d_arr_19_20=>
      d_arr_19_20, d_arr_19_19=>d_arr_19_19, d_arr_19_18=>d_arr_19_18, 
      d_arr_19_17=>d_arr_19_17, d_arr_19_16=>d_arr_19_16, d_arr_19_15=>
      d_arr_19_15, d_arr_19_14=>d_arr_19_14, d_arr_19_13=>d_arr_19_13, 
      d_arr_19_12=>d_arr_19_12, d_arr_19_11=>d_arr_19_11, d_arr_19_10=>
      d_arr_19_10, d_arr_19_9=>d_arr_19_9, d_arr_19_8=>d_arr_19_8, 
      d_arr_19_7=>d_arr_19_7, d_arr_19_6=>d_arr_19_6, d_arr_19_5=>d_arr_19_5, 
      d_arr_19_4=>d_arr_19_4, d_arr_19_3=>d_arr_19_3, d_arr_19_2=>d_arr_19_2, 
      d_arr_19_1=>d_arr_19_1, d_arr_19_0=>d_arr_19_0, d_arr_20_31=>
      d_arr_20_31, d_arr_20_30=>d_arr_20_30, d_arr_20_29=>d_arr_20_29, 
      d_arr_20_28=>d_arr_20_28, d_arr_20_27=>d_arr_20_27, d_arr_20_26=>
      d_arr_20_26, d_arr_20_25=>d_arr_20_25, d_arr_20_24=>d_arr_20_24, 
      d_arr_20_23=>d_arr_20_23, d_arr_20_22=>d_arr_20_22, d_arr_20_21=>
      d_arr_20_21, d_arr_20_20=>d_arr_20_20, d_arr_20_19=>d_arr_20_19, 
      d_arr_20_18=>d_arr_20_18, d_arr_20_17=>d_arr_20_17, d_arr_20_16=>
      d_arr_20_16, d_arr_20_15=>d_arr_20_15, d_arr_20_14=>d_arr_20_14, 
      d_arr_20_13=>d_arr_20_13, d_arr_20_12=>d_arr_20_12, d_arr_20_11=>
      d_arr_20_11, d_arr_20_10=>d_arr_20_10, d_arr_20_9=>d_arr_20_9, 
      d_arr_20_8=>d_arr_20_8, d_arr_20_7=>d_arr_20_7, d_arr_20_6=>d_arr_20_6, 
      d_arr_20_5=>d_arr_20_5, d_arr_20_4=>d_arr_20_4, d_arr_20_3=>d_arr_20_3, 
      d_arr_20_2=>d_arr_20_2, d_arr_20_1=>d_arr_20_1, d_arr_20_0=>d_arr_20_0, 
      d_arr_21_31=>d_arr_21_31, d_arr_21_30=>d_arr_21_30, d_arr_21_29=>
      d_arr_21_29, d_arr_21_28=>d_arr_21_28, d_arr_21_27=>d_arr_21_27, 
      d_arr_21_26=>d_arr_21_26, d_arr_21_25=>d_arr_21_25, d_arr_21_24=>
      d_arr_21_24, d_arr_21_23=>d_arr_21_23, d_arr_21_22=>d_arr_21_22, 
      d_arr_21_21=>d_arr_21_21, d_arr_21_20=>d_arr_21_20, d_arr_21_19=>
      d_arr_21_19, d_arr_21_18=>d_arr_21_18, d_arr_21_17=>d_arr_21_17, 
      d_arr_21_16=>d_arr_21_16, d_arr_21_15=>d_arr_21_15, d_arr_21_14=>
      d_arr_21_14, d_arr_21_13=>d_arr_21_13, d_arr_21_12=>d_arr_21_12, 
      d_arr_21_11=>d_arr_21_11, d_arr_21_10=>d_arr_21_10, d_arr_21_9=>
      d_arr_21_9, d_arr_21_8=>d_arr_21_8, d_arr_21_7=>d_arr_21_7, d_arr_21_6
      =>d_arr_21_6, d_arr_21_5=>d_arr_21_5, d_arr_21_4=>d_arr_21_4, 
      d_arr_21_3=>d_arr_21_3, d_arr_21_2=>d_arr_21_2, d_arr_21_1=>d_arr_21_1, 
      d_arr_21_0=>d_arr_21_0, d_arr_22_31=>d_arr_22_31, d_arr_22_30=>
      d_arr_22_30, d_arr_22_29=>d_arr_22_29, d_arr_22_28=>d_arr_22_28, 
      d_arr_22_27=>d_arr_22_27, d_arr_22_26=>d_arr_22_26, d_arr_22_25=>
      d_arr_22_25, d_arr_22_24=>d_arr_22_24, d_arr_22_23=>d_arr_22_23, 
      d_arr_22_22=>d_arr_22_22, d_arr_22_21=>d_arr_22_21, d_arr_22_20=>
      d_arr_22_20, d_arr_22_19=>d_arr_22_19, d_arr_22_18=>d_arr_22_18, 
      d_arr_22_17=>d_arr_22_17, d_arr_22_16=>d_arr_22_16, d_arr_22_15=>
      d_arr_22_15, d_arr_22_14=>d_arr_22_14, d_arr_22_13=>d_arr_22_13, 
      d_arr_22_12=>d_arr_22_12, d_arr_22_11=>d_arr_22_11, d_arr_22_10=>
      d_arr_22_10, d_arr_22_9=>d_arr_22_9, d_arr_22_8=>d_arr_22_8, 
      d_arr_22_7=>d_arr_22_7, d_arr_22_6=>d_arr_22_6, d_arr_22_5=>d_arr_22_5, 
      d_arr_22_4=>d_arr_22_4, d_arr_22_3=>d_arr_22_3, d_arr_22_2=>d_arr_22_2, 
      d_arr_22_1=>d_arr_22_1, d_arr_22_0=>d_arr_22_0, d_arr_23_31=>
      d_arr_23_31, d_arr_23_30=>d_arr_23_30, d_arr_23_29=>d_arr_23_29, 
      d_arr_23_28=>d_arr_23_28, d_arr_23_27=>d_arr_23_27, d_arr_23_26=>
      d_arr_23_26, d_arr_23_25=>d_arr_23_25, d_arr_23_24=>d_arr_23_24, 
      d_arr_23_23=>d_arr_23_23, d_arr_23_22=>d_arr_23_22, d_arr_23_21=>
      d_arr_23_21, d_arr_23_20=>d_arr_23_20, d_arr_23_19=>d_arr_23_19, 
      d_arr_23_18=>d_arr_23_18, d_arr_23_17=>d_arr_23_17, d_arr_23_16=>
      d_arr_23_16, d_arr_23_15=>d_arr_23_15, d_arr_23_14=>d_arr_23_14, 
      d_arr_23_13=>d_arr_23_13, d_arr_23_12=>d_arr_23_12, d_arr_23_11=>
      d_arr_23_11, d_arr_23_10=>d_arr_23_10, d_arr_23_9=>d_arr_23_9, 
      d_arr_23_8=>d_arr_23_8, d_arr_23_7=>d_arr_23_7, d_arr_23_6=>d_arr_23_6, 
      d_arr_23_5=>d_arr_23_5, d_arr_23_4=>d_arr_23_4, d_arr_23_3=>d_arr_23_3, 
      d_arr_23_2=>d_arr_23_2, d_arr_23_1=>d_arr_23_1, d_arr_23_0=>d_arr_23_0, 
      d_arr_24_31=>d_arr_24_31, d_arr_24_30=>d_arr_24_30, d_arr_24_29=>
      d_arr_24_29, d_arr_24_28=>d_arr_24_28, d_arr_24_27=>d_arr_24_27, 
      d_arr_24_26=>d_arr_24_26, d_arr_24_25=>d_arr_24_25, d_arr_24_24=>
      d_arr_24_24, d_arr_24_23=>d_arr_24_23, d_arr_24_22=>d_arr_24_22, 
      d_arr_24_21=>d_arr_24_21, d_arr_24_20=>d_arr_24_20, d_arr_24_19=>
      d_arr_24_19, d_arr_24_18=>d_arr_24_18, d_arr_24_17=>d_arr_24_17, 
      d_arr_24_16=>d_arr_24_16, d_arr_24_15=>d_arr_24_15, d_arr_24_14=>
      d_arr_24_14, d_arr_24_13=>d_arr_24_13, d_arr_24_12=>d_arr_24_12, 
      d_arr_24_11=>d_arr_24_11, d_arr_24_10=>d_arr_24_10, d_arr_24_9=>
      d_arr_24_9, d_arr_24_8=>d_arr_24_8, d_arr_24_7=>d_arr_24_7, d_arr_24_6
      =>d_arr_24_6, d_arr_24_5=>d_arr_24_5, d_arr_24_4=>d_arr_24_4, 
      d_arr_24_3=>d_arr_24_3, d_arr_24_2=>d_arr_24_2, d_arr_24_1=>d_arr_24_1, 
      d_arr_24_0=>d_arr_24_0);
   mux_layer_gen : MuxLayer port map ( img_data_0_31=>GND0, img_data_0_30=>
      GND0, img_data_0_29=>GND0, img_data_0_28=>GND0, img_data_0_27=>GND0, 
      img_data_0_26=>GND0, img_data_0_25=>GND0, img_data_0_24=>GND0, 
      img_data_0_23=>GND0, img_data_0_22=>GND0, img_data_0_21=>GND0, 
      img_data_0_20=>GND0, img_data_0_19=>GND0, img_data_0_18=>GND0, 
      img_data_0_17=>GND0, img_data_0_16=>GND0, img_data_0_15=>GND0, 
      img_data_0_14=>GND0, img_data_0_13=>GND0, img_data_0_12=>GND0, 
      img_data_0_11=>GND0, img_data_0_10=>GND0, img_data_0_9=>GND0, 
      img_data_0_8=>GND0, img_data_0_7=>GND0, img_data_0_6=>GND0, 
      img_data_0_5=>GND0, img_data_0_4=>GND0, img_data_0_3=>GND0, 
      img_data_0_2=>GND0, img_data_0_1=>GND0, img_data_0_0=>GND0, 
      img_data_1_31=>img_data_1_15, img_data_1_30=>GND0, img_data_1_29=>GND0, 
      img_data_1_28=>GND0, img_data_1_27=>GND0, img_data_1_26=>GND0, 
      img_data_1_25=>GND0, img_data_1_24=>GND0, img_data_1_23=>GND0, 
      img_data_1_22=>GND0, img_data_1_21=>GND0, img_data_1_20=>GND0, 
      img_data_1_19=>GND0, img_data_1_18=>GND0, img_data_1_17=>GND0, 
      img_data_1_16=>GND0, img_data_1_15=>GND0, img_data_1_14=>nx19398, 
      img_data_1_13=>img_data_1_13, img_data_1_12=>img_data_1_12, 
      img_data_1_11=>img_data_1_11, img_data_1_10=>nx19402, img_data_1_9=>
      img_data_1_9, img_data_1_8=>img_data_1_8, img_data_1_7=>img_data_1_7, 
      img_data_1_6=>img_data_1_6, img_data_1_5=>img_data_1_5, img_data_1_4=>
      img_data_1_4, img_data_1_3=>img_data_1_3, img_data_1_2=>img_data_1_2, 
      img_data_1_1=>img_data_1_1, img_data_1_0=>img_data_1_0, img_data_2_31
      =>img_data_2_15, img_data_2_30=>GND0, img_data_2_29=>GND0, 
      img_data_2_28=>GND0, img_data_2_27=>GND0, img_data_2_26=>GND0, 
      img_data_2_25=>GND0, img_data_2_24=>GND0, img_data_2_23=>GND0, 
      img_data_2_22=>GND0, img_data_2_21=>GND0, img_data_2_20=>GND0, 
      img_data_2_19=>GND0, img_data_2_18=>GND0, img_data_2_17=>GND0, 
      img_data_2_16=>GND0, img_data_2_15=>GND0, img_data_2_14=>nx19404, 
      img_data_2_13=>img_data_2_13, img_data_2_12=>img_data_2_12, 
      img_data_2_11=>img_data_2_11, img_data_2_10=>nx19408, img_data_2_9=>
      img_data_2_9, img_data_2_8=>img_data_2_8, img_data_2_7=>img_data_2_7, 
      img_data_2_6=>img_data_2_6, img_data_2_5=>img_data_2_5, img_data_2_4=>
      img_data_2_4, img_data_2_3=>img_data_2_3, img_data_2_2=>img_data_2_2, 
      img_data_2_1=>img_data_2_1, img_data_2_0=>img_data_2_0, img_data_3_31
      =>img_data_3_15, img_data_3_30=>GND0, img_data_3_29=>GND0, 
      img_data_3_28=>GND0, img_data_3_27=>GND0, img_data_3_26=>GND0, 
      img_data_3_25=>GND0, img_data_3_24=>GND0, img_data_3_23=>GND0, 
      img_data_3_22=>GND0, img_data_3_21=>GND0, img_data_3_20=>GND0, 
      img_data_3_19=>GND0, img_data_3_18=>GND0, img_data_3_17=>GND0, 
      img_data_3_16=>GND0, img_data_3_15=>GND0, img_data_3_14=>img_data_3_14, 
      img_data_3_13=>img_data_3_13, img_data_3_12=>img_data_3_12, 
      img_data_3_11=>img_data_3_11, img_data_3_10=>img_data_3_10, 
      img_data_3_9=>img_data_3_9, img_data_3_8=>img_data_3_8, img_data_3_7=>
      img_data_3_7, img_data_3_6=>img_data_3_6, img_data_3_5=>img_data_3_5, 
      img_data_3_4=>img_data_3_4, img_data_3_3=>img_data_3_3, img_data_3_2=>
      img_data_3_2, img_data_3_1=>img_data_3_1, img_data_3_0=>img_data_3_0, 
      img_data_4_31=>img_data_4_15, img_data_4_30=>GND0, img_data_4_29=>GND0, 
      img_data_4_28=>GND0, img_data_4_27=>GND0, img_data_4_26=>GND0, 
      img_data_4_25=>GND0, img_data_4_24=>GND0, img_data_4_23=>GND0, 
      img_data_4_22=>GND0, img_data_4_21=>GND0, img_data_4_20=>GND0, 
      img_data_4_19=>GND0, img_data_4_18=>GND0, img_data_4_17=>GND0, 
      img_data_4_16=>GND0, img_data_4_15=>GND0, img_data_4_14=>img_data_4_14, 
      img_data_4_13=>img_data_4_13, img_data_4_12=>img_data_4_12, 
      img_data_4_11=>img_data_4_11, img_data_4_10=>img_data_4_10, 
      img_data_4_9=>img_data_4_9, img_data_4_8=>img_data_4_8, img_data_4_7=>
      img_data_4_7, img_data_4_6=>img_data_4_6, img_data_4_5=>img_data_4_5, 
      img_data_4_4=>img_data_4_4, img_data_4_3=>img_data_4_3, img_data_4_2=>
      img_data_4_2, img_data_4_1=>img_data_4_1, img_data_4_0=>img_data_4_0, 
      img_data_5_31=>GND0, img_data_5_30=>GND0, img_data_5_29=>GND0, 
      img_data_5_28=>GND0, img_data_5_27=>GND0, img_data_5_26=>GND0, 
      img_data_5_25=>GND0, img_data_5_24=>GND0, img_data_5_23=>GND0, 
      img_data_5_22=>GND0, img_data_5_21=>GND0, img_data_5_20=>GND0, 
      img_data_5_19=>GND0, img_data_5_18=>GND0, img_data_5_17=>GND0, 
      img_data_5_16=>GND0, img_data_5_15=>GND0, img_data_5_14=>GND0, 
      img_data_5_13=>GND0, img_data_5_12=>GND0, img_data_5_11=>GND0, 
      img_data_5_10=>GND0, img_data_5_9=>GND0, img_data_5_8=>GND0, 
      img_data_5_7=>GND0, img_data_5_6=>GND0, img_data_5_5=>GND0, 
      img_data_5_4=>GND0, img_data_5_3=>GND0, img_data_5_2=>GND0, 
      img_data_5_1=>GND0, img_data_5_0=>GND0, img_data_6_31=>img_data_6_15, 
      img_data_6_30=>GND0, img_data_6_29=>GND0, img_data_6_28=>GND0, 
      img_data_6_27=>GND0, img_data_6_26=>GND0, img_data_6_25=>GND0, 
      img_data_6_24=>GND0, img_data_6_23=>GND0, img_data_6_22=>GND0, 
      img_data_6_21=>GND0, img_data_6_20=>GND0, img_data_6_19=>GND0, 
      img_data_6_18=>GND0, img_data_6_17=>GND0, img_data_6_16=>GND0, 
      img_data_6_15=>GND0, img_data_6_14=>nx19412, img_data_6_13=>
      img_data_6_13, img_data_6_12=>img_data_6_12, img_data_6_11=>
      img_data_6_11, img_data_6_10=>nx19416, img_data_6_9=>img_data_6_9, 
      img_data_6_8=>img_data_6_8, img_data_6_7=>img_data_6_7, img_data_6_6=>
      img_data_6_6, img_data_6_5=>img_data_6_5, img_data_6_4=>img_data_6_4, 
      img_data_6_3=>img_data_6_3, img_data_6_2=>img_data_6_2, img_data_6_1=>
      img_data_6_1, img_data_6_0=>img_data_6_0, img_data_7_31=>nx16659, 
      img_data_7_30=>GND0, img_data_7_29=>GND0, img_data_7_28=>GND0, 
      img_data_7_27=>GND0, img_data_7_26=>GND0, img_data_7_25=>GND0, 
      img_data_7_24=>GND0, img_data_7_23=>GND0, img_data_7_22=>GND0, 
      img_data_7_21=>GND0, img_data_7_20=>GND0, img_data_7_19=>GND0, 
      img_data_7_18=>GND0, img_data_7_17=>GND0, img_data_7_16=>GND0, 
      img_data_7_15=>GND0, img_data_7_14=>nx19418, img_data_7_13=>
      img_data_7_13, img_data_7_12=>img_data_7_12, img_data_7_11=>
      img_data_7_11, img_data_7_10=>nx19422, img_data_7_9=>img_data_7_9, 
      img_data_7_8=>img_data_7_8, img_data_7_7=>img_data_7_7, img_data_7_6=>
      img_data_7_6, img_data_7_5=>img_data_7_5, img_data_7_4=>img_data_7_4, 
      img_data_7_3=>img_data_7_3, img_data_7_2=>img_data_7_2, img_data_7_1=>
      img_data_7_1, img_data_7_0=>img_data_7_0, img_data_8_31=>img_data_8_15, 
      img_data_8_30=>GND0, img_data_8_29=>GND0, img_data_8_28=>GND0, 
      img_data_8_27=>GND0, img_data_8_26=>GND0, img_data_8_25=>GND0, 
      img_data_8_24=>GND0, img_data_8_23=>GND0, img_data_8_22=>GND0, 
      img_data_8_21=>GND0, img_data_8_20=>GND0, img_data_8_19=>GND0, 
      img_data_8_18=>GND0, img_data_8_17=>GND0, img_data_8_16=>GND0, 
      img_data_8_15=>GND0, img_data_8_14=>img_data_8_14, img_data_8_13=>
      img_data_8_13, img_data_8_12=>img_data_8_12, img_data_8_11=>
      img_data_8_11, img_data_8_10=>img_data_8_10, img_data_8_9=>
      img_data_8_9, img_data_8_8=>img_data_8_8, img_data_8_7=>img_data_8_7, 
      img_data_8_6=>img_data_8_6, img_data_8_5=>img_data_8_5, img_data_8_4=>
      img_data_8_4, img_data_8_3=>img_data_8_3, img_data_8_2=>img_data_8_2, 
      img_data_8_1=>img_data_8_1, img_data_8_0=>img_data_8_0, img_data_9_31
      =>img_data_9_15, img_data_9_30=>GND0, img_data_9_29=>GND0, 
      img_data_9_28=>GND0, img_data_9_27=>GND0, img_data_9_26=>GND0, 
      img_data_9_25=>GND0, img_data_9_24=>GND0, img_data_9_23=>GND0, 
      img_data_9_22=>GND0, img_data_9_21=>GND0, img_data_9_20=>GND0, 
      img_data_9_19=>GND0, img_data_9_18=>GND0, img_data_9_17=>GND0, 
      img_data_9_16=>GND0, img_data_9_15=>GND0, img_data_9_14=>img_data_9_14, 
      img_data_9_13=>img_data_9_13, img_data_9_12=>img_data_9_12, 
      img_data_9_11=>img_data_9_11, img_data_9_10=>img_data_9_10, 
      img_data_9_9=>img_data_9_9, img_data_9_8=>img_data_9_8, img_data_9_7=>
      img_data_9_7, img_data_9_6=>img_data_9_6, img_data_9_5=>img_data_9_5, 
      img_data_9_4=>img_data_9_4, img_data_9_3=>img_data_9_3, img_data_9_2=>
      img_data_9_2, img_data_9_1=>img_data_9_1, img_data_9_0=>img_data_9_0, 
      img_data_10_31=>GND0, img_data_10_30=>GND0, img_data_10_29=>GND0, 
      img_data_10_28=>GND0, img_data_10_27=>GND0, img_data_10_26=>GND0, 
      img_data_10_25=>GND0, img_data_10_24=>GND0, img_data_10_23=>GND0, 
      img_data_10_22=>GND0, img_data_10_21=>GND0, img_data_10_20=>GND0, 
      img_data_10_19=>GND0, img_data_10_18=>GND0, img_data_10_17=>GND0, 
      img_data_10_16=>GND0, img_data_10_15=>GND0, img_data_10_14=>GND0, 
      img_data_10_13=>GND0, img_data_10_12=>GND0, img_data_10_11=>GND0, 
      img_data_10_10=>GND0, img_data_10_9=>GND0, img_data_10_8=>GND0, 
      img_data_10_7=>GND0, img_data_10_6=>GND0, img_data_10_5=>GND0, 
      img_data_10_4=>GND0, img_data_10_3=>GND0, img_data_10_2=>GND0, 
      img_data_10_1=>GND0, img_data_10_0=>GND0, img_data_11_31=>nx16661, 
      img_data_11_30=>GND0, img_data_11_29=>GND0, img_data_11_28=>GND0, 
      img_data_11_27=>GND0, img_data_11_26=>GND0, img_data_11_25=>GND0, 
      img_data_11_24=>GND0, img_data_11_23=>GND0, img_data_11_22=>GND0, 
      img_data_11_21=>GND0, img_data_11_20=>GND0, img_data_11_19=>GND0, 
      img_data_11_18=>GND0, img_data_11_17=>GND0, img_data_11_16=>GND0, 
      img_data_11_15=>GND0, img_data_11_14=>nx19426, img_data_11_13=>
      img_data_11_13, img_data_11_12=>img_data_11_12, img_data_11_11=>
      img_data_11_11, img_data_11_10=>nx19430, img_data_11_9=>img_data_11_9, 
      img_data_11_8=>img_data_11_8, img_data_11_7=>img_data_11_7, 
      img_data_11_6=>img_data_11_6, img_data_11_5=>img_data_11_5, 
      img_data_11_4=>img_data_11_4, img_data_11_3=>img_data_11_3, 
      img_data_11_2=>img_data_11_2, img_data_11_1=>img_data_11_1, 
      img_data_11_0=>img_data_11_0, img_data_12_31=>nx16663, img_data_12_30
      =>GND0, img_data_12_29=>GND0, img_data_12_28=>GND0, img_data_12_27=>
      GND0, img_data_12_26=>GND0, img_data_12_25=>GND0, img_data_12_24=>GND0, 
      img_data_12_23=>GND0, img_data_12_22=>GND0, img_data_12_21=>GND0, 
      img_data_12_20=>GND0, img_data_12_19=>GND0, img_data_12_18=>GND0, 
      img_data_12_17=>GND0, img_data_12_16=>GND0, img_data_12_15=>GND0, 
      img_data_12_14=>nx19432, img_data_12_13=>img_data_12_13, 
      img_data_12_12=>img_data_12_12, img_data_12_11=>img_data_12_11, 
      img_data_12_10=>nx19436, img_data_12_9=>img_data_12_9, img_data_12_8=>
      img_data_12_8, img_data_12_7=>img_data_12_7, img_data_12_6=>
      img_data_12_6, img_data_12_5=>img_data_12_5, img_data_12_4=>
      img_data_12_4, img_data_12_3=>img_data_12_3, img_data_12_2=>
      img_data_12_2, img_data_12_1=>img_data_12_1, img_data_12_0=>
      img_data_12_0, img_data_13_31=>img_data_13_15, img_data_13_30=>GND0, 
      img_data_13_29=>GND0, img_data_13_28=>GND0, img_data_13_27=>GND0, 
      img_data_13_26=>GND0, img_data_13_25=>GND0, img_data_13_24=>GND0, 
      img_data_13_23=>GND0, img_data_13_22=>GND0, img_data_13_21=>GND0, 
      img_data_13_20=>GND0, img_data_13_19=>GND0, img_data_13_18=>GND0, 
      img_data_13_17=>GND0, img_data_13_16=>GND0, img_data_13_15=>GND0, 
      img_data_13_14=>img_data_13_14, img_data_13_13=>img_data_13_13, 
      img_data_13_12=>img_data_13_12, img_data_13_11=>img_data_13_11, 
      img_data_13_10=>img_data_13_10, img_data_13_9=>img_data_13_9, 
      img_data_13_8=>img_data_13_8, img_data_13_7=>img_data_13_7, 
      img_data_13_6=>img_data_13_6, img_data_13_5=>img_data_13_5, 
      img_data_13_4=>img_data_13_4, img_data_13_3=>img_data_13_3, 
      img_data_13_2=>img_data_13_2, img_data_13_1=>img_data_13_1, 
      img_data_13_0=>img_data_13_0, img_data_14_31=>img_data_14_15, 
      img_data_14_30=>GND0, img_data_14_29=>GND0, img_data_14_28=>GND0, 
      img_data_14_27=>GND0, img_data_14_26=>GND0, img_data_14_25=>GND0, 
      img_data_14_24=>GND0, img_data_14_23=>GND0, img_data_14_22=>GND0, 
      img_data_14_21=>GND0, img_data_14_20=>GND0, img_data_14_19=>GND0, 
      img_data_14_18=>GND0, img_data_14_17=>GND0, img_data_14_16=>GND0, 
      img_data_14_15=>GND0, img_data_14_14=>img_data_14_14, img_data_14_13=>
      img_data_14_13, img_data_14_12=>img_data_14_12, img_data_14_11=>
      img_data_14_11, img_data_14_10=>img_data_14_10, img_data_14_9=>
      img_data_14_9, img_data_14_8=>img_data_14_8, img_data_14_7=>
      img_data_14_7, img_data_14_6=>img_data_14_6, img_data_14_5=>
      img_data_14_5, img_data_14_4=>img_data_14_4, img_data_14_3=>
      img_data_14_3, img_data_14_2=>img_data_14_2, img_data_14_1=>
      img_data_14_1, img_data_14_0=>img_data_14_0, img_data_15_31=>
      img_data_15_15, img_data_15_30=>GND0, img_data_15_29=>GND0, 
      img_data_15_28=>GND0, img_data_15_27=>GND0, img_data_15_26=>GND0, 
      img_data_15_25=>GND0, img_data_15_24=>GND0, img_data_15_23=>GND0, 
      img_data_15_22=>GND0, img_data_15_21=>GND0, img_data_15_20=>GND0, 
      img_data_15_19=>GND0, img_data_15_18=>GND0, img_data_15_17=>GND0, 
      img_data_15_16=>GND0, img_data_15_15=>GND0, img_data_15_14=>
      img_data_15_14, img_data_15_13=>img_data_15_13, img_data_15_12=>
      img_data_15_12, img_data_15_11=>img_data_15_11, img_data_15_10=>
      img_data_15_10, img_data_15_9=>img_data_15_9, img_data_15_8=>
      img_data_15_8, img_data_15_7=>img_data_15_7, img_data_15_6=>
      img_data_15_6, img_data_15_5=>img_data_15_5, img_data_15_4=>
      img_data_15_4, img_data_15_3=>img_data_15_3, img_data_15_2=>
      img_data_15_2, img_data_15_1=>img_data_15_1, img_data_15_0=>
      img_data_15_0, img_data_16_31=>img_data_16_15, img_data_16_30=>GND0, 
      img_data_16_29=>GND0, img_data_16_28=>GND0, img_data_16_27=>GND0, 
      img_data_16_26=>GND0, img_data_16_25=>GND0, img_data_16_24=>GND0, 
      img_data_16_23=>GND0, img_data_16_22=>GND0, img_data_16_21=>GND0, 
      img_data_16_20=>GND0, img_data_16_19=>GND0, img_data_16_18=>GND0, 
      img_data_16_17=>GND0, img_data_16_16=>GND0, img_data_16_15=>GND0, 
      img_data_16_14=>img_data_16_14, img_data_16_13=>img_data_16_13, 
      img_data_16_12=>img_data_16_12, img_data_16_11=>img_data_16_11, 
      img_data_16_10=>img_data_16_10, img_data_16_9=>img_data_16_9, 
      img_data_16_8=>img_data_16_8, img_data_16_7=>img_data_16_7, 
      img_data_16_6=>img_data_16_6, img_data_16_5=>img_data_16_5, 
      img_data_16_4=>img_data_16_4, img_data_16_3=>img_data_16_3, 
      img_data_16_2=>img_data_16_2, img_data_16_1=>img_data_16_1, 
      img_data_16_0=>img_data_16_0, img_data_17_31=>img_data_17_15, 
      img_data_17_30=>GND0, img_data_17_29=>GND0, img_data_17_28=>GND0, 
      img_data_17_27=>GND0, img_data_17_26=>GND0, img_data_17_25=>GND0, 
      img_data_17_24=>GND0, img_data_17_23=>GND0, img_data_17_22=>GND0, 
      img_data_17_21=>GND0, img_data_17_20=>GND0, img_data_17_19=>GND0, 
      img_data_17_18=>GND0, img_data_17_17=>GND0, img_data_17_16=>GND0, 
      img_data_17_15=>GND0, img_data_17_14=>img_data_17_14, img_data_17_13=>
      img_data_17_13, img_data_17_12=>img_data_17_12, img_data_17_11=>
      img_data_17_11, img_data_17_10=>img_data_17_10, img_data_17_9=>
      img_data_17_9, img_data_17_8=>img_data_17_8, img_data_17_7=>
      img_data_17_7, img_data_17_6=>img_data_17_6, img_data_17_5=>
      img_data_17_5, img_data_17_4=>img_data_17_4, img_data_17_3=>
      img_data_17_3, img_data_17_2=>img_data_17_2, img_data_17_1=>
      img_data_17_1, img_data_17_0=>img_data_17_0, img_data_18_31=>GND0, 
      img_data_18_30=>GND0, img_data_18_29=>GND0, img_data_18_28=>GND0, 
      img_data_18_27=>GND0, img_data_18_26=>GND0, img_data_18_25=>GND0, 
      img_data_18_24=>GND0, img_data_18_23=>GND0, img_data_18_22=>GND0, 
      img_data_18_21=>GND0, img_data_18_20=>GND0, img_data_18_19=>GND0, 
      img_data_18_18=>GND0, img_data_18_17=>GND0, img_data_18_16=>GND0, 
      img_data_18_15=>GND0, img_data_18_14=>GND0, img_data_18_13=>GND0, 
      img_data_18_12=>GND0, img_data_18_11=>GND0, img_data_18_10=>GND0, 
      img_data_18_9=>GND0, img_data_18_8=>GND0, img_data_18_7=>GND0, 
      img_data_18_6=>GND0, img_data_18_5=>GND0, img_data_18_4=>GND0, 
      img_data_18_3=>GND0, img_data_18_2=>GND0, img_data_18_1=>GND0, 
      img_data_18_0=>GND0, img_data_19_31=>GND0, img_data_19_30=>GND0, 
      img_data_19_29=>GND0, img_data_19_28=>GND0, img_data_19_27=>GND0, 
      img_data_19_26=>GND0, img_data_19_25=>GND0, img_data_19_24=>GND0, 
      img_data_19_23=>GND0, img_data_19_22=>GND0, img_data_19_21=>GND0, 
      img_data_19_20=>GND0, img_data_19_19=>GND0, img_data_19_18=>GND0, 
      img_data_19_17=>GND0, img_data_19_16=>GND0, img_data_19_15=>GND0, 
      img_data_19_14=>GND0, img_data_19_13=>GND0, img_data_19_12=>GND0, 
      img_data_19_11=>GND0, img_data_19_10=>GND0, img_data_19_9=>GND0, 
      img_data_19_8=>GND0, img_data_19_7=>GND0, img_data_19_6=>GND0, 
      img_data_19_5=>GND0, img_data_19_4=>GND0, img_data_19_3=>GND0, 
      img_data_19_2=>GND0, img_data_19_1=>GND0, img_data_19_0=>GND0, 
      img_data_20_31=>GND0, img_data_20_30=>GND0, img_data_20_29=>GND0, 
      img_data_20_28=>GND0, img_data_20_27=>GND0, img_data_20_26=>GND0, 
      img_data_20_25=>GND0, img_data_20_24=>GND0, img_data_20_23=>GND0, 
      img_data_20_22=>GND0, img_data_20_21=>GND0, img_data_20_20=>GND0, 
      img_data_20_19=>GND0, img_data_20_18=>GND0, img_data_20_17=>GND0, 
      img_data_20_16=>GND0, img_data_20_15=>GND0, img_data_20_14=>GND0, 
      img_data_20_13=>GND0, img_data_20_12=>GND0, img_data_20_11=>GND0, 
      img_data_20_10=>GND0, img_data_20_9=>GND0, img_data_20_8=>GND0, 
      img_data_20_7=>GND0, img_data_20_6=>GND0, img_data_20_5=>GND0, 
      img_data_20_4=>GND0, img_data_20_3=>GND0, img_data_20_2=>GND0, 
      img_data_20_1=>GND0, img_data_20_0=>GND0, img_data_21_31=>GND0, 
      img_data_21_30=>GND0, img_data_21_29=>GND0, img_data_21_28=>GND0, 
      img_data_21_27=>GND0, img_data_21_26=>GND0, img_data_21_25=>GND0, 
      img_data_21_24=>GND0, img_data_21_23=>GND0, img_data_21_22=>GND0, 
      img_data_21_21=>GND0, img_data_21_20=>GND0, img_data_21_19=>GND0, 
      img_data_21_18=>GND0, img_data_21_17=>GND0, img_data_21_16=>GND0, 
      img_data_21_15=>GND0, img_data_21_14=>GND0, img_data_21_13=>GND0, 
      img_data_21_12=>GND0, img_data_21_11=>GND0, img_data_21_10=>GND0, 
      img_data_21_9=>GND0, img_data_21_8=>GND0, img_data_21_7=>GND0, 
      img_data_21_6=>GND0, img_data_21_5=>GND0, img_data_21_4=>GND0, 
      img_data_21_3=>GND0, img_data_21_2=>GND0, img_data_21_1=>GND0, 
      img_data_21_0=>GND0, img_data_22_31=>GND0, img_data_22_30=>GND0, 
      img_data_22_29=>GND0, img_data_22_28=>GND0, img_data_22_27=>GND0, 
      img_data_22_26=>GND0, img_data_22_25=>GND0, img_data_22_24=>GND0, 
      img_data_22_23=>GND0, img_data_22_22=>GND0, img_data_22_21=>GND0, 
      img_data_22_20=>GND0, img_data_22_19=>GND0, img_data_22_18=>GND0, 
      img_data_22_17=>GND0, img_data_22_16=>GND0, img_data_22_15=>GND0, 
      img_data_22_14=>GND0, img_data_22_13=>GND0, img_data_22_12=>GND0, 
      img_data_22_11=>GND0, img_data_22_10=>GND0, img_data_22_9=>GND0, 
      img_data_22_8=>GND0, img_data_22_7=>GND0, img_data_22_6=>GND0, 
      img_data_22_5=>GND0, img_data_22_4=>GND0, img_data_22_3=>GND0, 
      img_data_22_2=>GND0, img_data_22_1=>GND0, img_data_22_0=>GND0, 
      img_data_23_31=>GND0, img_data_23_30=>GND0, img_data_23_29=>GND0, 
      img_data_23_28=>GND0, img_data_23_27=>GND0, img_data_23_26=>GND0, 
      img_data_23_25=>GND0, img_data_23_24=>GND0, img_data_23_23=>GND0, 
      img_data_23_22=>GND0, img_data_23_21=>GND0, img_data_23_20=>GND0, 
      img_data_23_19=>GND0, img_data_23_18=>GND0, img_data_23_17=>GND0, 
      img_data_23_16=>GND0, img_data_23_15=>GND0, img_data_23_14=>GND0, 
      img_data_23_13=>GND0, img_data_23_12=>GND0, img_data_23_11=>GND0, 
      img_data_23_10=>GND0, img_data_23_9=>GND0, img_data_23_8=>GND0, 
      img_data_23_7=>GND0, img_data_23_6=>GND0, img_data_23_5=>GND0, 
      img_data_23_4=>GND0, img_data_23_3=>GND0, img_data_23_2=>GND0, 
      img_data_23_1=>GND0, img_data_23_0=>GND0, img_data_24_31=>GND0, 
      img_data_24_30=>GND0, img_data_24_29=>GND0, img_data_24_28=>GND0, 
      img_data_24_27=>GND0, img_data_24_26=>GND0, img_data_24_25=>GND0, 
      img_data_24_24=>GND0, img_data_24_23=>GND0, img_data_24_22=>GND0, 
      img_data_24_21=>GND0, img_data_24_20=>GND0, img_data_24_19=>GND0, 
      img_data_24_18=>GND0, img_data_24_17=>GND0, img_data_24_16=>GND0, 
      img_data_24_15=>GND0, img_data_24_14=>GND0, img_data_24_13=>GND0, 
      img_data_24_12=>GND0, img_data_24_11=>GND0, img_data_24_10=>GND0, 
      img_data_24_9=>GND0, img_data_24_8=>GND0, img_data_24_7=>GND0, 
      img_data_24_6=>GND0, img_data_24_5=>GND0, img_data_24_4=>GND0, 
      img_data_24_3=>GND0, img_data_24_2=>GND0, img_data_24_1=>GND0, 
      img_data_24_0=>GND0, filter_data_0_31=>filter_data_0_15, 
      filter_data_0_30=>GND0, filter_data_0_29=>GND0, filter_data_0_28=>GND0, 
      filter_data_0_27=>GND0, filter_data_0_26=>GND0, filter_data_0_25=>GND0, 
      filter_data_0_24=>GND0, filter_data_0_23=>GND0, filter_data_0_22=>GND0, 
      filter_data_0_21=>GND0, filter_data_0_20=>GND0, filter_data_0_19=>GND0, 
      filter_data_0_18=>GND0, filter_data_0_17=>GND0, filter_data_0_16=>GND0, 
      filter_data_0_15=>GND0, filter_data_0_14=>filter_data_0_14, 
      filter_data_0_13=>filter_data_0_13, filter_data_0_12=>filter_data_0_12, 
      filter_data_0_11=>filter_data_0_11, filter_data_0_10=>filter_data_0_10, 
      filter_data_0_9=>filter_data_0_9, filter_data_0_8=>filter_data_0_8, 
      filter_data_0_7=>filter_data_0_7, filter_data_0_6=>filter_data_0_6, 
      filter_data_0_5=>filter_data_0_5, filter_data_0_4=>filter_data_0_4, 
      filter_data_0_3=>filter_data_0_3, filter_data_0_2=>filter_data_0_2, 
      filter_data_0_1=>filter_data_0_1, filter_data_0_0=>filter_data_0_0, 
      filter_data_1_31=>filter_data_1_15, filter_data_1_30=>GND0, 
      filter_data_1_29=>GND0, filter_data_1_28=>GND0, filter_data_1_27=>GND0, 
      filter_data_1_26=>GND0, filter_data_1_25=>GND0, filter_data_1_24=>GND0, 
      filter_data_1_23=>GND0, filter_data_1_22=>GND0, filter_data_1_21=>GND0, 
      filter_data_1_20=>GND0, filter_data_1_19=>GND0, filter_data_1_18=>GND0, 
      filter_data_1_17=>GND0, filter_data_1_16=>GND0, filter_data_1_15=>GND0, 
      filter_data_1_14=>filter_data_1_14, filter_data_1_13=>filter_data_1_13, 
      filter_data_1_12=>filter_data_1_12, filter_data_1_11=>filter_data_1_11, 
      filter_data_1_10=>filter_data_1_10, filter_data_1_9=>filter_data_1_9, 
      filter_data_1_8=>filter_data_1_8, filter_data_1_7=>filter_data_1_7, 
      filter_data_1_6=>filter_data_1_6, filter_data_1_5=>filter_data_1_5, 
      filter_data_1_4=>filter_data_1_4, filter_data_1_3=>filter_data_1_3, 
      filter_data_1_2=>filter_data_1_2, filter_data_1_1=>filter_data_1_1, 
      filter_data_1_0=>filter_data_1_0, filter_data_2_31=>filter_data_2_15, 
      filter_data_2_30=>GND0, filter_data_2_29=>GND0, filter_data_2_28=>GND0, 
      filter_data_2_27=>GND0, filter_data_2_26=>GND0, filter_data_2_25=>GND0, 
      filter_data_2_24=>GND0, filter_data_2_23=>GND0, filter_data_2_22=>GND0, 
      filter_data_2_21=>GND0, filter_data_2_20=>GND0, filter_data_2_19=>GND0, 
      filter_data_2_18=>GND0, filter_data_2_17=>GND0, filter_data_2_16=>GND0, 
      filter_data_2_15=>GND0, filter_data_2_14=>filter_data_2_14, 
      filter_data_2_13=>filter_data_2_13, filter_data_2_12=>filter_data_2_12, 
      filter_data_2_11=>filter_data_2_11, filter_data_2_10=>filter_data_2_10, 
      filter_data_2_9=>filter_data_2_9, filter_data_2_8=>filter_data_2_8, 
      filter_data_2_7=>filter_data_2_7, filter_data_2_6=>filter_data_2_6, 
      filter_data_2_5=>filter_data_2_5, filter_data_2_4=>filter_data_2_4, 
      filter_data_2_3=>filter_data_2_3, filter_data_2_2=>filter_data_2_2, 
      filter_data_2_1=>filter_data_2_1, filter_data_2_0=>filter_data_2_0, 
      filter_data_3_31=>filter_data_3_15, filter_data_3_30=>GND0, 
      filter_data_3_29=>GND0, filter_data_3_28=>GND0, filter_data_3_27=>GND0, 
      filter_data_3_26=>GND0, filter_data_3_25=>GND0, filter_data_3_24=>GND0, 
      filter_data_3_23=>GND0, filter_data_3_22=>GND0, filter_data_3_21=>GND0, 
      filter_data_3_20=>GND0, filter_data_3_19=>GND0, filter_data_3_18=>GND0, 
      filter_data_3_17=>GND0, filter_data_3_16=>GND0, filter_data_3_15=>GND0, 
      filter_data_3_14=>filter_data_3_14, filter_data_3_13=>filter_data_3_13, 
      filter_data_3_12=>filter_data_3_12, filter_data_3_11=>filter_data_3_11, 
      filter_data_3_10=>filter_data_3_10, filter_data_3_9=>filter_data_3_9, 
      filter_data_3_8=>filter_data_3_8, filter_data_3_7=>filter_data_3_7, 
      filter_data_3_6=>filter_data_3_6, filter_data_3_5=>filter_data_3_5, 
      filter_data_3_4=>filter_data_3_4, filter_data_3_3=>filter_data_3_3, 
      filter_data_3_2=>filter_data_3_2, filter_data_3_1=>filter_data_3_1, 
      filter_data_3_0=>filter_data_3_0, filter_data_4_31=>filter_data_4_15, 
      filter_data_4_30=>GND0, filter_data_4_29=>GND0, filter_data_4_28=>GND0, 
      filter_data_4_27=>GND0, filter_data_4_26=>GND0, filter_data_4_25=>GND0, 
      filter_data_4_24=>GND0, filter_data_4_23=>GND0, filter_data_4_22=>GND0, 
      filter_data_4_21=>GND0, filter_data_4_20=>GND0, filter_data_4_19=>GND0, 
      filter_data_4_18=>GND0, filter_data_4_17=>GND0, filter_data_4_16=>GND0, 
      filter_data_4_15=>GND0, filter_data_4_14=>filter_data_4_14, 
      filter_data_4_13=>filter_data_4_13, filter_data_4_12=>filter_data_4_12, 
      filter_data_4_11=>filter_data_4_11, filter_data_4_10=>filter_data_4_10, 
      filter_data_4_9=>filter_data_4_9, filter_data_4_8=>filter_data_4_8, 
      filter_data_4_7=>filter_data_4_7, filter_data_4_6=>filter_data_4_6, 
      filter_data_4_5=>filter_data_4_5, filter_data_4_4=>filter_data_4_4, 
      filter_data_4_3=>filter_data_4_3, filter_data_4_2=>filter_data_4_2, 
      filter_data_4_1=>filter_data_4_1, filter_data_4_0=>filter_data_4_0, 
      filter_data_5_31=>filter_data_5_15, filter_data_5_30=>GND0, 
      filter_data_5_29=>GND0, filter_data_5_28=>GND0, filter_data_5_27=>GND0, 
      filter_data_5_26=>GND0, filter_data_5_25=>GND0, filter_data_5_24=>GND0, 
      filter_data_5_23=>GND0, filter_data_5_22=>GND0, filter_data_5_21=>GND0, 
      filter_data_5_20=>GND0, filter_data_5_19=>GND0, filter_data_5_18=>GND0, 
      filter_data_5_17=>GND0, filter_data_5_16=>GND0, filter_data_5_15=>GND0, 
      filter_data_5_14=>filter_data_5_14, filter_data_5_13=>filter_data_5_13, 
      filter_data_5_12=>filter_data_5_12, filter_data_5_11=>filter_data_5_11, 
      filter_data_5_10=>filter_data_5_10, filter_data_5_9=>filter_data_5_9, 
      filter_data_5_8=>filter_data_5_8, filter_data_5_7=>filter_data_5_7, 
      filter_data_5_6=>filter_data_5_6, filter_data_5_5=>filter_data_5_5, 
      filter_data_5_4=>filter_data_5_4, filter_data_5_3=>filter_data_5_3, 
      filter_data_5_2=>filter_data_5_2, filter_data_5_1=>filter_data_5_1, 
      filter_data_5_0=>filter_data_5_0, filter_data_6_31=>filter_data_6_15, 
      filter_data_6_30=>GND0, filter_data_6_29=>GND0, filter_data_6_28=>GND0, 
      filter_data_6_27=>GND0, filter_data_6_26=>GND0, filter_data_6_25=>GND0, 
      filter_data_6_24=>GND0, filter_data_6_23=>GND0, filter_data_6_22=>GND0, 
      filter_data_6_21=>GND0, filter_data_6_20=>GND0, filter_data_6_19=>GND0, 
      filter_data_6_18=>GND0, filter_data_6_17=>GND0, filter_data_6_16=>GND0, 
      filter_data_6_15=>GND0, filter_data_6_14=>filter_data_6_14, 
      filter_data_6_13=>filter_data_6_13, filter_data_6_12=>filter_data_6_12, 
      filter_data_6_11=>filter_data_6_11, filter_data_6_10=>filter_data_6_10, 
      filter_data_6_9=>filter_data_6_9, filter_data_6_8=>filter_data_6_8, 
      filter_data_6_7=>filter_data_6_7, filter_data_6_6=>filter_data_6_6, 
      filter_data_6_5=>filter_data_6_5, filter_data_6_4=>filter_data_6_4, 
      filter_data_6_3=>filter_data_6_3, filter_data_6_2=>filter_data_6_2, 
      filter_data_6_1=>filter_data_6_1, filter_data_6_0=>filter_data_6_0, 
      filter_data_7_31=>filter_data_7_15, filter_data_7_30=>GND0, 
      filter_data_7_29=>GND0, filter_data_7_28=>GND0, filter_data_7_27=>GND0, 
      filter_data_7_26=>GND0, filter_data_7_25=>GND0, filter_data_7_24=>GND0, 
      filter_data_7_23=>GND0, filter_data_7_22=>GND0, filter_data_7_21=>GND0, 
      filter_data_7_20=>GND0, filter_data_7_19=>GND0, filter_data_7_18=>GND0, 
      filter_data_7_17=>GND0, filter_data_7_16=>GND0, filter_data_7_15=>GND0, 
      filter_data_7_14=>filter_data_7_14, filter_data_7_13=>filter_data_7_13, 
      filter_data_7_12=>filter_data_7_12, filter_data_7_11=>filter_data_7_11, 
      filter_data_7_10=>filter_data_7_10, filter_data_7_9=>filter_data_7_9, 
      filter_data_7_8=>filter_data_7_8, filter_data_7_7=>filter_data_7_7, 
      filter_data_7_6=>filter_data_7_6, filter_data_7_5=>filter_data_7_5, 
      filter_data_7_4=>filter_data_7_4, filter_data_7_3=>filter_data_7_3, 
      filter_data_7_2=>filter_data_7_2, filter_data_7_1=>filter_data_7_1, 
      filter_data_7_0=>filter_data_7_0, filter_data_8_31=>filter_data_8_15, 
      filter_data_8_30=>GND0, filter_data_8_29=>GND0, filter_data_8_28=>GND0, 
      filter_data_8_27=>GND0, filter_data_8_26=>GND0, filter_data_8_25=>GND0, 
      filter_data_8_24=>GND0, filter_data_8_23=>GND0, filter_data_8_22=>GND0, 
      filter_data_8_21=>GND0, filter_data_8_20=>GND0, filter_data_8_19=>GND0, 
      filter_data_8_18=>GND0, filter_data_8_17=>GND0, filter_data_8_16=>GND0, 
      filter_data_8_15=>GND0, filter_data_8_14=>filter_data_8_14, 
      filter_data_8_13=>filter_data_8_13, filter_data_8_12=>filter_data_8_12, 
      filter_data_8_11=>filter_data_8_11, filter_data_8_10=>filter_data_8_10, 
      filter_data_8_9=>filter_data_8_9, filter_data_8_8=>filter_data_8_8, 
      filter_data_8_7=>filter_data_8_7, filter_data_8_6=>filter_data_8_6, 
      filter_data_8_5=>filter_data_8_5, filter_data_8_4=>filter_data_8_4, 
      filter_data_8_3=>filter_data_8_3, filter_data_8_2=>filter_data_8_2, 
      filter_data_8_1=>filter_data_8_1, filter_data_8_0=>filter_data_8_0, 
      filter_data_9_31=>filter_data_9_15, filter_data_9_30=>GND0, 
      filter_data_9_29=>GND0, filter_data_9_28=>GND0, filter_data_9_27=>GND0, 
      filter_data_9_26=>GND0, filter_data_9_25=>GND0, filter_data_9_24=>GND0, 
      filter_data_9_23=>GND0, filter_data_9_22=>GND0, filter_data_9_21=>GND0, 
      filter_data_9_20=>GND0, filter_data_9_19=>GND0, filter_data_9_18=>GND0, 
      filter_data_9_17=>GND0, filter_data_9_16=>GND0, filter_data_9_15=>GND0, 
      filter_data_9_14=>filter_data_9_14, filter_data_9_13=>filter_data_9_13, 
      filter_data_9_12=>filter_data_9_12, filter_data_9_11=>filter_data_9_11, 
      filter_data_9_10=>filter_data_9_10, filter_data_9_9=>filter_data_9_9, 
      filter_data_9_8=>filter_data_9_8, filter_data_9_7=>filter_data_9_7, 
      filter_data_9_6=>filter_data_9_6, filter_data_9_5=>filter_data_9_5, 
      filter_data_9_4=>filter_data_9_4, filter_data_9_3=>filter_data_9_3, 
      filter_data_9_2=>filter_data_9_2, filter_data_9_1=>filter_data_9_1, 
      filter_data_9_0=>filter_data_9_0, filter_data_10_31=>filter_data_10_15, 
      filter_data_10_30=>GND0, filter_data_10_29=>GND0, filter_data_10_28=>
      GND0, filter_data_10_27=>GND0, filter_data_10_26=>GND0, 
      filter_data_10_25=>GND0, filter_data_10_24=>GND0, filter_data_10_23=>
      GND0, filter_data_10_22=>GND0, filter_data_10_21=>GND0, 
      filter_data_10_20=>GND0, filter_data_10_19=>GND0, filter_data_10_18=>
      GND0, filter_data_10_17=>GND0, filter_data_10_16=>GND0, 
      filter_data_10_15=>GND0, filter_data_10_14=>filter_data_10_14, 
      filter_data_10_13=>filter_data_10_13, filter_data_10_12=>
      filter_data_10_12, filter_data_10_11=>filter_data_10_11, 
      filter_data_10_10=>filter_data_10_10, filter_data_10_9=>
      filter_data_10_9, filter_data_10_8=>filter_data_10_8, filter_data_10_7
      =>filter_data_10_7, filter_data_10_6=>filter_data_10_6, 
      filter_data_10_5=>filter_data_10_5, filter_data_10_4=>filter_data_10_4, 
      filter_data_10_3=>filter_data_10_3, filter_data_10_2=>filter_data_10_2, 
      filter_data_10_1=>filter_data_10_1, filter_data_10_0=>filter_data_10_0, 
      filter_data_11_31=>filter_data_11_15, filter_data_11_30=>GND0, 
      filter_data_11_29=>GND0, filter_data_11_28=>GND0, filter_data_11_27=>
      GND0, filter_data_11_26=>GND0, filter_data_11_25=>GND0, 
      filter_data_11_24=>GND0, filter_data_11_23=>GND0, filter_data_11_22=>
      GND0, filter_data_11_21=>GND0, filter_data_11_20=>GND0, 
      filter_data_11_19=>GND0, filter_data_11_18=>GND0, filter_data_11_17=>
      GND0, filter_data_11_16=>GND0, filter_data_11_15=>GND0, 
      filter_data_11_14=>filter_data_11_14, filter_data_11_13=>
      filter_data_11_13, filter_data_11_12=>filter_data_11_12, 
      filter_data_11_11=>filter_data_11_11, filter_data_11_10=>
      filter_data_11_10, filter_data_11_9=>filter_data_11_9, 
      filter_data_11_8=>filter_data_11_8, filter_data_11_7=>filter_data_11_7, 
      filter_data_11_6=>filter_data_11_6, filter_data_11_5=>filter_data_11_5, 
      filter_data_11_4=>filter_data_11_4, filter_data_11_3=>filter_data_11_3, 
      filter_data_11_2=>filter_data_11_2, filter_data_11_1=>filter_data_11_1, 
      filter_data_11_0=>filter_data_11_0, filter_data_12_31=>
      filter_data_12_15, filter_data_12_30=>GND0, filter_data_12_29=>GND0, 
      filter_data_12_28=>GND0, filter_data_12_27=>GND0, filter_data_12_26=>
      GND0, filter_data_12_25=>GND0, filter_data_12_24=>GND0, 
      filter_data_12_23=>GND0, filter_data_12_22=>GND0, filter_data_12_21=>
      GND0, filter_data_12_20=>GND0, filter_data_12_19=>GND0, 
      filter_data_12_18=>GND0, filter_data_12_17=>GND0, filter_data_12_16=>
      GND0, filter_data_12_15=>GND0, filter_data_12_14=>filter_data_12_14, 
      filter_data_12_13=>filter_data_12_13, filter_data_12_12=>
      filter_data_12_12, filter_data_12_11=>filter_data_12_11, 
      filter_data_12_10=>filter_data_12_10, filter_data_12_9=>
      filter_data_12_9, filter_data_12_8=>filter_data_12_8, filter_data_12_7
      =>filter_data_12_7, filter_data_12_6=>filter_data_12_6, 
      filter_data_12_5=>filter_data_12_5, filter_data_12_4=>filter_data_12_4, 
      filter_data_12_3=>filter_data_12_3, filter_data_12_2=>filter_data_12_2, 
      filter_data_12_1=>filter_data_12_1, filter_data_12_0=>filter_data_12_0, 
      filter_data_13_31=>filter_data_13_15, filter_data_13_30=>GND0, 
      filter_data_13_29=>GND0, filter_data_13_28=>GND0, filter_data_13_27=>
      GND0, filter_data_13_26=>GND0, filter_data_13_25=>GND0, 
      filter_data_13_24=>GND0, filter_data_13_23=>GND0, filter_data_13_22=>
      GND0, filter_data_13_21=>GND0, filter_data_13_20=>GND0, 
      filter_data_13_19=>GND0, filter_data_13_18=>GND0, filter_data_13_17=>
      GND0, filter_data_13_16=>GND0, filter_data_13_15=>GND0, 
      filter_data_13_14=>filter_data_13_14, filter_data_13_13=>
      filter_data_13_13, filter_data_13_12=>filter_data_13_12, 
      filter_data_13_11=>filter_data_13_11, filter_data_13_10=>
      filter_data_13_10, filter_data_13_9=>filter_data_13_9, 
      filter_data_13_8=>filter_data_13_8, filter_data_13_7=>filter_data_13_7, 
      filter_data_13_6=>filter_data_13_6, filter_data_13_5=>filter_data_13_5, 
      filter_data_13_4=>filter_data_13_4, filter_data_13_3=>filter_data_13_3, 
      filter_data_13_2=>filter_data_13_2, filter_data_13_1=>filter_data_13_1, 
      filter_data_13_0=>filter_data_13_0, filter_data_14_31=>
      filter_data_14_15, filter_data_14_30=>GND0, filter_data_14_29=>GND0, 
      filter_data_14_28=>GND0, filter_data_14_27=>GND0, filter_data_14_26=>
      GND0, filter_data_14_25=>GND0, filter_data_14_24=>GND0, 
      filter_data_14_23=>GND0, filter_data_14_22=>GND0, filter_data_14_21=>
      GND0, filter_data_14_20=>GND0, filter_data_14_19=>GND0, 
      filter_data_14_18=>GND0, filter_data_14_17=>GND0, filter_data_14_16=>
      GND0, filter_data_14_15=>GND0, filter_data_14_14=>filter_data_14_14, 
      filter_data_14_13=>filter_data_14_13, filter_data_14_12=>
      filter_data_14_12, filter_data_14_11=>filter_data_14_11, 
      filter_data_14_10=>filter_data_14_10, filter_data_14_9=>
      filter_data_14_9, filter_data_14_8=>filter_data_14_8, filter_data_14_7
      =>filter_data_14_7, filter_data_14_6=>filter_data_14_6, 
      filter_data_14_5=>filter_data_14_5, filter_data_14_4=>filter_data_14_4, 
      filter_data_14_3=>filter_data_14_3, filter_data_14_2=>filter_data_14_2, 
      filter_data_14_1=>filter_data_14_1, filter_data_14_0=>filter_data_14_0, 
      filter_data_15_31=>filter_data_15_15, filter_data_15_30=>GND0, 
      filter_data_15_29=>GND0, filter_data_15_28=>GND0, filter_data_15_27=>
      GND0, filter_data_15_26=>GND0, filter_data_15_25=>GND0, 
      filter_data_15_24=>GND0, filter_data_15_23=>GND0, filter_data_15_22=>
      GND0, filter_data_15_21=>GND0, filter_data_15_20=>GND0, 
      filter_data_15_19=>GND0, filter_data_15_18=>GND0, filter_data_15_17=>
      GND0, filter_data_15_16=>GND0, filter_data_15_15=>GND0, 
      filter_data_15_14=>filter_data_15_14, filter_data_15_13=>
      filter_data_15_13, filter_data_15_12=>filter_data_15_12, 
      filter_data_15_11=>filter_data_15_11, filter_data_15_10=>
      filter_data_15_10, filter_data_15_9=>filter_data_15_9, 
      filter_data_15_8=>filter_data_15_8, filter_data_15_7=>filter_data_15_7, 
      filter_data_15_6=>filter_data_15_6, filter_data_15_5=>filter_data_15_5, 
      filter_data_15_4=>filter_data_15_4, filter_data_15_3=>filter_data_15_3, 
      filter_data_15_2=>filter_data_15_2, filter_data_15_1=>filter_data_15_1, 
      filter_data_15_0=>filter_data_15_0, filter_data_16_31=>
      filter_data_16_15, filter_data_16_30=>GND0, filter_data_16_29=>GND0, 
      filter_data_16_28=>GND0, filter_data_16_27=>GND0, filter_data_16_26=>
      GND0, filter_data_16_25=>GND0, filter_data_16_24=>GND0, 
      filter_data_16_23=>GND0, filter_data_16_22=>GND0, filter_data_16_21=>
      GND0, filter_data_16_20=>GND0, filter_data_16_19=>GND0, 
      filter_data_16_18=>GND0, filter_data_16_17=>GND0, filter_data_16_16=>
      GND0, filter_data_16_15=>GND0, filter_data_16_14=>filter_data_16_14, 
      filter_data_16_13=>filter_data_16_13, filter_data_16_12=>
      filter_data_16_12, filter_data_16_11=>filter_data_16_11, 
      filter_data_16_10=>filter_data_16_10, filter_data_16_9=>
      filter_data_16_9, filter_data_16_8=>filter_data_16_8, filter_data_16_7
      =>filter_data_16_7, filter_data_16_6=>filter_data_16_6, 
      filter_data_16_5=>filter_data_16_5, filter_data_16_4=>filter_data_16_4, 
      filter_data_16_3=>filter_data_16_3, filter_data_16_2=>filter_data_16_2, 
      filter_data_16_1=>filter_data_16_1, filter_data_16_0=>filter_data_16_0, 
      filter_data_17_31=>filter_data_17_15, filter_data_17_30=>GND0, 
      filter_data_17_29=>GND0, filter_data_17_28=>GND0, filter_data_17_27=>
      GND0, filter_data_17_26=>GND0, filter_data_17_25=>GND0, 
      filter_data_17_24=>GND0, filter_data_17_23=>GND0, filter_data_17_22=>
      GND0, filter_data_17_21=>GND0, filter_data_17_20=>GND0, 
      filter_data_17_19=>GND0, filter_data_17_18=>GND0, filter_data_17_17=>
      GND0, filter_data_17_16=>GND0, filter_data_17_15=>GND0, 
      filter_data_17_14=>filter_data_17_14, filter_data_17_13=>
      filter_data_17_13, filter_data_17_12=>filter_data_17_12, 
      filter_data_17_11=>filter_data_17_11, filter_data_17_10=>
      filter_data_17_10, filter_data_17_9=>filter_data_17_9, 
      filter_data_17_8=>filter_data_17_8, filter_data_17_7=>filter_data_17_7, 
      filter_data_17_6=>filter_data_17_6, filter_data_17_5=>filter_data_17_5, 
      filter_data_17_4=>filter_data_17_4, filter_data_17_3=>filter_data_17_3, 
      filter_data_17_2=>filter_data_17_2, filter_data_17_1=>filter_data_17_1, 
      filter_data_17_0=>filter_data_17_0, filter_data_18_31=>GND0, 
      filter_data_18_30=>GND0, filter_data_18_29=>GND0, filter_data_18_28=>
      GND0, filter_data_18_27=>GND0, filter_data_18_26=>GND0, 
      filter_data_18_25=>GND0, filter_data_18_24=>GND0, filter_data_18_23=>
      GND0, filter_data_18_22=>GND0, filter_data_18_21=>GND0, 
      filter_data_18_20=>GND0, filter_data_18_19=>GND0, filter_data_18_18=>
      GND0, filter_data_18_17=>GND0, filter_data_18_16=>GND0, 
      filter_data_18_15=>GND0, filter_data_18_14=>GND0, filter_data_18_13=>
      GND0, filter_data_18_12=>GND0, filter_data_18_11=>GND0, 
      filter_data_18_10=>GND0, filter_data_18_9=>GND0, filter_data_18_8=>
      GND0, filter_data_18_7=>GND0, filter_data_18_6=>GND0, filter_data_18_5
      =>GND0, filter_data_18_4=>GND0, filter_data_18_3=>GND0, 
      filter_data_18_2=>GND0, filter_data_18_1=>GND0, filter_data_18_0=>GND0, 
      filter_data_19_31=>GND0, filter_data_19_30=>GND0, filter_data_19_29=>
      GND0, filter_data_19_28=>GND0, filter_data_19_27=>GND0, 
      filter_data_19_26=>GND0, filter_data_19_25=>GND0, filter_data_19_24=>
      GND0, filter_data_19_23=>GND0, filter_data_19_22=>GND0, 
      filter_data_19_21=>GND0, filter_data_19_20=>GND0, filter_data_19_19=>
      GND0, filter_data_19_18=>GND0, filter_data_19_17=>GND0, 
      filter_data_19_16=>GND0, filter_data_19_15=>GND0, filter_data_19_14=>
      GND0, filter_data_19_13=>GND0, filter_data_19_12=>GND0, 
      filter_data_19_11=>GND0, filter_data_19_10=>GND0, filter_data_19_9=>
      GND0, filter_data_19_8=>GND0, filter_data_19_7=>GND0, filter_data_19_6
      =>GND0, filter_data_19_5=>GND0, filter_data_19_4=>GND0, 
      filter_data_19_3=>GND0, filter_data_19_2=>GND0, filter_data_19_1=>GND0, 
      filter_data_19_0=>GND0, filter_data_20_31=>GND0, filter_data_20_30=>
      GND0, filter_data_20_29=>GND0, filter_data_20_28=>GND0, 
      filter_data_20_27=>GND0, filter_data_20_26=>GND0, filter_data_20_25=>
      GND0, filter_data_20_24=>GND0, filter_data_20_23=>GND0, 
      filter_data_20_22=>GND0, filter_data_20_21=>GND0, filter_data_20_20=>
      GND0, filter_data_20_19=>GND0, filter_data_20_18=>GND0, 
      filter_data_20_17=>GND0, filter_data_20_16=>GND0, filter_data_20_15=>
      GND0, filter_data_20_14=>GND0, filter_data_20_13=>GND0, 
      filter_data_20_12=>GND0, filter_data_20_11=>GND0, filter_data_20_10=>
      GND0, filter_data_20_9=>GND0, filter_data_20_8=>GND0, filter_data_20_7
      =>GND0, filter_data_20_6=>GND0, filter_data_20_5=>GND0, 
      filter_data_20_4=>GND0, filter_data_20_3=>GND0, filter_data_20_2=>GND0, 
      filter_data_20_1=>GND0, filter_data_20_0=>GND0, filter_data_21_31=>
      GND0, filter_data_21_30=>GND0, filter_data_21_29=>GND0, 
      filter_data_21_28=>GND0, filter_data_21_27=>GND0, filter_data_21_26=>
      GND0, filter_data_21_25=>GND0, filter_data_21_24=>GND0, 
      filter_data_21_23=>GND0, filter_data_21_22=>GND0, filter_data_21_21=>
      GND0, filter_data_21_20=>GND0, filter_data_21_19=>GND0, 
      filter_data_21_18=>GND0, filter_data_21_17=>GND0, filter_data_21_16=>
      GND0, filter_data_21_15=>GND0, filter_data_21_14=>GND0, 
      filter_data_21_13=>GND0, filter_data_21_12=>GND0, filter_data_21_11=>
      GND0, filter_data_21_10=>GND0, filter_data_21_9=>GND0, 
      filter_data_21_8=>GND0, filter_data_21_7=>GND0, filter_data_21_6=>GND0, 
      filter_data_21_5=>GND0, filter_data_21_4=>GND0, filter_data_21_3=>GND0, 
      filter_data_21_2=>GND0, filter_data_21_1=>GND0, filter_data_21_0=>GND0, 
      filter_data_22_31=>GND0, filter_data_22_30=>GND0, filter_data_22_29=>
      GND0, filter_data_22_28=>GND0, filter_data_22_27=>GND0, 
      filter_data_22_26=>GND0, filter_data_22_25=>GND0, filter_data_22_24=>
      GND0, filter_data_22_23=>GND0, filter_data_22_22=>GND0, 
      filter_data_22_21=>GND0, filter_data_22_20=>GND0, filter_data_22_19=>
      GND0, filter_data_22_18=>GND0, filter_data_22_17=>GND0, 
      filter_data_22_16=>GND0, filter_data_22_15=>GND0, filter_data_22_14=>
      GND0, filter_data_22_13=>GND0, filter_data_22_12=>GND0, 
      filter_data_22_11=>GND0, filter_data_22_10=>GND0, filter_data_22_9=>
      GND0, filter_data_22_8=>GND0, filter_data_22_7=>GND0, filter_data_22_6
      =>GND0, filter_data_22_5=>GND0, filter_data_22_4=>GND0, 
      filter_data_22_3=>GND0, filter_data_22_2=>GND0, filter_data_22_1=>GND0, 
      filter_data_22_0=>GND0, filter_data_23_31=>GND0, filter_data_23_30=>
      GND0, filter_data_23_29=>GND0, filter_data_23_28=>GND0, 
      filter_data_23_27=>GND0, filter_data_23_26=>GND0, filter_data_23_25=>
      GND0, filter_data_23_24=>GND0, filter_data_23_23=>GND0, 
      filter_data_23_22=>GND0, filter_data_23_21=>GND0, filter_data_23_20=>
      GND0, filter_data_23_19=>GND0, filter_data_23_18=>GND0, 
      filter_data_23_17=>GND0, filter_data_23_16=>GND0, filter_data_23_15=>
      GND0, filter_data_23_14=>GND0, filter_data_23_13=>GND0, 
      filter_data_23_12=>GND0, filter_data_23_11=>GND0, filter_data_23_10=>
      GND0, filter_data_23_9=>GND0, filter_data_23_8=>GND0, filter_data_23_7
      =>GND0, filter_data_23_6=>GND0, filter_data_23_5=>GND0, 
      filter_data_23_4=>GND0, filter_data_23_3=>GND0, filter_data_23_2=>GND0, 
      filter_data_23_1=>GND0, filter_data_23_0=>GND0, filter_data_24_31=>
      GND0, filter_data_24_30=>GND0, filter_data_24_29=>GND0, 
      filter_data_24_28=>GND0, filter_data_24_27=>GND0, filter_data_24_26=>
      GND0, filter_data_24_25=>GND0, filter_data_24_24=>GND0, 
      filter_data_24_23=>GND0, filter_data_24_22=>GND0, filter_data_24_21=>
      GND0, filter_data_24_20=>GND0, filter_data_24_19=>GND0, 
      filter_data_24_18=>GND0, filter_data_24_17=>GND0, filter_data_24_16=>
      GND0, filter_data_24_15=>GND0, filter_data_24_14=>GND0, 
      filter_data_24_13=>GND0, filter_data_24_12=>GND0, filter_data_24_11=>
      GND0, filter_data_24_10=>GND0, filter_data_24_9=>GND0, 
      filter_data_24_8=>GND0, filter_data_24_7=>GND0, filter_data_24_6=>GND0, 
      filter_data_24_5=>GND0, filter_data_24_4=>GND0, filter_data_24_3=>GND0, 
      filter_data_24_2=>GND0, filter_data_24_1=>GND0, filter_data_24_0=>GND0, 
      filter_size=>nx16665, ordered_img_data_0_31=>DANGLING(0), 
      ordered_img_data_0_30=>DANGLING(1), ordered_img_data_0_29=>DANGLING(2), 
      ordered_img_data_0_28=>DANGLING(3), ordered_img_data_0_27=>DANGLING(4), 
      ordered_img_data_0_26=>DANGLING(5), ordered_img_data_0_25=>DANGLING(6), 
      ordered_img_data_0_24=>DANGLING(7), ordered_img_data_0_23=>DANGLING(8), 
      ordered_img_data_0_22=>DANGLING(9), ordered_img_data_0_21=>DANGLING(10
      ), ordered_img_data_0_20=>DANGLING(11), ordered_img_data_0_19=>
      DANGLING(12), ordered_img_data_0_18=>DANGLING(13), 
      ordered_img_data_0_17=>DANGLING(14), ordered_img_data_0_16=>DANGLING(
      15), ordered_img_data_0_15=>DANGLING(16), ordered_img_data_0_14=>
      DANGLING(17), ordered_img_data_0_13=>DANGLING(18), 
      ordered_img_data_0_12=>DANGLING(19), ordered_img_data_0_11=>DANGLING(
      20), ordered_img_data_0_10=>DANGLING(21), ordered_img_data_0_9=>
      DANGLING(22), ordered_img_data_0_8=>DANGLING(23), ordered_img_data_0_7
      =>DANGLING(24), ordered_img_data_0_6=>DANGLING(25), 
      ordered_img_data_0_5=>DANGLING(26), ordered_img_data_0_4=>DANGLING(27), 
      ordered_img_data_0_3=>DANGLING(28), ordered_img_data_0_2=>DANGLING(29), 
      ordered_img_data_0_1=>DANGLING(30), ordered_img_data_0_0=>DANGLING(31), 
      ordered_img_data_1_31=>DANGLING(32), ordered_img_data_1_30=>DANGLING(
      33), ordered_img_data_1_29=>DANGLING(34), ordered_img_data_1_28=>
      DANGLING(35), ordered_img_data_1_27=>DANGLING(36), 
      ordered_img_data_1_26=>DANGLING(37), ordered_img_data_1_25=>DANGLING(
      38), ordered_img_data_1_24=>DANGLING(39), ordered_img_data_1_23=>
      DANGLING(40), ordered_img_data_1_22=>DANGLING(41), 
      ordered_img_data_1_21=>DANGLING(42), ordered_img_data_1_20=>DANGLING(
      43), ordered_img_data_1_19=>DANGLING(44), ordered_img_data_1_18=>
      DANGLING(45), ordered_img_data_1_17=>DANGLING(46), 
      ordered_img_data_1_16=>DANGLING(47), ordered_img_data_1_15=>DANGLING(
      48), ordered_img_data_1_14=>DANGLING(49), ordered_img_data_1_13=>
      DANGLING(50), ordered_img_data_1_12=>DANGLING(51), 
      ordered_img_data_1_11=>DANGLING(52), ordered_img_data_1_10=>DANGLING(
      53), ordered_img_data_1_9=>DANGLING(54), ordered_img_data_1_8=>
      DANGLING(55), ordered_img_data_1_7=>DANGLING(56), ordered_img_data_1_6
      =>DANGLING(57), ordered_img_data_1_5=>DANGLING(58), 
      ordered_img_data_1_4=>DANGLING(59), ordered_img_data_1_3=>DANGLING(60), 
      ordered_img_data_1_2=>DANGLING(61), ordered_img_data_1_1=>DANGLING(62), 
      ordered_img_data_1_0=>DANGLING(63), ordered_img_data_2_31=>DANGLING(64
      ), ordered_img_data_2_30=>DANGLING(65), ordered_img_data_2_29=>
      DANGLING(66), ordered_img_data_2_28=>DANGLING(67), 
      ordered_img_data_2_27=>DANGLING(68), ordered_img_data_2_26=>DANGLING(
      69), ordered_img_data_2_25=>DANGLING(70), ordered_img_data_2_24=>
      DANGLING(71), ordered_img_data_2_23=>DANGLING(72), 
      ordered_img_data_2_22=>DANGLING(73), ordered_img_data_2_21=>DANGLING(
      74), ordered_img_data_2_20=>DANGLING(75), ordered_img_data_2_19=>
      DANGLING(76), ordered_img_data_2_18=>DANGLING(77), 
      ordered_img_data_2_17=>DANGLING(78), ordered_img_data_2_16=>DANGLING(
      79), ordered_img_data_2_15=>DANGLING(80), ordered_img_data_2_14=>
      DANGLING(81), ordered_img_data_2_13=>DANGLING(82), 
      ordered_img_data_2_12=>DANGLING(83), ordered_img_data_2_11=>DANGLING(
      84), ordered_img_data_2_10=>DANGLING(85), ordered_img_data_2_9=>
      DANGLING(86), ordered_img_data_2_8=>DANGLING(87), ordered_img_data_2_7
      =>DANGLING(88), ordered_img_data_2_6=>DANGLING(89), 
      ordered_img_data_2_5=>DANGLING(90), ordered_img_data_2_4=>DANGLING(91), 
      ordered_img_data_2_3=>DANGLING(92), ordered_img_data_2_2=>DANGLING(93), 
      ordered_img_data_2_1=>DANGLING(94), ordered_img_data_2_0=>DANGLING(95), 
      ordered_img_data_3_31=>DANGLING(96), ordered_img_data_3_30=>DANGLING(
      97), ordered_img_data_3_29=>DANGLING(98), ordered_img_data_3_28=>
      DANGLING(99), ordered_img_data_3_27=>DANGLING(100), 
      ordered_img_data_3_26=>DANGLING(101), ordered_img_data_3_25=>DANGLING(
      102), ordered_img_data_3_24=>DANGLING(103), ordered_img_data_3_23=>
      DANGLING(104), ordered_img_data_3_22=>DANGLING(105), 
      ordered_img_data_3_21=>DANGLING(106), ordered_img_data_3_20=>DANGLING(
      107), ordered_img_data_3_19=>DANGLING(108), ordered_img_data_3_18=>
      DANGLING(109), ordered_img_data_3_17=>DANGLING(110), 
      ordered_img_data_3_16=>DANGLING(111), ordered_img_data_3_15=>DANGLING(
      112), ordered_img_data_3_14=>DANGLING(113), ordered_img_data_3_13=>
      DANGLING(114), ordered_img_data_3_12=>DANGLING(115), 
      ordered_img_data_3_11=>DANGLING(116), ordered_img_data_3_10=>DANGLING(
      117), ordered_img_data_3_9=>DANGLING(118), ordered_img_data_3_8=>
      DANGLING(119), ordered_img_data_3_7=>DANGLING(120), 
      ordered_img_data_3_6=>DANGLING(121), ordered_img_data_3_5=>DANGLING(
      122), ordered_img_data_3_4=>DANGLING(123), ordered_img_data_3_3=>
      DANGLING(124), ordered_img_data_3_2=>DANGLING(125), 
      ordered_img_data_3_1=>DANGLING(126), ordered_img_data_3_0=>DANGLING(
      127), ordered_img_data_4_31=>DANGLING(128), ordered_img_data_4_30=>
      DANGLING(129), ordered_img_data_4_29=>DANGLING(130), 
      ordered_img_data_4_28=>DANGLING(131), ordered_img_data_4_27=>DANGLING(
      132), ordered_img_data_4_26=>DANGLING(133), ordered_img_data_4_25=>
      DANGLING(134), ordered_img_data_4_24=>DANGLING(135), 
      ordered_img_data_4_23=>DANGLING(136), ordered_img_data_4_22=>DANGLING(
      137), ordered_img_data_4_21=>DANGLING(138), ordered_img_data_4_20=>
      DANGLING(139), ordered_img_data_4_19=>DANGLING(140), 
      ordered_img_data_4_18=>DANGLING(141), ordered_img_data_4_17=>DANGLING(
      142), ordered_img_data_4_16=>DANGLING(143), ordered_img_data_4_15=>
      DANGLING(144), ordered_img_data_4_14=>DANGLING(145), 
      ordered_img_data_4_13=>DANGLING(146), ordered_img_data_4_12=>DANGLING(
      147), ordered_img_data_4_11=>DANGLING(148), ordered_img_data_4_10=>
      DANGLING(149), ordered_img_data_4_9=>DANGLING(150), 
      ordered_img_data_4_8=>DANGLING(151), ordered_img_data_4_7=>DANGLING(
      152), ordered_img_data_4_6=>DANGLING(153), ordered_img_data_4_5=>
      DANGLING(154), ordered_img_data_4_4=>DANGLING(155), 
      ordered_img_data_4_3=>DANGLING(156), ordered_img_data_4_2=>DANGLING(
      157), ordered_img_data_4_1=>DANGLING(158), ordered_img_data_4_0=>
      DANGLING(159), ordered_img_data_5_31=>DANGLING(160), 
      ordered_img_data_5_30=>DANGLING(161), ordered_img_data_5_29=>DANGLING(
      162), ordered_img_data_5_28=>DANGLING(163), ordered_img_data_5_27=>
      DANGLING(164), ordered_img_data_5_26=>DANGLING(165), 
      ordered_img_data_5_25=>DANGLING(166), ordered_img_data_5_24=>DANGLING(
      167), ordered_img_data_5_23=>DANGLING(168), ordered_img_data_5_22=>
      DANGLING(169), ordered_img_data_5_21=>DANGLING(170), 
      ordered_img_data_5_20=>DANGLING(171), ordered_img_data_5_19=>DANGLING(
      172), ordered_img_data_5_18=>DANGLING(173), ordered_img_data_5_17=>
      DANGLING(174), ordered_img_data_5_16=>DANGLING(175), 
      ordered_img_data_5_15=>DANGLING(176), ordered_img_data_5_14=>DANGLING(
      177), ordered_img_data_5_13=>DANGLING(178), ordered_img_data_5_12=>
      DANGLING(179), ordered_img_data_5_11=>DANGLING(180), 
      ordered_img_data_5_10=>DANGLING(181), ordered_img_data_5_9=>DANGLING(
      182), ordered_img_data_5_8=>DANGLING(183), ordered_img_data_5_7=>
      DANGLING(184), ordered_img_data_5_6=>DANGLING(185), 
      ordered_img_data_5_5=>DANGLING(186), ordered_img_data_5_4=>DANGLING(
      187), ordered_img_data_5_3=>DANGLING(188), ordered_img_data_5_2=>
      DANGLING(189), ordered_img_data_5_1=>DANGLING(190), 
      ordered_img_data_5_0=>DANGLING(191), ordered_img_data_6_31=>DANGLING(
      192), ordered_img_data_6_30=>DANGLING(193), ordered_img_data_6_29=>
      DANGLING(194), ordered_img_data_6_28=>DANGLING(195), 
      ordered_img_data_6_27=>DANGLING(196), ordered_img_data_6_26=>DANGLING(
      197), ordered_img_data_6_25=>DANGLING(198), ordered_img_data_6_24=>
      DANGLING(199), ordered_img_data_6_23=>DANGLING(200), 
      ordered_img_data_6_22=>DANGLING(201), ordered_img_data_6_21=>DANGLING(
      202), ordered_img_data_6_20=>DANGLING(203), ordered_img_data_6_19=>
      DANGLING(204), ordered_img_data_6_18=>DANGLING(205), 
      ordered_img_data_6_17=>DANGLING(206), ordered_img_data_6_16=>DANGLING(
      207), ordered_img_data_6_15=>DANGLING(208), ordered_img_data_6_14=>
      DANGLING(209), ordered_img_data_6_13=>DANGLING(210), 
      ordered_img_data_6_12=>DANGLING(211), ordered_img_data_6_11=>DANGLING(
      212), ordered_img_data_6_10=>DANGLING(213), ordered_img_data_6_9=>
      DANGLING(214), ordered_img_data_6_8=>DANGLING(215), 
      ordered_img_data_6_7=>DANGLING(216), ordered_img_data_6_6=>DANGLING(
      217), ordered_img_data_6_5=>DANGLING(218), ordered_img_data_6_4=>
      DANGLING(219), ordered_img_data_6_3=>DANGLING(220), 
      ordered_img_data_6_2=>DANGLING(221), ordered_img_data_6_1=>DANGLING(
      222), ordered_img_data_6_0=>DANGLING(223), ordered_img_data_7_31=>
      DANGLING(224), ordered_img_data_7_30=>DANGLING(225), 
      ordered_img_data_7_29=>DANGLING(226), ordered_img_data_7_28=>DANGLING(
      227), ordered_img_data_7_27=>DANGLING(228), ordered_img_data_7_26=>
      DANGLING(229), ordered_img_data_7_25=>DANGLING(230), 
      ordered_img_data_7_24=>DANGLING(231), ordered_img_data_7_23=>DANGLING(
      232), ordered_img_data_7_22=>DANGLING(233), ordered_img_data_7_21=>
      DANGLING(234), ordered_img_data_7_20=>DANGLING(235), 
      ordered_img_data_7_19=>DANGLING(236), ordered_img_data_7_18=>DANGLING(
      237), ordered_img_data_7_17=>DANGLING(238), ordered_img_data_7_16=>
      DANGLING(239), ordered_img_data_7_15=>DANGLING(240), 
      ordered_img_data_7_14=>DANGLING(241), ordered_img_data_7_13=>DANGLING(
      242), ordered_img_data_7_12=>DANGLING(243), ordered_img_data_7_11=>
      DANGLING(244), ordered_img_data_7_10=>DANGLING(245), 
      ordered_img_data_7_9=>DANGLING(246), ordered_img_data_7_8=>DANGLING(
      247), ordered_img_data_7_7=>DANGLING(248), ordered_img_data_7_6=>
      DANGLING(249), ordered_img_data_7_5=>DANGLING(250), 
      ordered_img_data_7_4=>DANGLING(251), ordered_img_data_7_3=>DANGLING(
      252), ordered_img_data_7_2=>DANGLING(253), ordered_img_data_7_1=>
      DANGLING(254), ordered_img_data_7_0=>DANGLING(255), 
      ordered_img_data_8_31=>DANGLING(256), ordered_img_data_8_30=>DANGLING(
      257), ordered_img_data_8_29=>DANGLING(258), ordered_img_data_8_28=>
      DANGLING(259), ordered_img_data_8_27=>DANGLING(260), 
      ordered_img_data_8_26=>DANGLING(261), ordered_img_data_8_25=>DANGLING(
      262), ordered_img_data_8_24=>DANGLING(263), ordered_img_data_8_23=>
      DANGLING(264), ordered_img_data_8_22=>DANGLING(265), 
      ordered_img_data_8_21=>DANGLING(266), ordered_img_data_8_20=>DANGLING(
      267), ordered_img_data_8_19=>DANGLING(268), ordered_img_data_8_18=>
      DANGLING(269), ordered_img_data_8_17=>DANGLING(270), 
      ordered_img_data_8_16=>DANGLING(271), ordered_img_data_8_15=>DANGLING(
      272), ordered_img_data_8_14=>DANGLING(273), ordered_img_data_8_13=>
      DANGLING(274), ordered_img_data_8_12=>DANGLING(275), 
      ordered_img_data_8_11=>DANGLING(276), ordered_img_data_8_10=>DANGLING(
      277), ordered_img_data_8_9=>DANGLING(278), ordered_img_data_8_8=>
      DANGLING(279), ordered_img_data_8_7=>DANGLING(280), 
      ordered_img_data_8_6=>DANGLING(281), ordered_img_data_8_5=>DANGLING(
      282), ordered_img_data_8_4=>DANGLING(283), ordered_img_data_8_3=>
      DANGLING(284), ordered_img_data_8_2=>DANGLING(285), 
      ordered_img_data_8_1=>DANGLING(286), ordered_img_data_8_0=>DANGLING(
      287), ordered_img_data_9_31=>ordered_img_data_9_31, 
      ordered_img_data_9_30=>DANGLING(288), ordered_img_data_9_29=>DANGLING(
      289), ordered_img_data_9_28=>DANGLING(290), ordered_img_data_9_27=>
      DANGLING(291), ordered_img_data_9_26=>DANGLING(292), 
      ordered_img_data_9_25=>DANGLING(293), ordered_img_data_9_24=>DANGLING(
      294), ordered_img_data_9_23=>DANGLING(295), ordered_img_data_9_22=>
      DANGLING(296), ordered_img_data_9_21=>DANGLING(297), 
      ordered_img_data_9_20=>DANGLING(298), ordered_img_data_9_19=>DANGLING(
      299), ordered_img_data_9_18=>DANGLING(300), ordered_img_data_9_17=>
      DANGLING(301), ordered_img_data_9_16=>DANGLING(302), 
      ordered_img_data_9_15=>DANGLING(303), ordered_img_data_9_14=>
      ordered_img_data_9_14, ordered_img_data_9_13=>ordered_img_data_9_13, 
      ordered_img_data_9_12=>ordered_img_data_9_12, ordered_img_data_9_11=>
      ordered_img_data_9_11, ordered_img_data_9_10=>ordered_img_data_9_10, 
      ordered_img_data_9_9=>ordered_img_data_9_9, ordered_img_data_9_8=>
      ordered_img_data_9_8, ordered_img_data_9_7=>ordered_img_data_9_7, 
      ordered_img_data_9_6=>ordered_img_data_9_6, ordered_img_data_9_5=>
      ordered_img_data_9_5, ordered_img_data_9_4=>ordered_img_data_9_4, 
      ordered_img_data_9_3=>ordered_img_data_9_3, ordered_img_data_9_2=>
      ordered_img_data_9_2, ordered_img_data_9_1=>ordered_img_data_9_1, 
      ordered_img_data_9_0=>ordered_img_data_9_0, ordered_img_data_10_31=>
      ordered_img_data_10_31, ordered_img_data_10_30=>DANGLING(304), 
      ordered_img_data_10_29=>DANGLING(305), ordered_img_data_10_28=>
      DANGLING(306), ordered_img_data_10_27=>DANGLING(307), 
      ordered_img_data_10_26=>DANGLING(308), ordered_img_data_10_25=>
      DANGLING(309), ordered_img_data_10_24=>DANGLING(310), 
      ordered_img_data_10_23=>DANGLING(311), ordered_img_data_10_22=>
      DANGLING(312), ordered_img_data_10_21=>DANGLING(313), 
      ordered_img_data_10_20=>DANGLING(314), ordered_img_data_10_19=>
      DANGLING(315), ordered_img_data_10_18=>DANGLING(316), 
      ordered_img_data_10_17=>DANGLING(317), ordered_img_data_10_16=>
      DANGLING(318), ordered_img_data_10_15=>DANGLING(319), 
      ordered_img_data_10_14=>ordered_img_data_10_14, ordered_img_data_10_13
      =>ordered_img_data_10_13, ordered_img_data_10_12=>
      ordered_img_data_10_12, ordered_img_data_10_11=>ordered_img_data_10_11, 
      ordered_img_data_10_10=>ordered_img_data_10_10, ordered_img_data_10_9
      =>ordered_img_data_10_9, ordered_img_data_10_8=>ordered_img_data_10_8, 
      ordered_img_data_10_7=>ordered_img_data_10_7, ordered_img_data_10_6=>
      ordered_img_data_10_6, ordered_img_data_10_5=>ordered_img_data_10_5, 
      ordered_img_data_10_4=>ordered_img_data_10_4, ordered_img_data_10_3=>
      ordered_img_data_10_3, ordered_img_data_10_2=>ordered_img_data_10_2, 
      ordered_img_data_10_1=>ordered_img_data_10_1, ordered_img_data_10_0=>
      ordered_img_data_10_0, ordered_img_data_11_31=>ordered_img_data_11_31, 
      ordered_img_data_11_30=>DANGLING(320), ordered_img_data_11_29=>
      DANGLING(321), ordered_img_data_11_28=>DANGLING(322), 
      ordered_img_data_11_27=>DANGLING(323), ordered_img_data_11_26=>
      DANGLING(324), ordered_img_data_11_25=>DANGLING(325), 
      ordered_img_data_11_24=>DANGLING(326), ordered_img_data_11_23=>
      DANGLING(327), ordered_img_data_11_22=>DANGLING(328), 
      ordered_img_data_11_21=>DANGLING(329), ordered_img_data_11_20=>
      DANGLING(330), ordered_img_data_11_19=>DANGLING(331), 
      ordered_img_data_11_18=>DANGLING(332), ordered_img_data_11_17=>
      DANGLING(333), ordered_img_data_11_16=>DANGLING(334), 
      ordered_img_data_11_15=>DANGLING(335), ordered_img_data_11_14=>
      ordered_img_data_11_14, ordered_img_data_11_13=>ordered_img_data_11_13, 
      ordered_img_data_11_12=>ordered_img_data_11_12, ordered_img_data_11_11
      =>ordered_img_data_11_11, ordered_img_data_11_10=>
      ordered_img_data_11_10, ordered_img_data_11_9=>ordered_img_data_11_9, 
      ordered_img_data_11_8=>ordered_img_data_11_8, ordered_img_data_11_7=>
      ordered_img_data_11_7, ordered_img_data_11_6=>ordered_img_data_11_6, 
      ordered_img_data_11_5=>ordered_img_data_11_5, ordered_img_data_11_4=>
      ordered_img_data_11_4, ordered_img_data_11_3=>ordered_img_data_11_3, 
      ordered_img_data_11_2=>ordered_img_data_11_2, ordered_img_data_11_1=>
      ordered_img_data_11_1, ordered_img_data_11_0=>ordered_img_data_11_0, 
      ordered_img_data_12_31=>ordered_img_data_12_31, ordered_img_data_12_30
      =>DANGLING(336), ordered_img_data_12_29=>DANGLING(337), 
      ordered_img_data_12_28=>DANGLING(338), ordered_img_data_12_27=>
      DANGLING(339), ordered_img_data_12_26=>DANGLING(340), 
      ordered_img_data_12_25=>DANGLING(341), ordered_img_data_12_24=>
      DANGLING(342), ordered_img_data_12_23=>DANGLING(343), 
      ordered_img_data_12_22=>DANGLING(344), ordered_img_data_12_21=>
      DANGLING(345), ordered_img_data_12_20=>DANGLING(346), 
      ordered_img_data_12_19=>DANGLING(347), ordered_img_data_12_18=>
      DANGLING(348), ordered_img_data_12_17=>DANGLING(349), 
      ordered_img_data_12_16=>DANGLING(350), ordered_img_data_12_15=>
      DANGLING(351), ordered_img_data_12_14=>ordered_img_data_12_14, 
      ordered_img_data_12_13=>ordered_img_data_12_13, ordered_img_data_12_12
      =>ordered_img_data_12_12, ordered_img_data_12_11=>
      ordered_img_data_12_11, ordered_img_data_12_10=>ordered_img_data_12_10, 
      ordered_img_data_12_9=>ordered_img_data_12_9, ordered_img_data_12_8=>
      ordered_img_data_12_8, ordered_img_data_12_7=>ordered_img_data_12_7, 
      ordered_img_data_12_6=>ordered_img_data_12_6, ordered_img_data_12_5=>
      ordered_img_data_12_5, ordered_img_data_12_4=>ordered_img_data_12_4, 
      ordered_img_data_12_3=>ordered_img_data_12_3, ordered_img_data_12_2=>
      ordered_img_data_12_2, ordered_img_data_12_1=>ordered_img_data_12_1, 
      ordered_img_data_12_0=>ordered_img_data_12_0, ordered_img_data_13_31=>
      ordered_img_data_13_31, ordered_img_data_13_30=>DANGLING(352), 
      ordered_img_data_13_29=>DANGLING(353), ordered_img_data_13_28=>
      DANGLING(354), ordered_img_data_13_27=>DANGLING(355), 
      ordered_img_data_13_26=>DANGLING(356), ordered_img_data_13_25=>
      DANGLING(357), ordered_img_data_13_24=>DANGLING(358), 
      ordered_img_data_13_23=>DANGLING(359), ordered_img_data_13_22=>
      DANGLING(360), ordered_img_data_13_21=>DANGLING(361), 
      ordered_img_data_13_20=>DANGLING(362), ordered_img_data_13_19=>
      DANGLING(363), ordered_img_data_13_18=>DANGLING(364), 
      ordered_img_data_13_17=>DANGLING(365), ordered_img_data_13_16=>
      DANGLING(366), ordered_img_data_13_15=>DANGLING(367), 
      ordered_img_data_13_14=>ordered_img_data_13_14, ordered_img_data_13_13
      =>ordered_img_data_13_13, ordered_img_data_13_12=>
      ordered_img_data_13_12, ordered_img_data_13_11=>ordered_img_data_13_11, 
      ordered_img_data_13_10=>ordered_img_data_13_10, ordered_img_data_13_9
      =>ordered_img_data_13_9, ordered_img_data_13_8=>ordered_img_data_13_8, 
      ordered_img_data_13_7=>ordered_img_data_13_7, ordered_img_data_13_6=>
      ordered_img_data_13_6, ordered_img_data_13_5=>ordered_img_data_13_5, 
      ordered_img_data_13_4=>ordered_img_data_13_4, ordered_img_data_13_3=>
      ordered_img_data_13_3, ordered_img_data_13_2=>ordered_img_data_13_2, 
      ordered_img_data_13_1=>ordered_img_data_13_1, ordered_img_data_13_0=>
      ordered_img_data_13_0, ordered_img_data_14_31=>ordered_img_data_14_31, 
      ordered_img_data_14_30=>DANGLING(368), ordered_img_data_14_29=>
      DANGLING(369), ordered_img_data_14_28=>DANGLING(370), 
      ordered_img_data_14_27=>DANGLING(371), ordered_img_data_14_26=>
      DANGLING(372), ordered_img_data_14_25=>DANGLING(373), 
      ordered_img_data_14_24=>DANGLING(374), ordered_img_data_14_23=>
      DANGLING(375), ordered_img_data_14_22=>DANGLING(376), 
      ordered_img_data_14_21=>DANGLING(377), ordered_img_data_14_20=>
      DANGLING(378), ordered_img_data_14_19=>DANGLING(379), 
      ordered_img_data_14_18=>DANGLING(380), ordered_img_data_14_17=>
      DANGLING(381), ordered_img_data_14_16=>DANGLING(382), 
      ordered_img_data_14_15=>DANGLING(383), ordered_img_data_14_14=>
      ordered_img_data_14_14, ordered_img_data_14_13=>ordered_img_data_14_13, 
      ordered_img_data_14_12=>ordered_img_data_14_12, ordered_img_data_14_11
      =>ordered_img_data_14_11, ordered_img_data_14_10=>
      ordered_img_data_14_10, ordered_img_data_14_9=>ordered_img_data_14_9, 
      ordered_img_data_14_8=>ordered_img_data_14_8, ordered_img_data_14_7=>
      ordered_img_data_14_7, ordered_img_data_14_6=>ordered_img_data_14_6, 
      ordered_img_data_14_5=>ordered_img_data_14_5, ordered_img_data_14_4=>
      ordered_img_data_14_4, ordered_img_data_14_3=>ordered_img_data_14_3, 
      ordered_img_data_14_2=>ordered_img_data_14_2, ordered_img_data_14_1=>
      ordered_img_data_14_1, ordered_img_data_14_0=>ordered_img_data_14_0, 
      ordered_img_data_15_31=>ordered_img_data_15_31, ordered_img_data_15_30
      =>DANGLING(384), ordered_img_data_15_29=>DANGLING(385), 
      ordered_img_data_15_28=>DANGLING(386), ordered_img_data_15_27=>
      DANGLING(387), ordered_img_data_15_26=>DANGLING(388), 
      ordered_img_data_15_25=>DANGLING(389), ordered_img_data_15_24=>
      DANGLING(390), ordered_img_data_15_23=>DANGLING(391), 
      ordered_img_data_15_22=>DANGLING(392), ordered_img_data_15_21=>
      DANGLING(393), ordered_img_data_15_20=>DANGLING(394), 
      ordered_img_data_15_19=>DANGLING(395), ordered_img_data_15_18=>
      DANGLING(396), ordered_img_data_15_17=>DANGLING(397), 
      ordered_img_data_15_16=>DANGLING(398), ordered_img_data_15_15=>
      DANGLING(399), ordered_img_data_15_14=>ordered_img_data_15_14, 
      ordered_img_data_15_13=>ordered_img_data_15_13, ordered_img_data_15_12
      =>ordered_img_data_15_12, ordered_img_data_15_11=>
      ordered_img_data_15_11, ordered_img_data_15_10=>ordered_img_data_15_10, 
      ordered_img_data_15_9=>ordered_img_data_15_9, ordered_img_data_15_8=>
      ordered_img_data_15_8, ordered_img_data_15_7=>ordered_img_data_15_7, 
      ordered_img_data_15_6=>ordered_img_data_15_6, ordered_img_data_15_5=>
      ordered_img_data_15_5, ordered_img_data_15_4=>ordered_img_data_15_4, 
      ordered_img_data_15_3=>ordered_img_data_15_3, ordered_img_data_15_2=>
      ordered_img_data_15_2, ordered_img_data_15_1=>ordered_img_data_15_1, 
      ordered_img_data_15_0=>ordered_img_data_15_0, ordered_img_data_16_31=>
      ordered_img_data_16_31, ordered_img_data_16_30=>DANGLING(400), 
      ordered_img_data_16_29=>DANGLING(401), ordered_img_data_16_28=>
      DANGLING(402), ordered_img_data_16_27=>DANGLING(403), 
      ordered_img_data_16_26=>DANGLING(404), ordered_img_data_16_25=>
      DANGLING(405), ordered_img_data_16_24=>DANGLING(406), 
      ordered_img_data_16_23=>DANGLING(407), ordered_img_data_16_22=>
      DANGLING(408), ordered_img_data_16_21=>DANGLING(409), 
      ordered_img_data_16_20=>DANGLING(410), ordered_img_data_16_19=>
      DANGLING(411), ordered_img_data_16_18=>DANGLING(412), 
      ordered_img_data_16_17=>DANGLING(413), ordered_img_data_16_16=>
      DANGLING(414), ordered_img_data_16_15=>DANGLING(415), 
      ordered_img_data_16_14=>ordered_img_data_16_14, ordered_img_data_16_13
      =>ordered_img_data_16_13, ordered_img_data_16_12=>
      ordered_img_data_16_12, ordered_img_data_16_11=>ordered_img_data_16_11, 
      ordered_img_data_16_10=>ordered_img_data_16_10, ordered_img_data_16_9
      =>ordered_img_data_16_9, ordered_img_data_16_8=>ordered_img_data_16_8, 
      ordered_img_data_16_7=>ordered_img_data_16_7, ordered_img_data_16_6=>
      ordered_img_data_16_6, ordered_img_data_16_5=>ordered_img_data_16_5, 
      ordered_img_data_16_4=>ordered_img_data_16_4, ordered_img_data_16_3=>
      ordered_img_data_16_3, ordered_img_data_16_2=>ordered_img_data_16_2, 
      ordered_img_data_16_1=>ordered_img_data_16_1, ordered_img_data_16_0=>
      ordered_img_data_16_0, ordered_img_data_17_31=>ordered_img_data_17_31, 
      ordered_img_data_17_30=>DANGLING(416), ordered_img_data_17_29=>
      DANGLING(417), ordered_img_data_17_28=>DANGLING(418), 
      ordered_img_data_17_27=>DANGLING(419), ordered_img_data_17_26=>
      DANGLING(420), ordered_img_data_17_25=>DANGLING(421), 
      ordered_img_data_17_24=>DANGLING(422), ordered_img_data_17_23=>
      DANGLING(423), ordered_img_data_17_22=>DANGLING(424), 
      ordered_img_data_17_21=>DANGLING(425), ordered_img_data_17_20=>
      DANGLING(426), ordered_img_data_17_19=>DANGLING(427), 
      ordered_img_data_17_18=>DANGLING(428), ordered_img_data_17_17=>
      DANGLING(429), ordered_img_data_17_16=>DANGLING(430), 
      ordered_img_data_17_15=>DANGLING(431), ordered_img_data_17_14=>
      ordered_img_data_17_14, ordered_img_data_17_13=>ordered_img_data_17_13, 
      ordered_img_data_17_12=>ordered_img_data_17_12, ordered_img_data_17_11
      =>ordered_img_data_17_11, ordered_img_data_17_10=>
      ordered_img_data_17_10, ordered_img_data_17_9=>ordered_img_data_17_9, 
      ordered_img_data_17_8=>ordered_img_data_17_8, ordered_img_data_17_7=>
      ordered_img_data_17_7, ordered_img_data_17_6=>ordered_img_data_17_6, 
      ordered_img_data_17_5=>ordered_img_data_17_5, ordered_img_data_17_4=>
      ordered_img_data_17_4, ordered_img_data_17_3=>ordered_img_data_17_3, 
      ordered_img_data_17_2=>ordered_img_data_17_2, ordered_img_data_17_1=>
      ordered_img_data_17_1, ordered_img_data_17_0=>ordered_img_data_17_0, 
      ordered_img_data_18_31=>DANGLING(432), ordered_img_data_18_30=>
      DANGLING(433), ordered_img_data_18_29=>DANGLING(434), 
      ordered_img_data_18_28=>DANGLING(435), ordered_img_data_18_27=>
      DANGLING(436), ordered_img_data_18_26=>DANGLING(437), 
      ordered_img_data_18_25=>DANGLING(438), ordered_img_data_18_24=>
      DANGLING(439), ordered_img_data_18_23=>DANGLING(440), 
      ordered_img_data_18_22=>DANGLING(441), ordered_img_data_18_21=>
      DANGLING(442), ordered_img_data_18_20=>DANGLING(443), 
      ordered_img_data_18_19=>DANGLING(444), ordered_img_data_18_18=>
      DANGLING(445), ordered_img_data_18_17=>DANGLING(446), 
      ordered_img_data_18_16=>DANGLING(447), ordered_img_data_18_15=>
      DANGLING(448), ordered_img_data_18_14=>DANGLING(449), 
      ordered_img_data_18_13=>DANGLING(450), ordered_img_data_18_12=>
      DANGLING(451), ordered_img_data_18_11=>DANGLING(452), 
      ordered_img_data_18_10=>DANGLING(453), ordered_img_data_18_9=>DANGLING
      (454), ordered_img_data_18_8=>DANGLING(455), ordered_img_data_18_7=>
      DANGLING(456), ordered_img_data_18_6=>DANGLING(457), 
      ordered_img_data_18_5=>DANGLING(458), ordered_img_data_18_4=>DANGLING(
      459), ordered_img_data_18_3=>DANGLING(460), ordered_img_data_18_2=>
      DANGLING(461), ordered_img_data_18_1=>DANGLING(462), 
      ordered_img_data_18_0=>DANGLING(463), ordered_img_data_19_31=>DANGLING
      (464), ordered_img_data_19_30=>DANGLING(465), ordered_img_data_19_29=>
      DANGLING(466), ordered_img_data_19_28=>DANGLING(467), 
      ordered_img_data_19_27=>DANGLING(468), ordered_img_data_19_26=>
      DANGLING(469), ordered_img_data_19_25=>DANGLING(470), 
      ordered_img_data_19_24=>DANGLING(471), ordered_img_data_19_23=>
      DANGLING(472), ordered_img_data_19_22=>DANGLING(473), 
      ordered_img_data_19_21=>DANGLING(474), ordered_img_data_19_20=>
      DANGLING(475), ordered_img_data_19_19=>DANGLING(476), 
      ordered_img_data_19_18=>DANGLING(477), ordered_img_data_19_17=>
      DANGLING(478), ordered_img_data_19_16=>DANGLING(479), 
      ordered_img_data_19_15=>DANGLING(480), ordered_img_data_19_14=>
      DANGLING(481), ordered_img_data_19_13=>DANGLING(482), 
      ordered_img_data_19_12=>DANGLING(483), ordered_img_data_19_11=>
      DANGLING(484), ordered_img_data_19_10=>DANGLING(485), 
      ordered_img_data_19_9=>DANGLING(486), ordered_img_data_19_8=>DANGLING(
      487), ordered_img_data_19_7=>DANGLING(488), ordered_img_data_19_6=>
      DANGLING(489), ordered_img_data_19_5=>DANGLING(490), 
      ordered_img_data_19_4=>DANGLING(491), ordered_img_data_19_3=>DANGLING(
      492), ordered_img_data_19_2=>DANGLING(493), ordered_img_data_19_1=>
      DANGLING(494), ordered_img_data_19_0=>DANGLING(495), 
      ordered_img_data_20_31=>DANGLING(496), ordered_img_data_20_30=>
      DANGLING(497), ordered_img_data_20_29=>DANGLING(498), 
      ordered_img_data_20_28=>DANGLING(499), ordered_img_data_20_27=>
      DANGLING(500), ordered_img_data_20_26=>DANGLING(501), 
      ordered_img_data_20_25=>DANGLING(502), ordered_img_data_20_24=>
      DANGLING(503), ordered_img_data_20_23=>DANGLING(504), 
      ordered_img_data_20_22=>DANGLING(505), ordered_img_data_20_21=>
      DANGLING(506), ordered_img_data_20_20=>DANGLING(507), 
      ordered_img_data_20_19=>DANGLING(508), ordered_img_data_20_18=>
      DANGLING(509), ordered_img_data_20_17=>DANGLING(510), 
      ordered_img_data_20_16=>DANGLING(511), ordered_img_data_20_15=>
      DANGLING(512), ordered_img_data_20_14=>DANGLING(513), 
      ordered_img_data_20_13=>DANGLING(514), ordered_img_data_20_12=>
      DANGLING(515), ordered_img_data_20_11=>DANGLING(516), 
      ordered_img_data_20_10=>DANGLING(517), ordered_img_data_20_9=>DANGLING
      (518), ordered_img_data_20_8=>DANGLING(519), ordered_img_data_20_7=>
      DANGLING(520), ordered_img_data_20_6=>DANGLING(521), 
      ordered_img_data_20_5=>DANGLING(522), ordered_img_data_20_4=>DANGLING(
      523), ordered_img_data_20_3=>DANGLING(524), ordered_img_data_20_2=>
      DANGLING(525), ordered_img_data_20_1=>DANGLING(526), 
      ordered_img_data_20_0=>DANGLING(527), ordered_img_data_21_31=>DANGLING
      (528), ordered_img_data_21_30=>DANGLING(529), ordered_img_data_21_29=>
      DANGLING(530), ordered_img_data_21_28=>DANGLING(531), 
      ordered_img_data_21_27=>DANGLING(532), ordered_img_data_21_26=>
      DANGLING(533), ordered_img_data_21_25=>DANGLING(534), 
      ordered_img_data_21_24=>DANGLING(535), ordered_img_data_21_23=>
      DANGLING(536), ordered_img_data_21_22=>DANGLING(537), 
      ordered_img_data_21_21=>DANGLING(538), ordered_img_data_21_20=>
      DANGLING(539), ordered_img_data_21_19=>DANGLING(540), 
      ordered_img_data_21_18=>DANGLING(541), ordered_img_data_21_17=>
      DANGLING(542), ordered_img_data_21_16=>DANGLING(543), 
      ordered_img_data_21_15=>DANGLING(544), ordered_img_data_21_14=>
      DANGLING(545), ordered_img_data_21_13=>DANGLING(546), 
      ordered_img_data_21_12=>DANGLING(547), ordered_img_data_21_11=>
      DANGLING(548), ordered_img_data_21_10=>DANGLING(549), 
      ordered_img_data_21_9=>DANGLING(550), ordered_img_data_21_8=>DANGLING(
      551), ordered_img_data_21_7=>DANGLING(552), ordered_img_data_21_6=>
      DANGLING(553), ordered_img_data_21_5=>DANGLING(554), 
      ordered_img_data_21_4=>DANGLING(555), ordered_img_data_21_3=>DANGLING(
      556), ordered_img_data_21_2=>DANGLING(557), ordered_img_data_21_1=>
      DANGLING(558), ordered_img_data_21_0=>DANGLING(559), 
      ordered_img_data_22_31=>DANGLING(560), ordered_img_data_22_30=>
      DANGLING(561), ordered_img_data_22_29=>DANGLING(562), 
      ordered_img_data_22_28=>DANGLING(563), ordered_img_data_22_27=>
      DANGLING(564), ordered_img_data_22_26=>DANGLING(565), 
      ordered_img_data_22_25=>DANGLING(566), ordered_img_data_22_24=>
      DANGLING(567), ordered_img_data_22_23=>DANGLING(568), 
      ordered_img_data_22_22=>DANGLING(569), ordered_img_data_22_21=>
      DANGLING(570), ordered_img_data_22_20=>DANGLING(571), 
      ordered_img_data_22_19=>DANGLING(572), ordered_img_data_22_18=>
      DANGLING(573), ordered_img_data_22_17=>DANGLING(574), 
      ordered_img_data_22_16=>DANGLING(575), ordered_img_data_22_15=>
      DANGLING(576), ordered_img_data_22_14=>DANGLING(577), 
      ordered_img_data_22_13=>DANGLING(578), ordered_img_data_22_12=>
      DANGLING(579), ordered_img_data_22_11=>DANGLING(580), 
      ordered_img_data_22_10=>DANGLING(581), ordered_img_data_22_9=>DANGLING
      (582), ordered_img_data_22_8=>DANGLING(583), ordered_img_data_22_7=>
      DANGLING(584), ordered_img_data_22_6=>DANGLING(585), 
      ordered_img_data_22_5=>DANGLING(586), ordered_img_data_22_4=>DANGLING(
      587), ordered_img_data_22_3=>DANGLING(588), ordered_img_data_22_2=>
      DANGLING(589), ordered_img_data_22_1=>DANGLING(590), 
      ordered_img_data_22_0=>DANGLING(591), ordered_img_data_23_31=>DANGLING
      (592), ordered_img_data_23_30=>DANGLING(593), ordered_img_data_23_29=>
      DANGLING(594), ordered_img_data_23_28=>DANGLING(595), 
      ordered_img_data_23_27=>DANGLING(596), ordered_img_data_23_26=>
      DANGLING(597), ordered_img_data_23_25=>DANGLING(598), 
      ordered_img_data_23_24=>DANGLING(599), ordered_img_data_23_23=>
      DANGLING(600), ordered_img_data_23_22=>DANGLING(601), 
      ordered_img_data_23_21=>DANGLING(602), ordered_img_data_23_20=>
      DANGLING(603), ordered_img_data_23_19=>DANGLING(604), 
      ordered_img_data_23_18=>DANGLING(605), ordered_img_data_23_17=>
      DANGLING(606), ordered_img_data_23_16=>DANGLING(607), 
      ordered_img_data_23_15=>DANGLING(608), ordered_img_data_23_14=>
      DANGLING(609), ordered_img_data_23_13=>DANGLING(610), 
      ordered_img_data_23_12=>DANGLING(611), ordered_img_data_23_11=>
      DANGLING(612), ordered_img_data_23_10=>DANGLING(613), 
      ordered_img_data_23_9=>DANGLING(614), ordered_img_data_23_8=>DANGLING(
      615), ordered_img_data_23_7=>DANGLING(616), ordered_img_data_23_6=>
      DANGLING(617), ordered_img_data_23_5=>DANGLING(618), 
      ordered_img_data_23_4=>DANGLING(619), ordered_img_data_23_3=>DANGLING(
      620), ordered_img_data_23_2=>DANGLING(621), ordered_img_data_23_1=>
      DANGLING(622), ordered_img_data_23_0=>DANGLING(623), 
      ordered_img_data_24_31=>DANGLING(624), ordered_img_data_24_30=>
      DANGLING(625), ordered_img_data_24_29=>DANGLING(626), 
      ordered_img_data_24_28=>DANGLING(627), ordered_img_data_24_27=>
      DANGLING(628), ordered_img_data_24_26=>DANGLING(629), 
      ordered_img_data_24_25=>DANGLING(630), ordered_img_data_24_24=>
      DANGLING(631), ordered_img_data_24_23=>DANGLING(632), 
      ordered_img_data_24_22=>DANGLING(633), ordered_img_data_24_21=>
      DANGLING(634), ordered_img_data_24_20=>DANGLING(635), 
      ordered_img_data_24_19=>DANGLING(636), ordered_img_data_24_18=>
      DANGLING(637), ordered_img_data_24_17=>DANGLING(638), 
      ordered_img_data_24_16=>DANGLING(639), ordered_img_data_24_15=>
      DANGLING(640), ordered_img_data_24_14=>DANGLING(641), 
      ordered_img_data_24_13=>DANGLING(642), ordered_img_data_24_12=>
      DANGLING(643), ordered_img_data_24_11=>DANGLING(644), 
      ordered_img_data_24_10=>DANGLING(645), ordered_img_data_24_9=>DANGLING
      (646), ordered_img_data_24_8=>DANGLING(647), ordered_img_data_24_7=>
      DANGLING(648), ordered_img_data_24_6=>DANGLING(649), 
      ordered_img_data_24_5=>DANGLING(650), ordered_img_data_24_4=>DANGLING(
      651), ordered_img_data_24_3=>DANGLING(652), ordered_img_data_24_2=>
      DANGLING(653), ordered_img_data_24_1=>DANGLING(654), 
      ordered_img_data_24_0=>DANGLING(655), ordered_filter_data_0_31=>
      DANGLING(656), ordered_filter_data_0_30=>DANGLING(657), 
      ordered_filter_data_0_29=>DANGLING(658), ordered_filter_data_0_28=>
      DANGLING(659), ordered_filter_data_0_27=>DANGLING(660), 
      ordered_filter_data_0_26=>DANGLING(661), ordered_filter_data_0_25=>
      DANGLING(662), ordered_filter_data_0_24=>DANGLING(663), 
      ordered_filter_data_0_23=>DANGLING(664), ordered_filter_data_0_22=>
      DANGLING(665), ordered_filter_data_0_21=>DANGLING(666), 
      ordered_filter_data_0_20=>DANGLING(667), ordered_filter_data_0_19=>
      DANGLING(668), ordered_filter_data_0_18=>DANGLING(669), 
      ordered_filter_data_0_17=>DANGLING(670), ordered_filter_data_0_16=>
      DANGLING(671), ordered_filter_data_0_15=>DANGLING(672), 
      ordered_filter_data_0_14=>DANGLING(673), ordered_filter_data_0_13=>
      DANGLING(674), ordered_filter_data_0_12=>DANGLING(675), 
      ordered_filter_data_0_11=>DANGLING(676), ordered_filter_data_0_10=>
      DANGLING(677), ordered_filter_data_0_9=>DANGLING(678), 
      ordered_filter_data_0_8=>DANGLING(679), ordered_filter_data_0_7=>
      DANGLING(680), ordered_filter_data_0_6=>DANGLING(681), 
      ordered_filter_data_0_5=>DANGLING(682), ordered_filter_data_0_4=>
      DANGLING(683), ordered_filter_data_0_3=>DANGLING(684), 
      ordered_filter_data_0_2=>DANGLING(685), ordered_filter_data_0_1=>
      DANGLING(686), ordered_filter_data_0_0=>DANGLING(687), 
      ordered_filter_data_1_31=>DANGLING(688), ordered_filter_data_1_30=>
      DANGLING(689), ordered_filter_data_1_29=>DANGLING(690), 
      ordered_filter_data_1_28=>DANGLING(691), ordered_filter_data_1_27=>
      DANGLING(692), ordered_filter_data_1_26=>DANGLING(693), 
      ordered_filter_data_1_25=>DANGLING(694), ordered_filter_data_1_24=>
      DANGLING(695), ordered_filter_data_1_23=>DANGLING(696), 
      ordered_filter_data_1_22=>DANGLING(697), ordered_filter_data_1_21=>
      DANGLING(698), ordered_filter_data_1_20=>DANGLING(699), 
      ordered_filter_data_1_19=>DANGLING(700), ordered_filter_data_1_18=>
      DANGLING(701), ordered_filter_data_1_17=>DANGLING(702), 
      ordered_filter_data_1_16=>DANGLING(703), ordered_filter_data_1_15=>
      DANGLING(704), ordered_filter_data_1_14=>DANGLING(705), 
      ordered_filter_data_1_13=>DANGLING(706), ordered_filter_data_1_12=>
      DANGLING(707), ordered_filter_data_1_11=>DANGLING(708), 
      ordered_filter_data_1_10=>DANGLING(709), ordered_filter_data_1_9=>
      DANGLING(710), ordered_filter_data_1_8=>DANGLING(711), 
      ordered_filter_data_1_7=>DANGLING(712), ordered_filter_data_1_6=>
      DANGLING(713), ordered_filter_data_1_5=>DANGLING(714), 
      ordered_filter_data_1_4=>DANGLING(715), ordered_filter_data_1_3=>
      DANGLING(716), ordered_filter_data_1_2=>DANGLING(717), 
      ordered_filter_data_1_1=>DANGLING(718), ordered_filter_data_1_0=>
      DANGLING(719), ordered_filter_data_2_31=>DANGLING(720), 
      ordered_filter_data_2_30=>DANGLING(721), ordered_filter_data_2_29=>
      DANGLING(722), ordered_filter_data_2_28=>DANGLING(723), 
      ordered_filter_data_2_27=>DANGLING(724), ordered_filter_data_2_26=>
      DANGLING(725), ordered_filter_data_2_25=>DANGLING(726), 
      ordered_filter_data_2_24=>DANGLING(727), ordered_filter_data_2_23=>
      DANGLING(728), ordered_filter_data_2_22=>DANGLING(729), 
      ordered_filter_data_2_21=>DANGLING(730), ordered_filter_data_2_20=>
      DANGLING(731), ordered_filter_data_2_19=>DANGLING(732), 
      ordered_filter_data_2_18=>DANGLING(733), ordered_filter_data_2_17=>
      DANGLING(734), ordered_filter_data_2_16=>DANGLING(735), 
      ordered_filter_data_2_15=>DANGLING(736), ordered_filter_data_2_14=>
      DANGLING(737), ordered_filter_data_2_13=>DANGLING(738), 
      ordered_filter_data_2_12=>DANGLING(739), ordered_filter_data_2_11=>
      DANGLING(740), ordered_filter_data_2_10=>DANGLING(741), 
      ordered_filter_data_2_9=>DANGLING(742), ordered_filter_data_2_8=>
      DANGLING(743), ordered_filter_data_2_7=>DANGLING(744), 
      ordered_filter_data_2_6=>DANGLING(745), ordered_filter_data_2_5=>
      DANGLING(746), ordered_filter_data_2_4=>DANGLING(747), 
      ordered_filter_data_2_3=>DANGLING(748), ordered_filter_data_2_2=>
      DANGLING(749), ordered_filter_data_2_1=>DANGLING(750), 
      ordered_filter_data_2_0=>DANGLING(751), ordered_filter_data_3_31=>
      DANGLING(752), ordered_filter_data_3_30=>DANGLING(753), 
      ordered_filter_data_3_29=>DANGLING(754), ordered_filter_data_3_28=>
      DANGLING(755), ordered_filter_data_3_27=>DANGLING(756), 
      ordered_filter_data_3_26=>DANGLING(757), ordered_filter_data_3_25=>
      DANGLING(758), ordered_filter_data_3_24=>DANGLING(759), 
      ordered_filter_data_3_23=>DANGLING(760), ordered_filter_data_3_22=>
      DANGLING(761), ordered_filter_data_3_21=>DANGLING(762), 
      ordered_filter_data_3_20=>DANGLING(763), ordered_filter_data_3_19=>
      DANGLING(764), ordered_filter_data_3_18=>DANGLING(765), 
      ordered_filter_data_3_17=>DANGLING(766), ordered_filter_data_3_16=>
      DANGLING(767), ordered_filter_data_3_15=>ordered_filter_data_3_15, 
      ordered_filter_data_3_14=>ordered_filter_data_3_14, 
      ordered_filter_data_3_13=>ordered_filter_data_3_13, 
      ordered_filter_data_3_12=>ordered_filter_data_3_12, 
      ordered_filter_data_3_11=>ordered_filter_data_3_11, 
      ordered_filter_data_3_10=>ordered_filter_data_3_10, 
      ordered_filter_data_3_9=>ordered_filter_data_3_9, 
      ordered_filter_data_3_8=>ordered_filter_data_3_8, 
      ordered_filter_data_3_7=>ordered_filter_data_3_7, 
      ordered_filter_data_3_6=>ordered_filter_data_3_6, 
      ordered_filter_data_3_5=>ordered_filter_data_3_5, 
      ordered_filter_data_3_4=>ordered_filter_data_3_4, 
      ordered_filter_data_3_3=>ordered_filter_data_3_3, 
      ordered_filter_data_3_2=>ordered_filter_data_3_2, 
      ordered_filter_data_3_1=>ordered_filter_data_3_1, 
      ordered_filter_data_3_0=>ordered_filter_data_3_0, 
      ordered_filter_data_4_31=>DANGLING(768), ordered_filter_data_4_30=>
      DANGLING(769), ordered_filter_data_4_29=>DANGLING(770), 
      ordered_filter_data_4_28=>DANGLING(771), ordered_filter_data_4_27=>
      DANGLING(772), ordered_filter_data_4_26=>DANGLING(773), 
      ordered_filter_data_4_25=>DANGLING(774), ordered_filter_data_4_24=>
      DANGLING(775), ordered_filter_data_4_23=>DANGLING(776), 
      ordered_filter_data_4_22=>DANGLING(777), ordered_filter_data_4_21=>
      DANGLING(778), ordered_filter_data_4_20=>DANGLING(779), 
      ordered_filter_data_4_19=>DANGLING(780), ordered_filter_data_4_18=>
      DANGLING(781), ordered_filter_data_4_17=>DANGLING(782), 
      ordered_filter_data_4_16=>DANGLING(783), ordered_filter_data_4_15=>
      ordered_filter_data_4_15, ordered_filter_data_4_14=>
      ordered_filter_data_4_14, ordered_filter_data_4_13=>
      ordered_filter_data_4_13, ordered_filter_data_4_12=>
      ordered_filter_data_4_12, ordered_filter_data_4_11=>
      ordered_filter_data_4_11, ordered_filter_data_4_10=>
      ordered_filter_data_4_10, ordered_filter_data_4_9=>
      ordered_filter_data_4_9, ordered_filter_data_4_8=>
      ordered_filter_data_4_8, ordered_filter_data_4_7=>
      ordered_filter_data_4_7, ordered_filter_data_4_6=>
      ordered_filter_data_4_6, ordered_filter_data_4_5=>
      ordered_filter_data_4_5, ordered_filter_data_4_4=>
      ordered_filter_data_4_4, ordered_filter_data_4_3=>
      ordered_filter_data_4_3, ordered_filter_data_4_2=>
      ordered_filter_data_4_2, ordered_filter_data_4_1=>
      ordered_filter_data_4_1, ordered_filter_data_4_0=>
      ordered_filter_data_4_0, ordered_filter_data_5_31=>DANGLING(784), 
      ordered_filter_data_5_30=>DANGLING(785), ordered_filter_data_5_29=>
      DANGLING(786), ordered_filter_data_5_28=>DANGLING(787), 
      ordered_filter_data_5_27=>DANGLING(788), ordered_filter_data_5_26=>
      DANGLING(789), ordered_filter_data_5_25=>DANGLING(790), 
      ordered_filter_data_5_24=>DANGLING(791), ordered_filter_data_5_23=>
      DANGLING(792), ordered_filter_data_5_22=>DANGLING(793), 
      ordered_filter_data_5_21=>DANGLING(794), ordered_filter_data_5_20=>
      DANGLING(795), ordered_filter_data_5_19=>DANGLING(796), 
      ordered_filter_data_5_18=>DANGLING(797), ordered_filter_data_5_17=>
      DANGLING(798), ordered_filter_data_5_16=>DANGLING(799), 
      ordered_filter_data_5_15=>ordered_filter_data_5_15, 
      ordered_filter_data_5_14=>ordered_filter_data_5_14, 
      ordered_filter_data_5_13=>ordered_filter_data_5_13, 
      ordered_filter_data_5_12=>ordered_filter_data_5_12, 
      ordered_filter_data_5_11=>ordered_filter_data_5_11, 
      ordered_filter_data_5_10=>ordered_filter_data_5_10, 
      ordered_filter_data_5_9=>ordered_filter_data_5_9, 
      ordered_filter_data_5_8=>ordered_filter_data_5_8, 
      ordered_filter_data_5_7=>ordered_filter_data_5_7, 
      ordered_filter_data_5_6=>ordered_filter_data_5_6, 
      ordered_filter_data_5_5=>ordered_filter_data_5_5, 
      ordered_filter_data_5_4=>ordered_filter_data_5_4, 
      ordered_filter_data_5_3=>ordered_filter_data_5_3, 
      ordered_filter_data_5_2=>ordered_filter_data_5_2, 
      ordered_filter_data_5_1=>ordered_filter_data_5_1, 
      ordered_filter_data_5_0=>ordered_filter_data_5_0, 
      ordered_filter_data_6_31=>DANGLING(800), ordered_filter_data_6_30=>
      DANGLING(801), ordered_filter_data_6_29=>DANGLING(802), 
      ordered_filter_data_6_28=>DANGLING(803), ordered_filter_data_6_27=>
      DANGLING(804), ordered_filter_data_6_26=>DANGLING(805), 
      ordered_filter_data_6_25=>DANGLING(806), ordered_filter_data_6_24=>
      DANGLING(807), ordered_filter_data_6_23=>DANGLING(808), 
      ordered_filter_data_6_22=>DANGLING(809), ordered_filter_data_6_21=>
      DANGLING(810), ordered_filter_data_6_20=>DANGLING(811), 
      ordered_filter_data_6_19=>DANGLING(812), ordered_filter_data_6_18=>
      DANGLING(813), ordered_filter_data_6_17=>DANGLING(814), 
      ordered_filter_data_6_16=>DANGLING(815), ordered_filter_data_6_15=>
      ordered_filter_data_6_15, ordered_filter_data_6_14=>
      ordered_filter_data_6_14, ordered_filter_data_6_13=>
      ordered_filter_data_6_13, ordered_filter_data_6_12=>
      ordered_filter_data_6_12, ordered_filter_data_6_11=>
      ordered_filter_data_6_11, ordered_filter_data_6_10=>
      ordered_filter_data_6_10, ordered_filter_data_6_9=>
      ordered_filter_data_6_9, ordered_filter_data_6_8=>
      ordered_filter_data_6_8, ordered_filter_data_6_7=>
      ordered_filter_data_6_7, ordered_filter_data_6_6=>
      ordered_filter_data_6_6, ordered_filter_data_6_5=>
      ordered_filter_data_6_5, ordered_filter_data_6_4=>
      ordered_filter_data_6_4, ordered_filter_data_6_3=>
      ordered_filter_data_6_3, ordered_filter_data_6_2=>
      ordered_filter_data_6_2, ordered_filter_data_6_1=>
      ordered_filter_data_6_1, ordered_filter_data_6_0=>
      ordered_filter_data_6_0, ordered_filter_data_7_31=>DANGLING(816), 
      ordered_filter_data_7_30=>DANGLING(817), ordered_filter_data_7_29=>
      DANGLING(818), ordered_filter_data_7_28=>DANGLING(819), 
      ordered_filter_data_7_27=>DANGLING(820), ordered_filter_data_7_26=>
      DANGLING(821), ordered_filter_data_7_25=>DANGLING(822), 
      ordered_filter_data_7_24=>DANGLING(823), ordered_filter_data_7_23=>
      DANGLING(824), ordered_filter_data_7_22=>DANGLING(825), 
      ordered_filter_data_7_21=>DANGLING(826), ordered_filter_data_7_20=>
      DANGLING(827), ordered_filter_data_7_19=>DANGLING(828), 
      ordered_filter_data_7_18=>DANGLING(829), ordered_filter_data_7_17=>
      DANGLING(830), ordered_filter_data_7_16=>DANGLING(831), 
      ordered_filter_data_7_15=>ordered_filter_data_7_15, 
      ordered_filter_data_7_14=>ordered_filter_data_7_14, 
      ordered_filter_data_7_13=>ordered_filter_data_7_13, 
      ordered_filter_data_7_12=>ordered_filter_data_7_12, 
      ordered_filter_data_7_11=>ordered_filter_data_7_11, 
      ordered_filter_data_7_10=>ordered_filter_data_7_10, 
      ordered_filter_data_7_9=>ordered_filter_data_7_9, 
      ordered_filter_data_7_8=>ordered_filter_data_7_8, 
      ordered_filter_data_7_7=>ordered_filter_data_7_7, 
      ordered_filter_data_7_6=>ordered_filter_data_7_6, 
      ordered_filter_data_7_5=>ordered_filter_data_7_5, 
      ordered_filter_data_7_4=>ordered_filter_data_7_4, 
      ordered_filter_data_7_3=>ordered_filter_data_7_3, 
      ordered_filter_data_7_2=>ordered_filter_data_7_2, 
      ordered_filter_data_7_1=>ordered_filter_data_7_1, 
      ordered_filter_data_7_0=>ordered_filter_data_7_0, 
      ordered_filter_data_8_31=>DANGLING(832), ordered_filter_data_8_30=>
      DANGLING(833), ordered_filter_data_8_29=>DANGLING(834), 
      ordered_filter_data_8_28=>DANGLING(835), ordered_filter_data_8_27=>
      DANGLING(836), ordered_filter_data_8_26=>DANGLING(837), 
      ordered_filter_data_8_25=>DANGLING(838), ordered_filter_data_8_24=>
      DANGLING(839), ordered_filter_data_8_23=>DANGLING(840), 
      ordered_filter_data_8_22=>DANGLING(841), ordered_filter_data_8_21=>
      DANGLING(842), ordered_filter_data_8_20=>DANGLING(843), 
      ordered_filter_data_8_19=>DANGLING(844), ordered_filter_data_8_18=>
      DANGLING(845), ordered_filter_data_8_17=>DANGLING(846), 
      ordered_filter_data_8_16=>DANGLING(847), ordered_filter_data_8_15=>
      ordered_filter_data_8_15, ordered_filter_data_8_14=>
      ordered_filter_data_8_14, ordered_filter_data_8_13=>
      ordered_filter_data_8_13, ordered_filter_data_8_12=>
      ordered_filter_data_8_12, ordered_filter_data_8_11=>
      ordered_filter_data_8_11, ordered_filter_data_8_10=>
      ordered_filter_data_8_10, ordered_filter_data_8_9=>
      ordered_filter_data_8_9, ordered_filter_data_8_8=>
      ordered_filter_data_8_8, ordered_filter_data_8_7=>
      ordered_filter_data_8_7, ordered_filter_data_8_6=>
      ordered_filter_data_8_6, ordered_filter_data_8_5=>
      ordered_filter_data_8_5, ordered_filter_data_8_4=>
      ordered_filter_data_8_4, ordered_filter_data_8_3=>
      ordered_filter_data_8_3, ordered_filter_data_8_2=>
      ordered_filter_data_8_2, ordered_filter_data_8_1=>
      ordered_filter_data_8_1, ordered_filter_data_8_0=>
      ordered_filter_data_8_0, ordered_filter_data_9_31=>DANGLING(848), 
      ordered_filter_data_9_30=>DANGLING(849), ordered_filter_data_9_29=>
      DANGLING(850), ordered_filter_data_9_28=>DANGLING(851), 
      ordered_filter_data_9_27=>DANGLING(852), ordered_filter_data_9_26=>
      DANGLING(853), ordered_filter_data_9_25=>DANGLING(854), 
      ordered_filter_data_9_24=>DANGLING(855), ordered_filter_data_9_23=>
      DANGLING(856), ordered_filter_data_9_22=>DANGLING(857), 
      ordered_filter_data_9_21=>DANGLING(858), ordered_filter_data_9_20=>
      DANGLING(859), ordered_filter_data_9_19=>DANGLING(860), 
      ordered_filter_data_9_18=>DANGLING(861), ordered_filter_data_9_17=>
      DANGLING(862), ordered_filter_data_9_16=>DANGLING(863), 
      ordered_filter_data_9_15=>ordered_filter_data_9_15, 
      ordered_filter_data_9_14=>ordered_filter_data_9_14, 
      ordered_filter_data_9_13=>ordered_filter_data_9_13, 
      ordered_filter_data_9_12=>ordered_filter_data_9_12, 
      ordered_filter_data_9_11=>ordered_filter_data_9_11, 
      ordered_filter_data_9_10=>ordered_filter_data_9_10, 
      ordered_filter_data_9_9=>ordered_filter_data_9_9, 
      ordered_filter_data_9_8=>ordered_filter_data_9_8, 
      ordered_filter_data_9_7=>ordered_filter_data_9_7, 
      ordered_filter_data_9_6=>ordered_filter_data_9_6, 
      ordered_filter_data_9_5=>ordered_filter_data_9_5, 
      ordered_filter_data_9_4=>ordered_filter_data_9_4, 
      ordered_filter_data_9_3=>ordered_filter_data_9_3, 
      ordered_filter_data_9_2=>ordered_filter_data_9_2, 
      ordered_filter_data_9_1=>ordered_filter_data_9_1, 
      ordered_filter_data_9_0=>ordered_filter_data_9_0, 
      ordered_filter_data_10_31=>DANGLING(864), ordered_filter_data_10_30=>
      DANGLING(865), ordered_filter_data_10_29=>DANGLING(866), 
      ordered_filter_data_10_28=>DANGLING(867), ordered_filter_data_10_27=>
      DANGLING(868), ordered_filter_data_10_26=>DANGLING(869), 
      ordered_filter_data_10_25=>DANGLING(870), ordered_filter_data_10_24=>
      DANGLING(871), ordered_filter_data_10_23=>DANGLING(872), 
      ordered_filter_data_10_22=>DANGLING(873), ordered_filter_data_10_21=>
      DANGLING(874), ordered_filter_data_10_20=>DANGLING(875), 
      ordered_filter_data_10_19=>DANGLING(876), ordered_filter_data_10_18=>
      DANGLING(877), ordered_filter_data_10_17=>DANGLING(878), 
      ordered_filter_data_10_16=>DANGLING(879), ordered_filter_data_10_15=>
      ordered_filter_data_10_15, ordered_filter_data_10_14=>
      ordered_filter_data_10_14, ordered_filter_data_10_13=>
      ordered_filter_data_10_13, ordered_filter_data_10_12=>
      ordered_filter_data_10_12, ordered_filter_data_10_11=>
      ordered_filter_data_10_11, ordered_filter_data_10_10=>
      ordered_filter_data_10_10, ordered_filter_data_10_9=>
      ordered_filter_data_10_9, ordered_filter_data_10_8=>
      ordered_filter_data_10_8, ordered_filter_data_10_7=>
      ordered_filter_data_10_7, ordered_filter_data_10_6=>
      ordered_filter_data_10_6, ordered_filter_data_10_5=>
      ordered_filter_data_10_5, ordered_filter_data_10_4=>
      ordered_filter_data_10_4, ordered_filter_data_10_3=>
      ordered_filter_data_10_3, ordered_filter_data_10_2=>
      ordered_filter_data_10_2, ordered_filter_data_10_1=>
      ordered_filter_data_10_1, ordered_filter_data_10_0=>
      ordered_filter_data_10_0, ordered_filter_data_11_31=>DANGLING(880), 
      ordered_filter_data_11_30=>DANGLING(881), ordered_filter_data_11_29=>
      DANGLING(882), ordered_filter_data_11_28=>DANGLING(883), 
      ordered_filter_data_11_27=>DANGLING(884), ordered_filter_data_11_26=>
      DANGLING(885), ordered_filter_data_11_25=>DANGLING(886), 
      ordered_filter_data_11_24=>DANGLING(887), ordered_filter_data_11_23=>
      DANGLING(888), ordered_filter_data_11_22=>DANGLING(889), 
      ordered_filter_data_11_21=>DANGLING(890), ordered_filter_data_11_20=>
      DANGLING(891), ordered_filter_data_11_19=>DANGLING(892), 
      ordered_filter_data_11_18=>DANGLING(893), ordered_filter_data_11_17=>
      DANGLING(894), ordered_filter_data_11_16=>DANGLING(895), 
      ordered_filter_data_11_15=>ordered_filter_data_11_15, 
      ordered_filter_data_11_14=>ordered_filter_data_11_14, 
      ordered_filter_data_11_13=>ordered_filter_data_11_13, 
      ordered_filter_data_11_12=>ordered_filter_data_11_12, 
      ordered_filter_data_11_11=>ordered_filter_data_11_11, 
      ordered_filter_data_11_10=>ordered_filter_data_11_10, 
      ordered_filter_data_11_9=>ordered_filter_data_11_9, 
      ordered_filter_data_11_8=>ordered_filter_data_11_8, 
      ordered_filter_data_11_7=>ordered_filter_data_11_7, 
      ordered_filter_data_11_6=>ordered_filter_data_11_6, 
      ordered_filter_data_11_5=>ordered_filter_data_11_5, 
      ordered_filter_data_11_4=>ordered_filter_data_11_4, 
      ordered_filter_data_11_3=>ordered_filter_data_11_3, 
      ordered_filter_data_11_2=>ordered_filter_data_11_2, 
      ordered_filter_data_11_1=>ordered_filter_data_11_1, 
      ordered_filter_data_11_0=>ordered_filter_data_11_0, 
      ordered_filter_data_12_31=>DANGLING(896), ordered_filter_data_12_30=>
      DANGLING(897), ordered_filter_data_12_29=>DANGLING(898), 
      ordered_filter_data_12_28=>DANGLING(899), ordered_filter_data_12_27=>
      DANGLING(900), ordered_filter_data_12_26=>DANGLING(901), 
      ordered_filter_data_12_25=>DANGLING(902), ordered_filter_data_12_24=>
      DANGLING(903), ordered_filter_data_12_23=>DANGLING(904), 
      ordered_filter_data_12_22=>DANGLING(905), ordered_filter_data_12_21=>
      DANGLING(906), ordered_filter_data_12_20=>DANGLING(907), 
      ordered_filter_data_12_19=>DANGLING(908), ordered_filter_data_12_18=>
      DANGLING(909), ordered_filter_data_12_17=>DANGLING(910), 
      ordered_filter_data_12_16=>DANGLING(911), ordered_filter_data_12_15=>
      ordered_filter_data_12_15, ordered_filter_data_12_14=>
      ordered_filter_data_12_14, ordered_filter_data_12_13=>
      ordered_filter_data_12_13, ordered_filter_data_12_12=>
      ordered_filter_data_12_12, ordered_filter_data_12_11=>
      ordered_filter_data_12_11, ordered_filter_data_12_10=>
      ordered_filter_data_12_10, ordered_filter_data_12_9=>
      ordered_filter_data_12_9, ordered_filter_data_12_8=>
      ordered_filter_data_12_8, ordered_filter_data_12_7=>
      ordered_filter_data_12_7, ordered_filter_data_12_6=>
      ordered_filter_data_12_6, ordered_filter_data_12_5=>
      ordered_filter_data_12_5, ordered_filter_data_12_4=>
      ordered_filter_data_12_4, ordered_filter_data_12_3=>
      ordered_filter_data_12_3, ordered_filter_data_12_2=>
      ordered_filter_data_12_2, ordered_filter_data_12_1=>
      ordered_filter_data_12_1, ordered_filter_data_12_0=>
      ordered_filter_data_12_0, ordered_filter_data_13_31=>DANGLING(912), 
      ordered_filter_data_13_30=>DANGLING(913), ordered_filter_data_13_29=>
      DANGLING(914), ordered_filter_data_13_28=>DANGLING(915), 
      ordered_filter_data_13_27=>DANGLING(916), ordered_filter_data_13_26=>
      DANGLING(917), ordered_filter_data_13_25=>DANGLING(918), 
      ordered_filter_data_13_24=>DANGLING(919), ordered_filter_data_13_23=>
      DANGLING(920), ordered_filter_data_13_22=>DANGLING(921), 
      ordered_filter_data_13_21=>DANGLING(922), ordered_filter_data_13_20=>
      DANGLING(923), ordered_filter_data_13_19=>DANGLING(924), 
      ordered_filter_data_13_18=>DANGLING(925), ordered_filter_data_13_17=>
      DANGLING(926), ordered_filter_data_13_16=>DANGLING(927), 
      ordered_filter_data_13_15=>ordered_filter_data_13_15, 
      ordered_filter_data_13_14=>ordered_filter_data_13_14, 
      ordered_filter_data_13_13=>ordered_filter_data_13_13, 
      ordered_filter_data_13_12=>ordered_filter_data_13_12, 
      ordered_filter_data_13_11=>ordered_filter_data_13_11, 
      ordered_filter_data_13_10=>ordered_filter_data_13_10, 
      ordered_filter_data_13_9=>ordered_filter_data_13_9, 
      ordered_filter_data_13_8=>ordered_filter_data_13_8, 
      ordered_filter_data_13_7=>ordered_filter_data_13_7, 
      ordered_filter_data_13_6=>ordered_filter_data_13_6, 
      ordered_filter_data_13_5=>ordered_filter_data_13_5, 
      ordered_filter_data_13_4=>ordered_filter_data_13_4, 
      ordered_filter_data_13_3=>ordered_filter_data_13_3, 
      ordered_filter_data_13_2=>ordered_filter_data_13_2, 
      ordered_filter_data_13_1=>ordered_filter_data_13_1, 
      ordered_filter_data_13_0=>ordered_filter_data_13_0, 
      ordered_filter_data_14_31=>DANGLING(928), ordered_filter_data_14_30=>
      DANGLING(929), ordered_filter_data_14_29=>DANGLING(930), 
      ordered_filter_data_14_28=>DANGLING(931), ordered_filter_data_14_27=>
      DANGLING(932), ordered_filter_data_14_26=>DANGLING(933), 
      ordered_filter_data_14_25=>DANGLING(934), ordered_filter_data_14_24=>
      DANGLING(935), ordered_filter_data_14_23=>DANGLING(936), 
      ordered_filter_data_14_22=>DANGLING(937), ordered_filter_data_14_21=>
      DANGLING(938), ordered_filter_data_14_20=>DANGLING(939), 
      ordered_filter_data_14_19=>DANGLING(940), ordered_filter_data_14_18=>
      DANGLING(941), ordered_filter_data_14_17=>DANGLING(942), 
      ordered_filter_data_14_16=>DANGLING(943), ordered_filter_data_14_15=>
      ordered_filter_data_14_15, ordered_filter_data_14_14=>
      ordered_filter_data_14_14, ordered_filter_data_14_13=>
      ordered_filter_data_14_13, ordered_filter_data_14_12=>
      ordered_filter_data_14_12, ordered_filter_data_14_11=>
      ordered_filter_data_14_11, ordered_filter_data_14_10=>
      ordered_filter_data_14_10, ordered_filter_data_14_9=>
      ordered_filter_data_14_9, ordered_filter_data_14_8=>
      ordered_filter_data_14_8, ordered_filter_data_14_7=>
      ordered_filter_data_14_7, ordered_filter_data_14_6=>
      ordered_filter_data_14_6, ordered_filter_data_14_5=>
      ordered_filter_data_14_5, ordered_filter_data_14_4=>
      ordered_filter_data_14_4, ordered_filter_data_14_3=>
      ordered_filter_data_14_3, ordered_filter_data_14_2=>
      ordered_filter_data_14_2, ordered_filter_data_14_1=>
      ordered_filter_data_14_1, ordered_filter_data_14_0=>
      ordered_filter_data_14_0, ordered_filter_data_15_31=>DANGLING(944), 
      ordered_filter_data_15_30=>DANGLING(945), ordered_filter_data_15_29=>
      DANGLING(946), ordered_filter_data_15_28=>DANGLING(947), 
      ordered_filter_data_15_27=>DANGLING(948), ordered_filter_data_15_26=>
      DANGLING(949), ordered_filter_data_15_25=>DANGLING(950), 
      ordered_filter_data_15_24=>DANGLING(951), ordered_filter_data_15_23=>
      DANGLING(952), ordered_filter_data_15_22=>DANGLING(953), 
      ordered_filter_data_15_21=>DANGLING(954), ordered_filter_data_15_20=>
      DANGLING(955), ordered_filter_data_15_19=>DANGLING(956), 
      ordered_filter_data_15_18=>DANGLING(957), ordered_filter_data_15_17=>
      DANGLING(958), ordered_filter_data_15_16=>DANGLING(959), 
      ordered_filter_data_15_15=>ordered_filter_data_15_15, 
      ordered_filter_data_15_14=>ordered_filter_data_15_14, 
      ordered_filter_data_15_13=>ordered_filter_data_15_13, 
      ordered_filter_data_15_12=>ordered_filter_data_15_12, 
      ordered_filter_data_15_11=>ordered_filter_data_15_11, 
      ordered_filter_data_15_10=>ordered_filter_data_15_10, 
      ordered_filter_data_15_9=>ordered_filter_data_15_9, 
      ordered_filter_data_15_8=>ordered_filter_data_15_8, 
      ordered_filter_data_15_7=>ordered_filter_data_15_7, 
      ordered_filter_data_15_6=>ordered_filter_data_15_6, 
      ordered_filter_data_15_5=>ordered_filter_data_15_5, 
      ordered_filter_data_15_4=>ordered_filter_data_15_4, 
      ordered_filter_data_15_3=>ordered_filter_data_15_3, 
      ordered_filter_data_15_2=>ordered_filter_data_15_2, 
      ordered_filter_data_15_1=>ordered_filter_data_15_1, 
      ordered_filter_data_15_0=>ordered_filter_data_15_0, 
      ordered_filter_data_16_31=>DANGLING(960), ordered_filter_data_16_30=>
      DANGLING(961), ordered_filter_data_16_29=>DANGLING(962), 
      ordered_filter_data_16_28=>DANGLING(963), ordered_filter_data_16_27=>
      DANGLING(964), ordered_filter_data_16_26=>DANGLING(965), 
      ordered_filter_data_16_25=>DANGLING(966), ordered_filter_data_16_24=>
      DANGLING(967), ordered_filter_data_16_23=>DANGLING(968), 
      ordered_filter_data_16_22=>DANGLING(969), ordered_filter_data_16_21=>
      DANGLING(970), ordered_filter_data_16_20=>DANGLING(971), 
      ordered_filter_data_16_19=>DANGLING(972), ordered_filter_data_16_18=>
      DANGLING(973), ordered_filter_data_16_17=>DANGLING(974), 
      ordered_filter_data_16_16=>DANGLING(975), ordered_filter_data_16_15=>
      ordered_filter_data_16_15, ordered_filter_data_16_14=>
      ordered_filter_data_16_14, ordered_filter_data_16_13=>
      ordered_filter_data_16_13, ordered_filter_data_16_12=>
      ordered_filter_data_16_12, ordered_filter_data_16_11=>
      ordered_filter_data_16_11, ordered_filter_data_16_10=>
      ordered_filter_data_16_10, ordered_filter_data_16_9=>
      ordered_filter_data_16_9, ordered_filter_data_16_8=>
      ordered_filter_data_16_8, ordered_filter_data_16_7=>
      ordered_filter_data_16_7, ordered_filter_data_16_6=>
      ordered_filter_data_16_6, ordered_filter_data_16_5=>
      ordered_filter_data_16_5, ordered_filter_data_16_4=>
      ordered_filter_data_16_4, ordered_filter_data_16_3=>
      ordered_filter_data_16_3, ordered_filter_data_16_2=>
      ordered_filter_data_16_2, ordered_filter_data_16_1=>
      ordered_filter_data_16_1, ordered_filter_data_16_0=>
      ordered_filter_data_16_0, ordered_filter_data_17_31=>DANGLING(976), 
      ordered_filter_data_17_30=>DANGLING(977), ordered_filter_data_17_29=>
      DANGLING(978), ordered_filter_data_17_28=>DANGLING(979), 
      ordered_filter_data_17_27=>DANGLING(980), ordered_filter_data_17_26=>
      DANGLING(981), ordered_filter_data_17_25=>DANGLING(982), 
      ordered_filter_data_17_24=>DANGLING(983), ordered_filter_data_17_23=>
      DANGLING(984), ordered_filter_data_17_22=>DANGLING(985), 
      ordered_filter_data_17_21=>DANGLING(986), ordered_filter_data_17_20=>
      DANGLING(987), ordered_filter_data_17_19=>DANGLING(988), 
      ordered_filter_data_17_18=>DANGLING(989), ordered_filter_data_17_17=>
      DANGLING(990), ordered_filter_data_17_16=>DANGLING(991), 
      ordered_filter_data_17_15=>ordered_filter_data_17_15, 
      ordered_filter_data_17_14=>ordered_filter_data_17_14, 
      ordered_filter_data_17_13=>ordered_filter_data_17_13, 
      ordered_filter_data_17_12=>ordered_filter_data_17_12, 
      ordered_filter_data_17_11=>ordered_filter_data_17_11, 
      ordered_filter_data_17_10=>ordered_filter_data_17_10, 
      ordered_filter_data_17_9=>ordered_filter_data_17_9, 
      ordered_filter_data_17_8=>ordered_filter_data_17_8, 
      ordered_filter_data_17_7=>ordered_filter_data_17_7, 
      ordered_filter_data_17_6=>ordered_filter_data_17_6, 
      ordered_filter_data_17_5=>ordered_filter_data_17_5, 
      ordered_filter_data_17_4=>ordered_filter_data_17_4, 
      ordered_filter_data_17_3=>ordered_filter_data_17_3, 
      ordered_filter_data_17_2=>ordered_filter_data_17_2, 
      ordered_filter_data_17_1=>ordered_filter_data_17_1, 
      ordered_filter_data_17_0=>ordered_filter_data_17_0, 
      ordered_filter_data_18_31=>DANGLING(992), ordered_filter_data_18_30=>
      DANGLING(993), ordered_filter_data_18_29=>DANGLING(994), 
      ordered_filter_data_18_28=>DANGLING(995), ordered_filter_data_18_27=>
      DANGLING(996), ordered_filter_data_18_26=>DANGLING(997), 
      ordered_filter_data_18_25=>DANGLING(998), ordered_filter_data_18_24=>
      DANGLING(999), ordered_filter_data_18_23=>DANGLING(1000), 
      ordered_filter_data_18_22=>DANGLING(1001), ordered_filter_data_18_21=>
      DANGLING(1002), ordered_filter_data_18_20=>DANGLING(1003), 
      ordered_filter_data_18_19=>DANGLING(1004), ordered_filter_data_18_18=>
      DANGLING(1005), ordered_filter_data_18_17=>DANGLING(1006), 
      ordered_filter_data_18_16=>DANGLING(1007), ordered_filter_data_18_15=>
      DANGLING(1008), ordered_filter_data_18_14=>DANGLING(1009), 
      ordered_filter_data_18_13=>DANGLING(1010), ordered_filter_data_18_12=>
      DANGLING(1011), ordered_filter_data_18_11=>DANGLING(1012), 
      ordered_filter_data_18_10=>DANGLING(1013), ordered_filter_data_18_9=>
      DANGLING(1014), ordered_filter_data_18_8=>DANGLING(1015), 
      ordered_filter_data_18_7=>DANGLING(1016), ordered_filter_data_18_6=>
      DANGLING(1017), ordered_filter_data_18_5=>DANGLING(1018), 
      ordered_filter_data_18_4=>DANGLING(1019), ordered_filter_data_18_3=>
      DANGLING(1020), ordered_filter_data_18_2=>DANGLING(1021), 
      ordered_filter_data_18_1=>DANGLING(1022), ordered_filter_data_18_0=>
      DANGLING(1023), ordered_filter_data_19_31=>DANGLING(1024), 
      ordered_filter_data_19_30=>DANGLING(1025), ordered_filter_data_19_29=>
      DANGLING(1026), ordered_filter_data_19_28=>DANGLING(1027), 
      ordered_filter_data_19_27=>DANGLING(1028), ordered_filter_data_19_26=>
      DANGLING(1029), ordered_filter_data_19_25=>DANGLING(1030), 
      ordered_filter_data_19_24=>DANGLING(1031), ordered_filter_data_19_23=>
      DANGLING(1032), ordered_filter_data_19_22=>DANGLING(1033), 
      ordered_filter_data_19_21=>DANGLING(1034), ordered_filter_data_19_20=>
      DANGLING(1035), ordered_filter_data_19_19=>DANGLING(1036), 
      ordered_filter_data_19_18=>DANGLING(1037), ordered_filter_data_19_17=>
      DANGLING(1038), ordered_filter_data_19_16=>DANGLING(1039), 
      ordered_filter_data_19_15=>DANGLING(1040), ordered_filter_data_19_14=>
      DANGLING(1041), ordered_filter_data_19_13=>DANGLING(1042), 
      ordered_filter_data_19_12=>DANGLING(1043), ordered_filter_data_19_11=>
      DANGLING(1044), ordered_filter_data_19_10=>DANGLING(1045), 
      ordered_filter_data_19_9=>DANGLING(1046), ordered_filter_data_19_8=>
      DANGLING(1047), ordered_filter_data_19_7=>DANGLING(1048), 
      ordered_filter_data_19_6=>DANGLING(1049), ordered_filter_data_19_5=>
      DANGLING(1050), ordered_filter_data_19_4=>DANGLING(1051), 
      ordered_filter_data_19_3=>DANGLING(1052), ordered_filter_data_19_2=>
      DANGLING(1053), ordered_filter_data_19_1=>DANGLING(1054), 
      ordered_filter_data_19_0=>DANGLING(1055), ordered_filter_data_20_31=>
      DANGLING(1056), ordered_filter_data_20_30=>DANGLING(1057), 
      ordered_filter_data_20_29=>DANGLING(1058), ordered_filter_data_20_28=>
      DANGLING(1059), ordered_filter_data_20_27=>DANGLING(1060), 
      ordered_filter_data_20_26=>DANGLING(1061), ordered_filter_data_20_25=>
      DANGLING(1062), ordered_filter_data_20_24=>DANGLING(1063), 
      ordered_filter_data_20_23=>DANGLING(1064), ordered_filter_data_20_22=>
      DANGLING(1065), ordered_filter_data_20_21=>DANGLING(1066), 
      ordered_filter_data_20_20=>DANGLING(1067), ordered_filter_data_20_19=>
      DANGLING(1068), ordered_filter_data_20_18=>DANGLING(1069), 
      ordered_filter_data_20_17=>DANGLING(1070), ordered_filter_data_20_16=>
      DANGLING(1071), ordered_filter_data_20_15=>DANGLING(1072), 
      ordered_filter_data_20_14=>DANGLING(1073), ordered_filter_data_20_13=>
      DANGLING(1074), ordered_filter_data_20_12=>DANGLING(1075), 
      ordered_filter_data_20_11=>DANGLING(1076), ordered_filter_data_20_10=>
      DANGLING(1077), ordered_filter_data_20_9=>DANGLING(1078), 
      ordered_filter_data_20_8=>DANGLING(1079), ordered_filter_data_20_7=>
      DANGLING(1080), ordered_filter_data_20_6=>DANGLING(1081), 
      ordered_filter_data_20_5=>DANGLING(1082), ordered_filter_data_20_4=>
      DANGLING(1083), ordered_filter_data_20_3=>DANGLING(1084), 
      ordered_filter_data_20_2=>DANGLING(1085), ordered_filter_data_20_1=>
      DANGLING(1086), ordered_filter_data_20_0=>DANGLING(1087), 
      ordered_filter_data_21_31=>DANGLING(1088), ordered_filter_data_21_30=>
      DANGLING(1089), ordered_filter_data_21_29=>DANGLING(1090), 
      ordered_filter_data_21_28=>DANGLING(1091), ordered_filter_data_21_27=>
      DANGLING(1092), ordered_filter_data_21_26=>DANGLING(1093), 
      ordered_filter_data_21_25=>DANGLING(1094), ordered_filter_data_21_24=>
      DANGLING(1095), ordered_filter_data_21_23=>DANGLING(1096), 
      ordered_filter_data_21_22=>DANGLING(1097), ordered_filter_data_21_21=>
      DANGLING(1098), ordered_filter_data_21_20=>DANGLING(1099), 
      ordered_filter_data_21_19=>DANGLING(1100), ordered_filter_data_21_18=>
      DANGLING(1101), ordered_filter_data_21_17=>DANGLING(1102), 
      ordered_filter_data_21_16=>DANGLING(1103), ordered_filter_data_21_15=>
      DANGLING(1104), ordered_filter_data_21_14=>DANGLING(1105), 
      ordered_filter_data_21_13=>DANGLING(1106), ordered_filter_data_21_12=>
      DANGLING(1107), ordered_filter_data_21_11=>DANGLING(1108), 
      ordered_filter_data_21_10=>DANGLING(1109), ordered_filter_data_21_9=>
      DANGLING(1110), ordered_filter_data_21_8=>DANGLING(1111), 
      ordered_filter_data_21_7=>DANGLING(1112), ordered_filter_data_21_6=>
      DANGLING(1113), ordered_filter_data_21_5=>DANGLING(1114), 
      ordered_filter_data_21_4=>DANGLING(1115), ordered_filter_data_21_3=>
      DANGLING(1116), ordered_filter_data_21_2=>DANGLING(1117), 
      ordered_filter_data_21_1=>DANGLING(1118), ordered_filter_data_21_0=>
      DANGLING(1119), ordered_filter_data_22_31=>DANGLING(1120), 
      ordered_filter_data_22_30=>DANGLING(1121), ordered_filter_data_22_29=>
      DANGLING(1122), ordered_filter_data_22_28=>DANGLING(1123), 
      ordered_filter_data_22_27=>DANGLING(1124), ordered_filter_data_22_26=>
      DANGLING(1125), ordered_filter_data_22_25=>DANGLING(1126), 
      ordered_filter_data_22_24=>DANGLING(1127), ordered_filter_data_22_23=>
      DANGLING(1128), ordered_filter_data_22_22=>DANGLING(1129), 
      ordered_filter_data_22_21=>DANGLING(1130), ordered_filter_data_22_20=>
      DANGLING(1131), ordered_filter_data_22_19=>DANGLING(1132), 
      ordered_filter_data_22_18=>DANGLING(1133), ordered_filter_data_22_17=>
      DANGLING(1134), ordered_filter_data_22_16=>DANGLING(1135), 
      ordered_filter_data_22_15=>DANGLING(1136), ordered_filter_data_22_14=>
      DANGLING(1137), ordered_filter_data_22_13=>DANGLING(1138), 
      ordered_filter_data_22_12=>DANGLING(1139), ordered_filter_data_22_11=>
      DANGLING(1140), ordered_filter_data_22_10=>DANGLING(1141), 
      ordered_filter_data_22_9=>DANGLING(1142), ordered_filter_data_22_8=>
      DANGLING(1143), ordered_filter_data_22_7=>DANGLING(1144), 
      ordered_filter_data_22_6=>DANGLING(1145), ordered_filter_data_22_5=>
      DANGLING(1146), ordered_filter_data_22_4=>DANGLING(1147), 
      ordered_filter_data_22_3=>DANGLING(1148), ordered_filter_data_22_2=>
      DANGLING(1149), ordered_filter_data_22_1=>DANGLING(1150), 
      ordered_filter_data_22_0=>DANGLING(1151), ordered_filter_data_23_31=>
      DANGLING(1152), ordered_filter_data_23_30=>DANGLING(1153), 
      ordered_filter_data_23_29=>DANGLING(1154), ordered_filter_data_23_28=>
      DANGLING(1155), ordered_filter_data_23_27=>DANGLING(1156), 
      ordered_filter_data_23_26=>DANGLING(1157), ordered_filter_data_23_25=>
      DANGLING(1158), ordered_filter_data_23_24=>DANGLING(1159), 
      ordered_filter_data_23_23=>DANGLING(1160), ordered_filter_data_23_22=>
      DANGLING(1161), ordered_filter_data_23_21=>DANGLING(1162), 
      ordered_filter_data_23_20=>DANGLING(1163), ordered_filter_data_23_19=>
      DANGLING(1164), ordered_filter_data_23_18=>DANGLING(1165), 
      ordered_filter_data_23_17=>DANGLING(1166), ordered_filter_data_23_16=>
      DANGLING(1167), ordered_filter_data_23_15=>DANGLING(1168), 
      ordered_filter_data_23_14=>DANGLING(1169), ordered_filter_data_23_13=>
      DANGLING(1170), ordered_filter_data_23_12=>DANGLING(1171), 
      ordered_filter_data_23_11=>DANGLING(1172), ordered_filter_data_23_10=>
      DANGLING(1173), ordered_filter_data_23_9=>DANGLING(1174), 
      ordered_filter_data_23_8=>DANGLING(1175), ordered_filter_data_23_7=>
      DANGLING(1176), ordered_filter_data_23_6=>DANGLING(1177), 
      ordered_filter_data_23_5=>DANGLING(1178), ordered_filter_data_23_4=>
      DANGLING(1179), ordered_filter_data_23_3=>DANGLING(1180), 
      ordered_filter_data_23_2=>DANGLING(1181), ordered_filter_data_23_1=>
      DANGLING(1182), ordered_filter_data_23_0=>DANGLING(1183), 
      ordered_filter_data_24_31=>DANGLING(1184), ordered_filter_data_24_30=>
      DANGLING(1185), ordered_filter_data_24_29=>DANGLING(1186), 
      ordered_filter_data_24_28=>DANGLING(1187), ordered_filter_data_24_27=>
      DANGLING(1188), ordered_filter_data_24_26=>DANGLING(1189), 
      ordered_filter_data_24_25=>DANGLING(1190), ordered_filter_data_24_24=>
      DANGLING(1191), ordered_filter_data_24_23=>DANGLING(1192), 
      ordered_filter_data_24_22=>DANGLING(1193), ordered_filter_data_24_21=>
      DANGLING(1194), ordered_filter_data_24_20=>DANGLING(1195), 
      ordered_filter_data_24_19=>DANGLING(1196), ordered_filter_data_24_18=>
      DANGLING(1197), ordered_filter_data_24_17=>DANGLING(1198), 
      ordered_filter_data_24_16=>DANGLING(1199), ordered_filter_data_24_15=>
      DANGLING(1200), ordered_filter_data_24_14=>DANGLING(1201), 
      ordered_filter_data_24_13=>DANGLING(1202), ordered_filter_data_24_12=>
      DANGLING(1203), ordered_filter_data_24_11=>DANGLING(1204), 
      ordered_filter_data_24_10=>DANGLING(1205), ordered_filter_data_24_9=>
      DANGLING(1206), ordered_filter_data_24_8=>DANGLING(1207), 
      ordered_filter_data_24_7=>DANGLING(1208), ordered_filter_data_24_6=>
      DANGLING(1209), ordered_filter_data_24_5=>DANGLING(1210), 
      ordered_filter_data_24_4=>DANGLING(1211), ordered_filter_data_24_3=>
      DANGLING(1212), ordered_filter_data_24_2=>DANGLING(1213), 
      ordered_filter_data_24_1=>DANGLING(1214), ordered_filter_data_24_0=>
      DANGLING(1215));
   merge_layer1_gen : MergeLayer port map ( d_arr_0_31=>d_arr_merge1_0_31, 
      d_arr_0_30=>d_arr_merge1_0_30, d_arr_0_29=>d_arr_merge1_0_29, 
      d_arr_0_28=>d_arr_merge1_0_28, d_arr_0_27=>d_arr_merge1_0_27, 
      d_arr_0_26=>d_arr_merge1_0_26, d_arr_0_25=>d_arr_merge1_0_25, 
      d_arr_0_24=>d_arr_merge1_0_24, d_arr_0_23=>d_arr_merge1_0_23, 
      d_arr_0_22=>d_arr_merge1_0_22, d_arr_0_21=>d_arr_merge1_0_21, 
      d_arr_0_20=>d_arr_merge1_0_20, d_arr_0_19=>d_arr_merge1_0_19, 
      d_arr_0_18=>d_arr_merge1_0_18, d_arr_0_17=>d_arr_merge1_0_17, 
      d_arr_0_16=>d_arr_merge1_0_16, d_arr_0_15=>d_arr_merge1_0_15, 
      d_arr_0_14=>d_arr_merge1_0_14, d_arr_0_13=>d_arr_merge1_0_13, 
      d_arr_0_12=>d_arr_merge1_0_12, d_arr_0_11=>d_arr_merge1_0_11, 
      d_arr_0_10=>d_arr_merge1_0_10, d_arr_0_9=>d_arr_merge1_0_9, d_arr_0_8
      =>d_arr_merge1_0_8, d_arr_0_7=>d_arr_merge1_0_7, d_arr_0_6=>
      d_arr_merge1_0_6, d_arr_0_5=>d_arr_merge1_0_5, d_arr_0_4=>
      d_arr_merge1_0_4, d_arr_0_3=>d_arr_merge1_0_3, d_arr_0_2=>
      d_arr_merge1_0_2, d_arr_0_1=>d_arr_merge1_0_1, d_arr_0_0=>
      d_arr_merge1_0_0, d_arr_1_31=>d_arr_merge1_1_31, d_arr_1_30=>
      d_arr_merge1_1_30, d_arr_1_29=>d_arr_merge1_1_29, d_arr_1_28=>
      d_arr_merge1_1_28, d_arr_1_27=>d_arr_merge1_1_27, d_arr_1_26=>
      d_arr_merge1_1_26, d_arr_1_25=>d_arr_merge1_1_25, d_arr_1_24=>
      d_arr_merge1_1_24, d_arr_1_23=>d_arr_merge1_1_23, d_arr_1_22=>
      d_arr_merge1_1_22, d_arr_1_21=>d_arr_merge1_1_21, d_arr_1_20=>
      d_arr_merge1_1_20, d_arr_1_19=>d_arr_merge1_1_19, d_arr_1_18=>
      d_arr_merge1_1_18, d_arr_1_17=>d_arr_merge1_1_17, d_arr_1_16=>
      d_arr_merge1_1_16, d_arr_1_15=>d_arr_merge1_1_15, d_arr_1_14=>
      d_arr_merge1_1_14, d_arr_1_13=>d_arr_merge1_1_13, d_arr_1_12=>
      d_arr_merge1_1_12, d_arr_1_11=>d_arr_merge1_1_11, d_arr_1_10=>
      d_arr_merge1_1_10, d_arr_1_9=>d_arr_merge1_1_9, d_arr_1_8=>
      d_arr_merge1_1_8, d_arr_1_7=>d_arr_merge1_1_7, d_arr_1_6=>
      d_arr_merge1_1_6, d_arr_1_5=>d_arr_merge1_1_5, d_arr_1_4=>
      d_arr_merge1_1_4, d_arr_1_3=>d_arr_merge1_1_3, d_arr_1_2=>
      d_arr_merge1_1_2, d_arr_1_1=>d_arr_merge1_1_1, d_arr_1_0=>
      d_arr_merge1_1_0, d_arr_2_31=>DANGLING(1216), d_arr_2_30=>DANGLING(
      1217), d_arr_2_29=>DANGLING(1218), d_arr_2_28=>DANGLING(1219), 
      d_arr_2_27=>DANGLING(1220), d_arr_2_26=>DANGLING(1221), d_arr_2_25=>
      DANGLING(1222), d_arr_2_24=>DANGLING(1223), d_arr_2_23=>DANGLING(1224), 
      d_arr_2_22=>DANGLING(1225), d_arr_2_21=>DANGLING(1226), d_arr_2_20=>
      DANGLING(1227), d_arr_2_19=>DANGLING(1228), d_arr_2_18=>DANGLING(1229), 
      d_arr_2_17=>DANGLING(1230), d_arr_2_16=>DANGLING(1231), d_arr_2_15=>
      DANGLING(1232), d_arr_2_14=>DANGLING(1233), d_arr_2_13=>DANGLING(1234), 
      d_arr_2_12=>DANGLING(1235), d_arr_2_11=>DANGLING(1236), d_arr_2_10=>
      DANGLING(1237), d_arr_2_9=>DANGLING(1238), d_arr_2_8=>DANGLING(1239), 
      d_arr_2_7=>DANGLING(1240), d_arr_2_6=>DANGLING(1241), d_arr_2_5=>
      DANGLING(1242), d_arr_2_4=>DANGLING(1243), d_arr_2_3=>DANGLING(1244), 
      d_arr_2_2=>DANGLING(1245), d_arr_2_1=>DANGLING(1246), d_arr_2_0=>
      DANGLING(1247), d_arr_3_31=>DANGLING(1248), d_arr_3_30=>DANGLING(1249), 
      d_arr_3_29=>DANGLING(1250), d_arr_3_28=>DANGLING(1251), d_arr_3_27=>
      DANGLING(1252), d_arr_3_26=>DANGLING(1253), d_arr_3_25=>DANGLING(1254), 
      d_arr_3_24=>DANGLING(1255), d_arr_3_23=>DANGLING(1256), d_arr_3_22=>
      DANGLING(1257), d_arr_3_21=>DANGLING(1258), d_arr_3_20=>DANGLING(1259), 
      d_arr_3_19=>DANGLING(1260), d_arr_3_18=>DANGLING(1261), d_arr_3_17=>
      DANGLING(1262), d_arr_3_16=>DANGLING(1263), d_arr_3_15=>DANGLING(1264), 
      d_arr_3_14=>DANGLING(1265), d_arr_3_13=>DANGLING(1266), d_arr_3_12=>
      DANGLING(1267), d_arr_3_11=>DANGLING(1268), d_arr_3_10=>DANGLING(1269), 
      d_arr_3_9=>DANGLING(1270), d_arr_3_8=>DANGLING(1271), d_arr_3_7=>
      DANGLING(1272), d_arr_3_6=>DANGLING(1273), d_arr_3_5=>DANGLING(1274), 
      d_arr_3_4=>DANGLING(1275), d_arr_3_3=>DANGLING(1276), d_arr_3_2=>
      DANGLING(1277), d_arr_3_1=>DANGLING(1278), d_arr_3_0=>DANGLING(1279), 
      d_arr_4_31=>DANGLING(1280), d_arr_4_30=>DANGLING(1281), d_arr_4_29=>
      DANGLING(1282), d_arr_4_28=>DANGLING(1283), d_arr_4_27=>DANGLING(1284), 
      d_arr_4_26=>DANGLING(1285), d_arr_4_25=>DANGLING(1286), d_arr_4_24=>
      DANGLING(1287), d_arr_4_23=>DANGLING(1288), d_arr_4_22=>DANGLING(1289), 
      d_arr_4_21=>DANGLING(1290), d_arr_4_20=>DANGLING(1291), d_arr_4_19=>
      DANGLING(1292), d_arr_4_18=>DANGLING(1293), d_arr_4_17=>DANGLING(1294), 
      d_arr_4_16=>DANGLING(1295), d_arr_4_15=>DANGLING(1296), d_arr_4_14=>
      DANGLING(1297), d_arr_4_13=>DANGLING(1298), d_arr_4_12=>DANGLING(1299), 
      d_arr_4_11=>DANGLING(1300), d_arr_4_10=>DANGLING(1301), d_arr_4_9=>
      DANGLING(1302), d_arr_4_8=>DANGLING(1303), d_arr_4_7=>DANGLING(1304), 
      d_arr_4_6=>DANGLING(1305), d_arr_4_5=>DANGLING(1306), d_arr_4_4=>
      DANGLING(1307), d_arr_4_3=>DANGLING(1308), d_arr_4_2=>DANGLING(1309), 
      d_arr_4_1=>DANGLING(1310), d_arr_4_0=>DANGLING(1311), d_arr_5_31=>
      DANGLING(1312), d_arr_5_30=>DANGLING(1313), d_arr_5_29=>DANGLING(1314), 
      d_arr_5_28=>DANGLING(1315), d_arr_5_27=>DANGLING(1316), d_arr_5_26=>
      DANGLING(1317), d_arr_5_25=>DANGLING(1318), d_arr_5_24=>DANGLING(1319), 
      d_arr_5_23=>DANGLING(1320), d_arr_5_22=>DANGLING(1321), d_arr_5_21=>
      DANGLING(1322), d_arr_5_20=>DANGLING(1323), d_arr_5_19=>DANGLING(1324), 
      d_arr_5_18=>DANGLING(1325), d_arr_5_17=>DANGLING(1326), d_arr_5_16=>
      DANGLING(1327), d_arr_5_15=>DANGLING(1328), d_arr_5_14=>DANGLING(1329), 
      d_arr_5_13=>DANGLING(1330), d_arr_5_12=>DANGLING(1331), d_arr_5_11=>
      DANGLING(1332), d_arr_5_10=>DANGLING(1333), d_arr_5_9=>DANGLING(1334), 
      d_arr_5_8=>DANGLING(1335), d_arr_5_7=>DANGLING(1336), d_arr_5_6=>
      DANGLING(1337), d_arr_5_5=>DANGLING(1338), d_arr_5_4=>DANGLING(1339), 
      d_arr_5_3=>DANGLING(1340), d_arr_5_2=>DANGLING(1341), d_arr_5_1=>
      DANGLING(1342), d_arr_5_0=>DANGLING(1343), d_arr_6_31=>DANGLING(1344), 
      d_arr_6_30=>DANGLING(1345), d_arr_6_29=>DANGLING(1346), d_arr_6_28=>
      DANGLING(1347), d_arr_6_27=>DANGLING(1348), d_arr_6_26=>DANGLING(1349), 
      d_arr_6_25=>DANGLING(1350), d_arr_6_24=>DANGLING(1351), d_arr_6_23=>
      DANGLING(1352), d_arr_6_22=>DANGLING(1353), d_arr_6_21=>DANGLING(1354), 
      d_arr_6_20=>DANGLING(1355), d_arr_6_19=>DANGLING(1356), d_arr_6_18=>
      DANGLING(1357), d_arr_6_17=>DANGLING(1358), d_arr_6_16=>DANGLING(1359), 
      d_arr_6_15=>DANGLING(1360), d_arr_6_14=>DANGLING(1361), d_arr_6_13=>
      DANGLING(1362), d_arr_6_12=>DANGLING(1363), d_arr_6_11=>DANGLING(1364), 
      d_arr_6_10=>DANGLING(1365), d_arr_6_9=>DANGLING(1366), d_arr_6_8=>
      DANGLING(1367), d_arr_6_7=>DANGLING(1368), d_arr_6_6=>DANGLING(1369), 
      d_arr_6_5=>DANGLING(1370), d_arr_6_4=>DANGLING(1371), d_arr_6_3=>
      DANGLING(1372), d_arr_6_2=>DANGLING(1373), d_arr_6_1=>DANGLING(1374), 
      d_arr_6_0=>DANGLING(1375), d_arr_7_31=>DANGLING(1376), d_arr_7_30=>
      DANGLING(1377), d_arr_7_29=>DANGLING(1378), d_arr_7_28=>DANGLING(1379), 
      d_arr_7_27=>DANGLING(1380), d_arr_7_26=>DANGLING(1381), d_arr_7_25=>
      DANGLING(1382), d_arr_7_24=>DANGLING(1383), d_arr_7_23=>DANGLING(1384), 
      d_arr_7_22=>DANGLING(1385), d_arr_7_21=>DANGLING(1386), d_arr_7_20=>
      DANGLING(1387), d_arr_7_19=>DANGLING(1388), d_arr_7_18=>DANGLING(1389), 
      d_arr_7_17=>DANGLING(1390), d_arr_7_16=>DANGLING(1391), d_arr_7_15=>
      DANGLING(1392), d_arr_7_14=>DANGLING(1393), d_arr_7_13=>DANGLING(1394), 
      d_arr_7_12=>DANGLING(1395), d_arr_7_11=>DANGLING(1396), d_arr_7_10=>
      DANGLING(1397), d_arr_7_9=>DANGLING(1398), d_arr_7_8=>DANGLING(1399), 
      d_arr_7_7=>DANGLING(1400), d_arr_7_6=>DANGLING(1401), d_arr_7_5=>
      DANGLING(1402), d_arr_7_4=>DANGLING(1403), d_arr_7_3=>DANGLING(1404), 
      d_arr_7_2=>DANGLING(1405), d_arr_7_1=>DANGLING(1406), d_arr_7_0=>
      DANGLING(1407), d_arr_8_31=>DANGLING(1408), d_arr_8_30=>DANGLING(1409), 
      d_arr_8_29=>DANGLING(1410), d_arr_8_28=>DANGLING(1411), d_arr_8_27=>
      DANGLING(1412), d_arr_8_26=>DANGLING(1413), d_arr_8_25=>DANGLING(1414), 
      d_arr_8_24=>DANGLING(1415), d_arr_8_23=>DANGLING(1416), d_arr_8_22=>
      DANGLING(1417), d_arr_8_21=>DANGLING(1418), d_arr_8_20=>DANGLING(1419), 
      d_arr_8_19=>DANGLING(1420), d_arr_8_18=>DANGLING(1421), d_arr_8_17=>
      DANGLING(1422), d_arr_8_16=>DANGLING(1423), d_arr_8_15=>DANGLING(1424), 
      d_arr_8_14=>DANGLING(1425), d_arr_8_13=>DANGLING(1426), d_arr_8_12=>
      DANGLING(1427), d_arr_8_11=>DANGLING(1428), d_arr_8_10=>DANGLING(1429), 
      d_arr_8_9=>DANGLING(1430), d_arr_8_8=>DANGLING(1431), d_arr_8_7=>
      DANGLING(1432), d_arr_8_6=>DANGLING(1433), d_arr_8_5=>DANGLING(1434), 
      d_arr_8_4=>DANGLING(1435), d_arr_8_3=>DANGLING(1436), d_arr_8_2=>
      DANGLING(1437), d_arr_8_1=>DANGLING(1438), d_arr_8_0=>DANGLING(1439), 
      d_arr_9_31=>DANGLING(1440), d_arr_9_30=>DANGLING(1441), d_arr_9_29=>
      DANGLING(1442), d_arr_9_28=>DANGLING(1443), d_arr_9_27=>DANGLING(1444), 
      d_arr_9_26=>DANGLING(1445), d_arr_9_25=>DANGLING(1446), d_arr_9_24=>
      DANGLING(1447), d_arr_9_23=>DANGLING(1448), d_arr_9_22=>DANGLING(1449), 
      d_arr_9_21=>DANGLING(1450), d_arr_9_20=>DANGLING(1451), d_arr_9_19=>
      DANGLING(1452), d_arr_9_18=>DANGLING(1453), d_arr_9_17=>DANGLING(1454), 
      d_arr_9_16=>DANGLING(1455), d_arr_9_15=>DANGLING(1456), d_arr_9_14=>
      DANGLING(1457), d_arr_9_13=>DANGLING(1458), d_arr_9_12=>DANGLING(1459), 
      d_arr_9_11=>DANGLING(1460), d_arr_9_10=>DANGLING(1461), d_arr_9_9=>
      DANGLING(1462), d_arr_9_8=>DANGLING(1463), d_arr_9_7=>DANGLING(1464), 
      d_arr_9_6=>DANGLING(1465), d_arr_9_5=>DANGLING(1466), d_arr_9_4=>
      DANGLING(1467), d_arr_9_3=>DANGLING(1468), d_arr_9_2=>DANGLING(1469), 
      d_arr_9_1=>DANGLING(1470), d_arr_9_0=>DANGLING(1471), d_arr_10_31=>
      DANGLING(1472), d_arr_10_30=>DANGLING(1473), d_arr_10_29=>DANGLING(
      1474), d_arr_10_28=>DANGLING(1475), d_arr_10_27=>DANGLING(1476), 
      d_arr_10_26=>DANGLING(1477), d_arr_10_25=>DANGLING(1478), d_arr_10_24
      =>DANGLING(1479), d_arr_10_23=>DANGLING(1480), d_arr_10_22=>DANGLING(
      1481), d_arr_10_21=>DANGLING(1482), d_arr_10_20=>DANGLING(1483), 
      d_arr_10_19=>DANGLING(1484), d_arr_10_18=>DANGLING(1485), d_arr_10_17
      =>DANGLING(1486), d_arr_10_16=>DANGLING(1487), d_arr_10_15=>DANGLING(
      1488), d_arr_10_14=>DANGLING(1489), d_arr_10_13=>DANGLING(1490), 
      d_arr_10_12=>DANGLING(1491), d_arr_10_11=>DANGLING(1492), d_arr_10_10
      =>DANGLING(1493), d_arr_10_9=>DANGLING(1494), d_arr_10_8=>DANGLING(
      1495), d_arr_10_7=>DANGLING(1496), d_arr_10_6=>DANGLING(1497), 
      d_arr_10_5=>DANGLING(1498), d_arr_10_4=>DANGLING(1499), d_arr_10_3=>
      DANGLING(1500), d_arr_10_2=>DANGLING(1501), d_arr_10_1=>DANGLING(1502), 
      d_arr_10_0=>DANGLING(1503), d_arr_11_31=>DANGLING(1504), d_arr_11_30=>
      DANGLING(1505), d_arr_11_29=>DANGLING(1506), d_arr_11_28=>DANGLING(
      1507), d_arr_11_27=>DANGLING(1508), d_arr_11_26=>DANGLING(1509), 
      d_arr_11_25=>DANGLING(1510), d_arr_11_24=>DANGLING(1511), d_arr_11_23
      =>DANGLING(1512), d_arr_11_22=>DANGLING(1513), d_arr_11_21=>DANGLING(
      1514), d_arr_11_20=>DANGLING(1515), d_arr_11_19=>DANGLING(1516), 
      d_arr_11_18=>DANGLING(1517), d_arr_11_17=>DANGLING(1518), d_arr_11_16
      =>DANGLING(1519), d_arr_11_15=>DANGLING(1520), d_arr_11_14=>DANGLING(
      1521), d_arr_11_13=>DANGLING(1522), d_arr_11_12=>DANGLING(1523), 
      d_arr_11_11=>DANGLING(1524), d_arr_11_10=>DANGLING(1525), d_arr_11_9=>
      DANGLING(1526), d_arr_11_8=>DANGLING(1527), d_arr_11_7=>DANGLING(1528), 
      d_arr_11_6=>DANGLING(1529), d_arr_11_5=>DANGLING(1530), d_arr_11_4=>
      DANGLING(1531), d_arr_11_3=>DANGLING(1532), d_arr_11_2=>DANGLING(1533), 
      d_arr_11_1=>DANGLING(1534), d_arr_11_0=>DANGLING(1535), d_arr_12_31=>
      DANGLING(1536), d_arr_12_30=>DANGLING(1537), d_arr_12_29=>DANGLING(
      1538), d_arr_12_28=>DANGLING(1539), d_arr_12_27=>DANGLING(1540), 
      d_arr_12_26=>DANGLING(1541), d_arr_12_25=>DANGLING(1542), d_arr_12_24
      =>DANGLING(1543), d_arr_12_23=>DANGLING(1544), d_arr_12_22=>DANGLING(
      1545), d_arr_12_21=>DANGLING(1546), d_arr_12_20=>DANGLING(1547), 
      d_arr_12_19=>DANGLING(1548), d_arr_12_18=>DANGLING(1549), d_arr_12_17
      =>DANGLING(1550), d_arr_12_16=>DANGLING(1551), d_arr_12_15=>DANGLING(
      1552), d_arr_12_14=>DANGLING(1553), d_arr_12_13=>DANGLING(1554), 
      d_arr_12_12=>DANGLING(1555), d_arr_12_11=>DANGLING(1556), d_arr_12_10
      =>DANGLING(1557), d_arr_12_9=>DANGLING(1558), d_arr_12_8=>DANGLING(
      1559), d_arr_12_7=>DANGLING(1560), d_arr_12_6=>DANGLING(1561), 
      d_arr_12_5=>DANGLING(1562), d_arr_12_4=>DANGLING(1563), d_arr_12_3=>
      DANGLING(1564), d_arr_12_2=>DANGLING(1565), d_arr_12_1=>DANGLING(1566), 
      d_arr_12_0=>DANGLING(1567), d_arr_13_31=>DANGLING(1568), d_arr_13_30=>
      DANGLING(1569), d_arr_13_29=>DANGLING(1570), d_arr_13_28=>DANGLING(
      1571), d_arr_13_27=>DANGLING(1572), d_arr_13_26=>DANGLING(1573), 
      d_arr_13_25=>DANGLING(1574), d_arr_13_24=>DANGLING(1575), d_arr_13_23
      =>DANGLING(1576), d_arr_13_22=>DANGLING(1577), d_arr_13_21=>DANGLING(
      1578), d_arr_13_20=>DANGLING(1579), d_arr_13_19=>DANGLING(1580), 
      d_arr_13_18=>DANGLING(1581), d_arr_13_17=>DANGLING(1582), d_arr_13_16
      =>DANGLING(1583), d_arr_13_15=>DANGLING(1584), d_arr_13_14=>DANGLING(
      1585), d_arr_13_13=>DANGLING(1586), d_arr_13_12=>DANGLING(1587), 
      d_arr_13_11=>DANGLING(1588), d_arr_13_10=>DANGLING(1589), d_arr_13_9=>
      DANGLING(1590), d_arr_13_8=>DANGLING(1591), d_arr_13_7=>DANGLING(1592), 
      d_arr_13_6=>DANGLING(1593), d_arr_13_5=>DANGLING(1594), d_arr_13_4=>
      DANGLING(1595), d_arr_13_3=>DANGLING(1596), d_arr_13_2=>DANGLING(1597), 
      d_arr_13_1=>DANGLING(1598), d_arr_13_0=>DANGLING(1599), d_arr_14_31=>
      DANGLING(1600), d_arr_14_30=>DANGLING(1601), d_arr_14_29=>DANGLING(
      1602), d_arr_14_28=>DANGLING(1603), d_arr_14_27=>DANGLING(1604), 
      d_arr_14_26=>DANGLING(1605), d_arr_14_25=>DANGLING(1606), d_arr_14_24
      =>DANGLING(1607), d_arr_14_23=>DANGLING(1608), d_arr_14_22=>DANGLING(
      1609), d_arr_14_21=>DANGLING(1610), d_arr_14_20=>DANGLING(1611), 
      d_arr_14_19=>DANGLING(1612), d_arr_14_18=>DANGLING(1613), d_arr_14_17
      =>DANGLING(1614), d_arr_14_16=>DANGLING(1615), d_arr_14_15=>DANGLING(
      1616), d_arr_14_14=>DANGLING(1617), d_arr_14_13=>DANGLING(1618), 
      d_arr_14_12=>DANGLING(1619), d_arr_14_11=>DANGLING(1620), d_arr_14_10
      =>DANGLING(1621), d_arr_14_9=>DANGLING(1622), d_arr_14_8=>DANGLING(
      1623), d_arr_14_7=>DANGLING(1624), d_arr_14_6=>DANGLING(1625), 
      d_arr_14_5=>DANGLING(1626), d_arr_14_4=>DANGLING(1627), d_arr_14_3=>
      DANGLING(1628), d_arr_14_2=>DANGLING(1629), d_arr_14_1=>DANGLING(1630), 
      d_arr_14_0=>DANGLING(1631), d_arr_15_31=>DANGLING(1632), d_arr_15_30=>
      DANGLING(1633), d_arr_15_29=>DANGLING(1634), d_arr_15_28=>DANGLING(
      1635), d_arr_15_27=>DANGLING(1636), d_arr_15_26=>DANGLING(1637), 
      d_arr_15_25=>DANGLING(1638), d_arr_15_24=>DANGLING(1639), d_arr_15_23
      =>DANGLING(1640), d_arr_15_22=>DANGLING(1641), d_arr_15_21=>DANGLING(
      1642), d_arr_15_20=>DANGLING(1643), d_arr_15_19=>DANGLING(1644), 
      d_arr_15_18=>DANGLING(1645), d_arr_15_17=>DANGLING(1646), d_arr_15_16
      =>DANGLING(1647), d_arr_15_15=>DANGLING(1648), d_arr_15_14=>DANGLING(
      1649), d_arr_15_13=>DANGLING(1650), d_arr_15_12=>DANGLING(1651), 
      d_arr_15_11=>DANGLING(1652), d_arr_15_10=>DANGLING(1653), d_arr_15_9=>
      DANGLING(1654), d_arr_15_8=>DANGLING(1655), d_arr_15_7=>DANGLING(1656), 
      d_arr_15_6=>DANGLING(1657), d_arr_15_5=>DANGLING(1658), d_arr_15_4=>
      DANGLING(1659), d_arr_15_3=>DANGLING(1660), d_arr_15_2=>DANGLING(1661), 
      d_arr_15_1=>DANGLING(1662), d_arr_15_0=>DANGLING(1663), d_arr_16_31=>
      DANGLING(1664), d_arr_16_30=>DANGLING(1665), d_arr_16_29=>DANGLING(
      1666), d_arr_16_28=>DANGLING(1667), d_arr_16_27=>DANGLING(1668), 
      d_arr_16_26=>DANGLING(1669), d_arr_16_25=>DANGLING(1670), d_arr_16_24
      =>DANGLING(1671), d_arr_16_23=>DANGLING(1672), d_arr_16_22=>DANGLING(
      1673), d_arr_16_21=>DANGLING(1674), d_arr_16_20=>DANGLING(1675), 
      d_arr_16_19=>DANGLING(1676), d_arr_16_18=>DANGLING(1677), d_arr_16_17
      =>DANGLING(1678), d_arr_16_16=>DANGLING(1679), d_arr_16_15=>DANGLING(
      1680), d_arr_16_14=>DANGLING(1681), d_arr_16_13=>DANGLING(1682), 
      d_arr_16_12=>DANGLING(1683), d_arr_16_11=>DANGLING(1684), d_arr_16_10
      =>DANGLING(1685), d_arr_16_9=>DANGLING(1686), d_arr_16_8=>DANGLING(
      1687), d_arr_16_7=>DANGLING(1688), d_arr_16_6=>DANGLING(1689), 
      d_arr_16_5=>DANGLING(1690), d_arr_16_4=>DANGLING(1691), d_arr_16_3=>
      DANGLING(1692), d_arr_16_2=>DANGLING(1693), d_arr_16_1=>DANGLING(1694), 
      d_arr_16_0=>DANGLING(1695), d_arr_17_31=>DANGLING(1696), d_arr_17_30=>
      DANGLING(1697), d_arr_17_29=>DANGLING(1698), d_arr_17_28=>DANGLING(
      1699), d_arr_17_27=>DANGLING(1700), d_arr_17_26=>DANGLING(1701), 
      d_arr_17_25=>DANGLING(1702), d_arr_17_24=>DANGLING(1703), d_arr_17_23
      =>DANGLING(1704), d_arr_17_22=>DANGLING(1705), d_arr_17_21=>DANGLING(
      1706), d_arr_17_20=>DANGLING(1707), d_arr_17_19=>DANGLING(1708), 
      d_arr_17_18=>DANGLING(1709), d_arr_17_17=>DANGLING(1710), d_arr_17_16
      =>DANGLING(1711), d_arr_17_15=>DANGLING(1712), d_arr_17_14=>DANGLING(
      1713), d_arr_17_13=>DANGLING(1714), d_arr_17_12=>DANGLING(1715), 
      d_arr_17_11=>DANGLING(1716), d_arr_17_10=>DANGLING(1717), d_arr_17_9=>
      DANGLING(1718), d_arr_17_8=>DANGLING(1719), d_arr_17_7=>DANGLING(1720), 
      d_arr_17_6=>DANGLING(1721), d_arr_17_5=>DANGLING(1722), d_arr_17_4=>
      DANGLING(1723), d_arr_17_3=>DANGLING(1724), d_arr_17_2=>DANGLING(1725), 
      d_arr_17_1=>DANGLING(1726), d_arr_17_0=>DANGLING(1727), d_arr_18_31=>
      DANGLING(1728), d_arr_18_30=>DANGLING(1729), d_arr_18_29=>DANGLING(
      1730), d_arr_18_28=>DANGLING(1731), d_arr_18_27=>DANGLING(1732), 
      d_arr_18_26=>DANGLING(1733), d_arr_18_25=>DANGLING(1734), d_arr_18_24
      =>DANGLING(1735), d_arr_18_23=>DANGLING(1736), d_arr_18_22=>DANGLING(
      1737), d_arr_18_21=>DANGLING(1738), d_arr_18_20=>DANGLING(1739), 
      d_arr_18_19=>DANGLING(1740), d_arr_18_18=>DANGLING(1741), d_arr_18_17
      =>DANGLING(1742), d_arr_18_16=>DANGLING(1743), d_arr_18_15=>DANGLING(
      1744), d_arr_18_14=>DANGLING(1745), d_arr_18_13=>DANGLING(1746), 
      d_arr_18_12=>DANGLING(1747), d_arr_18_11=>DANGLING(1748), d_arr_18_10
      =>DANGLING(1749), d_arr_18_9=>DANGLING(1750), d_arr_18_8=>DANGLING(
      1751), d_arr_18_7=>DANGLING(1752), d_arr_18_6=>DANGLING(1753), 
      d_arr_18_5=>DANGLING(1754), d_arr_18_4=>DANGLING(1755), d_arr_18_3=>
      DANGLING(1756), d_arr_18_2=>DANGLING(1757), d_arr_18_1=>DANGLING(1758), 
      d_arr_18_0=>DANGLING(1759), d_arr_19_31=>DANGLING(1760), d_arr_19_30=>
      DANGLING(1761), d_arr_19_29=>DANGLING(1762), d_arr_19_28=>DANGLING(
      1763), d_arr_19_27=>DANGLING(1764), d_arr_19_26=>DANGLING(1765), 
      d_arr_19_25=>DANGLING(1766), d_arr_19_24=>DANGLING(1767), d_arr_19_23
      =>DANGLING(1768), d_arr_19_22=>DANGLING(1769), d_arr_19_21=>DANGLING(
      1770), d_arr_19_20=>DANGLING(1771), d_arr_19_19=>DANGLING(1772), 
      d_arr_19_18=>DANGLING(1773), d_arr_19_17=>DANGLING(1774), d_arr_19_16
      =>DANGLING(1775), d_arr_19_15=>DANGLING(1776), d_arr_19_14=>DANGLING(
      1777), d_arr_19_13=>DANGLING(1778), d_arr_19_12=>DANGLING(1779), 
      d_arr_19_11=>DANGLING(1780), d_arr_19_10=>DANGLING(1781), d_arr_19_9=>
      DANGLING(1782), d_arr_19_8=>DANGLING(1783), d_arr_19_7=>DANGLING(1784), 
      d_arr_19_6=>DANGLING(1785), d_arr_19_5=>DANGLING(1786), d_arr_19_4=>
      DANGLING(1787), d_arr_19_3=>DANGLING(1788), d_arr_19_2=>DANGLING(1789), 
      d_arr_19_1=>DANGLING(1790), d_arr_19_0=>DANGLING(1791), d_arr_20_31=>
      DANGLING(1792), d_arr_20_30=>DANGLING(1793), d_arr_20_29=>DANGLING(
      1794), d_arr_20_28=>DANGLING(1795), d_arr_20_27=>DANGLING(1796), 
      d_arr_20_26=>DANGLING(1797), d_arr_20_25=>DANGLING(1798), d_arr_20_24
      =>DANGLING(1799), d_arr_20_23=>DANGLING(1800), d_arr_20_22=>DANGLING(
      1801), d_arr_20_21=>DANGLING(1802), d_arr_20_20=>DANGLING(1803), 
      d_arr_20_19=>DANGLING(1804), d_arr_20_18=>DANGLING(1805), d_arr_20_17
      =>DANGLING(1806), d_arr_20_16=>DANGLING(1807), d_arr_20_15=>DANGLING(
      1808), d_arr_20_14=>DANGLING(1809), d_arr_20_13=>DANGLING(1810), 
      d_arr_20_12=>DANGLING(1811), d_arr_20_11=>DANGLING(1812), d_arr_20_10
      =>DANGLING(1813), d_arr_20_9=>DANGLING(1814), d_arr_20_8=>DANGLING(
      1815), d_arr_20_7=>DANGLING(1816), d_arr_20_6=>DANGLING(1817), 
      d_arr_20_5=>DANGLING(1818), d_arr_20_4=>DANGLING(1819), d_arr_20_3=>
      DANGLING(1820), d_arr_20_2=>DANGLING(1821), d_arr_20_1=>DANGLING(1822), 
      d_arr_20_0=>DANGLING(1823), d_arr_21_31=>DANGLING(1824), d_arr_21_30=>
      DANGLING(1825), d_arr_21_29=>DANGLING(1826), d_arr_21_28=>DANGLING(
      1827), d_arr_21_27=>DANGLING(1828), d_arr_21_26=>DANGLING(1829), 
      d_arr_21_25=>DANGLING(1830), d_arr_21_24=>DANGLING(1831), d_arr_21_23
      =>DANGLING(1832), d_arr_21_22=>DANGLING(1833), d_arr_21_21=>DANGLING(
      1834), d_arr_21_20=>DANGLING(1835), d_arr_21_19=>DANGLING(1836), 
      d_arr_21_18=>DANGLING(1837), d_arr_21_17=>DANGLING(1838), d_arr_21_16
      =>DANGLING(1839), d_arr_21_15=>DANGLING(1840), d_arr_21_14=>DANGLING(
      1841), d_arr_21_13=>DANGLING(1842), d_arr_21_12=>DANGLING(1843), 
      d_arr_21_11=>DANGLING(1844), d_arr_21_10=>DANGLING(1845), d_arr_21_9=>
      DANGLING(1846), d_arr_21_8=>DANGLING(1847), d_arr_21_7=>DANGLING(1848), 
      d_arr_21_6=>DANGLING(1849), d_arr_21_5=>DANGLING(1850), d_arr_21_4=>
      DANGLING(1851), d_arr_21_3=>DANGLING(1852), d_arr_21_2=>DANGLING(1853), 
      d_arr_21_1=>DANGLING(1854), d_arr_21_0=>DANGLING(1855), d_arr_22_31=>
      DANGLING(1856), d_arr_22_30=>DANGLING(1857), d_arr_22_29=>DANGLING(
      1858), d_arr_22_28=>DANGLING(1859), d_arr_22_27=>DANGLING(1860), 
      d_arr_22_26=>DANGLING(1861), d_arr_22_25=>DANGLING(1862), d_arr_22_24
      =>DANGLING(1863), d_arr_22_23=>DANGLING(1864), d_arr_22_22=>DANGLING(
      1865), d_arr_22_21=>DANGLING(1866), d_arr_22_20=>DANGLING(1867), 
      d_arr_22_19=>DANGLING(1868), d_arr_22_18=>DANGLING(1869), d_arr_22_17
      =>DANGLING(1870), d_arr_22_16=>DANGLING(1871), d_arr_22_15=>DANGLING(
      1872), d_arr_22_14=>DANGLING(1873), d_arr_22_13=>DANGLING(1874), 
      d_arr_22_12=>DANGLING(1875), d_arr_22_11=>DANGLING(1876), d_arr_22_10
      =>DANGLING(1877), d_arr_22_9=>DANGLING(1878), d_arr_22_8=>DANGLING(
      1879), d_arr_22_7=>DANGLING(1880), d_arr_22_6=>DANGLING(1881), 
      d_arr_22_5=>DANGLING(1882), d_arr_22_4=>DANGLING(1883), d_arr_22_3=>
      DANGLING(1884), d_arr_22_2=>DANGLING(1885), d_arr_22_1=>DANGLING(1886), 
      d_arr_22_0=>DANGLING(1887), d_arr_23_31=>DANGLING(1888), d_arr_23_30=>
      DANGLING(1889), d_arr_23_29=>DANGLING(1890), d_arr_23_28=>DANGLING(
      1891), d_arr_23_27=>DANGLING(1892), d_arr_23_26=>DANGLING(1893), 
      d_arr_23_25=>DANGLING(1894), d_arr_23_24=>DANGLING(1895), d_arr_23_23
      =>DANGLING(1896), d_arr_23_22=>DANGLING(1897), d_arr_23_21=>DANGLING(
      1898), d_arr_23_20=>DANGLING(1899), d_arr_23_19=>DANGLING(1900), 
      d_arr_23_18=>DANGLING(1901), d_arr_23_17=>DANGLING(1902), d_arr_23_16
      =>DANGLING(1903), d_arr_23_15=>DANGLING(1904), d_arr_23_14=>DANGLING(
      1905), d_arr_23_13=>DANGLING(1906), d_arr_23_12=>DANGLING(1907), 
      d_arr_23_11=>DANGLING(1908), d_arr_23_10=>DANGLING(1909), d_arr_23_9=>
      DANGLING(1910), d_arr_23_8=>DANGLING(1911), d_arr_23_7=>DANGLING(1912), 
      d_arr_23_6=>DANGLING(1913), d_arr_23_5=>DANGLING(1914), d_arr_23_4=>
      DANGLING(1915), d_arr_23_3=>DANGLING(1916), d_arr_23_2=>DANGLING(1917), 
      d_arr_23_1=>DANGLING(1918), d_arr_23_0=>DANGLING(1919), d_arr_24_31=>
      DANGLING(1920), d_arr_24_30=>DANGLING(1921), d_arr_24_29=>DANGLING(
      1922), d_arr_24_28=>DANGLING(1923), d_arr_24_27=>DANGLING(1924), 
      d_arr_24_26=>DANGLING(1925), d_arr_24_25=>DANGLING(1926), d_arr_24_24
      =>DANGLING(1927), d_arr_24_23=>DANGLING(1928), d_arr_24_22=>DANGLING(
      1929), d_arr_24_21=>DANGLING(1930), d_arr_24_20=>DANGLING(1931), 
      d_arr_24_19=>DANGLING(1932), d_arr_24_18=>DANGLING(1933), d_arr_24_17
      =>DANGLING(1934), d_arr_24_16=>DANGLING(1935), d_arr_24_15=>DANGLING(
      1936), d_arr_24_14=>DANGLING(1937), d_arr_24_13=>DANGLING(1938), 
      d_arr_24_12=>DANGLING(1939), d_arr_24_11=>DANGLING(1940), d_arr_24_10
      =>DANGLING(1941), d_arr_24_9=>DANGLING(1942), d_arr_24_8=>DANGLING(
      1943), d_arr_24_7=>DANGLING(1944), d_arr_24_6=>DANGLING(1945), 
      d_arr_24_5=>DANGLING(1946), d_arr_24_4=>DANGLING(1947), d_arr_24_3=>
      DANGLING(1948), d_arr_24_2=>DANGLING(1949), d_arr_24_1=>DANGLING(1950), 
      d_arr_24_0=>DANGLING(1951), q_arr_0_31=>nx19448, q_arr_0_30=>nx16499, 
      q_arr_0_29=>nx16503, q_arr_0_28=>nx16507, q_arr_0_27=>nx19388, 
      q_arr_0_26=>nx16515, q_arr_0_25=>nx16519, q_arr_0_24=>nx19390, 
      q_arr_0_23=>nx16527, q_arr_0_22=>nx16531, q_arr_0_21=>nx16535, 
      q_arr_0_20=>nx16539, q_arr_0_19=>nx16543, q_arr_0_18=>nx16547, 
      q_arr_0_17=>nx16551, q_arr_0_16=>nx16555, q_arr_0_15=>nx16559, 
      q_arr_0_14=>nx16563, q_arr_0_13=>nx16567, q_arr_0_12=>nx16571, 
      q_arr_0_11=>nx16575, q_arr_0_10=>nx16579, q_arr_0_9=>nx16583, 
      q_arr_0_8=>nx16587, q_arr_0_7=>nx16591, q_arr_0_6=>nx16595, q_arr_0_5
      =>nx16599, q_arr_0_4=>nx16601, q_arr_0_3=>nx16603, q_arr_0_2=>
      q_arr_0_2, q_arr_0_1=>q_arr_0_1, q_arr_0_0=>nx16605, q_arr_1_31=>GND0, 
      q_arr_1_30=>GND0, q_arr_1_29=>GND0, q_arr_1_28=>GND0, q_arr_1_27=>GND0, 
      q_arr_1_26=>GND0, q_arr_1_25=>GND0, q_arr_1_24=>GND0, q_arr_1_23=>GND0, 
      q_arr_1_22=>GND0, q_arr_1_21=>GND0, q_arr_1_20=>GND0, q_arr_1_19=>GND0, 
      q_arr_1_18=>GND0, q_arr_1_17=>GND0, q_arr_1_16=>GND0, q_arr_1_15=>GND0, 
      q_arr_1_14=>GND0, q_arr_1_13=>GND0, q_arr_1_12=>GND0, q_arr_1_11=>GND0, 
      q_arr_1_10=>GND0, q_arr_1_9=>GND0, q_arr_1_8=>GND0, q_arr_1_7=>GND0, 
      q_arr_1_6=>GND0, q_arr_1_5=>GND0, q_arr_1_4=>GND0, q_arr_1_3=>GND0, 
      q_arr_1_2=>GND0, q_arr_1_1=>GND0, q_arr_1_0=>GND0, q_arr_2_31=>GND0, 
      q_arr_2_30=>GND0, q_arr_2_29=>GND0, q_arr_2_28=>GND0, q_arr_2_27=>GND0, 
      q_arr_2_26=>GND0, q_arr_2_25=>GND0, q_arr_2_24=>GND0, q_arr_2_23=>GND0, 
      q_arr_2_22=>GND0, q_arr_2_21=>GND0, q_arr_2_20=>GND0, q_arr_2_19=>GND0, 
      q_arr_2_18=>GND0, q_arr_2_17=>GND0, q_arr_2_16=>GND0, q_arr_2_15=>GND0, 
      q_arr_2_14=>GND0, q_arr_2_13=>GND0, q_arr_2_12=>GND0, q_arr_2_11=>GND0, 
      q_arr_2_10=>GND0, q_arr_2_9=>GND0, q_arr_2_8=>GND0, q_arr_2_7=>GND0, 
      q_arr_2_6=>GND0, q_arr_2_5=>GND0, q_arr_2_4=>GND0, q_arr_2_3=>GND0, 
      q_arr_2_2=>GND0, q_arr_2_1=>GND0, q_arr_2_0=>GND0, q_arr_3_31=>GND0, 
      q_arr_3_30=>GND0, q_arr_3_29=>GND0, q_arr_3_28=>GND0, q_arr_3_27=>GND0, 
      q_arr_3_26=>GND0, q_arr_3_25=>GND0, q_arr_3_24=>GND0, q_arr_3_23=>GND0, 
      q_arr_3_22=>GND0, q_arr_3_21=>GND0, q_arr_3_20=>GND0, q_arr_3_19=>GND0, 
      q_arr_3_18=>GND0, q_arr_3_17=>GND0, q_arr_3_16=>GND0, q_arr_3_15=>GND0, 
      q_arr_3_14=>GND0, q_arr_3_13=>GND0, q_arr_3_12=>GND0, q_arr_3_11=>GND0, 
      q_arr_3_10=>GND0, q_arr_3_9=>GND0, q_arr_3_8=>GND0, q_arr_3_7=>GND0, 
      q_arr_3_6=>GND0, q_arr_3_5=>GND0, q_arr_3_4=>GND0, q_arr_3_3=>GND0, 
      q_arr_3_2=>GND0, q_arr_3_1=>GND0, q_arr_3_0=>GND0, q_arr_4_31=>GND0, 
      q_arr_4_30=>GND0, q_arr_4_29=>GND0, q_arr_4_28=>GND0, q_arr_4_27=>GND0, 
      q_arr_4_26=>GND0, q_arr_4_25=>GND0, q_arr_4_24=>GND0, q_arr_4_23=>GND0, 
      q_arr_4_22=>GND0, q_arr_4_21=>GND0, q_arr_4_20=>GND0, q_arr_4_19=>GND0, 
      q_arr_4_18=>GND0, q_arr_4_17=>GND0, q_arr_4_16=>GND0, q_arr_4_15=>GND0, 
      q_arr_4_14=>GND0, q_arr_4_13=>GND0, q_arr_4_12=>GND0, q_arr_4_11=>GND0, 
      q_arr_4_10=>GND0, q_arr_4_9=>GND0, q_arr_4_8=>GND0, q_arr_4_7=>GND0, 
      q_arr_4_6=>GND0, q_arr_4_5=>GND0, q_arr_4_4=>GND0, q_arr_4_3=>GND0, 
      q_arr_4_2=>GND0, q_arr_4_1=>GND0, q_arr_4_0=>GND0, q_arr_5_31=>GND0, 
      q_arr_5_30=>GND0, q_arr_5_29=>GND0, q_arr_5_28=>GND0, q_arr_5_27=>GND0, 
      q_arr_5_26=>GND0, q_arr_5_25=>GND0, q_arr_5_24=>GND0, q_arr_5_23=>GND0, 
      q_arr_5_22=>GND0, q_arr_5_21=>GND0, q_arr_5_20=>GND0, q_arr_5_19=>GND0, 
      q_arr_5_18=>GND0, q_arr_5_17=>GND0, q_arr_5_16=>GND0, q_arr_5_15=>GND0, 
      q_arr_5_14=>GND0, q_arr_5_13=>GND0, q_arr_5_12=>GND0, q_arr_5_11=>GND0, 
      q_arr_5_10=>GND0, q_arr_5_9=>GND0, q_arr_5_8=>GND0, q_arr_5_7=>GND0, 
      q_arr_5_6=>GND0, q_arr_5_5=>GND0, q_arr_5_4=>GND0, q_arr_5_3=>GND0, 
      q_arr_5_2=>GND0, q_arr_5_1=>GND0, q_arr_5_0=>GND0, q_arr_6_31=>GND0, 
      q_arr_6_30=>GND0, q_arr_6_29=>GND0, q_arr_6_28=>GND0, q_arr_6_27=>GND0, 
      q_arr_6_26=>GND0, q_arr_6_25=>GND0, q_arr_6_24=>GND0, q_arr_6_23=>GND0, 
      q_arr_6_22=>GND0, q_arr_6_21=>GND0, q_arr_6_20=>GND0, q_arr_6_19=>GND0, 
      q_arr_6_18=>GND0, q_arr_6_17=>GND0, q_arr_6_16=>GND0, q_arr_6_15=>GND0, 
      q_arr_6_14=>GND0, q_arr_6_13=>GND0, q_arr_6_12=>GND0, q_arr_6_11=>GND0, 
      q_arr_6_10=>GND0, q_arr_6_9=>GND0, q_arr_6_8=>GND0, q_arr_6_7=>GND0, 
      q_arr_6_6=>GND0, q_arr_6_5=>GND0, q_arr_6_4=>GND0, q_arr_6_3=>GND0, 
      q_arr_6_2=>GND0, q_arr_6_1=>GND0, q_arr_6_0=>GND0, q_arr_7_31=>GND0, 
      q_arr_7_30=>GND0, q_arr_7_29=>GND0, q_arr_7_28=>GND0, q_arr_7_27=>GND0, 
      q_arr_7_26=>GND0, q_arr_7_25=>GND0, q_arr_7_24=>GND0, q_arr_7_23=>GND0, 
      q_arr_7_22=>GND0, q_arr_7_21=>GND0, q_arr_7_20=>GND0, q_arr_7_19=>GND0, 
      q_arr_7_18=>GND0, q_arr_7_17=>GND0, q_arr_7_16=>GND0, q_arr_7_15=>GND0, 
      q_arr_7_14=>GND0, q_arr_7_13=>GND0, q_arr_7_12=>GND0, q_arr_7_11=>GND0, 
      q_arr_7_10=>GND0, q_arr_7_9=>GND0, q_arr_7_8=>GND0, q_arr_7_7=>GND0, 
      q_arr_7_6=>GND0, q_arr_7_5=>GND0, q_arr_7_4=>GND0, q_arr_7_3=>GND0, 
      q_arr_7_2=>GND0, q_arr_7_1=>GND0, q_arr_7_0=>GND0, q_arr_8_31=>GND0, 
      q_arr_8_30=>GND0, q_arr_8_29=>GND0, q_arr_8_28=>GND0, q_arr_8_27=>GND0, 
      q_arr_8_26=>GND0, q_arr_8_25=>GND0, q_arr_8_24=>GND0, q_arr_8_23=>GND0, 
      q_arr_8_22=>GND0, q_arr_8_21=>GND0, q_arr_8_20=>GND0, q_arr_8_19=>GND0, 
      q_arr_8_18=>GND0, q_arr_8_17=>GND0, q_arr_8_16=>GND0, q_arr_8_15=>GND0, 
      q_arr_8_14=>GND0, q_arr_8_13=>GND0, q_arr_8_12=>GND0, q_arr_8_11=>GND0, 
      q_arr_8_10=>GND0, q_arr_8_9=>GND0, q_arr_8_8=>GND0, q_arr_8_7=>GND0, 
      q_arr_8_6=>GND0, q_arr_8_5=>GND0, q_arr_8_4=>GND0, q_arr_8_3=>GND0, 
      q_arr_8_2=>GND0, q_arr_8_1=>GND0, q_arr_8_0=>GND0, q_arr_9_31=>
      q_arr_9_31, q_arr_9_30=>q_arr_9_30, q_arr_9_29=>q_arr_9_29, q_arr_9_28
      =>q_arr_9_28, q_arr_9_27=>q_arr_9_27, q_arr_9_26=>q_arr_9_26, 
      q_arr_9_25=>q_arr_9_25, q_arr_9_24=>q_arr_9_24, q_arr_9_23=>q_arr_9_23, 
      q_arr_9_22=>q_arr_9_22, q_arr_9_21=>q_arr_9_21, q_arr_9_20=>q_arr_9_20, 
      q_arr_9_19=>q_arr_9_19, q_arr_9_18=>q_arr_9_18, q_arr_9_17=>q_arr_9_17, 
      q_arr_9_16=>q_arr_9_16, q_arr_9_15=>q_arr_9_15, q_arr_9_14=>q_arr_9_14, 
      q_arr_9_13=>q_arr_9_13, q_arr_9_12=>q_arr_9_12, q_arr_9_11=>q_arr_9_11, 
      q_arr_9_10=>q_arr_9_10, q_arr_9_9=>q_arr_9_9, q_arr_9_8=>q_arr_9_8, 
      q_arr_9_7=>q_arr_9_7, q_arr_9_6=>q_arr_9_6, q_arr_9_5=>q_arr_9_5, 
      q_arr_9_4=>q_arr_9_4, q_arr_9_3=>q_arr_9_3, q_arr_9_2=>q_arr_9_2, 
      q_arr_9_1=>q_arr_9_1, q_arr_9_0=>q_arr_9_0, q_arr_10_31=>GND0, 
      q_arr_10_30=>GND0, q_arr_10_29=>GND0, q_arr_10_28=>GND0, q_arr_10_27=>
      GND0, q_arr_10_26=>GND0, q_arr_10_25=>GND0, q_arr_10_24=>GND0, 
      q_arr_10_23=>GND0, q_arr_10_22=>GND0, q_arr_10_21=>GND0, q_arr_10_20=>
      GND0, q_arr_10_19=>GND0, q_arr_10_18=>GND0, q_arr_10_17=>GND0, 
      q_arr_10_16=>GND0, q_arr_10_15=>GND0, q_arr_10_14=>GND0, q_arr_10_13=>
      GND0, q_arr_10_12=>GND0, q_arr_10_11=>GND0, q_arr_10_10=>GND0, 
      q_arr_10_9=>GND0, q_arr_10_8=>GND0, q_arr_10_7=>GND0, q_arr_10_6=>GND0, 
      q_arr_10_5=>GND0, q_arr_10_4=>GND0, q_arr_10_3=>GND0, q_arr_10_2=>GND0, 
      q_arr_10_1=>GND0, q_arr_10_0=>GND0, q_arr_11_31=>GND0, q_arr_11_30=>
      GND0, q_arr_11_29=>GND0, q_arr_11_28=>GND0, q_arr_11_27=>GND0, 
      q_arr_11_26=>GND0, q_arr_11_25=>GND0, q_arr_11_24=>GND0, q_arr_11_23=>
      GND0, q_arr_11_22=>GND0, q_arr_11_21=>GND0, q_arr_11_20=>GND0, 
      q_arr_11_19=>GND0, q_arr_11_18=>GND0, q_arr_11_17=>GND0, q_arr_11_16=>
      GND0, q_arr_11_15=>GND0, q_arr_11_14=>GND0, q_arr_11_13=>GND0, 
      q_arr_11_12=>GND0, q_arr_11_11=>GND0, q_arr_11_10=>GND0, q_arr_11_9=>
      GND0, q_arr_11_8=>GND0, q_arr_11_7=>GND0, q_arr_11_6=>GND0, q_arr_11_5
      =>GND0, q_arr_11_4=>GND0, q_arr_11_3=>GND0, q_arr_11_2=>GND0, 
      q_arr_11_1=>GND0, q_arr_11_0=>GND0, q_arr_12_31=>GND0, q_arr_12_30=>
      GND0, q_arr_12_29=>GND0, q_arr_12_28=>GND0, q_arr_12_27=>GND0, 
      q_arr_12_26=>GND0, q_arr_12_25=>GND0, q_arr_12_24=>GND0, q_arr_12_23=>
      GND0, q_arr_12_22=>GND0, q_arr_12_21=>GND0, q_arr_12_20=>GND0, 
      q_arr_12_19=>GND0, q_arr_12_18=>GND0, q_arr_12_17=>GND0, q_arr_12_16=>
      GND0, q_arr_12_15=>GND0, q_arr_12_14=>GND0, q_arr_12_13=>GND0, 
      q_arr_12_12=>GND0, q_arr_12_11=>GND0, q_arr_12_10=>GND0, q_arr_12_9=>
      GND0, q_arr_12_8=>GND0, q_arr_12_7=>GND0, q_arr_12_6=>GND0, q_arr_12_5
      =>GND0, q_arr_12_4=>GND0, q_arr_12_3=>GND0, q_arr_12_2=>GND0, 
      q_arr_12_1=>GND0, q_arr_12_0=>GND0, q_arr_13_31=>GND0, q_arr_13_30=>
      GND0, q_arr_13_29=>GND0, q_arr_13_28=>GND0, q_arr_13_27=>GND0, 
      q_arr_13_26=>GND0, q_arr_13_25=>GND0, q_arr_13_24=>GND0, q_arr_13_23=>
      GND0, q_arr_13_22=>GND0, q_arr_13_21=>GND0, q_arr_13_20=>GND0, 
      q_arr_13_19=>GND0, q_arr_13_18=>GND0, q_arr_13_17=>GND0, q_arr_13_16=>
      GND0, q_arr_13_15=>GND0, q_arr_13_14=>GND0, q_arr_13_13=>GND0, 
      q_arr_13_12=>GND0, q_arr_13_11=>GND0, q_arr_13_10=>GND0, q_arr_13_9=>
      GND0, q_arr_13_8=>GND0, q_arr_13_7=>GND0, q_arr_13_6=>GND0, q_arr_13_5
      =>GND0, q_arr_13_4=>GND0, q_arr_13_3=>GND0, q_arr_13_2=>GND0, 
      q_arr_13_1=>GND0, q_arr_13_0=>GND0, q_arr_14_31=>GND0, q_arr_14_30=>
      GND0, q_arr_14_29=>GND0, q_arr_14_28=>GND0, q_arr_14_27=>GND0, 
      q_arr_14_26=>GND0, q_arr_14_25=>GND0, q_arr_14_24=>GND0, q_arr_14_23=>
      GND0, q_arr_14_22=>GND0, q_arr_14_21=>GND0, q_arr_14_20=>GND0, 
      q_arr_14_19=>GND0, q_arr_14_18=>GND0, q_arr_14_17=>GND0, q_arr_14_16=>
      GND0, q_arr_14_15=>GND0, q_arr_14_14=>GND0, q_arr_14_13=>GND0, 
      q_arr_14_12=>GND0, q_arr_14_11=>GND0, q_arr_14_10=>GND0, q_arr_14_9=>
      GND0, q_arr_14_8=>GND0, q_arr_14_7=>GND0, q_arr_14_6=>GND0, q_arr_14_5
      =>GND0, q_arr_14_4=>GND0, q_arr_14_3=>GND0, q_arr_14_2=>GND0, 
      q_arr_14_1=>GND0, q_arr_14_0=>GND0, q_arr_15_31=>GND0, q_arr_15_30=>
      GND0, q_arr_15_29=>GND0, q_arr_15_28=>GND0, q_arr_15_27=>GND0, 
      q_arr_15_26=>GND0, q_arr_15_25=>GND0, q_arr_15_24=>GND0, q_arr_15_23=>
      GND0, q_arr_15_22=>GND0, q_arr_15_21=>GND0, q_arr_15_20=>GND0, 
      q_arr_15_19=>GND0, q_arr_15_18=>GND0, q_arr_15_17=>GND0, q_arr_15_16=>
      GND0, q_arr_15_15=>GND0, q_arr_15_14=>GND0, q_arr_15_13=>GND0, 
      q_arr_15_12=>GND0, q_arr_15_11=>GND0, q_arr_15_10=>GND0, q_arr_15_9=>
      GND0, q_arr_15_8=>GND0, q_arr_15_7=>GND0, q_arr_15_6=>GND0, q_arr_15_5
      =>GND0, q_arr_15_4=>GND0, q_arr_15_3=>GND0, q_arr_15_2=>GND0, 
      q_arr_15_1=>GND0, q_arr_15_0=>GND0, q_arr_16_31=>GND0, q_arr_16_30=>
      GND0, q_arr_16_29=>GND0, q_arr_16_28=>GND0, q_arr_16_27=>GND0, 
      q_arr_16_26=>GND0, q_arr_16_25=>GND0, q_arr_16_24=>GND0, q_arr_16_23=>
      GND0, q_arr_16_22=>GND0, q_arr_16_21=>GND0, q_arr_16_20=>GND0, 
      q_arr_16_19=>GND0, q_arr_16_18=>GND0, q_arr_16_17=>GND0, q_arr_16_16=>
      GND0, q_arr_16_15=>GND0, q_arr_16_14=>GND0, q_arr_16_13=>GND0, 
      q_arr_16_12=>GND0, q_arr_16_11=>GND0, q_arr_16_10=>GND0, q_arr_16_9=>
      GND0, q_arr_16_8=>GND0, q_arr_16_7=>GND0, q_arr_16_6=>GND0, q_arr_16_5
      =>GND0, q_arr_16_4=>GND0, q_arr_16_3=>GND0, q_arr_16_2=>GND0, 
      q_arr_16_1=>GND0, q_arr_16_0=>GND0, q_arr_17_31=>GND0, q_arr_17_30=>
      GND0, q_arr_17_29=>GND0, q_arr_17_28=>GND0, q_arr_17_27=>GND0, 
      q_arr_17_26=>GND0, q_arr_17_25=>GND0, q_arr_17_24=>GND0, q_arr_17_23=>
      GND0, q_arr_17_22=>GND0, q_arr_17_21=>GND0, q_arr_17_20=>GND0, 
      q_arr_17_19=>GND0, q_arr_17_18=>GND0, q_arr_17_17=>GND0, q_arr_17_16=>
      GND0, q_arr_17_15=>GND0, q_arr_17_14=>GND0, q_arr_17_13=>GND0, 
      q_arr_17_12=>GND0, q_arr_17_11=>GND0, q_arr_17_10=>GND0, q_arr_17_9=>
      GND0, q_arr_17_8=>GND0, q_arr_17_7=>GND0, q_arr_17_6=>GND0, q_arr_17_5
      =>GND0, q_arr_17_4=>GND0, q_arr_17_3=>GND0, q_arr_17_2=>GND0, 
      q_arr_17_1=>GND0, q_arr_17_0=>GND0, q_arr_18_31=>q_arr_18_31, 
      q_arr_18_30=>q_arr_18_30, q_arr_18_29=>q_arr_18_29, q_arr_18_28=>
      q_arr_18_28, q_arr_18_27=>nx19488, q_arr_18_26=>q_arr_18_26, 
      q_arr_18_25=>q_arr_18_25, q_arr_18_24=>nx19492, q_arr_18_23=>
      q_arr_18_23, q_arr_18_22=>q_arr_18_22, q_arr_18_21=>q_arr_18_21, 
      q_arr_18_20=>q_arr_18_20, q_arr_18_19=>q_arr_18_19, q_arr_18_18=>
      q_arr_18_18, q_arr_18_17=>q_arr_18_17, q_arr_18_16=>q_arr_18_16, 
      q_arr_18_15=>q_arr_18_15, q_arr_18_14=>q_arr_18_14, q_arr_18_13=>
      q_arr_18_13, q_arr_18_12=>q_arr_18_12, q_arr_18_11=>q_arr_18_11, 
      q_arr_18_10=>q_arr_18_10, q_arr_18_9=>q_arr_18_9, q_arr_18_8=>
      q_arr_18_8, q_arr_18_7=>q_arr_18_7, q_arr_18_6=>q_arr_18_6, q_arr_18_5
      =>q_arr_18_5, q_arr_18_4=>q_arr_18_4, q_arr_18_3=>q_arr_18_3, 
      q_arr_18_2=>q_arr_18_2, q_arr_18_1=>q_arr_18_1, q_arr_18_0=>q_arr_18_0, 
      q_arr_19_31=>GND0, q_arr_19_30=>GND0, q_arr_19_29=>GND0, q_arr_19_28=>
      GND0, q_arr_19_27=>GND0, q_arr_19_26=>GND0, q_arr_19_25=>GND0, 
      q_arr_19_24=>GND0, q_arr_19_23=>GND0, q_arr_19_22=>GND0, q_arr_19_21=>
      GND0, q_arr_19_20=>GND0, q_arr_19_19=>GND0, q_arr_19_18=>GND0, 
      q_arr_19_17=>GND0, q_arr_19_16=>GND0, q_arr_19_15=>GND0, q_arr_19_14=>
      GND0, q_arr_19_13=>GND0, q_arr_19_12=>GND0, q_arr_19_11=>GND0, 
      q_arr_19_10=>GND0, q_arr_19_9=>GND0, q_arr_19_8=>GND0, q_arr_19_7=>
      GND0, q_arr_19_6=>GND0, q_arr_19_5=>GND0, q_arr_19_4=>GND0, q_arr_19_3
      =>GND0, q_arr_19_2=>GND0, q_arr_19_1=>GND0, q_arr_19_0=>GND0, 
      q_arr_20_31=>GND0, q_arr_20_30=>GND0, q_arr_20_29=>GND0, q_arr_20_28=>
      GND0, q_arr_20_27=>GND0, q_arr_20_26=>GND0, q_arr_20_25=>GND0, 
      q_arr_20_24=>GND0, q_arr_20_23=>GND0, q_arr_20_22=>GND0, q_arr_20_21=>
      GND0, q_arr_20_20=>GND0, q_arr_20_19=>GND0, q_arr_20_18=>GND0, 
      q_arr_20_17=>GND0, q_arr_20_16=>GND0, q_arr_20_15=>GND0, q_arr_20_14=>
      GND0, q_arr_20_13=>GND0, q_arr_20_12=>GND0, q_arr_20_11=>GND0, 
      q_arr_20_10=>GND0, q_arr_20_9=>GND0, q_arr_20_8=>GND0, q_arr_20_7=>
      GND0, q_arr_20_6=>GND0, q_arr_20_5=>GND0, q_arr_20_4=>GND0, q_arr_20_3
      =>GND0, q_arr_20_2=>GND0, q_arr_20_1=>GND0, q_arr_20_0=>GND0, 
      q_arr_21_31=>GND0, q_arr_21_30=>GND0, q_arr_21_29=>GND0, q_arr_21_28=>
      GND0, q_arr_21_27=>GND0, q_arr_21_26=>GND0, q_arr_21_25=>GND0, 
      q_arr_21_24=>GND0, q_arr_21_23=>GND0, q_arr_21_22=>GND0, q_arr_21_21=>
      GND0, q_arr_21_20=>GND0, q_arr_21_19=>GND0, q_arr_21_18=>GND0, 
      q_arr_21_17=>GND0, q_arr_21_16=>GND0, q_arr_21_15=>GND0, q_arr_21_14=>
      GND0, q_arr_21_13=>GND0, q_arr_21_12=>GND0, q_arr_21_11=>GND0, 
      q_arr_21_10=>GND0, q_arr_21_9=>GND0, q_arr_21_8=>GND0, q_arr_21_7=>
      GND0, q_arr_21_6=>GND0, q_arr_21_5=>GND0, q_arr_21_4=>GND0, q_arr_21_3
      =>GND0, q_arr_21_2=>GND0, q_arr_21_1=>GND0, q_arr_21_0=>GND0, 
      q_arr_22_31=>GND0, q_arr_22_30=>GND0, q_arr_22_29=>GND0, q_arr_22_28=>
      GND0, q_arr_22_27=>GND0, q_arr_22_26=>GND0, q_arr_22_25=>GND0, 
      q_arr_22_24=>GND0, q_arr_22_23=>GND0, q_arr_22_22=>GND0, q_arr_22_21=>
      GND0, q_arr_22_20=>GND0, q_arr_22_19=>GND0, q_arr_22_18=>GND0, 
      q_arr_22_17=>GND0, q_arr_22_16=>GND0, q_arr_22_15=>GND0, q_arr_22_14=>
      GND0, q_arr_22_13=>GND0, q_arr_22_12=>GND0, q_arr_22_11=>GND0, 
      q_arr_22_10=>GND0, q_arr_22_9=>GND0, q_arr_22_8=>GND0, q_arr_22_7=>
      GND0, q_arr_22_6=>GND0, q_arr_22_5=>GND0, q_arr_22_4=>GND0, q_arr_22_3
      =>GND0, q_arr_22_2=>GND0, q_arr_22_1=>GND0, q_arr_22_0=>GND0, 
      q_arr_23_31=>GND0, q_arr_23_30=>GND0, q_arr_23_29=>GND0, q_arr_23_28=>
      GND0, q_arr_23_27=>GND0, q_arr_23_26=>GND0, q_arr_23_25=>GND0, 
      q_arr_23_24=>GND0, q_arr_23_23=>GND0, q_arr_23_22=>GND0, q_arr_23_21=>
      GND0, q_arr_23_20=>GND0, q_arr_23_19=>GND0, q_arr_23_18=>GND0, 
      q_arr_23_17=>GND0, q_arr_23_16=>GND0, q_arr_23_15=>GND0, q_arr_23_14=>
      GND0, q_arr_23_13=>GND0, q_arr_23_12=>GND0, q_arr_23_11=>GND0, 
      q_arr_23_10=>GND0, q_arr_23_9=>GND0, q_arr_23_8=>GND0, q_arr_23_7=>
      GND0, q_arr_23_6=>GND0, q_arr_23_5=>GND0, q_arr_23_4=>GND0, q_arr_23_3
      =>GND0, q_arr_23_2=>GND0, q_arr_23_1=>GND0, q_arr_23_0=>GND0, 
      q_arr_24_31=>GND0, q_arr_24_30=>GND0, q_arr_24_29=>GND0, q_arr_24_28=>
      GND0, q_arr_24_27=>GND0, q_arr_24_26=>GND0, q_arr_24_25=>GND0, 
      q_arr_24_24=>GND0, q_arr_24_23=>GND0, q_arr_24_22=>GND0, q_arr_24_21=>
      GND0, q_arr_24_20=>GND0, q_arr_24_19=>GND0, q_arr_24_18=>GND0, 
      q_arr_24_17=>GND0, q_arr_24_16=>GND0, q_arr_24_15=>GND0, q_arr_24_14=>
      GND0, q_arr_24_13=>GND0, q_arr_24_12=>GND0, q_arr_24_11=>GND0, 
      q_arr_24_10=>GND0, q_arr_24_9=>GND0, q_arr_24_8=>GND0, q_arr_24_7=>
      GND0, q_arr_24_6=>GND0, q_arr_24_5=>GND0, q_arr_24_4=>GND0, q_arr_24_3
      =>GND0, q_arr_24_2=>GND0, q_arr_24_1=>GND0, q_arr_24_0=>GND0, 
      operation=>operation, filter_size=>nx16667);
   relu_layer_gen : ReluLayer port map ( d_arr_0_31=>d_arr_relu_0_31, 
      d_arr_0_30=>d_arr_relu_0_30, d_arr_0_29=>d_arr_relu_0_29, d_arr_0_28=>
      d_arr_relu_0_28, d_arr_0_27=>d_arr_relu_0_27, d_arr_0_26=>
      d_arr_relu_0_26, d_arr_0_25=>d_arr_relu_0_25, d_arr_0_24=>
      d_arr_relu_0_24, d_arr_0_23=>d_arr_relu_0_23, d_arr_0_22=>
      d_arr_relu_0_22, d_arr_0_21=>d_arr_relu_0_21, d_arr_0_20=>
      d_arr_relu_0_20, d_arr_0_19=>d_arr_relu_0_19, d_arr_0_18=>
      d_arr_relu_0_18, d_arr_0_17=>d_arr_relu_0_17, d_arr_0_16=>
      d_arr_relu_0_16, d_arr_0_15=>DANGLING(1952), d_arr_0_14=>
      d_arr_relu_0_14, d_arr_0_13=>d_arr_relu_0_13, d_arr_0_12=>
      d_arr_relu_0_12, d_arr_0_11=>d_arr_relu_0_11, d_arr_0_10=>
      d_arr_relu_0_10, d_arr_0_9=>d_arr_relu_0_9, d_arr_0_8=>d_arr_relu_0_8, 
      d_arr_0_7=>d_arr_relu_0_7, d_arr_0_6=>d_arr_relu_0_6, d_arr_0_5=>
      d_arr_relu_0_5, d_arr_0_4=>d_arr_relu_0_4, d_arr_0_3=>d_arr_relu_0_3, 
      d_arr_0_2=>d_arr_relu_0_2, d_arr_0_1=>d_arr_relu_0_1, d_arr_0_0=>
      d_arr_relu_0_0, d_arr_1_31=>d_arr_relu_1_31, d_arr_1_30=>
      d_arr_relu_1_30, d_arr_1_29=>d_arr_relu_1_29, d_arr_1_28=>
      d_arr_relu_1_28, d_arr_1_27=>d_arr_relu_1_27, d_arr_1_26=>
      d_arr_relu_1_26, d_arr_1_25=>d_arr_relu_1_25, d_arr_1_24=>
      d_arr_relu_1_24, d_arr_1_23=>d_arr_relu_1_23, d_arr_1_22=>
      d_arr_relu_1_22, d_arr_1_21=>d_arr_relu_1_21, d_arr_1_20=>
      d_arr_relu_1_20, d_arr_1_19=>d_arr_relu_1_19, d_arr_1_18=>
      d_arr_relu_1_18, d_arr_1_17=>d_arr_relu_1_17, d_arr_1_16=>
      d_arr_relu_1_16, d_arr_1_15=>DANGLING(1953), d_arr_1_14=>
      d_arr_relu_1_14, d_arr_1_13=>d_arr_relu_1_13, d_arr_1_12=>
      d_arr_relu_1_12, d_arr_1_11=>d_arr_relu_1_11, d_arr_1_10=>
      d_arr_relu_1_10, d_arr_1_9=>d_arr_relu_1_9, d_arr_1_8=>d_arr_relu_1_8, 
      d_arr_1_7=>d_arr_relu_1_7, d_arr_1_6=>d_arr_relu_1_6, d_arr_1_5=>
      d_arr_relu_1_5, d_arr_1_4=>d_arr_relu_1_4, d_arr_1_3=>d_arr_relu_1_3, 
      d_arr_1_2=>d_arr_relu_1_2, d_arr_1_1=>d_arr_relu_1_1, d_arr_1_0=>
      d_arr_relu_1_0, d_arr_2_31=>DANGLING(1954), d_arr_2_30=>DANGLING(1955), 
      d_arr_2_29=>DANGLING(1956), d_arr_2_28=>DANGLING(1957), d_arr_2_27=>
      DANGLING(1958), d_arr_2_26=>DANGLING(1959), d_arr_2_25=>DANGLING(1960), 
      d_arr_2_24=>DANGLING(1961), d_arr_2_23=>DANGLING(1962), d_arr_2_22=>
      DANGLING(1963), d_arr_2_21=>DANGLING(1964), d_arr_2_20=>DANGLING(1965), 
      d_arr_2_19=>DANGLING(1966), d_arr_2_18=>DANGLING(1967), d_arr_2_17=>
      DANGLING(1968), d_arr_2_16=>DANGLING(1969), d_arr_2_15=>DANGLING(1970), 
      d_arr_2_14=>DANGLING(1971), d_arr_2_13=>DANGLING(1972), d_arr_2_12=>
      DANGLING(1973), d_arr_2_11=>DANGLING(1974), d_arr_2_10=>DANGLING(1975), 
      d_arr_2_9=>DANGLING(1976), d_arr_2_8=>DANGLING(1977), d_arr_2_7=>
      DANGLING(1978), d_arr_2_6=>DANGLING(1979), d_arr_2_5=>DANGLING(1980), 
      d_arr_2_4=>DANGLING(1981), d_arr_2_3=>DANGLING(1982), d_arr_2_2=>
      DANGLING(1983), d_arr_2_1=>DANGLING(1984), d_arr_2_0=>DANGLING(1985), 
      d_arr_3_31=>DANGLING(1986), d_arr_3_30=>DANGLING(1987), d_arr_3_29=>
      DANGLING(1988), d_arr_3_28=>DANGLING(1989), d_arr_3_27=>DANGLING(1990), 
      d_arr_3_26=>DANGLING(1991), d_arr_3_25=>DANGLING(1992), d_arr_3_24=>
      DANGLING(1993), d_arr_3_23=>DANGLING(1994), d_arr_3_22=>DANGLING(1995), 
      d_arr_3_21=>DANGLING(1996), d_arr_3_20=>DANGLING(1997), d_arr_3_19=>
      DANGLING(1998), d_arr_3_18=>DANGLING(1999), d_arr_3_17=>DANGLING(2000), 
      d_arr_3_16=>DANGLING(2001), d_arr_3_15=>DANGLING(2002), d_arr_3_14=>
      DANGLING(2003), d_arr_3_13=>DANGLING(2004), d_arr_3_12=>DANGLING(2005), 
      d_arr_3_11=>DANGLING(2006), d_arr_3_10=>DANGLING(2007), d_arr_3_9=>
      DANGLING(2008), d_arr_3_8=>DANGLING(2009), d_arr_3_7=>DANGLING(2010), 
      d_arr_3_6=>DANGLING(2011), d_arr_3_5=>DANGLING(2012), d_arr_3_4=>
      DANGLING(2013), d_arr_3_3=>DANGLING(2014), d_arr_3_2=>DANGLING(2015), 
      d_arr_3_1=>DANGLING(2016), d_arr_3_0=>DANGLING(2017), d_arr_4_31=>
      DANGLING(2018), d_arr_4_30=>DANGLING(2019), d_arr_4_29=>DANGLING(2020), 
      d_arr_4_28=>DANGLING(2021), d_arr_4_27=>DANGLING(2022), d_arr_4_26=>
      DANGLING(2023), d_arr_4_25=>DANGLING(2024), d_arr_4_24=>DANGLING(2025), 
      d_arr_4_23=>DANGLING(2026), d_arr_4_22=>DANGLING(2027), d_arr_4_21=>
      DANGLING(2028), d_arr_4_20=>DANGLING(2029), d_arr_4_19=>DANGLING(2030), 
      d_arr_4_18=>DANGLING(2031), d_arr_4_17=>DANGLING(2032), d_arr_4_16=>
      DANGLING(2033), d_arr_4_15=>DANGLING(2034), d_arr_4_14=>DANGLING(2035), 
      d_arr_4_13=>DANGLING(2036), d_arr_4_12=>DANGLING(2037), d_arr_4_11=>
      DANGLING(2038), d_arr_4_10=>DANGLING(2039), d_arr_4_9=>DANGLING(2040), 
      d_arr_4_8=>DANGLING(2041), d_arr_4_7=>DANGLING(2042), d_arr_4_6=>
      DANGLING(2043), d_arr_4_5=>DANGLING(2044), d_arr_4_4=>DANGLING(2045), 
      d_arr_4_3=>DANGLING(2046), d_arr_4_2=>DANGLING(2047), d_arr_4_1=>
      DANGLING(2048), d_arr_4_0=>DANGLING(2049), d_arr_5_31=>DANGLING(2050), 
      d_arr_5_30=>DANGLING(2051), d_arr_5_29=>DANGLING(2052), d_arr_5_28=>
      DANGLING(2053), d_arr_5_27=>DANGLING(2054), d_arr_5_26=>DANGLING(2055), 
      d_arr_5_25=>DANGLING(2056), d_arr_5_24=>DANGLING(2057), d_arr_5_23=>
      DANGLING(2058), d_arr_5_22=>DANGLING(2059), d_arr_5_21=>DANGLING(2060), 
      d_arr_5_20=>DANGLING(2061), d_arr_5_19=>DANGLING(2062), d_arr_5_18=>
      DANGLING(2063), d_arr_5_17=>DANGLING(2064), d_arr_5_16=>DANGLING(2065), 
      d_arr_5_15=>DANGLING(2066), d_arr_5_14=>DANGLING(2067), d_arr_5_13=>
      DANGLING(2068), d_arr_5_12=>DANGLING(2069), d_arr_5_11=>DANGLING(2070), 
      d_arr_5_10=>DANGLING(2071), d_arr_5_9=>DANGLING(2072), d_arr_5_8=>
      DANGLING(2073), d_arr_5_7=>DANGLING(2074), d_arr_5_6=>DANGLING(2075), 
      d_arr_5_5=>DANGLING(2076), d_arr_5_4=>DANGLING(2077), d_arr_5_3=>
      DANGLING(2078), d_arr_5_2=>DANGLING(2079), d_arr_5_1=>DANGLING(2080), 
      d_arr_5_0=>DANGLING(2081), d_arr_6_31=>DANGLING(2082), d_arr_6_30=>
      DANGLING(2083), d_arr_6_29=>DANGLING(2084), d_arr_6_28=>DANGLING(2085), 
      d_arr_6_27=>DANGLING(2086), d_arr_6_26=>DANGLING(2087), d_arr_6_25=>
      DANGLING(2088), d_arr_6_24=>DANGLING(2089), d_arr_6_23=>DANGLING(2090), 
      d_arr_6_22=>DANGLING(2091), d_arr_6_21=>DANGLING(2092), d_arr_6_20=>
      DANGLING(2093), d_arr_6_19=>DANGLING(2094), d_arr_6_18=>DANGLING(2095), 
      d_arr_6_17=>DANGLING(2096), d_arr_6_16=>DANGLING(2097), d_arr_6_15=>
      DANGLING(2098), d_arr_6_14=>DANGLING(2099), d_arr_6_13=>DANGLING(2100), 
      d_arr_6_12=>DANGLING(2101), d_arr_6_11=>DANGLING(2102), d_arr_6_10=>
      DANGLING(2103), d_arr_6_9=>DANGLING(2104), d_arr_6_8=>DANGLING(2105), 
      d_arr_6_7=>DANGLING(2106), d_arr_6_6=>DANGLING(2107), d_arr_6_5=>
      DANGLING(2108), d_arr_6_4=>DANGLING(2109), d_arr_6_3=>DANGLING(2110), 
      d_arr_6_2=>DANGLING(2111), d_arr_6_1=>DANGLING(2112), d_arr_6_0=>
      DANGLING(2113), d_arr_7_31=>DANGLING(2114), d_arr_7_30=>DANGLING(2115), 
      d_arr_7_29=>DANGLING(2116), d_arr_7_28=>DANGLING(2117), d_arr_7_27=>
      DANGLING(2118), d_arr_7_26=>DANGLING(2119), d_arr_7_25=>DANGLING(2120), 
      d_arr_7_24=>DANGLING(2121), d_arr_7_23=>DANGLING(2122), d_arr_7_22=>
      DANGLING(2123), d_arr_7_21=>DANGLING(2124), d_arr_7_20=>DANGLING(2125), 
      d_arr_7_19=>DANGLING(2126), d_arr_7_18=>DANGLING(2127), d_arr_7_17=>
      DANGLING(2128), d_arr_7_16=>DANGLING(2129), d_arr_7_15=>DANGLING(2130), 
      d_arr_7_14=>DANGLING(2131), d_arr_7_13=>DANGLING(2132), d_arr_7_12=>
      DANGLING(2133), d_arr_7_11=>DANGLING(2134), d_arr_7_10=>DANGLING(2135), 
      d_arr_7_9=>DANGLING(2136), d_arr_7_8=>DANGLING(2137), d_arr_7_7=>
      DANGLING(2138), d_arr_7_6=>DANGLING(2139), d_arr_7_5=>DANGLING(2140), 
      d_arr_7_4=>DANGLING(2141), d_arr_7_3=>DANGLING(2142), d_arr_7_2=>
      DANGLING(2143), d_arr_7_1=>DANGLING(2144), d_arr_7_0=>DANGLING(2145), 
      d_arr_8_31=>DANGLING(2146), d_arr_8_30=>DANGLING(2147), d_arr_8_29=>
      DANGLING(2148), d_arr_8_28=>DANGLING(2149), d_arr_8_27=>DANGLING(2150), 
      d_arr_8_26=>DANGLING(2151), d_arr_8_25=>DANGLING(2152), d_arr_8_24=>
      DANGLING(2153), d_arr_8_23=>DANGLING(2154), d_arr_8_22=>DANGLING(2155), 
      d_arr_8_21=>DANGLING(2156), d_arr_8_20=>DANGLING(2157), d_arr_8_19=>
      DANGLING(2158), d_arr_8_18=>DANGLING(2159), d_arr_8_17=>DANGLING(2160), 
      d_arr_8_16=>DANGLING(2161), d_arr_8_15=>DANGLING(2162), d_arr_8_14=>
      DANGLING(2163), d_arr_8_13=>DANGLING(2164), d_arr_8_12=>DANGLING(2165), 
      d_arr_8_11=>DANGLING(2166), d_arr_8_10=>DANGLING(2167), d_arr_8_9=>
      DANGLING(2168), d_arr_8_8=>DANGLING(2169), d_arr_8_7=>DANGLING(2170), 
      d_arr_8_6=>DANGLING(2171), d_arr_8_5=>DANGLING(2172), d_arr_8_4=>
      DANGLING(2173), d_arr_8_3=>DANGLING(2174), d_arr_8_2=>DANGLING(2175), 
      d_arr_8_1=>DANGLING(2176), d_arr_8_0=>DANGLING(2177), d_arr_9_31=>
      DANGLING(2178), d_arr_9_30=>DANGLING(2179), d_arr_9_29=>DANGLING(2180), 
      d_arr_9_28=>DANGLING(2181), d_arr_9_27=>DANGLING(2182), d_arr_9_26=>
      DANGLING(2183), d_arr_9_25=>DANGLING(2184), d_arr_9_24=>DANGLING(2185), 
      d_arr_9_23=>DANGLING(2186), d_arr_9_22=>DANGLING(2187), d_arr_9_21=>
      DANGLING(2188), d_arr_9_20=>DANGLING(2189), d_arr_9_19=>DANGLING(2190), 
      d_arr_9_18=>DANGLING(2191), d_arr_9_17=>DANGLING(2192), d_arr_9_16=>
      DANGLING(2193), d_arr_9_15=>DANGLING(2194), d_arr_9_14=>DANGLING(2195), 
      d_arr_9_13=>DANGLING(2196), d_arr_9_12=>DANGLING(2197), d_arr_9_11=>
      DANGLING(2198), d_arr_9_10=>DANGLING(2199), d_arr_9_9=>DANGLING(2200), 
      d_arr_9_8=>DANGLING(2201), d_arr_9_7=>DANGLING(2202), d_arr_9_6=>
      DANGLING(2203), d_arr_9_5=>DANGLING(2204), d_arr_9_4=>DANGLING(2205), 
      d_arr_9_3=>DANGLING(2206), d_arr_9_2=>DANGLING(2207), d_arr_9_1=>
      DANGLING(2208), d_arr_9_0=>DANGLING(2209), d_arr_10_31=>DANGLING(2210), 
      d_arr_10_30=>DANGLING(2211), d_arr_10_29=>DANGLING(2212), d_arr_10_28
      =>DANGLING(2213), d_arr_10_27=>DANGLING(2214), d_arr_10_26=>DANGLING(
      2215), d_arr_10_25=>DANGLING(2216), d_arr_10_24=>DANGLING(2217), 
      d_arr_10_23=>DANGLING(2218), d_arr_10_22=>DANGLING(2219), d_arr_10_21
      =>DANGLING(2220), d_arr_10_20=>DANGLING(2221), d_arr_10_19=>DANGLING(
      2222), d_arr_10_18=>DANGLING(2223), d_arr_10_17=>DANGLING(2224), 
      d_arr_10_16=>DANGLING(2225), d_arr_10_15=>DANGLING(2226), d_arr_10_14
      =>DANGLING(2227), d_arr_10_13=>DANGLING(2228), d_arr_10_12=>DANGLING(
      2229), d_arr_10_11=>DANGLING(2230), d_arr_10_10=>DANGLING(2231), 
      d_arr_10_9=>DANGLING(2232), d_arr_10_8=>DANGLING(2233), d_arr_10_7=>
      DANGLING(2234), d_arr_10_6=>DANGLING(2235), d_arr_10_5=>DANGLING(2236), 
      d_arr_10_4=>DANGLING(2237), d_arr_10_3=>DANGLING(2238), d_arr_10_2=>
      DANGLING(2239), d_arr_10_1=>DANGLING(2240), d_arr_10_0=>DANGLING(2241), 
      d_arr_11_31=>DANGLING(2242), d_arr_11_30=>DANGLING(2243), d_arr_11_29
      =>DANGLING(2244), d_arr_11_28=>DANGLING(2245), d_arr_11_27=>DANGLING(
      2246), d_arr_11_26=>DANGLING(2247), d_arr_11_25=>DANGLING(2248), 
      d_arr_11_24=>DANGLING(2249), d_arr_11_23=>DANGLING(2250), d_arr_11_22
      =>DANGLING(2251), d_arr_11_21=>DANGLING(2252), d_arr_11_20=>DANGLING(
      2253), d_arr_11_19=>DANGLING(2254), d_arr_11_18=>DANGLING(2255), 
      d_arr_11_17=>DANGLING(2256), d_arr_11_16=>DANGLING(2257), d_arr_11_15
      =>DANGLING(2258), d_arr_11_14=>DANGLING(2259), d_arr_11_13=>DANGLING(
      2260), d_arr_11_12=>DANGLING(2261), d_arr_11_11=>DANGLING(2262), 
      d_arr_11_10=>DANGLING(2263), d_arr_11_9=>DANGLING(2264), d_arr_11_8=>
      DANGLING(2265), d_arr_11_7=>DANGLING(2266), d_arr_11_6=>DANGLING(2267), 
      d_arr_11_5=>DANGLING(2268), d_arr_11_4=>DANGLING(2269), d_arr_11_3=>
      DANGLING(2270), d_arr_11_2=>DANGLING(2271), d_arr_11_1=>DANGLING(2272), 
      d_arr_11_0=>DANGLING(2273), d_arr_12_31=>DANGLING(2274), d_arr_12_30=>
      DANGLING(2275), d_arr_12_29=>DANGLING(2276), d_arr_12_28=>DANGLING(
      2277), d_arr_12_27=>DANGLING(2278), d_arr_12_26=>DANGLING(2279), 
      d_arr_12_25=>DANGLING(2280), d_arr_12_24=>DANGLING(2281), d_arr_12_23
      =>DANGLING(2282), d_arr_12_22=>DANGLING(2283), d_arr_12_21=>DANGLING(
      2284), d_arr_12_20=>DANGLING(2285), d_arr_12_19=>DANGLING(2286), 
      d_arr_12_18=>DANGLING(2287), d_arr_12_17=>DANGLING(2288), d_arr_12_16
      =>DANGLING(2289), d_arr_12_15=>DANGLING(2290), d_arr_12_14=>DANGLING(
      2291), d_arr_12_13=>DANGLING(2292), d_arr_12_12=>DANGLING(2293), 
      d_arr_12_11=>DANGLING(2294), d_arr_12_10=>DANGLING(2295), d_arr_12_9=>
      DANGLING(2296), d_arr_12_8=>DANGLING(2297), d_arr_12_7=>DANGLING(2298), 
      d_arr_12_6=>DANGLING(2299), d_arr_12_5=>DANGLING(2300), d_arr_12_4=>
      DANGLING(2301), d_arr_12_3=>DANGLING(2302), d_arr_12_2=>DANGLING(2303), 
      d_arr_12_1=>DANGLING(2304), d_arr_12_0=>DANGLING(2305), d_arr_13_31=>
      DANGLING(2306), d_arr_13_30=>DANGLING(2307), d_arr_13_29=>DANGLING(
      2308), d_arr_13_28=>DANGLING(2309), d_arr_13_27=>DANGLING(2310), 
      d_arr_13_26=>DANGLING(2311), d_arr_13_25=>DANGLING(2312), d_arr_13_24
      =>DANGLING(2313), d_arr_13_23=>DANGLING(2314), d_arr_13_22=>DANGLING(
      2315), d_arr_13_21=>DANGLING(2316), d_arr_13_20=>DANGLING(2317), 
      d_arr_13_19=>DANGLING(2318), d_arr_13_18=>DANGLING(2319), d_arr_13_17
      =>DANGLING(2320), d_arr_13_16=>DANGLING(2321), d_arr_13_15=>DANGLING(
      2322), d_arr_13_14=>DANGLING(2323), d_arr_13_13=>DANGLING(2324), 
      d_arr_13_12=>DANGLING(2325), d_arr_13_11=>DANGLING(2326), d_arr_13_10
      =>DANGLING(2327), d_arr_13_9=>DANGLING(2328), d_arr_13_8=>DANGLING(
      2329), d_arr_13_7=>DANGLING(2330), d_arr_13_6=>DANGLING(2331), 
      d_arr_13_5=>DANGLING(2332), d_arr_13_4=>DANGLING(2333), d_arr_13_3=>
      DANGLING(2334), d_arr_13_2=>DANGLING(2335), d_arr_13_1=>DANGLING(2336), 
      d_arr_13_0=>DANGLING(2337), d_arr_14_31=>DANGLING(2338), d_arr_14_30=>
      DANGLING(2339), d_arr_14_29=>DANGLING(2340), d_arr_14_28=>DANGLING(
      2341), d_arr_14_27=>DANGLING(2342), d_arr_14_26=>DANGLING(2343), 
      d_arr_14_25=>DANGLING(2344), d_arr_14_24=>DANGLING(2345), d_arr_14_23
      =>DANGLING(2346), d_arr_14_22=>DANGLING(2347), d_arr_14_21=>DANGLING(
      2348), d_arr_14_20=>DANGLING(2349), d_arr_14_19=>DANGLING(2350), 
      d_arr_14_18=>DANGLING(2351), d_arr_14_17=>DANGLING(2352), d_arr_14_16
      =>DANGLING(2353), d_arr_14_15=>DANGLING(2354), d_arr_14_14=>DANGLING(
      2355), d_arr_14_13=>DANGLING(2356), d_arr_14_12=>DANGLING(2357), 
      d_arr_14_11=>DANGLING(2358), d_arr_14_10=>DANGLING(2359), d_arr_14_9=>
      DANGLING(2360), d_arr_14_8=>DANGLING(2361), d_arr_14_7=>DANGLING(2362), 
      d_arr_14_6=>DANGLING(2363), d_arr_14_5=>DANGLING(2364), d_arr_14_4=>
      DANGLING(2365), d_arr_14_3=>DANGLING(2366), d_arr_14_2=>DANGLING(2367), 
      d_arr_14_1=>DANGLING(2368), d_arr_14_0=>DANGLING(2369), d_arr_15_31=>
      DANGLING(2370), d_arr_15_30=>DANGLING(2371), d_arr_15_29=>DANGLING(
      2372), d_arr_15_28=>DANGLING(2373), d_arr_15_27=>DANGLING(2374), 
      d_arr_15_26=>DANGLING(2375), d_arr_15_25=>DANGLING(2376), d_arr_15_24
      =>DANGLING(2377), d_arr_15_23=>DANGLING(2378), d_arr_15_22=>DANGLING(
      2379), d_arr_15_21=>DANGLING(2380), d_arr_15_20=>DANGLING(2381), 
      d_arr_15_19=>DANGLING(2382), d_arr_15_18=>DANGLING(2383), d_arr_15_17
      =>DANGLING(2384), d_arr_15_16=>DANGLING(2385), d_arr_15_15=>DANGLING(
      2386), d_arr_15_14=>DANGLING(2387), d_arr_15_13=>DANGLING(2388), 
      d_arr_15_12=>DANGLING(2389), d_arr_15_11=>DANGLING(2390), d_arr_15_10
      =>DANGLING(2391), d_arr_15_9=>DANGLING(2392), d_arr_15_8=>DANGLING(
      2393), d_arr_15_7=>DANGLING(2394), d_arr_15_6=>DANGLING(2395), 
      d_arr_15_5=>DANGLING(2396), d_arr_15_4=>DANGLING(2397), d_arr_15_3=>
      DANGLING(2398), d_arr_15_2=>DANGLING(2399), d_arr_15_1=>DANGLING(2400), 
      d_arr_15_0=>DANGLING(2401), d_arr_16_31=>DANGLING(2402), d_arr_16_30=>
      DANGLING(2403), d_arr_16_29=>DANGLING(2404), d_arr_16_28=>DANGLING(
      2405), d_arr_16_27=>DANGLING(2406), d_arr_16_26=>DANGLING(2407), 
      d_arr_16_25=>DANGLING(2408), d_arr_16_24=>DANGLING(2409), d_arr_16_23
      =>DANGLING(2410), d_arr_16_22=>DANGLING(2411), d_arr_16_21=>DANGLING(
      2412), d_arr_16_20=>DANGLING(2413), d_arr_16_19=>DANGLING(2414), 
      d_arr_16_18=>DANGLING(2415), d_arr_16_17=>DANGLING(2416), d_arr_16_16
      =>DANGLING(2417), d_arr_16_15=>DANGLING(2418), d_arr_16_14=>DANGLING(
      2419), d_arr_16_13=>DANGLING(2420), d_arr_16_12=>DANGLING(2421), 
      d_arr_16_11=>DANGLING(2422), d_arr_16_10=>DANGLING(2423), d_arr_16_9=>
      DANGLING(2424), d_arr_16_8=>DANGLING(2425), d_arr_16_7=>DANGLING(2426), 
      d_arr_16_6=>DANGLING(2427), d_arr_16_5=>DANGLING(2428), d_arr_16_4=>
      DANGLING(2429), d_arr_16_3=>DANGLING(2430), d_arr_16_2=>DANGLING(2431), 
      d_arr_16_1=>DANGLING(2432), d_arr_16_0=>DANGLING(2433), d_arr_17_31=>
      DANGLING(2434), d_arr_17_30=>DANGLING(2435), d_arr_17_29=>DANGLING(
      2436), d_arr_17_28=>DANGLING(2437), d_arr_17_27=>DANGLING(2438), 
      d_arr_17_26=>DANGLING(2439), d_arr_17_25=>DANGLING(2440), d_arr_17_24
      =>DANGLING(2441), d_arr_17_23=>DANGLING(2442), d_arr_17_22=>DANGLING(
      2443), d_arr_17_21=>DANGLING(2444), d_arr_17_20=>DANGLING(2445), 
      d_arr_17_19=>DANGLING(2446), d_arr_17_18=>DANGLING(2447), d_arr_17_17
      =>DANGLING(2448), d_arr_17_16=>DANGLING(2449), d_arr_17_15=>DANGLING(
      2450), d_arr_17_14=>DANGLING(2451), d_arr_17_13=>DANGLING(2452), 
      d_arr_17_12=>DANGLING(2453), d_arr_17_11=>DANGLING(2454), d_arr_17_10
      =>DANGLING(2455), d_arr_17_9=>DANGLING(2456), d_arr_17_8=>DANGLING(
      2457), d_arr_17_7=>DANGLING(2458), d_arr_17_6=>DANGLING(2459), 
      d_arr_17_5=>DANGLING(2460), d_arr_17_4=>DANGLING(2461), d_arr_17_3=>
      DANGLING(2462), d_arr_17_2=>DANGLING(2463), d_arr_17_1=>DANGLING(2464), 
      d_arr_17_0=>DANGLING(2465), d_arr_18_31=>DANGLING(2466), d_arr_18_30=>
      DANGLING(2467), d_arr_18_29=>DANGLING(2468), d_arr_18_28=>DANGLING(
      2469), d_arr_18_27=>DANGLING(2470), d_arr_18_26=>DANGLING(2471), 
      d_arr_18_25=>DANGLING(2472), d_arr_18_24=>DANGLING(2473), d_arr_18_23
      =>DANGLING(2474), d_arr_18_22=>DANGLING(2475), d_arr_18_21=>DANGLING(
      2476), d_arr_18_20=>DANGLING(2477), d_arr_18_19=>DANGLING(2478), 
      d_arr_18_18=>DANGLING(2479), d_arr_18_17=>DANGLING(2480), d_arr_18_16
      =>DANGLING(2481), d_arr_18_15=>DANGLING(2482), d_arr_18_14=>DANGLING(
      2483), d_arr_18_13=>DANGLING(2484), d_arr_18_12=>DANGLING(2485), 
      d_arr_18_11=>DANGLING(2486), d_arr_18_10=>DANGLING(2487), d_arr_18_9=>
      DANGLING(2488), d_arr_18_8=>DANGLING(2489), d_arr_18_7=>DANGLING(2490), 
      d_arr_18_6=>DANGLING(2491), d_arr_18_5=>DANGLING(2492), d_arr_18_4=>
      DANGLING(2493), d_arr_18_3=>DANGLING(2494), d_arr_18_2=>DANGLING(2495), 
      d_arr_18_1=>DANGLING(2496), d_arr_18_0=>DANGLING(2497), d_arr_19_31=>
      DANGLING(2498), d_arr_19_30=>DANGLING(2499), d_arr_19_29=>DANGLING(
      2500), d_arr_19_28=>DANGLING(2501), d_arr_19_27=>DANGLING(2502), 
      d_arr_19_26=>DANGLING(2503), d_arr_19_25=>DANGLING(2504), d_arr_19_24
      =>DANGLING(2505), d_arr_19_23=>DANGLING(2506), d_arr_19_22=>DANGLING(
      2507), d_arr_19_21=>DANGLING(2508), d_arr_19_20=>DANGLING(2509), 
      d_arr_19_19=>DANGLING(2510), d_arr_19_18=>DANGLING(2511), d_arr_19_17
      =>DANGLING(2512), d_arr_19_16=>DANGLING(2513), d_arr_19_15=>DANGLING(
      2514), d_arr_19_14=>DANGLING(2515), d_arr_19_13=>DANGLING(2516), 
      d_arr_19_12=>DANGLING(2517), d_arr_19_11=>DANGLING(2518), d_arr_19_10
      =>DANGLING(2519), d_arr_19_9=>DANGLING(2520), d_arr_19_8=>DANGLING(
      2521), d_arr_19_7=>DANGLING(2522), d_arr_19_6=>DANGLING(2523), 
      d_arr_19_5=>DANGLING(2524), d_arr_19_4=>DANGLING(2525), d_arr_19_3=>
      DANGLING(2526), d_arr_19_2=>DANGLING(2527), d_arr_19_1=>DANGLING(2528), 
      d_arr_19_0=>DANGLING(2529), d_arr_20_31=>DANGLING(2530), d_arr_20_30=>
      DANGLING(2531), d_arr_20_29=>DANGLING(2532), d_arr_20_28=>DANGLING(
      2533), d_arr_20_27=>DANGLING(2534), d_arr_20_26=>DANGLING(2535), 
      d_arr_20_25=>DANGLING(2536), d_arr_20_24=>DANGLING(2537), d_arr_20_23
      =>DANGLING(2538), d_arr_20_22=>DANGLING(2539), d_arr_20_21=>DANGLING(
      2540), d_arr_20_20=>DANGLING(2541), d_arr_20_19=>DANGLING(2542), 
      d_arr_20_18=>DANGLING(2543), d_arr_20_17=>DANGLING(2544), d_arr_20_16
      =>DANGLING(2545), d_arr_20_15=>DANGLING(2546), d_arr_20_14=>DANGLING(
      2547), d_arr_20_13=>DANGLING(2548), d_arr_20_12=>DANGLING(2549), 
      d_arr_20_11=>DANGLING(2550), d_arr_20_10=>DANGLING(2551), d_arr_20_9=>
      DANGLING(2552), d_arr_20_8=>DANGLING(2553), d_arr_20_7=>DANGLING(2554), 
      d_arr_20_6=>DANGLING(2555), d_arr_20_5=>DANGLING(2556), d_arr_20_4=>
      DANGLING(2557), d_arr_20_3=>DANGLING(2558), d_arr_20_2=>DANGLING(2559), 
      d_arr_20_1=>DANGLING(2560), d_arr_20_0=>DANGLING(2561), d_arr_21_31=>
      DANGLING(2562), d_arr_21_30=>DANGLING(2563), d_arr_21_29=>DANGLING(
      2564), d_arr_21_28=>DANGLING(2565), d_arr_21_27=>DANGLING(2566), 
      d_arr_21_26=>DANGLING(2567), d_arr_21_25=>DANGLING(2568), d_arr_21_24
      =>DANGLING(2569), d_arr_21_23=>DANGLING(2570), d_arr_21_22=>DANGLING(
      2571), d_arr_21_21=>DANGLING(2572), d_arr_21_20=>DANGLING(2573), 
      d_arr_21_19=>DANGLING(2574), d_arr_21_18=>DANGLING(2575), d_arr_21_17
      =>DANGLING(2576), d_arr_21_16=>DANGLING(2577), d_arr_21_15=>DANGLING(
      2578), d_arr_21_14=>DANGLING(2579), d_arr_21_13=>DANGLING(2580), 
      d_arr_21_12=>DANGLING(2581), d_arr_21_11=>DANGLING(2582), d_arr_21_10
      =>DANGLING(2583), d_arr_21_9=>DANGLING(2584), d_arr_21_8=>DANGLING(
      2585), d_arr_21_7=>DANGLING(2586), d_arr_21_6=>DANGLING(2587), 
      d_arr_21_5=>DANGLING(2588), d_arr_21_4=>DANGLING(2589), d_arr_21_3=>
      DANGLING(2590), d_arr_21_2=>DANGLING(2591), d_arr_21_1=>DANGLING(2592), 
      d_arr_21_0=>DANGLING(2593), d_arr_22_31=>DANGLING(2594), d_arr_22_30=>
      DANGLING(2595), d_arr_22_29=>DANGLING(2596), d_arr_22_28=>DANGLING(
      2597), d_arr_22_27=>DANGLING(2598), d_arr_22_26=>DANGLING(2599), 
      d_arr_22_25=>DANGLING(2600), d_arr_22_24=>DANGLING(2601), d_arr_22_23
      =>DANGLING(2602), d_arr_22_22=>DANGLING(2603), d_arr_22_21=>DANGLING(
      2604), d_arr_22_20=>DANGLING(2605), d_arr_22_19=>DANGLING(2606), 
      d_arr_22_18=>DANGLING(2607), d_arr_22_17=>DANGLING(2608), d_arr_22_16
      =>DANGLING(2609), d_arr_22_15=>DANGLING(2610), d_arr_22_14=>DANGLING(
      2611), d_arr_22_13=>DANGLING(2612), d_arr_22_12=>DANGLING(2613), 
      d_arr_22_11=>DANGLING(2614), d_arr_22_10=>DANGLING(2615), d_arr_22_9=>
      DANGLING(2616), d_arr_22_8=>DANGLING(2617), d_arr_22_7=>DANGLING(2618), 
      d_arr_22_6=>DANGLING(2619), d_arr_22_5=>DANGLING(2620), d_arr_22_4=>
      DANGLING(2621), d_arr_22_3=>DANGLING(2622), d_arr_22_2=>DANGLING(2623), 
      d_arr_22_1=>DANGLING(2624), d_arr_22_0=>DANGLING(2625), d_arr_23_31=>
      DANGLING(2626), d_arr_23_30=>DANGLING(2627), d_arr_23_29=>DANGLING(
      2628), d_arr_23_28=>DANGLING(2629), d_arr_23_27=>DANGLING(2630), 
      d_arr_23_26=>DANGLING(2631), d_arr_23_25=>DANGLING(2632), d_arr_23_24
      =>DANGLING(2633), d_arr_23_23=>DANGLING(2634), d_arr_23_22=>DANGLING(
      2635), d_arr_23_21=>DANGLING(2636), d_arr_23_20=>DANGLING(2637), 
      d_arr_23_19=>DANGLING(2638), d_arr_23_18=>DANGLING(2639), d_arr_23_17
      =>DANGLING(2640), d_arr_23_16=>DANGLING(2641), d_arr_23_15=>DANGLING(
      2642), d_arr_23_14=>DANGLING(2643), d_arr_23_13=>DANGLING(2644), 
      d_arr_23_12=>DANGLING(2645), d_arr_23_11=>DANGLING(2646), d_arr_23_10
      =>DANGLING(2647), d_arr_23_9=>DANGLING(2648), d_arr_23_8=>DANGLING(
      2649), d_arr_23_7=>DANGLING(2650), d_arr_23_6=>DANGLING(2651), 
      d_arr_23_5=>DANGLING(2652), d_arr_23_4=>DANGLING(2653), d_arr_23_3=>
      DANGLING(2654), d_arr_23_2=>DANGLING(2655), d_arr_23_1=>DANGLING(2656), 
      d_arr_23_0=>DANGLING(2657), d_arr_24_31=>DANGLING(2658), d_arr_24_30=>
      DANGLING(2659), d_arr_24_29=>DANGLING(2660), d_arr_24_28=>DANGLING(
      2661), d_arr_24_27=>DANGLING(2662), d_arr_24_26=>DANGLING(2663), 
      d_arr_24_25=>DANGLING(2664), d_arr_24_24=>DANGLING(2665), d_arr_24_23
      =>DANGLING(2666), d_arr_24_22=>DANGLING(2667), d_arr_24_21=>DANGLING(
      2668), d_arr_24_20=>DANGLING(2669), d_arr_24_19=>DANGLING(2670), 
      d_arr_24_18=>DANGLING(2671), d_arr_24_17=>DANGLING(2672), d_arr_24_16
      =>DANGLING(2673), d_arr_24_15=>DANGLING(2674), d_arr_24_14=>DANGLING(
      2675), d_arr_24_13=>DANGLING(2676), d_arr_24_12=>DANGLING(2677), 
      d_arr_24_11=>DANGLING(2678), d_arr_24_10=>DANGLING(2679), d_arr_24_9=>
      DANGLING(2680), d_arr_24_8=>DANGLING(2681), d_arr_24_7=>DANGLING(2682), 
      d_arr_24_6=>DANGLING(2683), d_arr_24_5=>DANGLING(2684), d_arr_24_4=>
      DANGLING(2685), d_arr_24_3=>DANGLING(2686), d_arr_24_2=>DANGLING(2687), 
      d_arr_24_1=>DANGLING(2688), d_arr_24_0=>DANGLING(2689), q_arr_0_31=>
      nx19448, q_arr_0_30=>nx16499, q_arr_0_29=>nx16503, q_arr_0_28=>nx16507, 
      q_arr_0_27=>nx16511, q_arr_0_26=>nx16515, q_arr_0_25=>nx16519, 
      q_arr_0_24=>nx19390, q_arr_0_23=>nx16527, q_arr_0_22=>nx16531, 
      q_arr_0_21=>nx16535, q_arr_0_20=>nx16539, q_arr_0_19=>nx16543, 
      q_arr_0_18=>nx16547, q_arr_0_17=>nx16551, q_arr_0_16=>nx16555, 
      q_arr_0_15=>nx16559, q_arr_0_14=>nx16563, q_arr_0_13=>nx16567, 
      q_arr_0_12=>nx16571, q_arr_0_11=>nx16575, q_arr_0_10=>nx16579, 
      q_arr_0_9=>nx16583, q_arr_0_8=>nx16587, q_arr_0_7=>nx16591, q_arr_0_6
      =>nx16595, q_arr_0_5=>nx16599, q_arr_0_4=>nx16601, q_arr_0_3=>nx16603, 
      q_arr_0_2=>q_arr_0_2, q_arr_0_1=>q_arr_0_1, q_arr_0_0=>nx16605, 
      q_arr_1_31=>q_arr_1_31, q_arr_1_30=>q_arr_1_30, q_arr_1_29=>q_arr_1_29, 
      q_arr_1_28=>q_arr_1_28, q_arr_1_27=>nx19450, q_arr_1_26=>nx19454, 
      q_arr_1_25=>q_arr_1_25, q_arr_1_24=>nx19458, q_arr_1_23=>q_arr_1_23, 
      q_arr_1_22=>q_arr_1_22, q_arr_1_21=>q_arr_1_21, q_arr_1_20=>q_arr_1_20, 
      q_arr_1_19=>q_arr_1_19, q_arr_1_18=>nx19462, q_arr_1_17=>nx19466, 
      q_arr_1_16=>nx19470, q_arr_1_15=>q_arr_1_15, q_arr_1_14=>nx19474, 
      q_arr_1_13=>q_arr_1_13, q_arr_1_12=>nx19476, q_arr_1_11=>q_arr_1_11, 
      q_arr_1_10=>nx19478, q_arr_1_9=>q_arr_1_9, q_arr_1_8=>nx19482, 
      q_arr_1_7=>nx19486, q_arr_1_6=>q_arr_1_6, q_arr_1_5=>q_arr_1_5, 
      q_arr_1_4=>q_arr_1_4, q_arr_1_3=>q_arr_1_3, q_arr_1_2=>q_arr_1_2, 
      q_arr_1_1=>q_arr_1_1, q_arr_1_0=>q_arr_1_0, q_arr_2_31=>GND0, 
      q_arr_2_30=>GND0, q_arr_2_29=>GND0, q_arr_2_28=>GND0, q_arr_2_27=>GND0, 
      q_arr_2_26=>GND0, q_arr_2_25=>GND0, q_arr_2_24=>GND0, q_arr_2_23=>GND0, 
      q_arr_2_22=>GND0, q_arr_2_21=>GND0, q_arr_2_20=>GND0, q_arr_2_19=>GND0, 
      q_arr_2_18=>GND0, q_arr_2_17=>GND0, q_arr_2_16=>GND0, q_arr_2_15=>GND0, 
      q_arr_2_14=>GND0, q_arr_2_13=>GND0, q_arr_2_12=>GND0, q_arr_2_11=>GND0, 
      q_arr_2_10=>GND0, q_arr_2_9=>GND0, q_arr_2_8=>GND0, q_arr_2_7=>GND0, 
      q_arr_2_6=>GND0, q_arr_2_5=>GND0, q_arr_2_4=>GND0, q_arr_2_3=>GND0, 
      q_arr_2_2=>GND0, q_arr_2_1=>GND0, q_arr_2_0=>GND0, q_arr_3_31=>GND0, 
      q_arr_3_30=>GND0, q_arr_3_29=>GND0, q_arr_3_28=>GND0, q_arr_3_27=>GND0, 
      q_arr_3_26=>GND0, q_arr_3_25=>GND0, q_arr_3_24=>GND0, q_arr_3_23=>GND0, 
      q_arr_3_22=>GND0, q_arr_3_21=>GND0, q_arr_3_20=>GND0, q_arr_3_19=>GND0, 
      q_arr_3_18=>GND0, q_arr_3_17=>GND0, q_arr_3_16=>GND0, q_arr_3_15=>GND0, 
      q_arr_3_14=>GND0, q_arr_3_13=>GND0, q_arr_3_12=>GND0, q_arr_3_11=>GND0, 
      q_arr_3_10=>GND0, q_arr_3_9=>GND0, q_arr_3_8=>GND0, q_arr_3_7=>GND0, 
      q_arr_3_6=>GND0, q_arr_3_5=>GND0, q_arr_3_4=>GND0, q_arr_3_3=>GND0, 
      q_arr_3_2=>GND0, q_arr_3_1=>GND0, q_arr_3_0=>GND0, q_arr_4_31=>GND0, 
      q_arr_4_30=>GND0, q_arr_4_29=>GND0, q_arr_4_28=>GND0, q_arr_4_27=>GND0, 
      q_arr_4_26=>GND0, q_arr_4_25=>GND0, q_arr_4_24=>GND0, q_arr_4_23=>GND0, 
      q_arr_4_22=>GND0, q_arr_4_21=>GND0, q_arr_4_20=>GND0, q_arr_4_19=>GND0, 
      q_arr_4_18=>GND0, q_arr_4_17=>GND0, q_arr_4_16=>GND0, q_arr_4_15=>GND0, 
      q_arr_4_14=>GND0, q_arr_4_13=>GND0, q_arr_4_12=>GND0, q_arr_4_11=>GND0, 
      q_arr_4_10=>GND0, q_arr_4_9=>GND0, q_arr_4_8=>GND0, q_arr_4_7=>GND0, 
      q_arr_4_6=>GND0, q_arr_4_5=>GND0, q_arr_4_4=>GND0, q_arr_4_3=>GND0, 
      q_arr_4_2=>GND0, q_arr_4_1=>GND0, q_arr_4_0=>GND0, q_arr_5_31=>GND0, 
      q_arr_5_30=>GND0, q_arr_5_29=>GND0, q_arr_5_28=>GND0, q_arr_5_27=>GND0, 
      q_arr_5_26=>GND0, q_arr_5_25=>GND0, q_arr_5_24=>GND0, q_arr_5_23=>GND0, 
      q_arr_5_22=>GND0, q_arr_5_21=>GND0, q_arr_5_20=>GND0, q_arr_5_19=>GND0, 
      q_arr_5_18=>GND0, q_arr_5_17=>GND0, q_arr_5_16=>GND0, q_arr_5_15=>GND0, 
      q_arr_5_14=>GND0, q_arr_5_13=>GND0, q_arr_5_12=>GND0, q_arr_5_11=>GND0, 
      q_arr_5_10=>GND0, q_arr_5_9=>GND0, q_arr_5_8=>GND0, q_arr_5_7=>GND0, 
      q_arr_5_6=>GND0, q_arr_5_5=>GND0, q_arr_5_4=>GND0, q_arr_5_3=>GND0, 
      q_arr_5_2=>GND0, q_arr_5_1=>GND0, q_arr_5_0=>GND0, q_arr_6_31=>GND0, 
      q_arr_6_30=>GND0, q_arr_6_29=>GND0, q_arr_6_28=>GND0, q_arr_6_27=>GND0, 
      q_arr_6_26=>GND0, q_arr_6_25=>GND0, q_arr_6_24=>GND0, q_arr_6_23=>GND0, 
      q_arr_6_22=>GND0, q_arr_6_21=>GND0, q_arr_6_20=>GND0, q_arr_6_19=>GND0, 
      q_arr_6_18=>GND0, q_arr_6_17=>GND0, q_arr_6_16=>GND0, q_arr_6_15=>GND0, 
      q_arr_6_14=>GND0, q_arr_6_13=>GND0, q_arr_6_12=>GND0, q_arr_6_11=>GND0, 
      q_arr_6_10=>GND0, q_arr_6_9=>GND0, q_arr_6_8=>GND0, q_arr_6_7=>GND0, 
      q_arr_6_6=>GND0, q_arr_6_5=>GND0, q_arr_6_4=>GND0, q_arr_6_3=>GND0, 
      q_arr_6_2=>GND0, q_arr_6_1=>GND0, q_arr_6_0=>GND0, q_arr_7_31=>GND0, 
      q_arr_7_30=>GND0, q_arr_7_29=>GND0, q_arr_7_28=>GND0, q_arr_7_27=>GND0, 
      q_arr_7_26=>GND0, q_arr_7_25=>GND0, q_arr_7_24=>GND0, q_arr_7_23=>GND0, 
      q_arr_7_22=>GND0, q_arr_7_21=>GND0, q_arr_7_20=>GND0, q_arr_7_19=>GND0, 
      q_arr_7_18=>GND0, q_arr_7_17=>GND0, q_arr_7_16=>GND0, q_arr_7_15=>GND0, 
      q_arr_7_14=>GND0, q_arr_7_13=>GND0, q_arr_7_12=>GND0, q_arr_7_11=>GND0, 
      q_arr_7_10=>GND0, q_arr_7_9=>GND0, q_arr_7_8=>GND0, q_arr_7_7=>GND0, 
      q_arr_7_6=>GND0, q_arr_7_5=>GND0, q_arr_7_4=>GND0, q_arr_7_3=>GND0, 
      q_arr_7_2=>GND0, q_arr_7_1=>GND0, q_arr_7_0=>GND0, q_arr_8_31=>GND0, 
      q_arr_8_30=>GND0, q_arr_8_29=>GND0, q_arr_8_28=>GND0, q_arr_8_27=>GND0, 
      q_arr_8_26=>GND0, q_arr_8_25=>GND0, q_arr_8_24=>GND0, q_arr_8_23=>GND0, 
      q_arr_8_22=>GND0, q_arr_8_21=>GND0, q_arr_8_20=>GND0, q_arr_8_19=>GND0, 
      q_arr_8_18=>GND0, q_arr_8_17=>GND0, q_arr_8_16=>GND0, q_arr_8_15=>GND0, 
      q_arr_8_14=>GND0, q_arr_8_13=>GND0, q_arr_8_12=>GND0, q_arr_8_11=>GND0, 
      q_arr_8_10=>GND0, q_arr_8_9=>GND0, q_arr_8_8=>GND0, q_arr_8_7=>GND0, 
      q_arr_8_6=>GND0, q_arr_8_5=>GND0, q_arr_8_4=>GND0, q_arr_8_3=>GND0, 
      q_arr_8_2=>GND0, q_arr_8_1=>GND0, q_arr_8_0=>GND0, q_arr_9_31=>GND0, 
      q_arr_9_30=>GND0, q_arr_9_29=>GND0, q_arr_9_28=>GND0, q_arr_9_27=>GND0, 
      q_arr_9_26=>GND0, q_arr_9_25=>GND0, q_arr_9_24=>GND0, q_arr_9_23=>GND0, 
      q_arr_9_22=>GND0, q_arr_9_21=>GND0, q_arr_9_20=>GND0, q_arr_9_19=>GND0, 
      q_arr_9_18=>GND0, q_arr_9_17=>GND0, q_arr_9_16=>GND0, q_arr_9_15=>GND0, 
      q_arr_9_14=>GND0, q_arr_9_13=>GND0, q_arr_9_12=>GND0, q_arr_9_11=>GND0, 
      q_arr_9_10=>GND0, q_arr_9_9=>GND0, q_arr_9_8=>GND0, q_arr_9_7=>GND0, 
      q_arr_9_6=>GND0, q_arr_9_5=>GND0, q_arr_9_4=>GND0, q_arr_9_3=>GND0, 
      q_arr_9_2=>GND0, q_arr_9_1=>GND0, q_arr_9_0=>GND0, q_arr_10_31=>GND0, 
      q_arr_10_30=>GND0, q_arr_10_29=>GND0, q_arr_10_28=>GND0, q_arr_10_27=>
      GND0, q_arr_10_26=>GND0, q_arr_10_25=>GND0, q_arr_10_24=>GND0, 
      q_arr_10_23=>GND0, q_arr_10_22=>GND0, q_arr_10_21=>GND0, q_arr_10_20=>
      GND0, q_arr_10_19=>GND0, q_arr_10_18=>GND0, q_arr_10_17=>GND0, 
      q_arr_10_16=>GND0, q_arr_10_15=>GND0, q_arr_10_14=>GND0, q_arr_10_13=>
      GND0, q_arr_10_12=>GND0, q_arr_10_11=>GND0, q_arr_10_10=>GND0, 
      q_arr_10_9=>GND0, q_arr_10_8=>GND0, q_arr_10_7=>GND0, q_arr_10_6=>GND0, 
      q_arr_10_5=>GND0, q_arr_10_4=>GND0, q_arr_10_3=>GND0, q_arr_10_2=>GND0, 
      q_arr_10_1=>GND0, q_arr_10_0=>GND0, q_arr_11_31=>GND0, q_arr_11_30=>
      GND0, q_arr_11_29=>GND0, q_arr_11_28=>GND0, q_arr_11_27=>GND0, 
      q_arr_11_26=>GND0, q_arr_11_25=>GND0, q_arr_11_24=>GND0, q_arr_11_23=>
      GND0, q_arr_11_22=>GND0, q_arr_11_21=>GND0, q_arr_11_20=>GND0, 
      q_arr_11_19=>GND0, q_arr_11_18=>GND0, q_arr_11_17=>GND0, q_arr_11_16=>
      GND0, q_arr_11_15=>GND0, q_arr_11_14=>GND0, q_arr_11_13=>GND0, 
      q_arr_11_12=>GND0, q_arr_11_11=>GND0, q_arr_11_10=>GND0, q_arr_11_9=>
      GND0, q_arr_11_8=>GND0, q_arr_11_7=>GND0, q_arr_11_6=>GND0, q_arr_11_5
      =>GND0, q_arr_11_4=>GND0, q_arr_11_3=>GND0, q_arr_11_2=>GND0, 
      q_arr_11_1=>GND0, q_arr_11_0=>GND0, q_arr_12_31=>GND0, q_arr_12_30=>
      GND0, q_arr_12_29=>GND0, q_arr_12_28=>GND0, q_arr_12_27=>GND0, 
      q_arr_12_26=>GND0, q_arr_12_25=>GND0, q_arr_12_24=>GND0, q_arr_12_23=>
      GND0, q_arr_12_22=>GND0, q_arr_12_21=>GND0, q_arr_12_20=>GND0, 
      q_arr_12_19=>GND0, q_arr_12_18=>GND0, q_arr_12_17=>GND0, q_arr_12_16=>
      GND0, q_arr_12_15=>GND0, q_arr_12_14=>GND0, q_arr_12_13=>GND0, 
      q_arr_12_12=>GND0, q_arr_12_11=>GND0, q_arr_12_10=>GND0, q_arr_12_9=>
      GND0, q_arr_12_8=>GND0, q_arr_12_7=>GND0, q_arr_12_6=>GND0, q_arr_12_5
      =>GND0, q_arr_12_4=>GND0, q_arr_12_3=>GND0, q_arr_12_2=>GND0, 
      q_arr_12_1=>GND0, q_arr_12_0=>GND0, q_arr_13_31=>GND0, q_arr_13_30=>
      GND0, q_arr_13_29=>GND0, q_arr_13_28=>GND0, q_arr_13_27=>GND0, 
      q_arr_13_26=>GND0, q_arr_13_25=>GND0, q_arr_13_24=>GND0, q_arr_13_23=>
      GND0, q_arr_13_22=>GND0, q_arr_13_21=>GND0, q_arr_13_20=>GND0, 
      q_arr_13_19=>GND0, q_arr_13_18=>GND0, q_arr_13_17=>GND0, q_arr_13_16=>
      GND0, q_arr_13_15=>GND0, q_arr_13_14=>GND0, q_arr_13_13=>GND0, 
      q_arr_13_12=>GND0, q_arr_13_11=>GND0, q_arr_13_10=>GND0, q_arr_13_9=>
      GND0, q_arr_13_8=>GND0, q_arr_13_7=>GND0, q_arr_13_6=>GND0, q_arr_13_5
      =>GND0, q_arr_13_4=>GND0, q_arr_13_3=>GND0, q_arr_13_2=>GND0, 
      q_arr_13_1=>GND0, q_arr_13_0=>GND0, q_arr_14_31=>GND0, q_arr_14_30=>
      GND0, q_arr_14_29=>GND0, q_arr_14_28=>GND0, q_arr_14_27=>GND0, 
      q_arr_14_26=>GND0, q_arr_14_25=>GND0, q_arr_14_24=>GND0, q_arr_14_23=>
      GND0, q_arr_14_22=>GND0, q_arr_14_21=>GND0, q_arr_14_20=>GND0, 
      q_arr_14_19=>GND0, q_arr_14_18=>GND0, q_arr_14_17=>GND0, q_arr_14_16=>
      GND0, q_arr_14_15=>GND0, q_arr_14_14=>GND0, q_arr_14_13=>GND0, 
      q_arr_14_12=>GND0, q_arr_14_11=>GND0, q_arr_14_10=>GND0, q_arr_14_9=>
      GND0, q_arr_14_8=>GND0, q_arr_14_7=>GND0, q_arr_14_6=>GND0, q_arr_14_5
      =>GND0, q_arr_14_4=>GND0, q_arr_14_3=>GND0, q_arr_14_2=>GND0, 
      q_arr_14_1=>GND0, q_arr_14_0=>GND0, q_arr_15_31=>GND0, q_arr_15_30=>
      GND0, q_arr_15_29=>GND0, q_arr_15_28=>GND0, q_arr_15_27=>GND0, 
      q_arr_15_26=>GND0, q_arr_15_25=>GND0, q_arr_15_24=>GND0, q_arr_15_23=>
      GND0, q_arr_15_22=>GND0, q_arr_15_21=>GND0, q_arr_15_20=>GND0, 
      q_arr_15_19=>GND0, q_arr_15_18=>GND0, q_arr_15_17=>GND0, q_arr_15_16=>
      GND0, q_arr_15_15=>GND0, q_arr_15_14=>GND0, q_arr_15_13=>GND0, 
      q_arr_15_12=>GND0, q_arr_15_11=>GND0, q_arr_15_10=>GND0, q_arr_15_9=>
      GND0, q_arr_15_8=>GND0, q_arr_15_7=>GND0, q_arr_15_6=>GND0, q_arr_15_5
      =>GND0, q_arr_15_4=>GND0, q_arr_15_3=>GND0, q_arr_15_2=>GND0, 
      q_arr_15_1=>GND0, q_arr_15_0=>GND0, q_arr_16_31=>GND0, q_arr_16_30=>
      GND0, q_arr_16_29=>GND0, q_arr_16_28=>GND0, q_arr_16_27=>GND0, 
      q_arr_16_26=>GND0, q_arr_16_25=>GND0, q_arr_16_24=>GND0, q_arr_16_23=>
      GND0, q_arr_16_22=>GND0, q_arr_16_21=>GND0, q_arr_16_20=>GND0, 
      q_arr_16_19=>GND0, q_arr_16_18=>GND0, q_arr_16_17=>GND0, q_arr_16_16=>
      GND0, q_arr_16_15=>GND0, q_arr_16_14=>GND0, q_arr_16_13=>GND0, 
      q_arr_16_12=>GND0, q_arr_16_11=>GND0, q_arr_16_10=>GND0, q_arr_16_9=>
      GND0, q_arr_16_8=>GND0, q_arr_16_7=>GND0, q_arr_16_6=>GND0, q_arr_16_5
      =>GND0, q_arr_16_4=>GND0, q_arr_16_3=>GND0, q_arr_16_2=>GND0, 
      q_arr_16_1=>GND0, q_arr_16_0=>GND0, q_arr_17_31=>GND0, q_arr_17_30=>
      GND0, q_arr_17_29=>GND0, q_arr_17_28=>GND0, q_arr_17_27=>GND0, 
      q_arr_17_26=>GND0, q_arr_17_25=>GND0, q_arr_17_24=>GND0, q_arr_17_23=>
      GND0, q_arr_17_22=>GND0, q_arr_17_21=>GND0, q_arr_17_20=>GND0, 
      q_arr_17_19=>GND0, q_arr_17_18=>GND0, q_arr_17_17=>GND0, q_arr_17_16=>
      GND0, q_arr_17_15=>GND0, q_arr_17_14=>GND0, q_arr_17_13=>GND0, 
      q_arr_17_12=>GND0, q_arr_17_11=>GND0, q_arr_17_10=>GND0, q_arr_17_9=>
      GND0, q_arr_17_8=>GND0, q_arr_17_7=>GND0, q_arr_17_6=>GND0, q_arr_17_5
      =>GND0, q_arr_17_4=>GND0, q_arr_17_3=>GND0, q_arr_17_2=>GND0, 
      q_arr_17_1=>GND0, q_arr_17_0=>GND0, q_arr_18_31=>GND0, q_arr_18_30=>
      GND0, q_arr_18_29=>GND0, q_arr_18_28=>GND0, q_arr_18_27=>GND0, 
      q_arr_18_26=>GND0, q_arr_18_25=>GND0, q_arr_18_24=>GND0, q_arr_18_23=>
      GND0, q_arr_18_22=>GND0, q_arr_18_21=>GND0, q_arr_18_20=>GND0, 
      q_arr_18_19=>GND0, q_arr_18_18=>GND0, q_arr_18_17=>GND0, q_arr_18_16=>
      GND0, q_arr_18_15=>GND0, q_arr_18_14=>GND0, q_arr_18_13=>GND0, 
      q_arr_18_12=>GND0, q_arr_18_11=>GND0, q_arr_18_10=>GND0, q_arr_18_9=>
      GND0, q_arr_18_8=>GND0, q_arr_18_7=>GND0, q_arr_18_6=>GND0, q_arr_18_5
      =>GND0, q_arr_18_4=>GND0, q_arr_18_3=>GND0, q_arr_18_2=>GND0, 
      q_arr_18_1=>GND0, q_arr_18_0=>GND0, q_arr_19_31=>GND0, q_arr_19_30=>
      GND0, q_arr_19_29=>GND0, q_arr_19_28=>GND0, q_arr_19_27=>GND0, 
      q_arr_19_26=>GND0, q_arr_19_25=>GND0, q_arr_19_24=>GND0, q_arr_19_23=>
      GND0, q_arr_19_22=>GND0, q_arr_19_21=>GND0, q_arr_19_20=>GND0, 
      q_arr_19_19=>GND0, q_arr_19_18=>GND0, q_arr_19_17=>GND0, q_arr_19_16=>
      GND0, q_arr_19_15=>GND0, q_arr_19_14=>GND0, q_arr_19_13=>GND0, 
      q_arr_19_12=>GND0, q_arr_19_11=>GND0, q_arr_19_10=>GND0, q_arr_19_9=>
      GND0, q_arr_19_8=>GND0, q_arr_19_7=>GND0, q_arr_19_6=>GND0, q_arr_19_5
      =>GND0, q_arr_19_4=>GND0, q_arr_19_3=>GND0, q_arr_19_2=>GND0, 
      q_arr_19_1=>GND0, q_arr_19_0=>GND0, q_arr_20_31=>GND0, q_arr_20_30=>
      GND0, q_arr_20_29=>GND0, q_arr_20_28=>GND0, q_arr_20_27=>GND0, 
      q_arr_20_26=>GND0, q_arr_20_25=>GND0, q_arr_20_24=>GND0, q_arr_20_23=>
      GND0, q_arr_20_22=>GND0, q_arr_20_21=>GND0, q_arr_20_20=>GND0, 
      q_arr_20_19=>GND0, q_arr_20_18=>GND0, q_arr_20_17=>GND0, q_arr_20_16=>
      GND0, q_arr_20_15=>GND0, q_arr_20_14=>GND0, q_arr_20_13=>GND0, 
      q_arr_20_12=>GND0, q_arr_20_11=>GND0, q_arr_20_10=>GND0, q_arr_20_9=>
      GND0, q_arr_20_8=>GND0, q_arr_20_7=>GND0, q_arr_20_6=>GND0, q_arr_20_5
      =>GND0, q_arr_20_4=>GND0, q_arr_20_3=>GND0, q_arr_20_2=>GND0, 
      q_arr_20_1=>GND0, q_arr_20_0=>GND0, q_arr_21_31=>GND0, q_arr_21_30=>
      GND0, q_arr_21_29=>GND0, q_arr_21_28=>GND0, q_arr_21_27=>GND0, 
      q_arr_21_26=>GND0, q_arr_21_25=>GND0, q_arr_21_24=>GND0, q_arr_21_23=>
      GND0, q_arr_21_22=>GND0, q_arr_21_21=>GND0, q_arr_21_20=>GND0, 
      q_arr_21_19=>GND0, q_arr_21_18=>GND0, q_arr_21_17=>GND0, q_arr_21_16=>
      GND0, q_arr_21_15=>GND0, q_arr_21_14=>GND0, q_arr_21_13=>GND0, 
      q_arr_21_12=>GND0, q_arr_21_11=>GND0, q_arr_21_10=>GND0, q_arr_21_9=>
      GND0, q_arr_21_8=>GND0, q_arr_21_7=>GND0, q_arr_21_6=>GND0, q_arr_21_5
      =>GND0, q_arr_21_4=>GND0, q_arr_21_3=>GND0, q_arr_21_2=>GND0, 
      q_arr_21_1=>GND0, q_arr_21_0=>GND0, q_arr_22_31=>GND0, q_arr_22_30=>
      GND0, q_arr_22_29=>GND0, q_arr_22_28=>GND0, q_arr_22_27=>GND0, 
      q_arr_22_26=>GND0, q_arr_22_25=>GND0, q_arr_22_24=>GND0, q_arr_22_23=>
      GND0, q_arr_22_22=>GND0, q_arr_22_21=>GND0, q_arr_22_20=>GND0, 
      q_arr_22_19=>GND0, q_arr_22_18=>GND0, q_arr_22_17=>GND0, q_arr_22_16=>
      GND0, q_arr_22_15=>GND0, q_arr_22_14=>GND0, q_arr_22_13=>GND0, 
      q_arr_22_12=>GND0, q_arr_22_11=>GND0, q_arr_22_10=>GND0, q_arr_22_9=>
      GND0, q_arr_22_8=>GND0, q_arr_22_7=>GND0, q_arr_22_6=>GND0, q_arr_22_5
      =>GND0, q_arr_22_4=>GND0, q_arr_22_3=>GND0, q_arr_22_2=>GND0, 
      q_arr_22_1=>GND0, q_arr_22_0=>GND0, q_arr_23_31=>GND0, q_arr_23_30=>
      GND0, q_arr_23_29=>GND0, q_arr_23_28=>GND0, q_arr_23_27=>GND0, 
      q_arr_23_26=>GND0, q_arr_23_25=>GND0, q_arr_23_24=>GND0, q_arr_23_23=>
      GND0, q_arr_23_22=>GND0, q_arr_23_21=>GND0, q_arr_23_20=>GND0, 
      q_arr_23_19=>GND0, q_arr_23_18=>GND0, q_arr_23_17=>GND0, q_arr_23_16=>
      GND0, q_arr_23_15=>GND0, q_arr_23_14=>GND0, q_arr_23_13=>GND0, 
      q_arr_23_12=>GND0, q_arr_23_11=>GND0, q_arr_23_10=>GND0, q_arr_23_9=>
      GND0, q_arr_23_8=>GND0, q_arr_23_7=>GND0, q_arr_23_6=>GND0, q_arr_23_5
      =>GND0, q_arr_23_4=>GND0, q_arr_23_3=>GND0, q_arr_23_2=>GND0, 
      q_arr_23_1=>GND0, q_arr_23_0=>GND0, q_arr_24_31=>GND0, q_arr_24_30=>
      GND0, q_arr_24_29=>GND0, q_arr_24_28=>GND0, q_arr_24_27=>GND0, 
      q_arr_24_26=>GND0, q_arr_24_25=>GND0, q_arr_24_24=>GND0, q_arr_24_23=>
      GND0, q_arr_24_22=>GND0, q_arr_24_21=>GND0, q_arr_24_20=>GND0, 
      q_arr_24_19=>GND0, q_arr_24_18=>GND0, q_arr_24_17=>GND0, q_arr_24_16=>
      GND0, q_arr_24_15=>GND0, q_arr_24_14=>GND0, q_arr_24_13=>GND0, 
      q_arr_24_12=>GND0, q_arr_24_11=>GND0, q_arr_24_10=>GND0, q_arr_24_9=>
      GND0, q_arr_24_8=>GND0, q_arr_24_7=>GND0, q_arr_24_6=>GND0, q_arr_24_5
      =>GND0, q_arr_24_4=>GND0, q_arr_24_3=>GND0, q_arr_24_2=>GND0, 
      q_arr_24_1=>GND0, q_arr_24_0=>GND0);
   mul_layer_gen_multipliers_gen_0_mul_gen_mul_gen : ModifiedBoothMultiplier
       port map ( M(15)=>img_data_0_15, M(14)=>nx19396, M(13)=>img_data_0_13, 
      M(12)=>img_data_0_12, M(11)=>img_data_0_11, M(10)=>img_data_0_10, M(9)
      =>img_data_0_9, M(8)=>img_data_0_8, M(7)=>img_data_0_7, M(6)=>
      img_data_0_6, M(5)=>img_data_0_5, M(4)=>img_data_0_4, M(3)=>
      img_data_0_3, M(2)=>img_data_0_2, M(1)=>img_data_0_1, M(0)=>
      img_data_0_0, R(15)=>filter_data_0_15, R(14)=>filter_data_0_14, R(13)
      =>filter_data_0_13, R(12)=>filter_data_0_12, R(11)=>filter_data_0_11, 
      R(10)=>filter_data_0_10, R(9)=>filter_data_0_9, R(8)=>filter_data_0_8, 
      R(7)=>filter_data_0_7, R(6)=>filter_data_0_6, R(5)=>filter_data_0_5, 
      R(4)=>filter_data_0_4, R(3)=>filter_data_0_3, R(2)=>filter_data_0_2, 
      R(1)=>filter_data_0_1, R(0)=>filter_data_0_0, cnt_enable=>nx16627, 
      product(31)=>d_arr_mul_0_31, product(30)=>d_arr_mul_0_30, product(29)
      =>d_arr_mul_0_29, product(28)=>d_arr_mul_0_28, product(27)=>
      d_arr_mul_0_27, product(26)=>d_arr_mul_0_26, product(25)=>
      d_arr_mul_0_25, product(24)=>d_arr_mul_0_24, product(23)=>
      d_arr_mul_0_23, product(22)=>d_arr_mul_0_22, product(21)=>
      d_arr_mul_0_21, product(20)=>d_arr_mul_0_20, product(19)=>
      d_arr_mul_0_19, product(18)=>d_arr_mul_0_18, product(17)=>
      d_arr_mul_0_17, product(16)=>d_arr_mul_0_16, product(15)=>
      d_arr_mul_0_15, product(14)=>d_arr_mul_0_14, product(13)=>
      d_arr_mul_0_13, product(12)=>d_arr_mul_0_12, product(11)=>
      d_arr_mul_0_11, product(10)=>d_arr_mul_0_10, product(9)=>d_arr_mul_0_9, 
      product(8)=>d_arr_mul_0_8, product(7)=>d_arr_mul_0_7, product(6)=>
      d_arr_mul_0_6, product(5)=>d_arr_mul_0_5, product(4)=>d_arr_mul_0_4, 
      product(3)=>d_arr_mul_0_3, product(2)=>d_arr_mul_0_2, product(1)=>
      d_arr_mul_0_1, product(0)=>d_arr_mul_0_0, clk=>clk);
   mul_layer_gen_multipliers_gen_1_mul_gen_mul_gen : ModifiedBoothMultiplier
       port map ( M(15)=>img_data_1_15, M(14)=>nx19400, M(13)=>img_data_1_13, 
      M(12)=>img_data_1_12, M(11)=>img_data_1_11, M(10)=>nx19402, M(9)=>
      img_data_1_9, M(8)=>img_data_1_8, M(7)=>img_data_1_7, M(6)=>
      img_data_1_6, M(5)=>img_data_1_5, M(4)=>img_data_1_4, M(3)=>
      img_data_1_3, M(2)=>img_data_1_2, M(1)=>img_data_1_1, M(0)=>
      img_data_1_0, R(15)=>filter_data_1_15, R(14)=>filter_data_1_14, R(13)
      =>filter_data_1_13, R(12)=>filter_data_1_12, R(11)=>filter_data_1_11, 
      R(10)=>filter_data_1_10, R(9)=>filter_data_1_9, R(8)=>filter_data_1_8, 
      R(7)=>filter_data_1_7, R(6)=>filter_data_1_6, R(5)=>filter_data_1_5, 
      R(4)=>filter_data_1_4, R(3)=>filter_data_1_3, R(2)=>filter_data_1_2, 
      R(1)=>filter_data_1_1, R(0)=>filter_data_1_0, cnt_enable=>nx16473, 
      product(31)=>d_arr_mul_1_31, product(30)=>d_arr_mul_1_30, product(29)
      =>d_arr_mul_1_29, product(28)=>d_arr_mul_1_28, product(27)=>
      d_arr_mul_1_27, product(26)=>d_arr_mul_1_26, product(25)=>
      d_arr_mul_1_25, product(24)=>d_arr_mul_1_24, product(23)=>
      d_arr_mul_1_23, product(22)=>d_arr_mul_1_22, product(21)=>
      d_arr_mul_1_21, product(20)=>d_arr_mul_1_20, product(19)=>
      d_arr_mul_1_19, product(18)=>d_arr_mul_1_18, product(17)=>
      d_arr_mul_1_17, product(16)=>d_arr_mul_1_16, product(15)=>
      d_arr_mul_1_15, product(14)=>d_arr_mul_1_14, product(13)=>
      d_arr_mul_1_13, product(12)=>d_arr_mul_1_12, product(11)=>
      d_arr_mul_1_11, product(10)=>d_arr_mul_1_10, product(9)=>d_arr_mul_1_9, 
      product(8)=>d_arr_mul_1_8, product(7)=>d_arr_mul_1_7, product(6)=>
      d_arr_mul_1_6, product(5)=>d_arr_mul_1_5, product(4)=>d_arr_mul_1_4, 
      product(3)=>d_arr_mul_1_3, product(2)=>d_arr_mul_1_2, product(1)=>
      d_arr_mul_1_1, product(0)=>d_arr_mul_1_0, clk=>clk);
   mul_layer_gen_multipliers_gen_2_mul_gen_mul_gen : ModifiedBoothMultiplier
       port map ( M(15)=>img_data_2_15, M(14)=>nx19406, M(13)=>img_data_2_13, 
      M(12)=>img_data_2_12, M(11)=>img_data_2_11, M(10)=>nx19408, M(9)=>
      img_data_2_9, M(8)=>img_data_2_8, M(7)=>img_data_2_7, M(6)=>
      img_data_2_6, M(5)=>img_data_2_5, M(4)=>img_data_2_4, M(3)=>
      img_data_2_3, M(2)=>img_data_2_2, M(1)=>img_data_2_1, M(0)=>
      img_data_2_0, R(15)=>filter_data_2_15, R(14)=>filter_data_2_14, R(13)
      =>filter_data_2_13, R(12)=>filter_data_2_12, R(11)=>filter_data_2_11, 
      R(10)=>filter_data_2_10, R(9)=>filter_data_2_9, R(8)=>filter_data_2_8, 
      R(7)=>filter_data_2_7, R(6)=>filter_data_2_6, R(5)=>filter_data_2_5, 
      R(4)=>filter_data_2_4, R(3)=>filter_data_2_3, R(2)=>filter_data_2_2, 
      R(1)=>filter_data_2_1, R(0)=>filter_data_2_0, cnt_enable=>nx16473, 
      product(31)=>d_arr_mul_2_31, product(30)=>d_arr_mul_2_30, product(29)
      =>d_arr_mul_2_29, product(28)=>d_arr_mul_2_28, product(27)=>
      d_arr_mul_2_27, product(26)=>d_arr_mul_2_26, product(25)=>
      d_arr_mul_2_25, product(24)=>d_arr_mul_2_24, product(23)=>
      d_arr_mul_2_23, product(22)=>d_arr_mul_2_22, product(21)=>
      d_arr_mul_2_21, product(20)=>d_arr_mul_2_20, product(19)=>
      d_arr_mul_2_19, product(18)=>d_arr_mul_2_18, product(17)=>
      d_arr_mul_2_17, product(16)=>d_arr_mul_2_16, product(15)=>
      d_arr_mul_2_15, product(14)=>d_arr_mul_2_14, product(13)=>
      d_arr_mul_2_13, product(12)=>d_arr_mul_2_12, product(11)=>
      d_arr_mul_2_11, product(10)=>d_arr_mul_2_10, product(9)=>d_arr_mul_2_9, 
      product(8)=>d_arr_mul_2_8, product(7)=>d_arr_mul_2_7, product(6)=>
      d_arr_mul_2_6, product(5)=>d_arr_mul_2_5, product(4)=>d_arr_mul_2_4, 
      product(3)=>d_arr_mul_2_3, product(2)=>d_arr_mul_2_2, product(1)=>
      d_arr_mul_2_1, product(0)=>d_arr_mul_2_0, clk=>clk);
   mul_layer_gen_multipliers_gen_3_mul_gen_mul_gen : ModifiedBoothMultiplier
       port map ( M(15)=>img_data_5_15, M(14)=>nx19410, M(13)=>img_data_5_13, 
      M(12)=>img_data_5_12, M(11)=>img_data_5_11, M(10)=>img_data_5_10, M(9)
      =>img_data_5_9, M(8)=>img_data_5_8, M(7)=>img_data_5_7, M(6)=>
      img_data_5_6, M(5)=>img_data_5_5, M(4)=>img_data_5_4, M(3)=>
      img_data_5_3, M(2)=>img_data_5_2, M(1)=>img_data_5_1, M(0)=>
      img_data_5_0, R(15)=>ordered_filter_data_3_15, R(14)=>
      ordered_filter_data_3_14, R(13)=>ordered_filter_data_3_13, R(12)=>
      ordered_filter_data_3_12, R(11)=>ordered_filter_data_3_11, R(10)=>
      ordered_filter_data_3_10, R(9)=>ordered_filter_data_3_9, R(8)=>
      ordered_filter_data_3_8, R(7)=>ordered_filter_data_3_7, R(6)=>
      ordered_filter_data_3_6, R(5)=>ordered_filter_data_3_5, R(4)=>
      ordered_filter_data_3_4, R(3)=>ordered_filter_data_3_3, R(2)=>
      ordered_filter_data_3_2, R(1)=>ordered_filter_data_3_1, R(0)=>
      ordered_filter_data_3_0, cnt_enable=>nx16629, product(31)=>
      d_arr_mul_3_31, product(30)=>d_arr_mul_3_30, product(29)=>
      d_arr_mul_3_29, product(28)=>d_arr_mul_3_28, product(27)=>
      d_arr_mul_3_27, product(26)=>d_arr_mul_3_26, product(25)=>
      d_arr_mul_3_25, product(24)=>d_arr_mul_3_24, product(23)=>
      d_arr_mul_3_23, product(22)=>d_arr_mul_3_22, product(21)=>
      d_arr_mul_3_21, product(20)=>d_arr_mul_3_20, product(19)=>
      d_arr_mul_3_19, product(18)=>d_arr_mul_3_18, product(17)=>
      d_arr_mul_3_17, product(16)=>d_arr_mul_3_16, product(15)=>
      d_arr_mul_3_15, product(14)=>d_arr_mul_3_14, product(13)=>
      d_arr_mul_3_13, product(12)=>d_arr_mul_3_12, product(11)=>
      d_arr_mul_3_11, product(10)=>d_arr_mul_3_10, product(9)=>d_arr_mul_3_9, 
      product(8)=>d_arr_mul_3_8, product(7)=>d_arr_mul_3_7, product(6)=>
      d_arr_mul_3_6, product(5)=>d_arr_mul_3_5, product(4)=>d_arr_mul_3_4, 
      product(3)=>d_arr_mul_3_3, product(2)=>d_arr_mul_3_2, product(1)=>
      d_arr_mul_3_1, product(0)=>d_arr_mul_3_0, clk=>clk);
   mul_layer_gen_multipliers_gen_4_mul_gen_mul_gen : ModifiedBoothMultiplier
       port map ( M(15)=>img_data_6_15, M(14)=>nx19414, M(13)=>img_data_6_13, 
      M(12)=>img_data_6_12, M(11)=>img_data_6_11, M(10)=>nx19416, M(9)=>
      img_data_6_9, M(8)=>img_data_6_8, M(7)=>img_data_6_7, M(6)=>
      img_data_6_6, M(5)=>img_data_6_5, M(4)=>img_data_6_4, M(3)=>
      img_data_6_3, M(2)=>img_data_6_2, M(1)=>img_data_6_1, M(0)=>
      img_data_6_0, R(15)=>ordered_filter_data_4_15, R(14)=>
      ordered_filter_data_4_14, R(13)=>ordered_filter_data_4_13, R(12)=>
      ordered_filter_data_4_12, R(11)=>ordered_filter_data_4_11, R(10)=>
      ordered_filter_data_4_10, R(9)=>ordered_filter_data_4_9, R(8)=>
      ordered_filter_data_4_8, R(7)=>ordered_filter_data_4_7, R(6)=>
      ordered_filter_data_4_6, R(5)=>ordered_filter_data_4_5, R(4)=>
      ordered_filter_data_4_4, R(3)=>ordered_filter_data_4_3, R(2)=>
      ordered_filter_data_4_2, R(1)=>ordered_filter_data_4_1, R(0)=>
      ordered_filter_data_4_0, cnt_enable=>nx16629, product(31)=>
      d_arr_mul_4_31, product(30)=>d_arr_mul_4_30, product(29)=>
      d_arr_mul_4_29, product(28)=>d_arr_mul_4_28, product(27)=>
      d_arr_mul_4_27, product(26)=>d_arr_mul_4_26, product(25)=>
      d_arr_mul_4_25, product(24)=>d_arr_mul_4_24, product(23)=>
      d_arr_mul_4_23, product(22)=>d_arr_mul_4_22, product(21)=>
      d_arr_mul_4_21, product(20)=>d_arr_mul_4_20, product(19)=>
      d_arr_mul_4_19, product(18)=>d_arr_mul_4_18, product(17)=>
      d_arr_mul_4_17, product(16)=>d_arr_mul_4_16, product(15)=>
      d_arr_mul_4_15, product(14)=>d_arr_mul_4_14, product(13)=>
      d_arr_mul_4_13, product(12)=>d_arr_mul_4_12, product(11)=>
      d_arr_mul_4_11, product(10)=>d_arr_mul_4_10, product(9)=>d_arr_mul_4_9, 
      product(8)=>d_arr_mul_4_8, product(7)=>d_arr_mul_4_7, product(6)=>
      d_arr_mul_4_6, product(5)=>d_arr_mul_4_5, product(4)=>d_arr_mul_4_4, 
      product(3)=>d_arr_mul_4_3, product(2)=>d_arr_mul_4_2, product(1)=>
      d_arr_mul_4_1, product(0)=>d_arr_mul_4_0, clk=>clk);
   mul_layer_gen_multipliers_gen_5_mul_gen_mul_gen : ModifiedBoothMultiplier
       port map ( M(15)=>nx16659, M(14)=>nx19420, M(13)=>img_data_7_13, 
      M(12)=>img_data_7_12, M(11)=>img_data_7_11, M(10)=>nx19422, M(9)=>
      img_data_7_9, M(8)=>img_data_7_8, M(7)=>img_data_7_7, M(6)=>
      img_data_7_6, M(5)=>img_data_7_5, M(4)=>img_data_7_4, M(3)=>
      img_data_7_3, M(2)=>img_data_7_2, M(1)=>img_data_7_1, M(0)=>
      img_data_7_0, R(15)=>ordered_filter_data_5_15, R(14)=>
      ordered_filter_data_5_14, R(13)=>ordered_filter_data_5_13, R(12)=>
      ordered_filter_data_5_12, R(11)=>ordered_filter_data_5_11, R(10)=>
      ordered_filter_data_5_10, R(9)=>ordered_filter_data_5_9, R(8)=>
      ordered_filter_data_5_8, R(7)=>ordered_filter_data_5_7, R(6)=>
      ordered_filter_data_5_6, R(5)=>ordered_filter_data_5_5, R(4)=>
      ordered_filter_data_5_4, R(3)=>ordered_filter_data_5_3, R(2)=>
      ordered_filter_data_5_2, R(1)=>ordered_filter_data_5_1, R(0)=>
      ordered_filter_data_5_0, cnt_enable=>nx16631, product(31)=>
      d_arr_mul_5_31, product(30)=>d_arr_mul_5_30, product(29)=>
      d_arr_mul_5_29, product(28)=>d_arr_mul_5_28, product(27)=>
      d_arr_mul_5_27, product(26)=>d_arr_mul_5_26, product(25)=>
      d_arr_mul_5_25, product(24)=>d_arr_mul_5_24, product(23)=>
      d_arr_mul_5_23, product(22)=>d_arr_mul_5_22, product(21)=>
      d_arr_mul_5_21, product(20)=>d_arr_mul_5_20, product(19)=>
      d_arr_mul_5_19, product(18)=>d_arr_mul_5_18, product(17)=>
      d_arr_mul_5_17, product(16)=>d_arr_mul_5_16, product(15)=>
      d_arr_mul_5_15, product(14)=>d_arr_mul_5_14, product(13)=>
      d_arr_mul_5_13, product(12)=>d_arr_mul_5_12, product(11)=>
      d_arr_mul_5_11, product(10)=>d_arr_mul_5_10, product(9)=>d_arr_mul_5_9, 
      product(8)=>d_arr_mul_5_8, product(7)=>d_arr_mul_5_7, product(6)=>
      d_arr_mul_5_6, product(5)=>d_arr_mul_5_5, product(4)=>d_arr_mul_5_4, 
      product(3)=>d_arr_mul_5_3, product(2)=>d_arr_mul_5_2, product(1)=>
      d_arr_mul_5_1, product(0)=>d_arr_mul_5_0, clk=>clk);
   mul_layer_gen_multipliers_gen_6_mul_gen_mul_gen : ModifiedBoothMultiplier
       port map ( M(15)=>img_data_10_15, M(14)=>nx19424, M(13)=>
      img_data_10_13, M(12)=>img_data_10_12, M(11)=>img_data_10_11, M(10)=>
      img_data_10_10, M(9)=>img_data_10_9, M(8)=>img_data_10_8, M(7)=>
      img_data_10_7, M(6)=>img_data_10_6, M(5)=>img_data_10_5, M(4)=>
      img_data_10_4, M(3)=>img_data_10_3, M(2)=>img_data_10_2, M(1)=>
      img_data_10_1, M(0)=>img_data_10_0, R(15)=>ordered_filter_data_6_15, 
      R(14)=>ordered_filter_data_6_14, R(13)=>ordered_filter_data_6_13, 
      R(12)=>ordered_filter_data_6_12, R(11)=>ordered_filter_data_6_11, 
      R(10)=>ordered_filter_data_6_10, R(9)=>ordered_filter_data_6_9, R(8)=>
      ordered_filter_data_6_8, R(7)=>ordered_filter_data_6_7, R(6)=>
      ordered_filter_data_6_6, R(5)=>ordered_filter_data_6_5, R(4)=>
      ordered_filter_data_6_4, R(3)=>ordered_filter_data_6_3, R(2)=>
      ordered_filter_data_6_2, R(1)=>ordered_filter_data_6_1, R(0)=>
      ordered_filter_data_6_0, cnt_enable=>nx16631, product(31)=>
      d_arr_mul_6_31, product(30)=>d_arr_mul_6_30, product(29)=>
      d_arr_mul_6_29, product(28)=>d_arr_mul_6_28, product(27)=>
      d_arr_mul_6_27, product(26)=>d_arr_mul_6_26, product(25)=>
      d_arr_mul_6_25, product(24)=>d_arr_mul_6_24, product(23)=>
      d_arr_mul_6_23, product(22)=>d_arr_mul_6_22, product(21)=>
      d_arr_mul_6_21, product(20)=>d_arr_mul_6_20, product(19)=>
      d_arr_mul_6_19, product(18)=>d_arr_mul_6_18, product(17)=>
      d_arr_mul_6_17, product(16)=>d_arr_mul_6_16, product(15)=>
      d_arr_mul_6_15, product(14)=>d_arr_mul_6_14, product(13)=>
      d_arr_mul_6_13, product(12)=>d_arr_mul_6_12, product(11)=>
      d_arr_mul_6_11, product(10)=>d_arr_mul_6_10, product(9)=>d_arr_mul_6_9, 
      product(8)=>d_arr_mul_6_8, product(7)=>d_arr_mul_6_7, product(6)=>
      d_arr_mul_6_6, product(5)=>d_arr_mul_6_5, product(4)=>d_arr_mul_6_4, 
      product(3)=>d_arr_mul_6_3, product(2)=>d_arr_mul_6_2, product(1)=>
      d_arr_mul_6_1, product(0)=>d_arr_mul_6_0, clk=>clk);
   mul_layer_gen_multipliers_gen_7_mul_gen_mul_gen : ModifiedBoothMultiplier
       port map ( M(15)=>nx16661, M(14)=>nx19428, M(13)=>img_data_11_13, 
      M(12)=>img_data_11_12, M(11)=>img_data_11_11, M(10)=>nx19430, M(9)=>
      img_data_11_9, M(8)=>img_data_11_8, M(7)=>img_data_11_7, M(6)=>
      img_data_11_6, M(5)=>img_data_11_5, M(4)=>img_data_11_4, M(3)=>
      img_data_11_3, M(2)=>img_data_11_2, M(1)=>img_data_11_1, M(0)=>
      img_data_11_0, R(15)=>ordered_filter_data_7_15, R(14)=>
      ordered_filter_data_7_14, R(13)=>ordered_filter_data_7_13, R(12)=>
      ordered_filter_data_7_12, R(11)=>ordered_filter_data_7_11, R(10)=>
      ordered_filter_data_7_10, R(9)=>ordered_filter_data_7_9, R(8)=>
      ordered_filter_data_7_8, R(7)=>ordered_filter_data_7_7, R(6)=>
      ordered_filter_data_7_6, R(5)=>ordered_filter_data_7_5, R(4)=>
      ordered_filter_data_7_4, R(3)=>ordered_filter_data_7_3, R(2)=>
      ordered_filter_data_7_2, R(1)=>ordered_filter_data_7_1, R(0)=>
      ordered_filter_data_7_0, cnt_enable=>nx16633, product(31)=>
      d_arr_mul_7_31, product(30)=>d_arr_mul_7_30, product(29)=>
      d_arr_mul_7_29, product(28)=>d_arr_mul_7_28, product(27)=>
      d_arr_mul_7_27, product(26)=>d_arr_mul_7_26, product(25)=>
      d_arr_mul_7_25, product(24)=>d_arr_mul_7_24, product(23)=>
      d_arr_mul_7_23, product(22)=>d_arr_mul_7_22, product(21)=>
      d_arr_mul_7_21, product(20)=>d_arr_mul_7_20, product(19)=>
      d_arr_mul_7_19, product(18)=>d_arr_mul_7_18, product(17)=>
      d_arr_mul_7_17, product(16)=>d_arr_mul_7_16, product(15)=>
      d_arr_mul_7_15, product(14)=>d_arr_mul_7_14, product(13)=>
      d_arr_mul_7_13, product(12)=>d_arr_mul_7_12, product(11)=>
      d_arr_mul_7_11, product(10)=>d_arr_mul_7_10, product(9)=>d_arr_mul_7_9, 
      product(8)=>d_arr_mul_7_8, product(7)=>d_arr_mul_7_7, product(6)=>
      d_arr_mul_7_6, product(5)=>d_arr_mul_7_5, product(4)=>d_arr_mul_7_4, 
      product(3)=>d_arr_mul_7_3, product(2)=>d_arr_mul_7_2, product(1)=>
      d_arr_mul_7_1, product(0)=>d_arr_mul_7_0, clk=>clk);
   mul_layer_gen_multipliers_gen_8_mul_gen_mul_gen : ModifiedBoothMultiplier
       port map ( M(15)=>nx16663, M(14)=>nx19434, M(13)=>img_data_12_13, 
      M(12)=>img_data_12_12, M(11)=>img_data_12_11, M(10)=>nx19436, M(9)=>
      img_data_12_9, M(8)=>img_data_12_8, M(7)=>img_data_12_7, M(6)=>
      img_data_12_6, M(5)=>img_data_12_5, M(4)=>img_data_12_4, M(3)=>
      img_data_12_3, M(2)=>img_data_12_2, M(1)=>img_data_12_1, M(0)=>
      img_data_12_0, R(15)=>ordered_filter_data_8_15, R(14)=>
      ordered_filter_data_8_14, R(13)=>ordered_filter_data_8_13, R(12)=>
      ordered_filter_data_8_12, R(11)=>ordered_filter_data_8_11, R(10)=>
      ordered_filter_data_8_10, R(9)=>ordered_filter_data_8_9, R(8)=>
      ordered_filter_data_8_8, R(7)=>ordered_filter_data_8_7, R(6)=>
      ordered_filter_data_8_6, R(5)=>ordered_filter_data_8_5, R(4)=>
      ordered_filter_data_8_4, R(3)=>ordered_filter_data_8_3, R(2)=>
      ordered_filter_data_8_2, R(1)=>ordered_filter_data_8_1, R(0)=>
      ordered_filter_data_8_0, cnt_enable=>nx16633, product(31)=>
      d_arr_mul_8_31, product(30)=>d_arr_mul_8_30, product(29)=>
      d_arr_mul_8_29, product(28)=>d_arr_mul_8_28, product(27)=>
      d_arr_mul_8_27, product(26)=>d_arr_mul_8_26, product(25)=>
      d_arr_mul_8_25, product(24)=>d_arr_mul_8_24, product(23)=>
      d_arr_mul_8_23, product(22)=>d_arr_mul_8_22, product(21)=>
      d_arr_mul_8_21, product(20)=>d_arr_mul_8_20, product(19)=>
      d_arr_mul_8_19, product(18)=>d_arr_mul_8_18, product(17)=>
      d_arr_mul_8_17, product(16)=>d_arr_mul_8_16, product(15)=>
      d_arr_mul_8_15, product(14)=>d_arr_mul_8_14, product(13)=>
      d_arr_mul_8_13, product(12)=>d_arr_mul_8_12, product(11)=>
      d_arr_mul_8_11, product(10)=>d_arr_mul_8_10, product(9)=>d_arr_mul_8_9, 
      product(8)=>d_arr_mul_8_8, product(7)=>d_arr_mul_8_7, product(6)=>
      d_arr_mul_8_6, product(5)=>d_arr_mul_8_5, product(4)=>d_arr_mul_8_4, 
      product(3)=>d_arr_mul_8_3, product(2)=>d_arr_mul_8_2, product(1)=>
      d_arr_mul_8_1, product(0)=>d_arr_mul_8_0, clk=>clk);
   mul_layer_gen_multipliers_gen_9_mul_gen_mul_gen : ModifiedBoothMultiplier
       port map ( M(15)=>nx16405, M(14)=>ordered_img_data_9_14, M(13)=>
      ordered_img_data_9_13, M(12)=>ordered_img_data_9_12, M(11)=>
      ordered_img_data_9_11, M(10)=>ordered_img_data_9_10, M(9)=>
      ordered_img_data_9_9, M(8)=>ordered_img_data_9_8, M(7)=>
      ordered_img_data_9_7, M(6)=>ordered_img_data_9_6, M(5)=>
      ordered_img_data_9_5, M(4)=>ordered_img_data_9_4, M(3)=>
      ordered_img_data_9_3, M(2)=>ordered_img_data_9_2, M(1)=>
      ordered_img_data_9_1, M(0)=>ordered_img_data_9_0, R(15)=>
      ordered_filter_data_9_15, R(14)=>ordered_filter_data_9_14, R(13)=>
      ordered_filter_data_9_13, R(12)=>ordered_filter_data_9_12, R(11)=>
      ordered_filter_data_9_11, R(10)=>ordered_filter_data_9_10, R(9)=>
      ordered_filter_data_9_9, R(8)=>ordered_filter_data_9_8, R(7)=>
      ordered_filter_data_9_7, R(6)=>ordered_filter_data_9_6, R(5)=>
      ordered_filter_data_9_5, R(4)=>ordered_filter_data_9_4, R(3)=>
      ordered_filter_data_9_3, R(2)=>ordered_filter_data_9_2, R(1)=>
      ordered_filter_data_9_1, R(0)=>ordered_filter_data_9_0, cnt_enable=>
      nx16475, product(31)=>d_arr_mul_9_31, product(30)=>d_arr_mul_9_30, 
      product(29)=>d_arr_mul_9_29, product(28)=>d_arr_mul_9_28, product(27)
      =>d_arr_mul_9_27, product(26)=>d_arr_mul_9_26, product(25)=>
      d_arr_mul_9_25, product(24)=>d_arr_mul_9_24, product(23)=>
      d_arr_mul_9_23, product(22)=>d_arr_mul_9_22, product(21)=>
      d_arr_mul_9_21, product(20)=>d_arr_mul_9_20, product(19)=>
      d_arr_mul_9_19, product(18)=>d_arr_mul_9_18, product(17)=>
      d_arr_mul_9_17, product(16)=>d_arr_mul_9_16, product(15)=>
      d_arr_mul_9_15, product(14)=>d_arr_mul_9_14, product(13)=>
      d_arr_mul_9_13, product(12)=>d_arr_mul_9_12, product(11)=>
      d_arr_mul_9_11, product(10)=>d_arr_mul_9_10, product(9)=>d_arr_mul_9_9, 
      product(8)=>d_arr_mul_9_8, product(7)=>d_arr_mul_9_7, product(6)=>
      d_arr_mul_9_6, product(5)=>d_arr_mul_9_5, product(4)=>d_arr_mul_9_4, 
      product(3)=>d_arr_mul_9_3, product(2)=>d_arr_mul_9_2, product(1)=>
      d_arr_mul_9_1, product(0)=>d_arr_mul_9_0, clk=>clk);
   mul_layer_gen_multipliers_gen_10_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>nx16413, M(14)=>
      ordered_img_data_10_14, M(13)=>ordered_img_data_10_13, M(12)=>
      ordered_img_data_10_12, M(11)=>ordered_img_data_10_11, M(10)=>
      ordered_img_data_10_10, M(9)=>ordered_img_data_10_9, M(8)=>
      ordered_img_data_10_8, M(7)=>ordered_img_data_10_7, M(6)=>
      ordered_img_data_10_6, M(5)=>ordered_img_data_10_5, M(4)=>
      ordered_img_data_10_4, M(3)=>ordered_img_data_10_3, M(2)=>
      ordered_img_data_10_2, M(1)=>ordered_img_data_10_1, M(0)=>
      ordered_img_data_10_0, R(15)=>ordered_filter_data_10_15, R(14)=>
      ordered_filter_data_10_14, R(13)=>ordered_filter_data_10_13, R(12)=>
      ordered_filter_data_10_12, R(11)=>ordered_filter_data_10_11, R(10)=>
      ordered_filter_data_10_10, R(9)=>ordered_filter_data_10_9, R(8)=>
      ordered_filter_data_10_8, R(7)=>ordered_filter_data_10_7, R(6)=>
      ordered_filter_data_10_6, R(5)=>ordered_filter_data_10_5, R(4)=>
      ordered_filter_data_10_4, R(3)=>ordered_filter_data_10_3, R(2)=>
      ordered_filter_data_10_2, R(1)=>ordered_filter_data_10_1, R(0)=>
      ordered_filter_data_10_0, cnt_enable=>nx16635, product(31)=>
      d_arr_mul_10_31, product(30)=>d_arr_mul_10_30, product(29)=>
      d_arr_mul_10_29, product(28)=>d_arr_mul_10_28, product(27)=>
      d_arr_mul_10_27, product(26)=>d_arr_mul_10_26, product(25)=>
      d_arr_mul_10_25, product(24)=>d_arr_mul_10_24, product(23)=>
      d_arr_mul_10_23, product(22)=>d_arr_mul_10_22, product(21)=>
      d_arr_mul_10_21, product(20)=>d_arr_mul_10_20, product(19)=>
      d_arr_mul_10_19, product(18)=>d_arr_mul_10_18, product(17)=>
      d_arr_mul_10_17, product(16)=>d_arr_mul_10_16, product(15)=>
      d_arr_mul_10_15, product(14)=>d_arr_mul_10_14, product(13)=>
      d_arr_mul_10_13, product(12)=>d_arr_mul_10_12, product(11)=>
      d_arr_mul_10_11, product(10)=>d_arr_mul_10_10, product(9)=>
      d_arr_mul_10_9, product(8)=>d_arr_mul_10_8, product(7)=>d_arr_mul_10_7, 
      product(6)=>d_arr_mul_10_6, product(5)=>d_arr_mul_10_5, product(4)=>
      d_arr_mul_10_4, product(3)=>d_arr_mul_10_3, product(2)=>d_arr_mul_10_2, 
      product(1)=>d_arr_mul_10_1, product(0)=>d_arr_mul_10_0, clk=>clk);
   mul_layer_gen_multipliers_gen_11_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>nx16421, M(14)=>
      ordered_img_data_11_14, M(13)=>ordered_img_data_11_13, M(12)=>
      ordered_img_data_11_12, M(11)=>ordered_img_data_11_11, M(10)=>
      ordered_img_data_11_10, M(9)=>ordered_img_data_11_9, M(8)=>
      ordered_img_data_11_8, M(7)=>ordered_img_data_11_7, M(6)=>
      ordered_img_data_11_6, M(5)=>ordered_img_data_11_5, M(4)=>
      ordered_img_data_11_4, M(3)=>ordered_img_data_11_3, M(2)=>
      ordered_img_data_11_2, M(1)=>ordered_img_data_11_1, M(0)=>
      ordered_img_data_11_0, R(15)=>ordered_filter_data_11_15, R(14)=>
      ordered_filter_data_11_14, R(13)=>ordered_filter_data_11_13, R(12)=>
      ordered_filter_data_11_12, R(11)=>ordered_filter_data_11_11, R(10)=>
      ordered_filter_data_11_10, R(9)=>ordered_filter_data_11_9, R(8)=>
      ordered_filter_data_11_8, R(7)=>ordered_filter_data_11_7, R(6)=>
      ordered_filter_data_11_6, R(5)=>ordered_filter_data_11_5, R(4)=>
      ordered_filter_data_11_4, R(3)=>ordered_filter_data_11_3, R(2)=>
      ordered_filter_data_11_2, R(1)=>ordered_filter_data_11_1, R(0)=>
      ordered_filter_data_11_0, cnt_enable=>nx16635, product(31)=>
      d_arr_mul_11_31, product(30)=>d_arr_mul_11_30, product(29)=>
      d_arr_mul_11_29, product(28)=>d_arr_mul_11_28, product(27)=>
      d_arr_mul_11_27, product(26)=>d_arr_mul_11_26, product(25)=>
      d_arr_mul_11_25, product(24)=>d_arr_mul_11_24, product(23)=>
      d_arr_mul_11_23, product(22)=>d_arr_mul_11_22, product(21)=>
      d_arr_mul_11_21, product(20)=>d_arr_mul_11_20, product(19)=>
      d_arr_mul_11_19, product(18)=>d_arr_mul_11_18, product(17)=>
      d_arr_mul_11_17, product(16)=>d_arr_mul_11_16, product(15)=>
      d_arr_mul_11_15, product(14)=>d_arr_mul_11_14, product(13)=>
      d_arr_mul_11_13, product(12)=>d_arr_mul_11_12, product(11)=>
      d_arr_mul_11_11, product(10)=>d_arr_mul_11_10, product(9)=>
      d_arr_mul_11_9, product(8)=>d_arr_mul_11_8, product(7)=>d_arr_mul_11_7, 
      product(6)=>d_arr_mul_11_6, product(5)=>d_arr_mul_11_5, product(4)=>
      d_arr_mul_11_4, product(3)=>d_arr_mul_11_3, product(2)=>d_arr_mul_11_2, 
      product(1)=>d_arr_mul_11_1, product(0)=>d_arr_mul_11_0, clk=>clk);
   mul_layer_gen_multipliers_gen_12_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>nx16429, M(14)=>
      ordered_img_data_12_14, M(13)=>ordered_img_data_12_13, M(12)=>
      ordered_img_data_12_12, M(11)=>ordered_img_data_12_11, M(10)=>
      ordered_img_data_12_10, M(9)=>ordered_img_data_12_9, M(8)=>
      ordered_img_data_12_8, M(7)=>ordered_img_data_12_7, M(6)=>
      ordered_img_data_12_6, M(5)=>ordered_img_data_12_5, M(4)=>
      ordered_img_data_12_4, M(3)=>ordered_img_data_12_3, M(2)=>
      ordered_img_data_12_2, M(1)=>ordered_img_data_12_1, M(0)=>
      ordered_img_data_12_0, R(15)=>ordered_filter_data_12_15, R(14)=>
      ordered_filter_data_12_14, R(13)=>ordered_filter_data_12_13, R(12)=>
      ordered_filter_data_12_12, R(11)=>ordered_filter_data_12_11, R(10)=>
      ordered_filter_data_12_10, R(9)=>ordered_filter_data_12_9, R(8)=>
      ordered_filter_data_12_8, R(7)=>ordered_filter_data_12_7, R(6)=>
      ordered_filter_data_12_6, R(5)=>ordered_filter_data_12_5, R(4)=>
      ordered_filter_data_12_4, R(3)=>ordered_filter_data_12_3, R(2)=>
      ordered_filter_data_12_2, R(1)=>ordered_filter_data_12_1, R(0)=>
      ordered_filter_data_12_0, cnt_enable=>nx16637, product(31)=>
      d_arr_mul_12_31, product(30)=>d_arr_mul_12_30, product(29)=>
      d_arr_mul_12_29, product(28)=>d_arr_mul_12_28, product(27)=>
      d_arr_mul_12_27, product(26)=>d_arr_mul_12_26, product(25)=>
      d_arr_mul_12_25, product(24)=>d_arr_mul_12_24, product(23)=>
      d_arr_mul_12_23, product(22)=>d_arr_mul_12_22, product(21)=>
      d_arr_mul_12_21, product(20)=>d_arr_mul_12_20, product(19)=>
      d_arr_mul_12_19, product(18)=>d_arr_mul_12_18, product(17)=>
      d_arr_mul_12_17, product(16)=>d_arr_mul_12_16, product(15)=>
      d_arr_mul_12_15, product(14)=>d_arr_mul_12_14, product(13)=>
      d_arr_mul_12_13, product(12)=>d_arr_mul_12_12, product(11)=>
      d_arr_mul_12_11, product(10)=>d_arr_mul_12_10, product(9)=>
      d_arr_mul_12_9, product(8)=>d_arr_mul_12_8, product(7)=>d_arr_mul_12_7, 
      product(6)=>d_arr_mul_12_6, product(5)=>d_arr_mul_12_5, product(4)=>
      d_arr_mul_12_4, product(3)=>d_arr_mul_12_3, product(2)=>d_arr_mul_12_2, 
      product(1)=>d_arr_mul_12_1, product(0)=>d_arr_mul_12_0, clk=>clk);
   mul_layer_gen_multipliers_gen_13_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>nx16437, M(14)=>
      ordered_img_data_13_14, M(13)=>ordered_img_data_13_13, M(12)=>
      ordered_img_data_13_12, M(11)=>ordered_img_data_13_11, M(10)=>
      ordered_img_data_13_10, M(9)=>ordered_img_data_13_9, M(8)=>
      ordered_img_data_13_8, M(7)=>ordered_img_data_13_7, M(6)=>
      ordered_img_data_13_6, M(5)=>ordered_img_data_13_5, M(4)=>
      ordered_img_data_13_4, M(3)=>ordered_img_data_13_3, M(2)=>
      ordered_img_data_13_2, M(1)=>ordered_img_data_13_1, M(0)=>
      ordered_img_data_13_0, R(15)=>ordered_filter_data_13_15, R(14)=>
      ordered_filter_data_13_14, R(13)=>ordered_filter_data_13_13, R(12)=>
      ordered_filter_data_13_12, R(11)=>ordered_filter_data_13_11, R(10)=>
      ordered_filter_data_13_10, R(9)=>ordered_filter_data_13_9, R(8)=>
      ordered_filter_data_13_8, R(7)=>ordered_filter_data_13_7, R(6)=>
      ordered_filter_data_13_6, R(5)=>ordered_filter_data_13_5, R(4)=>
      ordered_filter_data_13_4, R(3)=>ordered_filter_data_13_3, R(2)=>
      ordered_filter_data_13_2, R(1)=>ordered_filter_data_13_1, R(0)=>
      ordered_filter_data_13_0, cnt_enable=>nx16637, product(31)=>
      d_arr_mul_13_31, product(30)=>d_arr_mul_13_30, product(29)=>
      d_arr_mul_13_29, product(28)=>d_arr_mul_13_28, product(27)=>
      d_arr_mul_13_27, product(26)=>d_arr_mul_13_26, product(25)=>
      d_arr_mul_13_25, product(24)=>d_arr_mul_13_24, product(23)=>
      d_arr_mul_13_23, product(22)=>d_arr_mul_13_22, product(21)=>
      d_arr_mul_13_21, product(20)=>d_arr_mul_13_20, product(19)=>
      d_arr_mul_13_19, product(18)=>d_arr_mul_13_18, product(17)=>
      d_arr_mul_13_17, product(16)=>d_arr_mul_13_16, product(15)=>
      d_arr_mul_13_15, product(14)=>d_arr_mul_13_14, product(13)=>
      d_arr_mul_13_13, product(12)=>d_arr_mul_13_12, product(11)=>
      d_arr_mul_13_11, product(10)=>d_arr_mul_13_10, product(9)=>
      d_arr_mul_13_9, product(8)=>d_arr_mul_13_8, product(7)=>d_arr_mul_13_7, 
      product(6)=>d_arr_mul_13_6, product(5)=>d_arr_mul_13_5, product(4)=>
      d_arr_mul_13_4, product(3)=>d_arr_mul_13_3, product(2)=>d_arr_mul_13_2, 
      product(1)=>d_arr_mul_13_1, product(0)=>d_arr_mul_13_0, clk=>clk);
   mul_layer_gen_multipliers_gen_14_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>nx16445, M(14)=>
      ordered_img_data_14_14, M(13)=>ordered_img_data_14_13, M(12)=>
      ordered_img_data_14_12, M(11)=>ordered_img_data_14_11, M(10)=>
      ordered_img_data_14_10, M(9)=>ordered_img_data_14_9, M(8)=>
      ordered_img_data_14_8, M(7)=>ordered_img_data_14_7, M(6)=>
      ordered_img_data_14_6, M(5)=>ordered_img_data_14_5, M(4)=>
      ordered_img_data_14_4, M(3)=>ordered_img_data_14_3, M(2)=>
      ordered_img_data_14_2, M(1)=>ordered_img_data_14_1, M(0)=>
      ordered_img_data_14_0, R(15)=>ordered_filter_data_14_15, R(14)=>
      ordered_filter_data_14_14, R(13)=>ordered_filter_data_14_13, R(12)=>
      ordered_filter_data_14_12, R(11)=>ordered_filter_data_14_11, R(10)=>
      ordered_filter_data_14_10, R(9)=>ordered_filter_data_14_9, R(8)=>
      ordered_filter_data_14_8, R(7)=>ordered_filter_data_14_7, R(6)=>
      ordered_filter_data_14_6, R(5)=>ordered_filter_data_14_5, R(4)=>
      ordered_filter_data_14_4, R(3)=>ordered_filter_data_14_3, R(2)=>
      ordered_filter_data_14_2, R(1)=>ordered_filter_data_14_1, R(0)=>
      ordered_filter_data_14_0, cnt_enable=>nx16639, product(31)=>
      d_arr_mul_14_31, product(30)=>d_arr_mul_14_30, product(29)=>
      d_arr_mul_14_29, product(28)=>d_arr_mul_14_28, product(27)=>
      d_arr_mul_14_27, product(26)=>d_arr_mul_14_26, product(25)=>
      d_arr_mul_14_25, product(24)=>d_arr_mul_14_24, product(23)=>
      d_arr_mul_14_23, product(22)=>d_arr_mul_14_22, product(21)=>
      d_arr_mul_14_21, product(20)=>d_arr_mul_14_20, product(19)=>
      d_arr_mul_14_19, product(18)=>d_arr_mul_14_18, product(17)=>
      d_arr_mul_14_17, product(16)=>d_arr_mul_14_16, product(15)=>
      d_arr_mul_14_15, product(14)=>d_arr_mul_14_14, product(13)=>
      d_arr_mul_14_13, product(12)=>d_arr_mul_14_12, product(11)=>
      d_arr_mul_14_11, product(10)=>d_arr_mul_14_10, product(9)=>
      d_arr_mul_14_9, product(8)=>d_arr_mul_14_8, product(7)=>d_arr_mul_14_7, 
      product(6)=>d_arr_mul_14_6, product(5)=>d_arr_mul_14_5, product(4)=>
      d_arr_mul_14_4, product(3)=>d_arr_mul_14_3, product(2)=>d_arr_mul_14_2, 
      product(1)=>d_arr_mul_14_1, product(0)=>d_arr_mul_14_0, clk=>clk);
   mul_layer_gen_multipliers_gen_15_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>nx16453, M(14)=>
      ordered_img_data_15_14, M(13)=>ordered_img_data_15_13, M(12)=>
      ordered_img_data_15_12, M(11)=>ordered_img_data_15_11, M(10)=>
      ordered_img_data_15_10, M(9)=>ordered_img_data_15_9, M(8)=>
      ordered_img_data_15_8, M(7)=>ordered_img_data_15_7, M(6)=>
      ordered_img_data_15_6, M(5)=>ordered_img_data_15_5, M(4)=>
      ordered_img_data_15_4, M(3)=>ordered_img_data_15_3, M(2)=>
      ordered_img_data_15_2, M(1)=>ordered_img_data_15_1, M(0)=>
      ordered_img_data_15_0, R(15)=>ordered_filter_data_15_15, R(14)=>
      ordered_filter_data_15_14, R(13)=>ordered_filter_data_15_13, R(12)=>
      ordered_filter_data_15_12, R(11)=>ordered_filter_data_15_11, R(10)=>
      ordered_filter_data_15_10, R(9)=>ordered_filter_data_15_9, R(8)=>
      ordered_filter_data_15_8, R(7)=>ordered_filter_data_15_7, R(6)=>
      ordered_filter_data_15_6, R(5)=>ordered_filter_data_15_5, R(4)=>
      ordered_filter_data_15_4, R(3)=>ordered_filter_data_15_3, R(2)=>
      ordered_filter_data_15_2, R(1)=>ordered_filter_data_15_1, R(0)=>
      ordered_filter_data_15_0, cnt_enable=>nx16639, product(31)=>
      d_arr_mul_15_31, product(30)=>d_arr_mul_15_30, product(29)=>
      d_arr_mul_15_29, product(28)=>d_arr_mul_15_28, product(27)=>
      d_arr_mul_15_27, product(26)=>d_arr_mul_15_26, product(25)=>
      d_arr_mul_15_25, product(24)=>d_arr_mul_15_24, product(23)=>
      d_arr_mul_15_23, product(22)=>d_arr_mul_15_22, product(21)=>
      d_arr_mul_15_21, product(20)=>d_arr_mul_15_20, product(19)=>
      d_arr_mul_15_19, product(18)=>d_arr_mul_15_18, product(17)=>
      d_arr_mul_15_17, product(16)=>d_arr_mul_15_16, product(15)=>
      d_arr_mul_15_15, product(14)=>d_arr_mul_15_14, product(13)=>
      d_arr_mul_15_13, product(12)=>d_arr_mul_15_12, product(11)=>
      d_arr_mul_15_11, product(10)=>d_arr_mul_15_10, product(9)=>
      d_arr_mul_15_9, product(8)=>d_arr_mul_15_8, product(7)=>d_arr_mul_15_7, 
      product(6)=>d_arr_mul_15_6, product(5)=>d_arr_mul_15_5, product(4)=>
      d_arr_mul_15_4, product(3)=>d_arr_mul_15_3, product(2)=>d_arr_mul_15_2, 
      product(1)=>d_arr_mul_15_1, product(0)=>d_arr_mul_15_0, clk=>clk);
   mul_layer_gen_multipliers_gen_16_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>nx16461, M(14)=>
      ordered_img_data_16_14, M(13)=>ordered_img_data_16_13, M(12)=>
      ordered_img_data_16_12, M(11)=>ordered_img_data_16_11, M(10)=>
      ordered_img_data_16_10, M(9)=>ordered_img_data_16_9, M(8)=>
      ordered_img_data_16_8, M(7)=>ordered_img_data_16_7, M(6)=>
      ordered_img_data_16_6, M(5)=>ordered_img_data_16_5, M(4)=>
      ordered_img_data_16_4, M(3)=>ordered_img_data_16_3, M(2)=>
      ordered_img_data_16_2, M(1)=>ordered_img_data_16_1, M(0)=>
      ordered_img_data_16_0, R(15)=>ordered_filter_data_16_15, R(14)=>
      ordered_filter_data_16_14, R(13)=>ordered_filter_data_16_13, R(12)=>
      ordered_filter_data_16_12, R(11)=>ordered_filter_data_16_11, R(10)=>
      ordered_filter_data_16_10, R(9)=>ordered_filter_data_16_9, R(8)=>
      ordered_filter_data_16_8, R(7)=>ordered_filter_data_16_7, R(6)=>
      ordered_filter_data_16_6, R(5)=>ordered_filter_data_16_5, R(4)=>
      ordered_filter_data_16_4, R(3)=>ordered_filter_data_16_3, R(2)=>
      ordered_filter_data_16_2, R(1)=>ordered_filter_data_16_1, R(0)=>
      ordered_filter_data_16_0, cnt_enable=>nx16477, product(31)=>
      d_arr_mul_16_31, product(30)=>d_arr_mul_16_30, product(29)=>
      d_arr_mul_16_29, product(28)=>d_arr_mul_16_28, product(27)=>
      d_arr_mul_16_27, product(26)=>d_arr_mul_16_26, product(25)=>
      d_arr_mul_16_25, product(24)=>d_arr_mul_16_24, product(23)=>
      d_arr_mul_16_23, product(22)=>d_arr_mul_16_22, product(21)=>
      d_arr_mul_16_21, product(20)=>d_arr_mul_16_20, product(19)=>
      d_arr_mul_16_19, product(18)=>d_arr_mul_16_18, product(17)=>
      d_arr_mul_16_17, product(16)=>d_arr_mul_16_16, product(15)=>
      d_arr_mul_16_15, product(14)=>d_arr_mul_16_14, product(13)=>
      d_arr_mul_16_13, product(12)=>d_arr_mul_16_12, product(11)=>
      d_arr_mul_16_11, product(10)=>d_arr_mul_16_10, product(9)=>
      d_arr_mul_16_9, product(8)=>d_arr_mul_16_8, product(7)=>d_arr_mul_16_7, 
      product(6)=>d_arr_mul_16_6, product(5)=>d_arr_mul_16_5, product(4)=>
      d_arr_mul_16_4, product(3)=>d_arr_mul_16_3, product(2)=>d_arr_mul_16_2, 
      product(1)=>d_arr_mul_16_1, product(0)=>d_arr_mul_16_0, clk=>clk);
   mul_layer_gen_multipliers_gen_17_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>nx16469, M(14)=>
      ordered_img_data_17_14, M(13)=>ordered_img_data_17_13, M(12)=>
      ordered_img_data_17_12, M(11)=>ordered_img_data_17_11, M(10)=>
      ordered_img_data_17_10, M(9)=>ordered_img_data_17_9, M(8)=>
      ordered_img_data_17_8, M(7)=>ordered_img_data_17_7, M(6)=>
      ordered_img_data_17_6, M(5)=>ordered_img_data_17_5, M(4)=>
      ordered_img_data_17_4, M(3)=>ordered_img_data_17_3, M(2)=>
      ordered_img_data_17_2, M(1)=>ordered_img_data_17_1, M(0)=>
      ordered_img_data_17_0, R(15)=>ordered_filter_data_17_15, R(14)=>
      ordered_filter_data_17_14, R(13)=>ordered_filter_data_17_13, R(12)=>
      ordered_filter_data_17_12, R(11)=>ordered_filter_data_17_11, R(10)=>
      ordered_filter_data_17_10, R(9)=>ordered_filter_data_17_9, R(8)=>
      ordered_filter_data_17_8, R(7)=>ordered_filter_data_17_7, R(6)=>
      ordered_filter_data_17_6, R(5)=>ordered_filter_data_17_5, R(4)=>
      ordered_filter_data_17_4, R(3)=>ordered_filter_data_17_3, R(2)=>
      ordered_filter_data_17_2, R(1)=>ordered_filter_data_17_1, R(0)=>
      ordered_filter_data_17_0, cnt_enable=>nx16641, product(31)=>
      d_arr_mul_17_31, product(30)=>d_arr_mul_17_30, product(29)=>
      d_arr_mul_17_29, product(28)=>d_arr_mul_17_28, product(27)=>
      d_arr_mul_17_27, product(26)=>d_arr_mul_17_26, product(25)=>
      d_arr_mul_17_25, product(24)=>d_arr_mul_17_24, product(23)=>
      d_arr_mul_17_23, product(22)=>d_arr_mul_17_22, product(21)=>
      d_arr_mul_17_21, product(20)=>d_arr_mul_17_20, product(19)=>
      d_arr_mul_17_19, product(18)=>d_arr_mul_17_18, product(17)=>
      d_arr_mul_17_17, product(16)=>d_arr_mul_17_16, product(15)=>
      d_arr_mul_17_15, product(14)=>d_arr_mul_17_14, product(13)=>
      d_arr_mul_17_13, product(12)=>d_arr_mul_17_12, product(11)=>
      d_arr_mul_17_11, product(10)=>d_arr_mul_17_10, product(9)=>
      d_arr_mul_17_9, product(8)=>d_arr_mul_17_8, product(7)=>d_arr_mul_17_7, 
      product(6)=>d_arr_mul_17_6, product(5)=>d_arr_mul_17_5, product(4)=>
      d_arr_mul_17_4, product(3)=>d_arr_mul_17_3, product(2)=>d_arr_mul_17_2, 
      product(1)=>d_arr_mul_17_1, product(0)=>d_arr_mul_17_0, clk=>clk);
   mul_layer_gen_multipliers_gen_18_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>img_data_18_15, M(14)=>
      nx19438, M(13)=>img_data_18_13, M(12)=>img_data_18_12, M(11)=>
      img_data_18_11, M(10)=>img_data_18_10, M(9)=>img_data_18_9, M(8)=>
      img_data_18_8, M(7)=>img_data_18_7, M(6)=>img_data_18_6, M(5)=>
      img_data_18_5, M(4)=>img_data_18_4, M(3)=>img_data_18_3, M(2)=>
      img_data_18_2, M(1)=>img_data_18_1, M(0)=>img_data_18_0, R(15)=>
      filter_data_18_15, R(14)=>filter_data_18_14, R(13)=>filter_data_18_13, 
      R(12)=>filter_data_18_12, R(11)=>filter_data_18_11, R(10)=>
      filter_data_18_10, R(9)=>filter_data_18_9, R(8)=>filter_data_18_8, 
      R(7)=>filter_data_18_7, R(6)=>filter_data_18_6, R(5)=>filter_data_18_5, 
      R(4)=>filter_data_18_4, R(3)=>filter_data_18_3, R(2)=>filter_data_18_2, 
      R(1)=>filter_data_18_1, R(0)=>filter_data_18_0, cnt_enable=>nx16641, 
      product(31)=>d_arr_mul_18_31, product(30)=>d_arr_mul_18_30, 
      product(29)=>d_arr_mul_18_29, product(28)=>d_arr_mul_18_28, 
      product(27)=>d_arr_mul_18_27, product(26)=>d_arr_mul_18_26, 
      product(25)=>d_arr_mul_18_25, product(24)=>d_arr_mul_18_24, 
      product(23)=>d_arr_mul_18_23, product(22)=>d_arr_mul_18_22, 
      product(21)=>d_arr_mul_18_21, product(20)=>d_arr_mul_18_20, 
      product(19)=>d_arr_mul_18_19, product(18)=>d_arr_mul_18_18, 
      product(17)=>d_arr_mul_18_17, product(16)=>d_arr_mul_18_16, 
      product(15)=>d_arr_mul_18_15, product(14)=>d_arr_mul_18_14, 
      product(13)=>d_arr_mul_18_13, product(12)=>d_arr_mul_18_12, 
      product(11)=>d_arr_mul_18_11, product(10)=>d_arr_mul_18_10, product(9)
      =>d_arr_mul_18_9, product(8)=>d_arr_mul_18_8, product(7)=>
      d_arr_mul_18_7, product(6)=>d_arr_mul_18_6, product(5)=>d_arr_mul_18_5, 
      product(4)=>d_arr_mul_18_4, product(3)=>d_arr_mul_18_3, product(2)=>
      d_arr_mul_18_2, product(1)=>d_arr_mul_18_1, product(0)=>d_arr_mul_18_0, 
      clk=>clk);
   mul_layer_gen_multipliers_gen_19_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>img_data_19_15, M(14)=>
      img_data_19_14, M(13)=>img_data_19_13, M(12)=>img_data_19_12, M(11)=>
      img_data_19_11, M(10)=>img_data_19_10, M(9)=>img_data_19_9, M(8)=>
      img_data_19_8, M(7)=>img_data_19_7, M(6)=>img_data_19_6, M(5)=>
      img_data_19_5, M(4)=>img_data_19_4, M(3)=>img_data_19_3, M(2)=>
      img_data_19_2, M(1)=>img_data_19_1, M(0)=>img_data_19_0, R(15)=>
      filter_data_19_15, R(14)=>filter_data_19_14, R(13)=>filter_data_19_13, 
      R(12)=>filter_data_19_12, R(11)=>filter_data_19_11, R(10)=>
      filter_data_19_10, R(9)=>filter_data_19_9, R(8)=>filter_data_19_8, 
      R(7)=>filter_data_19_7, R(6)=>filter_data_19_6, R(5)=>filter_data_19_5, 
      R(4)=>filter_data_19_4, R(3)=>filter_data_19_3, R(2)=>filter_data_19_2, 
      R(1)=>filter_data_19_1, R(0)=>filter_data_19_0, cnt_enable=>nx16643, 
      product(31)=>d_arr_mul_19_31, product(30)=>d_arr_mul_19_30, 
      product(29)=>d_arr_mul_19_29, product(28)=>d_arr_mul_19_28, 
      product(27)=>d_arr_mul_19_27, product(26)=>d_arr_mul_19_26, 
      product(25)=>d_arr_mul_19_25, product(24)=>d_arr_mul_19_24, 
      product(23)=>d_arr_mul_19_23, product(22)=>d_arr_mul_19_22, 
      product(21)=>d_arr_mul_19_21, product(20)=>d_arr_mul_19_20, 
      product(19)=>d_arr_mul_19_19, product(18)=>d_arr_mul_19_18, 
      product(17)=>d_arr_mul_19_17, product(16)=>d_arr_mul_19_16, 
      product(15)=>d_arr_mul_19_15, product(14)=>d_arr_mul_19_14, 
      product(13)=>d_arr_mul_19_13, product(12)=>d_arr_mul_19_12, 
      product(11)=>d_arr_mul_19_11, product(10)=>d_arr_mul_19_10, product(9)
      =>d_arr_mul_19_9, product(8)=>d_arr_mul_19_8, product(7)=>
      d_arr_mul_19_7, product(6)=>d_arr_mul_19_6, product(5)=>d_arr_mul_19_5, 
      product(4)=>d_arr_mul_19_4, product(3)=>d_arr_mul_19_3, product(2)=>
      d_arr_mul_19_2, product(1)=>d_arr_mul_19_1, product(0)=>d_arr_mul_19_0, 
      clk=>clk);
   mul_layer_gen_multipliers_gen_20_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>img_data_20_15, M(14)=>
      nx19440, M(13)=>img_data_20_13, M(12)=>img_data_20_12, M(11)=>
      img_data_20_11, M(10)=>img_data_20_10, M(9)=>img_data_20_9, M(8)=>
      img_data_20_8, M(7)=>img_data_20_7, M(6)=>img_data_20_6, M(5)=>
      img_data_20_5, M(4)=>img_data_20_4, M(3)=>img_data_20_3, M(2)=>
      img_data_20_2, M(1)=>img_data_20_1, M(0)=>img_data_20_0, R(15)=>
      filter_data_20_15, R(14)=>filter_data_20_14, R(13)=>filter_data_20_13, 
      R(12)=>filter_data_20_12, R(11)=>filter_data_20_11, R(10)=>
      filter_data_20_10, R(9)=>filter_data_20_9, R(8)=>filter_data_20_8, 
      R(7)=>filter_data_20_7, R(6)=>filter_data_20_6, R(5)=>filter_data_20_5, 
      R(4)=>filter_data_20_4, R(3)=>filter_data_20_3, R(2)=>filter_data_20_2, 
      R(1)=>filter_data_20_1, R(0)=>filter_data_20_0, cnt_enable=>nx16643, 
      product(31)=>d_arr_mul_20_31, product(30)=>d_arr_mul_20_30, 
      product(29)=>d_arr_mul_20_29, product(28)=>d_arr_mul_20_28, 
      product(27)=>d_arr_mul_20_27, product(26)=>d_arr_mul_20_26, 
      product(25)=>d_arr_mul_20_25, product(24)=>d_arr_mul_20_24, 
      product(23)=>d_arr_mul_20_23, product(22)=>d_arr_mul_20_22, 
      product(21)=>d_arr_mul_20_21, product(20)=>d_arr_mul_20_20, 
      product(19)=>d_arr_mul_20_19, product(18)=>d_arr_mul_20_18, 
      product(17)=>d_arr_mul_20_17, product(16)=>d_arr_mul_20_16, 
      product(15)=>d_arr_mul_20_15, product(14)=>d_arr_mul_20_14, 
      product(13)=>d_arr_mul_20_13, product(12)=>d_arr_mul_20_12, 
      product(11)=>d_arr_mul_20_11, product(10)=>d_arr_mul_20_10, product(9)
      =>d_arr_mul_20_9, product(8)=>d_arr_mul_20_8, product(7)=>
      d_arr_mul_20_7, product(6)=>d_arr_mul_20_6, product(5)=>d_arr_mul_20_5, 
      product(4)=>d_arr_mul_20_4, product(3)=>d_arr_mul_20_3, product(2)=>
      d_arr_mul_20_2, product(1)=>d_arr_mul_20_1, product(0)=>d_arr_mul_20_0, 
      clk=>clk);
   mul_layer_gen_multipliers_gen_21_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>img_data_21_15, M(14)=>
      nx19442, M(13)=>img_data_21_13, M(12)=>img_data_21_12, M(11)=>
      img_data_21_11, M(10)=>img_data_21_10, M(9)=>img_data_21_9, M(8)=>
      img_data_21_8, M(7)=>img_data_21_7, M(6)=>img_data_21_6, M(5)=>
      img_data_21_5, M(4)=>img_data_21_4, M(3)=>img_data_21_3, M(2)=>
      img_data_21_2, M(1)=>img_data_21_1, M(0)=>img_data_21_0, R(15)=>
      filter_data_21_15, R(14)=>filter_data_21_14, R(13)=>filter_data_21_13, 
      R(12)=>filter_data_21_12, R(11)=>filter_data_21_11, R(10)=>
      filter_data_21_10, R(9)=>filter_data_21_9, R(8)=>filter_data_21_8, 
      R(7)=>filter_data_21_7, R(6)=>filter_data_21_6, R(5)=>filter_data_21_5, 
      R(4)=>filter_data_21_4, R(3)=>filter_data_21_3, R(2)=>filter_data_21_2, 
      R(1)=>filter_data_21_1, R(0)=>filter_data_21_0, cnt_enable=>nx16645, 
      product(31)=>d_arr_mul_21_31, product(30)=>d_arr_mul_21_30, 
      product(29)=>d_arr_mul_21_29, product(28)=>d_arr_mul_21_28, 
      product(27)=>d_arr_mul_21_27, product(26)=>d_arr_mul_21_26, 
      product(25)=>d_arr_mul_21_25, product(24)=>d_arr_mul_21_24, 
      product(23)=>d_arr_mul_21_23, product(22)=>d_arr_mul_21_22, 
      product(21)=>d_arr_mul_21_21, product(20)=>d_arr_mul_21_20, 
      product(19)=>d_arr_mul_21_19, product(18)=>d_arr_mul_21_18, 
      product(17)=>d_arr_mul_21_17, product(16)=>d_arr_mul_21_16, 
      product(15)=>d_arr_mul_21_15, product(14)=>d_arr_mul_21_14, 
      product(13)=>d_arr_mul_21_13, product(12)=>d_arr_mul_21_12, 
      product(11)=>d_arr_mul_21_11, product(10)=>d_arr_mul_21_10, product(9)
      =>d_arr_mul_21_9, product(8)=>d_arr_mul_21_8, product(7)=>
      d_arr_mul_21_7, product(6)=>d_arr_mul_21_6, product(5)=>d_arr_mul_21_5, 
      product(4)=>d_arr_mul_21_4, product(3)=>d_arr_mul_21_3, product(2)=>
      d_arr_mul_21_2, product(1)=>d_arr_mul_21_1, product(0)=>d_arr_mul_21_0, 
      clk=>clk);
   mul_layer_gen_multipliers_gen_22_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>img_data_22_15, M(14)=>
      nx19444, M(13)=>img_data_22_13, M(12)=>img_data_22_12, M(11)=>
      img_data_22_11, M(10)=>img_data_22_10, M(9)=>img_data_22_9, M(8)=>
      img_data_22_8, M(7)=>img_data_22_7, M(6)=>img_data_22_6, M(5)=>
      img_data_22_5, M(4)=>img_data_22_4, M(3)=>img_data_22_3, M(2)=>
      img_data_22_2, M(1)=>img_data_22_1, M(0)=>img_data_22_0, R(15)=>
      filter_data_22_15, R(14)=>filter_data_22_14, R(13)=>filter_data_22_13, 
      R(12)=>filter_data_22_12, R(11)=>filter_data_22_11, R(10)=>
      filter_data_22_10, R(9)=>filter_data_22_9, R(8)=>filter_data_22_8, 
      R(7)=>filter_data_22_7, R(6)=>filter_data_22_6, R(5)=>filter_data_22_5, 
      R(4)=>filter_data_22_4, R(3)=>filter_data_22_3, R(2)=>filter_data_22_2, 
      R(1)=>filter_data_22_1, R(0)=>filter_data_22_0, cnt_enable=>nx16645, 
      product(31)=>d_arr_mul_22_31, product(30)=>d_arr_mul_22_30, 
      product(29)=>d_arr_mul_22_29, product(28)=>d_arr_mul_22_28, 
      product(27)=>d_arr_mul_22_27, product(26)=>d_arr_mul_22_26, 
      product(25)=>d_arr_mul_22_25, product(24)=>d_arr_mul_22_24, 
      product(23)=>d_arr_mul_22_23, product(22)=>d_arr_mul_22_22, 
      product(21)=>d_arr_mul_22_21, product(20)=>d_arr_mul_22_20, 
      product(19)=>d_arr_mul_22_19, product(18)=>d_arr_mul_22_18, 
      product(17)=>d_arr_mul_22_17, product(16)=>d_arr_mul_22_16, 
      product(15)=>d_arr_mul_22_15, product(14)=>d_arr_mul_22_14, 
      product(13)=>d_arr_mul_22_13, product(12)=>d_arr_mul_22_12, 
      product(11)=>d_arr_mul_22_11, product(10)=>d_arr_mul_22_10, product(9)
      =>d_arr_mul_22_9, product(8)=>d_arr_mul_22_8, product(7)=>
      d_arr_mul_22_7, product(6)=>d_arr_mul_22_6, product(5)=>d_arr_mul_22_5, 
      product(4)=>d_arr_mul_22_4, product(3)=>d_arr_mul_22_3, product(2)=>
      d_arr_mul_22_2, product(1)=>d_arr_mul_22_1, product(0)=>d_arr_mul_22_0, 
      clk=>clk);
   mul_layer_gen_multipliers_gen_23_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>img_data_23_15, M(14)=>
      nx19446, M(13)=>img_data_23_13, M(12)=>img_data_23_12, M(11)=>
      img_data_23_11, M(10)=>img_data_23_10, M(9)=>img_data_23_9, M(8)=>
      img_data_23_8, M(7)=>img_data_23_7, M(6)=>img_data_23_6, M(5)=>
      img_data_23_5, M(4)=>img_data_23_4, M(3)=>img_data_23_3, M(2)=>
      img_data_23_2, M(1)=>img_data_23_1, M(0)=>img_data_23_0, R(15)=>
      filter_data_23_15, R(14)=>filter_data_23_14, R(13)=>filter_data_23_13, 
      R(12)=>filter_data_23_12, R(11)=>filter_data_23_11, R(10)=>
      filter_data_23_10, R(9)=>filter_data_23_9, R(8)=>filter_data_23_8, 
      R(7)=>filter_data_23_7, R(6)=>filter_data_23_6, R(5)=>filter_data_23_5, 
      R(4)=>filter_data_23_4, R(3)=>filter_data_23_3, R(2)=>filter_data_23_2, 
      R(1)=>filter_data_23_1, R(0)=>filter_data_23_0, cnt_enable=>nx16479, 
      product(31)=>d_arr_mul_23_31, product(30)=>d_arr_mul_23_30, 
      product(29)=>d_arr_mul_23_29, product(28)=>d_arr_mul_23_28, 
      product(27)=>d_arr_mul_23_27, product(26)=>d_arr_mul_23_26, 
      product(25)=>d_arr_mul_23_25, product(24)=>d_arr_mul_23_24, 
      product(23)=>d_arr_mul_23_23, product(22)=>d_arr_mul_23_22, 
      product(21)=>d_arr_mul_23_21, product(20)=>d_arr_mul_23_20, 
      product(19)=>d_arr_mul_23_19, product(18)=>d_arr_mul_23_18, 
      product(17)=>d_arr_mul_23_17, product(16)=>d_arr_mul_23_16, 
      product(15)=>d_arr_mul_23_15, product(14)=>d_arr_mul_23_14, 
      product(13)=>d_arr_mul_23_13, product(12)=>d_arr_mul_23_12, 
      product(11)=>d_arr_mul_23_11, product(10)=>d_arr_mul_23_10, product(9)
      =>d_arr_mul_23_9, product(8)=>d_arr_mul_23_8, product(7)=>
      d_arr_mul_23_7, product(6)=>d_arr_mul_23_6, product(5)=>d_arr_mul_23_5, 
      product(4)=>d_arr_mul_23_4, product(3)=>d_arr_mul_23_3, product(2)=>
      d_arr_mul_23_2, product(1)=>d_arr_mul_23_1, product(0)=>d_arr_mul_23_0, 
      clk=>clk);
   mul_layer_gen_multipliers_gen_24_mul_gen_mul_gen : 
      ModifiedBoothMultiplier port map ( M(15)=>img_data_24_15, M(14)=>
      img_data_24_14, M(13)=>img_data_24_13, M(12)=>img_data_24_12, M(11)=>
      img_data_24_11, M(10)=>img_data_24_10, M(9)=>img_data_24_9, M(8)=>
      img_data_24_8, M(7)=>img_data_24_7, M(6)=>img_data_24_6, M(5)=>
      img_data_24_5, M(4)=>img_data_24_4, M(3)=>img_data_24_3, M(2)=>
      img_data_24_2, M(1)=>img_data_24_1, M(0)=>img_data_24_0, R(15)=>
      filter_data_24_15, R(14)=>filter_data_24_14, R(13)=>filter_data_24_13, 
      R(12)=>filter_data_24_12, R(11)=>filter_data_24_11, R(10)=>
      filter_data_24_10, R(9)=>filter_data_24_9, R(8)=>filter_data_24_8, 
      R(7)=>filter_data_24_7, R(6)=>filter_data_24_6, R(5)=>filter_data_24_5, 
      R(4)=>filter_data_24_4, R(3)=>filter_data_24_3, R(2)=>filter_data_24_2, 
      R(1)=>filter_data_24_1, R(0)=>filter_data_24_0, cnt_enable=>nx16481, 
      product(31)=>d_arr_mul_24_31, product(30)=>d_arr_mul_24_30, 
      product(29)=>d_arr_mul_24_29, product(28)=>d_arr_mul_24_28, 
      product(27)=>d_arr_mul_24_27, product(26)=>d_arr_mul_24_26, 
      product(25)=>d_arr_mul_24_25, product(24)=>d_arr_mul_24_24, 
      product(23)=>d_arr_mul_24_23, product(22)=>d_arr_mul_24_22, 
      product(21)=>d_arr_mul_24_21, product(20)=>d_arr_mul_24_20, 
      product(19)=>d_arr_mul_24_19, product(18)=>d_arr_mul_24_18, 
      product(17)=>d_arr_mul_24_17, product(16)=>d_arr_mul_24_16, 
      product(15)=>d_arr_mul_24_15, product(14)=>d_arr_mul_24_14, 
      product(13)=>d_arr_mul_24_13, product(12)=>d_arr_mul_24_12, 
      product(11)=>d_arr_mul_24_11, product(10)=>d_arr_mul_24_10, product(9)
      =>d_arr_mul_24_9, product(8)=>d_arr_mul_24_8, product(7)=>
      d_arr_mul_24_7, product(6)=>d_arr_mul_24_6, product(5)=>d_arr_mul_24_5, 
      product(4)=>d_arr_mul_24_4, product(3)=>d_arr_mul_24_3, product(2)=>
      d_arr_mul_24_2, product(1)=>d_arr_mul_24_1, product(0)=>d_arr_mul_24_0, 
      clk=>clk);
   add_layer_gen_op9tree1_gen_loop_0_adder_gen : NAdder_32 port map ( a(31)
      =>nx19448, a(30)=>nx16499, a(29)=>nx16503, a(28)=>nx16507, a(27)=>
      nx16511, a(26)=>nx16515, a(25)=>nx16519, a(24)=>nx16523, a(23)=>
      nx16527, a(22)=>nx16531, a(21)=>nx16535, a(20)=>nx16539, a(19)=>
      nx16543, a(18)=>nx16547, a(17)=>nx16551, a(16)=>nx16555, a(15)=>
      nx16559, a(14)=>nx16563, a(13)=>nx16567, a(12)=>nx16571, a(11)=>
      nx16575, a(10)=>nx16579, a(9)=>nx16583, a(8)=>nx16587, a(7)=>nx16591, 
      a(6)=>nx16595, a(5)=>nx16599, a(4)=>nx16601, a(3)=>nx16603, a(2)=>
      q_arr_0_2, a(1)=>q_arr_0_1, a(0)=>nx16607, b(31)=>q_arr_1_31, b(30)=>
      q_arr_1_30, b(29)=>q_arr_1_29, b(28)=>q_arr_1_28, b(27)=>nx19450, 
      b(26)=>nx19454, b(25)=>q_arr_1_25, b(24)=>nx19458, b(23)=>q_arr_1_23, 
      b(22)=>q_arr_1_22, b(21)=>q_arr_1_21, b(20)=>q_arr_1_20, b(19)=>
      q_arr_1_19, b(18)=>nx19462, b(17)=>nx19466, b(16)=>nx19470, b(15)=>
      q_arr_1_15, b(14)=>nx19474, b(13)=>q_arr_1_13, b(12)=>nx19476, b(11)=>
      q_arr_1_11, b(10)=>nx19478, b(9)=>q_arr_1_9, b(8)=>nx19482, b(7)=>
      nx19486, b(6)=>q_arr_1_6, b(5)=>q_arr_1_5, b(4)=>q_arr_1_4, b(3)=>
      q_arr_1_3, b(2)=>q_arr_1_2, b(1)=>q_arr_1_1, b(0)=>q_arr_1_0, cin=>
      GND0, s(31)=>d_arr_add_0_31, s(30)=>d_arr_add_0_30, s(29)=>
      d_arr_add_0_29, s(28)=>d_arr_add_0_28, s(27)=>d_arr_add_0_27, s(26)=>
      d_arr_add_0_26, s(25)=>d_arr_add_0_25, s(24)=>d_arr_add_0_24, s(23)=>
      d_arr_add_0_23, s(22)=>d_arr_add_0_22, s(21)=>d_arr_add_0_21, s(20)=>
      d_arr_add_0_20, s(19)=>d_arr_add_0_19, s(18)=>d_arr_add_0_18, s(17)=>
      d_arr_add_0_17, s(16)=>d_arr_add_0_16, s(15)=>d_arr_add_0_15, s(14)=>
      d_arr_add_0_14, s(13)=>d_arr_add_0_13, s(12)=>d_arr_add_0_12, s(11)=>
      d_arr_add_0_11, s(10)=>d_arr_add_0_10, s(9)=>d_arr_add_0_9, s(8)=>
      d_arr_add_0_8, s(7)=>d_arr_add_0_7, s(6)=>d_arr_add_0_6, s(5)=>
      d_arr_add_0_5, s(4)=>d_arr_add_0_4, s(3)=>d_arr_add_0_3, s(2)=>
      d_arr_add_0_2, s(1)=>d_arr_add_0_1, s(0)=>d_arr_add_0_0, cout=>
      DANGLING(2690));
   add_layer_gen_op9tree1_gen_loop_1_adder_gen : NAdder_32 port map ( a(31)
      =>q_arr_2_31, a(30)=>q_arr_2_30, a(29)=>q_arr_2_29, a(28)=>q_arr_2_28, 
      a(27)=>q_arr_2_27, a(26)=>q_arr_2_26, a(25)=>q_arr_2_25, a(24)=>
      q_arr_2_24, a(23)=>q_arr_2_23, a(22)=>q_arr_2_22, a(21)=>q_arr_2_21, 
      a(20)=>q_arr_2_20, a(19)=>q_arr_2_19, a(18)=>q_arr_2_18, a(17)=>
      q_arr_2_17, a(16)=>q_arr_2_16, a(15)=>q_arr_2_15, a(14)=>q_arr_2_14, 
      a(13)=>q_arr_2_13, a(12)=>q_arr_2_12, a(11)=>q_arr_2_11, a(10)=>
      q_arr_2_10, a(9)=>q_arr_2_9, a(8)=>q_arr_2_8, a(7)=>q_arr_2_7, a(6)=>
      q_arr_2_6, a(5)=>q_arr_2_5, a(4)=>q_arr_2_4, a(3)=>q_arr_2_3, a(2)=>
      q_arr_2_2, a(1)=>q_arr_2_1, a(0)=>q_arr_2_0, b(31)=>q_arr_3_31, b(30)
      =>q_arr_3_30, b(29)=>q_arr_3_29, b(28)=>q_arr_3_28, b(27)=>q_arr_3_27, 
      b(26)=>q_arr_3_26, b(25)=>q_arr_3_25, b(24)=>q_arr_3_24, b(23)=>
      q_arr_3_23, b(22)=>q_arr_3_22, b(21)=>q_arr_3_21, b(20)=>q_arr_3_20, 
      b(19)=>q_arr_3_19, b(18)=>q_arr_3_18, b(17)=>q_arr_3_17, b(16)=>
      q_arr_3_16, b(15)=>q_arr_3_15, b(14)=>q_arr_3_14, b(13)=>q_arr_3_13, 
      b(12)=>q_arr_3_12, b(11)=>q_arr_3_11, b(10)=>q_arr_3_10, b(9)=>
      q_arr_3_9, b(8)=>q_arr_3_8, b(7)=>q_arr_3_7, b(6)=>q_arr_3_6, b(5)=>
      q_arr_3_5, b(4)=>q_arr_3_4, b(3)=>q_arr_3_3, b(2)=>q_arr_3_2, b(1)=>
      q_arr_3_1, b(0)=>q_arr_3_0, cin=>GND0, s(31)=>d_arr_add_1_31, s(30)=>
      d_arr_add_1_30, s(29)=>d_arr_add_1_29, s(28)=>d_arr_add_1_28, s(27)=>
      d_arr_add_1_27, s(26)=>d_arr_add_1_26, s(25)=>d_arr_add_1_25, s(24)=>
      d_arr_add_1_24, s(23)=>d_arr_add_1_23, s(22)=>d_arr_add_1_22, s(21)=>
      d_arr_add_1_21, s(20)=>d_arr_add_1_20, s(19)=>d_arr_add_1_19, s(18)=>
      d_arr_add_1_18, s(17)=>d_arr_add_1_17, s(16)=>d_arr_add_1_16, s(15)=>
      d_arr_add_1_15, s(14)=>d_arr_add_1_14, s(13)=>d_arr_add_1_13, s(12)=>
      d_arr_add_1_12, s(11)=>d_arr_add_1_11, s(10)=>d_arr_add_1_10, s(9)=>
      d_arr_add_1_9, s(8)=>d_arr_add_1_8, s(7)=>d_arr_add_1_7, s(6)=>
      d_arr_add_1_6, s(5)=>d_arr_add_1_5, s(4)=>d_arr_add_1_4, s(3)=>
      d_arr_add_1_3, s(2)=>d_arr_add_1_2, s(1)=>d_arr_add_1_1, s(0)=>
      d_arr_add_1_0, cout=>DANGLING(2691));
   add_layer_gen_op9tree1_gen_loop_2_adder_gen : NAdder_32 port map ( a(31)
      =>q_arr_4_31, a(30)=>q_arr_4_30, a(29)=>q_arr_4_29, a(28)=>q_arr_4_28, 
      a(27)=>q_arr_4_27, a(26)=>q_arr_4_26, a(25)=>q_arr_4_25, a(24)=>
      q_arr_4_24, a(23)=>q_arr_4_23, a(22)=>q_arr_4_22, a(21)=>q_arr_4_21, 
      a(20)=>q_arr_4_20, a(19)=>q_arr_4_19, a(18)=>q_arr_4_18, a(17)=>
      q_arr_4_17, a(16)=>q_arr_4_16, a(15)=>q_arr_4_15, a(14)=>q_arr_4_14, 
      a(13)=>q_arr_4_13, a(12)=>q_arr_4_12, a(11)=>q_arr_4_11, a(10)=>
      q_arr_4_10, a(9)=>q_arr_4_9, a(8)=>q_arr_4_8, a(7)=>q_arr_4_7, a(6)=>
      q_arr_4_6, a(5)=>q_arr_4_5, a(4)=>q_arr_4_4, a(3)=>q_arr_4_3, a(2)=>
      q_arr_4_2, a(1)=>q_arr_4_1, a(0)=>q_arr_4_0, b(31)=>q_arr_5_31, b(30)
      =>q_arr_5_30, b(29)=>q_arr_5_29, b(28)=>q_arr_5_28, b(27)=>q_arr_5_27, 
      b(26)=>q_arr_5_26, b(25)=>q_arr_5_25, b(24)=>q_arr_5_24, b(23)=>
      q_arr_5_23, b(22)=>q_arr_5_22, b(21)=>q_arr_5_21, b(20)=>q_arr_5_20, 
      b(19)=>q_arr_5_19, b(18)=>q_arr_5_18, b(17)=>q_arr_5_17, b(16)=>
      q_arr_5_16, b(15)=>q_arr_5_15, b(14)=>q_arr_5_14, b(13)=>q_arr_5_13, 
      b(12)=>q_arr_5_12, b(11)=>q_arr_5_11, b(10)=>q_arr_5_10, b(9)=>
      q_arr_5_9, b(8)=>q_arr_5_8, b(7)=>q_arr_5_7, b(6)=>q_arr_5_6, b(5)=>
      q_arr_5_5, b(4)=>q_arr_5_4, b(3)=>q_arr_5_3, b(2)=>q_arr_5_2, b(1)=>
      q_arr_5_1, b(0)=>q_arr_5_0, cin=>GND0, s(31)=>d_arr_add_2_31, s(30)=>
      d_arr_add_2_30, s(29)=>d_arr_add_2_29, s(28)=>d_arr_add_2_28, s(27)=>
      d_arr_add_2_27, s(26)=>d_arr_add_2_26, s(25)=>d_arr_add_2_25, s(24)=>
      d_arr_add_2_24, s(23)=>d_arr_add_2_23, s(22)=>d_arr_add_2_22, s(21)=>
      d_arr_add_2_21, s(20)=>d_arr_add_2_20, s(19)=>d_arr_add_2_19, s(18)=>
      d_arr_add_2_18, s(17)=>d_arr_add_2_17, s(16)=>d_arr_add_2_16, s(15)=>
      d_arr_add_2_15, s(14)=>d_arr_add_2_14, s(13)=>d_arr_add_2_13, s(12)=>
      d_arr_add_2_12, s(11)=>d_arr_add_2_11, s(10)=>d_arr_add_2_10, s(9)=>
      d_arr_add_2_9, s(8)=>d_arr_add_2_8, s(7)=>d_arr_add_2_7, s(6)=>
      d_arr_add_2_6, s(5)=>d_arr_add_2_5, s(4)=>d_arr_add_2_4, s(3)=>
      d_arr_add_2_3, s(2)=>d_arr_add_2_2, s(1)=>d_arr_add_2_1, s(0)=>
      d_arr_add_2_0, cout=>DANGLING(2692));
   add_layer_gen_op9tree1_gen_loop_3_adder_gen : NAdder_32 port map ( a(31)
      =>q_arr_6_31, a(30)=>q_arr_6_30, a(29)=>q_arr_6_29, a(28)=>q_arr_6_28, 
      a(27)=>q_arr_6_27, a(26)=>q_arr_6_26, a(25)=>q_arr_6_25, a(24)=>
      q_arr_6_24, a(23)=>q_arr_6_23, a(22)=>q_arr_6_22, a(21)=>q_arr_6_21, 
      a(20)=>q_arr_6_20, a(19)=>q_arr_6_19, a(18)=>q_arr_6_18, a(17)=>
      q_arr_6_17, a(16)=>q_arr_6_16, a(15)=>q_arr_6_15, a(14)=>q_arr_6_14, 
      a(13)=>q_arr_6_13, a(12)=>q_arr_6_12, a(11)=>q_arr_6_11, a(10)=>
      q_arr_6_10, a(9)=>q_arr_6_9, a(8)=>q_arr_6_8, a(7)=>q_arr_6_7, a(6)=>
      q_arr_6_6, a(5)=>q_arr_6_5, a(4)=>q_arr_6_4, a(3)=>q_arr_6_3, a(2)=>
      q_arr_6_2, a(1)=>q_arr_6_1, a(0)=>q_arr_6_0, b(31)=>q_arr_7_31, b(30)
      =>q_arr_7_30, b(29)=>q_arr_7_29, b(28)=>q_arr_7_28, b(27)=>q_arr_7_27, 
      b(26)=>q_arr_7_26, b(25)=>q_arr_7_25, b(24)=>q_arr_7_24, b(23)=>
      q_arr_7_23, b(22)=>q_arr_7_22, b(21)=>q_arr_7_21, b(20)=>q_arr_7_20, 
      b(19)=>q_arr_7_19, b(18)=>q_arr_7_18, b(17)=>q_arr_7_17, b(16)=>
      q_arr_7_16, b(15)=>q_arr_7_15, b(14)=>q_arr_7_14, b(13)=>q_arr_7_13, 
      b(12)=>q_arr_7_12, b(11)=>q_arr_7_11, b(10)=>q_arr_7_10, b(9)=>
      q_arr_7_9, b(8)=>q_arr_7_8, b(7)=>q_arr_7_7, b(6)=>q_arr_7_6, b(5)=>
      q_arr_7_5, b(4)=>q_arr_7_4, b(3)=>q_arr_7_3, b(2)=>q_arr_7_2, b(1)=>
      q_arr_7_1, b(0)=>q_arr_7_0, cin=>GND0, s(31)=>d_arr_add_3_31, s(30)=>
      d_arr_add_3_30, s(29)=>d_arr_add_3_29, s(28)=>d_arr_add_3_28, s(27)=>
      d_arr_add_3_27, s(26)=>d_arr_add_3_26, s(25)=>d_arr_add_3_25, s(24)=>
      d_arr_add_3_24, s(23)=>d_arr_add_3_23, s(22)=>d_arr_add_3_22, s(21)=>
      d_arr_add_3_21, s(20)=>d_arr_add_3_20, s(19)=>d_arr_add_3_19, s(18)=>
      d_arr_add_3_18, s(17)=>d_arr_add_3_17, s(16)=>d_arr_add_3_16, s(15)=>
      d_arr_add_3_15, s(14)=>d_arr_add_3_14, s(13)=>d_arr_add_3_13, s(12)=>
      d_arr_add_3_12, s(11)=>d_arr_add_3_11, s(10)=>d_arr_add_3_10, s(9)=>
      d_arr_add_3_9, s(8)=>d_arr_add_3_8, s(7)=>d_arr_add_3_7, s(6)=>
      d_arr_add_3_6, s(5)=>d_arr_add_3_5, s(4)=>d_arr_add_3_4, s(3)=>
      d_arr_add_3_3, s(2)=>d_arr_add_3_2, s(1)=>d_arr_add_3_1, s(0)=>
      d_arr_add_3_0, cout=>DANGLING(2693));
   add_layer_gen_op9tree2_gen_loop_0_adder_gen : NAdder_32 port map ( a(31)
      =>q_arr_9_31, a(30)=>q_arr_9_30, a(29)=>q_arr_9_29, a(28)=>q_arr_9_28, 
      a(27)=>q_arr_9_27, a(26)=>q_arr_9_26, a(25)=>q_arr_9_25, a(24)=>
      q_arr_9_24, a(23)=>q_arr_9_23, a(22)=>q_arr_9_22, a(21)=>q_arr_9_21, 
      a(20)=>q_arr_9_20, a(19)=>q_arr_9_19, a(18)=>q_arr_9_18, a(17)=>
      q_arr_9_17, a(16)=>q_arr_9_16, a(15)=>q_arr_9_15, a(14)=>q_arr_9_14, 
      a(13)=>q_arr_9_13, a(12)=>q_arr_9_12, a(11)=>q_arr_9_11, a(10)=>
      q_arr_9_10, a(9)=>q_arr_9_9, a(8)=>q_arr_9_8, a(7)=>q_arr_9_7, a(6)=>
      q_arr_9_6, a(5)=>q_arr_9_5, a(4)=>q_arr_9_4, a(3)=>q_arr_9_3, a(2)=>
      q_arr_9_2, a(1)=>q_arr_9_1, a(0)=>q_arr_9_0, b(31)=>q_arr_10_31, b(30)
      =>q_arr_10_30, b(29)=>q_arr_10_29, b(28)=>q_arr_10_28, b(27)=>
      q_arr_10_27, b(26)=>q_arr_10_26, b(25)=>q_arr_10_25, b(24)=>
      q_arr_10_24, b(23)=>q_arr_10_23, b(22)=>q_arr_10_22, b(21)=>
      q_arr_10_21, b(20)=>q_arr_10_20, b(19)=>q_arr_10_19, b(18)=>
      q_arr_10_18, b(17)=>q_arr_10_17, b(16)=>q_arr_10_16, b(15)=>
      q_arr_10_15, b(14)=>q_arr_10_14, b(13)=>q_arr_10_13, b(12)=>
      q_arr_10_12, b(11)=>q_arr_10_11, b(10)=>q_arr_10_10, b(9)=>q_arr_10_9, 
      b(8)=>q_arr_10_8, b(7)=>q_arr_10_7, b(6)=>q_arr_10_6, b(5)=>q_arr_10_5, 
      b(4)=>q_arr_10_4, b(3)=>q_arr_10_3, b(2)=>q_arr_10_2, b(1)=>q_arr_10_1, 
      b(0)=>q_arr_10_0, cin=>GND0, s(31)=>d_arr_add_9_31, s(30)=>
      d_arr_add_9_30, s(29)=>d_arr_add_9_29, s(28)=>d_arr_add_9_28, s(27)=>
      d_arr_add_9_27, s(26)=>d_arr_add_9_26, s(25)=>d_arr_add_9_25, s(24)=>
      d_arr_add_9_24, s(23)=>d_arr_add_9_23, s(22)=>d_arr_add_9_22, s(21)=>
      d_arr_add_9_21, s(20)=>d_arr_add_9_20, s(19)=>d_arr_add_9_19, s(18)=>
      d_arr_add_9_18, s(17)=>d_arr_add_9_17, s(16)=>d_arr_add_9_16, s(15)=>
      d_arr_add_9_15, s(14)=>d_arr_add_9_14, s(13)=>d_arr_add_9_13, s(12)=>
      d_arr_add_9_12, s(11)=>d_arr_add_9_11, s(10)=>d_arr_add_9_10, s(9)=>
      d_arr_add_9_9, s(8)=>d_arr_add_9_8, s(7)=>d_arr_add_9_7, s(6)=>
      d_arr_add_9_6, s(5)=>d_arr_add_9_5, s(4)=>d_arr_add_9_4, s(3)=>
      d_arr_add_9_3, s(2)=>d_arr_add_9_2, s(1)=>d_arr_add_9_1, s(0)=>
      d_arr_add_9_0, cout=>DANGLING(2694));
   add_layer_gen_op9tree2_gen_loop_1_adder_gen : NAdder_32 port map ( a(31)
      =>q_arr_11_31, a(30)=>q_arr_11_30, a(29)=>q_arr_11_29, a(28)=>
      q_arr_11_28, a(27)=>q_arr_11_27, a(26)=>q_arr_11_26, a(25)=>
      q_arr_11_25, a(24)=>q_arr_11_24, a(23)=>q_arr_11_23, a(22)=>
      q_arr_11_22, a(21)=>q_arr_11_21, a(20)=>q_arr_11_20, a(19)=>
      q_arr_11_19, a(18)=>q_arr_11_18, a(17)=>q_arr_11_17, a(16)=>
      q_arr_11_16, a(15)=>q_arr_11_15, a(14)=>q_arr_11_14, a(13)=>
      q_arr_11_13, a(12)=>q_arr_11_12, a(11)=>q_arr_11_11, a(10)=>
      q_arr_11_10, a(9)=>q_arr_11_9, a(8)=>q_arr_11_8, a(7)=>q_arr_11_7, 
      a(6)=>q_arr_11_6, a(5)=>q_arr_11_5, a(4)=>q_arr_11_4, a(3)=>q_arr_11_3, 
      a(2)=>q_arr_11_2, a(1)=>q_arr_11_1, a(0)=>q_arr_11_0, b(31)=>
      q_arr_12_31, b(30)=>q_arr_12_30, b(29)=>q_arr_12_29, b(28)=>
      q_arr_12_28, b(27)=>q_arr_12_27, b(26)=>q_arr_12_26, b(25)=>
      q_arr_12_25, b(24)=>q_arr_12_24, b(23)=>q_arr_12_23, b(22)=>
      q_arr_12_22, b(21)=>q_arr_12_21, b(20)=>q_arr_12_20, b(19)=>
      q_arr_12_19, b(18)=>q_arr_12_18, b(17)=>q_arr_12_17, b(16)=>
      q_arr_12_16, b(15)=>q_arr_12_15, b(14)=>q_arr_12_14, b(13)=>
      q_arr_12_13, b(12)=>q_arr_12_12, b(11)=>q_arr_12_11, b(10)=>
      q_arr_12_10, b(9)=>q_arr_12_9, b(8)=>q_arr_12_8, b(7)=>q_arr_12_7, 
      b(6)=>q_arr_12_6, b(5)=>q_arr_12_5, b(4)=>q_arr_12_4, b(3)=>q_arr_12_3, 
      b(2)=>q_arr_12_2, b(1)=>q_arr_12_1, b(0)=>q_arr_12_0, cin=>GND0, s(31)
      =>d_arr_add_10_31, s(30)=>d_arr_add_10_30, s(29)=>d_arr_add_10_29, 
      s(28)=>d_arr_add_10_28, s(27)=>d_arr_add_10_27, s(26)=>d_arr_add_10_26, 
      s(25)=>d_arr_add_10_25, s(24)=>d_arr_add_10_24, s(23)=>d_arr_add_10_23, 
      s(22)=>d_arr_add_10_22, s(21)=>d_arr_add_10_21, s(20)=>d_arr_add_10_20, 
      s(19)=>d_arr_add_10_19, s(18)=>d_arr_add_10_18, s(17)=>d_arr_add_10_17, 
      s(16)=>d_arr_add_10_16, s(15)=>d_arr_add_10_15, s(14)=>d_arr_add_10_14, 
      s(13)=>d_arr_add_10_13, s(12)=>d_arr_add_10_12, s(11)=>d_arr_add_10_11, 
      s(10)=>d_arr_add_10_10, s(9)=>d_arr_add_10_9, s(8)=>d_arr_add_10_8, 
      s(7)=>d_arr_add_10_7, s(6)=>d_arr_add_10_6, s(5)=>d_arr_add_10_5, s(4)
      =>d_arr_add_10_4, s(3)=>d_arr_add_10_3, s(2)=>d_arr_add_10_2, s(1)=>
      d_arr_add_10_1, s(0)=>d_arr_add_10_0, cout=>DANGLING(2695));
   add_layer_gen_op9tree2_gen_loop_2_adder_gen : NAdder_32 port map ( a(31)
      =>q_arr_13_31, a(30)=>q_arr_13_30, a(29)=>q_arr_13_29, a(28)=>
      q_arr_13_28, a(27)=>q_arr_13_27, a(26)=>q_arr_13_26, a(25)=>
      q_arr_13_25, a(24)=>q_arr_13_24, a(23)=>q_arr_13_23, a(22)=>
      q_arr_13_22, a(21)=>q_arr_13_21, a(20)=>q_arr_13_20, a(19)=>
      q_arr_13_19, a(18)=>q_arr_13_18, a(17)=>q_arr_13_17, a(16)=>
      q_arr_13_16, a(15)=>q_arr_13_15, a(14)=>q_arr_13_14, a(13)=>
      q_arr_13_13, a(12)=>q_arr_13_12, a(11)=>q_arr_13_11, a(10)=>
      q_arr_13_10, a(9)=>q_arr_13_9, a(8)=>q_arr_13_8, a(7)=>q_arr_13_7, 
      a(6)=>q_arr_13_6, a(5)=>q_arr_13_5, a(4)=>q_arr_13_4, a(3)=>q_arr_13_3, 
      a(2)=>q_arr_13_2, a(1)=>q_arr_13_1, a(0)=>q_arr_13_0, b(31)=>
      q_arr_14_31, b(30)=>q_arr_14_30, b(29)=>q_arr_14_29, b(28)=>
      q_arr_14_28, b(27)=>q_arr_14_27, b(26)=>q_arr_14_26, b(25)=>
      q_arr_14_25, b(24)=>q_arr_14_24, b(23)=>q_arr_14_23, b(22)=>
      q_arr_14_22, b(21)=>q_arr_14_21, b(20)=>q_arr_14_20, b(19)=>
      q_arr_14_19, b(18)=>q_arr_14_18, b(17)=>q_arr_14_17, b(16)=>
      q_arr_14_16, b(15)=>q_arr_14_15, b(14)=>q_arr_14_14, b(13)=>
      q_arr_14_13, b(12)=>q_arr_14_12, b(11)=>q_arr_14_11, b(10)=>
      q_arr_14_10, b(9)=>q_arr_14_9, b(8)=>q_arr_14_8, b(7)=>q_arr_14_7, 
      b(6)=>q_arr_14_6, b(5)=>q_arr_14_5, b(4)=>q_arr_14_4, b(3)=>q_arr_14_3, 
      b(2)=>q_arr_14_2, b(1)=>q_arr_14_1, b(0)=>q_arr_14_0, cin=>GND0, s(31)
      =>d_arr_add_11_31, s(30)=>d_arr_add_11_30, s(29)=>d_arr_add_11_29, 
      s(28)=>d_arr_add_11_28, s(27)=>d_arr_add_11_27, s(26)=>d_arr_add_11_26, 
      s(25)=>d_arr_add_11_25, s(24)=>d_arr_add_11_24, s(23)=>d_arr_add_11_23, 
      s(22)=>d_arr_add_11_22, s(21)=>d_arr_add_11_21, s(20)=>d_arr_add_11_20, 
      s(19)=>d_arr_add_11_19, s(18)=>d_arr_add_11_18, s(17)=>d_arr_add_11_17, 
      s(16)=>d_arr_add_11_16, s(15)=>d_arr_add_11_15, s(14)=>d_arr_add_11_14, 
      s(13)=>d_arr_add_11_13, s(12)=>d_arr_add_11_12, s(11)=>d_arr_add_11_11, 
      s(10)=>d_arr_add_11_10, s(9)=>d_arr_add_11_9, s(8)=>d_arr_add_11_8, 
      s(7)=>d_arr_add_11_7, s(6)=>d_arr_add_11_6, s(5)=>d_arr_add_11_5, s(4)
      =>d_arr_add_11_4, s(3)=>d_arr_add_11_3, s(2)=>d_arr_add_11_2, s(1)=>
      d_arr_add_11_1, s(0)=>d_arr_add_11_0, cout=>DANGLING(2696));
   add_layer_gen_op9tree2_gen_loop_3_adder_gen : NAdder_32 port map ( a(31)
      =>q_arr_15_31, a(30)=>q_arr_15_30, a(29)=>q_arr_15_29, a(28)=>
      q_arr_15_28, a(27)=>q_arr_15_27, a(26)=>q_arr_15_26, a(25)=>
      q_arr_15_25, a(24)=>q_arr_15_24, a(23)=>q_arr_15_23, a(22)=>
      q_arr_15_22, a(21)=>q_arr_15_21, a(20)=>q_arr_15_20, a(19)=>
      q_arr_15_19, a(18)=>q_arr_15_18, a(17)=>q_arr_15_17, a(16)=>
      q_arr_15_16, a(15)=>q_arr_15_15, a(14)=>q_arr_15_14, a(13)=>
      q_arr_15_13, a(12)=>q_arr_15_12, a(11)=>q_arr_15_11, a(10)=>
      q_arr_15_10, a(9)=>q_arr_15_9, a(8)=>q_arr_15_8, a(7)=>q_arr_15_7, 
      a(6)=>q_arr_15_6, a(5)=>q_arr_15_5, a(4)=>q_arr_15_4, a(3)=>q_arr_15_3, 
      a(2)=>q_arr_15_2, a(1)=>q_arr_15_1, a(0)=>q_arr_15_0, b(31)=>
      q_arr_16_31, b(30)=>q_arr_16_30, b(29)=>q_arr_16_29, b(28)=>
      q_arr_16_28, b(27)=>q_arr_16_27, b(26)=>q_arr_16_26, b(25)=>
      q_arr_16_25, b(24)=>q_arr_16_24, b(23)=>q_arr_16_23, b(22)=>
      q_arr_16_22, b(21)=>q_arr_16_21, b(20)=>q_arr_16_20, b(19)=>
      q_arr_16_19, b(18)=>q_arr_16_18, b(17)=>q_arr_16_17, b(16)=>
      q_arr_16_16, b(15)=>q_arr_16_15, b(14)=>q_arr_16_14, b(13)=>
      q_arr_16_13, b(12)=>q_arr_16_12, b(11)=>q_arr_16_11, b(10)=>
      q_arr_16_10, b(9)=>q_arr_16_9, b(8)=>q_arr_16_8, b(7)=>q_arr_16_7, 
      b(6)=>q_arr_16_6, b(5)=>q_arr_16_5, b(4)=>q_arr_16_4, b(3)=>q_arr_16_3, 
      b(2)=>q_arr_16_2, b(1)=>q_arr_16_1, b(0)=>q_arr_16_0, cin=>GND0, s(31)
      =>d_arr_add_12_31, s(30)=>d_arr_add_12_30, s(29)=>d_arr_add_12_29, 
      s(28)=>d_arr_add_12_28, s(27)=>d_arr_add_12_27, s(26)=>d_arr_add_12_26, 
      s(25)=>d_arr_add_12_25, s(24)=>d_arr_add_12_24, s(23)=>d_arr_add_12_23, 
      s(22)=>d_arr_add_12_22, s(21)=>d_arr_add_12_21, s(20)=>d_arr_add_12_20, 
      s(19)=>d_arr_add_12_19, s(18)=>d_arr_add_12_18, s(17)=>d_arr_add_12_17, 
      s(16)=>d_arr_add_12_16, s(15)=>d_arr_add_12_15, s(14)=>d_arr_add_12_14, 
      s(13)=>d_arr_add_12_13, s(12)=>d_arr_add_12_12, s(11)=>d_arr_add_12_11, 
      s(10)=>d_arr_add_12_10, s(9)=>d_arr_add_12_9, s(8)=>d_arr_add_12_8, 
      s(7)=>d_arr_add_12_7, s(6)=>d_arr_add_12_6, s(5)=>d_arr_add_12_5, s(4)
      =>d_arr_add_12_4, s(3)=>d_arr_add_12_3, s(2)=>d_arr_add_12_2, s(1)=>
      d_arr_add_12_1, s(0)=>d_arr_add_12_0, cout=>DANGLING(2697));
   add_layer_gen_op7tree1_gen_loop_0_adder_gen : NAdder_32 port map ( a(31)
      =>q_arr_18_31, a(30)=>q_arr_18_30, a(29)=>q_arr_18_29, a(28)=>
      q_arr_18_28, a(27)=>nx19490, a(26)=>q_arr_18_26, a(25)=>q_arr_18_25, 
      a(24)=>nx19494, a(23)=>q_arr_18_23, a(22)=>q_arr_18_22, a(21)=>
      q_arr_18_21, a(20)=>q_arr_18_20, a(19)=>q_arr_18_19, a(18)=>
      q_arr_18_18, a(17)=>q_arr_18_17, a(16)=>q_arr_18_16, a(15)=>
      q_arr_18_15, a(14)=>q_arr_18_14, a(13)=>q_arr_18_13, a(12)=>
      q_arr_18_12, a(11)=>q_arr_18_11, a(10)=>q_arr_18_10, a(9)=>q_arr_18_9, 
      a(8)=>q_arr_18_8, a(7)=>q_arr_18_7, a(6)=>q_arr_18_6, a(5)=>q_arr_18_5, 
      a(4)=>q_arr_18_4, a(3)=>q_arr_18_3, a(2)=>q_arr_18_2, a(1)=>q_arr_18_1, 
      a(0)=>q_arr_18_0, b(31)=>q_arr_19_31, b(30)=>q_arr_19_30, b(29)=>
      q_arr_19_29, b(28)=>q_arr_19_28, b(27)=>q_arr_19_27, b(26)=>
      q_arr_19_26, b(25)=>q_arr_19_25, b(24)=>q_arr_19_24, b(23)=>
      q_arr_19_23, b(22)=>q_arr_19_22, b(21)=>q_arr_19_21, b(20)=>
      q_arr_19_20, b(19)=>q_arr_19_19, b(18)=>q_arr_19_18, b(17)=>
      q_arr_19_17, b(16)=>q_arr_19_16, b(15)=>q_arr_19_15, b(14)=>
      q_arr_19_14, b(13)=>q_arr_19_13, b(12)=>q_arr_19_12, b(11)=>
      q_arr_19_11, b(10)=>q_arr_19_10, b(9)=>q_arr_19_9, b(8)=>q_arr_19_8, 
      b(7)=>q_arr_19_7, b(6)=>q_arr_19_6, b(5)=>q_arr_19_5, b(4)=>q_arr_19_4, 
      b(3)=>q_arr_19_3, b(2)=>q_arr_19_2, b(1)=>q_arr_19_1, b(0)=>q_arr_19_0, 
      cin=>GND0, s(31)=>d_arr_add_18_31, s(30)=>d_arr_add_18_30, s(29)=>
      d_arr_add_18_29, s(28)=>d_arr_add_18_28, s(27)=>d_arr_add_18_27, s(26)
      =>d_arr_add_18_26, s(25)=>d_arr_add_18_25, s(24)=>d_arr_add_18_24, 
      s(23)=>d_arr_add_18_23, s(22)=>d_arr_add_18_22, s(21)=>d_arr_add_18_21, 
      s(20)=>d_arr_add_18_20, s(19)=>d_arr_add_18_19, s(18)=>d_arr_add_18_18, 
      s(17)=>d_arr_add_18_17, s(16)=>d_arr_add_18_16, s(15)=>d_arr_add_18_15, 
      s(14)=>d_arr_add_18_14, s(13)=>d_arr_add_18_13, s(12)=>d_arr_add_18_12, 
      s(11)=>d_arr_add_18_11, s(10)=>d_arr_add_18_10, s(9)=>d_arr_add_18_9, 
      s(8)=>d_arr_add_18_8, s(7)=>d_arr_add_18_7, s(6)=>d_arr_add_18_6, s(5)
      =>d_arr_add_18_5, s(4)=>d_arr_add_18_4, s(3)=>d_arr_add_18_3, s(2)=>
      d_arr_add_18_2, s(1)=>d_arr_add_18_1, s(0)=>d_arr_add_18_0, cout=>
      DANGLING(2698));
   add_layer_gen_op7tree1_gen_loop_1_adder_gen : NAdder_32 port map ( a(31)
      =>q_arr_20_31, a(30)=>q_arr_20_30, a(29)=>q_arr_20_29, a(28)=>
      q_arr_20_28, a(27)=>q_arr_20_27, a(26)=>q_arr_20_26, a(25)=>
      q_arr_20_25, a(24)=>q_arr_20_24, a(23)=>q_arr_20_23, a(22)=>
      q_arr_20_22, a(21)=>q_arr_20_21, a(20)=>q_arr_20_20, a(19)=>
      q_arr_20_19, a(18)=>q_arr_20_18, a(17)=>q_arr_20_17, a(16)=>
      q_arr_20_16, a(15)=>q_arr_20_15, a(14)=>q_arr_20_14, a(13)=>
      q_arr_20_13, a(12)=>q_arr_20_12, a(11)=>q_arr_20_11, a(10)=>
      q_arr_20_10, a(9)=>q_arr_20_9, a(8)=>q_arr_20_8, a(7)=>q_arr_20_7, 
      a(6)=>q_arr_20_6, a(5)=>q_arr_20_5, a(4)=>q_arr_20_4, a(3)=>q_arr_20_3, 
      a(2)=>q_arr_20_2, a(1)=>q_arr_20_1, a(0)=>q_arr_20_0, b(31)=>
      q_arr_21_31, b(30)=>q_arr_21_30, b(29)=>q_arr_21_29, b(28)=>
      q_arr_21_28, b(27)=>q_arr_21_27, b(26)=>q_arr_21_26, b(25)=>
      q_arr_21_25, b(24)=>q_arr_21_24, b(23)=>q_arr_21_23, b(22)=>
      q_arr_21_22, b(21)=>q_arr_21_21, b(20)=>q_arr_21_20, b(19)=>
      q_arr_21_19, b(18)=>q_arr_21_18, b(17)=>q_arr_21_17, b(16)=>
      q_arr_21_16, b(15)=>q_arr_21_15, b(14)=>q_arr_21_14, b(13)=>
      q_arr_21_13, b(12)=>q_arr_21_12, b(11)=>q_arr_21_11, b(10)=>
      q_arr_21_10, b(9)=>q_arr_21_9, b(8)=>q_arr_21_8, b(7)=>q_arr_21_7, 
      b(6)=>q_arr_21_6, b(5)=>q_arr_21_5, b(4)=>q_arr_21_4, b(3)=>q_arr_21_3, 
      b(2)=>q_arr_21_2, b(1)=>q_arr_21_1, b(0)=>q_arr_21_0, cin=>GND0, s(31)
      =>d_arr_add_19_31, s(30)=>d_arr_add_19_30, s(29)=>d_arr_add_19_29, 
      s(28)=>d_arr_add_19_28, s(27)=>d_arr_add_19_27, s(26)=>d_arr_add_19_26, 
      s(25)=>d_arr_add_19_25, s(24)=>d_arr_add_19_24, s(23)=>d_arr_add_19_23, 
      s(22)=>d_arr_add_19_22, s(21)=>d_arr_add_19_21, s(20)=>d_arr_add_19_20, 
      s(19)=>d_arr_add_19_19, s(18)=>d_arr_add_19_18, s(17)=>d_arr_add_19_17, 
      s(16)=>d_arr_add_19_16, s(15)=>d_arr_add_19_15, s(14)=>d_arr_add_19_14, 
      s(13)=>d_arr_add_19_13, s(12)=>d_arr_add_19_12, s(11)=>d_arr_add_19_11, 
      s(10)=>d_arr_add_19_10, s(9)=>d_arr_add_19_9, s(8)=>d_arr_add_19_8, 
      s(7)=>d_arr_add_19_7, s(6)=>d_arr_add_19_6, s(5)=>d_arr_add_19_5, s(4)
      =>d_arr_add_19_4, s(3)=>d_arr_add_19_3, s(2)=>d_arr_add_19_2, s(1)=>
      d_arr_add_19_1, s(0)=>d_arr_add_19_0, cout=>DANGLING(2699));
   add_layer_gen_op7tree1_gen_loop_2_adder_gen : NAdder_32 port map ( a(31)
      =>q_arr_22_31, a(30)=>q_arr_22_30, a(29)=>q_arr_22_29, a(28)=>
      q_arr_22_28, a(27)=>q_arr_22_27, a(26)=>q_arr_22_26, a(25)=>
      q_arr_22_25, a(24)=>q_arr_22_24, a(23)=>q_arr_22_23, a(22)=>
      q_arr_22_22, a(21)=>q_arr_22_21, a(20)=>q_arr_22_20, a(19)=>
      q_arr_22_19, a(18)=>q_arr_22_18, a(17)=>q_arr_22_17, a(16)=>
      q_arr_22_16, a(15)=>q_arr_22_15, a(14)=>q_arr_22_14, a(13)=>
      q_arr_22_13, a(12)=>q_arr_22_12, a(11)=>q_arr_22_11, a(10)=>
      q_arr_22_10, a(9)=>q_arr_22_9, a(8)=>q_arr_22_8, a(7)=>q_arr_22_7, 
      a(6)=>q_arr_22_6, a(5)=>q_arr_22_5, a(4)=>q_arr_22_4, a(3)=>q_arr_22_3, 
      a(2)=>q_arr_22_2, a(1)=>q_arr_22_1, a(0)=>q_arr_22_0, b(31)=>
      q_arr_23_31, b(30)=>q_arr_23_30, b(29)=>q_arr_23_29, b(28)=>
      q_arr_23_28, b(27)=>q_arr_23_27, b(26)=>q_arr_23_26, b(25)=>
      q_arr_23_25, b(24)=>q_arr_23_24, b(23)=>q_arr_23_23, b(22)=>
      q_arr_23_22, b(21)=>q_arr_23_21, b(20)=>q_arr_23_20, b(19)=>
      q_arr_23_19, b(18)=>q_arr_23_18, b(17)=>q_arr_23_17, b(16)=>
      q_arr_23_16, b(15)=>q_arr_23_15, b(14)=>q_arr_23_14, b(13)=>
      q_arr_23_13, b(12)=>q_arr_23_12, b(11)=>q_arr_23_11, b(10)=>
      q_arr_23_10, b(9)=>q_arr_23_9, b(8)=>q_arr_23_8, b(7)=>q_arr_23_7, 
      b(6)=>q_arr_23_6, b(5)=>q_arr_23_5, b(4)=>q_arr_23_4, b(3)=>q_arr_23_3, 
      b(2)=>q_arr_23_2, b(1)=>q_arr_23_1, b(0)=>q_arr_23_0, cin=>GND0, s(31)
      =>d_arr_add_20_31, s(30)=>d_arr_add_20_30, s(29)=>d_arr_add_20_29, 
      s(28)=>d_arr_add_20_28, s(27)=>d_arr_add_20_27, s(26)=>d_arr_add_20_26, 
      s(25)=>d_arr_add_20_25, s(24)=>d_arr_add_20_24, s(23)=>d_arr_add_20_23, 
      s(22)=>d_arr_add_20_22, s(21)=>d_arr_add_20_21, s(20)=>d_arr_add_20_20, 
      s(19)=>d_arr_add_20_19, s(18)=>d_arr_add_20_18, s(17)=>d_arr_add_20_17, 
      s(16)=>d_arr_add_20_16, s(15)=>d_arr_add_20_15, s(14)=>d_arr_add_20_14, 
      s(13)=>d_arr_add_20_13, s(12)=>d_arr_add_20_12, s(11)=>d_arr_add_20_11, 
      s(10)=>d_arr_add_20_10, s(9)=>d_arr_add_20_9, s(8)=>d_arr_add_20_8, 
      s(7)=>d_arr_add_20_7, s(6)=>d_arr_add_20_6, s(5)=>d_arr_add_20_5, s(4)
      =>d_arr_add_20_4, s(3)=>d_arr_add_20_3, s(2)=>d_arr_add_20_2, s(1)=>
      d_arr_add_20_1, s(0)=>d_arr_add_20_0, cout=>DANGLING(2700));
   merge_layer2_gen_adder1_gen : NAdder_32_unfolded0 port map ( a(31)=>GND0, 
      a(30)=>GND0, a(29)=>GND0, a(28)=>GND0, a(27)=>GND0, a(26)=>GND0, a(25)
      =>nx19448, a(24)=>nx16501, a(23)=>nx16505, a(22)=>nx16509, a(21)=>
      nx16513, a(20)=>nx16517, a(19)=>nx16521, a(18)=>nx16525, a(17)=>
      nx16529, a(16)=>nx16533, a(15)=>nx16537, a(14)=>nx16541, a(13)=>
      nx16545, a(12)=>nx16549, a(11)=>nx16553, a(10)=>nx16557, a(9)=>nx16561, 
      a(8)=>nx16565, a(7)=>nx16569, a(6)=>nx16573, a(5)=>nx16577, a(4)=>
      nx16581, a(3)=>nx16585, a(2)=>nx16589, a(1)=>nx16593, a(0)=>nx16597, 
      b(31)=>output1_init(15), b(30)=>GND0, b(29)=>GND0, b(28)=>GND0, b(27)
      =>GND0, b(26)=>GND0, b(25)=>GND0, b(24)=>GND0, b(23)=>GND0, b(22)=>
      GND0, b(21)=>GND0, b(20)=>GND0, b(19)=>GND0, b(18)=>GND0, b(17)=>GND0, 
      b(16)=>GND0, b(15)=>GND0, b(14)=>output1_init(14), b(13)=>
      output1_init(13), b(12)=>output1_init(12), b(11)=>output1_init(11), 
      b(10)=>output1_init(10), b(9)=>output1_init(9), b(8)=>output1_init(8), 
      b(7)=>output1_init(7), b(6)=>output1_init(6), b(5)=>output1_init(5), 
      b(4)=>output1_init(4), b(3)=>output1_init(3), b(2)=>output1_init(2), 
      b(1)=>output1_init(1), b(0)=>output1_init(0), cin=>GND0, s(31)=>
      d_arr_merge2_0_31, s(30)=>DANGLING(2701), s(29)=>DANGLING(2702), s(28)
      =>DANGLING(2703), s(27)=>DANGLING(2704), s(26)=>d_arr_merge2_0_26, 
      s(25)=>d_arr_merge2_0_25, s(24)=>d_arr_merge2_0_24, s(23)=>
      d_arr_merge2_0_23, s(22)=>d_arr_merge2_0_22, s(21)=>d_arr_merge2_0_21, 
      s(20)=>d_arr_merge2_0_20, s(19)=>d_arr_merge2_0_19, s(18)=>
      d_arr_merge2_0_18, s(17)=>d_arr_merge2_0_17, s(16)=>d_arr_merge2_0_16, 
      s(15)=>d_arr_merge2_0_15, s(14)=>d_arr_merge2_0_14, s(13)=>
      d_arr_merge2_0_13, s(12)=>d_arr_merge2_0_12, s(11)=>d_arr_merge2_0_11, 
      s(10)=>d_arr_merge2_0_10, s(9)=>d_arr_merge2_0_9, s(8)=>
      d_arr_merge2_0_8, s(7)=>d_arr_merge2_0_7, s(6)=>d_arr_merge2_0_6, s(5)
      =>d_arr_merge2_0_5, s(4)=>d_arr_merge2_0_4, s(3)=>d_arr_merge2_0_3, 
      s(2)=>d_arr_merge2_0_2, s(1)=>d_arr_merge2_0_1, s(0)=>d_arr_merge2_0_0, 
      cout=>DANGLING(2705));
   merge_layer2_gen_adder2_gen : NAdder_32_unfolded0 port map ( a(31)=>GND0, 
      a(30)=>GND0, a(29)=>GND0, a(28)=>GND0, a(27)=>GND0, a(26)=>GND0, a(25)
      =>q_arr_1_31, a(24)=>q_arr_1_30, a(23)=>q_arr_1_29, a(22)=>q_arr_1_28, 
      a(21)=>nx19452, a(20)=>nx19456, a(19)=>q_arr_1_25, a(18)=>nx19460, 
      a(17)=>q_arr_1_23, a(16)=>q_arr_1_22, a(15)=>q_arr_1_21, a(14)=>
      q_arr_1_20, a(13)=>q_arr_1_19, a(12)=>nx19464, a(11)=>nx19468, a(10)=>
      nx19472, a(9)=>q_arr_1_15, a(8)=>nx19474, a(7)=>q_arr_1_13, a(6)=>
      nx19476, a(5)=>q_arr_1_11, a(4)=>nx19480, a(3)=>q_arr_1_9, a(2)=>
      nx19484, a(1)=>nx19486, a(0)=>q_arr_1_6, b(31)=>output2_init(15), 
      b(30)=>GND0, b(29)=>GND0, b(28)=>GND0, b(27)=>GND0, b(26)=>GND0, b(25)
      =>GND0, b(24)=>GND0, b(23)=>GND0, b(22)=>GND0, b(21)=>GND0, b(20)=>
      GND0, b(19)=>GND0, b(18)=>GND0, b(17)=>GND0, b(16)=>GND0, b(15)=>GND0, 
      b(14)=>output2_init(14), b(13)=>output2_init(13), b(12)=>
      output2_init(12), b(11)=>output2_init(11), b(10)=>output2_init(10), 
      b(9)=>output2_init(9), b(8)=>output2_init(8), b(7)=>output2_init(7), 
      b(6)=>output2_init(6), b(5)=>output2_init(5), b(4)=>output2_init(4), 
      b(3)=>output2_init(3), b(2)=>output2_init(2), b(1)=>output2_init(1), 
      b(0)=>output2_init(0), cin=>GND0, s(31)=>d_arr_merge2_1_31, s(30)=>
      DANGLING(2706), s(29)=>DANGLING(2707), s(28)=>DANGLING(2708), s(27)=>
      DANGLING(2709), s(26)=>d_arr_merge2_1_26, s(25)=>d_arr_merge2_1_25, 
      s(24)=>d_arr_merge2_1_24, s(23)=>d_arr_merge2_1_23, s(22)=>
      d_arr_merge2_1_22, s(21)=>d_arr_merge2_1_21, s(20)=>d_arr_merge2_1_20, 
      s(19)=>d_arr_merge2_1_19, s(18)=>d_arr_merge2_1_18, s(17)=>
      d_arr_merge2_1_17, s(16)=>d_arr_merge2_1_16, s(15)=>d_arr_merge2_1_15, 
      s(14)=>d_arr_merge2_1_14, s(13)=>d_arr_merge2_1_13, s(12)=>
      d_arr_merge2_1_12, s(11)=>d_arr_merge2_1_11, s(10)=>d_arr_merge2_1_10, 
      s(9)=>d_arr_merge2_1_9, s(8)=>d_arr_merge2_1_8, s(7)=>d_arr_merge2_1_7, 
      s(6)=>d_arr_merge2_1_6, s(5)=>d_arr_merge2_1_5, s(4)=>d_arr_merge2_1_4, 
      s(3)=>d_arr_merge2_1_3, s(2)=>d_arr_merge2_1_2, s(1)=>d_arr_merge2_1_1, 
      s(0)=>d_arr_merge2_1_0, cout=>DANGLING(2710));
   ix16087 : fake_gnd port map ( Y=>GND0);
   ix201 : nand02 port map ( Y=>ready, A0=>nx16276, A1=>nx16625);
   ix16277 : nand04 port map ( Y=>nx16276, A0=>nx16278, A1=>
      buffer_ready_EXMPLR, A2=>nx16375, A3=>nx194);
   ix16246 : oai21 port map ( Y=>nx16245, A0=>nx16278, A1=>nx16617, B0=>
      nx16281);
   ix16282 : nand03 port map ( Y=>nx16281, A0=>counter_12, A1=>nx16491, A2=>
      nx16623);
   ix16236 : oai21 port map ( Y=>nx16235, A0=>nx16285, A1=>nx16617, B0=>
      nx16289);
   reg_counter_12 : dffr port map ( Q=>counter_12, QB=>nx16285, D=>nx16235, 
      CLK=>nx16483, R=>nx16611);
   ix16290 : nand03 port map ( Y=>nx16289, A0=>counter_11, A1=>nx16491, A2=>
      nx16623);
   ix16226 : oai21 port map ( Y=>nx16225, A0=>nx16293, A1=>nx16617, B0=>
      nx16295);
   reg_counter_11 : dffr port map ( Q=>counter_11, QB=>nx16293, D=>nx16225, 
      CLK=>nx16483, R=>nx16611);
   ix16296 : nand03 port map ( Y=>nx16295, A0=>counter_10, A1=>nx16491, A2=>
      nx16623);
   ix16216 : oai21 port map ( Y=>nx16215, A0=>nx16299, A1=>nx16617, B0=>
      nx16301);
   reg_counter_10 : dffr port map ( Q=>counter_10, QB=>nx16299, D=>nx16215, 
      CLK=>nx16483, R=>nx16611);
   ix16302 : nand03 port map ( Y=>nx16301, A0=>counter_9, A1=>nx16491, A2=>
      nx16623);
   reg_counter_9 : dffr port map ( Q=>counter_9, QB=>OPEN, D=>nx16205, CLK=>
      nx16487, R=>nx16615);
   ix16206 : mux21_ni port map ( Y=>nx16205, A0=>counter_9, A1=>nx92, S0=>
      nx16623);
   ix93 : oai21 port map ( Y=>nx92, A0=>nx16306, A1=>nx20, B0=>nx16366);
   reg_counter_8 : dffr port map ( Q=>OPEN, QB=>nx16306, D=>nx16195, CLK=>
      nx16485, R=>nx16613);
   ix16196 : oai21 port map ( Y=>nx16195, A0=>nx16306, A1=>nx16617, B0=>
      nx16309);
   ix16310 : nand03 port map ( Y=>nx16309, A0=>counter_7, A1=>nx16491, A2=>
      nx16623);
   ix16186 : oai21 port map ( Y=>nx16185, A0=>nx16313, A1=>nx16617, B0=>
      nx16315);
   reg_counter_7 : dffr port map ( Q=>counter_7, QB=>nx16313, D=>nx16185, 
      CLK=>nx16483, R=>nx16611);
   ix16316 : nand03 port map ( Y=>nx16315, A0=>counter_6, A1=>nx16491, A2=>
      nx16623);
   ix16176 : oai21 port map ( Y=>nx16175, A0=>nx16319, A1=>nx16617, B0=>
      nx16321);
   reg_counter_6 : dffr port map ( Q=>counter_6, QB=>nx16319, D=>nx16175, 
      CLK=>nx16483, R=>nx16611);
   ix16322 : nand03 port map ( Y=>nx16321, A0=>counter_5, A1=>nx16489, A2=>
      nx16621);
   ix16166 : oai21 port map ( Y=>nx16165, A0=>nx16325, A1=>nx16619, B0=>
      nx16327);
   reg_counter_5 : dffr port map ( Q=>counter_5, QB=>nx16325, D=>nx16165, 
      CLK=>nx16483, R=>nx16611);
   ix16328 : nand03 port map ( Y=>nx16327, A0=>counter_4, A1=>nx16489, A2=>
      nx16621);
   ix16156 : oai21 port map ( Y=>nx16155, A0=>nx16331, A1=>nx16619, B0=>
      nx16333);
   reg_counter_4 : dffr port map ( Q=>counter_4, QB=>nx16331, D=>nx16155, 
      CLK=>nx16483, R=>nx16611);
   ix16334 : nand03 port map ( Y=>nx16333, A0=>counter_3, A1=>nx16489, A2=>
      nx16621);
   ix16146 : oai21 port map ( Y=>nx16145, A0=>nx16337, A1=>nx16619, B0=>
      nx16339);
   reg_counter_3 : dffr port map ( Q=>counter_3, QB=>nx16337, D=>nx16145, 
      CLK=>nx16485, R=>nx16613);
   ix16340 : nand03 port map ( Y=>nx16339, A0=>counter_2, A1=>nx16489, A2=>
      nx16621);
   ix16136 : oai21 port map ( Y=>nx16135, A0=>nx16343, A1=>nx16619, B0=>
      nx16345);
   reg_counter_2 : dffr port map ( Q=>counter_2, QB=>nx16343, D=>nx16135, 
      CLK=>nx16485, R=>nx16613);
   ix16346 : nand03 port map ( Y=>nx16345, A0=>counter_1, A1=>nx16489, A2=>
      nx16621);
   ix16126 : oai21 port map ( Y=>nx16125, A0=>nx16349, A1=>nx16619, B0=>
      nx16351);
   reg_counter_1 : dffr port map ( Q=>counter_1, QB=>nx16349, D=>nx16125, 
      CLK=>nx16485, R=>nx16613);
   ix16352 : nand03 port map ( Y=>nx16351, A0=>nx16489, A1=>counter_0, A2=>
      nx16621);
   ix16354 : aoi21 port map ( Y=>nx16353, A0=>operation, A1=>counter_0, B0=>
      nx20);
   reg_counter_0 : dffs_ni port map ( Q=>counter_0, QB=>OPEN, D=>nx16101, 
      CLK=>nx16485, S=>nx16613);
   ix16102 : nor02ii port map ( Y=>nx16101, A0=>nx16619, A1=>counter_0);
   ix16116 : oai21 port map ( Y=>nx16115, A0=>nx16361, A1=>nx16619, B0=>
      nx16363);
   reg_counter_14 : dffr port map ( Q=>counter_14, QB=>nx16361, D=>nx16115, 
      CLK=>nx16485, R=>nx16613);
   ix16364 : nand03 port map ( Y=>nx16363, A0=>nx16489, A1=>counter_13, A2=>
      nx16621);
   reg_counter_13 : dffr port map ( Q=>counter_13, QB=>nx16278, D=>nx16245, 
      CLK=>nx16485, R=>nx16613);
   ix16367 : nand02 port map ( Y=>nx16366, A0=>operation, A1=>counter_0);
   ix153 : oai21 port map ( Y=>buffer_ready_EXMPLR, A0=>nx16481, A1=>
      counter_0, B0=>nx16625);
   ix143 : nand02 port map ( Y=>sel_mul, A0=>nx16371, A1=>nx16373);
   ix195 : nor03_2x port map ( Y=>nx194, A0=>counter_14, A1=>counter_15, A2
      =>semi_ready_EXMPLR);
   ix16256 : oai21 port map ( Y=>nx16255, A0=>nx16380, A1=>nx16625, B0=>
      nx16382);
   reg_counter_15 : dffr port map ( Q=>counter_15, QB=>nx16380, D=>nx16255, 
      CLK=>nx16487, R=>nx16615);
   ix16383 : nand03 port map ( Y=>nx16382, A0=>nx16491, A1=>counter_14, A2=>
      nx16625);
   reg_counter_16 : dffr port map ( Q=>semi_ready_EXMPLR, QB=>OPEN, D=>
      nx16265, CLK=>nx16487, R=>nx16615);
   ix16266 : oai21 port map ( Y=>nx16265, A0=>nx16386, A1=>nx16388, B0=>
      nx16390);
   ix16387 : oai21 port map ( Y=>nx16386, A0=>counter_15, A1=>nx20, B0=>
      nx16366);
   ix16389 : inv02 port map ( Y=>nx16388, A=>en);
   ix16391 : nand02 port map ( Y=>nx16390, A0=>semi_ready_EXMPLR, A1=>
      nx16388);
   ix159 : inv01 port map ( Y=>sel_add, A=>nx16375);
   ix16398 : inv01 port map ( Y=>nx16399, A=>ordered_img_data_9_31);
   ix16400 : inv02 port map ( Y=>nx16401, A=>nx16399);
   ix16402 : inv02 port map ( Y=>nx16403, A=>nx16399);
   ix16404 : inv02 port map ( Y=>nx16405, A=>nx16399);
   ix16406 : inv01 port map ( Y=>nx16407, A=>ordered_img_data_10_31);
   ix16408 : inv02 port map ( Y=>nx16409, A=>nx16407);
   ix16410 : inv02 port map ( Y=>nx16411, A=>nx16407);
   ix16412 : inv02 port map ( Y=>nx16413, A=>nx16407);
   ix16414 : inv01 port map ( Y=>nx16415, A=>ordered_img_data_11_31);
   ix16416 : inv02 port map ( Y=>nx16417, A=>nx16415);
   ix16418 : inv02 port map ( Y=>nx16419, A=>nx16415);
   ix16420 : inv02 port map ( Y=>nx16421, A=>nx16415);
   ix16422 : inv01 port map ( Y=>nx16423, A=>ordered_img_data_12_31);
   ix16424 : inv02 port map ( Y=>nx16425, A=>nx16423);
   ix16426 : inv02 port map ( Y=>nx16427, A=>nx16423);
   ix16428 : inv02 port map ( Y=>nx16429, A=>nx16423);
   ix16430 : inv01 port map ( Y=>nx16431, A=>ordered_img_data_13_31);
   ix16432 : inv02 port map ( Y=>nx16433, A=>nx16431);
   ix16434 : inv02 port map ( Y=>nx16435, A=>nx16431);
   ix16436 : inv02 port map ( Y=>nx16437, A=>nx16431);
   ix16438 : inv01 port map ( Y=>nx16439, A=>ordered_img_data_14_31);
   ix16440 : inv02 port map ( Y=>nx16441, A=>nx16439);
   ix16442 : inv02 port map ( Y=>nx16443, A=>nx16439);
   ix16444 : inv02 port map ( Y=>nx16445, A=>nx16439);
   ix16446 : inv01 port map ( Y=>nx16447, A=>ordered_img_data_15_31);
   ix16448 : inv02 port map ( Y=>nx16449, A=>nx16447);
   ix16450 : inv02 port map ( Y=>nx16451, A=>nx16447);
   ix16452 : inv02 port map ( Y=>nx16453, A=>nx16447);
   ix16454 : inv01 port map ( Y=>nx16455, A=>ordered_img_data_16_31);
   ix16456 : inv02 port map ( Y=>nx16457, A=>nx16455);
   ix16458 : inv02 port map ( Y=>nx16459, A=>nx16455);
   ix16460 : inv02 port map ( Y=>nx16461, A=>nx16455);
   ix16462 : inv01 port map ( Y=>nx16463, A=>ordered_img_data_17_31);
   ix16464 : inv02 port map ( Y=>nx16465, A=>nx16463);
   ix16466 : inv02 port map ( Y=>nx16467, A=>nx16463);
   ix16468 : inv02 port map ( Y=>nx16469, A=>nx16463);
   ix16470 : inv01 port map ( Y=>nx16471, A=>sel_mul);
   ix16472 : inv02 port map ( Y=>nx16473, A=>nx16651);
   ix16474 : inv02 port map ( Y=>nx16475, A=>nx16651);
   ix16476 : inv02 port map ( Y=>nx16477, A=>nx16651);
   ix16478 : inv02 port map ( Y=>nx16479, A=>nx16651);
   ix16480 : inv02 port map ( Y=>nx16481, A=>nx16651);
   ix16482 : inv02 port map ( Y=>nx16483, A=>clk);
   ix16484 : inv02 port map ( Y=>nx16485, A=>clk);
   ix16486 : inv02 port map ( Y=>nx16487, A=>clk);
   ix16488 : buf02 port map ( Y=>nx16489, A=>nx16353);
   ix16490 : buf02 port map ( Y=>nx16491, A=>nx16353);
   ix21 : nor02_2x port map ( Y=>nx20, A0=>compute_relu, A1=>nx16361);
   ix16372 : and04 port map ( Y=>nx16371, A0=>nx16349, A1=>nx16343, A2=>
      nx16337, A3=>nx16331);
   ix16374 : and04 port map ( Y=>nx16373, A0=>nx16325, A1=>nx16319, A2=>
      nx16313, A3=>nx16306);
   ix16376 : and04 port map ( Y=>nx16375, A0=>nx16497, A1=>nx16299, A2=>
      nx16293, A3=>nx16285);
   ix16496 : inv01 port map ( Y=>nx16497, A=>counter_9);
   ix16498 : buf02 port map ( Y=>nx16499, A=>q_arr_0_30);
   ix16500 : buf02 port map ( Y=>nx16501, A=>q_arr_0_30);
   ix16502 : buf02 port map ( Y=>nx16503, A=>q_arr_0_29);
   ix16504 : buf02 port map ( Y=>nx16505, A=>q_arr_0_29);
   ix16506 : buf02 port map ( Y=>nx16507, A=>q_arr_0_28);
   ix16508 : buf02 port map ( Y=>nx16509, A=>q_arr_0_28);
   ix16510 : buf02 port map ( Y=>nx16511, A=>q_arr_0_27);
   ix16512 : buf02 port map ( Y=>nx16513, A=>q_arr_0_27);
   ix16514 : buf02 port map ( Y=>nx16515, A=>q_arr_0_26);
   ix16516 : buf02 port map ( Y=>nx16517, A=>q_arr_0_26);
   ix16518 : buf02 port map ( Y=>nx16519, A=>q_arr_0_25);
   ix16520 : buf02 port map ( Y=>nx16521, A=>q_arr_0_25);
   ix16522 : buf02 port map ( Y=>nx16523, A=>q_arr_0_24);
   ix16524 : buf02 port map ( Y=>nx16525, A=>q_arr_0_24);
   ix16526 : buf02 port map ( Y=>nx16527, A=>q_arr_0_23);
   ix16528 : buf02 port map ( Y=>nx16529, A=>q_arr_0_23);
   ix16530 : buf02 port map ( Y=>nx16531, A=>q_arr_0_22);
   ix16532 : buf02 port map ( Y=>nx16533, A=>q_arr_0_22);
   ix16534 : buf02 port map ( Y=>nx16535, A=>q_arr_0_21);
   ix16536 : buf02 port map ( Y=>nx16537, A=>q_arr_0_21);
   ix16538 : buf02 port map ( Y=>nx16539, A=>q_arr_0_20);
   ix16540 : buf02 port map ( Y=>nx16541, A=>q_arr_0_20);
   ix16542 : buf02 port map ( Y=>nx16543, A=>q_arr_0_19);
   ix16544 : buf02 port map ( Y=>nx16545, A=>q_arr_0_19);
   ix16546 : buf02 port map ( Y=>nx16547, A=>q_arr_0_18);
   ix16548 : buf02 port map ( Y=>nx16549, A=>q_arr_0_18);
   ix16550 : buf02 port map ( Y=>nx16551, A=>q_arr_0_17);
   ix16552 : buf02 port map ( Y=>nx16553, A=>q_arr_0_17);
   ix16554 : buf02 port map ( Y=>nx16555, A=>q_arr_0_16);
   ix16556 : buf02 port map ( Y=>nx16557, A=>q_arr_0_16);
   ix16558 : buf02 port map ( Y=>nx16559, A=>q_arr_0_15);
   ix16560 : buf02 port map ( Y=>nx16561, A=>q_arr_0_15);
   ix16562 : buf02 port map ( Y=>nx16563, A=>q_arr_0_14);
   ix16564 : buf02 port map ( Y=>nx16565, A=>q_arr_0_14);
   ix16566 : buf02 port map ( Y=>nx16567, A=>q_arr_0_13);
   ix16568 : buf02 port map ( Y=>nx16569, A=>q_arr_0_13);
   ix16570 : buf02 port map ( Y=>nx16571, A=>q_arr_0_12);
   ix16572 : buf02 port map ( Y=>nx16573, A=>q_arr_0_12);
   ix16574 : buf02 port map ( Y=>nx16575, A=>q_arr_0_11);
   ix16576 : buf02 port map ( Y=>nx16577, A=>q_arr_0_11);
   ix16578 : buf02 port map ( Y=>nx16579, A=>q_arr_0_10);
   ix16580 : buf02 port map ( Y=>nx16581, A=>q_arr_0_10);
   ix16582 : buf02 port map ( Y=>nx16583, A=>q_arr_0_9);
   ix16584 : buf02 port map ( Y=>nx16585, A=>q_arr_0_9);
   ix16586 : buf02 port map ( Y=>nx16587, A=>q_arr_0_8);
   ix16588 : buf02 port map ( Y=>nx16589, A=>q_arr_0_8);
   ix16590 : buf02 port map ( Y=>nx16591, A=>q_arr_0_7);
   ix16592 : buf02 port map ( Y=>nx16593, A=>q_arr_0_7);
   ix16594 : buf02 port map ( Y=>nx16595, A=>q_arr_0_6);
   ix16596 : buf02 port map ( Y=>nx16597, A=>q_arr_0_6);
   ix16598 : buf02 port map ( Y=>nx16599, A=>q_arr_0_5);
   ix16600 : buf02 port map ( Y=>nx16601, A=>q_arr_0_4);
   ix16602 : buf02 port map ( Y=>nx16603, A=>q_arr_0_3);
   ix16604 : buf02 port map ( Y=>nx16605, A=>q_arr_0_0);
   ix16606 : buf02 port map ( Y=>nx16607, A=>q_arr_0_0);
   ix16608 : inv01 port map ( Y=>nx16609, A=>reset);
   ix16610 : inv02 port map ( Y=>nx16611, A=>nx16609);
   ix16612 : inv02 port map ( Y=>nx16613, A=>nx16609);
   ix16614 : inv02 port map ( Y=>nx16615, A=>nx16609);
   ix16616 : inv02 port map ( Y=>nx16617, A=>nx16388);
   ix16618 : inv02 port map ( Y=>nx16619, A=>nx16388);
   ix16620 : inv02 port map ( Y=>nx16621, A=>nx16388);
   ix16622 : inv02 port map ( Y=>nx16623, A=>nx16388);
   ix16624 : inv02 port map ( Y=>nx16625, A=>nx16388);
   ix16626 : inv02 port map ( Y=>nx16627, A=>nx16653);
   ix16628 : inv02 port map ( Y=>nx16629, A=>nx16653);
   ix16630 : inv02 port map ( Y=>nx16631, A=>nx16653);
   ix16632 : inv02 port map ( Y=>nx16633, A=>nx16653);
   ix16634 : inv02 port map ( Y=>nx16635, A=>nx16653);
   ix16636 : inv02 port map ( Y=>nx16637, A=>nx16471);
   ix16638 : inv02 port map ( Y=>nx16639, A=>nx16471);
   ix16640 : inv02 port map ( Y=>nx16641, A=>nx16471);
   ix16642 : inv02 port map ( Y=>nx16643, A=>nx16471);
   ix16644 : inv02 port map ( Y=>nx16645, A=>nx16471);
   ix16650 : inv01 port map ( Y=>nx16651, A=>sel_mul);
   ix16652 : inv01 port map ( Y=>nx16653, A=>sel_mul);
   ix16658 : buf02 port map ( Y=>nx16659, A=>img_data_7_15);
   ix16660 : buf02 port map ( Y=>nx16661, A=>img_data_11_15);
   ix16662 : buf02 port map ( Y=>nx16663, A=>img_data_12_15);
   ix16664 : buf02 port map ( Y=>nx16665, A=>filter_size);
   ix16666 : buf02 port map ( Y=>nx16667, A=>filter_size);
   ix19387 : buf02 port map ( Y=>nx19388, A=>q_arr_0_27);
   ix19389 : buf02 port map ( Y=>nx19390, A=>q_arr_0_24);
   ix19395 : buf02 port map ( Y=>nx19396, A=>img_data_0_14);
   ix19397 : buf02 port map ( Y=>nx19398, A=>img_data_1_14);
   ix19399 : buf02 port map ( Y=>nx19400, A=>img_data_1_14);
   ix19401 : buf02 port map ( Y=>nx19402, A=>img_data_1_10);
   ix19403 : buf02 port map ( Y=>nx19404, A=>img_data_2_14);
   ix19405 : buf02 port map ( Y=>nx19406, A=>img_data_2_14);
   ix19407 : buf02 port map ( Y=>nx19408, A=>img_data_2_10);
   ix19409 : buf02 port map ( Y=>nx19410, A=>img_data_5_14);
   ix19411 : buf02 port map ( Y=>nx19412, A=>img_data_6_14);
   ix19413 : buf02 port map ( Y=>nx19414, A=>img_data_6_14);
   ix19415 : buf02 port map ( Y=>nx19416, A=>img_data_6_10);
   ix19417 : buf02 port map ( Y=>nx19418, A=>img_data_7_14);
   ix19419 : buf02 port map ( Y=>nx19420, A=>img_data_7_14);
   ix19421 : buf02 port map ( Y=>nx19422, A=>img_data_7_10);
   ix19423 : buf02 port map ( Y=>nx19424, A=>img_data_10_14);
   ix19425 : buf02 port map ( Y=>nx19426, A=>img_data_11_14);
   ix19427 : buf02 port map ( Y=>nx19428, A=>img_data_11_14);
   ix19429 : buf02 port map ( Y=>nx19430, A=>img_data_11_10);
   ix19431 : buf02 port map ( Y=>nx19432, A=>img_data_12_14);
   ix19433 : buf02 port map ( Y=>nx19434, A=>img_data_12_14);
   ix19435 : buf02 port map ( Y=>nx19436, A=>img_data_12_10);
   ix19437 : buf02 port map ( Y=>nx19438, A=>img_data_18_14);
   ix19439 : buf02 port map ( Y=>nx19440, A=>img_data_20_14);
   ix19441 : buf02 port map ( Y=>nx19442, A=>img_data_21_14);
   ix19443 : buf02 port map ( Y=>nx19444, A=>img_data_22_14);
   ix19445 : buf02 port map ( Y=>nx19446, A=>img_data_23_14);
   ix19447 : buf02 port map ( Y=>nx19448, A=>q_arr_0_31);
   ix19449 : buf02 port map ( Y=>nx19450, A=>q_arr_1_27);
   ix19451 : buf02 port map ( Y=>nx19452, A=>q_arr_1_27);
   ix19453 : buf02 port map ( Y=>nx19454, A=>q_arr_1_26);
   ix19455 : buf02 port map ( Y=>nx19456, A=>q_arr_1_26);
   ix19457 : buf02 port map ( Y=>nx19458, A=>q_arr_1_24);
   ix19459 : buf02 port map ( Y=>nx19460, A=>q_arr_1_24);
   ix19461 : buf02 port map ( Y=>nx19462, A=>q_arr_1_18);
   ix19463 : buf02 port map ( Y=>nx19464, A=>q_arr_1_18);
   ix19465 : buf02 port map ( Y=>nx19466, A=>q_arr_1_17);
   ix19467 : buf02 port map ( Y=>nx19468, A=>q_arr_1_17);
   ix19469 : buf02 port map ( Y=>nx19470, A=>q_arr_1_16);
   ix19471 : buf02 port map ( Y=>nx19472, A=>q_arr_1_16);
   ix19473 : buf02 port map ( Y=>nx19474, A=>q_arr_1_14);
   ix19475 : buf02 port map ( Y=>nx19476, A=>q_arr_1_12);
   ix19477 : buf02 port map ( Y=>nx19478, A=>q_arr_1_10);
   ix19479 : buf02 port map ( Y=>nx19480, A=>q_arr_1_10);
   ix19481 : buf02 port map ( Y=>nx19482, A=>q_arr_1_8);
   ix19483 : buf02 port map ( Y=>nx19484, A=>q_arr_1_8);
   ix19485 : buf02 port map ( Y=>nx19486, A=>q_arr_1_7);
   ix19487 : buf02 port map ( Y=>nx19488, A=>q_arr_18_27);
   ix19489 : buf02 port map ( Y=>nx19490, A=>q_arr_18_27);
   ix19491 : buf02 port map ( Y=>nx19492, A=>q_arr_18_24);
   ix19493 : buf02 port map ( Y=>nx19494, A=>q_arr_18_24);
end Behavioral ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Queue_5_unfolded0 is
   port (
      d : IN std_logic_vector (15 DOWNTO 0) ;
      q_0_15 : OUT std_logic ;
      q_0_14 : OUT std_logic ;
      q_0_13 : OUT std_logic ;
      q_0_12 : OUT std_logic ;
      q_0_11 : OUT std_logic ;
      q_0_10 : OUT std_logic ;
      q_0_9 : OUT std_logic ;
      q_0_8 : OUT std_logic ;
      q_0_7 : OUT std_logic ;
      q_0_6 : OUT std_logic ;
      q_0_5 : OUT std_logic ;
      q_0_4 : OUT std_logic ;
      q_0_3 : OUT std_logic ;
      q_0_2 : OUT std_logic ;
      q_0_1 : OUT std_logic ;
      q_0_0 : OUT std_logic ;
      q_1_15 : OUT std_logic ;
      q_1_14 : OUT std_logic ;
      q_1_13 : OUT std_logic ;
      q_1_12 : OUT std_logic ;
      q_1_11 : OUT std_logic ;
      q_1_10 : OUT std_logic ;
      q_1_9 : OUT std_logic ;
      q_1_8 : OUT std_logic ;
      q_1_7 : OUT std_logic ;
      q_1_6 : OUT std_logic ;
      q_1_5 : OUT std_logic ;
      q_1_4 : OUT std_logic ;
      q_1_3 : OUT std_logic ;
      q_1_2 : OUT std_logic ;
      q_1_1 : OUT std_logic ;
      q_1_0 : OUT std_logic ;
      q_2_15 : OUT std_logic ;
      q_2_14 : OUT std_logic ;
      q_2_13 : OUT std_logic ;
      q_2_12 : OUT std_logic ;
      q_2_11 : OUT std_logic ;
      q_2_10 : OUT std_logic ;
      q_2_9 : OUT std_logic ;
      q_2_8 : OUT std_logic ;
      q_2_7 : OUT std_logic ;
      q_2_6 : OUT std_logic ;
      q_2_5 : OUT std_logic ;
      q_2_4 : OUT std_logic ;
      q_2_3 : OUT std_logic ;
      q_2_2 : OUT std_logic ;
      q_2_1 : OUT std_logic ;
      q_2_0 : OUT std_logic ;
      q_3_15 : OUT std_logic ;
      q_3_14 : OUT std_logic ;
      q_3_13 : OUT std_logic ;
      q_3_12 : OUT std_logic ;
      q_3_11 : OUT std_logic ;
      q_3_10 : OUT std_logic ;
      q_3_9 : OUT std_logic ;
      q_3_8 : OUT std_logic ;
      q_3_7 : OUT std_logic ;
      q_3_6 : OUT std_logic ;
      q_3_5 : OUT std_logic ;
      q_3_4 : OUT std_logic ;
      q_3_3 : OUT std_logic ;
      q_3_2 : OUT std_logic ;
      q_3_1 : OUT std_logic ;
      q_3_0 : OUT std_logic ;
      q_4_15 : OUT std_logic ;
      q_4_14 : OUT std_logic ;
      q_4_13 : OUT std_logic ;
      q_4_12 : OUT std_logic ;
      q_4_11 : OUT std_logic ;
      q_4_10 : OUT std_logic ;
      q_4_9 : OUT std_logic ;
      q_4_8 : OUT std_logic ;
      q_4_7 : OUT std_logic ;
      q_4_6 : OUT std_logic ;
      q_4_5 : OUT std_logic ;
      q_4_4 : OUT std_logic ;
      q_4_3 : OUT std_logic ;
      q_4_2 : OUT std_logic ;
      q_4_1 : OUT std_logic ;
      q_4_0 : OUT std_logic ;
      clk : IN std_logic ;
      load : IN std_logic ;
      reset : IN std_logic) ;
end Queue_5_unfolded0 ;

architecture Structural_unfold_3007 of Queue_5_unfolded0 is
   signal q_0_15_EXMPLR, q_0_14_EXMPLR, q_0_13_EXMPLR, q_0_12_EXMPLR, 
      q_0_11_EXMPLR, q_0_10_EXMPLR, q_0_9_EXMPLR, q_0_8_EXMPLR, q_0_7_EXMPLR, 
      q_0_6_EXMPLR, q_0_5_EXMPLR, q_0_4_EXMPLR, q_0_3_EXMPLR, q_0_2_EXMPLR, 
      q_0_1_EXMPLR, q_0_0_EXMPLR, q_1_15_EXMPLR, q_1_14_EXMPLR, 
      q_1_13_EXMPLR, q_1_12_EXMPLR, q_1_11_EXMPLR, q_1_10_EXMPLR, 
      q_1_9_EXMPLR, q_1_8_EXMPLR, q_1_7_EXMPLR, q_1_6_EXMPLR, q_1_5_EXMPLR, 
      q_1_4_EXMPLR, q_1_3_EXMPLR, q_1_2_EXMPLR, q_1_1_EXMPLR, q_1_0_EXMPLR, 
      q_2_15_EXMPLR, q_2_14_EXMPLR, q_2_13_EXMPLR, q_2_12_EXMPLR, 
      q_2_11_EXMPLR, q_2_10_EXMPLR, q_2_9_EXMPLR, q_2_8_EXMPLR, q_2_7_EXMPLR, 
      q_2_6_EXMPLR, q_2_5_EXMPLR, q_2_4_EXMPLR, q_2_3_EXMPLR, q_2_2_EXMPLR, 
      q_2_1_EXMPLR, q_2_0_EXMPLR, q_3_15_EXMPLR, q_3_14_EXMPLR, 
      q_3_13_EXMPLR, q_3_12_EXMPLR, q_3_11_EXMPLR, q_3_10_EXMPLR, 
      q_3_9_EXMPLR, q_3_8_EXMPLR, q_3_7_EXMPLR, q_3_6_EXMPLR, q_3_5_EXMPLR, 
      q_3_4_EXMPLR, q_3_3_EXMPLR, q_3_2_EXMPLR, q_3_1_EXMPLR, q_3_0_EXMPLR, 
      q_4_15_EXMPLR, q_4_14_EXMPLR, q_4_13_EXMPLR, q_4_12_EXMPLR, 
      q_4_11_EXMPLR, q_4_10_EXMPLR, q_4_9_EXMPLR, q_4_8_EXMPLR, q_4_7_EXMPLR, 
      q_4_6_EXMPLR, q_4_5_EXMPLR, q_4_4_EXMPLR, q_4_3_EXMPLR, q_4_2_EXMPLR, 
      q_4_1_EXMPLR, q_4_0_EXMPLR, nx240, nx250, nx260, nx270, nx280, nx290, 
      nx300, nx310, nx320, nx330, nx340, nx350, nx360, nx370, nx380, nx390, 
      nx400, nx410, nx420, nx430, nx440, nx450, nx460, nx470, nx480, nx490, 
      nx500, nx510, nx520, nx530, nx540, nx550, nx560, nx570, nx580, nx590, 
      nx600, nx610, nx620, nx630, nx640, nx650, nx660, nx670, nx680, nx690, 
      nx700, nx710, nx720, nx730, nx740, nx750, nx760, nx770, nx780, nx790, 
      nx800, nx810, nx820, nx830, nx840, nx850, nx860, nx870, nx880, nx890, 
      nx900, nx910, nx920, nx930, nx940, nx950, nx960, nx970, nx980, nx990, 
      nx1000, nx1010, nx1020, nx1030, nx1287, nx1289, nx1291, nx1293, nx1295, 
      nx1297, nx1299, nx1301, nx1303, nx1305, nx1307, nx1309, nx1313, nx1315, 
      nx1317, nx1319, nx1321, nx1323, nx1325, nx1327, nx1329, nx1331, nx1333, 
      nx1335, nx1337, nx1339, nx1341, nx1343: std_logic ;

begin
   q_0_15 <= q_0_15_EXMPLR ;
   q_0_14 <= q_0_14_EXMPLR ;
   q_0_13 <= q_0_13_EXMPLR ;
   q_0_12 <= q_0_12_EXMPLR ;
   q_0_11 <= q_0_11_EXMPLR ;
   q_0_10 <= q_0_10_EXMPLR ;
   q_0_9 <= q_0_9_EXMPLR ;
   q_0_8 <= q_0_8_EXMPLR ;
   q_0_7 <= q_0_7_EXMPLR ;
   q_0_6 <= q_0_6_EXMPLR ;
   q_0_5 <= q_0_5_EXMPLR ;
   q_0_4 <= q_0_4_EXMPLR ;
   q_0_3 <= q_0_3_EXMPLR ;
   q_0_2 <= q_0_2_EXMPLR ;
   q_0_1 <= q_0_1_EXMPLR ;
   q_0_0 <= q_0_0_EXMPLR ;
   q_1_15 <= q_1_15_EXMPLR ;
   q_1_14 <= q_1_14_EXMPLR ;
   q_1_13 <= q_1_13_EXMPLR ;
   q_1_12 <= q_1_12_EXMPLR ;
   q_1_11 <= q_1_11_EXMPLR ;
   q_1_10 <= q_1_10_EXMPLR ;
   q_1_9 <= q_1_9_EXMPLR ;
   q_1_8 <= q_1_8_EXMPLR ;
   q_1_7 <= q_1_7_EXMPLR ;
   q_1_6 <= q_1_6_EXMPLR ;
   q_1_5 <= q_1_5_EXMPLR ;
   q_1_4 <= q_1_4_EXMPLR ;
   q_1_3 <= q_1_3_EXMPLR ;
   q_1_2 <= q_1_2_EXMPLR ;
   q_1_1 <= q_1_1_EXMPLR ;
   q_1_0 <= q_1_0_EXMPLR ;
   q_2_15 <= q_2_15_EXMPLR ;
   q_2_14 <= q_2_14_EXMPLR ;
   q_2_13 <= q_2_13_EXMPLR ;
   q_2_12 <= q_2_12_EXMPLR ;
   q_2_11 <= q_2_11_EXMPLR ;
   q_2_10 <= q_2_10_EXMPLR ;
   q_2_9 <= q_2_9_EXMPLR ;
   q_2_8 <= q_2_8_EXMPLR ;
   q_2_7 <= q_2_7_EXMPLR ;
   q_2_6 <= q_2_6_EXMPLR ;
   q_2_5 <= q_2_5_EXMPLR ;
   q_2_4 <= q_2_4_EXMPLR ;
   q_2_3 <= q_2_3_EXMPLR ;
   q_2_2 <= q_2_2_EXMPLR ;
   q_2_1 <= q_2_1_EXMPLR ;
   q_2_0 <= q_2_0_EXMPLR ;
   q_3_15 <= q_3_15_EXMPLR ;
   q_3_14 <= q_3_14_EXMPLR ;
   q_3_13 <= q_3_13_EXMPLR ;
   q_3_12 <= q_3_12_EXMPLR ;
   q_3_11 <= q_3_11_EXMPLR ;
   q_3_10 <= q_3_10_EXMPLR ;
   q_3_9 <= q_3_9_EXMPLR ;
   q_3_8 <= q_3_8_EXMPLR ;
   q_3_7 <= q_3_7_EXMPLR ;
   q_3_6 <= q_3_6_EXMPLR ;
   q_3_5 <= q_3_5_EXMPLR ;
   q_3_4 <= q_3_4_EXMPLR ;
   q_3_3 <= q_3_3_EXMPLR ;
   q_3_2 <= q_3_2_EXMPLR ;
   q_3_1 <= q_3_1_EXMPLR ;
   q_3_0 <= q_3_0_EXMPLR ;
   q_4_15 <= q_4_15_EXMPLR ;
   q_4_14 <= q_4_14_EXMPLR ;
   q_4_13 <= q_4_13_EXMPLR ;
   q_4_12 <= q_4_12_EXMPLR ;
   q_4_11 <= q_4_11_EXMPLR ;
   q_4_10 <= q_4_10_EXMPLR ;
   q_4_9 <= q_4_9_EXMPLR ;
   q_4_8 <= q_4_8_EXMPLR ;
   q_4_7 <= q_4_7_EXMPLR ;
   q_4_6 <= q_4_6_EXMPLR ;
   q_4_5 <= q_4_5_EXMPLR ;
   q_4_4 <= q_4_4_EXMPLR ;
   q_4_3 <= q_4_3_EXMPLR ;
   q_4_2 <= q_4_2_EXMPLR ;
   q_4_1 <= q_4_1_EXMPLR ;
   q_4_0 <= q_4_0_EXMPLR ;
   gen_regs_4_regi_reg_q_0 : dff port map ( Q=>q_4_0_EXMPLR, QB=>OPEN, D=>
      nx280, CLK=>nx1313);
   ix281 : mux21_ni port map ( Y=>nx280, A0=>q_4_0_EXMPLR, A1=>q_3_0_EXMPLR, 
      S0=>nx1287);
   gen_regs_3_regi_reg_q_0 : dff port map ( Q=>q_3_0_EXMPLR, QB=>OPEN, D=>
      nx270, CLK=>nx1313);
   ix271 : mux21_ni port map ( Y=>nx270, A0=>q_3_0_EXMPLR, A1=>q_2_0_EXMPLR, 
      S0=>nx1287);
   gen_regs_2_regi_reg_q_0 : dff port map ( Q=>q_2_0_EXMPLR, QB=>OPEN, D=>
      nx260, CLK=>nx1313);
   ix261 : mux21_ni port map ( Y=>nx260, A0=>q_2_0_EXMPLR, A1=>q_1_0_EXMPLR, 
      S0=>nx1287);
   gen_regs_1_regi_reg_q_0 : dff port map ( Q=>q_1_0_EXMPLR, QB=>OPEN, D=>
      nx250, CLK=>nx1313);
   ix251 : mux21_ni port map ( Y=>nx250, A0=>q_1_0_EXMPLR, A1=>q_0_0_EXMPLR, 
      S0=>nx1287);
   reg0_reg_q_0 : dff port map ( Q=>q_0_0_EXMPLR, QB=>OPEN, D=>nx240, CLK=>
      nx1313);
   ix241 : mux21_ni port map ( Y=>nx240, A0=>q_0_0_EXMPLR, A1=>d(0), S0=>
      nx1287);
   gen_regs_4_regi_reg_q_1 : dff port map ( Q=>q_4_1_EXMPLR, QB=>OPEN, D=>
      nx330, CLK=>nx1315);
   ix331 : mux21_ni port map ( Y=>nx330, A0=>q_4_1_EXMPLR, A1=>q_3_1_EXMPLR, 
      S0=>nx1289);
   gen_regs_3_regi_reg_q_1 : dff port map ( Q=>q_3_1_EXMPLR, QB=>OPEN, D=>
      nx320, CLK=>nx1315);
   ix321 : mux21_ni port map ( Y=>nx320, A0=>q_3_1_EXMPLR, A1=>q_2_1_EXMPLR, 
      S0=>nx1289);
   gen_regs_2_regi_reg_q_1 : dff port map ( Q=>q_2_1_EXMPLR, QB=>OPEN, D=>
      nx310, CLK=>nx1315);
   ix311 : mux21_ni port map ( Y=>nx310, A0=>q_2_1_EXMPLR, A1=>q_1_1_EXMPLR, 
      S0=>nx1289);
   gen_regs_1_regi_reg_q_1 : dff port map ( Q=>q_1_1_EXMPLR, QB=>OPEN, D=>
      nx300, CLK=>nx1313);
   ix301 : mux21_ni port map ( Y=>nx300, A0=>q_1_1_EXMPLR, A1=>q_0_1_EXMPLR, 
      S0=>nx1287);
   reg0_reg_q_1 : dff port map ( Q=>q_0_1_EXMPLR, QB=>OPEN, D=>nx290, CLK=>
      nx1313);
   ix291 : mux21_ni port map ( Y=>nx290, A0=>q_0_1_EXMPLR, A1=>d(1), S0=>
      nx1287);
   gen_regs_4_regi_reg_q_2 : dff port map ( Q=>q_4_2_EXMPLR, QB=>OPEN, D=>
      nx380, CLK=>nx1317);
   ix381 : mux21_ni port map ( Y=>nx380, A0=>q_4_2_EXMPLR, A1=>q_3_2_EXMPLR, 
      S0=>nx1291);
   gen_regs_3_regi_reg_q_2 : dff port map ( Q=>q_3_2_EXMPLR, QB=>OPEN, D=>
      nx370, CLK=>nx1315);
   ix371 : mux21_ni port map ( Y=>nx370, A0=>q_3_2_EXMPLR, A1=>q_2_2_EXMPLR, 
      S0=>nx1289);
   gen_regs_2_regi_reg_q_2 : dff port map ( Q=>q_2_2_EXMPLR, QB=>OPEN, D=>
      nx360, CLK=>nx1315);
   ix361 : mux21_ni port map ( Y=>nx360, A0=>q_2_2_EXMPLR, A1=>q_1_2_EXMPLR, 
      S0=>nx1289);
   gen_regs_1_regi_reg_q_2 : dff port map ( Q=>q_1_2_EXMPLR, QB=>OPEN, D=>
      nx350, CLK=>nx1315);
   ix351 : mux21_ni port map ( Y=>nx350, A0=>q_1_2_EXMPLR, A1=>q_0_2_EXMPLR, 
      S0=>nx1289);
   reg0_reg_q_2 : dff port map ( Q=>q_0_2_EXMPLR, QB=>OPEN, D=>nx340, CLK=>
      nx1315);
   ix341 : mux21_ni port map ( Y=>nx340, A0=>q_0_2_EXMPLR, A1=>d(2), S0=>
      nx1289);
   gen_regs_4_regi_reg_q_3 : dff port map ( Q=>q_4_3_EXMPLR, QB=>OPEN, D=>
      nx430, CLK=>nx1317);
   ix431 : mux21_ni port map ( Y=>nx430, A0=>q_4_3_EXMPLR, A1=>q_3_3_EXMPLR, 
      S0=>nx1291);
   gen_regs_3_regi_reg_q_3 : dff port map ( Q=>q_3_3_EXMPLR, QB=>OPEN, D=>
      nx420, CLK=>nx1317);
   ix421 : mux21_ni port map ( Y=>nx420, A0=>q_3_3_EXMPLR, A1=>q_2_3_EXMPLR, 
      S0=>nx1291);
   gen_regs_2_regi_reg_q_3 : dff port map ( Q=>q_2_3_EXMPLR, QB=>OPEN, D=>
      nx410, CLK=>nx1317);
   ix411 : mux21_ni port map ( Y=>nx410, A0=>q_2_3_EXMPLR, A1=>q_1_3_EXMPLR, 
      S0=>nx1291);
   gen_regs_1_regi_reg_q_3 : dff port map ( Q=>q_1_3_EXMPLR, QB=>OPEN, D=>
      nx400, CLK=>nx1317);
   ix401 : mux21_ni port map ( Y=>nx400, A0=>q_1_3_EXMPLR, A1=>q_0_3_EXMPLR, 
      S0=>nx1291);
   reg0_reg_q_3 : dff port map ( Q=>q_0_3_EXMPLR, QB=>OPEN, D=>nx390, CLK=>
      nx1317);
   ix391 : mux21_ni port map ( Y=>nx390, A0=>q_0_3_EXMPLR, A1=>d(3), S0=>
      nx1291);
   gen_regs_4_regi_reg_q_4 : dff port map ( Q=>q_4_4_EXMPLR, QB=>OPEN, D=>
      nx480, CLK=>nx1319);
   ix481 : mux21_ni port map ( Y=>nx480, A0=>q_4_4_EXMPLR, A1=>q_3_4_EXMPLR, 
      S0=>nx1293);
   gen_regs_3_regi_reg_q_4 : dff port map ( Q=>q_3_4_EXMPLR, QB=>OPEN, D=>
      nx470, CLK=>nx1319);
   ix471 : mux21_ni port map ( Y=>nx470, A0=>q_3_4_EXMPLR, A1=>q_2_4_EXMPLR, 
      S0=>nx1293);
   gen_regs_2_regi_reg_q_4 : dff port map ( Q=>q_2_4_EXMPLR, QB=>OPEN, D=>
      nx460, CLK=>nx1319);
   ix461 : mux21_ni port map ( Y=>nx460, A0=>q_2_4_EXMPLR, A1=>q_1_4_EXMPLR, 
      S0=>nx1293);
   gen_regs_1_regi_reg_q_4 : dff port map ( Q=>q_1_4_EXMPLR, QB=>OPEN, D=>
      nx450, CLK=>nx1319);
   ix451 : mux21_ni port map ( Y=>nx450, A0=>q_1_4_EXMPLR, A1=>q_0_4_EXMPLR, 
      S0=>nx1293);
   reg0_reg_q_4 : dff port map ( Q=>q_0_4_EXMPLR, QB=>OPEN, D=>nx440, CLK=>
      nx1317);
   ix441 : mux21_ni port map ( Y=>nx440, A0=>q_0_4_EXMPLR, A1=>d(4), S0=>
      nx1291);
   gen_regs_4_regi_reg_q_5 : dff port map ( Q=>q_4_5_EXMPLR, QB=>OPEN, D=>
      nx530, CLK=>nx1321);
   ix531 : mux21_ni port map ( Y=>nx530, A0=>q_4_5_EXMPLR, A1=>q_3_5_EXMPLR, 
      S0=>nx1295);
   gen_regs_3_regi_reg_q_5 : dff port map ( Q=>q_3_5_EXMPLR, QB=>OPEN, D=>
      nx520, CLK=>nx1321);
   ix521 : mux21_ni port map ( Y=>nx520, A0=>q_3_5_EXMPLR, A1=>q_2_5_EXMPLR, 
      S0=>nx1295);
   gen_regs_2_regi_reg_q_5 : dff port map ( Q=>q_2_5_EXMPLR, QB=>OPEN, D=>
      nx510, CLK=>nx1319);
   ix511 : mux21_ni port map ( Y=>nx510, A0=>q_2_5_EXMPLR, A1=>q_1_5_EXMPLR, 
      S0=>nx1293);
   gen_regs_1_regi_reg_q_5 : dff port map ( Q=>q_1_5_EXMPLR, QB=>OPEN, D=>
      nx500, CLK=>nx1319);
   ix501 : mux21_ni port map ( Y=>nx500, A0=>q_1_5_EXMPLR, A1=>q_0_5_EXMPLR, 
      S0=>nx1293);
   reg0_reg_q_5 : dff port map ( Q=>q_0_5_EXMPLR, QB=>OPEN, D=>nx490, CLK=>
      nx1319);
   ix491 : mux21_ni port map ( Y=>nx490, A0=>q_0_5_EXMPLR, A1=>d(5), S0=>
      nx1293);
   gen_regs_4_regi_reg_q_6 : dff port map ( Q=>q_4_6_EXMPLR, QB=>OPEN, D=>
      nx580, CLK=>nx1321);
   ix581 : mux21_ni port map ( Y=>nx580, A0=>q_4_6_EXMPLR, A1=>q_3_6_EXMPLR, 
      S0=>nx1295);
   gen_regs_3_regi_reg_q_6 : dff port map ( Q=>q_3_6_EXMPLR, QB=>OPEN, D=>
      nx570, CLK=>nx1321);
   ix571 : mux21_ni port map ( Y=>nx570, A0=>q_3_6_EXMPLR, A1=>q_2_6_EXMPLR, 
      S0=>nx1295);
   gen_regs_2_regi_reg_q_6 : dff port map ( Q=>q_2_6_EXMPLR, QB=>OPEN, D=>
      nx560, CLK=>nx1321);
   ix561 : mux21_ni port map ( Y=>nx560, A0=>q_2_6_EXMPLR, A1=>q_1_6_EXMPLR, 
      S0=>nx1295);
   gen_regs_1_regi_reg_q_6 : dff port map ( Q=>q_1_6_EXMPLR, QB=>OPEN, D=>
      nx550, CLK=>nx1321);
   ix551 : mux21_ni port map ( Y=>nx550, A0=>q_1_6_EXMPLR, A1=>q_0_6_EXMPLR, 
      S0=>nx1295);
   reg0_reg_q_6 : dff port map ( Q=>q_0_6_EXMPLR, QB=>OPEN, D=>nx540, CLK=>
      nx1321);
   ix541 : mux21_ni port map ( Y=>nx540, A0=>q_0_6_EXMPLR, A1=>d(6), S0=>
      nx1295);
   gen_regs_4_regi_reg_q_7 : dff port map ( Q=>q_4_7_EXMPLR, QB=>OPEN, D=>
      nx630, CLK=>nx1323);
   ix631 : mux21_ni port map ( Y=>nx630, A0=>q_4_7_EXMPLR, A1=>q_3_7_EXMPLR, 
      S0=>nx1297);
   gen_regs_3_regi_reg_q_7 : dff port map ( Q=>q_3_7_EXMPLR, QB=>OPEN, D=>
      nx620, CLK=>nx1323);
   ix621 : mux21_ni port map ( Y=>nx620, A0=>q_3_7_EXMPLR, A1=>q_2_7_EXMPLR, 
      S0=>nx1297);
   gen_regs_2_regi_reg_q_7 : dff port map ( Q=>q_2_7_EXMPLR, QB=>OPEN, D=>
      nx610, CLK=>nx1323);
   ix611 : mux21_ni port map ( Y=>nx610, A0=>q_2_7_EXMPLR, A1=>q_1_7_EXMPLR, 
      S0=>nx1297);
   gen_regs_1_regi_reg_q_7 : dff port map ( Q=>q_1_7_EXMPLR, QB=>OPEN, D=>
      nx600, CLK=>nx1323);
   ix601 : mux21_ni port map ( Y=>nx600, A0=>q_1_7_EXMPLR, A1=>q_0_7_EXMPLR, 
      S0=>nx1297);
   reg0_reg_q_7 : dff port map ( Q=>q_0_7_EXMPLR, QB=>OPEN, D=>nx590, CLK=>
      nx1323);
   ix591 : mux21_ni port map ( Y=>nx590, A0=>q_0_7_EXMPLR, A1=>d(7), S0=>
      nx1297);
   gen_regs_4_regi_reg_q_8 : dff port map ( Q=>q_4_8_EXMPLR, QB=>OPEN, D=>
      nx680, CLK=>nx1325);
   ix681 : mux21_ni port map ( Y=>nx680, A0=>q_4_8_EXMPLR, A1=>q_3_8_EXMPLR, 
      S0=>nx1299);
   gen_regs_3_regi_reg_q_8 : dff port map ( Q=>q_3_8_EXMPLR, QB=>OPEN, D=>
      nx670, CLK=>nx1325);
   ix671 : mux21_ni port map ( Y=>nx670, A0=>q_3_8_EXMPLR, A1=>q_2_8_EXMPLR, 
      S0=>nx1299);
   gen_regs_2_regi_reg_q_8 : dff port map ( Q=>q_2_8_EXMPLR, QB=>OPEN, D=>
      nx660, CLK=>nx1325);
   ix661 : mux21_ni port map ( Y=>nx660, A0=>q_2_8_EXMPLR, A1=>q_1_8_EXMPLR, 
      S0=>nx1299);
   gen_regs_1_regi_reg_q_8 : dff port map ( Q=>q_1_8_EXMPLR, QB=>OPEN, D=>
      nx650, CLK=>nx1323);
   ix651 : mux21_ni port map ( Y=>nx650, A0=>q_1_8_EXMPLR, A1=>q_0_8_EXMPLR, 
      S0=>nx1297);
   reg0_reg_q_8 : dff port map ( Q=>q_0_8_EXMPLR, QB=>OPEN, D=>nx640, CLK=>
      nx1323);
   ix641 : mux21_ni port map ( Y=>nx640, A0=>q_0_8_EXMPLR, A1=>d(8), S0=>
      nx1297);
   gen_regs_4_regi_reg_q_9 : dff port map ( Q=>q_4_9_EXMPLR, QB=>OPEN, D=>
      nx730, CLK=>nx1327);
   ix731 : mux21_ni port map ( Y=>nx730, A0=>q_4_9_EXMPLR, A1=>q_3_9_EXMPLR, 
      S0=>nx1301);
   gen_regs_3_regi_reg_q_9 : dff port map ( Q=>q_3_9_EXMPLR, QB=>OPEN, D=>
      nx720, CLK=>nx1325);
   ix721 : mux21_ni port map ( Y=>nx720, A0=>q_3_9_EXMPLR, A1=>q_2_9_EXMPLR, 
      S0=>nx1299);
   gen_regs_2_regi_reg_q_9 : dff port map ( Q=>q_2_9_EXMPLR, QB=>OPEN, D=>
      nx710, CLK=>nx1325);
   ix711 : mux21_ni port map ( Y=>nx710, A0=>q_2_9_EXMPLR, A1=>q_1_9_EXMPLR, 
      S0=>nx1299);
   gen_regs_1_regi_reg_q_9 : dff port map ( Q=>q_1_9_EXMPLR, QB=>OPEN, D=>
      nx700, CLK=>nx1325);
   ix701 : mux21_ni port map ( Y=>nx700, A0=>q_1_9_EXMPLR, A1=>q_0_9_EXMPLR, 
      S0=>nx1299);
   reg0_reg_q_9 : dff port map ( Q=>q_0_9_EXMPLR, QB=>OPEN, D=>nx690, CLK=>
      nx1325);
   ix691 : mux21_ni port map ( Y=>nx690, A0=>q_0_9_EXMPLR, A1=>d(9), S0=>
      nx1299);
   gen_regs_4_regi_reg_q_10 : dff port map ( Q=>q_4_10_EXMPLR, QB=>OPEN, D=>
      nx780, CLK=>nx1327);
   ix781 : mux21_ni port map ( Y=>nx780, A0=>q_4_10_EXMPLR, A1=>
      q_3_10_EXMPLR, S0=>nx1301);
   gen_regs_3_regi_reg_q_10 : dff port map ( Q=>q_3_10_EXMPLR, QB=>OPEN, D=>
      nx770, CLK=>nx1327);
   ix771 : mux21_ni port map ( Y=>nx770, A0=>q_3_10_EXMPLR, A1=>
      q_2_10_EXMPLR, S0=>nx1301);
   gen_regs_2_regi_reg_q_10 : dff port map ( Q=>q_2_10_EXMPLR, QB=>OPEN, D=>
      nx760, CLK=>nx1327);
   ix761 : mux21_ni port map ( Y=>nx760, A0=>q_2_10_EXMPLR, A1=>
      q_1_10_EXMPLR, S0=>nx1301);
   gen_regs_1_regi_reg_q_10 : dff port map ( Q=>q_1_10_EXMPLR, QB=>OPEN, D=>
      nx750, CLK=>nx1327);
   ix751 : mux21_ni port map ( Y=>nx750, A0=>q_1_10_EXMPLR, A1=>
      q_0_10_EXMPLR, S0=>nx1301);
   reg0_reg_q_10 : dff port map ( Q=>q_0_10_EXMPLR, QB=>OPEN, D=>nx740, CLK
      =>nx1327);
   ix741 : mux21_ni port map ( Y=>nx740, A0=>q_0_10_EXMPLR, A1=>d(10), S0=>
      nx1301);
   gen_regs_4_regi_reg_q_11 : dff port map ( Q=>q_4_11_EXMPLR, QB=>OPEN, D=>
      nx830, CLK=>nx1329);
   ix831 : mux21_ni port map ( Y=>nx830, A0=>q_4_11_EXMPLR, A1=>
      q_3_11_EXMPLR, S0=>nx1303);
   gen_regs_3_regi_reg_q_11 : dff port map ( Q=>q_3_11_EXMPLR, QB=>OPEN, D=>
      nx820, CLK=>nx1329);
   ix821 : mux21_ni port map ( Y=>nx820, A0=>q_3_11_EXMPLR, A1=>
      q_2_11_EXMPLR, S0=>nx1303);
   gen_regs_2_regi_reg_q_11 : dff port map ( Q=>q_2_11_EXMPLR, QB=>OPEN, D=>
      nx810, CLK=>nx1329);
   ix811 : mux21_ni port map ( Y=>nx810, A0=>q_2_11_EXMPLR, A1=>
      q_1_11_EXMPLR, S0=>nx1303);
   gen_regs_1_regi_reg_q_11 : dff port map ( Q=>q_1_11_EXMPLR, QB=>OPEN, D=>
      nx800, CLK=>nx1329);
   ix801 : mux21_ni port map ( Y=>nx800, A0=>q_1_11_EXMPLR, A1=>
      q_0_11_EXMPLR, S0=>nx1303);
   reg0_reg_q_11 : dff port map ( Q=>q_0_11_EXMPLR, QB=>OPEN, D=>nx790, CLK
      =>nx1327);
   ix791 : mux21_ni port map ( Y=>nx790, A0=>q_0_11_EXMPLR, A1=>d(11), S0=>
      nx1301);
   gen_regs_4_regi_reg_q_12 : dff port map ( Q=>q_4_12_EXMPLR, QB=>OPEN, D=>
      nx880, CLK=>nx1331);
   ix881 : mux21_ni port map ( Y=>nx880, A0=>q_4_12_EXMPLR, A1=>
      q_3_12_EXMPLR, S0=>nx1305);
   gen_regs_3_regi_reg_q_12 : dff port map ( Q=>q_3_12_EXMPLR, QB=>OPEN, D=>
      nx870, CLK=>nx1331);
   ix871 : mux21_ni port map ( Y=>nx870, A0=>q_3_12_EXMPLR, A1=>
      q_2_12_EXMPLR, S0=>nx1305);
   gen_regs_2_regi_reg_q_12 : dff port map ( Q=>q_2_12_EXMPLR, QB=>OPEN, D=>
      nx860, CLK=>nx1329);
   ix861 : mux21_ni port map ( Y=>nx860, A0=>q_2_12_EXMPLR, A1=>
      q_1_12_EXMPLR, S0=>nx1303);
   gen_regs_1_regi_reg_q_12 : dff port map ( Q=>q_1_12_EXMPLR, QB=>OPEN, D=>
      nx850, CLK=>nx1329);
   ix851 : mux21_ni port map ( Y=>nx850, A0=>q_1_12_EXMPLR, A1=>
      q_0_12_EXMPLR, S0=>nx1303);
   reg0_reg_q_12 : dff port map ( Q=>q_0_12_EXMPLR, QB=>OPEN, D=>nx840, CLK
      =>nx1329);
   ix841 : mux21_ni port map ( Y=>nx840, A0=>q_0_12_EXMPLR, A1=>d(12), S0=>
      nx1303);
   gen_regs_4_regi_reg_q_13 : dff port map ( Q=>q_4_13_EXMPLR, QB=>OPEN, D=>
      nx930, CLK=>nx1331);
   ix931 : mux21_ni port map ( Y=>nx930, A0=>q_4_13_EXMPLR, A1=>
      q_3_13_EXMPLR, S0=>nx1305);
   gen_regs_3_regi_reg_q_13 : dff port map ( Q=>q_3_13_EXMPLR, QB=>OPEN, D=>
      nx920, CLK=>nx1331);
   ix921 : mux21_ni port map ( Y=>nx920, A0=>q_3_13_EXMPLR, A1=>
      q_2_13_EXMPLR, S0=>nx1305);
   gen_regs_2_regi_reg_q_13 : dff port map ( Q=>q_2_13_EXMPLR, QB=>OPEN, D=>
      nx910, CLK=>nx1331);
   ix911 : mux21_ni port map ( Y=>nx910, A0=>q_2_13_EXMPLR, A1=>
      q_1_13_EXMPLR, S0=>nx1305);
   gen_regs_1_regi_reg_q_13 : dff port map ( Q=>q_1_13_EXMPLR, QB=>OPEN, D=>
      nx900, CLK=>nx1331);
   ix901 : mux21_ni port map ( Y=>nx900, A0=>q_1_13_EXMPLR, A1=>
      q_0_13_EXMPLR, S0=>nx1305);
   reg0_reg_q_13 : dff port map ( Q=>q_0_13_EXMPLR, QB=>OPEN, D=>nx890, CLK
      =>nx1331);
   ix891 : mux21_ni port map ( Y=>nx890, A0=>q_0_13_EXMPLR, A1=>d(13), S0=>
      nx1305);
   gen_regs_4_regi_reg_q_14 : dff port map ( Q=>q_4_14_EXMPLR, QB=>OPEN, D=>
      nx980, CLK=>nx1333);
   ix981 : mux21_ni port map ( Y=>nx980, A0=>q_4_14_EXMPLR, A1=>
      q_3_14_EXMPLR, S0=>nx1307);
   gen_regs_3_regi_reg_q_14 : dff port map ( Q=>q_3_14_EXMPLR, QB=>OPEN, D=>
      nx970, CLK=>nx1333);
   ix971 : mux21_ni port map ( Y=>nx970, A0=>q_3_14_EXMPLR, A1=>
      q_2_14_EXMPLR, S0=>nx1307);
   gen_regs_2_regi_reg_q_14 : dff port map ( Q=>q_2_14_EXMPLR, QB=>OPEN, D=>
      nx960, CLK=>nx1333);
   ix961 : mux21_ni port map ( Y=>nx960, A0=>q_2_14_EXMPLR, A1=>
      q_1_14_EXMPLR, S0=>nx1307);
   gen_regs_1_regi_reg_q_14 : dff port map ( Q=>q_1_14_EXMPLR, QB=>OPEN, D=>
      nx950, CLK=>nx1333);
   ix951 : mux21_ni port map ( Y=>nx950, A0=>q_1_14_EXMPLR, A1=>
      q_0_14_EXMPLR, S0=>nx1307);
   reg0_reg_q_14 : dff port map ( Q=>q_0_14_EXMPLR, QB=>OPEN, D=>nx940, CLK
      =>nx1333);
   ix941 : mux21_ni port map ( Y=>nx940, A0=>q_0_14_EXMPLR, A1=>d(14), S0=>
      nx1307);
   gen_regs_4_regi_reg_q_15 : dff port map ( Q=>q_4_15_EXMPLR, QB=>OPEN, D=>
      nx1030, CLK=>nx1335);
   ix1031 : mux21_ni port map ( Y=>nx1030, A0=>q_4_15_EXMPLR, A1=>
      q_3_15_EXMPLR, S0=>nx1309);
   gen_regs_3_regi_reg_q_15 : dff port map ( Q=>q_3_15_EXMPLR, QB=>OPEN, D=>
      nx1020, CLK=>nx1335);
   ix1021 : mux21_ni port map ( Y=>nx1020, A0=>q_3_15_EXMPLR, A1=>
      q_2_15_EXMPLR, S0=>nx1309);
   gen_regs_2_regi_reg_q_15 : dff port map ( Q=>q_2_15_EXMPLR, QB=>OPEN, D=>
      nx1010, CLK=>nx1335);
   ix1011 : mux21_ni port map ( Y=>nx1010, A0=>q_2_15_EXMPLR, A1=>
      q_1_15_EXMPLR, S0=>nx1309);
   gen_regs_1_regi_reg_q_15 : dff port map ( Q=>q_1_15_EXMPLR, QB=>OPEN, D=>
      nx1000, CLK=>nx1333);
   ix1001 : mux21_ni port map ( Y=>nx1000, A0=>q_1_15_EXMPLR, A1=>
      q_0_15_EXMPLR, S0=>nx1307);
   reg0_reg_q_15 : dff port map ( Q=>q_0_15_EXMPLR, QB=>OPEN, D=>nx990, CLK
      =>nx1333);
   ix991 : mux21_ni port map ( Y=>nx990, A0=>q_0_15_EXMPLR, A1=>d(15), S0=>
      nx1307);
   ix1286 : inv02 port map ( Y=>nx1287, A=>nx1337);
   ix1288 : inv02 port map ( Y=>nx1289, A=>nx1337);
   ix1290 : inv02 port map ( Y=>nx1291, A=>nx1337);
   ix1292 : inv02 port map ( Y=>nx1293, A=>nx1337);
   ix1294 : inv02 port map ( Y=>nx1295, A=>nx1337);
   ix1296 : inv02 port map ( Y=>nx1297, A=>nx1337);
   ix1298 : inv02 port map ( Y=>nx1299, A=>nx1337);
   ix1300 : inv02 port map ( Y=>nx1301, A=>nx1339);
   ix1302 : inv02 port map ( Y=>nx1303, A=>nx1339);
   ix1304 : inv02 port map ( Y=>nx1305, A=>nx1339);
   ix1306 : inv02 port map ( Y=>nx1307, A=>nx1339);
   ix1308 : inv02 port map ( Y=>nx1309, A=>nx1339);
   ix1312 : inv02 port map ( Y=>nx1313, A=>nx1341);
   ix1314 : inv02 port map ( Y=>nx1315, A=>nx1341);
   ix1316 : inv02 port map ( Y=>nx1317, A=>nx1341);
   ix1318 : inv02 port map ( Y=>nx1319, A=>nx1341);
   ix1320 : inv02 port map ( Y=>nx1321, A=>nx1341);
   ix1322 : inv02 port map ( Y=>nx1323, A=>nx1341);
   ix1324 : inv02 port map ( Y=>nx1325, A=>nx1341);
   ix1326 : inv02 port map ( Y=>nx1327, A=>nx1343);
   ix1328 : inv02 port map ( Y=>nx1329, A=>nx1343);
   ix1330 : inv02 port map ( Y=>nx1331, A=>nx1343);
   ix1332 : inv02 port map ( Y=>nx1333, A=>nx1343);
   ix1334 : inv02 port map ( Y=>nx1335, A=>nx1343);
   ix1336 : inv02 port map ( Y=>nx1337, A=>load);
   ix1338 : inv02 port map ( Y=>nx1339, A=>load);
   ix1340 : inv02 port map ( Y=>nx1341, A=>clk);
   ix1342 : inv02 port map ( Y=>nx1343, A=>clk);
end Structural_unfold_3007 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Queue_25 is
   port (
      d : IN std_logic_vector (15 DOWNTO 0) ;
      q_0_15 : OUT std_logic ;
      q_0_14 : OUT std_logic ;
      q_0_13 : OUT std_logic ;
      q_0_12 : OUT std_logic ;
      q_0_11 : OUT std_logic ;
      q_0_10 : OUT std_logic ;
      q_0_9 : OUT std_logic ;
      q_0_8 : OUT std_logic ;
      q_0_7 : OUT std_logic ;
      q_0_6 : OUT std_logic ;
      q_0_5 : OUT std_logic ;
      q_0_4 : OUT std_logic ;
      q_0_3 : OUT std_logic ;
      q_0_2 : OUT std_logic ;
      q_0_1 : OUT std_logic ;
      q_0_0 : OUT std_logic ;
      q_1_15 : OUT std_logic ;
      q_1_14 : OUT std_logic ;
      q_1_13 : OUT std_logic ;
      q_1_12 : OUT std_logic ;
      q_1_11 : OUT std_logic ;
      q_1_10 : OUT std_logic ;
      q_1_9 : OUT std_logic ;
      q_1_8 : OUT std_logic ;
      q_1_7 : OUT std_logic ;
      q_1_6 : OUT std_logic ;
      q_1_5 : OUT std_logic ;
      q_1_4 : OUT std_logic ;
      q_1_3 : OUT std_logic ;
      q_1_2 : OUT std_logic ;
      q_1_1 : OUT std_logic ;
      q_1_0 : OUT std_logic ;
      q_2_15 : OUT std_logic ;
      q_2_14 : OUT std_logic ;
      q_2_13 : OUT std_logic ;
      q_2_12 : OUT std_logic ;
      q_2_11 : OUT std_logic ;
      q_2_10 : OUT std_logic ;
      q_2_9 : OUT std_logic ;
      q_2_8 : OUT std_logic ;
      q_2_7 : OUT std_logic ;
      q_2_6 : OUT std_logic ;
      q_2_5 : OUT std_logic ;
      q_2_4 : OUT std_logic ;
      q_2_3 : OUT std_logic ;
      q_2_2 : OUT std_logic ;
      q_2_1 : OUT std_logic ;
      q_2_0 : OUT std_logic ;
      q_3_15 : OUT std_logic ;
      q_3_14 : OUT std_logic ;
      q_3_13 : OUT std_logic ;
      q_3_12 : OUT std_logic ;
      q_3_11 : OUT std_logic ;
      q_3_10 : OUT std_logic ;
      q_3_9 : OUT std_logic ;
      q_3_8 : OUT std_logic ;
      q_3_7 : OUT std_logic ;
      q_3_6 : OUT std_logic ;
      q_3_5 : OUT std_logic ;
      q_3_4 : OUT std_logic ;
      q_3_3 : OUT std_logic ;
      q_3_2 : OUT std_logic ;
      q_3_1 : OUT std_logic ;
      q_3_0 : OUT std_logic ;
      q_4_15 : OUT std_logic ;
      q_4_14 : OUT std_logic ;
      q_4_13 : OUT std_logic ;
      q_4_12 : OUT std_logic ;
      q_4_11 : OUT std_logic ;
      q_4_10 : OUT std_logic ;
      q_4_9 : OUT std_logic ;
      q_4_8 : OUT std_logic ;
      q_4_7 : OUT std_logic ;
      q_4_6 : OUT std_logic ;
      q_4_5 : OUT std_logic ;
      q_4_4 : OUT std_logic ;
      q_4_3 : OUT std_logic ;
      q_4_2 : OUT std_logic ;
      q_4_1 : OUT std_logic ;
      q_4_0 : OUT std_logic ;
      q_5_15 : OUT std_logic ;
      q_5_14 : OUT std_logic ;
      q_5_13 : OUT std_logic ;
      q_5_12 : OUT std_logic ;
      q_5_11 : OUT std_logic ;
      q_5_10 : OUT std_logic ;
      q_5_9 : OUT std_logic ;
      q_5_8 : OUT std_logic ;
      q_5_7 : OUT std_logic ;
      q_5_6 : OUT std_logic ;
      q_5_5 : OUT std_logic ;
      q_5_4 : OUT std_logic ;
      q_5_3 : OUT std_logic ;
      q_5_2 : OUT std_logic ;
      q_5_1 : OUT std_logic ;
      q_5_0 : OUT std_logic ;
      q_6_15 : OUT std_logic ;
      q_6_14 : OUT std_logic ;
      q_6_13 : OUT std_logic ;
      q_6_12 : OUT std_logic ;
      q_6_11 : OUT std_logic ;
      q_6_10 : OUT std_logic ;
      q_6_9 : OUT std_logic ;
      q_6_8 : OUT std_logic ;
      q_6_7 : OUT std_logic ;
      q_6_6 : OUT std_logic ;
      q_6_5 : OUT std_logic ;
      q_6_4 : OUT std_logic ;
      q_6_3 : OUT std_logic ;
      q_6_2 : OUT std_logic ;
      q_6_1 : OUT std_logic ;
      q_6_0 : OUT std_logic ;
      q_7_15 : OUT std_logic ;
      q_7_14 : OUT std_logic ;
      q_7_13 : OUT std_logic ;
      q_7_12 : OUT std_logic ;
      q_7_11 : OUT std_logic ;
      q_7_10 : OUT std_logic ;
      q_7_9 : OUT std_logic ;
      q_7_8 : OUT std_logic ;
      q_7_7 : OUT std_logic ;
      q_7_6 : OUT std_logic ;
      q_7_5 : OUT std_logic ;
      q_7_4 : OUT std_logic ;
      q_7_3 : OUT std_logic ;
      q_7_2 : OUT std_logic ;
      q_7_1 : OUT std_logic ;
      q_7_0 : OUT std_logic ;
      q_8_15 : OUT std_logic ;
      q_8_14 : OUT std_logic ;
      q_8_13 : OUT std_logic ;
      q_8_12 : OUT std_logic ;
      q_8_11 : OUT std_logic ;
      q_8_10 : OUT std_logic ;
      q_8_9 : OUT std_logic ;
      q_8_8 : OUT std_logic ;
      q_8_7 : OUT std_logic ;
      q_8_6 : OUT std_logic ;
      q_8_5 : OUT std_logic ;
      q_8_4 : OUT std_logic ;
      q_8_3 : OUT std_logic ;
      q_8_2 : OUT std_logic ;
      q_8_1 : OUT std_logic ;
      q_8_0 : OUT std_logic ;
      q_9_15 : OUT std_logic ;
      q_9_14 : OUT std_logic ;
      q_9_13 : OUT std_logic ;
      q_9_12 : OUT std_logic ;
      q_9_11 : OUT std_logic ;
      q_9_10 : OUT std_logic ;
      q_9_9 : OUT std_logic ;
      q_9_8 : OUT std_logic ;
      q_9_7 : OUT std_logic ;
      q_9_6 : OUT std_logic ;
      q_9_5 : OUT std_logic ;
      q_9_4 : OUT std_logic ;
      q_9_3 : OUT std_logic ;
      q_9_2 : OUT std_logic ;
      q_9_1 : OUT std_logic ;
      q_9_0 : OUT std_logic ;
      q_10_15 : OUT std_logic ;
      q_10_14 : OUT std_logic ;
      q_10_13 : OUT std_logic ;
      q_10_12 : OUT std_logic ;
      q_10_11 : OUT std_logic ;
      q_10_10 : OUT std_logic ;
      q_10_9 : OUT std_logic ;
      q_10_8 : OUT std_logic ;
      q_10_7 : OUT std_logic ;
      q_10_6 : OUT std_logic ;
      q_10_5 : OUT std_logic ;
      q_10_4 : OUT std_logic ;
      q_10_3 : OUT std_logic ;
      q_10_2 : OUT std_logic ;
      q_10_1 : OUT std_logic ;
      q_10_0 : OUT std_logic ;
      q_11_15 : OUT std_logic ;
      q_11_14 : OUT std_logic ;
      q_11_13 : OUT std_logic ;
      q_11_12 : OUT std_logic ;
      q_11_11 : OUT std_logic ;
      q_11_10 : OUT std_logic ;
      q_11_9 : OUT std_logic ;
      q_11_8 : OUT std_logic ;
      q_11_7 : OUT std_logic ;
      q_11_6 : OUT std_logic ;
      q_11_5 : OUT std_logic ;
      q_11_4 : OUT std_logic ;
      q_11_3 : OUT std_logic ;
      q_11_2 : OUT std_logic ;
      q_11_1 : OUT std_logic ;
      q_11_0 : OUT std_logic ;
      q_12_15 : OUT std_logic ;
      q_12_14 : OUT std_logic ;
      q_12_13 : OUT std_logic ;
      q_12_12 : OUT std_logic ;
      q_12_11 : OUT std_logic ;
      q_12_10 : OUT std_logic ;
      q_12_9 : OUT std_logic ;
      q_12_8 : OUT std_logic ;
      q_12_7 : OUT std_logic ;
      q_12_6 : OUT std_logic ;
      q_12_5 : OUT std_logic ;
      q_12_4 : OUT std_logic ;
      q_12_3 : OUT std_logic ;
      q_12_2 : OUT std_logic ;
      q_12_1 : OUT std_logic ;
      q_12_0 : OUT std_logic ;
      q_13_15 : OUT std_logic ;
      q_13_14 : OUT std_logic ;
      q_13_13 : OUT std_logic ;
      q_13_12 : OUT std_logic ;
      q_13_11 : OUT std_logic ;
      q_13_10 : OUT std_logic ;
      q_13_9 : OUT std_logic ;
      q_13_8 : OUT std_logic ;
      q_13_7 : OUT std_logic ;
      q_13_6 : OUT std_logic ;
      q_13_5 : OUT std_logic ;
      q_13_4 : OUT std_logic ;
      q_13_3 : OUT std_logic ;
      q_13_2 : OUT std_logic ;
      q_13_1 : OUT std_logic ;
      q_13_0 : OUT std_logic ;
      q_14_15 : OUT std_logic ;
      q_14_14 : OUT std_logic ;
      q_14_13 : OUT std_logic ;
      q_14_12 : OUT std_logic ;
      q_14_11 : OUT std_logic ;
      q_14_10 : OUT std_logic ;
      q_14_9 : OUT std_logic ;
      q_14_8 : OUT std_logic ;
      q_14_7 : OUT std_logic ;
      q_14_6 : OUT std_logic ;
      q_14_5 : OUT std_logic ;
      q_14_4 : OUT std_logic ;
      q_14_3 : OUT std_logic ;
      q_14_2 : OUT std_logic ;
      q_14_1 : OUT std_logic ;
      q_14_0 : OUT std_logic ;
      q_15_15 : OUT std_logic ;
      q_15_14 : OUT std_logic ;
      q_15_13 : OUT std_logic ;
      q_15_12 : OUT std_logic ;
      q_15_11 : OUT std_logic ;
      q_15_10 : OUT std_logic ;
      q_15_9 : OUT std_logic ;
      q_15_8 : OUT std_logic ;
      q_15_7 : OUT std_logic ;
      q_15_6 : OUT std_logic ;
      q_15_5 : OUT std_logic ;
      q_15_4 : OUT std_logic ;
      q_15_3 : OUT std_logic ;
      q_15_2 : OUT std_logic ;
      q_15_1 : OUT std_logic ;
      q_15_0 : OUT std_logic ;
      q_16_15 : OUT std_logic ;
      q_16_14 : OUT std_logic ;
      q_16_13 : OUT std_logic ;
      q_16_12 : OUT std_logic ;
      q_16_11 : OUT std_logic ;
      q_16_10 : OUT std_logic ;
      q_16_9 : OUT std_logic ;
      q_16_8 : OUT std_logic ;
      q_16_7 : OUT std_logic ;
      q_16_6 : OUT std_logic ;
      q_16_5 : OUT std_logic ;
      q_16_4 : OUT std_logic ;
      q_16_3 : OUT std_logic ;
      q_16_2 : OUT std_logic ;
      q_16_1 : OUT std_logic ;
      q_16_0 : OUT std_logic ;
      q_17_15 : OUT std_logic ;
      q_17_14 : OUT std_logic ;
      q_17_13 : OUT std_logic ;
      q_17_12 : OUT std_logic ;
      q_17_11 : OUT std_logic ;
      q_17_10 : OUT std_logic ;
      q_17_9 : OUT std_logic ;
      q_17_8 : OUT std_logic ;
      q_17_7 : OUT std_logic ;
      q_17_6 : OUT std_logic ;
      q_17_5 : OUT std_logic ;
      q_17_4 : OUT std_logic ;
      q_17_3 : OUT std_logic ;
      q_17_2 : OUT std_logic ;
      q_17_1 : OUT std_logic ;
      q_17_0 : OUT std_logic ;
      q_18_15 : OUT std_logic ;
      q_18_14 : OUT std_logic ;
      q_18_13 : OUT std_logic ;
      q_18_12 : OUT std_logic ;
      q_18_11 : OUT std_logic ;
      q_18_10 : OUT std_logic ;
      q_18_9 : OUT std_logic ;
      q_18_8 : OUT std_logic ;
      q_18_7 : OUT std_logic ;
      q_18_6 : OUT std_logic ;
      q_18_5 : OUT std_logic ;
      q_18_4 : OUT std_logic ;
      q_18_3 : OUT std_logic ;
      q_18_2 : OUT std_logic ;
      q_18_1 : OUT std_logic ;
      q_18_0 : OUT std_logic ;
      q_19_15 : OUT std_logic ;
      q_19_14 : OUT std_logic ;
      q_19_13 : OUT std_logic ;
      q_19_12 : OUT std_logic ;
      q_19_11 : OUT std_logic ;
      q_19_10 : OUT std_logic ;
      q_19_9 : OUT std_logic ;
      q_19_8 : OUT std_logic ;
      q_19_7 : OUT std_logic ;
      q_19_6 : OUT std_logic ;
      q_19_5 : OUT std_logic ;
      q_19_4 : OUT std_logic ;
      q_19_3 : OUT std_logic ;
      q_19_2 : OUT std_logic ;
      q_19_1 : OUT std_logic ;
      q_19_0 : OUT std_logic ;
      q_20_15 : OUT std_logic ;
      q_20_14 : OUT std_logic ;
      q_20_13 : OUT std_logic ;
      q_20_12 : OUT std_logic ;
      q_20_11 : OUT std_logic ;
      q_20_10 : OUT std_logic ;
      q_20_9 : OUT std_logic ;
      q_20_8 : OUT std_logic ;
      q_20_7 : OUT std_logic ;
      q_20_6 : OUT std_logic ;
      q_20_5 : OUT std_logic ;
      q_20_4 : OUT std_logic ;
      q_20_3 : OUT std_logic ;
      q_20_2 : OUT std_logic ;
      q_20_1 : OUT std_logic ;
      q_20_0 : OUT std_logic ;
      q_21_15 : OUT std_logic ;
      q_21_14 : OUT std_logic ;
      q_21_13 : OUT std_logic ;
      q_21_12 : OUT std_logic ;
      q_21_11 : OUT std_logic ;
      q_21_10 : OUT std_logic ;
      q_21_9 : OUT std_logic ;
      q_21_8 : OUT std_logic ;
      q_21_7 : OUT std_logic ;
      q_21_6 : OUT std_logic ;
      q_21_5 : OUT std_logic ;
      q_21_4 : OUT std_logic ;
      q_21_3 : OUT std_logic ;
      q_21_2 : OUT std_logic ;
      q_21_1 : OUT std_logic ;
      q_21_0 : OUT std_logic ;
      q_22_15 : OUT std_logic ;
      q_22_14 : OUT std_logic ;
      q_22_13 : OUT std_logic ;
      q_22_12 : OUT std_logic ;
      q_22_11 : OUT std_logic ;
      q_22_10 : OUT std_logic ;
      q_22_9 : OUT std_logic ;
      q_22_8 : OUT std_logic ;
      q_22_7 : OUT std_logic ;
      q_22_6 : OUT std_logic ;
      q_22_5 : OUT std_logic ;
      q_22_4 : OUT std_logic ;
      q_22_3 : OUT std_logic ;
      q_22_2 : OUT std_logic ;
      q_22_1 : OUT std_logic ;
      q_22_0 : OUT std_logic ;
      q_23_15 : OUT std_logic ;
      q_23_14 : OUT std_logic ;
      q_23_13 : OUT std_logic ;
      q_23_12 : OUT std_logic ;
      q_23_11 : OUT std_logic ;
      q_23_10 : OUT std_logic ;
      q_23_9 : OUT std_logic ;
      q_23_8 : OUT std_logic ;
      q_23_7 : OUT std_logic ;
      q_23_6 : OUT std_logic ;
      q_23_5 : OUT std_logic ;
      q_23_4 : OUT std_logic ;
      q_23_3 : OUT std_logic ;
      q_23_2 : OUT std_logic ;
      q_23_1 : OUT std_logic ;
      q_23_0 : OUT std_logic ;
      q_24_15 : OUT std_logic ;
      q_24_14 : OUT std_logic ;
      q_24_13 : OUT std_logic ;
      q_24_12 : OUT std_logic ;
      q_24_11 : OUT std_logic ;
      q_24_10 : OUT std_logic ;
      q_24_9 : OUT std_logic ;
      q_24_8 : OUT std_logic ;
      q_24_7 : OUT std_logic ;
      q_24_6 : OUT std_logic ;
      q_24_5 : OUT std_logic ;
      q_24_4 : OUT std_logic ;
      q_24_3 : OUT std_logic ;
      q_24_2 : OUT std_logic ;
      q_24_1 : OUT std_logic ;
      q_24_0 : OUT std_logic ;
      clk : IN std_logic ;
      load : IN std_logic ;
      reset : IN std_logic) ;
end Queue_25 ;

architecture Structural of Queue_25 is
   signal q_0_15_EXMPLR, q_0_14_EXMPLR, q_0_13_EXMPLR, q_0_12_EXMPLR, 
      q_0_11_EXMPLR, q_0_10_EXMPLR, q_0_9_EXMPLR, q_0_8_EXMPLR, q_0_7_EXMPLR, 
      q_0_6_EXMPLR, q_0_5_EXMPLR, q_0_4_EXMPLR, q_0_3_EXMPLR, q_0_2_EXMPLR, 
      q_0_1_EXMPLR, q_0_0_EXMPLR, q_1_15_EXMPLR, q_1_14_EXMPLR, 
      q_1_13_EXMPLR, q_1_12_EXMPLR, q_1_11_EXMPLR, q_1_10_EXMPLR, 
      q_1_9_EXMPLR, q_1_8_EXMPLR, q_1_7_EXMPLR, q_1_6_EXMPLR, q_1_5_EXMPLR, 
      q_1_4_EXMPLR, q_1_3_EXMPLR, q_1_2_EXMPLR, q_1_1_EXMPLR, q_1_0_EXMPLR, 
      q_2_15_EXMPLR, q_2_14_EXMPLR, q_2_13_EXMPLR, q_2_12_EXMPLR, 
      q_2_11_EXMPLR, q_2_10_EXMPLR, q_2_9_EXMPLR, q_2_8_EXMPLR, q_2_7_EXMPLR, 
      q_2_6_EXMPLR, q_2_5_EXMPLR, q_2_4_EXMPLR, q_2_3_EXMPLR, q_2_2_EXMPLR, 
      q_2_1_EXMPLR, q_2_0_EXMPLR, q_3_15_EXMPLR, q_3_14_EXMPLR, 
      q_3_13_EXMPLR, q_3_12_EXMPLR, q_3_11_EXMPLR, q_3_10_EXMPLR, 
      q_3_9_EXMPLR, q_3_8_EXMPLR, q_3_7_EXMPLR, q_3_6_EXMPLR, q_3_5_EXMPLR, 
      q_3_4_EXMPLR, q_3_3_EXMPLR, q_3_2_EXMPLR, q_3_1_EXMPLR, q_3_0_EXMPLR, 
      q_4_15_EXMPLR, q_4_14_EXMPLR, q_4_13_EXMPLR, q_4_12_EXMPLR, 
      q_4_11_EXMPLR, q_4_10_EXMPLR, q_4_9_EXMPLR, q_4_8_EXMPLR, q_4_7_EXMPLR, 
      q_4_6_EXMPLR, q_4_5_EXMPLR, q_4_4_EXMPLR, q_4_3_EXMPLR, q_4_2_EXMPLR, 
      q_4_1_EXMPLR, q_4_0_EXMPLR, q_5_15_EXMPLR, q_5_14_EXMPLR, 
      q_5_13_EXMPLR, q_5_12_EXMPLR, q_5_11_EXMPLR, q_5_10_EXMPLR, 
      q_5_9_EXMPLR, q_5_8_EXMPLR, q_5_7_EXMPLR, q_5_6_EXMPLR, q_5_5_EXMPLR, 
      q_5_4_EXMPLR, q_5_3_EXMPLR, q_5_2_EXMPLR, q_5_1_EXMPLR, q_5_0_EXMPLR, 
      q_6_15_EXMPLR, q_6_14_EXMPLR, q_6_13_EXMPLR, q_6_12_EXMPLR, 
      q_6_11_EXMPLR, q_6_10_EXMPLR, q_6_9_EXMPLR, q_6_8_EXMPLR, q_6_7_EXMPLR, 
      q_6_6_EXMPLR, q_6_5_EXMPLR, q_6_4_EXMPLR, q_6_3_EXMPLR, q_6_2_EXMPLR, 
      q_6_1_EXMPLR, q_6_0_EXMPLR, q_7_15_EXMPLR, q_7_14_EXMPLR, 
      q_7_13_EXMPLR, q_7_12_EXMPLR, q_7_11_EXMPLR, q_7_10_EXMPLR, 
      q_7_9_EXMPLR, q_7_8_EXMPLR, q_7_7_EXMPLR, q_7_6_EXMPLR, q_7_5_EXMPLR, 
      q_7_4_EXMPLR, q_7_3_EXMPLR, q_7_2_EXMPLR, q_7_1_EXMPLR, q_7_0_EXMPLR, 
      q_8_15_EXMPLR, q_8_14_EXMPLR, q_8_13_EXMPLR, q_8_12_EXMPLR, 
      q_8_11_EXMPLR, q_8_10_EXMPLR, q_8_9_EXMPLR, q_8_8_EXMPLR, q_8_7_EXMPLR, 
      q_8_6_EXMPLR, q_8_5_EXMPLR, q_8_4_EXMPLR, q_8_3_EXMPLR, q_8_2_EXMPLR, 
      q_8_1_EXMPLR, q_8_0_EXMPLR, q_9_15_EXMPLR, q_9_14_EXMPLR, 
      q_9_13_EXMPLR, q_9_12_EXMPLR, q_9_11_EXMPLR, q_9_10_EXMPLR, 
      q_9_9_EXMPLR, q_9_8_EXMPLR, q_9_7_EXMPLR, q_9_6_EXMPLR, q_9_5_EXMPLR, 
      q_9_4_EXMPLR, q_9_3_EXMPLR, q_9_2_EXMPLR, q_9_1_EXMPLR, q_9_0_EXMPLR, 
      q_10_15_EXMPLR, q_10_14_EXMPLR, q_10_13_EXMPLR, q_10_12_EXMPLR, 
      q_10_11_EXMPLR, q_10_10_EXMPLR, q_10_9_EXMPLR, q_10_8_EXMPLR, 
      q_10_7_EXMPLR, q_10_6_EXMPLR, q_10_5_EXMPLR, q_10_4_EXMPLR, 
      q_10_3_EXMPLR, q_10_2_EXMPLR, q_10_1_EXMPLR, q_10_0_EXMPLR, 
      q_11_15_EXMPLR, q_11_14_EXMPLR, q_11_13_EXMPLR, q_11_12_EXMPLR, 
      q_11_11_EXMPLR, q_11_10_EXMPLR, q_11_9_EXMPLR, q_11_8_EXMPLR, 
      q_11_7_EXMPLR, q_11_6_EXMPLR, q_11_5_EXMPLR, q_11_4_EXMPLR, 
      q_11_3_EXMPLR, q_11_2_EXMPLR, q_11_1_EXMPLR, q_11_0_EXMPLR, 
      q_12_15_EXMPLR, q_12_14_EXMPLR, q_12_13_EXMPLR, q_12_12_EXMPLR, 
      q_12_11_EXMPLR, q_12_10_EXMPLR, q_12_9_EXMPLR, q_12_8_EXMPLR, 
      q_12_7_EXMPLR, q_12_6_EXMPLR, q_12_5_EXMPLR, q_12_4_EXMPLR, 
      q_12_3_EXMPLR, q_12_2_EXMPLR, q_12_1_EXMPLR, q_12_0_EXMPLR, 
      q_13_15_EXMPLR, q_13_14_EXMPLR, q_13_13_EXMPLR, q_13_12_EXMPLR, 
      q_13_11_EXMPLR, q_13_10_EXMPLR, q_13_9_EXMPLR, q_13_8_EXMPLR, 
      q_13_7_EXMPLR, q_13_6_EXMPLR, q_13_5_EXMPLR, q_13_4_EXMPLR, 
      q_13_3_EXMPLR, q_13_2_EXMPLR, q_13_1_EXMPLR, q_13_0_EXMPLR, 
      q_14_15_EXMPLR, q_14_14_EXMPLR, q_14_13_EXMPLR, q_14_12_EXMPLR, 
      q_14_11_EXMPLR, q_14_10_EXMPLR, q_14_9_EXMPLR, q_14_8_EXMPLR, 
      q_14_7_EXMPLR, q_14_6_EXMPLR, q_14_5_EXMPLR, q_14_4_EXMPLR, 
      q_14_3_EXMPLR, q_14_2_EXMPLR, q_14_1_EXMPLR, q_14_0_EXMPLR, 
      q_15_15_EXMPLR, q_15_14_EXMPLR, q_15_13_EXMPLR, q_15_12_EXMPLR, 
      q_15_11_EXMPLR, q_15_10_EXMPLR, q_15_9_EXMPLR, q_15_8_EXMPLR, 
      q_15_7_EXMPLR, q_15_6_EXMPLR, q_15_5_EXMPLR, q_15_4_EXMPLR, 
      q_15_3_EXMPLR, q_15_2_EXMPLR, q_15_1_EXMPLR, q_15_0_EXMPLR, 
      q_16_15_EXMPLR, q_16_14_EXMPLR, q_16_13_EXMPLR, q_16_12_EXMPLR, 
      q_16_11_EXMPLR, q_16_10_EXMPLR, q_16_9_EXMPLR, q_16_8_EXMPLR, 
      q_16_7_EXMPLR, q_16_6_EXMPLR, q_16_5_EXMPLR, q_16_4_EXMPLR, 
      q_16_3_EXMPLR, q_16_2_EXMPLR, q_16_1_EXMPLR, q_16_0_EXMPLR, 
      q_17_15_EXMPLR, q_17_14_EXMPLR, q_17_13_EXMPLR, q_17_12_EXMPLR, 
      q_17_11_EXMPLR, q_17_10_EXMPLR, q_17_9_EXMPLR, q_17_8_EXMPLR, 
      q_17_7_EXMPLR, q_17_6_EXMPLR, q_17_5_EXMPLR, q_17_4_EXMPLR, 
      q_17_3_EXMPLR, q_17_2_EXMPLR, q_17_1_EXMPLR, q_17_0_EXMPLR, 
      q_18_15_EXMPLR, q_18_14_EXMPLR, q_18_13_EXMPLR, q_18_12_EXMPLR, 
      q_18_11_EXMPLR, q_18_10_EXMPLR, q_18_9_EXMPLR, q_18_8_EXMPLR, 
      q_18_7_EXMPLR, q_18_6_EXMPLR, q_18_5_EXMPLR, q_18_4_EXMPLR, 
      q_18_3_EXMPLR, q_18_2_EXMPLR, q_18_1_EXMPLR, q_18_0_EXMPLR, 
      q_19_15_EXMPLR, q_19_14_EXMPLR, q_19_13_EXMPLR, q_19_12_EXMPLR, 
      q_19_11_EXMPLR, q_19_10_EXMPLR, q_19_9_EXMPLR, q_19_8_EXMPLR, 
      q_19_7_EXMPLR, q_19_6_EXMPLR, q_19_5_EXMPLR, q_19_4_EXMPLR, 
      q_19_3_EXMPLR, q_19_2_EXMPLR, q_19_1_EXMPLR, q_19_0_EXMPLR, 
      q_20_15_EXMPLR, q_20_14_EXMPLR, q_20_13_EXMPLR, q_20_12_EXMPLR, 
      q_20_11_EXMPLR, q_20_10_EXMPLR, q_20_9_EXMPLR, q_20_8_EXMPLR, 
      q_20_7_EXMPLR, q_20_6_EXMPLR, q_20_5_EXMPLR, q_20_4_EXMPLR, 
      q_20_3_EXMPLR, q_20_2_EXMPLR, q_20_1_EXMPLR, q_20_0_EXMPLR, 
      q_21_15_EXMPLR, q_21_14_EXMPLR, q_21_13_EXMPLR, q_21_12_EXMPLR, 
      q_21_11_EXMPLR, q_21_10_EXMPLR, q_21_9_EXMPLR, q_21_8_EXMPLR, 
      q_21_7_EXMPLR, q_21_6_EXMPLR, q_21_5_EXMPLR, q_21_4_EXMPLR, 
      q_21_3_EXMPLR, q_21_2_EXMPLR, q_21_1_EXMPLR, q_21_0_EXMPLR, 
      q_22_15_EXMPLR, q_22_14_EXMPLR, q_22_13_EXMPLR, q_22_12_EXMPLR, 
      q_22_11_EXMPLR, q_22_10_EXMPLR, q_22_9_EXMPLR, q_22_8_EXMPLR, 
      q_22_7_EXMPLR, q_22_6_EXMPLR, q_22_5_EXMPLR, q_22_4_EXMPLR, 
      q_22_3_EXMPLR, q_22_2_EXMPLR, q_22_1_EXMPLR, q_22_0_EXMPLR, 
      q_23_15_EXMPLR, q_23_14_EXMPLR, q_23_13_EXMPLR, q_23_12_EXMPLR, 
      q_23_11_EXMPLR, q_23_10_EXMPLR, q_23_9_EXMPLR, q_23_8_EXMPLR, 
      q_23_7_EXMPLR, q_23_6_EXMPLR, q_23_5_EXMPLR, q_23_4_EXMPLR, 
      q_23_3_EXMPLR, q_23_2_EXMPLR, q_23_1_EXMPLR, q_23_0_EXMPLR, 
      q_24_15_EXMPLR, q_24_14_EXMPLR, q_24_13_EXMPLR, q_24_12_EXMPLR, 
      q_24_11_EXMPLR, q_24_10_EXMPLR, q_24_9_EXMPLR, q_24_8_EXMPLR, 
      q_24_7_EXMPLR, q_24_6_EXMPLR, q_24_5_EXMPLR, q_24_4_EXMPLR, 
      q_24_3_EXMPLR, q_24_2_EXMPLR, q_24_1_EXMPLR, q_24_0_EXMPLR, nx1733, 
      nx1743, nx1753, nx1763, nx1773, nx1783, nx1793, nx1803, nx1813, nx1823, 
      nx1833, nx1843, nx1853, nx1863, nx1873, nx1883, nx1893, nx1903, nx1913, 
      nx1923, nx1933, nx1943, nx1953, nx1963, nx1973, nx1983, nx1993, nx2003, 
      nx2013, nx2023, nx2033, nx2043, nx2053, nx2063, nx2073, nx2083, nx2093, 
      nx2103, nx2113, nx2123, nx2133, nx2143, nx2153, nx2163, nx2173, nx2183, 
      nx2193, nx2203, nx2213, nx2223, nx2233, nx2243, nx2253, nx2263, nx2273, 
      nx2283, nx2293, nx2303, nx2313, nx2323, nx2333, nx2343, nx2353, nx2363, 
      nx2373, nx2383, nx2393, nx2403, nx2413, nx2423, nx2433, nx2443, nx2453, 
      nx2463, nx2473, nx2483, nx2493, nx2503, nx2513, nx2523, nx2533, nx2543, 
      nx2553, nx2563, nx2573, nx2583, nx2593, nx2603, nx2613, nx2623, nx2633, 
      nx2643, nx2653, nx2663, nx2673, nx2683, nx2693, nx2703, nx2713, nx2723, 
      nx2733, nx2743, nx2753, nx2763, nx2773, nx2783, nx2793, nx2803, nx2813, 
      nx2823, nx2833, nx2843, nx2853, nx2863, nx2873, nx2883, nx2893, nx2903, 
      nx2913, nx2923, nx2933, nx2943, nx2953, nx2963, nx2973, nx2983, nx2993, 
      nx3003, nx3013, nx3023, nx3033, nx3043, nx3053, nx3063, nx3073, nx3083, 
      nx3093, nx3103, nx3113, nx3123, nx3133, nx3143, nx3153, nx3163, nx3173, 
      nx3183, nx3193, nx3203, nx3213, nx3223, nx3233, nx3243, nx3253, nx3263, 
      nx3273, nx3283, nx3293, nx3303, nx3313, nx3323, nx3333, nx3343, nx3353, 
      nx3363, nx3373, nx3383, nx3393, nx3403, nx3413, nx3423, nx3433, nx3443, 
      nx3453, nx3463, nx3473, nx3483, nx3493, nx3503, nx3513, nx3523, nx3533, 
      nx3543, nx3553, nx3563, nx3573, nx3583, nx3593, nx3603, nx3613, nx3623, 
      nx3633, nx3643, nx3653, nx3663, nx3673, nx3683, nx3693, nx3703, nx3713, 
      nx3723, nx3733, nx3743, nx3753, nx3763, nx3773, nx3783, nx3793, nx3803, 
      nx3813, nx3823, nx3833, nx3843, nx3853, nx3863, nx3873, nx3883, nx3893, 
      nx3903, nx3913, nx3923, nx3933, nx3943, nx3953, nx3963, nx3973, nx3983, 
      nx3993, nx4003, nx4013, nx4023, nx4033, nx4043, nx4053, nx4063, nx4073, 
      nx4083, nx4093, nx4103, nx4113, nx4123, nx4133, nx4143, nx4153, nx4163, 
      nx4173, nx4183, nx4193, nx4203, nx4213, nx4223, nx4233, nx4243, nx4253, 
      nx4263, nx4273, nx4283, nx4293, nx4303, nx4313, nx4323, nx4333, nx4343, 
      nx4353, nx4363, nx4373, nx4383, nx4393, nx4403, nx4413, nx4423, nx4433, 
      nx4443, nx4453, nx4463, nx4473, nx4483, nx4493, nx4503, nx4513, nx4523, 
      nx4533, nx4543, nx4553, nx4563, nx4573, nx4583, nx4593, nx4603, nx4613, 
      nx4623, nx4633, nx4643, nx4653, nx4663, nx4673, nx4683, nx4693, nx4703, 
      nx4713, nx4723, nx4733, nx4743, nx4753, nx4763, nx4773, nx4783, nx4793, 
      nx4803, nx4813, nx4823, nx4833, nx4843, nx4853, nx4863, nx4873, nx4883, 
      nx4893, nx4903, nx4913, nx4923, nx4933, nx4943, nx4953, nx4963, nx4973, 
      nx4983, nx4993, nx5003, nx5013, nx5023, nx5033, nx5043, nx5053, nx5063, 
      nx5073, nx5083, nx5093, nx5103, nx5113, nx5123, nx5133, nx5143, nx5153, 
      nx5163, nx5173, nx5183, nx5193, nx5203, nx5213, nx5223, nx5233, nx5243, 
      nx5253, nx5263, nx5273, nx5283, nx5293, nx5303, nx5313, nx5323, nx5333, 
      nx5343, nx5353, nx5363, nx5373, nx5383, nx5393, nx5403, nx5413, nx5423, 
      nx5433, nx5443, nx5453, nx5463, nx5473, nx5483, nx5493, nx5503, nx5513, 
      nx5523, nx5533, nx5543, nx5553, nx5563, nx5573, nx5583, nx5593, nx5603, 
      nx5613, nx5623, nx5633, nx5643, nx5653, nx5663, nx5673, nx5683, nx5693, 
      nx5703, nx5713, nx5723, nx6940, nx6942, nx6944, nx6946, nx6948, nx6950, 
      nx6952, nx6954, nx6956, nx6958, nx6960, nx6962, nx6964, nx6966, nx6968, 
      nx6970, nx6972, nx6974, nx6976, nx6978, nx6980, nx6982, nx6984, nx6986, 
      nx6988, nx6990, nx6992, nx6994, nx6996, nx6998, nx7000, nx7002, nx7004, 
      nx7006, nx7008, nx7010, nx7012, nx7014, nx7016, nx7018, nx7020, nx7022, 
      nx7024, nx7026, nx7028, nx7030, nx7032, nx7034, nx7036, nx7038, nx7040, 
      nx7042, nx7044, nx7046, nx7048, nx7050, nx7052, nx7054, nx7058, nx7060, 
      nx7062, nx7064, nx7066, nx7068, nx7070, nx7072, nx7074, nx7076, nx7078, 
      nx7080, nx7082, nx7084, nx7086, nx7088, nx7090, nx7092, nx7094, nx7096, 
      nx7098, nx7100, nx7102, nx7104, nx7106, nx7108, nx7110, nx7112, nx7114, 
      nx7116, nx7118, nx7120, nx7122, nx7124, nx7126, nx7128, nx7130, nx7132, 
      nx7134, nx7136, nx7138, nx7140, nx7142, nx7144, nx7146, nx7148, nx7150, 
      nx7152, nx7154, nx7156, nx7158, nx7160, nx7162, nx7164, nx7166, nx7168, 
      nx7170, nx7172, nx7174, nx7176, nx7178, nx7180, nx7182, nx7184, nx7186, 
      nx7188, nx7190, nx7192, nx7194, nx7196, nx7198, nx7200, nx7202, nx7204, 
      nx7206, nx7208, nx7214, nx7216, nx7218, nx7220, nx7626, nx7628: 
   std_logic ;

begin
   q_0_15 <= q_0_15_EXMPLR ;
   q_0_14 <= q_0_14_EXMPLR ;
   q_0_13 <= q_0_13_EXMPLR ;
   q_0_12 <= q_0_12_EXMPLR ;
   q_0_11 <= q_0_11_EXMPLR ;
   q_0_10 <= q_0_10_EXMPLR ;
   q_0_9 <= q_0_9_EXMPLR ;
   q_0_8 <= q_0_8_EXMPLR ;
   q_0_7 <= q_0_7_EXMPLR ;
   q_0_6 <= q_0_6_EXMPLR ;
   q_0_5 <= q_0_5_EXMPLR ;
   q_0_4 <= q_0_4_EXMPLR ;
   q_0_3 <= q_0_3_EXMPLR ;
   q_0_2 <= q_0_2_EXMPLR ;
   q_0_1 <= q_0_1_EXMPLR ;
   q_0_0 <= q_0_0_EXMPLR ;
   q_1_15 <= q_1_15_EXMPLR ;
   q_1_14 <= q_1_14_EXMPLR ;
   q_1_13 <= q_1_13_EXMPLR ;
   q_1_12 <= q_1_12_EXMPLR ;
   q_1_11 <= q_1_11_EXMPLR ;
   q_1_10 <= q_1_10_EXMPLR ;
   q_1_9 <= q_1_9_EXMPLR ;
   q_1_8 <= q_1_8_EXMPLR ;
   q_1_7 <= q_1_7_EXMPLR ;
   q_1_6 <= q_1_6_EXMPLR ;
   q_1_5 <= q_1_5_EXMPLR ;
   q_1_4 <= q_1_4_EXMPLR ;
   q_1_3 <= q_1_3_EXMPLR ;
   q_1_2 <= q_1_2_EXMPLR ;
   q_1_1 <= q_1_1_EXMPLR ;
   q_1_0 <= q_1_0_EXMPLR ;
   q_2_15 <= q_2_15_EXMPLR ;
   q_2_14 <= q_2_14_EXMPLR ;
   q_2_13 <= q_2_13_EXMPLR ;
   q_2_12 <= q_2_12_EXMPLR ;
   q_2_11 <= q_2_11_EXMPLR ;
   q_2_10 <= q_2_10_EXMPLR ;
   q_2_9 <= q_2_9_EXMPLR ;
   q_2_8 <= q_2_8_EXMPLR ;
   q_2_7 <= q_2_7_EXMPLR ;
   q_2_6 <= q_2_6_EXMPLR ;
   q_2_5 <= q_2_5_EXMPLR ;
   q_2_4 <= q_2_4_EXMPLR ;
   q_2_3 <= q_2_3_EXMPLR ;
   q_2_2 <= q_2_2_EXMPLR ;
   q_2_1 <= q_2_1_EXMPLR ;
   q_2_0 <= q_2_0_EXMPLR ;
   q_3_15 <= q_3_15_EXMPLR ;
   q_3_14 <= q_3_14_EXMPLR ;
   q_3_13 <= q_3_13_EXMPLR ;
   q_3_12 <= q_3_12_EXMPLR ;
   q_3_11 <= q_3_11_EXMPLR ;
   q_3_10 <= q_3_10_EXMPLR ;
   q_3_9 <= q_3_9_EXMPLR ;
   q_3_8 <= q_3_8_EXMPLR ;
   q_3_7 <= q_3_7_EXMPLR ;
   q_3_6 <= q_3_6_EXMPLR ;
   q_3_5 <= q_3_5_EXMPLR ;
   q_3_4 <= q_3_4_EXMPLR ;
   q_3_3 <= q_3_3_EXMPLR ;
   q_3_2 <= q_3_2_EXMPLR ;
   q_3_1 <= q_3_1_EXMPLR ;
   q_3_0 <= q_3_0_EXMPLR ;
   q_4_15 <= q_4_15_EXMPLR ;
   q_4_14 <= q_4_14_EXMPLR ;
   q_4_13 <= q_4_13_EXMPLR ;
   q_4_12 <= q_4_12_EXMPLR ;
   q_4_11 <= q_4_11_EXMPLR ;
   q_4_10 <= q_4_10_EXMPLR ;
   q_4_9 <= q_4_9_EXMPLR ;
   q_4_8 <= q_4_8_EXMPLR ;
   q_4_7 <= q_4_7_EXMPLR ;
   q_4_6 <= q_4_6_EXMPLR ;
   q_4_5 <= q_4_5_EXMPLR ;
   q_4_4 <= q_4_4_EXMPLR ;
   q_4_3 <= q_4_3_EXMPLR ;
   q_4_2 <= q_4_2_EXMPLR ;
   q_4_1 <= q_4_1_EXMPLR ;
   q_4_0 <= q_4_0_EXMPLR ;
   q_5_15 <= q_5_15_EXMPLR ;
   q_5_14 <= q_5_14_EXMPLR ;
   q_5_13 <= q_5_13_EXMPLR ;
   q_5_12 <= q_5_12_EXMPLR ;
   q_5_11 <= q_5_11_EXMPLR ;
   q_5_10 <= q_5_10_EXMPLR ;
   q_5_9 <= q_5_9_EXMPLR ;
   q_5_8 <= q_5_8_EXMPLR ;
   q_5_7 <= q_5_7_EXMPLR ;
   q_5_6 <= q_5_6_EXMPLR ;
   q_5_5 <= q_5_5_EXMPLR ;
   q_5_4 <= q_5_4_EXMPLR ;
   q_5_3 <= q_5_3_EXMPLR ;
   q_5_2 <= q_5_2_EXMPLR ;
   q_5_1 <= q_5_1_EXMPLR ;
   q_5_0 <= q_5_0_EXMPLR ;
   q_6_15 <= q_6_15_EXMPLR ;
   q_6_14 <= q_6_14_EXMPLR ;
   q_6_13 <= q_6_13_EXMPLR ;
   q_6_12 <= q_6_12_EXMPLR ;
   q_6_11 <= q_6_11_EXMPLR ;
   q_6_10 <= q_6_10_EXMPLR ;
   q_6_9 <= q_6_9_EXMPLR ;
   q_6_8 <= q_6_8_EXMPLR ;
   q_6_7 <= q_6_7_EXMPLR ;
   q_6_6 <= q_6_6_EXMPLR ;
   q_6_5 <= q_6_5_EXMPLR ;
   q_6_4 <= q_6_4_EXMPLR ;
   q_6_3 <= q_6_3_EXMPLR ;
   q_6_2 <= q_6_2_EXMPLR ;
   q_6_1 <= q_6_1_EXMPLR ;
   q_6_0 <= q_6_0_EXMPLR ;
   q_7_15 <= q_7_15_EXMPLR ;
   q_7_14 <= q_7_14_EXMPLR ;
   q_7_13 <= q_7_13_EXMPLR ;
   q_7_12 <= q_7_12_EXMPLR ;
   q_7_11 <= q_7_11_EXMPLR ;
   q_7_10 <= q_7_10_EXMPLR ;
   q_7_9 <= q_7_9_EXMPLR ;
   q_7_8 <= q_7_8_EXMPLR ;
   q_7_7 <= q_7_7_EXMPLR ;
   q_7_6 <= q_7_6_EXMPLR ;
   q_7_5 <= q_7_5_EXMPLR ;
   q_7_4 <= q_7_4_EXMPLR ;
   q_7_3 <= q_7_3_EXMPLR ;
   q_7_2 <= q_7_2_EXMPLR ;
   q_7_1 <= q_7_1_EXMPLR ;
   q_7_0 <= q_7_0_EXMPLR ;
   q_8_15 <= q_8_15_EXMPLR ;
   q_8_14 <= q_8_14_EXMPLR ;
   q_8_13 <= q_8_13_EXMPLR ;
   q_8_12 <= q_8_12_EXMPLR ;
   q_8_11 <= q_8_11_EXMPLR ;
   q_8_10 <= q_8_10_EXMPLR ;
   q_8_9 <= q_8_9_EXMPLR ;
   q_8_8 <= q_8_8_EXMPLR ;
   q_8_7 <= q_8_7_EXMPLR ;
   q_8_6 <= q_8_6_EXMPLR ;
   q_8_5 <= q_8_5_EXMPLR ;
   q_8_4 <= q_8_4_EXMPLR ;
   q_8_3 <= q_8_3_EXMPLR ;
   q_8_2 <= q_8_2_EXMPLR ;
   q_8_1 <= q_8_1_EXMPLR ;
   q_8_0 <= q_8_0_EXMPLR ;
   q_9_15 <= q_9_15_EXMPLR ;
   q_9_14 <= q_9_14_EXMPLR ;
   q_9_13 <= q_9_13_EXMPLR ;
   q_9_12 <= q_9_12_EXMPLR ;
   q_9_11 <= q_9_11_EXMPLR ;
   q_9_10 <= q_9_10_EXMPLR ;
   q_9_9 <= q_9_9_EXMPLR ;
   q_9_8 <= q_9_8_EXMPLR ;
   q_9_7 <= q_9_7_EXMPLR ;
   q_9_6 <= q_9_6_EXMPLR ;
   q_9_5 <= q_9_5_EXMPLR ;
   q_9_4 <= q_9_4_EXMPLR ;
   q_9_3 <= q_9_3_EXMPLR ;
   q_9_2 <= q_9_2_EXMPLR ;
   q_9_1 <= q_9_1_EXMPLR ;
   q_9_0 <= q_9_0_EXMPLR ;
   q_10_15 <= q_10_15_EXMPLR ;
   q_10_14 <= q_10_14_EXMPLR ;
   q_10_13 <= q_10_13_EXMPLR ;
   q_10_12 <= q_10_12_EXMPLR ;
   q_10_11 <= q_10_11_EXMPLR ;
   q_10_10 <= q_10_10_EXMPLR ;
   q_10_9 <= q_10_9_EXMPLR ;
   q_10_8 <= q_10_8_EXMPLR ;
   q_10_7 <= q_10_7_EXMPLR ;
   q_10_6 <= q_10_6_EXMPLR ;
   q_10_5 <= q_10_5_EXMPLR ;
   q_10_4 <= q_10_4_EXMPLR ;
   q_10_3 <= q_10_3_EXMPLR ;
   q_10_2 <= q_10_2_EXMPLR ;
   q_10_1 <= q_10_1_EXMPLR ;
   q_10_0 <= q_10_0_EXMPLR ;
   q_11_15 <= q_11_15_EXMPLR ;
   q_11_14 <= q_11_14_EXMPLR ;
   q_11_13 <= q_11_13_EXMPLR ;
   q_11_12 <= q_11_12_EXMPLR ;
   q_11_11 <= q_11_11_EXMPLR ;
   q_11_10 <= q_11_10_EXMPLR ;
   q_11_9 <= q_11_9_EXMPLR ;
   q_11_8 <= q_11_8_EXMPLR ;
   q_11_7 <= q_11_7_EXMPLR ;
   q_11_6 <= q_11_6_EXMPLR ;
   q_11_5 <= q_11_5_EXMPLR ;
   q_11_4 <= q_11_4_EXMPLR ;
   q_11_3 <= q_11_3_EXMPLR ;
   q_11_2 <= q_11_2_EXMPLR ;
   q_11_1 <= q_11_1_EXMPLR ;
   q_11_0 <= q_11_0_EXMPLR ;
   q_12_15 <= q_12_15_EXMPLR ;
   q_12_14 <= q_12_14_EXMPLR ;
   q_12_13 <= q_12_13_EXMPLR ;
   q_12_12 <= q_12_12_EXMPLR ;
   q_12_11 <= q_12_11_EXMPLR ;
   q_12_10 <= q_12_10_EXMPLR ;
   q_12_9 <= q_12_9_EXMPLR ;
   q_12_8 <= q_12_8_EXMPLR ;
   q_12_7 <= q_12_7_EXMPLR ;
   q_12_6 <= q_12_6_EXMPLR ;
   q_12_5 <= q_12_5_EXMPLR ;
   q_12_4 <= q_12_4_EXMPLR ;
   q_12_3 <= q_12_3_EXMPLR ;
   q_12_2 <= q_12_2_EXMPLR ;
   q_12_1 <= q_12_1_EXMPLR ;
   q_12_0 <= q_12_0_EXMPLR ;
   q_13_15 <= q_13_15_EXMPLR ;
   q_13_14 <= q_13_14_EXMPLR ;
   q_13_13 <= q_13_13_EXMPLR ;
   q_13_12 <= q_13_12_EXMPLR ;
   q_13_11 <= q_13_11_EXMPLR ;
   q_13_10 <= q_13_10_EXMPLR ;
   q_13_9 <= q_13_9_EXMPLR ;
   q_13_8 <= q_13_8_EXMPLR ;
   q_13_7 <= q_13_7_EXMPLR ;
   q_13_6 <= q_13_6_EXMPLR ;
   q_13_5 <= q_13_5_EXMPLR ;
   q_13_4 <= q_13_4_EXMPLR ;
   q_13_3 <= q_13_3_EXMPLR ;
   q_13_2 <= q_13_2_EXMPLR ;
   q_13_1 <= q_13_1_EXMPLR ;
   q_13_0 <= q_13_0_EXMPLR ;
   q_14_15 <= q_14_15_EXMPLR ;
   q_14_14 <= q_14_14_EXMPLR ;
   q_14_13 <= q_14_13_EXMPLR ;
   q_14_12 <= q_14_12_EXMPLR ;
   q_14_11 <= q_14_11_EXMPLR ;
   q_14_10 <= q_14_10_EXMPLR ;
   q_14_9 <= q_14_9_EXMPLR ;
   q_14_8 <= q_14_8_EXMPLR ;
   q_14_7 <= q_14_7_EXMPLR ;
   q_14_6 <= q_14_6_EXMPLR ;
   q_14_5 <= q_14_5_EXMPLR ;
   q_14_4 <= q_14_4_EXMPLR ;
   q_14_3 <= q_14_3_EXMPLR ;
   q_14_2 <= q_14_2_EXMPLR ;
   q_14_1 <= q_14_1_EXMPLR ;
   q_14_0 <= q_14_0_EXMPLR ;
   q_15_15 <= q_15_15_EXMPLR ;
   q_15_14 <= q_15_14_EXMPLR ;
   q_15_13 <= q_15_13_EXMPLR ;
   q_15_12 <= q_15_12_EXMPLR ;
   q_15_11 <= q_15_11_EXMPLR ;
   q_15_10 <= q_15_10_EXMPLR ;
   q_15_9 <= q_15_9_EXMPLR ;
   q_15_8 <= q_15_8_EXMPLR ;
   q_15_7 <= q_15_7_EXMPLR ;
   q_15_6 <= q_15_6_EXMPLR ;
   q_15_5 <= q_15_5_EXMPLR ;
   q_15_4 <= q_15_4_EXMPLR ;
   q_15_3 <= q_15_3_EXMPLR ;
   q_15_2 <= q_15_2_EXMPLR ;
   q_15_1 <= q_15_1_EXMPLR ;
   q_15_0 <= q_15_0_EXMPLR ;
   q_16_15 <= q_16_15_EXMPLR ;
   q_16_14 <= q_16_14_EXMPLR ;
   q_16_13 <= q_16_13_EXMPLR ;
   q_16_12 <= q_16_12_EXMPLR ;
   q_16_11 <= q_16_11_EXMPLR ;
   q_16_10 <= q_16_10_EXMPLR ;
   q_16_9 <= q_16_9_EXMPLR ;
   q_16_8 <= q_16_8_EXMPLR ;
   q_16_7 <= q_16_7_EXMPLR ;
   q_16_6 <= q_16_6_EXMPLR ;
   q_16_5 <= q_16_5_EXMPLR ;
   q_16_4 <= q_16_4_EXMPLR ;
   q_16_3 <= q_16_3_EXMPLR ;
   q_16_2 <= q_16_2_EXMPLR ;
   q_16_1 <= q_16_1_EXMPLR ;
   q_16_0 <= q_16_0_EXMPLR ;
   q_17_15 <= q_17_15_EXMPLR ;
   q_17_14 <= q_17_14_EXMPLR ;
   q_17_13 <= q_17_13_EXMPLR ;
   q_17_12 <= q_17_12_EXMPLR ;
   q_17_11 <= q_17_11_EXMPLR ;
   q_17_10 <= q_17_10_EXMPLR ;
   q_17_9 <= q_17_9_EXMPLR ;
   q_17_8 <= q_17_8_EXMPLR ;
   q_17_7 <= q_17_7_EXMPLR ;
   q_17_6 <= q_17_6_EXMPLR ;
   q_17_5 <= q_17_5_EXMPLR ;
   q_17_4 <= q_17_4_EXMPLR ;
   q_17_3 <= q_17_3_EXMPLR ;
   q_17_2 <= q_17_2_EXMPLR ;
   q_17_1 <= q_17_1_EXMPLR ;
   q_17_0 <= q_17_0_EXMPLR ;
   q_18_15 <= q_18_15_EXMPLR ;
   q_18_14 <= q_18_14_EXMPLR ;
   q_18_13 <= q_18_13_EXMPLR ;
   q_18_12 <= q_18_12_EXMPLR ;
   q_18_11 <= q_18_11_EXMPLR ;
   q_18_10 <= q_18_10_EXMPLR ;
   q_18_9 <= q_18_9_EXMPLR ;
   q_18_8 <= q_18_8_EXMPLR ;
   q_18_7 <= q_18_7_EXMPLR ;
   q_18_6 <= q_18_6_EXMPLR ;
   q_18_5 <= q_18_5_EXMPLR ;
   q_18_4 <= q_18_4_EXMPLR ;
   q_18_3 <= q_18_3_EXMPLR ;
   q_18_2 <= q_18_2_EXMPLR ;
   q_18_1 <= q_18_1_EXMPLR ;
   q_18_0 <= q_18_0_EXMPLR ;
   q_19_15 <= q_19_15_EXMPLR ;
   q_19_14 <= q_19_14_EXMPLR ;
   q_19_13 <= q_19_13_EXMPLR ;
   q_19_12 <= q_19_12_EXMPLR ;
   q_19_11 <= q_19_11_EXMPLR ;
   q_19_10 <= q_19_10_EXMPLR ;
   q_19_9 <= q_19_9_EXMPLR ;
   q_19_8 <= q_19_8_EXMPLR ;
   q_19_7 <= q_19_7_EXMPLR ;
   q_19_6 <= q_19_6_EXMPLR ;
   q_19_5 <= q_19_5_EXMPLR ;
   q_19_4 <= q_19_4_EXMPLR ;
   q_19_3 <= q_19_3_EXMPLR ;
   q_19_2 <= q_19_2_EXMPLR ;
   q_19_1 <= q_19_1_EXMPLR ;
   q_19_0 <= q_19_0_EXMPLR ;
   q_20_15 <= q_20_15_EXMPLR ;
   q_20_14 <= q_20_14_EXMPLR ;
   q_20_13 <= q_20_13_EXMPLR ;
   q_20_12 <= q_20_12_EXMPLR ;
   q_20_11 <= q_20_11_EXMPLR ;
   q_20_10 <= q_20_10_EXMPLR ;
   q_20_9 <= q_20_9_EXMPLR ;
   q_20_8 <= q_20_8_EXMPLR ;
   q_20_7 <= q_20_7_EXMPLR ;
   q_20_6 <= q_20_6_EXMPLR ;
   q_20_5 <= q_20_5_EXMPLR ;
   q_20_4 <= q_20_4_EXMPLR ;
   q_20_3 <= q_20_3_EXMPLR ;
   q_20_2 <= q_20_2_EXMPLR ;
   q_20_1 <= q_20_1_EXMPLR ;
   q_20_0 <= q_20_0_EXMPLR ;
   q_21_15 <= q_21_15_EXMPLR ;
   q_21_14 <= q_21_14_EXMPLR ;
   q_21_13 <= q_21_13_EXMPLR ;
   q_21_12 <= q_21_12_EXMPLR ;
   q_21_11 <= q_21_11_EXMPLR ;
   q_21_10 <= q_21_10_EXMPLR ;
   q_21_9 <= q_21_9_EXMPLR ;
   q_21_8 <= q_21_8_EXMPLR ;
   q_21_7 <= q_21_7_EXMPLR ;
   q_21_6 <= q_21_6_EXMPLR ;
   q_21_5 <= q_21_5_EXMPLR ;
   q_21_4 <= q_21_4_EXMPLR ;
   q_21_3 <= q_21_3_EXMPLR ;
   q_21_2 <= q_21_2_EXMPLR ;
   q_21_1 <= q_21_1_EXMPLR ;
   q_21_0 <= q_21_0_EXMPLR ;
   q_22_15 <= q_22_15_EXMPLR ;
   q_22_14 <= q_22_14_EXMPLR ;
   q_22_13 <= q_22_13_EXMPLR ;
   q_22_12 <= q_22_12_EXMPLR ;
   q_22_11 <= q_22_11_EXMPLR ;
   q_22_10 <= q_22_10_EXMPLR ;
   q_22_9 <= q_22_9_EXMPLR ;
   q_22_8 <= q_22_8_EXMPLR ;
   q_22_7 <= q_22_7_EXMPLR ;
   q_22_6 <= q_22_6_EXMPLR ;
   q_22_5 <= q_22_5_EXMPLR ;
   q_22_4 <= q_22_4_EXMPLR ;
   q_22_3 <= q_22_3_EXMPLR ;
   q_22_2 <= q_22_2_EXMPLR ;
   q_22_1 <= q_22_1_EXMPLR ;
   q_22_0 <= q_22_0_EXMPLR ;
   q_23_15 <= q_23_15_EXMPLR ;
   q_23_14 <= q_23_14_EXMPLR ;
   q_23_13 <= q_23_13_EXMPLR ;
   q_23_12 <= q_23_12_EXMPLR ;
   q_23_11 <= q_23_11_EXMPLR ;
   q_23_10 <= q_23_10_EXMPLR ;
   q_23_9 <= q_23_9_EXMPLR ;
   q_23_8 <= q_23_8_EXMPLR ;
   q_23_7 <= q_23_7_EXMPLR ;
   q_23_6 <= q_23_6_EXMPLR ;
   q_23_5 <= q_23_5_EXMPLR ;
   q_23_4 <= q_23_4_EXMPLR ;
   q_23_3 <= q_23_3_EXMPLR ;
   q_23_2 <= q_23_2_EXMPLR ;
   q_23_1 <= q_23_1_EXMPLR ;
   q_23_0 <= q_23_0_EXMPLR ;
   q_24_15 <= q_24_15_EXMPLR ;
   q_24_14 <= q_24_14_EXMPLR ;
   q_24_13 <= q_24_13_EXMPLR ;
   q_24_12 <= q_24_12_EXMPLR ;
   q_24_11 <= q_24_11_EXMPLR ;
   q_24_10 <= q_24_10_EXMPLR ;
   q_24_9 <= q_24_9_EXMPLR ;
   q_24_8 <= q_24_8_EXMPLR ;
   q_24_7 <= q_24_7_EXMPLR ;
   q_24_6 <= q_24_6_EXMPLR ;
   q_24_5 <= q_24_5_EXMPLR ;
   q_24_4 <= q_24_4_EXMPLR ;
   q_24_3 <= q_24_3_EXMPLR ;
   q_24_2 <= q_24_2_EXMPLR ;
   q_24_1 <= q_24_1_EXMPLR ;
   q_24_0 <= q_24_0_EXMPLR ;
   gen_regs_24_regi_reg_q_0 : dffr port map ( Q=>q_24_0_EXMPLR, QB=>OPEN, D
      =>nx1973, CLK=>nx7064, R=>reset);
   ix1974 : mux21_ni port map ( Y=>nx1973, A0=>q_24_0_EXMPLR, A1=>
      q_23_0_EXMPLR, S0=>nx6946);
   gen_regs_23_regi_reg_q_0 : dffr port map ( Q=>q_23_0_EXMPLR, QB=>OPEN, D
      =>nx1963, CLK=>nx7064, R=>reset);
   ix1964 : mux21_ni port map ( Y=>nx1963, A0=>q_23_0_EXMPLR, A1=>
      q_22_0_EXMPLR, S0=>nx6946);
   gen_regs_22_regi_reg_q_0 : dffr port map ( Q=>q_22_0_EXMPLR, QB=>OPEN, D
      =>nx1953, CLK=>nx7064, R=>reset);
   ix1954 : mux21_ni port map ( Y=>nx1953, A0=>q_22_0_EXMPLR, A1=>
      q_21_0_EXMPLR, S0=>nx6946);
   gen_regs_21_regi_reg_q_0 : dffr port map ( Q=>q_21_0_EXMPLR, QB=>OPEN, D
      =>nx1943, CLK=>nx7064, R=>reset);
   ix1944 : mux21_ni port map ( Y=>nx1943, A0=>q_21_0_EXMPLR, A1=>
      q_20_0_EXMPLR, S0=>nx6946);
   gen_regs_20_regi_reg_q_0 : dffr port map ( Q=>q_20_0_EXMPLR, QB=>OPEN, D
      =>nx1933, CLK=>nx7062, R=>reset);
   ix1934 : mux21_ni port map ( Y=>nx1933, A0=>q_20_0_EXMPLR, A1=>
      q_19_0_EXMPLR, S0=>nx6944);
   gen_regs_19_regi_reg_q_0 : dffr port map ( Q=>q_19_0_EXMPLR, QB=>OPEN, D
      =>nx1923, CLK=>nx7062, R=>reset);
   ix1924 : mux21_ni port map ( Y=>nx1923, A0=>q_19_0_EXMPLR, A1=>
      q_18_0_EXMPLR, S0=>nx6944);
   gen_regs_18_regi_reg_q_0 : dffr port map ( Q=>q_18_0_EXMPLR, QB=>OPEN, D
      =>nx1913, CLK=>nx7062, R=>reset);
   ix1914 : mux21_ni port map ( Y=>nx1913, A0=>q_18_0_EXMPLR, A1=>
      q_17_0_EXMPLR, S0=>nx6944);
   gen_regs_17_regi_reg_q_0 : dffr port map ( Q=>q_17_0_EXMPLR, QB=>OPEN, D
      =>nx1903, CLK=>nx7062, R=>reset);
   ix1904 : mux21_ni port map ( Y=>nx1903, A0=>q_17_0_EXMPLR, A1=>
      q_16_0_EXMPLR, S0=>nx6944);
   gen_regs_16_regi_reg_q_0 : dffr port map ( Q=>q_16_0_EXMPLR, QB=>OPEN, D
      =>nx1893, CLK=>nx7062, R=>reset);
   ix1894 : mux21_ni port map ( Y=>nx1893, A0=>q_16_0_EXMPLR, A1=>
      q_15_0_EXMPLR, S0=>nx6944);
   gen_regs_15_regi_reg_q_0 : dffr port map ( Q=>q_15_0_EXMPLR, QB=>OPEN, D
      =>nx1883, CLK=>nx7062, R=>reset);
   ix1884 : mux21_ni port map ( Y=>nx1883, A0=>q_15_0_EXMPLR, A1=>
      q_14_0_EXMPLR, S0=>nx6944);
   gen_regs_14_regi_reg_q_0 : dffr port map ( Q=>q_14_0_EXMPLR, QB=>OPEN, D
      =>nx1873, CLK=>nx7062, R=>reset);
   ix1874 : mux21_ni port map ( Y=>nx1873, A0=>q_14_0_EXMPLR, A1=>
      q_13_0_EXMPLR, S0=>nx6944);
   gen_regs_13_regi_reg_q_0 : dffr port map ( Q=>q_13_0_EXMPLR, QB=>OPEN, D
      =>nx1863, CLK=>nx7060, R=>reset);
   ix1864 : mux21_ni port map ( Y=>nx1863, A0=>q_13_0_EXMPLR, A1=>
      q_12_0_EXMPLR, S0=>nx6942);
   gen_regs_12_regi_reg_q_0 : dffr port map ( Q=>q_12_0_EXMPLR, QB=>OPEN, D
      =>nx1853, CLK=>nx7060, R=>reset);
   ix1854 : mux21_ni port map ( Y=>nx1853, A0=>q_12_0_EXMPLR, A1=>
      q_11_0_EXMPLR, S0=>nx6942);
   gen_regs_11_regi_reg_q_0 : dffr port map ( Q=>q_11_0_EXMPLR, QB=>OPEN, D
      =>nx1843, CLK=>nx7060, R=>reset);
   ix1844 : mux21_ni port map ( Y=>nx1843, A0=>q_11_0_EXMPLR, A1=>
      q_10_0_EXMPLR, S0=>nx6942);
   gen_regs_10_regi_reg_q_0 : dffr port map ( Q=>q_10_0_EXMPLR, QB=>OPEN, D
      =>nx1833, CLK=>nx7060, R=>reset);
   ix1834 : mux21_ni port map ( Y=>nx1833, A0=>q_10_0_EXMPLR, A1=>
      q_9_0_EXMPLR, S0=>nx6942);
   gen_regs_9_regi_reg_q_0 : dffr port map ( Q=>q_9_0_EXMPLR, QB=>OPEN, D=>
      nx1823, CLK=>nx7060, R=>reset);
   ix1824 : mux21_ni port map ( Y=>nx1823, A0=>q_9_0_EXMPLR, A1=>
      q_8_0_EXMPLR, S0=>nx6942);
   gen_regs_8_regi_reg_q_0 : dffr port map ( Q=>q_8_0_EXMPLR, QB=>OPEN, D=>
      nx1813, CLK=>nx7060, R=>reset);
   ix1814 : mux21_ni port map ( Y=>nx1813, A0=>q_8_0_EXMPLR, A1=>
      q_7_0_EXMPLR, S0=>nx6942);
   gen_regs_7_regi_reg_q_0 : dffr port map ( Q=>q_7_0_EXMPLR, QB=>OPEN, D=>
      nx1803, CLK=>nx7060, R=>reset);
   ix1804 : mux21_ni port map ( Y=>nx1803, A0=>q_7_0_EXMPLR, A1=>
      q_6_0_EXMPLR, S0=>nx6942);
   gen_regs_6_regi_reg_q_0 : dffr port map ( Q=>q_6_0_EXMPLR, QB=>OPEN, D=>
      nx1793, CLK=>nx7058, R=>reset);
   ix1794 : mux21_ni port map ( Y=>nx1793, A0=>q_6_0_EXMPLR, A1=>
      q_5_0_EXMPLR, S0=>nx6940);
   gen_regs_5_regi_reg_q_0 : dffr port map ( Q=>q_5_0_EXMPLR, QB=>OPEN, D=>
      nx1783, CLK=>nx7058, R=>reset);
   ix1784 : mux21_ni port map ( Y=>nx1783, A0=>q_5_0_EXMPLR, A1=>
      q_4_0_EXMPLR, S0=>nx6940);
   gen_regs_4_regi_reg_q_0 : dffr port map ( Q=>q_4_0_EXMPLR, QB=>OPEN, D=>
      nx1773, CLK=>nx7058, R=>reset);
   ix1774 : mux21_ni port map ( Y=>nx1773, A0=>q_4_0_EXMPLR, A1=>
      q_3_0_EXMPLR, S0=>nx6940);
   gen_regs_3_regi_reg_q_0 : dffr port map ( Q=>q_3_0_EXMPLR, QB=>OPEN, D=>
      nx1763, CLK=>nx7058, R=>reset);
   ix1764 : mux21_ni port map ( Y=>nx1763, A0=>q_3_0_EXMPLR, A1=>
      q_2_0_EXMPLR, S0=>nx6940);
   gen_regs_2_regi_reg_q_0 : dffr port map ( Q=>q_2_0_EXMPLR, QB=>OPEN, D=>
      nx1753, CLK=>nx7058, R=>reset);
   ix1754 : mux21_ni port map ( Y=>nx1753, A0=>q_2_0_EXMPLR, A1=>
      q_1_0_EXMPLR, S0=>nx6940);
   gen_regs_1_regi_reg_q_0 : dffr port map ( Q=>q_1_0_EXMPLR, QB=>OPEN, D=>
      nx1743, CLK=>nx7058, R=>reset);
   ix1744 : mux21_ni port map ( Y=>nx1743, A0=>q_1_0_EXMPLR, A1=>
      q_0_0_EXMPLR, S0=>nx6940);
   reg0_reg_q_0 : dffr port map ( Q=>q_0_0_EXMPLR, QB=>OPEN, D=>nx1733, CLK
      =>nx7058, R=>reset);
   ix1734 : mux21_ni port map ( Y=>nx1733, A0=>q_0_0_EXMPLR, A1=>d(0), S0=>
      nx6940);
   gen_regs_24_regi_reg_q_1 : dffr port map ( Q=>q_24_1_EXMPLR, QB=>OPEN, D
      =>nx2223, CLK=>nx7072, R=>reset);
   ix2224 : mux21_ni port map ( Y=>nx2223, A0=>q_24_1_EXMPLR, A1=>
      q_23_1_EXMPLR, S0=>nx6954);
   gen_regs_23_regi_reg_q_1 : dffr port map ( Q=>q_23_1_EXMPLR, QB=>OPEN, D
      =>nx2213, CLK=>nx7070, R=>reset);
   ix2214 : mux21_ni port map ( Y=>nx2213, A0=>q_23_1_EXMPLR, A1=>
      q_22_1_EXMPLR, S0=>nx6952);
   gen_regs_22_regi_reg_q_1 : dffr port map ( Q=>q_22_1_EXMPLR, QB=>OPEN, D
      =>nx2203, CLK=>nx7070, R=>reset);
   ix2204 : mux21_ni port map ( Y=>nx2203, A0=>q_22_1_EXMPLR, A1=>
      q_21_1_EXMPLR, S0=>nx6952);
   gen_regs_21_regi_reg_q_1 : dffr port map ( Q=>q_21_1_EXMPLR, QB=>OPEN, D
      =>nx2193, CLK=>nx7070, R=>reset);
   ix2194 : mux21_ni port map ( Y=>nx2193, A0=>q_21_1_EXMPLR, A1=>
      q_20_1_EXMPLR, S0=>nx6952);
   gen_regs_20_regi_reg_q_1 : dffr port map ( Q=>q_20_1_EXMPLR, QB=>OPEN, D
      =>nx2183, CLK=>nx7070, R=>reset);
   ix2184 : mux21_ni port map ( Y=>nx2183, A0=>q_20_1_EXMPLR, A1=>
      q_19_1_EXMPLR, S0=>nx6952);
   gen_regs_19_regi_reg_q_1 : dffr port map ( Q=>q_19_1_EXMPLR, QB=>OPEN, D
      =>nx2173, CLK=>nx7070, R=>reset);
   ix2174 : mux21_ni port map ( Y=>nx2173, A0=>q_19_1_EXMPLR, A1=>
      q_18_1_EXMPLR, S0=>nx6952);
   gen_regs_18_regi_reg_q_1 : dffr port map ( Q=>q_18_1_EXMPLR, QB=>OPEN, D
      =>nx2163, CLK=>nx7070, R=>reset);
   ix2164 : mux21_ni port map ( Y=>nx2163, A0=>q_18_1_EXMPLR, A1=>
      q_17_1_EXMPLR, S0=>nx6952);
   gen_regs_17_regi_reg_q_1 : dffr port map ( Q=>q_17_1_EXMPLR, QB=>OPEN, D
      =>nx2153, CLK=>nx7070, R=>reset);
   ix2154 : mux21_ni port map ( Y=>nx2153, A0=>q_17_1_EXMPLR, A1=>
      q_16_1_EXMPLR, S0=>nx6952);
   gen_regs_16_regi_reg_q_1 : dffr port map ( Q=>q_16_1_EXMPLR, QB=>OPEN, D
      =>nx2143, CLK=>nx7068, R=>reset);
   ix2144 : mux21_ni port map ( Y=>nx2143, A0=>q_16_1_EXMPLR, A1=>
      q_15_1_EXMPLR, S0=>nx6950);
   gen_regs_15_regi_reg_q_1 : dffr port map ( Q=>q_15_1_EXMPLR, QB=>OPEN, D
      =>nx2133, CLK=>nx7068, R=>reset);
   ix2134 : mux21_ni port map ( Y=>nx2133, A0=>q_15_1_EXMPLR, A1=>
      q_14_1_EXMPLR, S0=>nx6950);
   gen_regs_14_regi_reg_q_1 : dffr port map ( Q=>q_14_1_EXMPLR, QB=>OPEN, D
      =>nx2123, CLK=>nx7068, R=>reset);
   ix2124 : mux21_ni port map ( Y=>nx2123, A0=>q_14_1_EXMPLR, A1=>
      q_13_1_EXMPLR, S0=>nx6950);
   gen_regs_13_regi_reg_q_1 : dffr port map ( Q=>q_13_1_EXMPLR, QB=>OPEN, D
      =>nx2113, CLK=>nx7068, R=>reset);
   ix2114 : mux21_ni port map ( Y=>nx2113, A0=>q_13_1_EXMPLR, A1=>
      q_12_1_EXMPLR, S0=>nx6950);
   gen_regs_12_regi_reg_q_1 : dffr port map ( Q=>q_12_1_EXMPLR, QB=>OPEN, D
      =>nx2103, CLK=>nx7068, R=>reset);
   ix2104 : mux21_ni port map ( Y=>nx2103, A0=>q_12_1_EXMPLR, A1=>
      q_11_1_EXMPLR, S0=>nx6950);
   gen_regs_11_regi_reg_q_1 : dffr port map ( Q=>q_11_1_EXMPLR, QB=>OPEN, D
      =>nx2093, CLK=>nx7068, R=>reset);
   ix2094 : mux21_ni port map ( Y=>nx2093, A0=>q_11_1_EXMPLR, A1=>
      q_10_1_EXMPLR, S0=>nx6950);
   gen_regs_10_regi_reg_q_1 : dffr port map ( Q=>q_10_1_EXMPLR, QB=>OPEN, D
      =>nx2083, CLK=>nx7068, R=>reset);
   ix2084 : mux21_ni port map ( Y=>nx2083, A0=>q_10_1_EXMPLR, A1=>
      q_9_1_EXMPLR, S0=>nx6950);
   gen_regs_9_regi_reg_q_1 : dffr port map ( Q=>q_9_1_EXMPLR, QB=>OPEN, D=>
      nx2073, CLK=>nx7066, R=>reset);
   ix2074 : mux21_ni port map ( Y=>nx2073, A0=>q_9_1_EXMPLR, A1=>
      q_8_1_EXMPLR, S0=>nx6948);
   gen_regs_8_regi_reg_q_1 : dffr port map ( Q=>q_8_1_EXMPLR, QB=>OPEN, D=>
      nx2063, CLK=>nx7066, R=>reset);
   ix2064 : mux21_ni port map ( Y=>nx2063, A0=>q_8_1_EXMPLR, A1=>
      q_7_1_EXMPLR, S0=>nx6948);
   gen_regs_7_regi_reg_q_1 : dffr port map ( Q=>q_7_1_EXMPLR, QB=>OPEN, D=>
      nx2053, CLK=>nx7066, R=>reset);
   ix2054 : mux21_ni port map ( Y=>nx2053, A0=>q_7_1_EXMPLR, A1=>
      q_6_1_EXMPLR, S0=>nx6948);
   gen_regs_6_regi_reg_q_1 : dffr port map ( Q=>q_6_1_EXMPLR, QB=>OPEN, D=>
      nx2043, CLK=>nx7066, R=>reset);
   ix2044 : mux21_ni port map ( Y=>nx2043, A0=>q_6_1_EXMPLR, A1=>
      q_5_1_EXMPLR, S0=>nx6948);
   gen_regs_5_regi_reg_q_1 : dffr port map ( Q=>q_5_1_EXMPLR, QB=>OPEN, D=>
      nx2033, CLK=>nx7066, R=>reset);
   ix2034 : mux21_ni port map ( Y=>nx2033, A0=>q_5_1_EXMPLR, A1=>
      q_4_1_EXMPLR, S0=>nx6948);
   gen_regs_4_regi_reg_q_1 : dffr port map ( Q=>q_4_1_EXMPLR, QB=>OPEN, D=>
      nx2023, CLK=>nx7066, R=>reset);
   ix2024 : mux21_ni port map ( Y=>nx2023, A0=>q_4_1_EXMPLR, A1=>
      q_3_1_EXMPLR, S0=>nx6948);
   gen_regs_3_regi_reg_q_1 : dffr port map ( Q=>q_3_1_EXMPLR, QB=>OPEN, D=>
      nx2013, CLK=>nx7066, R=>reset);
   ix2014 : mux21_ni port map ( Y=>nx2013, A0=>q_3_1_EXMPLR, A1=>
      q_2_1_EXMPLR, S0=>nx6948);
   gen_regs_2_regi_reg_q_1 : dffr port map ( Q=>q_2_1_EXMPLR, QB=>OPEN, D=>
      nx2003, CLK=>nx7064, R=>reset);
   ix2004 : mux21_ni port map ( Y=>nx2003, A0=>q_2_1_EXMPLR, A1=>
      q_1_1_EXMPLR, S0=>nx6946);
   gen_regs_1_regi_reg_q_1 : dffr port map ( Q=>q_1_1_EXMPLR, QB=>OPEN, D=>
      nx1993, CLK=>nx7064, R=>reset);
   ix1994 : mux21_ni port map ( Y=>nx1993, A0=>q_1_1_EXMPLR, A1=>
      q_0_1_EXMPLR, S0=>nx6946);
   reg0_reg_q_1 : dffr port map ( Q=>q_0_1_EXMPLR, QB=>OPEN, D=>nx1983, CLK
      =>nx7064, R=>reset);
   ix1984 : mux21_ni port map ( Y=>nx1983, A0=>q_0_1_EXMPLR, A1=>d(1), S0=>
      nx6946);
   gen_regs_24_regi_reg_q_2 : dffr port map ( Q=>q_24_2_EXMPLR, QB=>OPEN, D
      =>nx2473, CLK=>nx7078, R=>reset);
   ix2474 : mux21_ni port map ( Y=>nx2473, A0=>q_24_2_EXMPLR, A1=>
      q_23_2_EXMPLR, S0=>nx6960);
   gen_regs_23_regi_reg_q_2 : dffr port map ( Q=>q_23_2_EXMPLR, QB=>OPEN, D
      =>nx2463, CLK=>nx7078, R=>reset);
   ix2464 : mux21_ni port map ( Y=>nx2463, A0=>q_23_2_EXMPLR, A1=>
      q_22_2_EXMPLR, S0=>nx6960);
   gen_regs_22_regi_reg_q_2 : dffr port map ( Q=>q_22_2_EXMPLR, QB=>OPEN, D
      =>nx2453, CLK=>nx7078, R=>reset);
   ix2454 : mux21_ni port map ( Y=>nx2453, A0=>q_22_2_EXMPLR, A1=>
      q_21_2_EXMPLR, S0=>nx6960);
   gen_regs_21_regi_reg_q_2 : dffr port map ( Q=>q_21_2_EXMPLR, QB=>OPEN, D
      =>nx2443, CLK=>nx7078, R=>reset);
   ix2444 : mux21_ni port map ( Y=>nx2443, A0=>q_21_2_EXMPLR, A1=>
      q_20_2_EXMPLR, S0=>nx6960);
   gen_regs_20_regi_reg_q_2 : dffr port map ( Q=>q_20_2_EXMPLR, QB=>OPEN, D
      =>nx2433, CLK=>nx7078, R=>reset);
   ix2434 : mux21_ni port map ( Y=>nx2433, A0=>q_20_2_EXMPLR, A1=>
      q_19_2_EXMPLR, S0=>nx6960);
   gen_regs_19_regi_reg_q_2 : dffr port map ( Q=>q_19_2_EXMPLR, QB=>OPEN, D
      =>nx2423, CLK=>nx7076, R=>reset);
   ix2424 : mux21_ni port map ( Y=>nx2423, A0=>q_19_2_EXMPLR, A1=>
      q_18_2_EXMPLR, S0=>nx6958);
   gen_regs_18_regi_reg_q_2 : dffr port map ( Q=>q_18_2_EXMPLR, QB=>OPEN, D
      =>nx2413, CLK=>nx7076, R=>reset);
   ix2414 : mux21_ni port map ( Y=>nx2413, A0=>q_18_2_EXMPLR, A1=>
      q_17_2_EXMPLR, S0=>nx6958);
   gen_regs_17_regi_reg_q_2 : dffr port map ( Q=>q_17_2_EXMPLR, QB=>OPEN, D
      =>nx2403, CLK=>nx7076, R=>reset);
   ix2404 : mux21_ni port map ( Y=>nx2403, A0=>q_17_2_EXMPLR, A1=>
      q_16_2_EXMPLR, S0=>nx6958);
   gen_regs_16_regi_reg_q_2 : dffr port map ( Q=>q_16_2_EXMPLR, QB=>OPEN, D
      =>nx2393, CLK=>nx7076, R=>reset);
   ix2394 : mux21_ni port map ( Y=>nx2393, A0=>q_16_2_EXMPLR, A1=>
      q_15_2_EXMPLR, S0=>nx6958);
   gen_regs_15_regi_reg_q_2 : dffr port map ( Q=>q_15_2_EXMPLR, QB=>OPEN, D
      =>nx2383, CLK=>nx7076, R=>reset);
   ix2384 : mux21_ni port map ( Y=>nx2383, A0=>q_15_2_EXMPLR, A1=>
      q_14_2_EXMPLR, S0=>nx6958);
   gen_regs_14_regi_reg_q_2 : dffr port map ( Q=>q_14_2_EXMPLR, QB=>OPEN, D
      =>nx2373, CLK=>nx7076, R=>reset);
   ix2374 : mux21_ni port map ( Y=>nx2373, A0=>q_14_2_EXMPLR, A1=>
      q_13_2_EXMPLR, S0=>nx6958);
   gen_regs_13_regi_reg_q_2 : dffr port map ( Q=>q_13_2_EXMPLR, QB=>OPEN, D
      =>nx2363, CLK=>nx7076, R=>reset);
   ix2364 : mux21_ni port map ( Y=>nx2363, A0=>q_13_2_EXMPLR, A1=>
      q_12_2_EXMPLR, S0=>nx6958);
   gen_regs_12_regi_reg_q_2 : dffr port map ( Q=>q_12_2_EXMPLR, QB=>OPEN, D
      =>nx2353, CLK=>nx7074, R=>reset);
   ix2354 : mux21_ni port map ( Y=>nx2353, A0=>q_12_2_EXMPLR, A1=>
      q_11_2_EXMPLR, S0=>nx6956);
   gen_regs_11_regi_reg_q_2 : dffr port map ( Q=>q_11_2_EXMPLR, QB=>OPEN, D
      =>nx2343, CLK=>nx7074, R=>reset);
   ix2344 : mux21_ni port map ( Y=>nx2343, A0=>q_11_2_EXMPLR, A1=>
      q_10_2_EXMPLR, S0=>nx6956);
   gen_regs_10_regi_reg_q_2 : dffr port map ( Q=>q_10_2_EXMPLR, QB=>OPEN, D
      =>nx2333, CLK=>nx7074, R=>reset);
   ix2334 : mux21_ni port map ( Y=>nx2333, A0=>q_10_2_EXMPLR, A1=>
      q_9_2_EXMPLR, S0=>nx6956);
   gen_regs_9_regi_reg_q_2 : dffr port map ( Q=>q_9_2_EXMPLR, QB=>OPEN, D=>
      nx2323, CLK=>nx7074, R=>reset);
   ix2324 : mux21_ni port map ( Y=>nx2323, A0=>q_9_2_EXMPLR, A1=>
      q_8_2_EXMPLR, S0=>nx6956);
   gen_regs_8_regi_reg_q_2 : dffr port map ( Q=>q_8_2_EXMPLR, QB=>OPEN, D=>
      nx2313, CLK=>nx7074, R=>reset);
   ix2314 : mux21_ni port map ( Y=>nx2313, A0=>q_8_2_EXMPLR, A1=>
      q_7_2_EXMPLR, S0=>nx6956);
   gen_regs_7_regi_reg_q_2 : dffr port map ( Q=>q_7_2_EXMPLR, QB=>OPEN, D=>
      nx2303, CLK=>nx7074, R=>reset);
   ix2304 : mux21_ni port map ( Y=>nx2303, A0=>q_7_2_EXMPLR, A1=>
      q_6_2_EXMPLR, S0=>nx6956);
   gen_regs_6_regi_reg_q_2 : dffr port map ( Q=>q_6_2_EXMPLR, QB=>OPEN, D=>
      nx2293, CLK=>nx7074, R=>reset);
   ix2294 : mux21_ni port map ( Y=>nx2293, A0=>q_6_2_EXMPLR, A1=>
      q_5_2_EXMPLR, S0=>nx6956);
   gen_regs_5_regi_reg_q_2 : dffr port map ( Q=>q_5_2_EXMPLR, QB=>OPEN, D=>
      nx2283, CLK=>nx7072, R=>reset);
   ix2284 : mux21_ni port map ( Y=>nx2283, A0=>q_5_2_EXMPLR, A1=>
      q_4_2_EXMPLR, S0=>nx6954);
   gen_regs_4_regi_reg_q_2 : dffr port map ( Q=>q_4_2_EXMPLR, QB=>OPEN, D=>
      nx2273, CLK=>nx7072, R=>reset);
   ix2274 : mux21_ni port map ( Y=>nx2273, A0=>q_4_2_EXMPLR, A1=>
      q_3_2_EXMPLR, S0=>nx6954);
   gen_regs_3_regi_reg_q_2 : dffr port map ( Q=>q_3_2_EXMPLR, QB=>OPEN, D=>
      nx2263, CLK=>nx7072, R=>reset);
   ix2264 : mux21_ni port map ( Y=>nx2263, A0=>q_3_2_EXMPLR, A1=>
      q_2_2_EXMPLR, S0=>nx6954);
   gen_regs_2_regi_reg_q_2 : dffr port map ( Q=>q_2_2_EXMPLR, QB=>OPEN, D=>
      nx2253, CLK=>nx7072, R=>reset);
   ix2254 : mux21_ni port map ( Y=>nx2253, A0=>q_2_2_EXMPLR, A1=>
      q_1_2_EXMPLR, S0=>nx6954);
   gen_regs_1_regi_reg_q_2 : dffr port map ( Q=>q_1_2_EXMPLR, QB=>OPEN, D=>
      nx2243, CLK=>nx7072, R=>reset);
   ix2244 : mux21_ni port map ( Y=>nx2243, A0=>q_1_2_EXMPLR, A1=>
      q_0_2_EXMPLR, S0=>nx6954);
   reg0_reg_q_2 : dffr port map ( Q=>q_0_2_EXMPLR, QB=>OPEN, D=>nx2233, CLK
      =>nx7072, R=>reset);
   ix2234 : mux21_ni port map ( Y=>nx2233, A0=>q_0_2_EXMPLR, A1=>d(2), S0=>
      nx6954);
   gen_regs_24_regi_reg_q_3 : dffr port map ( Q=>q_24_3_EXMPLR, QB=>OPEN, D
      =>nx2723, CLK=>nx7086, R=>reset);
   ix2724 : mux21_ni port map ( Y=>nx2723, A0=>q_24_3_EXMPLR, A1=>
      q_23_3_EXMPLR, S0=>nx6968);
   gen_regs_23_regi_reg_q_3 : dffr port map ( Q=>q_23_3_EXMPLR, QB=>OPEN, D
      =>nx2713, CLK=>nx7086, R=>reset);
   ix2714 : mux21_ni port map ( Y=>nx2713, A0=>q_23_3_EXMPLR, A1=>
      q_22_3_EXMPLR, S0=>nx6968);
   gen_regs_22_regi_reg_q_3 : dffr port map ( Q=>q_22_3_EXMPLR, QB=>OPEN, D
      =>nx2703, CLK=>nx7084, R=>reset);
   ix2704 : mux21_ni port map ( Y=>nx2703, A0=>q_22_3_EXMPLR, A1=>
      q_21_3_EXMPLR, S0=>nx6966);
   gen_regs_21_regi_reg_q_3 : dffr port map ( Q=>q_21_3_EXMPLR, QB=>OPEN, D
      =>nx2693, CLK=>nx7084, R=>reset);
   ix2694 : mux21_ni port map ( Y=>nx2693, A0=>q_21_3_EXMPLR, A1=>
      q_20_3_EXMPLR, S0=>nx6966);
   gen_regs_20_regi_reg_q_3 : dffr port map ( Q=>q_20_3_EXMPLR, QB=>OPEN, D
      =>nx2683, CLK=>nx7084, R=>reset);
   ix2684 : mux21_ni port map ( Y=>nx2683, A0=>q_20_3_EXMPLR, A1=>
      q_19_3_EXMPLR, S0=>nx6966);
   gen_regs_19_regi_reg_q_3 : dffr port map ( Q=>q_19_3_EXMPLR, QB=>OPEN, D
      =>nx2673, CLK=>nx7084, R=>reset);
   ix2674 : mux21_ni port map ( Y=>nx2673, A0=>q_19_3_EXMPLR, A1=>
      q_18_3_EXMPLR, S0=>nx6966);
   gen_regs_18_regi_reg_q_3 : dffr port map ( Q=>q_18_3_EXMPLR, QB=>OPEN, D
      =>nx2663, CLK=>nx7084, R=>reset);
   ix2664 : mux21_ni port map ( Y=>nx2663, A0=>q_18_3_EXMPLR, A1=>
      q_17_3_EXMPLR, S0=>nx6966);
   gen_regs_17_regi_reg_q_3 : dffr port map ( Q=>q_17_3_EXMPLR, QB=>OPEN, D
      =>nx2653, CLK=>nx7084, R=>reset);
   ix2654 : mux21_ni port map ( Y=>nx2653, A0=>q_17_3_EXMPLR, A1=>
      q_16_3_EXMPLR, S0=>nx6966);
   gen_regs_16_regi_reg_q_3 : dffr port map ( Q=>q_16_3_EXMPLR, QB=>OPEN, D
      =>nx2643, CLK=>nx7084, R=>reset);
   ix2644 : mux21_ni port map ( Y=>nx2643, A0=>q_16_3_EXMPLR, A1=>
      q_15_3_EXMPLR, S0=>nx6966);
   gen_regs_15_regi_reg_q_3 : dffr port map ( Q=>q_15_3_EXMPLR, QB=>OPEN, D
      =>nx2633, CLK=>nx7082, R=>reset);
   ix2634 : mux21_ni port map ( Y=>nx2633, A0=>q_15_3_EXMPLR, A1=>
      q_14_3_EXMPLR, S0=>nx6964);
   gen_regs_14_regi_reg_q_3 : dffr port map ( Q=>q_14_3_EXMPLR, QB=>OPEN, D
      =>nx2623, CLK=>nx7082, R=>reset);
   ix2624 : mux21_ni port map ( Y=>nx2623, A0=>q_14_3_EXMPLR, A1=>
      q_13_3_EXMPLR, S0=>nx6964);
   gen_regs_13_regi_reg_q_3 : dffr port map ( Q=>q_13_3_EXMPLR, QB=>OPEN, D
      =>nx2613, CLK=>nx7082, R=>reset);
   ix2614 : mux21_ni port map ( Y=>nx2613, A0=>q_13_3_EXMPLR, A1=>
      q_12_3_EXMPLR, S0=>nx6964);
   gen_regs_12_regi_reg_q_3 : dffr port map ( Q=>q_12_3_EXMPLR, QB=>OPEN, D
      =>nx2603, CLK=>nx7082, R=>reset);
   ix2604 : mux21_ni port map ( Y=>nx2603, A0=>q_12_3_EXMPLR, A1=>
      q_11_3_EXMPLR, S0=>nx6964);
   gen_regs_11_regi_reg_q_3 : dffr port map ( Q=>q_11_3_EXMPLR, QB=>OPEN, D
      =>nx2593, CLK=>nx7082, R=>reset);
   ix2594 : mux21_ni port map ( Y=>nx2593, A0=>q_11_3_EXMPLR, A1=>
      q_10_3_EXMPLR, S0=>nx6964);
   gen_regs_10_regi_reg_q_3 : dffr port map ( Q=>q_10_3_EXMPLR, QB=>OPEN, D
      =>nx2583, CLK=>nx7082, R=>reset);
   ix2584 : mux21_ni port map ( Y=>nx2583, A0=>q_10_3_EXMPLR, A1=>
      q_9_3_EXMPLR, S0=>nx6964);
   gen_regs_9_regi_reg_q_3 : dffr port map ( Q=>q_9_3_EXMPLR, QB=>OPEN, D=>
      nx2573, CLK=>nx7082, R=>reset);
   ix2574 : mux21_ni port map ( Y=>nx2573, A0=>q_9_3_EXMPLR, A1=>
      q_8_3_EXMPLR, S0=>nx6964);
   gen_regs_8_regi_reg_q_3 : dffr port map ( Q=>q_8_3_EXMPLR, QB=>OPEN, D=>
      nx2563, CLK=>nx7080, R=>reset);
   ix2564 : mux21_ni port map ( Y=>nx2563, A0=>q_8_3_EXMPLR, A1=>
      q_7_3_EXMPLR, S0=>nx6962);
   gen_regs_7_regi_reg_q_3 : dffr port map ( Q=>q_7_3_EXMPLR, QB=>OPEN, D=>
      nx2553, CLK=>nx7080, R=>reset);
   ix2554 : mux21_ni port map ( Y=>nx2553, A0=>q_7_3_EXMPLR, A1=>
      q_6_3_EXMPLR, S0=>nx6962);
   gen_regs_6_regi_reg_q_3 : dffr port map ( Q=>q_6_3_EXMPLR, QB=>OPEN, D=>
      nx2543, CLK=>nx7080, R=>reset);
   ix2544 : mux21_ni port map ( Y=>nx2543, A0=>q_6_3_EXMPLR, A1=>
      q_5_3_EXMPLR, S0=>nx6962);
   gen_regs_5_regi_reg_q_3 : dffr port map ( Q=>q_5_3_EXMPLR, QB=>OPEN, D=>
      nx2533, CLK=>nx7080, R=>reset);
   ix2534 : mux21_ni port map ( Y=>nx2533, A0=>q_5_3_EXMPLR, A1=>
      q_4_3_EXMPLR, S0=>nx6962);
   gen_regs_4_regi_reg_q_3 : dffr port map ( Q=>q_4_3_EXMPLR, QB=>OPEN, D=>
      nx2523, CLK=>nx7080, R=>reset);
   ix2524 : mux21_ni port map ( Y=>nx2523, A0=>q_4_3_EXMPLR, A1=>
      q_3_3_EXMPLR, S0=>nx6962);
   gen_regs_3_regi_reg_q_3 : dffr port map ( Q=>q_3_3_EXMPLR, QB=>OPEN, D=>
      nx2513, CLK=>nx7080, R=>reset);
   ix2514 : mux21_ni port map ( Y=>nx2513, A0=>q_3_3_EXMPLR, A1=>
      q_2_3_EXMPLR, S0=>nx6962);
   gen_regs_2_regi_reg_q_3 : dffr port map ( Q=>q_2_3_EXMPLR, QB=>OPEN, D=>
      nx2503, CLK=>nx7080, R=>reset);
   ix2504 : mux21_ni port map ( Y=>nx2503, A0=>q_2_3_EXMPLR, A1=>
      q_1_3_EXMPLR, S0=>nx6962);
   gen_regs_1_regi_reg_q_3 : dffr port map ( Q=>q_1_3_EXMPLR, QB=>OPEN, D=>
      nx2493, CLK=>nx7078, R=>reset);
   ix2494 : mux21_ni port map ( Y=>nx2493, A0=>q_1_3_EXMPLR, A1=>
      q_0_3_EXMPLR, S0=>nx6960);
   reg0_reg_q_3 : dffr port map ( Q=>q_0_3_EXMPLR, QB=>OPEN, D=>nx2483, CLK
      =>nx7078, R=>reset);
   ix2484 : mux21_ni port map ( Y=>nx2483, A0=>q_0_3_EXMPLR, A1=>d(3), S0=>
      nx6960);
   gen_regs_24_regi_reg_q_4 : dffr port map ( Q=>q_24_4_EXMPLR, QB=>OPEN, D
      =>nx2973, CLK=>nx7092, R=>reset);
   ix2974 : mux21_ni port map ( Y=>nx2973, A0=>q_24_4_EXMPLR, A1=>
      q_23_4_EXMPLR, S0=>nx6974);
   gen_regs_23_regi_reg_q_4 : dffr port map ( Q=>q_23_4_EXMPLR, QB=>OPEN, D
      =>nx2963, CLK=>nx7092, R=>reset);
   ix2964 : mux21_ni port map ( Y=>nx2963, A0=>q_23_4_EXMPLR, A1=>
      q_22_4_EXMPLR, S0=>nx6974);
   gen_regs_22_regi_reg_q_4 : dffr port map ( Q=>q_22_4_EXMPLR, QB=>OPEN, D
      =>nx2953, CLK=>nx7092, R=>reset);
   ix2954 : mux21_ni port map ( Y=>nx2953, A0=>q_22_4_EXMPLR, A1=>
      q_21_4_EXMPLR, S0=>nx6974);
   gen_regs_21_regi_reg_q_4 : dffr port map ( Q=>q_21_4_EXMPLR, QB=>OPEN, D
      =>nx2943, CLK=>nx7092, R=>reset);
   ix2944 : mux21_ni port map ( Y=>nx2943, A0=>q_21_4_EXMPLR, A1=>
      q_20_4_EXMPLR, S0=>nx6974);
   gen_regs_20_regi_reg_q_4 : dffr port map ( Q=>q_20_4_EXMPLR, QB=>OPEN, D
      =>nx2933, CLK=>nx7092, R=>reset);
   ix2934 : mux21_ni port map ( Y=>nx2933, A0=>q_20_4_EXMPLR, A1=>
      q_19_4_EXMPLR, S0=>nx6974);
   gen_regs_19_regi_reg_q_4 : dffr port map ( Q=>q_19_4_EXMPLR, QB=>OPEN, D
      =>nx2923, CLK=>nx7092, R=>reset);
   ix2924 : mux21_ni port map ( Y=>nx2923, A0=>q_19_4_EXMPLR, A1=>
      q_18_4_EXMPLR, S0=>nx6974);
   gen_regs_18_regi_reg_q_4 : dffr port map ( Q=>q_18_4_EXMPLR, QB=>OPEN, D
      =>nx2913, CLK=>nx7090, R=>reset);
   ix2914 : mux21_ni port map ( Y=>nx2913, A0=>q_18_4_EXMPLR, A1=>
      q_17_4_EXMPLR, S0=>nx6972);
   gen_regs_17_regi_reg_q_4 : dffr port map ( Q=>q_17_4_EXMPLR, QB=>OPEN, D
      =>nx2903, CLK=>nx7090, R=>reset);
   ix2904 : mux21_ni port map ( Y=>nx2903, A0=>q_17_4_EXMPLR, A1=>
      q_16_4_EXMPLR, S0=>nx6972);
   gen_regs_16_regi_reg_q_4 : dffr port map ( Q=>q_16_4_EXMPLR, QB=>OPEN, D
      =>nx2893, CLK=>nx7090, R=>reset);
   ix2894 : mux21_ni port map ( Y=>nx2893, A0=>q_16_4_EXMPLR, A1=>
      q_15_4_EXMPLR, S0=>nx6972);
   gen_regs_15_regi_reg_q_4 : dffr port map ( Q=>q_15_4_EXMPLR, QB=>OPEN, D
      =>nx2883, CLK=>nx7090, R=>reset);
   ix2884 : mux21_ni port map ( Y=>nx2883, A0=>q_15_4_EXMPLR, A1=>
      q_14_4_EXMPLR, S0=>nx6972);
   gen_regs_14_regi_reg_q_4 : dffr port map ( Q=>q_14_4_EXMPLR, QB=>OPEN, D
      =>nx2873, CLK=>nx7090, R=>reset);
   ix2874 : mux21_ni port map ( Y=>nx2873, A0=>q_14_4_EXMPLR, A1=>
      q_13_4_EXMPLR, S0=>nx6972);
   gen_regs_13_regi_reg_q_4 : dffr port map ( Q=>q_13_4_EXMPLR, QB=>OPEN, D
      =>nx2863, CLK=>nx7090, R=>reset);
   ix2864 : mux21_ni port map ( Y=>nx2863, A0=>q_13_4_EXMPLR, A1=>
      q_12_4_EXMPLR, S0=>nx6972);
   gen_regs_12_regi_reg_q_4 : dffr port map ( Q=>q_12_4_EXMPLR, QB=>OPEN, D
      =>nx2853, CLK=>nx7090, R=>reset);
   ix2854 : mux21_ni port map ( Y=>nx2853, A0=>q_12_4_EXMPLR, A1=>
      q_11_4_EXMPLR, S0=>nx6972);
   gen_regs_11_regi_reg_q_4 : dffr port map ( Q=>q_11_4_EXMPLR, QB=>OPEN, D
      =>nx2843, CLK=>nx7088, R=>reset);
   ix2844 : mux21_ni port map ( Y=>nx2843, A0=>q_11_4_EXMPLR, A1=>
      q_10_4_EXMPLR, S0=>nx6970);
   gen_regs_10_regi_reg_q_4 : dffr port map ( Q=>q_10_4_EXMPLR, QB=>OPEN, D
      =>nx2833, CLK=>nx7088, R=>reset);
   ix2834 : mux21_ni port map ( Y=>nx2833, A0=>q_10_4_EXMPLR, A1=>
      q_9_4_EXMPLR, S0=>nx6970);
   gen_regs_9_regi_reg_q_4 : dffr port map ( Q=>q_9_4_EXMPLR, QB=>OPEN, D=>
      nx2823, CLK=>nx7088, R=>reset);
   ix2824 : mux21_ni port map ( Y=>nx2823, A0=>q_9_4_EXMPLR, A1=>
      q_8_4_EXMPLR, S0=>nx6970);
   gen_regs_8_regi_reg_q_4 : dffr port map ( Q=>q_8_4_EXMPLR, QB=>OPEN, D=>
      nx2813, CLK=>nx7088, R=>reset);
   ix2814 : mux21_ni port map ( Y=>nx2813, A0=>q_8_4_EXMPLR, A1=>
      q_7_4_EXMPLR, S0=>nx6970);
   gen_regs_7_regi_reg_q_4 : dffr port map ( Q=>q_7_4_EXMPLR, QB=>OPEN, D=>
      nx2803, CLK=>nx7088, R=>reset);
   ix2804 : mux21_ni port map ( Y=>nx2803, A0=>q_7_4_EXMPLR, A1=>
      q_6_4_EXMPLR, S0=>nx6970);
   gen_regs_6_regi_reg_q_4 : dffr port map ( Q=>q_6_4_EXMPLR, QB=>OPEN, D=>
      nx2793, CLK=>nx7088, R=>reset);
   ix2794 : mux21_ni port map ( Y=>nx2793, A0=>q_6_4_EXMPLR, A1=>
      q_5_4_EXMPLR, S0=>nx6970);
   gen_regs_5_regi_reg_q_4 : dffr port map ( Q=>q_5_4_EXMPLR, QB=>OPEN, D=>
      nx2783, CLK=>nx7088, R=>reset);
   ix2784 : mux21_ni port map ( Y=>nx2783, A0=>q_5_4_EXMPLR, A1=>
      q_4_4_EXMPLR, S0=>nx6970);
   gen_regs_4_regi_reg_q_4 : dffr port map ( Q=>q_4_4_EXMPLR, QB=>OPEN, D=>
      nx2773, CLK=>nx7086, R=>reset);
   ix2774 : mux21_ni port map ( Y=>nx2773, A0=>q_4_4_EXMPLR, A1=>
      q_3_4_EXMPLR, S0=>nx6968);
   gen_regs_3_regi_reg_q_4 : dffr port map ( Q=>q_3_4_EXMPLR, QB=>OPEN, D=>
      nx2763, CLK=>nx7086, R=>reset);
   ix2764 : mux21_ni port map ( Y=>nx2763, A0=>q_3_4_EXMPLR, A1=>
      q_2_4_EXMPLR, S0=>nx6968);
   gen_regs_2_regi_reg_q_4 : dffr port map ( Q=>q_2_4_EXMPLR, QB=>OPEN, D=>
      nx2753, CLK=>nx7086, R=>reset);
   ix2754 : mux21_ni port map ( Y=>nx2753, A0=>q_2_4_EXMPLR, A1=>
      q_1_4_EXMPLR, S0=>nx6968);
   gen_regs_1_regi_reg_q_4 : dffr port map ( Q=>q_1_4_EXMPLR, QB=>OPEN, D=>
      nx2743, CLK=>nx7086, R=>reset);
   ix2744 : mux21_ni port map ( Y=>nx2743, A0=>q_1_4_EXMPLR, A1=>
      q_0_4_EXMPLR, S0=>nx6968);
   reg0_reg_q_4 : dffr port map ( Q=>q_0_4_EXMPLR, QB=>OPEN, D=>nx2733, CLK
      =>nx7086, R=>reset);
   ix2734 : mux21_ni port map ( Y=>nx2733, A0=>q_0_4_EXMPLR, A1=>d(4), S0=>
      nx6968);
   gen_regs_24_regi_reg_q_5 : dffr port map ( Q=>q_24_5_EXMPLR, QB=>OPEN, D
      =>nx3223, CLK=>nx7100, R=>reset);
   ix3224 : mux21_ni port map ( Y=>nx3223, A0=>q_24_5_EXMPLR, A1=>
      q_23_5_EXMPLR, S0=>nx6982);
   gen_regs_23_regi_reg_q_5 : dffr port map ( Q=>q_23_5_EXMPLR, QB=>OPEN, D
      =>nx3213, CLK=>nx7100, R=>reset);
   ix3214 : mux21_ni port map ( Y=>nx3213, A0=>q_23_5_EXMPLR, A1=>
      q_22_5_EXMPLR, S0=>nx6982);
   gen_regs_22_regi_reg_q_5 : dffr port map ( Q=>q_22_5_EXMPLR, QB=>OPEN, D
      =>nx3203, CLK=>nx7100, R=>reset);
   ix3204 : mux21_ni port map ( Y=>nx3203, A0=>q_22_5_EXMPLR, A1=>
      q_21_5_EXMPLR, S0=>nx6982);
   gen_regs_21_regi_reg_q_5 : dffr port map ( Q=>q_21_5_EXMPLR, QB=>OPEN, D
      =>nx3193, CLK=>nx7098, R=>reset);
   ix3194 : mux21_ni port map ( Y=>nx3193, A0=>q_21_5_EXMPLR, A1=>
      q_20_5_EXMPLR, S0=>nx6980);
   gen_regs_20_regi_reg_q_5 : dffr port map ( Q=>q_20_5_EXMPLR, QB=>OPEN, D
      =>nx3183, CLK=>nx7098, R=>reset);
   ix3184 : mux21_ni port map ( Y=>nx3183, A0=>q_20_5_EXMPLR, A1=>
      q_19_5_EXMPLR, S0=>nx6980);
   gen_regs_19_regi_reg_q_5 : dffr port map ( Q=>q_19_5_EXMPLR, QB=>OPEN, D
      =>nx3173, CLK=>nx7098, R=>reset);
   ix3174 : mux21_ni port map ( Y=>nx3173, A0=>q_19_5_EXMPLR, A1=>
      q_18_5_EXMPLR, S0=>nx6980);
   gen_regs_18_regi_reg_q_5 : dffr port map ( Q=>q_18_5_EXMPLR, QB=>OPEN, D
      =>nx3163, CLK=>nx7098, R=>reset);
   ix3164 : mux21_ni port map ( Y=>nx3163, A0=>q_18_5_EXMPLR, A1=>
      q_17_5_EXMPLR, S0=>nx6980);
   gen_regs_17_regi_reg_q_5 : dffr port map ( Q=>q_17_5_EXMPLR, QB=>OPEN, D
      =>nx3153, CLK=>nx7098, R=>reset);
   ix3154 : mux21_ni port map ( Y=>nx3153, A0=>q_17_5_EXMPLR, A1=>
      q_16_5_EXMPLR, S0=>nx6980);
   gen_regs_16_regi_reg_q_5 : dffr port map ( Q=>q_16_5_EXMPLR, QB=>OPEN, D
      =>nx3143, CLK=>nx7098, R=>reset);
   ix3144 : mux21_ni port map ( Y=>nx3143, A0=>q_16_5_EXMPLR, A1=>
      q_15_5_EXMPLR, S0=>nx6980);
   gen_regs_15_regi_reg_q_5 : dffr port map ( Q=>q_15_5_EXMPLR, QB=>OPEN, D
      =>nx3133, CLK=>nx7098, R=>reset);
   ix3134 : mux21_ni port map ( Y=>nx3133, A0=>q_15_5_EXMPLR, A1=>
      q_14_5_EXMPLR, S0=>nx6980);
   gen_regs_14_regi_reg_q_5 : dffr port map ( Q=>q_14_5_EXMPLR, QB=>OPEN, D
      =>nx3123, CLK=>nx7096, R=>reset);
   ix3124 : mux21_ni port map ( Y=>nx3123, A0=>q_14_5_EXMPLR, A1=>
      q_13_5_EXMPLR, S0=>nx6978);
   gen_regs_13_regi_reg_q_5 : dffr port map ( Q=>q_13_5_EXMPLR, QB=>OPEN, D
      =>nx3113, CLK=>nx7096, R=>reset);
   ix3114 : mux21_ni port map ( Y=>nx3113, A0=>q_13_5_EXMPLR, A1=>
      q_12_5_EXMPLR, S0=>nx6978);
   gen_regs_12_regi_reg_q_5 : dffr port map ( Q=>q_12_5_EXMPLR, QB=>OPEN, D
      =>nx3103, CLK=>nx7096, R=>reset);
   ix3104 : mux21_ni port map ( Y=>nx3103, A0=>q_12_5_EXMPLR, A1=>
      q_11_5_EXMPLR, S0=>nx6978);
   gen_regs_11_regi_reg_q_5 : dffr port map ( Q=>q_11_5_EXMPLR, QB=>OPEN, D
      =>nx3093, CLK=>nx7096, R=>reset);
   ix3094 : mux21_ni port map ( Y=>nx3093, A0=>q_11_5_EXMPLR, A1=>
      q_10_5_EXMPLR, S0=>nx6978);
   gen_regs_10_regi_reg_q_5 : dffr port map ( Q=>q_10_5_EXMPLR, QB=>OPEN, D
      =>nx3083, CLK=>nx7096, R=>reset);
   ix3084 : mux21_ni port map ( Y=>nx3083, A0=>q_10_5_EXMPLR, A1=>
      q_9_5_EXMPLR, S0=>nx6978);
   gen_regs_9_regi_reg_q_5 : dffr port map ( Q=>q_9_5_EXMPLR, QB=>OPEN, D=>
      nx3073, CLK=>nx7096, R=>reset);
   ix3074 : mux21_ni port map ( Y=>nx3073, A0=>q_9_5_EXMPLR, A1=>
      q_8_5_EXMPLR, S0=>nx6978);
   gen_regs_8_regi_reg_q_5 : dffr port map ( Q=>q_8_5_EXMPLR, QB=>OPEN, D=>
      nx3063, CLK=>nx7096, R=>reset);
   ix3064 : mux21_ni port map ( Y=>nx3063, A0=>q_8_5_EXMPLR, A1=>
      q_7_5_EXMPLR, S0=>nx6978);
   gen_regs_7_regi_reg_q_5 : dffr port map ( Q=>q_7_5_EXMPLR, QB=>OPEN, D=>
      nx3053, CLK=>nx7094, R=>reset);
   ix3054 : mux21_ni port map ( Y=>nx3053, A0=>q_7_5_EXMPLR, A1=>
      q_6_5_EXMPLR, S0=>nx6976);
   gen_regs_6_regi_reg_q_5 : dffr port map ( Q=>q_6_5_EXMPLR, QB=>OPEN, D=>
      nx3043, CLK=>nx7094, R=>reset);
   ix3044 : mux21_ni port map ( Y=>nx3043, A0=>q_6_5_EXMPLR, A1=>
      q_5_5_EXMPLR, S0=>nx6976);
   gen_regs_5_regi_reg_q_5 : dffr port map ( Q=>q_5_5_EXMPLR, QB=>OPEN, D=>
      nx3033, CLK=>nx7094, R=>reset);
   ix3034 : mux21_ni port map ( Y=>nx3033, A0=>q_5_5_EXMPLR, A1=>
      q_4_5_EXMPLR, S0=>nx6976);
   gen_regs_4_regi_reg_q_5 : dffr port map ( Q=>q_4_5_EXMPLR, QB=>OPEN, D=>
      nx3023, CLK=>nx7094, R=>reset);
   ix3024 : mux21_ni port map ( Y=>nx3023, A0=>q_4_5_EXMPLR, A1=>
      q_3_5_EXMPLR, S0=>nx6976);
   gen_regs_3_regi_reg_q_5 : dffr port map ( Q=>q_3_5_EXMPLR, QB=>OPEN, D=>
      nx3013, CLK=>nx7094, R=>reset);
   ix3014 : mux21_ni port map ( Y=>nx3013, A0=>q_3_5_EXMPLR, A1=>
      q_2_5_EXMPLR, S0=>nx6976);
   gen_regs_2_regi_reg_q_5 : dffr port map ( Q=>q_2_5_EXMPLR, QB=>OPEN, D=>
      nx3003, CLK=>nx7094, R=>reset);
   ix3004 : mux21_ni port map ( Y=>nx3003, A0=>q_2_5_EXMPLR, A1=>
      q_1_5_EXMPLR, S0=>nx6976);
   gen_regs_1_regi_reg_q_5 : dffr port map ( Q=>q_1_5_EXMPLR, QB=>OPEN, D=>
      nx2993, CLK=>nx7094, R=>reset);
   ix2994 : mux21_ni port map ( Y=>nx2993, A0=>q_1_5_EXMPLR, A1=>
      q_0_5_EXMPLR, S0=>nx6976);
   reg0_reg_q_5 : dffr port map ( Q=>q_0_5_EXMPLR, QB=>OPEN, D=>nx2983, CLK
      =>nx7092, R=>reset);
   ix2984 : mux21_ni port map ( Y=>nx2983, A0=>q_0_5_EXMPLR, A1=>d(5), S0=>
      nx6974);
   gen_regs_24_regi_reg_q_6 : dffr port map ( Q=>q_24_6_EXMPLR, QB=>OPEN, D
      =>nx3473, CLK=>nx7106, R=>reset);
   ix3474 : mux21_ni port map ( Y=>nx3473, A0=>q_24_6_EXMPLR, A1=>
      q_23_6_EXMPLR, S0=>nx6988);
   gen_regs_23_regi_reg_q_6 : dffr port map ( Q=>q_23_6_EXMPLR, QB=>OPEN, D
      =>nx3463, CLK=>nx7106, R=>reset);
   ix3464 : mux21_ni port map ( Y=>nx3463, A0=>q_23_6_EXMPLR, A1=>
      q_22_6_EXMPLR, S0=>nx6988);
   gen_regs_22_regi_reg_q_6 : dffr port map ( Q=>q_22_6_EXMPLR, QB=>OPEN, D
      =>nx3453, CLK=>nx7106, R=>reset);
   ix3454 : mux21_ni port map ( Y=>nx3453, A0=>q_22_6_EXMPLR, A1=>
      q_21_6_EXMPLR, S0=>nx6988);
   gen_regs_21_regi_reg_q_6 : dffr port map ( Q=>q_21_6_EXMPLR, QB=>OPEN, D
      =>nx3443, CLK=>nx7106, R=>reset);
   ix3444 : mux21_ni port map ( Y=>nx3443, A0=>q_21_6_EXMPLR, A1=>
      q_20_6_EXMPLR, S0=>nx6988);
   gen_regs_20_regi_reg_q_6 : dffr port map ( Q=>q_20_6_EXMPLR, QB=>OPEN, D
      =>nx3433, CLK=>nx7106, R=>reset);
   ix3434 : mux21_ni port map ( Y=>nx3433, A0=>q_20_6_EXMPLR, A1=>
      q_19_6_EXMPLR, S0=>nx6988);
   gen_regs_19_regi_reg_q_6 : dffr port map ( Q=>q_19_6_EXMPLR, QB=>OPEN, D
      =>nx3423, CLK=>nx7106, R=>reset);
   ix3424 : mux21_ni port map ( Y=>nx3423, A0=>q_19_6_EXMPLR, A1=>
      q_18_6_EXMPLR, S0=>nx6988);
   gen_regs_18_regi_reg_q_6 : dffr port map ( Q=>q_18_6_EXMPLR, QB=>OPEN, D
      =>nx3413, CLK=>nx7106, R=>reset);
   ix3414 : mux21_ni port map ( Y=>nx3413, A0=>q_18_6_EXMPLR, A1=>
      q_17_6_EXMPLR, S0=>nx6988);
   gen_regs_17_regi_reg_q_6 : dffr port map ( Q=>q_17_6_EXMPLR, QB=>OPEN, D
      =>nx3403, CLK=>nx7104, R=>reset);
   ix3404 : mux21_ni port map ( Y=>nx3403, A0=>q_17_6_EXMPLR, A1=>
      q_16_6_EXMPLR, S0=>nx6986);
   gen_regs_16_regi_reg_q_6 : dffr port map ( Q=>q_16_6_EXMPLR, QB=>OPEN, D
      =>nx3393, CLK=>nx7104, R=>reset);
   ix3394 : mux21_ni port map ( Y=>nx3393, A0=>q_16_6_EXMPLR, A1=>
      q_15_6_EXMPLR, S0=>nx6986);
   gen_regs_15_regi_reg_q_6 : dffr port map ( Q=>q_15_6_EXMPLR, QB=>OPEN, D
      =>nx3383, CLK=>nx7104, R=>reset);
   ix3384 : mux21_ni port map ( Y=>nx3383, A0=>q_15_6_EXMPLR, A1=>
      q_14_6_EXMPLR, S0=>nx6986);
   gen_regs_14_regi_reg_q_6 : dffr port map ( Q=>q_14_6_EXMPLR, QB=>OPEN, D
      =>nx3373, CLK=>nx7104, R=>reset);
   ix3374 : mux21_ni port map ( Y=>nx3373, A0=>q_14_6_EXMPLR, A1=>
      q_13_6_EXMPLR, S0=>nx6986);
   gen_regs_13_regi_reg_q_6 : dffr port map ( Q=>q_13_6_EXMPLR, QB=>OPEN, D
      =>nx3363, CLK=>nx7104, R=>reset);
   ix3364 : mux21_ni port map ( Y=>nx3363, A0=>q_13_6_EXMPLR, A1=>
      q_12_6_EXMPLR, S0=>nx6986);
   gen_regs_12_regi_reg_q_6 : dffr port map ( Q=>q_12_6_EXMPLR, QB=>OPEN, D
      =>nx3353, CLK=>nx7104, R=>reset);
   ix3354 : mux21_ni port map ( Y=>nx3353, A0=>q_12_6_EXMPLR, A1=>
      q_11_6_EXMPLR, S0=>nx6986);
   gen_regs_11_regi_reg_q_6 : dffr port map ( Q=>q_11_6_EXMPLR, QB=>OPEN, D
      =>nx3343, CLK=>nx7104, R=>reset);
   ix3344 : mux21_ni port map ( Y=>nx3343, A0=>q_11_6_EXMPLR, A1=>
      q_10_6_EXMPLR, S0=>nx6986);
   gen_regs_10_regi_reg_q_6 : dffr port map ( Q=>q_10_6_EXMPLR, QB=>OPEN, D
      =>nx3333, CLK=>nx7102, R=>reset);
   ix3334 : mux21_ni port map ( Y=>nx3333, A0=>q_10_6_EXMPLR, A1=>
      q_9_6_EXMPLR, S0=>nx6984);
   gen_regs_9_regi_reg_q_6 : dffr port map ( Q=>q_9_6_EXMPLR, QB=>OPEN, D=>
      nx3323, CLK=>nx7102, R=>reset);
   ix3324 : mux21_ni port map ( Y=>nx3323, A0=>q_9_6_EXMPLR, A1=>
      q_8_6_EXMPLR, S0=>nx6984);
   gen_regs_8_regi_reg_q_6 : dffr port map ( Q=>q_8_6_EXMPLR, QB=>OPEN, D=>
      nx3313, CLK=>nx7102, R=>reset);
   ix3314 : mux21_ni port map ( Y=>nx3313, A0=>q_8_6_EXMPLR, A1=>
      q_7_6_EXMPLR, S0=>nx6984);
   gen_regs_7_regi_reg_q_6 : dffr port map ( Q=>q_7_6_EXMPLR, QB=>OPEN, D=>
      nx3303, CLK=>nx7102, R=>reset);
   ix3304 : mux21_ni port map ( Y=>nx3303, A0=>q_7_6_EXMPLR, A1=>
      q_6_6_EXMPLR, S0=>nx6984);
   gen_regs_6_regi_reg_q_6 : dffr port map ( Q=>q_6_6_EXMPLR, QB=>OPEN, D=>
      nx3293, CLK=>nx7102, R=>reset);
   ix3294 : mux21_ni port map ( Y=>nx3293, A0=>q_6_6_EXMPLR, A1=>
      q_5_6_EXMPLR, S0=>nx6984);
   gen_regs_5_regi_reg_q_6 : dffr port map ( Q=>q_5_6_EXMPLR, QB=>OPEN, D=>
      nx3283, CLK=>nx7102, R=>reset);
   ix3284 : mux21_ni port map ( Y=>nx3283, A0=>q_5_6_EXMPLR, A1=>
      q_4_6_EXMPLR, S0=>nx6984);
   gen_regs_4_regi_reg_q_6 : dffr port map ( Q=>q_4_6_EXMPLR, QB=>OPEN, D=>
      nx3273, CLK=>nx7102, R=>reset);
   ix3274 : mux21_ni port map ( Y=>nx3273, A0=>q_4_6_EXMPLR, A1=>
      q_3_6_EXMPLR, S0=>nx6984);
   gen_regs_3_regi_reg_q_6 : dffr port map ( Q=>q_3_6_EXMPLR, QB=>OPEN, D=>
      nx3263, CLK=>nx7100, R=>reset);
   ix3264 : mux21_ni port map ( Y=>nx3263, A0=>q_3_6_EXMPLR, A1=>
      q_2_6_EXMPLR, S0=>nx6982);
   gen_regs_2_regi_reg_q_6 : dffr port map ( Q=>q_2_6_EXMPLR, QB=>OPEN, D=>
      nx3253, CLK=>nx7100, R=>reset);
   ix3254 : mux21_ni port map ( Y=>nx3253, A0=>q_2_6_EXMPLR, A1=>
      q_1_6_EXMPLR, S0=>nx6982);
   gen_regs_1_regi_reg_q_6 : dffr port map ( Q=>q_1_6_EXMPLR, QB=>OPEN, D=>
      nx3243, CLK=>nx7100, R=>reset);
   ix3244 : mux21_ni port map ( Y=>nx3243, A0=>q_1_6_EXMPLR, A1=>
      q_0_6_EXMPLR, S0=>nx6982);
   reg0_reg_q_6 : dffr port map ( Q=>q_0_6_EXMPLR, QB=>OPEN, D=>nx3233, CLK
      =>nx7100, R=>reset);
   ix3234 : mux21_ni port map ( Y=>nx3233, A0=>q_0_6_EXMPLR, A1=>d(6), S0=>
      nx6982);
   gen_regs_24_regi_reg_q_7 : dffr port map ( Q=>q_24_7_EXMPLR, QB=>OPEN, D
      =>nx3723, CLK=>nx7114, R=>reset);
   ix3724 : mux21_ni port map ( Y=>nx3723, A0=>q_24_7_EXMPLR, A1=>
      q_23_7_EXMPLR, S0=>nx6996);
   gen_regs_23_regi_reg_q_7 : dffr port map ( Q=>q_23_7_EXMPLR, QB=>OPEN, D
      =>nx3713, CLK=>nx7114, R=>reset);
   ix3714 : mux21_ni port map ( Y=>nx3713, A0=>q_23_7_EXMPLR, A1=>
      q_22_7_EXMPLR, S0=>nx6996);
   gen_regs_22_regi_reg_q_7 : dffr port map ( Q=>q_22_7_EXMPLR, QB=>OPEN, D
      =>nx3703, CLK=>nx7114, R=>reset);
   ix3704 : mux21_ni port map ( Y=>nx3703, A0=>q_22_7_EXMPLR, A1=>
      q_21_7_EXMPLR, S0=>nx6996);
   gen_regs_21_regi_reg_q_7 : dffr port map ( Q=>q_21_7_EXMPLR, QB=>OPEN, D
      =>nx3693, CLK=>nx7114, R=>reset);
   ix3694 : mux21_ni port map ( Y=>nx3693, A0=>q_21_7_EXMPLR, A1=>
      q_20_7_EXMPLR, S0=>nx6996);
   gen_regs_20_regi_reg_q_7 : dffr port map ( Q=>q_20_7_EXMPLR, QB=>OPEN, D
      =>nx3683, CLK=>nx7112, R=>reset);
   ix3684 : mux21_ni port map ( Y=>nx3683, A0=>q_20_7_EXMPLR, A1=>
      q_19_7_EXMPLR, S0=>nx6994);
   gen_regs_19_regi_reg_q_7 : dffr port map ( Q=>q_19_7_EXMPLR, QB=>OPEN, D
      =>nx3673, CLK=>nx7112, R=>reset);
   ix3674 : mux21_ni port map ( Y=>nx3673, A0=>q_19_7_EXMPLR, A1=>
      q_18_7_EXMPLR, S0=>nx6994);
   gen_regs_18_regi_reg_q_7 : dffr port map ( Q=>q_18_7_EXMPLR, QB=>OPEN, D
      =>nx3663, CLK=>nx7112, R=>reset);
   ix3664 : mux21_ni port map ( Y=>nx3663, A0=>q_18_7_EXMPLR, A1=>
      q_17_7_EXMPLR, S0=>nx6994);
   gen_regs_17_regi_reg_q_7 : dffr port map ( Q=>q_17_7_EXMPLR, QB=>OPEN, D
      =>nx3653, CLK=>nx7112, R=>reset);
   ix3654 : mux21_ni port map ( Y=>nx3653, A0=>q_17_7_EXMPLR, A1=>
      q_16_7_EXMPLR, S0=>nx6994);
   gen_regs_16_regi_reg_q_7 : dffr port map ( Q=>q_16_7_EXMPLR, QB=>OPEN, D
      =>nx3643, CLK=>nx7112, R=>reset);
   ix3644 : mux21_ni port map ( Y=>nx3643, A0=>q_16_7_EXMPLR, A1=>
      q_15_7_EXMPLR, S0=>nx6994);
   gen_regs_15_regi_reg_q_7 : dffr port map ( Q=>q_15_7_EXMPLR, QB=>OPEN, D
      =>nx3633, CLK=>nx7112, R=>reset);
   ix3634 : mux21_ni port map ( Y=>nx3633, A0=>q_15_7_EXMPLR, A1=>
      q_14_7_EXMPLR, S0=>nx6994);
   gen_regs_14_regi_reg_q_7 : dffr port map ( Q=>q_14_7_EXMPLR, QB=>OPEN, D
      =>nx3623, CLK=>nx7112, R=>reset);
   ix3624 : mux21_ni port map ( Y=>nx3623, A0=>q_14_7_EXMPLR, A1=>
      q_13_7_EXMPLR, S0=>nx6994);
   gen_regs_13_regi_reg_q_7 : dffr port map ( Q=>q_13_7_EXMPLR, QB=>OPEN, D
      =>nx3613, CLK=>nx7110, R=>reset);
   ix3614 : mux21_ni port map ( Y=>nx3613, A0=>q_13_7_EXMPLR, A1=>
      q_12_7_EXMPLR, S0=>nx6992);
   gen_regs_12_regi_reg_q_7 : dffr port map ( Q=>q_12_7_EXMPLR, QB=>OPEN, D
      =>nx3603, CLK=>nx7110, R=>reset);
   ix3604 : mux21_ni port map ( Y=>nx3603, A0=>q_12_7_EXMPLR, A1=>
      q_11_7_EXMPLR, S0=>nx6992);
   gen_regs_11_regi_reg_q_7 : dffr port map ( Q=>q_11_7_EXMPLR, QB=>OPEN, D
      =>nx3593, CLK=>nx7110, R=>reset);
   ix3594 : mux21_ni port map ( Y=>nx3593, A0=>q_11_7_EXMPLR, A1=>
      q_10_7_EXMPLR, S0=>nx6992);
   gen_regs_10_regi_reg_q_7 : dffr port map ( Q=>q_10_7_EXMPLR, QB=>OPEN, D
      =>nx3583, CLK=>nx7110, R=>reset);
   ix3584 : mux21_ni port map ( Y=>nx3583, A0=>q_10_7_EXMPLR, A1=>
      q_9_7_EXMPLR, S0=>nx6992);
   gen_regs_9_regi_reg_q_7 : dffr port map ( Q=>q_9_7_EXMPLR, QB=>OPEN, D=>
      nx3573, CLK=>nx7110, R=>reset);
   ix3574 : mux21_ni port map ( Y=>nx3573, A0=>q_9_7_EXMPLR, A1=>
      q_8_7_EXMPLR, S0=>nx6992);
   gen_regs_8_regi_reg_q_7 : dffr port map ( Q=>q_8_7_EXMPLR, QB=>OPEN, D=>
      nx3563, CLK=>nx7110, R=>reset);
   ix3564 : mux21_ni port map ( Y=>nx3563, A0=>q_8_7_EXMPLR, A1=>
      q_7_7_EXMPLR, S0=>nx6992);
   gen_regs_7_regi_reg_q_7 : dffr port map ( Q=>q_7_7_EXMPLR, QB=>OPEN, D=>
      nx3553, CLK=>nx7110, R=>reset);
   ix3554 : mux21_ni port map ( Y=>nx3553, A0=>q_7_7_EXMPLR, A1=>
      q_6_7_EXMPLR, S0=>nx6992);
   gen_regs_6_regi_reg_q_7 : dffr port map ( Q=>q_6_7_EXMPLR, QB=>OPEN, D=>
      nx3543, CLK=>nx7108, R=>reset);
   ix3544 : mux21_ni port map ( Y=>nx3543, A0=>q_6_7_EXMPLR, A1=>
      q_5_7_EXMPLR, S0=>nx6990);
   gen_regs_5_regi_reg_q_7 : dffr port map ( Q=>q_5_7_EXMPLR, QB=>OPEN, D=>
      nx3533, CLK=>nx7108, R=>reset);
   ix3534 : mux21_ni port map ( Y=>nx3533, A0=>q_5_7_EXMPLR, A1=>
      q_4_7_EXMPLR, S0=>nx6990);
   gen_regs_4_regi_reg_q_7 : dffr port map ( Q=>q_4_7_EXMPLR, QB=>OPEN, D=>
      nx3523, CLK=>nx7108, R=>reset);
   ix3524 : mux21_ni port map ( Y=>nx3523, A0=>q_4_7_EXMPLR, A1=>
      q_3_7_EXMPLR, S0=>nx6990);
   gen_regs_3_regi_reg_q_7 : dffr port map ( Q=>q_3_7_EXMPLR, QB=>OPEN, D=>
      nx3513, CLK=>nx7108, R=>reset);
   ix3514 : mux21_ni port map ( Y=>nx3513, A0=>q_3_7_EXMPLR, A1=>
      q_2_7_EXMPLR, S0=>nx6990);
   gen_regs_2_regi_reg_q_7 : dffr port map ( Q=>q_2_7_EXMPLR, QB=>OPEN, D=>
      nx3503, CLK=>nx7108, R=>reset);
   ix3504 : mux21_ni port map ( Y=>nx3503, A0=>q_2_7_EXMPLR, A1=>
      q_1_7_EXMPLR, S0=>nx6990);
   gen_regs_1_regi_reg_q_7 : dffr port map ( Q=>q_1_7_EXMPLR, QB=>OPEN, D=>
      nx3493, CLK=>nx7108, R=>reset);
   ix3494 : mux21_ni port map ( Y=>nx3493, A0=>q_1_7_EXMPLR, A1=>
      q_0_7_EXMPLR, S0=>nx6990);
   reg0_reg_q_7 : dffr port map ( Q=>q_0_7_EXMPLR, QB=>OPEN, D=>nx3483, CLK
      =>nx7108, R=>reset);
   ix3484 : mux21_ni port map ( Y=>nx3483, A0=>q_0_7_EXMPLR, A1=>d(7), S0=>
      nx6990);
   gen_regs_24_regi_reg_q_8 : dffr port map ( Q=>q_24_8_EXMPLR, QB=>OPEN, D
      =>nx3973, CLK=>nx7122, R=>reset);
   ix3974 : mux21_ni port map ( Y=>nx3973, A0=>q_24_8_EXMPLR, A1=>
      q_23_8_EXMPLR, S0=>nx7004);
   gen_regs_23_regi_reg_q_8 : dffr port map ( Q=>q_23_8_EXMPLR, QB=>OPEN, D
      =>nx3963, CLK=>nx7120, R=>reset);
   ix3964 : mux21_ni port map ( Y=>nx3963, A0=>q_23_8_EXMPLR, A1=>
      q_22_8_EXMPLR, S0=>nx7002);
   gen_regs_22_regi_reg_q_8 : dffr port map ( Q=>q_22_8_EXMPLR, QB=>OPEN, D
      =>nx3953, CLK=>nx7120, R=>reset);
   ix3954 : mux21_ni port map ( Y=>nx3953, A0=>q_22_8_EXMPLR, A1=>
      q_21_8_EXMPLR, S0=>nx7002);
   gen_regs_21_regi_reg_q_8 : dffr port map ( Q=>q_21_8_EXMPLR, QB=>OPEN, D
      =>nx3943, CLK=>nx7120, R=>reset);
   ix3944 : mux21_ni port map ( Y=>nx3943, A0=>q_21_8_EXMPLR, A1=>
      q_20_8_EXMPLR, S0=>nx7002);
   gen_regs_20_regi_reg_q_8 : dffr port map ( Q=>q_20_8_EXMPLR, QB=>OPEN, D
      =>nx3933, CLK=>nx7120, R=>reset);
   ix3934 : mux21_ni port map ( Y=>nx3933, A0=>q_20_8_EXMPLR, A1=>
      q_19_8_EXMPLR, S0=>nx7002);
   gen_regs_19_regi_reg_q_8 : dffr port map ( Q=>q_19_8_EXMPLR, QB=>OPEN, D
      =>nx3923, CLK=>nx7120, R=>reset);
   ix3924 : mux21_ni port map ( Y=>nx3923, A0=>q_19_8_EXMPLR, A1=>
      q_18_8_EXMPLR, S0=>nx7002);
   gen_regs_18_regi_reg_q_8 : dffr port map ( Q=>q_18_8_EXMPLR, QB=>OPEN, D
      =>nx3913, CLK=>nx7120, R=>reset);
   ix3914 : mux21_ni port map ( Y=>nx3913, A0=>q_18_8_EXMPLR, A1=>
      q_17_8_EXMPLR, S0=>nx7002);
   gen_regs_17_regi_reg_q_8 : dffr port map ( Q=>q_17_8_EXMPLR, QB=>OPEN, D
      =>nx3903, CLK=>nx7120, R=>reset);
   ix3904 : mux21_ni port map ( Y=>nx3903, A0=>q_17_8_EXMPLR, A1=>
      q_16_8_EXMPLR, S0=>nx7002);
   gen_regs_16_regi_reg_q_8 : dffr port map ( Q=>q_16_8_EXMPLR, QB=>OPEN, D
      =>nx3893, CLK=>nx7118, R=>reset);
   ix3894 : mux21_ni port map ( Y=>nx3893, A0=>q_16_8_EXMPLR, A1=>
      q_15_8_EXMPLR, S0=>nx7000);
   gen_regs_15_regi_reg_q_8 : dffr port map ( Q=>q_15_8_EXMPLR, QB=>OPEN, D
      =>nx3883, CLK=>nx7118, R=>reset);
   ix3884 : mux21_ni port map ( Y=>nx3883, A0=>q_15_8_EXMPLR, A1=>
      q_14_8_EXMPLR, S0=>nx7000);
   gen_regs_14_regi_reg_q_8 : dffr port map ( Q=>q_14_8_EXMPLR, QB=>OPEN, D
      =>nx3873, CLK=>nx7118, R=>reset);
   ix3874 : mux21_ni port map ( Y=>nx3873, A0=>q_14_8_EXMPLR, A1=>
      q_13_8_EXMPLR, S0=>nx7000);
   gen_regs_13_regi_reg_q_8 : dffr port map ( Q=>q_13_8_EXMPLR, QB=>OPEN, D
      =>nx3863, CLK=>nx7118, R=>reset);
   ix3864 : mux21_ni port map ( Y=>nx3863, A0=>q_13_8_EXMPLR, A1=>
      q_12_8_EXMPLR, S0=>nx7000);
   gen_regs_12_regi_reg_q_8 : dffr port map ( Q=>q_12_8_EXMPLR, QB=>OPEN, D
      =>nx3853, CLK=>nx7118, R=>reset);
   ix3854 : mux21_ni port map ( Y=>nx3853, A0=>q_12_8_EXMPLR, A1=>
      q_11_8_EXMPLR, S0=>nx7000);
   gen_regs_11_regi_reg_q_8 : dffr port map ( Q=>q_11_8_EXMPLR, QB=>OPEN, D
      =>nx3843, CLK=>nx7118, R=>reset);
   ix3844 : mux21_ni port map ( Y=>nx3843, A0=>q_11_8_EXMPLR, A1=>
      q_10_8_EXMPLR, S0=>nx7000);
   gen_regs_10_regi_reg_q_8 : dffr port map ( Q=>q_10_8_EXMPLR, QB=>OPEN, D
      =>nx3833, CLK=>nx7118, R=>reset);
   ix3834 : mux21_ni port map ( Y=>nx3833, A0=>q_10_8_EXMPLR, A1=>
      q_9_8_EXMPLR, S0=>nx7000);
   gen_regs_9_regi_reg_q_8 : dffr port map ( Q=>q_9_8_EXMPLR, QB=>OPEN, D=>
      nx3823, CLK=>nx7116, R=>reset);
   ix3824 : mux21_ni port map ( Y=>nx3823, A0=>q_9_8_EXMPLR, A1=>
      q_8_8_EXMPLR, S0=>nx6998);
   gen_regs_8_regi_reg_q_8 : dffr port map ( Q=>q_8_8_EXMPLR, QB=>OPEN, D=>
      nx3813, CLK=>nx7116, R=>reset);
   ix3814 : mux21_ni port map ( Y=>nx3813, A0=>q_8_8_EXMPLR, A1=>
      q_7_8_EXMPLR, S0=>nx6998);
   gen_regs_7_regi_reg_q_8 : dffr port map ( Q=>q_7_8_EXMPLR, QB=>OPEN, D=>
      nx3803, CLK=>nx7116, R=>reset);
   ix3804 : mux21_ni port map ( Y=>nx3803, A0=>q_7_8_EXMPLR, A1=>
      q_6_8_EXMPLR, S0=>nx6998);
   gen_regs_6_regi_reg_q_8 : dffr port map ( Q=>q_6_8_EXMPLR, QB=>OPEN, D=>
      nx3793, CLK=>nx7116, R=>reset);
   ix3794 : mux21_ni port map ( Y=>nx3793, A0=>q_6_8_EXMPLR, A1=>
      q_5_8_EXMPLR, S0=>nx6998);
   gen_regs_5_regi_reg_q_8 : dffr port map ( Q=>q_5_8_EXMPLR, QB=>OPEN, D=>
      nx3783, CLK=>nx7116, R=>reset);
   ix3784 : mux21_ni port map ( Y=>nx3783, A0=>q_5_8_EXMPLR, A1=>
      q_4_8_EXMPLR, S0=>nx6998);
   gen_regs_4_regi_reg_q_8 : dffr port map ( Q=>q_4_8_EXMPLR, QB=>OPEN, D=>
      nx3773, CLK=>nx7116, R=>reset);
   ix3774 : mux21_ni port map ( Y=>nx3773, A0=>q_4_8_EXMPLR, A1=>
      q_3_8_EXMPLR, S0=>nx6998);
   gen_regs_3_regi_reg_q_8 : dffr port map ( Q=>q_3_8_EXMPLR, QB=>OPEN, D=>
      nx3763, CLK=>nx7116, R=>reset);
   ix3764 : mux21_ni port map ( Y=>nx3763, A0=>q_3_8_EXMPLR, A1=>
      q_2_8_EXMPLR, S0=>nx6998);
   gen_regs_2_regi_reg_q_8 : dffr port map ( Q=>q_2_8_EXMPLR, QB=>OPEN, D=>
      nx3753, CLK=>nx7114, R=>reset);
   ix3754 : mux21_ni port map ( Y=>nx3753, A0=>q_2_8_EXMPLR, A1=>
      q_1_8_EXMPLR, S0=>nx6996);
   gen_regs_1_regi_reg_q_8 : dffr port map ( Q=>q_1_8_EXMPLR, QB=>OPEN, D=>
      nx3743, CLK=>nx7114, R=>reset);
   ix3744 : mux21_ni port map ( Y=>nx3743, A0=>q_1_8_EXMPLR, A1=>
      q_0_8_EXMPLR, S0=>nx6996);
   reg0_reg_q_8 : dffr port map ( Q=>q_0_8_EXMPLR, QB=>OPEN, D=>nx3733, CLK
      =>nx7114, R=>reset);
   ix3734 : mux21_ni port map ( Y=>nx3733, A0=>q_0_8_EXMPLR, A1=>d(8), S0=>
      nx6996);
   gen_regs_24_regi_reg_q_9 : dffr port map ( Q=>q_24_9_EXMPLR, QB=>OPEN, D
      =>nx4223, CLK=>nx7128, R=>reset);
   ix4224 : mux21_ni port map ( Y=>nx4223, A0=>q_24_9_EXMPLR, A1=>
      q_23_9_EXMPLR, S0=>nx7010);
   gen_regs_23_regi_reg_q_9 : dffr port map ( Q=>q_23_9_EXMPLR, QB=>OPEN, D
      =>nx4213, CLK=>nx7128, R=>reset);
   ix4214 : mux21_ni port map ( Y=>nx4213, A0=>q_23_9_EXMPLR, A1=>
      q_22_9_EXMPLR, S0=>nx7010);
   gen_regs_22_regi_reg_q_9 : dffr port map ( Q=>q_22_9_EXMPLR, QB=>OPEN, D
      =>nx4203, CLK=>nx7128, R=>reset);
   ix4204 : mux21_ni port map ( Y=>nx4203, A0=>q_22_9_EXMPLR, A1=>
      q_21_9_EXMPLR, S0=>nx7010);
   gen_regs_21_regi_reg_q_9 : dffr port map ( Q=>q_21_9_EXMPLR, QB=>OPEN, D
      =>nx4193, CLK=>nx7128, R=>reset);
   ix4194 : mux21_ni port map ( Y=>nx4193, A0=>q_21_9_EXMPLR, A1=>
      q_20_9_EXMPLR, S0=>nx7010);
   gen_regs_20_regi_reg_q_9 : dffr port map ( Q=>q_20_9_EXMPLR, QB=>OPEN, D
      =>nx4183, CLK=>nx7128, R=>reset);
   ix4184 : mux21_ni port map ( Y=>nx4183, A0=>q_20_9_EXMPLR, A1=>
      q_19_9_EXMPLR, S0=>nx7010);
   gen_regs_19_regi_reg_q_9 : dffr port map ( Q=>q_19_9_EXMPLR, QB=>OPEN, D
      =>nx4173, CLK=>nx7126, R=>reset);
   ix4174 : mux21_ni port map ( Y=>nx4173, A0=>q_19_9_EXMPLR, A1=>
      q_18_9_EXMPLR, S0=>nx7008);
   gen_regs_18_regi_reg_q_9 : dffr port map ( Q=>q_18_9_EXMPLR, QB=>OPEN, D
      =>nx4163, CLK=>nx7126, R=>reset);
   ix4164 : mux21_ni port map ( Y=>nx4163, A0=>q_18_9_EXMPLR, A1=>
      q_17_9_EXMPLR, S0=>nx7008);
   gen_regs_17_regi_reg_q_9 : dffr port map ( Q=>q_17_9_EXMPLR, QB=>OPEN, D
      =>nx4153, CLK=>nx7126, R=>reset);
   ix4154 : mux21_ni port map ( Y=>nx4153, A0=>q_17_9_EXMPLR, A1=>
      q_16_9_EXMPLR, S0=>nx7008);
   gen_regs_16_regi_reg_q_9 : dffr port map ( Q=>q_16_9_EXMPLR, QB=>OPEN, D
      =>nx4143, CLK=>nx7126, R=>reset);
   ix4144 : mux21_ni port map ( Y=>nx4143, A0=>q_16_9_EXMPLR, A1=>
      q_15_9_EXMPLR, S0=>nx7008);
   gen_regs_15_regi_reg_q_9 : dffr port map ( Q=>q_15_9_EXMPLR, QB=>OPEN, D
      =>nx4133, CLK=>nx7126, R=>reset);
   ix4134 : mux21_ni port map ( Y=>nx4133, A0=>q_15_9_EXMPLR, A1=>
      q_14_9_EXMPLR, S0=>nx7008);
   gen_regs_14_regi_reg_q_9 : dffr port map ( Q=>q_14_9_EXMPLR, QB=>OPEN, D
      =>nx4123, CLK=>nx7126, R=>reset);
   ix4124 : mux21_ni port map ( Y=>nx4123, A0=>q_14_9_EXMPLR, A1=>
      q_13_9_EXMPLR, S0=>nx7008);
   gen_regs_13_regi_reg_q_9 : dffr port map ( Q=>q_13_9_EXMPLR, QB=>OPEN, D
      =>nx4113, CLK=>nx7126, R=>reset);
   ix4114 : mux21_ni port map ( Y=>nx4113, A0=>q_13_9_EXMPLR, A1=>
      q_12_9_EXMPLR, S0=>nx7008);
   gen_regs_12_regi_reg_q_9 : dffr port map ( Q=>q_12_9_EXMPLR, QB=>OPEN, D
      =>nx4103, CLK=>nx7124, R=>reset);
   ix4104 : mux21_ni port map ( Y=>nx4103, A0=>q_12_9_EXMPLR, A1=>
      q_11_9_EXMPLR, S0=>nx7006);
   gen_regs_11_regi_reg_q_9 : dffr port map ( Q=>q_11_9_EXMPLR, QB=>OPEN, D
      =>nx4093, CLK=>nx7124, R=>reset);
   ix4094 : mux21_ni port map ( Y=>nx4093, A0=>q_11_9_EXMPLR, A1=>
      q_10_9_EXMPLR, S0=>nx7006);
   gen_regs_10_regi_reg_q_9 : dffr port map ( Q=>q_10_9_EXMPLR, QB=>OPEN, D
      =>nx4083, CLK=>nx7124, R=>reset);
   ix4084 : mux21_ni port map ( Y=>nx4083, A0=>q_10_9_EXMPLR, A1=>
      q_9_9_EXMPLR, S0=>nx7006);
   gen_regs_9_regi_reg_q_9 : dffr port map ( Q=>q_9_9_EXMPLR, QB=>OPEN, D=>
      nx4073, CLK=>nx7124, R=>reset);
   ix4074 : mux21_ni port map ( Y=>nx4073, A0=>q_9_9_EXMPLR, A1=>
      q_8_9_EXMPLR, S0=>nx7006);
   gen_regs_8_regi_reg_q_9 : dffr port map ( Q=>q_8_9_EXMPLR, QB=>OPEN, D=>
      nx4063, CLK=>nx7124, R=>reset);
   ix4064 : mux21_ni port map ( Y=>nx4063, A0=>q_8_9_EXMPLR, A1=>
      q_7_9_EXMPLR, S0=>nx7006);
   gen_regs_7_regi_reg_q_9 : dffr port map ( Q=>q_7_9_EXMPLR, QB=>OPEN, D=>
      nx4053, CLK=>nx7124, R=>reset);
   ix4054 : mux21_ni port map ( Y=>nx4053, A0=>q_7_9_EXMPLR, A1=>
      q_6_9_EXMPLR, S0=>nx7006);
   gen_regs_6_regi_reg_q_9 : dffr port map ( Q=>q_6_9_EXMPLR, QB=>OPEN, D=>
      nx4043, CLK=>nx7124, R=>reset);
   ix4044 : mux21_ni port map ( Y=>nx4043, A0=>q_6_9_EXMPLR, A1=>
      q_5_9_EXMPLR, S0=>nx7006);
   gen_regs_5_regi_reg_q_9 : dffr port map ( Q=>q_5_9_EXMPLR, QB=>OPEN, D=>
      nx4033, CLK=>nx7122, R=>reset);
   ix4034 : mux21_ni port map ( Y=>nx4033, A0=>q_5_9_EXMPLR, A1=>
      q_4_9_EXMPLR, S0=>nx7004);
   gen_regs_4_regi_reg_q_9 : dffr port map ( Q=>q_4_9_EXMPLR, QB=>OPEN, D=>
      nx4023, CLK=>nx7122, R=>reset);
   ix4024 : mux21_ni port map ( Y=>nx4023, A0=>q_4_9_EXMPLR, A1=>
      q_3_9_EXMPLR, S0=>nx7004);
   gen_regs_3_regi_reg_q_9 : dffr port map ( Q=>q_3_9_EXMPLR, QB=>OPEN, D=>
      nx4013, CLK=>nx7122, R=>reset);
   ix4014 : mux21_ni port map ( Y=>nx4013, A0=>q_3_9_EXMPLR, A1=>
      q_2_9_EXMPLR, S0=>nx7004);
   gen_regs_2_regi_reg_q_9 : dffr port map ( Q=>q_2_9_EXMPLR, QB=>OPEN, D=>
      nx4003, CLK=>nx7122, R=>reset);
   ix4004 : mux21_ni port map ( Y=>nx4003, A0=>q_2_9_EXMPLR, A1=>
      q_1_9_EXMPLR, S0=>nx7004);
   gen_regs_1_regi_reg_q_9 : dffr port map ( Q=>q_1_9_EXMPLR, QB=>OPEN, D=>
      nx3993, CLK=>nx7122, R=>reset);
   ix3994 : mux21_ni port map ( Y=>nx3993, A0=>q_1_9_EXMPLR, A1=>
      q_0_9_EXMPLR, S0=>nx7004);
   reg0_reg_q_9 : dffr port map ( Q=>q_0_9_EXMPLR, QB=>OPEN, D=>nx3983, CLK
      =>nx7122, R=>reset);
   ix3984 : mux21_ni port map ( Y=>nx3983, A0=>q_0_9_EXMPLR, A1=>d(9), S0=>
      nx7004);
   gen_regs_24_regi_reg_q_10 : dffr port map ( Q=>q_24_10_EXMPLR, QB=>OPEN, 
      D=>nx4473, CLK=>nx7136, R=>reset);
   ix4474 : mux21_ni port map ( Y=>nx4473, A0=>q_24_10_EXMPLR, A1=>
      q_23_10_EXMPLR, S0=>nx7018);
   gen_regs_23_regi_reg_q_10 : dffr port map ( Q=>q_23_10_EXMPLR, QB=>OPEN, 
      D=>nx4463, CLK=>nx7136, R=>reset);
   ix4464 : mux21_ni port map ( Y=>nx4463, A0=>q_23_10_EXMPLR, A1=>
      q_22_10_EXMPLR, S0=>nx7018);
   gen_regs_22_regi_reg_q_10 : dffr port map ( Q=>q_22_10_EXMPLR, QB=>OPEN, 
      D=>nx4453, CLK=>nx7134, R=>reset);
   ix4454 : mux21_ni port map ( Y=>nx4453, A0=>q_22_10_EXMPLR, A1=>
      q_21_10_EXMPLR, S0=>nx7016);
   gen_regs_21_regi_reg_q_10 : dffr port map ( Q=>q_21_10_EXMPLR, QB=>OPEN, 
      D=>nx4443, CLK=>nx7134, R=>reset);
   ix4444 : mux21_ni port map ( Y=>nx4443, A0=>q_21_10_EXMPLR, A1=>
      q_20_10_EXMPLR, S0=>nx7016);
   gen_regs_20_regi_reg_q_10 : dffr port map ( Q=>q_20_10_EXMPLR, QB=>OPEN, 
      D=>nx4433, CLK=>nx7134, R=>reset);
   ix4434 : mux21_ni port map ( Y=>nx4433, A0=>q_20_10_EXMPLR, A1=>
      q_19_10_EXMPLR, S0=>nx7016);
   gen_regs_19_regi_reg_q_10 : dffr port map ( Q=>q_19_10_EXMPLR, QB=>OPEN, 
      D=>nx4423, CLK=>nx7134, R=>reset);
   ix4424 : mux21_ni port map ( Y=>nx4423, A0=>q_19_10_EXMPLR, A1=>
      q_18_10_EXMPLR, S0=>nx7016);
   gen_regs_18_regi_reg_q_10 : dffr port map ( Q=>q_18_10_EXMPLR, QB=>OPEN, 
      D=>nx4413, CLK=>nx7134, R=>reset);
   ix4414 : mux21_ni port map ( Y=>nx4413, A0=>q_18_10_EXMPLR, A1=>
      q_17_10_EXMPLR, S0=>nx7016);
   gen_regs_17_regi_reg_q_10 : dffr port map ( Q=>q_17_10_EXMPLR, QB=>OPEN, 
      D=>nx4403, CLK=>nx7134, R=>reset);
   ix4404 : mux21_ni port map ( Y=>nx4403, A0=>q_17_10_EXMPLR, A1=>
      q_16_10_EXMPLR, S0=>nx7016);
   gen_regs_16_regi_reg_q_10 : dffr port map ( Q=>q_16_10_EXMPLR, QB=>OPEN, 
      D=>nx4393, CLK=>nx7134, R=>reset);
   ix4394 : mux21_ni port map ( Y=>nx4393, A0=>q_16_10_EXMPLR, A1=>
      q_15_10_EXMPLR, S0=>nx7016);
   gen_regs_15_regi_reg_q_10 : dffr port map ( Q=>q_15_10_EXMPLR, QB=>OPEN, 
      D=>nx4383, CLK=>nx7132, R=>reset);
   ix4384 : mux21_ni port map ( Y=>nx4383, A0=>q_15_10_EXMPLR, A1=>
      q_14_10_EXMPLR, S0=>nx7014);
   gen_regs_14_regi_reg_q_10 : dffr port map ( Q=>q_14_10_EXMPLR, QB=>OPEN, 
      D=>nx4373, CLK=>nx7132, R=>reset);
   ix4374 : mux21_ni port map ( Y=>nx4373, A0=>q_14_10_EXMPLR, A1=>
      q_13_10_EXMPLR, S0=>nx7014);
   gen_regs_13_regi_reg_q_10 : dffr port map ( Q=>q_13_10_EXMPLR, QB=>OPEN, 
      D=>nx4363, CLK=>nx7132, R=>reset);
   ix4364 : mux21_ni port map ( Y=>nx4363, A0=>q_13_10_EXMPLR, A1=>
      q_12_10_EXMPLR, S0=>nx7014);
   gen_regs_12_regi_reg_q_10 : dffr port map ( Q=>q_12_10_EXMPLR, QB=>OPEN, 
      D=>nx4353, CLK=>nx7132, R=>reset);
   ix4354 : mux21_ni port map ( Y=>nx4353, A0=>q_12_10_EXMPLR, A1=>
      q_11_10_EXMPLR, S0=>nx7014);
   gen_regs_11_regi_reg_q_10 : dffr port map ( Q=>q_11_10_EXMPLR, QB=>OPEN, 
      D=>nx4343, CLK=>nx7132, R=>reset);
   ix4344 : mux21_ni port map ( Y=>nx4343, A0=>q_11_10_EXMPLR, A1=>
      q_10_10_EXMPLR, S0=>nx7014);
   gen_regs_10_regi_reg_q_10 : dffr port map ( Q=>q_10_10_EXMPLR, QB=>OPEN, 
      D=>nx4333, CLK=>nx7132, R=>reset);
   ix4334 : mux21_ni port map ( Y=>nx4333, A0=>q_10_10_EXMPLR, A1=>
      q_9_10_EXMPLR, S0=>nx7014);
   gen_regs_9_regi_reg_q_10 : dffr port map ( Q=>q_9_10_EXMPLR, QB=>OPEN, D
      =>nx4323, CLK=>nx7132, R=>reset);
   ix4324 : mux21_ni port map ( Y=>nx4323, A0=>q_9_10_EXMPLR, A1=>
      q_8_10_EXMPLR, S0=>nx7014);
   gen_regs_8_regi_reg_q_10 : dffr port map ( Q=>q_8_10_EXMPLR, QB=>OPEN, D
      =>nx4313, CLK=>nx7130, R=>reset);
   ix4314 : mux21_ni port map ( Y=>nx4313, A0=>q_8_10_EXMPLR, A1=>
      q_7_10_EXMPLR, S0=>nx7012);
   gen_regs_7_regi_reg_q_10 : dffr port map ( Q=>q_7_10_EXMPLR, QB=>OPEN, D
      =>nx4303, CLK=>nx7130, R=>reset);
   ix4304 : mux21_ni port map ( Y=>nx4303, A0=>q_7_10_EXMPLR, A1=>
      q_6_10_EXMPLR, S0=>nx7012);
   gen_regs_6_regi_reg_q_10 : dffr port map ( Q=>q_6_10_EXMPLR, QB=>OPEN, D
      =>nx4293, CLK=>nx7130, R=>reset);
   ix4294 : mux21_ni port map ( Y=>nx4293, A0=>q_6_10_EXMPLR, A1=>
      q_5_10_EXMPLR, S0=>nx7012);
   gen_regs_5_regi_reg_q_10 : dffr port map ( Q=>q_5_10_EXMPLR, QB=>OPEN, D
      =>nx4283, CLK=>nx7130, R=>reset);
   ix4284 : mux21_ni port map ( Y=>nx4283, A0=>q_5_10_EXMPLR, A1=>
      q_4_10_EXMPLR, S0=>nx7012);
   gen_regs_4_regi_reg_q_10 : dffr port map ( Q=>q_4_10_EXMPLR, QB=>OPEN, D
      =>nx4273, CLK=>nx7130, R=>reset);
   ix4274 : mux21_ni port map ( Y=>nx4273, A0=>q_4_10_EXMPLR, A1=>
      q_3_10_EXMPLR, S0=>nx7012);
   gen_regs_3_regi_reg_q_10 : dffr port map ( Q=>q_3_10_EXMPLR, QB=>OPEN, D
      =>nx4263, CLK=>nx7130, R=>reset);
   ix4264 : mux21_ni port map ( Y=>nx4263, A0=>q_3_10_EXMPLR, A1=>
      q_2_10_EXMPLR, S0=>nx7012);
   gen_regs_2_regi_reg_q_10 : dffr port map ( Q=>q_2_10_EXMPLR, QB=>OPEN, D
      =>nx4253, CLK=>nx7130, R=>reset);
   ix4254 : mux21_ni port map ( Y=>nx4253, A0=>q_2_10_EXMPLR, A1=>
      q_1_10_EXMPLR, S0=>nx7012);
   gen_regs_1_regi_reg_q_10 : dffr port map ( Q=>q_1_10_EXMPLR, QB=>OPEN, D
      =>nx4243, CLK=>nx7128, R=>reset);
   ix4244 : mux21_ni port map ( Y=>nx4243, A0=>q_1_10_EXMPLR, A1=>
      q_0_10_EXMPLR, S0=>nx7010);
   reg0_reg_q_10 : dffr port map ( Q=>q_0_10_EXMPLR, QB=>OPEN, D=>nx4233, 
      CLK=>nx7128, R=>reset);
   ix4234 : mux21_ni port map ( Y=>nx4233, A0=>q_0_10_EXMPLR, A1=>d(10), S0
      =>nx7010);
   gen_regs_24_regi_reg_q_11 : dffr port map ( Q=>q_24_11_EXMPLR, QB=>OPEN, 
      D=>nx4723, CLK=>nx7142, R=>reset);
   ix4724 : mux21_ni port map ( Y=>nx4723, A0=>q_24_11_EXMPLR, A1=>
      q_23_11_EXMPLR, S0=>nx7024);
   gen_regs_23_regi_reg_q_11 : dffr port map ( Q=>q_23_11_EXMPLR, QB=>OPEN, 
      D=>nx4713, CLK=>nx7142, R=>reset);
   ix4714 : mux21_ni port map ( Y=>nx4713, A0=>q_23_11_EXMPLR, A1=>
      q_22_11_EXMPLR, S0=>nx7024);
   gen_regs_22_regi_reg_q_11 : dffr port map ( Q=>q_22_11_EXMPLR, QB=>OPEN, 
      D=>nx4703, CLK=>nx7142, R=>reset);
   ix4704 : mux21_ni port map ( Y=>nx4703, A0=>q_22_11_EXMPLR, A1=>
      q_21_11_EXMPLR, S0=>nx7024);
   gen_regs_21_regi_reg_q_11 : dffr port map ( Q=>q_21_11_EXMPLR, QB=>OPEN, 
      D=>nx4693, CLK=>nx7142, R=>reset);
   ix4694 : mux21_ni port map ( Y=>nx4693, A0=>q_21_11_EXMPLR, A1=>
      q_20_11_EXMPLR, S0=>nx7024);
   gen_regs_20_regi_reg_q_11 : dffr port map ( Q=>q_20_11_EXMPLR, QB=>OPEN, 
      D=>nx4683, CLK=>nx7142, R=>reset);
   ix4684 : mux21_ni port map ( Y=>nx4683, A0=>q_20_11_EXMPLR, A1=>
      q_19_11_EXMPLR, S0=>nx7024);
   gen_regs_19_regi_reg_q_11 : dffr port map ( Q=>q_19_11_EXMPLR, QB=>OPEN, 
      D=>nx4673, CLK=>nx7142, R=>reset);
   ix4674 : mux21_ni port map ( Y=>nx4673, A0=>q_19_11_EXMPLR, A1=>
      q_18_11_EXMPLR, S0=>nx7024);
   gen_regs_18_regi_reg_q_11 : dffr port map ( Q=>q_18_11_EXMPLR, QB=>OPEN, 
      D=>nx4663, CLK=>nx7140, R=>reset);
   ix4664 : mux21_ni port map ( Y=>nx4663, A0=>q_18_11_EXMPLR, A1=>
      q_17_11_EXMPLR, S0=>nx7022);
   gen_regs_17_regi_reg_q_11 : dffr port map ( Q=>q_17_11_EXMPLR, QB=>OPEN, 
      D=>nx4653, CLK=>nx7140, R=>reset);
   ix4654 : mux21_ni port map ( Y=>nx4653, A0=>q_17_11_EXMPLR, A1=>
      q_16_11_EXMPLR, S0=>nx7022);
   gen_regs_16_regi_reg_q_11 : dffr port map ( Q=>q_16_11_EXMPLR, QB=>OPEN, 
      D=>nx4643, CLK=>nx7140, R=>reset);
   ix4644 : mux21_ni port map ( Y=>nx4643, A0=>q_16_11_EXMPLR, A1=>
      q_15_11_EXMPLR, S0=>nx7022);
   gen_regs_15_regi_reg_q_11 : dffr port map ( Q=>q_15_11_EXMPLR, QB=>OPEN, 
      D=>nx4633, CLK=>nx7140, R=>reset);
   ix4634 : mux21_ni port map ( Y=>nx4633, A0=>q_15_11_EXMPLR, A1=>
      q_14_11_EXMPLR, S0=>nx7022);
   gen_regs_14_regi_reg_q_11 : dffr port map ( Q=>q_14_11_EXMPLR, QB=>OPEN, 
      D=>nx4623, CLK=>nx7140, R=>reset);
   ix4624 : mux21_ni port map ( Y=>nx4623, A0=>q_14_11_EXMPLR, A1=>
      q_13_11_EXMPLR, S0=>nx7022);
   gen_regs_13_regi_reg_q_11 : dffr port map ( Q=>q_13_11_EXMPLR, QB=>OPEN, 
      D=>nx4613, CLK=>nx7140, R=>reset);
   ix4614 : mux21_ni port map ( Y=>nx4613, A0=>q_13_11_EXMPLR, A1=>
      q_12_11_EXMPLR, S0=>nx7022);
   gen_regs_12_regi_reg_q_11 : dffr port map ( Q=>q_12_11_EXMPLR, QB=>OPEN, 
      D=>nx4603, CLK=>nx7140, R=>reset);
   ix4604 : mux21_ni port map ( Y=>nx4603, A0=>q_12_11_EXMPLR, A1=>
      q_11_11_EXMPLR, S0=>nx7022);
   gen_regs_11_regi_reg_q_11 : dffr port map ( Q=>q_11_11_EXMPLR, QB=>OPEN, 
      D=>nx4593, CLK=>nx7138, R=>reset);
   ix4594 : mux21_ni port map ( Y=>nx4593, A0=>q_11_11_EXMPLR, A1=>
      q_10_11_EXMPLR, S0=>nx7020);
   gen_regs_10_regi_reg_q_11 : dffr port map ( Q=>q_10_11_EXMPLR, QB=>OPEN, 
      D=>nx4583, CLK=>nx7138, R=>reset);
   ix4584 : mux21_ni port map ( Y=>nx4583, A0=>q_10_11_EXMPLR, A1=>
      q_9_11_EXMPLR, S0=>nx7020);
   gen_regs_9_regi_reg_q_11 : dffr port map ( Q=>q_9_11_EXMPLR, QB=>OPEN, D
      =>nx4573, CLK=>nx7138, R=>reset);
   ix4574 : mux21_ni port map ( Y=>nx4573, A0=>q_9_11_EXMPLR, A1=>
      q_8_11_EXMPLR, S0=>nx7020);
   gen_regs_8_regi_reg_q_11 : dffr port map ( Q=>q_8_11_EXMPLR, QB=>OPEN, D
      =>nx4563, CLK=>nx7138, R=>reset);
   ix4564 : mux21_ni port map ( Y=>nx4563, A0=>q_8_11_EXMPLR, A1=>
      q_7_11_EXMPLR, S0=>nx7020);
   gen_regs_7_regi_reg_q_11 : dffr port map ( Q=>q_7_11_EXMPLR, QB=>OPEN, D
      =>nx4553, CLK=>nx7138, R=>reset);
   ix4554 : mux21_ni port map ( Y=>nx4553, A0=>q_7_11_EXMPLR, A1=>
      q_6_11_EXMPLR, S0=>nx7020);
   gen_regs_6_regi_reg_q_11 : dffr port map ( Q=>q_6_11_EXMPLR, QB=>OPEN, D
      =>nx4543, CLK=>nx7138, R=>reset);
   ix4544 : mux21_ni port map ( Y=>nx4543, A0=>q_6_11_EXMPLR, A1=>
      q_5_11_EXMPLR, S0=>nx7020);
   gen_regs_5_regi_reg_q_11 : dffr port map ( Q=>q_5_11_EXMPLR, QB=>OPEN, D
      =>nx4533, CLK=>nx7138, R=>reset);
   ix4534 : mux21_ni port map ( Y=>nx4533, A0=>q_5_11_EXMPLR, A1=>
      q_4_11_EXMPLR, S0=>nx7020);
   gen_regs_4_regi_reg_q_11 : dffr port map ( Q=>q_4_11_EXMPLR, QB=>OPEN, D
      =>nx4523, CLK=>nx7136, R=>reset);
   ix4524 : mux21_ni port map ( Y=>nx4523, A0=>q_4_11_EXMPLR, A1=>
      q_3_11_EXMPLR, S0=>nx7018);
   gen_regs_3_regi_reg_q_11 : dffr port map ( Q=>q_3_11_EXMPLR, QB=>OPEN, D
      =>nx4513, CLK=>nx7136, R=>reset);
   ix4514 : mux21_ni port map ( Y=>nx4513, A0=>q_3_11_EXMPLR, A1=>
      q_2_11_EXMPLR, S0=>nx7018);
   gen_regs_2_regi_reg_q_11 : dffr port map ( Q=>q_2_11_EXMPLR, QB=>OPEN, D
      =>nx4503, CLK=>nx7136, R=>reset);
   ix4504 : mux21_ni port map ( Y=>nx4503, A0=>q_2_11_EXMPLR, A1=>
      q_1_11_EXMPLR, S0=>nx7018);
   gen_regs_1_regi_reg_q_11 : dffr port map ( Q=>q_1_11_EXMPLR, QB=>OPEN, D
      =>nx4493, CLK=>nx7136, R=>reset);
   ix4494 : mux21_ni port map ( Y=>nx4493, A0=>q_1_11_EXMPLR, A1=>
      q_0_11_EXMPLR, S0=>nx7018);
   reg0_reg_q_11 : dffr port map ( Q=>q_0_11_EXMPLR, QB=>OPEN, D=>nx4483, 
      CLK=>nx7136, R=>reset);
   ix4484 : mux21_ni port map ( Y=>nx4483, A0=>q_0_11_EXMPLR, A1=>d(11), S0
      =>nx7018);
   gen_regs_24_regi_reg_q_12 : dffr port map ( Q=>q_24_12_EXMPLR, QB=>OPEN, 
      D=>nx4973, CLK=>nx7150, R=>reset);
   ix4974 : mux21_ni port map ( Y=>nx4973, A0=>q_24_12_EXMPLR, A1=>
      q_23_12_EXMPLR, S0=>nx7032);
   gen_regs_23_regi_reg_q_12 : dffr port map ( Q=>q_23_12_EXMPLR, QB=>OPEN, 
      D=>nx4963, CLK=>nx7150, R=>reset);
   ix4964 : mux21_ni port map ( Y=>nx4963, A0=>q_23_12_EXMPLR, A1=>
      q_22_12_EXMPLR, S0=>nx7032);
   gen_regs_22_regi_reg_q_12 : dffr port map ( Q=>q_22_12_EXMPLR, QB=>OPEN, 
      D=>nx4953, CLK=>nx7150, R=>reset);
   ix4954 : mux21_ni port map ( Y=>nx4953, A0=>q_22_12_EXMPLR, A1=>
      q_21_12_EXMPLR, S0=>nx7032);
   gen_regs_21_regi_reg_q_12 : dffr port map ( Q=>q_21_12_EXMPLR, QB=>OPEN, 
      D=>nx4943, CLK=>nx7148, R=>reset);
   ix4944 : mux21_ni port map ( Y=>nx4943, A0=>q_21_12_EXMPLR, A1=>
      q_20_12_EXMPLR, S0=>nx7030);
   gen_regs_20_regi_reg_q_12 : dffr port map ( Q=>q_20_12_EXMPLR, QB=>OPEN, 
      D=>nx4933, CLK=>nx7148, R=>reset);
   ix4934 : mux21_ni port map ( Y=>nx4933, A0=>q_20_12_EXMPLR, A1=>
      q_19_12_EXMPLR, S0=>nx7030);
   gen_regs_19_regi_reg_q_12 : dffr port map ( Q=>q_19_12_EXMPLR, QB=>OPEN, 
      D=>nx4923, CLK=>nx7148, R=>reset);
   ix4924 : mux21_ni port map ( Y=>nx4923, A0=>q_19_12_EXMPLR, A1=>
      q_18_12_EXMPLR, S0=>nx7030);
   gen_regs_18_regi_reg_q_12 : dffr port map ( Q=>q_18_12_EXMPLR, QB=>OPEN, 
      D=>nx4913, CLK=>nx7148, R=>reset);
   ix4914 : mux21_ni port map ( Y=>nx4913, A0=>q_18_12_EXMPLR, A1=>
      q_17_12_EXMPLR, S0=>nx7030);
   gen_regs_17_regi_reg_q_12 : dffr port map ( Q=>q_17_12_EXMPLR, QB=>OPEN, 
      D=>nx4903, CLK=>nx7148, R=>reset);
   ix4904 : mux21_ni port map ( Y=>nx4903, A0=>q_17_12_EXMPLR, A1=>
      q_16_12_EXMPLR, S0=>nx7030);
   gen_regs_16_regi_reg_q_12 : dffr port map ( Q=>q_16_12_EXMPLR, QB=>OPEN, 
      D=>nx4893, CLK=>nx7148, R=>reset);
   ix4894 : mux21_ni port map ( Y=>nx4893, A0=>q_16_12_EXMPLR, A1=>
      q_15_12_EXMPLR, S0=>nx7030);
   gen_regs_15_regi_reg_q_12 : dffr port map ( Q=>q_15_12_EXMPLR, QB=>OPEN, 
      D=>nx4883, CLK=>nx7148, R=>reset);
   ix4884 : mux21_ni port map ( Y=>nx4883, A0=>q_15_12_EXMPLR, A1=>
      q_14_12_EXMPLR, S0=>nx7030);
   gen_regs_14_regi_reg_q_12 : dffr port map ( Q=>q_14_12_EXMPLR, QB=>OPEN, 
      D=>nx4873, CLK=>nx7146, R=>reset);
   ix4874 : mux21_ni port map ( Y=>nx4873, A0=>q_14_12_EXMPLR, A1=>
      q_13_12_EXMPLR, S0=>nx7028);
   gen_regs_13_regi_reg_q_12 : dffr port map ( Q=>q_13_12_EXMPLR, QB=>OPEN, 
      D=>nx4863, CLK=>nx7146, R=>reset);
   ix4864 : mux21_ni port map ( Y=>nx4863, A0=>q_13_12_EXMPLR, A1=>
      q_12_12_EXMPLR, S0=>nx7028);
   gen_regs_12_regi_reg_q_12 : dffr port map ( Q=>q_12_12_EXMPLR, QB=>OPEN, 
      D=>nx4853, CLK=>nx7146, R=>reset);
   ix4854 : mux21_ni port map ( Y=>nx4853, A0=>q_12_12_EXMPLR, A1=>
      q_11_12_EXMPLR, S0=>nx7028);
   gen_regs_11_regi_reg_q_12 : dffr port map ( Q=>q_11_12_EXMPLR, QB=>OPEN, 
      D=>nx4843, CLK=>nx7146, R=>reset);
   ix4844 : mux21_ni port map ( Y=>nx4843, A0=>q_11_12_EXMPLR, A1=>
      q_10_12_EXMPLR, S0=>nx7028);
   gen_regs_10_regi_reg_q_12 : dffr port map ( Q=>q_10_12_EXMPLR, QB=>OPEN, 
      D=>nx4833, CLK=>nx7146, R=>reset);
   ix4834 : mux21_ni port map ( Y=>nx4833, A0=>q_10_12_EXMPLR, A1=>
      q_9_12_EXMPLR, S0=>nx7028);
   gen_regs_9_regi_reg_q_12 : dffr port map ( Q=>q_9_12_EXMPLR, QB=>OPEN, D
      =>nx4823, CLK=>nx7146, R=>reset);
   ix4824 : mux21_ni port map ( Y=>nx4823, A0=>q_9_12_EXMPLR, A1=>
      q_8_12_EXMPLR, S0=>nx7028);
   gen_regs_8_regi_reg_q_12 : dffr port map ( Q=>q_8_12_EXMPLR, QB=>OPEN, D
      =>nx4813, CLK=>nx7146, R=>reset);
   ix4814 : mux21_ni port map ( Y=>nx4813, A0=>q_8_12_EXMPLR, A1=>
      q_7_12_EXMPLR, S0=>nx7028);
   gen_regs_7_regi_reg_q_12 : dffr port map ( Q=>q_7_12_EXMPLR, QB=>OPEN, D
      =>nx4803, CLK=>nx7144, R=>reset);
   ix4804 : mux21_ni port map ( Y=>nx4803, A0=>q_7_12_EXMPLR, A1=>
      q_6_12_EXMPLR, S0=>nx7026);
   gen_regs_6_regi_reg_q_12 : dffr port map ( Q=>q_6_12_EXMPLR, QB=>OPEN, D
      =>nx4793, CLK=>nx7144, R=>reset);
   ix4794 : mux21_ni port map ( Y=>nx4793, A0=>q_6_12_EXMPLR, A1=>
      q_5_12_EXMPLR, S0=>nx7026);
   gen_regs_5_regi_reg_q_12 : dffr port map ( Q=>q_5_12_EXMPLR, QB=>OPEN, D
      =>nx4783, CLK=>nx7144, R=>reset);
   ix4784 : mux21_ni port map ( Y=>nx4783, A0=>q_5_12_EXMPLR, A1=>
      q_4_12_EXMPLR, S0=>nx7026);
   gen_regs_4_regi_reg_q_12 : dffr port map ( Q=>q_4_12_EXMPLR, QB=>OPEN, D
      =>nx4773, CLK=>nx7144, R=>reset);
   ix4774 : mux21_ni port map ( Y=>nx4773, A0=>q_4_12_EXMPLR, A1=>
      q_3_12_EXMPLR, S0=>nx7026);
   gen_regs_3_regi_reg_q_12 : dffr port map ( Q=>q_3_12_EXMPLR, QB=>OPEN, D
      =>nx4763, CLK=>nx7144, R=>reset);
   ix4764 : mux21_ni port map ( Y=>nx4763, A0=>q_3_12_EXMPLR, A1=>
      q_2_12_EXMPLR, S0=>nx7026);
   gen_regs_2_regi_reg_q_12 : dffr port map ( Q=>q_2_12_EXMPLR, QB=>OPEN, D
      =>nx4753, CLK=>nx7144, R=>reset);
   ix4754 : mux21_ni port map ( Y=>nx4753, A0=>q_2_12_EXMPLR, A1=>
      q_1_12_EXMPLR, S0=>nx7026);
   gen_regs_1_regi_reg_q_12 : dffr port map ( Q=>q_1_12_EXMPLR, QB=>OPEN, D
      =>nx4743, CLK=>nx7144, R=>reset);
   ix4744 : mux21_ni port map ( Y=>nx4743, A0=>q_1_12_EXMPLR, A1=>
      q_0_12_EXMPLR, S0=>nx7026);
   reg0_reg_q_12 : dffr port map ( Q=>q_0_12_EXMPLR, QB=>OPEN, D=>nx4733, 
      CLK=>nx7142, R=>reset);
   ix4734 : mux21_ni port map ( Y=>nx4733, A0=>q_0_12_EXMPLR, A1=>d(12), S0
      =>nx7024);
   gen_regs_24_regi_reg_q_13 : dffr port map ( Q=>q_24_13_EXMPLR, QB=>OPEN, 
      D=>nx5223, CLK=>nx7156, R=>reset);
   ix5224 : mux21_ni port map ( Y=>nx5223, A0=>q_24_13_EXMPLR, A1=>
      q_23_13_EXMPLR, S0=>nx7038);
   gen_regs_23_regi_reg_q_13 : dffr port map ( Q=>q_23_13_EXMPLR, QB=>OPEN, 
      D=>nx5213, CLK=>nx7156, R=>reset);
   ix5214 : mux21_ni port map ( Y=>nx5213, A0=>q_23_13_EXMPLR, A1=>
      q_22_13_EXMPLR, S0=>nx7038);
   gen_regs_22_regi_reg_q_13 : dffr port map ( Q=>q_22_13_EXMPLR, QB=>OPEN, 
      D=>nx5203, CLK=>nx7156, R=>reset);
   ix5204 : mux21_ni port map ( Y=>nx5203, A0=>q_22_13_EXMPLR, A1=>
      q_21_13_EXMPLR, S0=>nx7038);
   gen_regs_21_regi_reg_q_13 : dffr port map ( Q=>q_21_13_EXMPLR, QB=>OPEN, 
      D=>nx5193, CLK=>nx7156, R=>reset);
   ix5194 : mux21_ni port map ( Y=>nx5193, A0=>q_21_13_EXMPLR, A1=>
      q_20_13_EXMPLR, S0=>nx7038);
   gen_regs_20_regi_reg_q_13 : dffr port map ( Q=>q_20_13_EXMPLR, QB=>OPEN, 
      D=>nx5183, CLK=>nx7156, R=>reset);
   ix5184 : mux21_ni port map ( Y=>nx5183, A0=>q_20_13_EXMPLR, A1=>
      q_19_13_EXMPLR, S0=>nx7038);
   gen_regs_19_regi_reg_q_13 : dffr port map ( Q=>q_19_13_EXMPLR, QB=>OPEN, 
      D=>nx5173, CLK=>nx7156, R=>reset);
   ix5174 : mux21_ni port map ( Y=>nx5173, A0=>q_19_13_EXMPLR, A1=>
      q_18_13_EXMPLR, S0=>nx7038);
   gen_regs_18_regi_reg_q_13 : dffr port map ( Q=>q_18_13_EXMPLR, QB=>OPEN, 
      D=>nx5163, CLK=>nx7156, R=>reset);
   ix5164 : mux21_ni port map ( Y=>nx5163, A0=>q_18_13_EXMPLR, A1=>
      q_17_13_EXMPLR, S0=>nx7038);
   gen_regs_17_regi_reg_q_13 : dffr port map ( Q=>q_17_13_EXMPLR, QB=>OPEN, 
      D=>nx5153, CLK=>nx7154, R=>reset);
   ix5154 : mux21_ni port map ( Y=>nx5153, A0=>q_17_13_EXMPLR, A1=>
      q_16_13_EXMPLR, S0=>nx7036);
   gen_regs_16_regi_reg_q_13 : dffr port map ( Q=>q_16_13_EXMPLR, QB=>OPEN, 
      D=>nx5143, CLK=>nx7154, R=>reset);
   ix5144 : mux21_ni port map ( Y=>nx5143, A0=>q_16_13_EXMPLR, A1=>
      q_15_13_EXMPLR, S0=>nx7036);
   gen_regs_15_regi_reg_q_13 : dffr port map ( Q=>q_15_13_EXMPLR, QB=>OPEN, 
      D=>nx5133, CLK=>nx7154, R=>reset);
   ix5134 : mux21_ni port map ( Y=>nx5133, A0=>q_15_13_EXMPLR, A1=>
      q_14_13_EXMPLR, S0=>nx7036);
   gen_regs_14_regi_reg_q_13 : dffr port map ( Q=>q_14_13_EXMPLR, QB=>OPEN, 
      D=>nx5123, CLK=>nx7154, R=>reset);
   ix5124 : mux21_ni port map ( Y=>nx5123, A0=>q_14_13_EXMPLR, A1=>
      q_13_13_EXMPLR, S0=>nx7036);
   gen_regs_13_regi_reg_q_13 : dffr port map ( Q=>q_13_13_EXMPLR, QB=>OPEN, 
      D=>nx5113, CLK=>nx7154, R=>reset);
   ix5114 : mux21_ni port map ( Y=>nx5113, A0=>q_13_13_EXMPLR, A1=>
      q_12_13_EXMPLR, S0=>nx7036);
   gen_regs_12_regi_reg_q_13 : dffr port map ( Q=>q_12_13_EXMPLR, QB=>OPEN, 
      D=>nx5103, CLK=>nx7154, R=>reset);
   ix5104 : mux21_ni port map ( Y=>nx5103, A0=>q_12_13_EXMPLR, A1=>
      q_11_13_EXMPLR, S0=>nx7036);
   gen_regs_11_regi_reg_q_13 : dffr port map ( Q=>q_11_13_EXMPLR, QB=>OPEN, 
      D=>nx5093, CLK=>nx7154, R=>reset);
   ix5094 : mux21_ni port map ( Y=>nx5093, A0=>q_11_13_EXMPLR, A1=>
      q_10_13_EXMPLR, S0=>nx7036);
   gen_regs_10_regi_reg_q_13 : dffr port map ( Q=>q_10_13_EXMPLR, QB=>OPEN, 
      D=>nx5083, CLK=>nx7152, R=>reset);
   ix5084 : mux21_ni port map ( Y=>nx5083, A0=>q_10_13_EXMPLR, A1=>
      q_9_13_EXMPLR, S0=>nx7034);
   gen_regs_9_regi_reg_q_13 : dffr port map ( Q=>q_9_13_EXMPLR, QB=>OPEN, D
      =>nx5073, CLK=>nx7152, R=>reset);
   ix5074 : mux21_ni port map ( Y=>nx5073, A0=>q_9_13_EXMPLR, A1=>
      q_8_13_EXMPLR, S0=>nx7034);
   gen_regs_8_regi_reg_q_13 : dffr port map ( Q=>q_8_13_EXMPLR, QB=>OPEN, D
      =>nx5063, CLK=>nx7152, R=>reset);
   ix5064 : mux21_ni port map ( Y=>nx5063, A0=>q_8_13_EXMPLR, A1=>
      q_7_13_EXMPLR, S0=>nx7034);
   gen_regs_7_regi_reg_q_13 : dffr port map ( Q=>q_7_13_EXMPLR, QB=>OPEN, D
      =>nx5053, CLK=>nx7152, R=>reset);
   ix5054 : mux21_ni port map ( Y=>nx5053, A0=>q_7_13_EXMPLR, A1=>
      q_6_13_EXMPLR, S0=>nx7034);
   gen_regs_6_regi_reg_q_13 : dffr port map ( Q=>q_6_13_EXMPLR, QB=>OPEN, D
      =>nx5043, CLK=>nx7152, R=>reset);
   ix5044 : mux21_ni port map ( Y=>nx5043, A0=>q_6_13_EXMPLR, A1=>
      q_5_13_EXMPLR, S0=>nx7034);
   gen_regs_5_regi_reg_q_13 : dffr port map ( Q=>q_5_13_EXMPLR, QB=>OPEN, D
      =>nx5033, CLK=>nx7152, R=>reset);
   ix5034 : mux21_ni port map ( Y=>nx5033, A0=>q_5_13_EXMPLR, A1=>
      q_4_13_EXMPLR, S0=>nx7034);
   gen_regs_4_regi_reg_q_13 : dffr port map ( Q=>q_4_13_EXMPLR, QB=>OPEN, D
      =>nx5023, CLK=>nx7152, R=>reset);
   ix5024 : mux21_ni port map ( Y=>nx5023, A0=>q_4_13_EXMPLR, A1=>
      q_3_13_EXMPLR, S0=>nx7034);
   gen_regs_3_regi_reg_q_13 : dffr port map ( Q=>q_3_13_EXMPLR, QB=>OPEN, D
      =>nx5013, CLK=>nx7150, R=>reset);
   ix5014 : mux21_ni port map ( Y=>nx5013, A0=>q_3_13_EXMPLR, A1=>
      q_2_13_EXMPLR, S0=>nx7032);
   gen_regs_2_regi_reg_q_13 : dffr port map ( Q=>q_2_13_EXMPLR, QB=>OPEN, D
      =>nx5003, CLK=>nx7150, R=>reset);
   ix5004 : mux21_ni port map ( Y=>nx5003, A0=>q_2_13_EXMPLR, A1=>
      q_1_13_EXMPLR, S0=>nx7032);
   gen_regs_1_regi_reg_q_13 : dffr port map ( Q=>q_1_13_EXMPLR, QB=>OPEN, D
      =>nx4993, CLK=>nx7150, R=>reset);
   ix4994 : mux21_ni port map ( Y=>nx4993, A0=>q_1_13_EXMPLR, A1=>
      q_0_13_EXMPLR, S0=>nx7032);
   reg0_reg_q_13 : dffr port map ( Q=>q_0_13_EXMPLR, QB=>OPEN, D=>nx4983, 
      CLK=>nx7150, R=>reset);
   ix4984 : mux21_ni port map ( Y=>nx4983, A0=>q_0_13_EXMPLR, A1=>d(13), S0
      =>nx7032);
   gen_regs_24_regi_reg_q_14 : dffr port map ( Q=>q_24_14_EXMPLR, QB=>OPEN, 
      D=>nx5473, CLK=>nx7164, R=>reset);
   ix5474 : mux21_ni port map ( Y=>nx5473, A0=>q_24_14_EXMPLR, A1=>
      q_23_14_EXMPLR, S0=>nx7046);
   gen_regs_23_regi_reg_q_14 : dffr port map ( Q=>q_23_14_EXMPLR, QB=>OPEN, 
      D=>nx5463, CLK=>nx7164, R=>reset);
   ix5464 : mux21_ni port map ( Y=>nx5463, A0=>q_23_14_EXMPLR, A1=>
      q_22_14_EXMPLR, S0=>nx7046);
   gen_regs_22_regi_reg_q_14 : dffr port map ( Q=>q_22_14_EXMPLR, QB=>OPEN, 
      D=>nx5453, CLK=>nx7164, R=>reset);
   ix5454 : mux21_ni port map ( Y=>nx5453, A0=>q_22_14_EXMPLR, A1=>
      q_21_14_EXMPLR, S0=>nx7046);
   gen_regs_21_regi_reg_q_14 : dffr port map ( Q=>q_21_14_EXMPLR, QB=>OPEN, 
      D=>nx5443, CLK=>nx7164, R=>reset);
   ix5444 : mux21_ni port map ( Y=>nx5443, A0=>q_21_14_EXMPLR, A1=>
      q_20_14_EXMPLR, S0=>nx7046);
   gen_regs_20_regi_reg_q_14 : dffr port map ( Q=>q_20_14_EXMPLR, QB=>OPEN, 
      D=>nx5433, CLK=>nx7162, R=>reset);
   ix5434 : mux21_ni port map ( Y=>nx5433, A0=>q_20_14_EXMPLR, A1=>
      q_19_14_EXMPLR, S0=>nx7044);
   gen_regs_19_regi_reg_q_14 : dffr port map ( Q=>q_19_14_EXMPLR, QB=>OPEN, 
      D=>nx5423, CLK=>nx7162, R=>reset);
   ix5424 : mux21_ni port map ( Y=>nx5423, A0=>q_19_14_EXMPLR, A1=>
      q_18_14_EXMPLR, S0=>nx7044);
   gen_regs_18_regi_reg_q_14 : dffr port map ( Q=>q_18_14_EXMPLR, QB=>OPEN, 
      D=>nx5413, CLK=>nx7162, R=>reset);
   ix5414 : mux21_ni port map ( Y=>nx5413, A0=>q_18_14_EXMPLR, A1=>
      q_17_14_EXMPLR, S0=>nx7044);
   gen_regs_17_regi_reg_q_14 : dffr port map ( Q=>q_17_14_EXMPLR, QB=>OPEN, 
      D=>nx5403, CLK=>nx7162, R=>reset);
   ix5404 : mux21_ni port map ( Y=>nx5403, A0=>q_17_14_EXMPLR, A1=>
      q_16_14_EXMPLR, S0=>nx7044);
   gen_regs_16_regi_reg_q_14 : dffr port map ( Q=>q_16_14_EXMPLR, QB=>OPEN, 
      D=>nx5393, CLK=>nx7162, R=>reset);
   ix5394 : mux21_ni port map ( Y=>nx5393, A0=>q_16_14_EXMPLR, A1=>
      q_15_14_EXMPLR, S0=>nx7044);
   gen_regs_15_regi_reg_q_14 : dffr port map ( Q=>q_15_14_EXMPLR, QB=>OPEN, 
      D=>nx5383, CLK=>nx7162, R=>reset);
   ix5384 : mux21_ni port map ( Y=>nx5383, A0=>q_15_14_EXMPLR, A1=>
      q_14_14_EXMPLR, S0=>nx7044);
   gen_regs_14_regi_reg_q_14 : dffr port map ( Q=>q_14_14_EXMPLR, QB=>OPEN, 
      D=>nx5373, CLK=>nx7162, R=>reset);
   ix5374 : mux21_ni port map ( Y=>nx5373, A0=>q_14_14_EXMPLR, A1=>
      q_13_14_EXMPLR, S0=>nx7044);
   gen_regs_13_regi_reg_q_14 : dffr port map ( Q=>q_13_14_EXMPLR, QB=>OPEN, 
      D=>nx5363, CLK=>nx7160, R=>reset);
   ix5364 : mux21_ni port map ( Y=>nx5363, A0=>q_13_14_EXMPLR, A1=>
      q_12_14_EXMPLR, S0=>nx7042);
   gen_regs_12_regi_reg_q_14 : dffr port map ( Q=>q_12_14_EXMPLR, QB=>OPEN, 
      D=>nx5353, CLK=>nx7160, R=>reset);
   ix5354 : mux21_ni port map ( Y=>nx5353, A0=>q_12_14_EXMPLR, A1=>
      q_11_14_EXMPLR, S0=>nx7042);
   gen_regs_11_regi_reg_q_14 : dffr port map ( Q=>q_11_14_EXMPLR, QB=>OPEN, 
      D=>nx5343, CLK=>nx7160, R=>reset);
   ix5344 : mux21_ni port map ( Y=>nx5343, A0=>q_11_14_EXMPLR, A1=>
      q_10_14_EXMPLR, S0=>nx7042);
   gen_regs_10_regi_reg_q_14 : dffr port map ( Q=>q_10_14_EXMPLR, QB=>OPEN, 
      D=>nx5333, CLK=>nx7160, R=>reset);
   ix5334 : mux21_ni port map ( Y=>nx5333, A0=>q_10_14_EXMPLR, A1=>
      q_9_14_EXMPLR, S0=>nx7042);
   gen_regs_9_regi_reg_q_14 : dffr port map ( Q=>q_9_14_EXMPLR, QB=>OPEN, D
      =>nx5323, CLK=>nx7160, R=>reset);
   ix5324 : mux21_ni port map ( Y=>nx5323, A0=>q_9_14_EXMPLR, A1=>
      q_8_14_EXMPLR, S0=>nx7042);
   gen_regs_8_regi_reg_q_14 : dffr port map ( Q=>q_8_14_EXMPLR, QB=>OPEN, D
      =>nx5313, CLK=>nx7160, R=>reset);
   ix5314 : mux21_ni port map ( Y=>nx5313, A0=>q_8_14_EXMPLR, A1=>
      q_7_14_EXMPLR, S0=>nx7042);
   gen_regs_7_regi_reg_q_14 : dffr port map ( Q=>q_7_14_EXMPLR, QB=>OPEN, D
      =>nx5303, CLK=>nx7160, R=>reset);
   ix5304 : mux21_ni port map ( Y=>nx5303, A0=>q_7_14_EXMPLR, A1=>
      q_6_14_EXMPLR, S0=>nx7042);
   gen_regs_6_regi_reg_q_14 : dffr port map ( Q=>q_6_14_EXMPLR, QB=>OPEN, D
      =>nx5293, CLK=>nx7158, R=>reset);
   ix5294 : mux21_ni port map ( Y=>nx5293, A0=>q_6_14_EXMPLR, A1=>
      q_5_14_EXMPLR, S0=>nx7040);
   gen_regs_5_regi_reg_q_14 : dffr port map ( Q=>q_5_14_EXMPLR, QB=>OPEN, D
      =>nx5283, CLK=>nx7158, R=>reset);
   ix5284 : mux21_ni port map ( Y=>nx5283, A0=>q_5_14_EXMPLR, A1=>
      q_4_14_EXMPLR, S0=>nx7040);
   gen_regs_4_regi_reg_q_14 : dffr port map ( Q=>q_4_14_EXMPLR, QB=>OPEN, D
      =>nx5273, CLK=>nx7158, R=>reset);
   ix5274 : mux21_ni port map ( Y=>nx5273, A0=>q_4_14_EXMPLR, A1=>
      q_3_14_EXMPLR, S0=>nx7040);
   gen_regs_3_regi_reg_q_14 : dffr port map ( Q=>q_3_14_EXMPLR, QB=>OPEN, D
      =>nx5263, CLK=>nx7158, R=>reset);
   ix5264 : mux21_ni port map ( Y=>nx5263, A0=>q_3_14_EXMPLR, A1=>
      q_2_14_EXMPLR, S0=>nx7040);
   gen_regs_2_regi_reg_q_14 : dffr port map ( Q=>q_2_14_EXMPLR, QB=>OPEN, D
      =>nx5253, CLK=>nx7158, R=>reset);
   ix5254 : mux21_ni port map ( Y=>nx5253, A0=>q_2_14_EXMPLR, A1=>
      q_1_14_EXMPLR, S0=>nx7040);
   gen_regs_1_regi_reg_q_14 : dffr port map ( Q=>q_1_14_EXMPLR, QB=>OPEN, D
      =>nx5243, CLK=>nx7158, R=>reset);
   ix5244 : mux21_ni port map ( Y=>nx5243, A0=>q_1_14_EXMPLR, A1=>
      q_0_14_EXMPLR, S0=>nx7040);
   reg0_reg_q_14 : dffr port map ( Q=>q_0_14_EXMPLR, QB=>OPEN, D=>nx5233, 
      CLK=>nx7158, R=>reset);
   ix5234 : mux21_ni port map ( Y=>nx5233, A0=>q_0_14_EXMPLR, A1=>d(14), S0
      =>nx7040);
   gen_regs_24_regi_reg_q_15 : dffr port map ( Q=>q_24_15_EXMPLR, QB=>OPEN, 
      D=>nx5723, CLK=>nx7172, R=>reset);
   ix5724 : mux21_ni port map ( Y=>nx5723, A0=>q_24_15_EXMPLR, A1=>
      q_23_15_EXMPLR, S0=>nx7054);
   gen_regs_23_regi_reg_q_15 : dffr port map ( Q=>q_23_15_EXMPLR, QB=>OPEN, 
      D=>nx5713, CLK=>nx7170, R=>reset);
   ix5714 : mux21_ni port map ( Y=>nx5713, A0=>q_23_15_EXMPLR, A1=>
      q_22_15_EXMPLR, S0=>nx7052);
   gen_regs_22_regi_reg_q_15 : dffr port map ( Q=>q_22_15_EXMPLR, QB=>OPEN, 
      D=>nx5703, CLK=>nx7170, R=>reset);
   ix5704 : mux21_ni port map ( Y=>nx5703, A0=>q_22_15_EXMPLR, A1=>
      q_21_15_EXMPLR, S0=>nx7052);
   gen_regs_21_regi_reg_q_15 : dffr port map ( Q=>q_21_15_EXMPLR, QB=>OPEN, 
      D=>nx5693, CLK=>nx7170, R=>reset);
   ix5694 : mux21_ni port map ( Y=>nx5693, A0=>q_21_15_EXMPLR, A1=>
      q_20_15_EXMPLR, S0=>nx7052);
   gen_regs_20_regi_reg_q_15 : dffr port map ( Q=>q_20_15_EXMPLR, QB=>OPEN, 
      D=>nx5683, CLK=>nx7170, R=>reset);
   ix5684 : mux21_ni port map ( Y=>nx5683, A0=>q_20_15_EXMPLR, A1=>
      q_19_15_EXMPLR, S0=>nx7052);
   gen_regs_19_regi_reg_q_15 : dffr port map ( Q=>q_19_15_EXMPLR, QB=>OPEN, 
      D=>nx5673, CLK=>nx7170, R=>reset);
   ix5674 : mux21_ni port map ( Y=>nx5673, A0=>q_19_15_EXMPLR, A1=>
      q_18_15_EXMPLR, S0=>nx7052);
   gen_regs_18_regi_reg_q_15 : dffr port map ( Q=>q_18_15_EXMPLR, QB=>OPEN, 
      D=>nx5663, CLK=>nx7170, R=>reset);
   ix5664 : mux21_ni port map ( Y=>nx5663, A0=>q_18_15_EXMPLR, A1=>
      q_17_15_EXMPLR, S0=>nx7052);
   gen_regs_17_regi_reg_q_15 : dffr port map ( Q=>q_17_15_EXMPLR, QB=>OPEN, 
      D=>nx5653, CLK=>nx7170, R=>reset);
   ix5654 : mux21_ni port map ( Y=>nx5653, A0=>q_17_15_EXMPLR, A1=>
      q_16_15_EXMPLR, S0=>nx7052);
   gen_regs_16_regi_reg_q_15 : dffr port map ( Q=>q_16_15_EXMPLR, QB=>OPEN, 
      D=>nx5643, CLK=>nx7168, R=>reset);
   ix5644 : mux21_ni port map ( Y=>nx5643, A0=>q_16_15_EXMPLR, A1=>
      q_15_15_EXMPLR, S0=>nx7050);
   gen_regs_15_regi_reg_q_15 : dffr port map ( Q=>q_15_15_EXMPLR, QB=>OPEN, 
      D=>nx5633, CLK=>nx7168, R=>reset);
   ix5634 : mux21_ni port map ( Y=>nx5633, A0=>q_15_15_EXMPLR, A1=>
      q_14_15_EXMPLR, S0=>nx7050);
   gen_regs_14_regi_reg_q_15 : dffr port map ( Q=>q_14_15_EXMPLR, QB=>OPEN, 
      D=>nx5623, CLK=>nx7168, R=>reset);
   ix5624 : mux21_ni port map ( Y=>nx5623, A0=>q_14_15_EXMPLR, A1=>
      q_13_15_EXMPLR, S0=>nx7050);
   gen_regs_13_regi_reg_q_15 : dffr port map ( Q=>q_13_15_EXMPLR, QB=>OPEN, 
      D=>nx5613, CLK=>nx7168, R=>reset);
   ix5614 : mux21_ni port map ( Y=>nx5613, A0=>q_13_15_EXMPLR, A1=>
      q_12_15_EXMPLR, S0=>nx7050);
   gen_regs_12_regi_reg_q_15 : dffr port map ( Q=>q_12_15_EXMPLR, QB=>OPEN, 
      D=>nx5603, CLK=>nx7168, R=>reset);
   ix5604 : mux21_ni port map ( Y=>nx5603, A0=>q_12_15_EXMPLR, A1=>
      q_11_15_EXMPLR, S0=>nx7050);
   gen_regs_11_regi_reg_q_15 : dffr port map ( Q=>q_11_15_EXMPLR, QB=>OPEN, 
      D=>nx5593, CLK=>nx7168, R=>reset);
   ix5594 : mux21_ni port map ( Y=>nx5593, A0=>q_11_15_EXMPLR, A1=>
      q_10_15_EXMPLR, S0=>nx7050);
   gen_regs_10_regi_reg_q_15 : dffr port map ( Q=>q_10_15_EXMPLR, QB=>OPEN, 
      D=>nx5583, CLK=>nx7168, R=>reset);
   ix5584 : mux21_ni port map ( Y=>nx5583, A0=>q_10_15_EXMPLR, A1=>
      q_9_15_EXMPLR, S0=>nx7050);
   gen_regs_9_regi_reg_q_15 : dffr port map ( Q=>q_9_15_EXMPLR, QB=>OPEN, D
      =>nx5573, CLK=>nx7166, R=>reset);
   ix5574 : mux21_ni port map ( Y=>nx5573, A0=>q_9_15_EXMPLR, A1=>
      q_8_15_EXMPLR, S0=>nx7048);
   gen_regs_8_regi_reg_q_15 : dffr port map ( Q=>q_8_15_EXMPLR, QB=>OPEN, D
      =>nx5563, CLK=>nx7166, R=>reset);
   ix5564 : mux21_ni port map ( Y=>nx5563, A0=>q_8_15_EXMPLR, A1=>
      q_7_15_EXMPLR, S0=>nx7048);
   gen_regs_7_regi_reg_q_15 : dffr port map ( Q=>q_7_15_EXMPLR, QB=>OPEN, D
      =>nx5553, CLK=>nx7166, R=>reset);
   ix5554 : mux21_ni port map ( Y=>nx5553, A0=>q_7_15_EXMPLR, A1=>
      q_6_15_EXMPLR, S0=>nx7048);
   gen_regs_6_regi_reg_q_15 : dffr port map ( Q=>q_6_15_EXMPLR, QB=>OPEN, D
      =>nx5543, CLK=>nx7166, R=>reset);
   ix5544 : mux21_ni port map ( Y=>nx5543, A0=>q_6_15_EXMPLR, A1=>
      q_5_15_EXMPLR, S0=>nx7048);
   gen_regs_5_regi_reg_q_15 : dffr port map ( Q=>q_5_15_EXMPLR, QB=>OPEN, D
      =>nx5533, CLK=>nx7166, R=>reset);
   ix5534 : mux21_ni port map ( Y=>nx5533, A0=>q_5_15_EXMPLR, A1=>
      q_4_15_EXMPLR, S0=>nx7048);
   gen_regs_4_regi_reg_q_15 : dffr port map ( Q=>q_4_15_EXMPLR, QB=>OPEN, D
      =>nx5523, CLK=>nx7166, R=>reset);
   ix5524 : mux21_ni port map ( Y=>nx5523, A0=>q_4_15_EXMPLR, A1=>
      q_3_15_EXMPLR, S0=>nx7048);
   gen_regs_3_regi_reg_q_15 : dffr port map ( Q=>q_3_15_EXMPLR, QB=>OPEN, D
      =>nx5513, CLK=>nx7166, R=>reset);
   ix5514 : mux21_ni port map ( Y=>nx5513, A0=>q_3_15_EXMPLR, A1=>
      q_2_15_EXMPLR, S0=>nx7048);
   gen_regs_2_regi_reg_q_15 : dffr port map ( Q=>q_2_15_EXMPLR, QB=>OPEN, D
      =>nx5503, CLK=>nx7164, R=>reset);
   ix5504 : mux21_ni port map ( Y=>nx5503, A0=>q_2_15_EXMPLR, A1=>
      q_1_15_EXMPLR, S0=>nx7046);
   gen_regs_1_regi_reg_q_15 : dffr port map ( Q=>q_1_15_EXMPLR, QB=>OPEN, D
      =>nx5493, CLK=>nx7164, R=>reset);
   ix5494 : mux21_ni port map ( Y=>nx5493, A0=>q_1_15_EXMPLR, A1=>
      q_0_15_EXMPLR, S0=>nx7046);
   reg0_reg_q_15 : dffr port map ( Q=>q_0_15_EXMPLR, QB=>OPEN, D=>nx5483, 
      CLK=>nx7164, R=>reset);
   ix5484 : mux21_ni port map ( Y=>nx5483, A0=>q_0_15_EXMPLR, A1=>d(15), S0
      =>nx7046);
   ix6939 : inv02 port map ( Y=>nx6940, A=>nx7626);
   ix6941 : inv02 port map ( Y=>nx6942, A=>nx7626);
   ix6943 : inv02 port map ( Y=>nx6944, A=>nx7626);
   ix6945 : inv02 port map ( Y=>nx6946, A=>nx7626);
   ix6947 : inv02 port map ( Y=>nx6948, A=>nx7626);
   ix6949 : inv02 port map ( Y=>nx6950, A=>nx7626);
   ix6951 : inv02 port map ( Y=>nx6952, A=>nx7174);
   ix6953 : inv02 port map ( Y=>nx6954, A=>nx7176);
   ix6955 : inv02 port map ( Y=>nx6956, A=>nx7176);
   ix6957 : inv02 port map ( Y=>nx6958, A=>nx7176);
   ix6959 : inv02 port map ( Y=>nx6960, A=>nx7176);
   ix6961 : inv02 port map ( Y=>nx6962, A=>nx7176);
   ix6963 : inv02 port map ( Y=>nx6964, A=>nx7176);
   ix6965 : inv02 port map ( Y=>nx6966, A=>nx7176);
   ix6967 : inv02 port map ( Y=>nx6968, A=>nx7178);
   ix6969 : inv02 port map ( Y=>nx6970, A=>nx7178);
   ix6971 : inv02 port map ( Y=>nx6972, A=>nx7178);
   ix6973 : inv02 port map ( Y=>nx6974, A=>nx7178);
   ix6975 : inv02 port map ( Y=>nx6976, A=>nx7178);
   ix6977 : inv02 port map ( Y=>nx6978, A=>nx7178);
   ix6979 : inv02 port map ( Y=>nx6980, A=>nx7178);
   ix6981 : inv02 port map ( Y=>nx6982, A=>nx7180);
   ix6983 : inv02 port map ( Y=>nx6984, A=>nx7180);
   ix6985 : inv02 port map ( Y=>nx6986, A=>nx7180);
   ix6987 : inv02 port map ( Y=>nx6988, A=>nx7180);
   ix6989 : inv02 port map ( Y=>nx6990, A=>nx7180);
   ix6991 : inv02 port map ( Y=>nx6992, A=>nx7180);
   ix6993 : inv02 port map ( Y=>nx6994, A=>nx7180);
   ix6995 : inv02 port map ( Y=>nx6996, A=>nx7182);
   ix6997 : inv02 port map ( Y=>nx6998, A=>nx7182);
   ix6999 : inv02 port map ( Y=>nx7000, A=>nx7182);
   ix7001 : inv02 port map ( Y=>nx7002, A=>nx7182);
   ix7003 : inv02 port map ( Y=>nx7004, A=>nx7182);
   ix7005 : inv02 port map ( Y=>nx7006, A=>nx7182);
   ix7007 : inv02 port map ( Y=>nx7008, A=>nx7182);
   ix7009 : inv02 port map ( Y=>nx7010, A=>nx7184);
   ix7011 : inv02 port map ( Y=>nx7012, A=>nx7184);
   ix7013 : inv02 port map ( Y=>nx7014, A=>nx7184);
   ix7015 : inv02 port map ( Y=>nx7016, A=>nx7184);
   ix7017 : inv02 port map ( Y=>nx7018, A=>nx7184);
   ix7019 : inv02 port map ( Y=>nx7020, A=>nx7184);
   ix7021 : inv02 port map ( Y=>nx7022, A=>nx7184);
   ix7023 : inv02 port map ( Y=>nx7024, A=>nx7186);
   ix7025 : inv02 port map ( Y=>nx7026, A=>nx7186);
   ix7027 : inv02 port map ( Y=>nx7028, A=>nx7186);
   ix7029 : inv02 port map ( Y=>nx7030, A=>nx7186);
   ix7031 : inv02 port map ( Y=>nx7032, A=>nx7186);
   ix7033 : inv02 port map ( Y=>nx7034, A=>nx7186);
   ix7035 : inv02 port map ( Y=>nx7036, A=>nx7186);
   ix7037 : inv02 port map ( Y=>nx7038, A=>nx7188);
   ix7039 : inv02 port map ( Y=>nx7040, A=>nx7188);
   ix7041 : inv02 port map ( Y=>nx7042, A=>nx7188);
   ix7043 : inv02 port map ( Y=>nx7044, A=>nx7188);
   ix7045 : inv02 port map ( Y=>nx7046, A=>nx7188);
   ix7047 : inv02 port map ( Y=>nx7048, A=>nx7188);
   ix7049 : inv02 port map ( Y=>nx7050, A=>nx7188);
   ix7051 : inv02 port map ( Y=>nx7052, A=>nx7190);
   ix7053 : inv02 port map ( Y=>nx7054, A=>nx7190);
   ix7057 : inv02 port map ( Y=>nx7058, A=>nx7628);
   ix7059 : inv02 port map ( Y=>nx7060, A=>nx7628);
   ix7061 : inv02 port map ( Y=>nx7062, A=>nx7628);
   ix7063 : inv02 port map ( Y=>nx7064, A=>nx7628);
   ix7065 : inv02 port map ( Y=>nx7066, A=>nx7628);
   ix7067 : inv02 port map ( Y=>nx7068, A=>nx7628);
   ix7069 : inv02 port map ( Y=>nx7070, A=>nx7192);
   ix7071 : inv02 port map ( Y=>nx7072, A=>nx7194);
   ix7073 : inv02 port map ( Y=>nx7074, A=>nx7194);
   ix7075 : inv02 port map ( Y=>nx7076, A=>nx7194);
   ix7077 : inv02 port map ( Y=>nx7078, A=>nx7194);
   ix7079 : inv02 port map ( Y=>nx7080, A=>nx7194);
   ix7081 : inv02 port map ( Y=>nx7082, A=>nx7194);
   ix7083 : inv02 port map ( Y=>nx7084, A=>nx7194);
   ix7085 : inv02 port map ( Y=>nx7086, A=>nx7196);
   ix7087 : inv02 port map ( Y=>nx7088, A=>nx7196);
   ix7089 : inv02 port map ( Y=>nx7090, A=>nx7196);
   ix7091 : inv02 port map ( Y=>nx7092, A=>nx7196);
   ix7093 : inv02 port map ( Y=>nx7094, A=>nx7196);
   ix7095 : inv02 port map ( Y=>nx7096, A=>nx7196);
   ix7097 : inv02 port map ( Y=>nx7098, A=>nx7196);
   ix7099 : inv02 port map ( Y=>nx7100, A=>nx7198);
   ix7101 : inv02 port map ( Y=>nx7102, A=>nx7198);
   ix7103 : inv02 port map ( Y=>nx7104, A=>nx7198);
   ix7105 : inv02 port map ( Y=>nx7106, A=>nx7198);
   ix7107 : inv02 port map ( Y=>nx7108, A=>nx7198);
   ix7109 : inv02 port map ( Y=>nx7110, A=>nx7198);
   ix7111 : inv02 port map ( Y=>nx7112, A=>nx7198);
   ix7113 : inv02 port map ( Y=>nx7114, A=>nx7200);
   ix7115 : inv02 port map ( Y=>nx7116, A=>nx7200);
   ix7117 : inv02 port map ( Y=>nx7118, A=>nx7200);
   ix7119 : inv02 port map ( Y=>nx7120, A=>nx7200);
   ix7121 : inv02 port map ( Y=>nx7122, A=>nx7200);
   ix7123 : inv02 port map ( Y=>nx7124, A=>nx7200);
   ix7125 : inv02 port map ( Y=>nx7126, A=>nx7200);
   ix7127 : inv02 port map ( Y=>nx7128, A=>nx7202);
   ix7129 : inv02 port map ( Y=>nx7130, A=>nx7202);
   ix7131 : inv02 port map ( Y=>nx7132, A=>nx7202);
   ix7133 : inv02 port map ( Y=>nx7134, A=>nx7202);
   ix7135 : inv02 port map ( Y=>nx7136, A=>nx7202);
   ix7137 : inv02 port map ( Y=>nx7138, A=>nx7202);
   ix7139 : inv02 port map ( Y=>nx7140, A=>nx7202);
   ix7141 : inv02 port map ( Y=>nx7142, A=>nx7204);
   ix7143 : inv02 port map ( Y=>nx7144, A=>nx7204);
   ix7145 : inv02 port map ( Y=>nx7146, A=>nx7204);
   ix7147 : inv02 port map ( Y=>nx7148, A=>nx7204);
   ix7149 : inv02 port map ( Y=>nx7150, A=>nx7204);
   ix7151 : inv02 port map ( Y=>nx7152, A=>nx7204);
   ix7153 : inv02 port map ( Y=>nx7154, A=>nx7204);
   ix7155 : inv02 port map ( Y=>nx7156, A=>nx7206);
   ix7157 : inv02 port map ( Y=>nx7158, A=>nx7206);
   ix7159 : inv02 port map ( Y=>nx7160, A=>nx7206);
   ix7161 : inv02 port map ( Y=>nx7162, A=>nx7206);
   ix7163 : inv02 port map ( Y=>nx7164, A=>nx7206);
   ix7165 : inv02 port map ( Y=>nx7166, A=>nx7206);
   ix7167 : inv02 port map ( Y=>nx7168, A=>nx7206);
   ix7169 : inv02 port map ( Y=>nx7170, A=>nx7208);
   ix7171 : inv02 port map ( Y=>nx7172, A=>nx7208);
   ix7173 : inv02 port map ( Y=>nx7174, A=>load);
   ix7175 : inv02 port map ( Y=>nx7176, A=>nx7214);
   ix7177 : inv02 port map ( Y=>nx7178, A=>nx7214);
   ix7179 : inv02 port map ( Y=>nx7180, A=>nx7214);
   ix7181 : inv02 port map ( Y=>nx7182, A=>nx7214);
   ix7183 : inv02 port map ( Y=>nx7184, A=>nx7214);
   ix7185 : inv02 port map ( Y=>nx7186, A=>nx7216);
   ix7187 : inv02 port map ( Y=>nx7188, A=>nx7216);
   ix7189 : inv02 port map ( Y=>nx7190, A=>nx7216);
   ix7191 : inv02 port map ( Y=>nx7192, A=>clk);
   ix7193 : inv02 port map ( Y=>nx7194, A=>nx7218);
   ix7195 : inv02 port map ( Y=>nx7196, A=>nx7218);
   ix7197 : inv02 port map ( Y=>nx7198, A=>nx7218);
   ix7199 : inv02 port map ( Y=>nx7200, A=>nx7218);
   ix7201 : inv02 port map ( Y=>nx7202, A=>nx7218);
   ix7203 : inv02 port map ( Y=>nx7204, A=>nx7220);
   ix7205 : inv02 port map ( Y=>nx7206, A=>nx7220);
   ix7207 : inv02 port map ( Y=>nx7208, A=>nx7220);
   ix7213 : inv01 port map ( Y=>nx7214, A=>nx7626);
   ix7215 : inv01 port map ( Y=>nx7216, A=>nx7174);
   ix7217 : inv01 port map ( Y=>nx7218, A=>nx7628);
   ix7219 : inv01 port map ( Y=>nx7220, A=>nx7192);
   ix7625 : inv02 port map ( Y=>nx7626, A=>load);
   ix7627 : inv02 port map ( Y=>nx7628, A=>clk);
end Structural ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Reg_32 is
   port (
      d : IN std_logic_vector (31 DOWNTO 0) ;
      q : OUT std_logic_vector (31 DOWNTO 0) ;
      rst_data : IN std_logic_vector (31 DOWNTO 0) ;
      clk : IN std_logic ;
      load : IN std_logic ;
      reset : IN std_logic) ;
end Reg_32 ;

architecture Behavioral_unfold_3258 of Reg_32 is
   signal q_31_EXMPLR, q_30_EXMPLR, q_29_EXMPLR, q_28_EXMPLR, q_27_EXMPLR, 
      q_26_EXMPLR, q_25_EXMPLR, q_24_EXMPLR, q_23_EXMPLR, q_22_EXMPLR, 
      q_21_EXMPLR, q_20_EXMPLR, q_19_EXMPLR, q_18_EXMPLR, q_17_EXMPLR, 
      q_16_EXMPLR, q_15_EXMPLR, q_14_EXMPLR, q_13_EXMPLR, q_12_EXMPLR, 
      q_11_EXMPLR, q_10_EXMPLR, q_9_EXMPLR, q_8_EXMPLR, q_7_EXMPLR, 
      q_6_EXMPLR, q_5_EXMPLR, q_4_EXMPLR, q_3_EXMPLR, q_2_EXMPLR, q_1_EXMPLR, 
      q_0_EXMPLR, nx114, nx124, nx134, nx144, nx154, nx164, nx174, nx184, 
      nx194, nx204, nx214, nx224, nx234, nx244, nx254, nx264, nx274, nx284, 
      nx294, nx304, nx314, nx324, nx334, nx344, nx354, nx364, nx374, nx384, 
      nx394, nx404, nx414, nx424, nx535, nx537, nx539, nx541, nx543, nx545: 
   std_logic ;

begin
   q(31) <= q_31_EXMPLR ;
   q(30) <= q_30_EXMPLR ;
   q(29) <= q_29_EXMPLR ;
   q(28) <= q_28_EXMPLR ;
   q(27) <= q_27_EXMPLR ;
   q(26) <= q_26_EXMPLR ;
   q(25) <= q_25_EXMPLR ;
   q(24) <= q_24_EXMPLR ;
   q(23) <= q_23_EXMPLR ;
   q(22) <= q_22_EXMPLR ;
   q(21) <= q_21_EXMPLR ;
   q(20) <= q_20_EXMPLR ;
   q(19) <= q_19_EXMPLR ;
   q(18) <= q_18_EXMPLR ;
   q(17) <= q_17_EXMPLR ;
   q(16) <= q_16_EXMPLR ;
   q(15) <= q_15_EXMPLR ;
   q(14) <= q_14_EXMPLR ;
   q(13) <= q_13_EXMPLR ;
   q(12) <= q_12_EXMPLR ;
   q(11) <= q_11_EXMPLR ;
   q(10) <= q_10_EXMPLR ;
   q(9) <= q_9_EXMPLR ;
   q(8) <= q_8_EXMPLR ;
   q(7) <= q_7_EXMPLR ;
   q(6) <= q_6_EXMPLR ;
   q(5) <= q_5_EXMPLR ;
   q(4) <= q_4_EXMPLR ;
   q(3) <= q_3_EXMPLR ;
   q(2) <= q_2_EXMPLR ;
   q(1) <= q_1_EXMPLR ;
   q(0) <= q_0_EXMPLR ;
   reg_q_0 : dffr port map ( Q=>q_0_EXMPLR, QB=>OPEN, D=>nx114, CLK=>clk, R
      =>reset);
   ix115 : mux21_ni port map ( Y=>nx114, A0=>q_0_EXMPLR, A1=>d(0), S0=>nx537
   );
   reg_q_1 : dffr port map ( Q=>q_1_EXMPLR, QB=>OPEN, D=>nx124, CLK=>clk, R
      =>reset);
   ix125 : mux21_ni port map ( Y=>nx124, A0=>q_1_EXMPLR, A1=>d(1), S0=>nx537
   );
   reg_q_2 : dffr port map ( Q=>q_2_EXMPLR, QB=>OPEN, D=>nx134, CLK=>clk, R
      =>reset);
   ix135 : mux21_ni port map ( Y=>nx134, A0=>q_2_EXMPLR, A1=>d(2), S0=>nx537
   );
   reg_q_3 : dffr port map ( Q=>q_3_EXMPLR, QB=>OPEN, D=>nx144, CLK=>clk, R
      =>reset);
   ix145 : mux21_ni port map ( Y=>nx144, A0=>q_3_EXMPLR, A1=>d(3), S0=>nx537
   );
   reg_q_4 : dffr port map ( Q=>q_4_EXMPLR, QB=>OPEN, D=>nx154, CLK=>clk, R
      =>reset);
   ix155 : mux21_ni port map ( Y=>nx154, A0=>q_4_EXMPLR, A1=>d(4), S0=>nx537
   );
   reg_q_5 : dffr port map ( Q=>q_5_EXMPLR, QB=>OPEN, D=>nx164, CLK=>clk, R
      =>reset);
   ix165 : mux21_ni port map ( Y=>nx164, A0=>q_5_EXMPLR, A1=>d(5), S0=>nx537
   );
   reg_q_6 : dffr port map ( Q=>q_6_EXMPLR, QB=>OPEN, D=>nx174, CLK=>clk, R
      =>reset);
   ix175 : mux21_ni port map ( Y=>nx174, A0=>q_6_EXMPLR, A1=>d(6), S0=>nx537
   );
   reg_q_7 : dffr port map ( Q=>q_7_EXMPLR, QB=>OPEN, D=>nx184, CLK=>clk, R
      =>reset);
   ix185 : mux21_ni port map ( Y=>nx184, A0=>q_7_EXMPLR, A1=>d(7), S0=>nx539
   );
   reg_q_8 : dffr port map ( Q=>q_8_EXMPLR, QB=>OPEN, D=>nx194, CLK=>clk, R
      =>reset);
   ix195 : mux21_ni port map ( Y=>nx194, A0=>q_8_EXMPLR, A1=>d(8), S0=>nx539
   );
   reg_q_9 : dffr port map ( Q=>q_9_EXMPLR, QB=>OPEN, D=>nx204, CLK=>clk, R
      =>reset);
   ix205 : mux21_ni port map ( Y=>nx204, A0=>q_9_EXMPLR, A1=>d(9), S0=>nx539
   );
   reg_q_10 : dffr port map ( Q=>q_10_EXMPLR, QB=>OPEN, D=>nx214, CLK=>clk, 
      R=>reset);
   ix215 : mux21_ni port map ( Y=>nx214, A0=>q_10_EXMPLR, A1=>d(10), S0=>
      nx539);
   reg_q_11 : dffr port map ( Q=>q_11_EXMPLR, QB=>OPEN, D=>nx224, CLK=>clk, 
      R=>reset);
   ix225 : mux21_ni port map ( Y=>nx224, A0=>q_11_EXMPLR, A1=>d(11), S0=>
      nx539);
   reg_q_12 : dffr port map ( Q=>q_12_EXMPLR, QB=>OPEN, D=>nx234, CLK=>clk, 
      R=>reset);
   ix235 : mux21_ni port map ( Y=>nx234, A0=>q_12_EXMPLR, A1=>d(12), S0=>
      nx539);
   reg_q_13 : dffr port map ( Q=>q_13_EXMPLR, QB=>OPEN, D=>nx244, CLK=>clk, 
      R=>reset);
   ix245 : mux21_ni port map ( Y=>nx244, A0=>q_13_EXMPLR, A1=>d(13), S0=>
      nx539);
   reg_q_14 : dffr port map ( Q=>q_14_EXMPLR, QB=>OPEN, D=>nx254, CLK=>clk, 
      R=>reset);
   ix255 : mux21_ni port map ( Y=>nx254, A0=>q_14_EXMPLR, A1=>d(14), S0=>
      nx541);
   reg_q_15 : dffr port map ( Q=>q_15_EXMPLR, QB=>OPEN, D=>nx264, CLK=>clk, 
      R=>reset);
   ix265 : mux21_ni port map ( Y=>nx264, A0=>q_15_EXMPLR, A1=>d(15), S0=>
      nx541);
   reg_q_16 : dffr port map ( Q=>q_16_EXMPLR, QB=>OPEN, D=>nx274, CLK=>clk, 
      R=>reset);
   ix275 : mux21_ni port map ( Y=>nx274, A0=>q_16_EXMPLR, A1=>d(16), S0=>
      nx541);
   reg_q_17 : dffr port map ( Q=>q_17_EXMPLR, QB=>OPEN, D=>nx284, CLK=>clk, 
      R=>reset);
   ix285 : mux21_ni port map ( Y=>nx284, A0=>q_17_EXMPLR, A1=>d(17), S0=>
      nx541);
   reg_q_18 : dffr port map ( Q=>q_18_EXMPLR, QB=>OPEN, D=>nx294, CLK=>clk, 
      R=>reset);
   ix295 : mux21_ni port map ( Y=>nx294, A0=>q_18_EXMPLR, A1=>d(18), S0=>
      nx541);
   reg_q_19 : dffr port map ( Q=>q_19_EXMPLR, QB=>OPEN, D=>nx304, CLK=>clk, 
      R=>reset);
   ix305 : mux21_ni port map ( Y=>nx304, A0=>q_19_EXMPLR, A1=>d(19), S0=>
      nx541);
   reg_q_20 : dffr port map ( Q=>q_20_EXMPLR, QB=>OPEN, D=>nx314, CLK=>clk, 
      R=>reset);
   ix315 : mux21_ni port map ( Y=>nx314, A0=>q_20_EXMPLR, A1=>d(20), S0=>
      nx541);
   reg_q_21 : dffr port map ( Q=>q_21_EXMPLR, QB=>OPEN, D=>nx324, CLK=>clk, 
      R=>reset);
   ix325 : mux21_ni port map ( Y=>nx324, A0=>q_21_EXMPLR, A1=>d(21), S0=>
      nx543);
   reg_q_22 : dffr port map ( Q=>q_22_EXMPLR, QB=>OPEN, D=>nx334, CLK=>clk, 
      R=>reset);
   ix335 : mux21_ni port map ( Y=>nx334, A0=>q_22_EXMPLR, A1=>d(22), S0=>
      nx543);
   reg_q_23 : dffr port map ( Q=>q_23_EXMPLR, QB=>OPEN, D=>nx344, CLK=>clk, 
      R=>reset);
   ix345 : mux21_ni port map ( Y=>nx344, A0=>q_23_EXMPLR, A1=>d(23), S0=>
      nx543);
   reg_q_24 : dffr port map ( Q=>q_24_EXMPLR, QB=>OPEN, D=>nx354, CLK=>clk, 
      R=>reset);
   ix355 : mux21_ni port map ( Y=>nx354, A0=>q_24_EXMPLR, A1=>d(24), S0=>
      nx543);
   reg_q_25 : dffr port map ( Q=>q_25_EXMPLR, QB=>OPEN, D=>nx364, CLK=>clk, 
      R=>reset);
   ix365 : mux21_ni port map ( Y=>nx364, A0=>q_25_EXMPLR, A1=>d(25), S0=>
      nx543);
   reg_q_26 : dffr port map ( Q=>q_26_EXMPLR, QB=>OPEN, D=>nx374, CLK=>clk, 
      R=>reset);
   ix375 : mux21_ni port map ( Y=>nx374, A0=>q_26_EXMPLR, A1=>d(26), S0=>
      nx543);
   reg_q_27 : dffr port map ( Q=>q_27_EXMPLR, QB=>OPEN, D=>nx384, CLK=>clk, 
      R=>reset);
   ix385 : mux21_ni port map ( Y=>nx384, A0=>q_27_EXMPLR, A1=>d(27), S0=>
      nx543);
   reg_q_28 : dffr port map ( Q=>q_28_EXMPLR, QB=>OPEN, D=>nx394, CLK=>clk, 
      R=>reset);
   ix395 : mux21_ni port map ( Y=>nx394, A0=>q_28_EXMPLR, A1=>d(28), S0=>
      nx545);
   reg_q_29 : dffr port map ( Q=>q_29_EXMPLR, QB=>OPEN, D=>nx404, CLK=>clk, 
      R=>reset);
   ix405 : mux21_ni port map ( Y=>nx404, A0=>q_29_EXMPLR, A1=>d(29), S0=>
      nx545);
   reg_q_30 : dffr port map ( Q=>q_30_EXMPLR, QB=>OPEN, D=>nx414, CLK=>clk, 
      R=>reset);
   ix415 : mux21_ni port map ( Y=>nx414, A0=>q_30_EXMPLR, A1=>d(30), S0=>
      nx545);
   reg_q_31 : dffr port map ( Q=>q_31_EXMPLR, QB=>OPEN, D=>nx424, CLK=>clk, 
      R=>reset);
   ix425 : mux21_ni port map ( Y=>nx424, A0=>q_31_EXMPLR, A1=>d(31), S0=>
      nx545);
   ix534 : inv01 port map ( Y=>nx535, A=>load);
   ix536 : inv02 port map ( Y=>nx537, A=>nx535);
   ix538 : inv02 port map ( Y=>nx539, A=>nx535);
   ix540 : inv02 port map ( Y=>nx541, A=>nx535);
   ix542 : inv02 port map ( Y=>nx543, A=>nx535);
   ix544 : inv02 port map ( Y=>nx545, A=>nx535);
end Behavioral_unfold_3258 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity ComputationBlock is
   port (
      img_data_col_0 : IN std_logic_vector (15 DOWNTO 0) ;
      img_data_col_1 : IN std_logic_vector (15 DOWNTO 0) ;
      img_data_col_2 : IN std_logic_vector (15 DOWNTO 0) ;
      img_data_col_3 : IN std_logic_vector (15 DOWNTO 0) ;
      img_data_col_4 : IN std_logic_vector (15 DOWNTO 0) ;
      img_load : IN std_logic ;
      img_reset : IN std_logic ;
      filter_data_word : IN std_logic_vector (15 DOWNTO 0) ;
      filter_load : IN std_logic ;
      filter_reset : IN std_logic ;
      start : IN std_logic ;
      operation : IN std_logic ;
      compute_relu : IN std_logic ;
      filter_size : IN std_logic ;
      output1_init : IN std_logic_vector (15 DOWNTO 0) ;
      output2_init : IN std_logic_vector (15 DOWNTO 0) ;
      output1 : OUT std_logic_vector (15 DOWNTO 0) ;
      output2 : OUT std_logic_vector (15 DOWNTO 0) ;
      buffer_ready : OUT std_logic ;
      ready : OUT std_logic ;
      clk : IN std_logic ;
      en : IN std_logic ;
      reset : IN std_logic) ;
end ComputationBlock ;

architecture Structural_unfold_2968_0 of ComputationBlock is
   component ComputationPipeline
      port (
         img_data_0_15 : IN std_logic ;
         img_data_0_14 : IN std_logic ;
         img_data_0_13 : IN std_logic ;
         img_data_0_12 : IN std_logic ;
         img_data_0_11 : IN std_logic ;
         img_data_0_10 : IN std_logic ;
         img_data_0_9 : IN std_logic ;
         img_data_0_8 : IN std_logic ;
         img_data_0_7 : IN std_logic ;
         img_data_0_6 : IN std_logic ;
         img_data_0_5 : IN std_logic ;
         img_data_0_4 : IN std_logic ;
         img_data_0_3 : IN std_logic ;
         img_data_0_2 : IN std_logic ;
         img_data_0_1 : IN std_logic ;
         img_data_0_0 : IN std_logic ;
         img_data_1_15 : IN std_logic ;
         img_data_1_14 : IN std_logic ;
         img_data_1_13 : IN std_logic ;
         img_data_1_12 : IN std_logic ;
         img_data_1_11 : IN std_logic ;
         img_data_1_10 : IN std_logic ;
         img_data_1_9 : IN std_logic ;
         img_data_1_8 : IN std_logic ;
         img_data_1_7 : IN std_logic ;
         img_data_1_6 : IN std_logic ;
         img_data_1_5 : IN std_logic ;
         img_data_1_4 : IN std_logic ;
         img_data_1_3 : IN std_logic ;
         img_data_1_2 : IN std_logic ;
         img_data_1_1 : IN std_logic ;
         img_data_1_0 : IN std_logic ;
         img_data_2_15 : IN std_logic ;
         img_data_2_14 : IN std_logic ;
         img_data_2_13 : IN std_logic ;
         img_data_2_12 : IN std_logic ;
         img_data_2_11 : IN std_logic ;
         img_data_2_10 : IN std_logic ;
         img_data_2_9 : IN std_logic ;
         img_data_2_8 : IN std_logic ;
         img_data_2_7 : IN std_logic ;
         img_data_2_6 : IN std_logic ;
         img_data_2_5 : IN std_logic ;
         img_data_2_4 : IN std_logic ;
         img_data_2_3 : IN std_logic ;
         img_data_2_2 : IN std_logic ;
         img_data_2_1 : IN std_logic ;
         img_data_2_0 : IN std_logic ;
         img_data_3_15 : IN std_logic ;
         img_data_3_14 : IN std_logic ;
         img_data_3_13 : IN std_logic ;
         img_data_3_12 : IN std_logic ;
         img_data_3_11 : IN std_logic ;
         img_data_3_10 : IN std_logic ;
         img_data_3_9 : IN std_logic ;
         img_data_3_8 : IN std_logic ;
         img_data_3_7 : IN std_logic ;
         img_data_3_6 : IN std_logic ;
         img_data_3_5 : IN std_logic ;
         img_data_3_4 : IN std_logic ;
         img_data_3_3 : IN std_logic ;
         img_data_3_2 : IN std_logic ;
         img_data_3_1 : IN std_logic ;
         img_data_3_0 : IN std_logic ;
         img_data_4_15 : IN std_logic ;
         img_data_4_14 : IN std_logic ;
         img_data_4_13 : IN std_logic ;
         img_data_4_12 : IN std_logic ;
         img_data_4_11 : IN std_logic ;
         img_data_4_10 : IN std_logic ;
         img_data_4_9 : IN std_logic ;
         img_data_4_8 : IN std_logic ;
         img_data_4_7 : IN std_logic ;
         img_data_4_6 : IN std_logic ;
         img_data_4_5 : IN std_logic ;
         img_data_4_4 : IN std_logic ;
         img_data_4_3 : IN std_logic ;
         img_data_4_2 : IN std_logic ;
         img_data_4_1 : IN std_logic ;
         img_data_4_0 : IN std_logic ;
         img_data_5_15 : IN std_logic ;
         img_data_5_14 : IN std_logic ;
         img_data_5_13 : IN std_logic ;
         img_data_5_12 : IN std_logic ;
         img_data_5_11 : IN std_logic ;
         img_data_5_10 : IN std_logic ;
         img_data_5_9 : IN std_logic ;
         img_data_5_8 : IN std_logic ;
         img_data_5_7 : IN std_logic ;
         img_data_5_6 : IN std_logic ;
         img_data_5_5 : IN std_logic ;
         img_data_5_4 : IN std_logic ;
         img_data_5_3 : IN std_logic ;
         img_data_5_2 : IN std_logic ;
         img_data_5_1 : IN std_logic ;
         img_data_5_0 : IN std_logic ;
         img_data_6_15 : IN std_logic ;
         img_data_6_14 : IN std_logic ;
         img_data_6_13 : IN std_logic ;
         img_data_6_12 : IN std_logic ;
         img_data_6_11 : IN std_logic ;
         img_data_6_10 : IN std_logic ;
         img_data_6_9 : IN std_logic ;
         img_data_6_8 : IN std_logic ;
         img_data_6_7 : IN std_logic ;
         img_data_6_6 : IN std_logic ;
         img_data_6_5 : IN std_logic ;
         img_data_6_4 : IN std_logic ;
         img_data_6_3 : IN std_logic ;
         img_data_6_2 : IN std_logic ;
         img_data_6_1 : IN std_logic ;
         img_data_6_0 : IN std_logic ;
         img_data_7_15 : IN std_logic ;
         img_data_7_14 : IN std_logic ;
         img_data_7_13 : IN std_logic ;
         img_data_7_12 : IN std_logic ;
         img_data_7_11 : IN std_logic ;
         img_data_7_10 : IN std_logic ;
         img_data_7_9 : IN std_logic ;
         img_data_7_8 : IN std_logic ;
         img_data_7_7 : IN std_logic ;
         img_data_7_6 : IN std_logic ;
         img_data_7_5 : IN std_logic ;
         img_data_7_4 : IN std_logic ;
         img_data_7_3 : IN std_logic ;
         img_data_7_2 : IN std_logic ;
         img_data_7_1 : IN std_logic ;
         img_data_7_0 : IN std_logic ;
         img_data_8_15 : IN std_logic ;
         img_data_8_14 : IN std_logic ;
         img_data_8_13 : IN std_logic ;
         img_data_8_12 : IN std_logic ;
         img_data_8_11 : IN std_logic ;
         img_data_8_10 : IN std_logic ;
         img_data_8_9 : IN std_logic ;
         img_data_8_8 : IN std_logic ;
         img_data_8_7 : IN std_logic ;
         img_data_8_6 : IN std_logic ;
         img_data_8_5 : IN std_logic ;
         img_data_8_4 : IN std_logic ;
         img_data_8_3 : IN std_logic ;
         img_data_8_2 : IN std_logic ;
         img_data_8_1 : IN std_logic ;
         img_data_8_0 : IN std_logic ;
         img_data_9_15 : IN std_logic ;
         img_data_9_14 : IN std_logic ;
         img_data_9_13 : IN std_logic ;
         img_data_9_12 : IN std_logic ;
         img_data_9_11 : IN std_logic ;
         img_data_9_10 : IN std_logic ;
         img_data_9_9 : IN std_logic ;
         img_data_9_8 : IN std_logic ;
         img_data_9_7 : IN std_logic ;
         img_data_9_6 : IN std_logic ;
         img_data_9_5 : IN std_logic ;
         img_data_9_4 : IN std_logic ;
         img_data_9_3 : IN std_logic ;
         img_data_9_2 : IN std_logic ;
         img_data_9_1 : IN std_logic ;
         img_data_9_0 : IN std_logic ;
         img_data_10_15 : IN std_logic ;
         img_data_10_14 : IN std_logic ;
         img_data_10_13 : IN std_logic ;
         img_data_10_12 : IN std_logic ;
         img_data_10_11 : IN std_logic ;
         img_data_10_10 : IN std_logic ;
         img_data_10_9 : IN std_logic ;
         img_data_10_8 : IN std_logic ;
         img_data_10_7 : IN std_logic ;
         img_data_10_6 : IN std_logic ;
         img_data_10_5 : IN std_logic ;
         img_data_10_4 : IN std_logic ;
         img_data_10_3 : IN std_logic ;
         img_data_10_2 : IN std_logic ;
         img_data_10_1 : IN std_logic ;
         img_data_10_0 : IN std_logic ;
         img_data_11_15 : IN std_logic ;
         img_data_11_14 : IN std_logic ;
         img_data_11_13 : IN std_logic ;
         img_data_11_12 : IN std_logic ;
         img_data_11_11 : IN std_logic ;
         img_data_11_10 : IN std_logic ;
         img_data_11_9 : IN std_logic ;
         img_data_11_8 : IN std_logic ;
         img_data_11_7 : IN std_logic ;
         img_data_11_6 : IN std_logic ;
         img_data_11_5 : IN std_logic ;
         img_data_11_4 : IN std_logic ;
         img_data_11_3 : IN std_logic ;
         img_data_11_2 : IN std_logic ;
         img_data_11_1 : IN std_logic ;
         img_data_11_0 : IN std_logic ;
         img_data_12_15 : IN std_logic ;
         img_data_12_14 : IN std_logic ;
         img_data_12_13 : IN std_logic ;
         img_data_12_12 : IN std_logic ;
         img_data_12_11 : IN std_logic ;
         img_data_12_10 : IN std_logic ;
         img_data_12_9 : IN std_logic ;
         img_data_12_8 : IN std_logic ;
         img_data_12_7 : IN std_logic ;
         img_data_12_6 : IN std_logic ;
         img_data_12_5 : IN std_logic ;
         img_data_12_4 : IN std_logic ;
         img_data_12_3 : IN std_logic ;
         img_data_12_2 : IN std_logic ;
         img_data_12_1 : IN std_logic ;
         img_data_12_0 : IN std_logic ;
         img_data_13_15 : IN std_logic ;
         img_data_13_14 : IN std_logic ;
         img_data_13_13 : IN std_logic ;
         img_data_13_12 : IN std_logic ;
         img_data_13_11 : IN std_logic ;
         img_data_13_10 : IN std_logic ;
         img_data_13_9 : IN std_logic ;
         img_data_13_8 : IN std_logic ;
         img_data_13_7 : IN std_logic ;
         img_data_13_6 : IN std_logic ;
         img_data_13_5 : IN std_logic ;
         img_data_13_4 : IN std_logic ;
         img_data_13_3 : IN std_logic ;
         img_data_13_2 : IN std_logic ;
         img_data_13_1 : IN std_logic ;
         img_data_13_0 : IN std_logic ;
         img_data_14_15 : IN std_logic ;
         img_data_14_14 : IN std_logic ;
         img_data_14_13 : IN std_logic ;
         img_data_14_12 : IN std_logic ;
         img_data_14_11 : IN std_logic ;
         img_data_14_10 : IN std_logic ;
         img_data_14_9 : IN std_logic ;
         img_data_14_8 : IN std_logic ;
         img_data_14_7 : IN std_logic ;
         img_data_14_6 : IN std_logic ;
         img_data_14_5 : IN std_logic ;
         img_data_14_4 : IN std_logic ;
         img_data_14_3 : IN std_logic ;
         img_data_14_2 : IN std_logic ;
         img_data_14_1 : IN std_logic ;
         img_data_14_0 : IN std_logic ;
         img_data_15_15 : IN std_logic ;
         img_data_15_14 : IN std_logic ;
         img_data_15_13 : IN std_logic ;
         img_data_15_12 : IN std_logic ;
         img_data_15_11 : IN std_logic ;
         img_data_15_10 : IN std_logic ;
         img_data_15_9 : IN std_logic ;
         img_data_15_8 : IN std_logic ;
         img_data_15_7 : IN std_logic ;
         img_data_15_6 : IN std_logic ;
         img_data_15_5 : IN std_logic ;
         img_data_15_4 : IN std_logic ;
         img_data_15_3 : IN std_logic ;
         img_data_15_2 : IN std_logic ;
         img_data_15_1 : IN std_logic ;
         img_data_15_0 : IN std_logic ;
         img_data_16_15 : IN std_logic ;
         img_data_16_14 : IN std_logic ;
         img_data_16_13 : IN std_logic ;
         img_data_16_12 : IN std_logic ;
         img_data_16_11 : IN std_logic ;
         img_data_16_10 : IN std_logic ;
         img_data_16_9 : IN std_logic ;
         img_data_16_8 : IN std_logic ;
         img_data_16_7 : IN std_logic ;
         img_data_16_6 : IN std_logic ;
         img_data_16_5 : IN std_logic ;
         img_data_16_4 : IN std_logic ;
         img_data_16_3 : IN std_logic ;
         img_data_16_2 : IN std_logic ;
         img_data_16_1 : IN std_logic ;
         img_data_16_0 : IN std_logic ;
         img_data_17_15 : IN std_logic ;
         img_data_17_14 : IN std_logic ;
         img_data_17_13 : IN std_logic ;
         img_data_17_12 : IN std_logic ;
         img_data_17_11 : IN std_logic ;
         img_data_17_10 : IN std_logic ;
         img_data_17_9 : IN std_logic ;
         img_data_17_8 : IN std_logic ;
         img_data_17_7 : IN std_logic ;
         img_data_17_6 : IN std_logic ;
         img_data_17_5 : IN std_logic ;
         img_data_17_4 : IN std_logic ;
         img_data_17_3 : IN std_logic ;
         img_data_17_2 : IN std_logic ;
         img_data_17_1 : IN std_logic ;
         img_data_17_0 : IN std_logic ;
         img_data_18_15 : IN std_logic ;
         img_data_18_14 : IN std_logic ;
         img_data_18_13 : IN std_logic ;
         img_data_18_12 : IN std_logic ;
         img_data_18_11 : IN std_logic ;
         img_data_18_10 : IN std_logic ;
         img_data_18_9 : IN std_logic ;
         img_data_18_8 : IN std_logic ;
         img_data_18_7 : IN std_logic ;
         img_data_18_6 : IN std_logic ;
         img_data_18_5 : IN std_logic ;
         img_data_18_4 : IN std_logic ;
         img_data_18_3 : IN std_logic ;
         img_data_18_2 : IN std_logic ;
         img_data_18_1 : IN std_logic ;
         img_data_18_0 : IN std_logic ;
         img_data_19_15 : IN std_logic ;
         img_data_19_14 : IN std_logic ;
         img_data_19_13 : IN std_logic ;
         img_data_19_12 : IN std_logic ;
         img_data_19_11 : IN std_logic ;
         img_data_19_10 : IN std_logic ;
         img_data_19_9 : IN std_logic ;
         img_data_19_8 : IN std_logic ;
         img_data_19_7 : IN std_logic ;
         img_data_19_6 : IN std_logic ;
         img_data_19_5 : IN std_logic ;
         img_data_19_4 : IN std_logic ;
         img_data_19_3 : IN std_logic ;
         img_data_19_2 : IN std_logic ;
         img_data_19_1 : IN std_logic ;
         img_data_19_0 : IN std_logic ;
         img_data_20_15 : IN std_logic ;
         img_data_20_14 : IN std_logic ;
         img_data_20_13 : IN std_logic ;
         img_data_20_12 : IN std_logic ;
         img_data_20_11 : IN std_logic ;
         img_data_20_10 : IN std_logic ;
         img_data_20_9 : IN std_logic ;
         img_data_20_8 : IN std_logic ;
         img_data_20_7 : IN std_logic ;
         img_data_20_6 : IN std_logic ;
         img_data_20_5 : IN std_logic ;
         img_data_20_4 : IN std_logic ;
         img_data_20_3 : IN std_logic ;
         img_data_20_2 : IN std_logic ;
         img_data_20_1 : IN std_logic ;
         img_data_20_0 : IN std_logic ;
         img_data_21_15 : IN std_logic ;
         img_data_21_14 : IN std_logic ;
         img_data_21_13 : IN std_logic ;
         img_data_21_12 : IN std_logic ;
         img_data_21_11 : IN std_logic ;
         img_data_21_10 : IN std_logic ;
         img_data_21_9 : IN std_logic ;
         img_data_21_8 : IN std_logic ;
         img_data_21_7 : IN std_logic ;
         img_data_21_6 : IN std_logic ;
         img_data_21_5 : IN std_logic ;
         img_data_21_4 : IN std_logic ;
         img_data_21_3 : IN std_logic ;
         img_data_21_2 : IN std_logic ;
         img_data_21_1 : IN std_logic ;
         img_data_21_0 : IN std_logic ;
         img_data_22_15 : IN std_logic ;
         img_data_22_14 : IN std_logic ;
         img_data_22_13 : IN std_logic ;
         img_data_22_12 : IN std_logic ;
         img_data_22_11 : IN std_logic ;
         img_data_22_10 : IN std_logic ;
         img_data_22_9 : IN std_logic ;
         img_data_22_8 : IN std_logic ;
         img_data_22_7 : IN std_logic ;
         img_data_22_6 : IN std_logic ;
         img_data_22_5 : IN std_logic ;
         img_data_22_4 : IN std_logic ;
         img_data_22_3 : IN std_logic ;
         img_data_22_2 : IN std_logic ;
         img_data_22_1 : IN std_logic ;
         img_data_22_0 : IN std_logic ;
         img_data_23_15 : IN std_logic ;
         img_data_23_14 : IN std_logic ;
         img_data_23_13 : IN std_logic ;
         img_data_23_12 : IN std_logic ;
         img_data_23_11 : IN std_logic ;
         img_data_23_10 : IN std_logic ;
         img_data_23_9 : IN std_logic ;
         img_data_23_8 : IN std_logic ;
         img_data_23_7 : IN std_logic ;
         img_data_23_6 : IN std_logic ;
         img_data_23_5 : IN std_logic ;
         img_data_23_4 : IN std_logic ;
         img_data_23_3 : IN std_logic ;
         img_data_23_2 : IN std_logic ;
         img_data_23_1 : IN std_logic ;
         img_data_23_0 : IN std_logic ;
         img_data_24_15 : IN std_logic ;
         img_data_24_14 : IN std_logic ;
         img_data_24_13 : IN std_logic ;
         img_data_24_12 : IN std_logic ;
         img_data_24_11 : IN std_logic ;
         img_data_24_10 : IN std_logic ;
         img_data_24_9 : IN std_logic ;
         img_data_24_8 : IN std_logic ;
         img_data_24_7 : IN std_logic ;
         img_data_24_6 : IN std_logic ;
         img_data_24_5 : IN std_logic ;
         img_data_24_4 : IN std_logic ;
         img_data_24_3 : IN std_logic ;
         img_data_24_2 : IN std_logic ;
         img_data_24_1 : IN std_logic ;
         img_data_24_0 : IN std_logic ;
         filter_data_0_15 : IN std_logic ;
         filter_data_0_14 : IN std_logic ;
         filter_data_0_13 : IN std_logic ;
         filter_data_0_12 : IN std_logic ;
         filter_data_0_11 : IN std_logic ;
         filter_data_0_10 : IN std_logic ;
         filter_data_0_9 : IN std_logic ;
         filter_data_0_8 : IN std_logic ;
         filter_data_0_7 : IN std_logic ;
         filter_data_0_6 : IN std_logic ;
         filter_data_0_5 : IN std_logic ;
         filter_data_0_4 : IN std_logic ;
         filter_data_0_3 : IN std_logic ;
         filter_data_0_2 : IN std_logic ;
         filter_data_0_1 : IN std_logic ;
         filter_data_0_0 : IN std_logic ;
         filter_data_1_15 : IN std_logic ;
         filter_data_1_14 : IN std_logic ;
         filter_data_1_13 : IN std_logic ;
         filter_data_1_12 : IN std_logic ;
         filter_data_1_11 : IN std_logic ;
         filter_data_1_10 : IN std_logic ;
         filter_data_1_9 : IN std_logic ;
         filter_data_1_8 : IN std_logic ;
         filter_data_1_7 : IN std_logic ;
         filter_data_1_6 : IN std_logic ;
         filter_data_1_5 : IN std_logic ;
         filter_data_1_4 : IN std_logic ;
         filter_data_1_3 : IN std_logic ;
         filter_data_1_2 : IN std_logic ;
         filter_data_1_1 : IN std_logic ;
         filter_data_1_0 : IN std_logic ;
         filter_data_2_15 : IN std_logic ;
         filter_data_2_14 : IN std_logic ;
         filter_data_2_13 : IN std_logic ;
         filter_data_2_12 : IN std_logic ;
         filter_data_2_11 : IN std_logic ;
         filter_data_2_10 : IN std_logic ;
         filter_data_2_9 : IN std_logic ;
         filter_data_2_8 : IN std_logic ;
         filter_data_2_7 : IN std_logic ;
         filter_data_2_6 : IN std_logic ;
         filter_data_2_5 : IN std_logic ;
         filter_data_2_4 : IN std_logic ;
         filter_data_2_3 : IN std_logic ;
         filter_data_2_2 : IN std_logic ;
         filter_data_2_1 : IN std_logic ;
         filter_data_2_0 : IN std_logic ;
         filter_data_3_15 : IN std_logic ;
         filter_data_3_14 : IN std_logic ;
         filter_data_3_13 : IN std_logic ;
         filter_data_3_12 : IN std_logic ;
         filter_data_3_11 : IN std_logic ;
         filter_data_3_10 : IN std_logic ;
         filter_data_3_9 : IN std_logic ;
         filter_data_3_8 : IN std_logic ;
         filter_data_3_7 : IN std_logic ;
         filter_data_3_6 : IN std_logic ;
         filter_data_3_5 : IN std_logic ;
         filter_data_3_4 : IN std_logic ;
         filter_data_3_3 : IN std_logic ;
         filter_data_3_2 : IN std_logic ;
         filter_data_3_1 : IN std_logic ;
         filter_data_3_0 : IN std_logic ;
         filter_data_4_15 : IN std_logic ;
         filter_data_4_14 : IN std_logic ;
         filter_data_4_13 : IN std_logic ;
         filter_data_4_12 : IN std_logic ;
         filter_data_4_11 : IN std_logic ;
         filter_data_4_10 : IN std_logic ;
         filter_data_4_9 : IN std_logic ;
         filter_data_4_8 : IN std_logic ;
         filter_data_4_7 : IN std_logic ;
         filter_data_4_6 : IN std_logic ;
         filter_data_4_5 : IN std_logic ;
         filter_data_4_4 : IN std_logic ;
         filter_data_4_3 : IN std_logic ;
         filter_data_4_2 : IN std_logic ;
         filter_data_4_1 : IN std_logic ;
         filter_data_4_0 : IN std_logic ;
         filter_data_5_15 : IN std_logic ;
         filter_data_5_14 : IN std_logic ;
         filter_data_5_13 : IN std_logic ;
         filter_data_5_12 : IN std_logic ;
         filter_data_5_11 : IN std_logic ;
         filter_data_5_10 : IN std_logic ;
         filter_data_5_9 : IN std_logic ;
         filter_data_5_8 : IN std_logic ;
         filter_data_5_7 : IN std_logic ;
         filter_data_5_6 : IN std_logic ;
         filter_data_5_5 : IN std_logic ;
         filter_data_5_4 : IN std_logic ;
         filter_data_5_3 : IN std_logic ;
         filter_data_5_2 : IN std_logic ;
         filter_data_5_1 : IN std_logic ;
         filter_data_5_0 : IN std_logic ;
         filter_data_6_15 : IN std_logic ;
         filter_data_6_14 : IN std_logic ;
         filter_data_6_13 : IN std_logic ;
         filter_data_6_12 : IN std_logic ;
         filter_data_6_11 : IN std_logic ;
         filter_data_6_10 : IN std_logic ;
         filter_data_6_9 : IN std_logic ;
         filter_data_6_8 : IN std_logic ;
         filter_data_6_7 : IN std_logic ;
         filter_data_6_6 : IN std_logic ;
         filter_data_6_5 : IN std_logic ;
         filter_data_6_4 : IN std_logic ;
         filter_data_6_3 : IN std_logic ;
         filter_data_6_2 : IN std_logic ;
         filter_data_6_1 : IN std_logic ;
         filter_data_6_0 : IN std_logic ;
         filter_data_7_15 : IN std_logic ;
         filter_data_7_14 : IN std_logic ;
         filter_data_7_13 : IN std_logic ;
         filter_data_7_12 : IN std_logic ;
         filter_data_7_11 : IN std_logic ;
         filter_data_7_10 : IN std_logic ;
         filter_data_7_9 : IN std_logic ;
         filter_data_7_8 : IN std_logic ;
         filter_data_7_7 : IN std_logic ;
         filter_data_7_6 : IN std_logic ;
         filter_data_7_5 : IN std_logic ;
         filter_data_7_4 : IN std_logic ;
         filter_data_7_3 : IN std_logic ;
         filter_data_7_2 : IN std_logic ;
         filter_data_7_1 : IN std_logic ;
         filter_data_7_0 : IN std_logic ;
         filter_data_8_15 : IN std_logic ;
         filter_data_8_14 : IN std_logic ;
         filter_data_8_13 : IN std_logic ;
         filter_data_8_12 : IN std_logic ;
         filter_data_8_11 : IN std_logic ;
         filter_data_8_10 : IN std_logic ;
         filter_data_8_9 : IN std_logic ;
         filter_data_8_8 : IN std_logic ;
         filter_data_8_7 : IN std_logic ;
         filter_data_8_6 : IN std_logic ;
         filter_data_8_5 : IN std_logic ;
         filter_data_8_4 : IN std_logic ;
         filter_data_8_3 : IN std_logic ;
         filter_data_8_2 : IN std_logic ;
         filter_data_8_1 : IN std_logic ;
         filter_data_8_0 : IN std_logic ;
         filter_data_9_15 : IN std_logic ;
         filter_data_9_14 : IN std_logic ;
         filter_data_9_13 : IN std_logic ;
         filter_data_9_12 : IN std_logic ;
         filter_data_9_11 : IN std_logic ;
         filter_data_9_10 : IN std_logic ;
         filter_data_9_9 : IN std_logic ;
         filter_data_9_8 : IN std_logic ;
         filter_data_9_7 : IN std_logic ;
         filter_data_9_6 : IN std_logic ;
         filter_data_9_5 : IN std_logic ;
         filter_data_9_4 : IN std_logic ;
         filter_data_9_3 : IN std_logic ;
         filter_data_9_2 : IN std_logic ;
         filter_data_9_1 : IN std_logic ;
         filter_data_9_0 : IN std_logic ;
         filter_data_10_15 : IN std_logic ;
         filter_data_10_14 : IN std_logic ;
         filter_data_10_13 : IN std_logic ;
         filter_data_10_12 : IN std_logic ;
         filter_data_10_11 : IN std_logic ;
         filter_data_10_10 : IN std_logic ;
         filter_data_10_9 : IN std_logic ;
         filter_data_10_8 : IN std_logic ;
         filter_data_10_7 : IN std_logic ;
         filter_data_10_6 : IN std_logic ;
         filter_data_10_5 : IN std_logic ;
         filter_data_10_4 : IN std_logic ;
         filter_data_10_3 : IN std_logic ;
         filter_data_10_2 : IN std_logic ;
         filter_data_10_1 : IN std_logic ;
         filter_data_10_0 : IN std_logic ;
         filter_data_11_15 : IN std_logic ;
         filter_data_11_14 : IN std_logic ;
         filter_data_11_13 : IN std_logic ;
         filter_data_11_12 : IN std_logic ;
         filter_data_11_11 : IN std_logic ;
         filter_data_11_10 : IN std_logic ;
         filter_data_11_9 : IN std_logic ;
         filter_data_11_8 : IN std_logic ;
         filter_data_11_7 : IN std_logic ;
         filter_data_11_6 : IN std_logic ;
         filter_data_11_5 : IN std_logic ;
         filter_data_11_4 : IN std_logic ;
         filter_data_11_3 : IN std_logic ;
         filter_data_11_2 : IN std_logic ;
         filter_data_11_1 : IN std_logic ;
         filter_data_11_0 : IN std_logic ;
         filter_data_12_15 : IN std_logic ;
         filter_data_12_14 : IN std_logic ;
         filter_data_12_13 : IN std_logic ;
         filter_data_12_12 : IN std_logic ;
         filter_data_12_11 : IN std_logic ;
         filter_data_12_10 : IN std_logic ;
         filter_data_12_9 : IN std_logic ;
         filter_data_12_8 : IN std_logic ;
         filter_data_12_7 : IN std_logic ;
         filter_data_12_6 : IN std_logic ;
         filter_data_12_5 : IN std_logic ;
         filter_data_12_4 : IN std_logic ;
         filter_data_12_3 : IN std_logic ;
         filter_data_12_2 : IN std_logic ;
         filter_data_12_1 : IN std_logic ;
         filter_data_12_0 : IN std_logic ;
         filter_data_13_15 : IN std_logic ;
         filter_data_13_14 : IN std_logic ;
         filter_data_13_13 : IN std_logic ;
         filter_data_13_12 : IN std_logic ;
         filter_data_13_11 : IN std_logic ;
         filter_data_13_10 : IN std_logic ;
         filter_data_13_9 : IN std_logic ;
         filter_data_13_8 : IN std_logic ;
         filter_data_13_7 : IN std_logic ;
         filter_data_13_6 : IN std_logic ;
         filter_data_13_5 : IN std_logic ;
         filter_data_13_4 : IN std_logic ;
         filter_data_13_3 : IN std_logic ;
         filter_data_13_2 : IN std_logic ;
         filter_data_13_1 : IN std_logic ;
         filter_data_13_0 : IN std_logic ;
         filter_data_14_15 : IN std_logic ;
         filter_data_14_14 : IN std_logic ;
         filter_data_14_13 : IN std_logic ;
         filter_data_14_12 : IN std_logic ;
         filter_data_14_11 : IN std_logic ;
         filter_data_14_10 : IN std_logic ;
         filter_data_14_9 : IN std_logic ;
         filter_data_14_8 : IN std_logic ;
         filter_data_14_7 : IN std_logic ;
         filter_data_14_6 : IN std_logic ;
         filter_data_14_5 : IN std_logic ;
         filter_data_14_4 : IN std_logic ;
         filter_data_14_3 : IN std_logic ;
         filter_data_14_2 : IN std_logic ;
         filter_data_14_1 : IN std_logic ;
         filter_data_14_0 : IN std_logic ;
         filter_data_15_15 : IN std_logic ;
         filter_data_15_14 : IN std_logic ;
         filter_data_15_13 : IN std_logic ;
         filter_data_15_12 : IN std_logic ;
         filter_data_15_11 : IN std_logic ;
         filter_data_15_10 : IN std_logic ;
         filter_data_15_9 : IN std_logic ;
         filter_data_15_8 : IN std_logic ;
         filter_data_15_7 : IN std_logic ;
         filter_data_15_6 : IN std_logic ;
         filter_data_15_5 : IN std_logic ;
         filter_data_15_4 : IN std_logic ;
         filter_data_15_3 : IN std_logic ;
         filter_data_15_2 : IN std_logic ;
         filter_data_15_1 : IN std_logic ;
         filter_data_15_0 : IN std_logic ;
         filter_data_16_15 : IN std_logic ;
         filter_data_16_14 : IN std_logic ;
         filter_data_16_13 : IN std_logic ;
         filter_data_16_12 : IN std_logic ;
         filter_data_16_11 : IN std_logic ;
         filter_data_16_10 : IN std_logic ;
         filter_data_16_9 : IN std_logic ;
         filter_data_16_8 : IN std_logic ;
         filter_data_16_7 : IN std_logic ;
         filter_data_16_6 : IN std_logic ;
         filter_data_16_5 : IN std_logic ;
         filter_data_16_4 : IN std_logic ;
         filter_data_16_3 : IN std_logic ;
         filter_data_16_2 : IN std_logic ;
         filter_data_16_1 : IN std_logic ;
         filter_data_16_0 : IN std_logic ;
         filter_data_17_15 : IN std_logic ;
         filter_data_17_14 : IN std_logic ;
         filter_data_17_13 : IN std_logic ;
         filter_data_17_12 : IN std_logic ;
         filter_data_17_11 : IN std_logic ;
         filter_data_17_10 : IN std_logic ;
         filter_data_17_9 : IN std_logic ;
         filter_data_17_8 : IN std_logic ;
         filter_data_17_7 : IN std_logic ;
         filter_data_17_6 : IN std_logic ;
         filter_data_17_5 : IN std_logic ;
         filter_data_17_4 : IN std_logic ;
         filter_data_17_3 : IN std_logic ;
         filter_data_17_2 : IN std_logic ;
         filter_data_17_1 : IN std_logic ;
         filter_data_17_0 : IN std_logic ;
         filter_data_18_15 : IN std_logic ;
         filter_data_18_14 : IN std_logic ;
         filter_data_18_13 : IN std_logic ;
         filter_data_18_12 : IN std_logic ;
         filter_data_18_11 : IN std_logic ;
         filter_data_18_10 : IN std_logic ;
         filter_data_18_9 : IN std_logic ;
         filter_data_18_8 : IN std_logic ;
         filter_data_18_7 : IN std_logic ;
         filter_data_18_6 : IN std_logic ;
         filter_data_18_5 : IN std_logic ;
         filter_data_18_4 : IN std_logic ;
         filter_data_18_3 : IN std_logic ;
         filter_data_18_2 : IN std_logic ;
         filter_data_18_1 : IN std_logic ;
         filter_data_18_0 : IN std_logic ;
         filter_data_19_15 : IN std_logic ;
         filter_data_19_14 : IN std_logic ;
         filter_data_19_13 : IN std_logic ;
         filter_data_19_12 : IN std_logic ;
         filter_data_19_11 : IN std_logic ;
         filter_data_19_10 : IN std_logic ;
         filter_data_19_9 : IN std_logic ;
         filter_data_19_8 : IN std_logic ;
         filter_data_19_7 : IN std_logic ;
         filter_data_19_6 : IN std_logic ;
         filter_data_19_5 : IN std_logic ;
         filter_data_19_4 : IN std_logic ;
         filter_data_19_3 : IN std_logic ;
         filter_data_19_2 : IN std_logic ;
         filter_data_19_1 : IN std_logic ;
         filter_data_19_0 : IN std_logic ;
         filter_data_20_15 : IN std_logic ;
         filter_data_20_14 : IN std_logic ;
         filter_data_20_13 : IN std_logic ;
         filter_data_20_12 : IN std_logic ;
         filter_data_20_11 : IN std_logic ;
         filter_data_20_10 : IN std_logic ;
         filter_data_20_9 : IN std_logic ;
         filter_data_20_8 : IN std_logic ;
         filter_data_20_7 : IN std_logic ;
         filter_data_20_6 : IN std_logic ;
         filter_data_20_5 : IN std_logic ;
         filter_data_20_4 : IN std_logic ;
         filter_data_20_3 : IN std_logic ;
         filter_data_20_2 : IN std_logic ;
         filter_data_20_1 : IN std_logic ;
         filter_data_20_0 : IN std_logic ;
         filter_data_21_15 : IN std_logic ;
         filter_data_21_14 : IN std_logic ;
         filter_data_21_13 : IN std_logic ;
         filter_data_21_12 : IN std_logic ;
         filter_data_21_11 : IN std_logic ;
         filter_data_21_10 : IN std_logic ;
         filter_data_21_9 : IN std_logic ;
         filter_data_21_8 : IN std_logic ;
         filter_data_21_7 : IN std_logic ;
         filter_data_21_6 : IN std_logic ;
         filter_data_21_5 : IN std_logic ;
         filter_data_21_4 : IN std_logic ;
         filter_data_21_3 : IN std_logic ;
         filter_data_21_2 : IN std_logic ;
         filter_data_21_1 : IN std_logic ;
         filter_data_21_0 : IN std_logic ;
         filter_data_22_15 : IN std_logic ;
         filter_data_22_14 : IN std_logic ;
         filter_data_22_13 : IN std_logic ;
         filter_data_22_12 : IN std_logic ;
         filter_data_22_11 : IN std_logic ;
         filter_data_22_10 : IN std_logic ;
         filter_data_22_9 : IN std_logic ;
         filter_data_22_8 : IN std_logic ;
         filter_data_22_7 : IN std_logic ;
         filter_data_22_6 : IN std_logic ;
         filter_data_22_5 : IN std_logic ;
         filter_data_22_4 : IN std_logic ;
         filter_data_22_3 : IN std_logic ;
         filter_data_22_2 : IN std_logic ;
         filter_data_22_1 : IN std_logic ;
         filter_data_22_0 : IN std_logic ;
         filter_data_23_15 : IN std_logic ;
         filter_data_23_14 : IN std_logic ;
         filter_data_23_13 : IN std_logic ;
         filter_data_23_12 : IN std_logic ;
         filter_data_23_11 : IN std_logic ;
         filter_data_23_10 : IN std_logic ;
         filter_data_23_9 : IN std_logic ;
         filter_data_23_8 : IN std_logic ;
         filter_data_23_7 : IN std_logic ;
         filter_data_23_6 : IN std_logic ;
         filter_data_23_5 : IN std_logic ;
         filter_data_23_4 : IN std_logic ;
         filter_data_23_3 : IN std_logic ;
         filter_data_23_2 : IN std_logic ;
         filter_data_23_1 : IN std_logic ;
         filter_data_23_0 : IN std_logic ;
         filter_data_24_15 : IN std_logic ;
         filter_data_24_14 : IN std_logic ;
         filter_data_24_13 : IN std_logic ;
         filter_data_24_12 : IN std_logic ;
         filter_data_24_11 : IN std_logic ;
         filter_data_24_10 : IN std_logic ;
         filter_data_24_9 : IN std_logic ;
         filter_data_24_8 : IN std_logic ;
         filter_data_24_7 : IN std_logic ;
         filter_data_24_6 : IN std_logic ;
         filter_data_24_5 : IN std_logic ;
         filter_data_24_4 : IN std_logic ;
         filter_data_24_3 : IN std_logic ;
         filter_data_24_2 : IN std_logic ;
         filter_data_24_1 : IN std_logic ;
         filter_data_24_0 : IN std_logic ;
         d_arr_0_31 : OUT std_logic ;
         d_arr_0_30 : OUT std_logic ;
         d_arr_0_29 : OUT std_logic ;
         d_arr_0_28 : OUT std_logic ;
         d_arr_0_27 : OUT std_logic ;
         d_arr_0_26 : OUT std_logic ;
         d_arr_0_25 : OUT std_logic ;
         d_arr_0_24 : OUT std_logic ;
         d_arr_0_23 : OUT std_logic ;
         d_arr_0_22 : OUT std_logic ;
         d_arr_0_21 : OUT std_logic ;
         d_arr_0_20 : OUT std_logic ;
         d_arr_0_19 : OUT std_logic ;
         d_arr_0_18 : OUT std_logic ;
         d_arr_0_17 : OUT std_logic ;
         d_arr_0_16 : OUT std_logic ;
         d_arr_0_15 : OUT std_logic ;
         d_arr_0_14 : OUT std_logic ;
         d_arr_0_13 : OUT std_logic ;
         d_arr_0_12 : OUT std_logic ;
         d_arr_0_11 : OUT std_logic ;
         d_arr_0_10 : OUT std_logic ;
         d_arr_0_9 : OUT std_logic ;
         d_arr_0_8 : OUT std_logic ;
         d_arr_0_7 : OUT std_logic ;
         d_arr_0_6 : OUT std_logic ;
         d_arr_0_5 : OUT std_logic ;
         d_arr_0_4 : OUT std_logic ;
         d_arr_0_3 : OUT std_logic ;
         d_arr_0_2 : OUT std_logic ;
         d_arr_0_1 : OUT std_logic ;
         d_arr_0_0 : OUT std_logic ;
         d_arr_1_31 : OUT std_logic ;
         d_arr_1_30 : OUT std_logic ;
         d_arr_1_29 : OUT std_logic ;
         d_arr_1_28 : OUT std_logic ;
         d_arr_1_27 : OUT std_logic ;
         d_arr_1_26 : OUT std_logic ;
         d_arr_1_25 : OUT std_logic ;
         d_arr_1_24 : OUT std_logic ;
         d_arr_1_23 : OUT std_logic ;
         d_arr_1_22 : OUT std_logic ;
         d_arr_1_21 : OUT std_logic ;
         d_arr_1_20 : OUT std_logic ;
         d_arr_1_19 : OUT std_logic ;
         d_arr_1_18 : OUT std_logic ;
         d_arr_1_17 : OUT std_logic ;
         d_arr_1_16 : OUT std_logic ;
         d_arr_1_15 : OUT std_logic ;
         d_arr_1_14 : OUT std_logic ;
         d_arr_1_13 : OUT std_logic ;
         d_arr_1_12 : OUT std_logic ;
         d_arr_1_11 : OUT std_logic ;
         d_arr_1_10 : OUT std_logic ;
         d_arr_1_9 : OUT std_logic ;
         d_arr_1_8 : OUT std_logic ;
         d_arr_1_7 : OUT std_logic ;
         d_arr_1_6 : OUT std_logic ;
         d_arr_1_5 : OUT std_logic ;
         d_arr_1_4 : OUT std_logic ;
         d_arr_1_3 : OUT std_logic ;
         d_arr_1_2 : OUT std_logic ;
         d_arr_1_1 : OUT std_logic ;
         d_arr_1_0 : OUT std_logic ;
         d_arr_2_31 : OUT std_logic ;
         d_arr_2_30 : OUT std_logic ;
         d_arr_2_29 : OUT std_logic ;
         d_arr_2_28 : OUT std_logic ;
         d_arr_2_27 : OUT std_logic ;
         d_arr_2_26 : OUT std_logic ;
         d_arr_2_25 : OUT std_logic ;
         d_arr_2_24 : OUT std_logic ;
         d_arr_2_23 : OUT std_logic ;
         d_arr_2_22 : OUT std_logic ;
         d_arr_2_21 : OUT std_logic ;
         d_arr_2_20 : OUT std_logic ;
         d_arr_2_19 : OUT std_logic ;
         d_arr_2_18 : OUT std_logic ;
         d_arr_2_17 : OUT std_logic ;
         d_arr_2_16 : OUT std_logic ;
         d_arr_2_15 : OUT std_logic ;
         d_arr_2_14 : OUT std_logic ;
         d_arr_2_13 : OUT std_logic ;
         d_arr_2_12 : OUT std_logic ;
         d_arr_2_11 : OUT std_logic ;
         d_arr_2_10 : OUT std_logic ;
         d_arr_2_9 : OUT std_logic ;
         d_arr_2_8 : OUT std_logic ;
         d_arr_2_7 : OUT std_logic ;
         d_arr_2_6 : OUT std_logic ;
         d_arr_2_5 : OUT std_logic ;
         d_arr_2_4 : OUT std_logic ;
         d_arr_2_3 : OUT std_logic ;
         d_arr_2_2 : OUT std_logic ;
         d_arr_2_1 : OUT std_logic ;
         d_arr_2_0 : OUT std_logic ;
         d_arr_3_31 : OUT std_logic ;
         d_arr_3_30 : OUT std_logic ;
         d_arr_3_29 : OUT std_logic ;
         d_arr_3_28 : OUT std_logic ;
         d_arr_3_27 : OUT std_logic ;
         d_arr_3_26 : OUT std_logic ;
         d_arr_3_25 : OUT std_logic ;
         d_arr_3_24 : OUT std_logic ;
         d_arr_3_23 : OUT std_logic ;
         d_arr_3_22 : OUT std_logic ;
         d_arr_3_21 : OUT std_logic ;
         d_arr_3_20 : OUT std_logic ;
         d_arr_3_19 : OUT std_logic ;
         d_arr_3_18 : OUT std_logic ;
         d_arr_3_17 : OUT std_logic ;
         d_arr_3_16 : OUT std_logic ;
         d_arr_3_15 : OUT std_logic ;
         d_arr_3_14 : OUT std_logic ;
         d_arr_3_13 : OUT std_logic ;
         d_arr_3_12 : OUT std_logic ;
         d_arr_3_11 : OUT std_logic ;
         d_arr_3_10 : OUT std_logic ;
         d_arr_3_9 : OUT std_logic ;
         d_arr_3_8 : OUT std_logic ;
         d_arr_3_7 : OUT std_logic ;
         d_arr_3_6 : OUT std_logic ;
         d_arr_3_5 : OUT std_logic ;
         d_arr_3_4 : OUT std_logic ;
         d_arr_3_3 : OUT std_logic ;
         d_arr_3_2 : OUT std_logic ;
         d_arr_3_1 : OUT std_logic ;
         d_arr_3_0 : OUT std_logic ;
         d_arr_4_31 : OUT std_logic ;
         d_arr_4_30 : OUT std_logic ;
         d_arr_4_29 : OUT std_logic ;
         d_arr_4_28 : OUT std_logic ;
         d_arr_4_27 : OUT std_logic ;
         d_arr_4_26 : OUT std_logic ;
         d_arr_4_25 : OUT std_logic ;
         d_arr_4_24 : OUT std_logic ;
         d_arr_4_23 : OUT std_logic ;
         d_arr_4_22 : OUT std_logic ;
         d_arr_4_21 : OUT std_logic ;
         d_arr_4_20 : OUT std_logic ;
         d_arr_4_19 : OUT std_logic ;
         d_arr_4_18 : OUT std_logic ;
         d_arr_4_17 : OUT std_logic ;
         d_arr_4_16 : OUT std_logic ;
         d_arr_4_15 : OUT std_logic ;
         d_arr_4_14 : OUT std_logic ;
         d_arr_4_13 : OUT std_logic ;
         d_arr_4_12 : OUT std_logic ;
         d_arr_4_11 : OUT std_logic ;
         d_arr_4_10 : OUT std_logic ;
         d_arr_4_9 : OUT std_logic ;
         d_arr_4_8 : OUT std_logic ;
         d_arr_4_7 : OUT std_logic ;
         d_arr_4_6 : OUT std_logic ;
         d_arr_4_5 : OUT std_logic ;
         d_arr_4_4 : OUT std_logic ;
         d_arr_4_3 : OUT std_logic ;
         d_arr_4_2 : OUT std_logic ;
         d_arr_4_1 : OUT std_logic ;
         d_arr_4_0 : OUT std_logic ;
         d_arr_5_31 : OUT std_logic ;
         d_arr_5_30 : OUT std_logic ;
         d_arr_5_29 : OUT std_logic ;
         d_arr_5_28 : OUT std_logic ;
         d_arr_5_27 : OUT std_logic ;
         d_arr_5_26 : OUT std_logic ;
         d_arr_5_25 : OUT std_logic ;
         d_arr_5_24 : OUT std_logic ;
         d_arr_5_23 : OUT std_logic ;
         d_arr_5_22 : OUT std_logic ;
         d_arr_5_21 : OUT std_logic ;
         d_arr_5_20 : OUT std_logic ;
         d_arr_5_19 : OUT std_logic ;
         d_arr_5_18 : OUT std_logic ;
         d_arr_5_17 : OUT std_logic ;
         d_arr_5_16 : OUT std_logic ;
         d_arr_5_15 : OUT std_logic ;
         d_arr_5_14 : OUT std_logic ;
         d_arr_5_13 : OUT std_logic ;
         d_arr_5_12 : OUT std_logic ;
         d_arr_5_11 : OUT std_logic ;
         d_arr_5_10 : OUT std_logic ;
         d_arr_5_9 : OUT std_logic ;
         d_arr_5_8 : OUT std_logic ;
         d_arr_5_7 : OUT std_logic ;
         d_arr_5_6 : OUT std_logic ;
         d_arr_5_5 : OUT std_logic ;
         d_arr_5_4 : OUT std_logic ;
         d_arr_5_3 : OUT std_logic ;
         d_arr_5_2 : OUT std_logic ;
         d_arr_5_1 : OUT std_logic ;
         d_arr_5_0 : OUT std_logic ;
         d_arr_6_31 : OUT std_logic ;
         d_arr_6_30 : OUT std_logic ;
         d_arr_6_29 : OUT std_logic ;
         d_arr_6_28 : OUT std_logic ;
         d_arr_6_27 : OUT std_logic ;
         d_arr_6_26 : OUT std_logic ;
         d_arr_6_25 : OUT std_logic ;
         d_arr_6_24 : OUT std_logic ;
         d_arr_6_23 : OUT std_logic ;
         d_arr_6_22 : OUT std_logic ;
         d_arr_6_21 : OUT std_logic ;
         d_arr_6_20 : OUT std_logic ;
         d_arr_6_19 : OUT std_logic ;
         d_arr_6_18 : OUT std_logic ;
         d_arr_6_17 : OUT std_logic ;
         d_arr_6_16 : OUT std_logic ;
         d_arr_6_15 : OUT std_logic ;
         d_arr_6_14 : OUT std_logic ;
         d_arr_6_13 : OUT std_logic ;
         d_arr_6_12 : OUT std_logic ;
         d_arr_6_11 : OUT std_logic ;
         d_arr_6_10 : OUT std_logic ;
         d_arr_6_9 : OUT std_logic ;
         d_arr_6_8 : OUT std_logic ;
         d_arr_6_7 : OUT std_logic ;
         d_arr_6_6 : OUT std_logic ;
         d_arr_6_5 : OUT std_logic ;
         d_arr_6_4 : OUT std_logic ;
         d_arr_6_3 : OUT std_logic ;
         d_arr_6_2 : OUT std_logic ;
         d_arr_6_1 : OUT std_logic ;
         d_arr_6_0 : OUT std_logic ;
         d_arr_7_31 : OUT std_logic ;
         d_arr_7_30 : OUT std_logic ;
         d_arr_7_29 : OUT std_logic ;
         d_arr_7_28 : OUT std_logic ;
         d_arr_7_27 : OUT std_logic ;
         d_arr_7_26 : OUT std_logic ;
         d_arr_7_25 : OUT std_logic ;
         d_arr_7_24 : OUT std_logic ;
         d_arr_7_23 : OUT std_logic ;
         d_arr_7_22 : OUT std_logic ;
         d_arr_7_21 : OUT std_logic ;
         d_arr_7_20 : OUT std_logic ;
         d_arr_7_19 : OUT std_logic ;
         d_arr_7_18 : OUT std_logic ;
         d_arr_7_17 : OUT std_logic ;
         d_arr_7_16 : OUT std_logic ;
         d_arr_7_15 : OUT std_logic ;
         d_arr_7_14 : OUT std_logic ;
         d_arr_7_13 : OUT std_logic ;
         d_arr_7_12 : OUT std_logic ;
         d_arr_7_11 : OUT std_logic ;
         d_arr_7_10 : OUT std_logic ;
         d_arr_7_9 : OUT std_logic ;
         d_arr_7_8 : OUT std_logic ;
         d_arr_7_7 : OUT std_logic ;
         d_arr_7_6 : OUT std_logic ;
         d_arr_7_5 : OUT std_logic ;
         d_arr_7_4 : OUT std_logic ;
         d_arr_7_3 : OUT std_logic ;
         d_arr_7_2 : OUT std_logic ;
         d_arr_7_1 : OUT std_logic ;
         d_arr_7_0 : OUT std_logic ;
         d_arr_8_31 : OUT std_logic ;
         d_arr_8_30 : OUT std_logic ;
         d_arr_8_29 : OUT std_logic ;
         d_arr_8_28 : OUT std_logic ;
         d_arr_8_27 : OUT std_logic ;
         d_arr_8_26 : OUT std_logic ;
         d_arr_8_25 : OUT std_logic ;
         d_arr_8_24 : OUT std_logic ;
         d_arr_8_23 : OUT std_logic ;
         d_arr_8_22 : OUT std_logic ;
         d_arr_8_21 : OUT std_logic ;
         d_arr_8_20 : OUT std_logic ;
         d_arr_8_19 : OUT std_logic ;
         d_arr_8_18 : OUT std_logic ;
         d_arr_8_17 : OUT std_logic ;
         d_arr_8_16 : OUT std_logic ;
         d_arr_8_15 : OUT std_logic ;
         d_arr_8_14 : OUT std_logic ;
         d_arr_8_13 : OUT std_logic ;
         d_arr_8_12 : OUT std_logic ;
         d_arr_8_11 : OUT std_logic ;
         d_arr_8_10 : OUT std_logic ;
         d_arr_8_9 : OUT std_logic ;
         d_arr_8_8 : OUT std_logic ;
         d_arr_8_7 : OUT std_logic ;
         d_arr_8_6 : OUT std_logic ;
         d_arr_8_5 : OUT std_logic ;
         d_arr_8_4 : OUT std_logic ;
         d_arr_8_3 : OUT std_logic ;
         d_arr_8_2 : OUT std_logic ;
         d_arr_8_1 : OUT std_logic ;
         d_arr_8_0 : OUT std_logic ;
         d_arr_9_31 : OUT std_logic ;
         d_arr_9_30 : OUT std_logic ;
         d_arr_9_29 : OUT std_logic ;
         d_arr_9_28 : OUT std_logic ;
         d_arr_9_27 : OUT std_logic ;
         d_arr_9_26 : OUT std_logic ;
         d_arr_9_25 : OUT std_logic ;
         d_arr_9_24 : OUT std_logic ;
         d_arr_9_23 : OUT std_logic ;
         d_arr_9_22 : OUT std_logic ;
         d_arr_9_21 : OUT std_logic ;
         d_arr_9_20 : OUT std_logic ;
         d_arr_9_19 : OUT std_logic ;
         d_arr_9_18 : OUT std_logic ;
         d_arr_9_17 : OUT std_logic ;
         d_arr_9_16 : OUT std_logic ;
         d_arr_9_15 : OUT std_logic ;
         d_arr_9_14 : OUT std_logic ;
         d_arr_9_13 : OUT std_logic ;
         d_arr_9_12 : OUT std_logic ;
         d_arr_9_11 : OUT std_logic ;
         d_arr_9_10 : OUT std_logic ;
         d_arr_9_9 : OUT std_logic ;
         d_arr_9_8 : OUT std_logic ;
         d_arr_9_7 : OUT std_logic ;
         d_arr_9_6 : OUT std_logic ;
         d_arr_9_5 : OUT std_logic ;
         d_arr_9_4 : OUT std_logic ;
         d_arr_9_3 : OUT std_logic ;
         d_arr_9_2 : OUT std_logic ;
         d_arr_9_1 : OUT std_logic ;
         d_arr_9_0 : OUT std_logic ;
         d_arr_10_31 : OUT std_logic ;
         d_arr_10_30 : OUT std_logic ;
         d_arr_10_29 : OUT std_logic ;
         d_arr_10_28 : OUT std_logic ;
         d_arr_10_27 : OUT std_logic ;
         d_arr_10_26 : OUT std_logic ;
         d_arr_10_25 : OUT std_logic ;
         d_arr_10_24 : OUT std_logic ;
         d_arr_10_23 : OUT std_logic ;
         d_arr_10_22 : OUT std_logic ;
         d_arr_10_21 : OUT std_logic ;
         d_arr_10_20 : OUT std_logic ;
         d_arr_10_19 : OUT std_logic ;
         d_arr_10_18 : OUT std_logic ;
         d_arr_10_17 : OUT std_logic ;
         d_arr_10_16 : OUT std_logic ;
         d_arr_10_15 : OUT std_logic ;
         d_arr_10_14 : OUT std_logic ;
         d_arr_10_13 : OUT std_logic ;
         d_arr_10_12 : OUT std_logic ;
         d_arr_10_11 : OUT std_logic ;
         d_arr_10_10 : OUT std_logic ;
         d_arr_10_9 : OUT std_logic ;
         d_arr_10_8 : OUT std_logic ;
         d_arr_10_7 : OUT std_logic ;
         d_arr_10_6 : OUT std_logic ;
         d_arr_10_5 : OUT std_logic ;
         d_arr_10_4 : OUT std_logic ;
         d_arr_10_3 : OUT std_logic ;
         d_arr_10_2 : OUT std_logic ;
         d_arr_10_1 : OUT std_logic ;
         d_arr_10_0 : OUT std_logic ;
         d_arr_11_31 : OUT std_logic ;
         d_arr_11_30 : OUT std_logic ;
         d_arr_11_29 : OUT std_logic ;
         d_arr_11_28 : OUT std_logic ;
         d_arr_11_27 : OUT std_logic ;
         d_arr_11_26 : OUT std_logic ;
         d_arr_11_25 : OUT std_logic ;
         d_arr_11_24 : OUT std_logic ;
         d_arr_11_23 : OUT std_logic ;
         d_arr_11_22 : OUT std_logic ;
         d_arr_11_21 : OUT std_logic ;
         d_arr_11_20 : OUT std_logic ;
         d_arr_11_19 : OUT std_logic ;
         d_arr_11_18 : OUT std_logic ;
         d_arr_11_17 : OUT std_logic ;
         d_arr_11_16 : OUT std_logic ;
         d_arr_11_15 : OUT std_logic ;
         d_arr_11_14 : OUT std_logic ;
         d_arr_11_13 : OUT std_logic ;
         d_arr_11_12 : OUT std_logic ;
         d_arr_11_11 : OUT std_logic ;
         d_arr_11_10 : OUT std_logic ;
         d_arr_11_9 : OUT std_logic ;
         d_arr_11_8 : OUT std_logic ;
         d_arr_11_7 : OUT std_logic ;
         d_arr_11_6 : OUT std_logic ;
         d_arr_11_5 : OUT std_logic ;
         d_arr_11_4 : OUT std_logic ;
         d_arr_11_3 : OUT std_logic ;
         d_arr_11_2 : OUT std_logic ;
         d_arr_11_1 : OUT std_logic ;
         d_arr_11_0 : OUT std_logic ;
         d_arr_12_31 : OUT std_logic ;
         d_arr_12_30 : OUT std_logic ;
         d_arr_12_29 : OUT std_logic ;
         d_arr_12_28 : OUT std_logic ;
         d_arr_12_27 : OUT std_logic ;
         d_arr_12_26 : OUT std_logic ;
         d_arr_12_25 : OUT std_logic ;
         d_arr_12_24 : OUT std_logic ;
         d_arr_12_23 : OUT std_logic ;
         d_arr_12_22 : OUT std_logic ;
         d_arr_12_21 : OUT std_logic ;
         d_arr_12_20 : OUT std_logic ;
         d_arr_12_19 : OUT std_logic ;
         d_arr_12_18 : OUT std_logic ;
         d_arr_12_17 : OUT std_logic ;
         d_arr_12_16 : OUT std_logic ;
         d_arr_12_15 : OUT std_logic ;
         d_arr_12_14 : OUT std_logic ;
         d_arr_12_13 : OUT std_logic ;
         d_arr_12_12 : OUT std_logic ;
         d_arr_12_11 : OUT std_logic ;
         d_arr_12_10 : OUT std_logic ;
         d_arr_12_9 : OUT std_logic ;
         d_arr_12_8 : OUT std_logic ;
         d_arr_12_7 : OUT std_logic ;
         d_arr_12_6 : OUT std_logic ;
         d_arr_12_5 : OUT std_logic ;
         d_arr_12_4 : OUT std_logic ;
         d_arr_12_3 : OUT std_logic ;
         d_arr_12_2 : OUT std_logic ;
         d_arr_12_1 : OUT std_logic ;
         d_arr_12_0 : OUT std_logic ;
         d_arr_13_31 : OUT std_logic ;
         d_arr_13_30 : OUT std_logic ;
         d_arr_13_29 : OUT std_logic ;
         d_arr_13_28 : OUT std_logic ;
         d_arr_13_27 : OUT std_logic ;
         d_arr_13_26 : OUT std_logic ;
         d_arr_13_25 : OUT std_logic ;
         d_arr_13_24 : OUT std_logic ;
         d_arr_13_23 : OUT std_logic ;
         d_arr_13_22 : OUT std_logic ;
         d_arr_13_21 : OUT std_logic ;
         d_arr_13_20 : OUT std_logic ;
         d_arr_13_19 : OUT std_logic ;
         d_arr_13_18 : OUT std_logic ;
         d_arr_13_17 : OUT std_logic ;
         d_arr_13_16 : OUT std_logic ;
         d_arr_13_15 : OUT std_logic ;
         d_arr_13_14 : OUT std_logic ;
         d_arr_13_13 : OUT std_logic ;
         d_arr_13_12 : OUT std_logic ;
         d_arr_13_11 : OUT std_logic ;
         d_arr_13_10 : OUT std_logic ;
         d_arr_13_9 : OUT std_logic ;
         d_arr_13_8 : OUT std_logic ;
         d_arr_13_7 : OUT std_logic ;
         d_arr_13_6 : OUT std_logic ;
         d_arr_13_5 : OUT std_logic ;
         d_arr_13_4 : OUT std_logic ;
         d_arr_13_3 : OUT std_logic ;
         d_arr_13_2 : OUT std_logic ;
         d_arr_13_1 : OUT std_logic ;
         d_arr_13_0 : OUT std_logic ;
         d_arr_14_31 : OUT std_logic ;
         d_arr_14_30 : OUT std_logic ;
         d_arr_14_29 : OUT std_logic ;
         d_arr_14_28 : OUT std_logic ;
         d_arr_14_27 : OUT std_logic ;
         d_arr_14_26 : OUT std_logic ;
         d_arr_14_25 : OUT std_logic ;
         d_arr_14_24 : OUT std_logic ;
         d_arr_14_23 : OUT std_logic ;
         d_arr_14_22 : OUT std_logic ;
         d_arr_14_21 : OUT std_logic ;
         d_arr_14_20 : OUT std_logic ;
         d_arr_14_19 : OUT std_logic ;
         d_arr_14_18 : OUT std_logic ;
         d_arr_14_17 : OUT std_logic ;
         d_arr_14_16 : OUT std_logic ;
         d_arr_14_15 : OUT std_logic ;
         d_arr_14_14 : OUT std_logic ;
         d_arr_14_13 : OUT std_logic ;
         d_arr_14_12 : OUT std_logic ;
         d_arr_14_11 : OUT std_logic ;
         d_arr_14_10 : OUT std_logic ;
         d_arr_14_9 : OUT std_logic ;
         d_arr_14_8 : OUT std_logic ;
         d_arr_14_7 : OUT std_logic ;
         d_arr_14_6 : OUT std_logic ;
         d_arr_14_5 : OUT std_logic ;
         d_arr_14_4 : OUT std_logic ;
         d_arr_14_3 : OUT std_logic ;
         d_arr_14_2 : OUT std_logic ;
         d_arr_14_1 : OUT std_logic ;
         d_arr_14_0 : OUT std_logic ;
         d_arr_15_31 : OUT std_logic ;
         d_arr_15_30 : OUT std_logic ;
         d_arr_15_29 : OUT std_logic ;
         d_arr_15_28 : OUT std_logic ;
         d_arr_15_27 : OUT std_logic ;
         d_arr_15_26 : OUT std_logic ;
         d_arr_15_25 : OUT std_logic ;
         d_arr_15_24 : OUT std_logic ;
         d_arr_15_23 : OUT std_logic ;
         d_arr_15_22 : OUT std_logic ;
         d_arr_15_21 : OUT std_logic ;
         d_arr_15_20 : OUT std_logic ;
         d_arr_15_19 : OUT std_logic ;
         d_arr_15_18 : OUT std_logic ;
         d_arr_15_17 : OUT std_logic ;
         d_arr_15_16 : OUT std_logic ;
         d_arr_15_15 : OUT std_logic ;
         d_arr_15_14 : OUT std_logic ;
         d_arr_15_13 : OUT std_logic ;
         d_arr_15_12 : OUT std_logic ;
         d_arr_15_11 : OUT std_logic ;
         d_arr_15_10 : OUT std_logic ;
         d_arr_15_9 : OUT std_logic ;
         d_arr_15_8 : OUT std_logic ;
         d_arr_15_7 : OUT std_logic ;
         d_arr_15_6 : OUT std_logic ;
         d_arr_15_5 : OUT std_logic ;
         d_arr_15_4 : OUT std_logic ;
         d_arr_15_3 : OUT std_logic ;
         d_arr_15_2 : OUT std_logic ;
         d_arr_15_1 : OUT std_logic ;
         d_arr_15_0 : OUT std_logic ;
         d_arr_16_31 : OUT std_logic ;
         d_arr_16_30 : OUT std_logic ;
         d_arr_16_29 : OUT std_logic ;
         d_arr_16_28 : OUT std_logic ;
         d_arr_16_27 : OUT std_logic ;
         d_arr_16_26 : OUT std_logic ;
         d_arr_16_25 : OUT std_logic ;
         d_arr_16_24 : OUT std_logic ;
         d_arr_16_23 : OUT std_logic ;
         d_arr_16_22 : OUT std_logic ;
         d_arr_16_21 : OUT std_logic ;
         d_arr_16_20 : OUT std_logic ;
         d_arr_16_19 : OUT std_logic ;
         d_arr_16_18 : OUT std_logic ;
         d_arr_16_17 : OUT std_logic ;
         d_arr_16_16 : OUT std_logic ;
         d_arr_16_15 : OUT std_logic ;
         d_arr_16_14 : OUT std_logic ;
         d_arr_16_13 : OUT std_logic ;
         d_arr_16_12 : OUT std_logic ;
         d_arr_16_11 : OUT std_logic ;
         d_arr_16_10 : OUT std_logic ;
         d_arr_16_9 : OUT std_logic ;
         d_arr_16_8 : OUT std_logic ;
         d_arr_16_7 : OUT std_logic ;
         d_arr_16_6 : OUT std_logic ;
         d_arr_16_5 : OUT std_logic ;
         d_arr_16_4 : OUT std_logic ;
         d_arr_16_3 : OUT std_logic ;
         d_arr_16_2 : OUT std_logic ;
         d_arr_16_1 : OUT std_logic ;
         d_arr_16_0 : OUT std_logic ;
         d_arr_17_31 : OUT std_logic ;
         d_arr_17_30 : OUT std_logic ;
         d_arr_17_29 : OUT std_logic ;
         d_arr_17_28 : OUT std_logic ;
         d_arr_17_27 : OUT std_logic ;
         d_arr_17_26 : OUT std_logic ;
         d_arr_17_25 : OUT std_logic ;
         d_arr_17_24 : OUT std_logic ;
         d_arr_17_23 : OUT std_logic ;
         d_arr_17_22 : OUT std_logic ;
         d_arr_17_21 : OUT std_logic ;
         d_arr_17_20 : OUT std_logic ;
         d_arr_17_19 : OUT std_logic ;
         d_arr_17_18 : OUT std_logic ;
         d_arr_17_17 : OUT std_logic ;
         d_arr_17_16 : OUT std_logic ;
         d_arr_17_15 : OUT std_logic ;
         d_arr_17_14 : OUT std_logic ;
         d_arr_17_13 : OUT std_logic ;
         d_arr_17_12 : OUT std_logic ;
         d_arr_17_11 : OUT std_logic ;
         d_arr_17_10 : OUT std_logic ;
         d_arr_17_9 : OUT std_logic ;
         d_arr_17_8 : OUT std_logic ;
         d_arr_17_7 : OUT std_logic ;
         d_arr_17_6 : OUT std_logic ;
         d_arr_17_5 : OUT std_logic ;
         d_arr_17_4 : OUT std_logic ;
         d_arr_17_3 : OUT std_logic ;
         d_arr_17_2 : OUT std_logic ;
         d_arr_17_1 : OUT std_logic ;
         d_arr_17_0 : OUT std_logic ;
         d_arr_18_31 : OUT std_logic ;
         d_arr_18_30 : OUT std_logic ;
         d_arr_18_29 : OUT std_logic ;
         d_arr_18_28 : OUT std_logic ;
         d_arr_18_27 : OUT std_logic ;
         d_arr_18_26 : OUT std_logic ;
         d_arr_18_25 : OUT std_logic ;
         d_arr_18_24 : OUT std_logic ;
         d_arr_18_23 : OUT std_logic ;
         d_arr_18_22 : OUT std_logic ;
         d_arr_18_21 : OUT std_logic ;
         d_arr_18_20 : OUT std_logic ;
         d_arr_18_19 : OUT std_logic ;
         d_arr_18_18 : OUT std_logic ;
         d_arr_18_17 : OUT std_logic ;
         d_arr_18_16 : OUT std_logic ;
         d_arr_18_15 : OUT std_logic ;
         d_arr_18_14 : OUT std_logic ;
         d_arr_18_13 : OUT std_logic ;
         d_arr_18_12 : OUT std_logic ;
         d_arr_18_11 : OUT std_logic ;
         d_arr_18_10 : OUT std_logic ;
         d_arr_18_9 : OUT std_logic ;
         d_arr_18_8 : OUT std_logic ;
         d_arr_18_7 : OUT std_logic ;
         d_arr_18_6 : OUT std_logic ;
         d_arr_18_5 : OUT std_logic ;
         d_arr_18_4 : OUT std_logic ;
         d_arr_18_3 : OUT std_logic ;
         d_arr_18_2 : OUT std_logic ;
         d_arr_18_1 : OUT std_logic ;
         d_arr_18_0 : OUT std_logic ;
         d_arr_19_31 : OUT std_logic ;
         d_arr_19_30 : OUT std_logic ;
         d_arr_19_29 : OUT std_logic ;
         d_arr_19_28 : OUT std_logic ;
         d_arr_19_27 : OUT std_logic ;
         d_arr_19_26 : OUT std_logic ;
         d_arr_19_25 : OUT std_logic ;
         d_arr_19_24 : OUT std_logic ;
         d_arr_19_23 : OUT std_logic ;
         d_arr_19_22 : OUT std_logic ;
         d_arr_19_21 : OUT std_logic ;
         d_arr_19_20 : OUT std_logic ;
         d_arr_19_19 : OUT std_logic ;
         d_arr_19_18 : OUT std_logic ;
         d_arr_19_17 : OUT std_logic ;
         d_arr_19_16 : OUT std_logic ;
         d_arr_19_15 : OUT std_logic ;
         d_arr_19_14 : OUT std_logic ;
         d_arr_19_13 : OUT std_logic ;
         d_arr_19_12 : OUT std_logic ;
         d_arr_19_11 : OUT std_logic ;
         d_arr_19_10 : OUT std_logic ;
         d_arr_19_9 : OUT std_logic ;
         d_arr_19_8 : OUT std_logic ;
         d_arr_19_7 : OUT std_logic ;
         d_arr_19_6 : OUT std_logic ;
         d_arr_19_5 : OUT std_logic ;
         d_arr_19_4 : OUT std_logic ;
         d_arr_19_3 : OUT std_logic ;
         d_arr_19_2 : OUT std_logic ;
         d_arr_19_1 : OUT std_logic ;
         d_arr_19_0 : OUT std_logic ;
         d_arr_20_31 : OUT std_logic ;
         d_arr_20_30 : OUT std_logic ;
         d_arr_20_29 : OUT std_logic ;
         d_arr_20_28 : OUT std_logic ;
         d_arr_20_27 : OUT std_logic ;
         d_arr_20_26 : OUT std_logic ;
         d_arr_20_25 : OUT std_logic ;
         d_arr_20_24 : OUT std_logic ;
         d_arr_20_23 : OUT std_logic ;
         d_arr_20_22 : OUT std_logic ;
         d_arr_20_21 : OUT std_logic ;
         d_arr_20_20 : OUT std_logic ;
         d_arr_20_19 : OUT std_logic ;
         d_arr_20_18 : OUT std_logic ;
         d_arr_20_17 : OUT std_logic ;
         d_arr_20_16 : OUT std_logic ;
         d_arr_20_15 : OUT std_logic ;
         d_arr_20_14 : OUT std_logic ;
         d_arr_20_13 : OUT std_logic ;
         d_arr_20_12 : OUT std_logic ;
         d_arr_20_11 : OUT std_logic ;
         d_arr_20_10 : OUT std_logic ;
         d_arr_20_9 : OUT std_logic ;
         d_arr_20_8 : OUT std_logic ;
         d_arr_20_7 : OUT std_logic ;
         d_arr_20_6 : OUT std_logic ;
         d_arr_20_5 : OUT std_logic ;
         d_arr_20_4 : OUT std_logic ;
         d_arr_20_3 : OUT std_logic ;
         d_arr_20_2 : OUT std_logic ;
         d_arr_20_1 : OUT std_logic ;
         d_arr_20_0 : OUT std_logic ;
         d_arr_21_31 : OUT std_logic ;
         d_arr_21_30 : OUT std_logic ;
         d_arr_21_29 : OUT std_logic ;
         d_arr_21_28 : OUT std_logic ;
         d_arr_21_27 : OUT std_logic ;
         d_arr_21_26 : OUT std_logic ;
         d_arr_21_25 : OUT std_logic ;
         d_arr_21_24 : OUT std_logic ;
         d_arr_21_23 : OUT std_logic ;
         d_arr_21_22 : OUT std_logic ;
         d_arr_21_21 : OUT std_logic ;
         d_arr_21_20 : OUT std_logic ;
         d_arr_21_19 : OUT std_logic ;
         d_arr_21_18 : OUT std_logic ;
         d_arr_21_17 : OUT std_logic ;
         d_arr_21_16 : OUT std_logic ;
         d_arr_21_15 : OUT std_logic ;
         d_arr_21_14 : OUT std_logic ;
         d_arr_21_13 : OUT std_logic ;
         d_arr_21_12 : OUT std_logic ;
         d_arr_21_11 : OUT std_logic ;
         d_arr_21_10 : OUT std_logic ;
         d_arr_21_9 : OUT std_logic ;
         d_arr_21_8 : OUT std_logic ;
         d_arr_21_7 : OUT std_logic ;
         d_arr_21_6 : OUT std_logic ;
         d_arr_21_5 : OUT std_logic ;
         d_arr_21_4 : OUT std_logic ;
         d_arr_21_3 : OUT std_logic ;
         d_arr_21_2 : OUT std_logic ;
         d_arr_21_1 : OUT std_logic ;
         d_arr_21_0 : OUT std_logic ;
         d_arr_22_31 : OUT std_logic ;
         d_arr_22_30 : OUT std_logic ;
         d_arr_22_29 : OUT std_logic ;
         d_arr_22_28 : OUT std_logic ;
         d_arr_22_27 : OUT std_logic ;
         d_arr_22_26 : OUT std_logic ;
         d_arr_22_25 : OUT std_logic ;
         d_arr_22_24 : OUT std_logic ;
         d_arr_22_23 : OUT std_logic ;
         d_arr_22_22 : OUT std_logic ;
         d_arr_22_21 : OUT std_logic ;
         d_arr_22_20 : OUT std_logic ;
         d_arr_22_19 : OUT std_logic ;
         d_arr_22_18 : OUT std_logic ;
         d_arr_22_17 : OUT std_logic ;
         d_arr_22_16 : OUT std_logic ;
         d_arr_22_15 : OUT std_logic ;
         d_arr_22_14 : OUT std_logic ;
         d_arr_22_13 : OUT std_logic ;
         d_arr_22_12 : OUT std_logic ;
         d_arr_22_11 : OUT std_logic ;
         d_arr_22_10 : OUT std_logic ;
         d_arr_22_9 : OUT std_logic ;
         d_arr_22_8 : OUT std_logic ;
         d_arr_22_7 : OUT std_logic ;
         d_arr_22_6 : OUT std_logic ;
         d_arr_22_5 : OUT std_logic ;
         d_arr_22_4 : OUT std_logic ;
         d_arr_22_3 : OUT std_logic ;
         d_arr_22_2 : OUT std_logic ;
         d_arr_22_1 : OUT std_logic ;
         d_arr_22_0 : OUT std_logic ;
         d_arr_23_31 : OUT std_logic ;
         d_arr_23_30 : OUT std_logic ;
         d_arr_23_29 : OUT std_logic ;
         d_arr_23_28 : OUT std_logic ;
         d_arr_23_27 : OUT std_logic ;
         d_arr_23_26 : OUT std_logic ;
         d_arr_23_25 : OUT std_logic ;
         d_arr_23_24 : OUT std_logic ;
         d_arr_23_23 : OUT std_logic ;
         d_arr_23_22 : OUT std_logic ;
         d_arr_23_21 : OUT std_logic ;
         d_arr_23_20 : OUT std_logic ;
         d_arr_23_19 : OUT std_logic ;
         d_arr_23_18 : OUT std_logic ;
         d_arr_23_17 : OUT std_logic ;
         d_arr_23_16 : OUT std_logic ;
         d_arr_23_15 : OUT std_logic ;
         d_arr_23_14 : OUT std_logic ;
         d_arr_23_13 : OUT std_logic ;
         d_arr_23_12 : OUT std_logic ;
         d_arr_23_11 : OUT std_logic ;
         d_arr_23_10 : OUT std_logic ;
         d_arr_23_9 : OUT std_logic ;
         d_arr_23_8 : OUT std_logic ;
         d_arr_23_7 : OUT std_logic ;
         d_arr_23_6 : OUT std_logic ;
         d_arr_23_5 : OUT std_logic ;
         d_arr_23_4 : OUT std_logic ;
         d_arr_23_3 : OUT std_logic ;
         d_arr_23_2 : OUT std_logic ;
         d_arr_23_1 : OUT std_logic ;
         d_arr_23_0 : OUT std_logic ;
         d_arr_24_31 : OUT std_logic ;
         d_arr_24_30 : OUT std_logic ;
         d_arr_24_29 : OUT std_logic ;
         d_arr_24_28 : OUT std_logic ;
         d_arr_24_27 : OUT std_logic ;
         d_arr_24_26 : OUT std_logic ;
         d_arr_24_25 : OUT std_logic ;
         d_arr_24_24 : OUT std_logic ;
         d_arr_24_23 : OUT std_logic ;
         d_arr_24_22 : OUT std_logic ;
         d_arr_24_21 : OUT std_logic ;
         d_arr_24_20 : OUT std_logic ;
         d_arr_24_19 : OUT std_logic ;
         d_arr_24_18 : OUT std_logic ;
         d_arr_24_17 : OUT std_logic ;
         d_arr_24_16 : OUT std_logic ;
         d_arr_24_15 : OUT std_logic ;
         d_arr_24_14 : OUT std_logic ;
         d_arr_24_13 : OUT std_logic ;
         d_arr_24_12 : OUT std_logic ;
         d_arr_24_11 : OUT std_logic ;
         d_arr_24_10 : OUT std_logic ;
         d_arr_24_9 : OUT std_logic ;
         d_arr_24_8 : OUT std_logic ;
         d_arr_24_7 : OUT std_logic ;
         d_arr_24_6 : OUT std_logic ;
         d_arr_24_5 : OUT std_logic ;
         d_arr_24_4 : OUT std_logic ;
         d_arr_24_3 : OUT std_logic ;
         d_arr_24_2 : OUT std_logic ;
         d_arr_24_1 : OUT std_logic ;
         d_arr_24_0 : OUT std_logic ;
         q_arr_0_31 : IN std_logic ;
         q_arr_0_30 : IN std_logic ;
         q_arr_0_29 : IN std_logic ;
         q_arr_0_28 : IN std_logic ;
         q_arr_0_27 : IN std_logic ;
         q_arr_0_26 : IN std_logic ;
         q_arr_0_25 : IN std_logic ;
         q_arr_0_24 : IN std_logic ;
         q_arr_0_23 : IN std_logic ;
         q_arr_0_22 : IN std_logic ;
         q_arr_0_21 : IN std_logic ;
         q_arr_0_20 : IN std_logic ;
         q_arr_0_19 : IN std_logic ;
         q_arr_0_18 : IN std_logic ;
         q_arr_0_17 : IN std_logic ;
         q_arr_0_16 : IN std_logic ;
         q_arr_0_15 : IN std_logic ;
         q_arr_0_14 : IN std_logic ;
         q_arr_0_13 : IN std_logic ;
         q_arr_0_12 : IN std_logic ;
         q_arr_0_11 : IN std_logic ;
         q_arr_0_10 : IN std_logic ;
         q_arr_0_9 : IN std_logic ;
         q_arr_0_8 : IN std_logic ;
         q_arr_0_7 : IN std_logic ;
         q_arr_0_6 : IN std_logic ;
         q_arr_0_5 : IN std_logic ;
         q_arr_0_4 : IN std_logic ;
         q_arr_0_3 : IN std_logic ;
         q_arr_0_2 : IN std_logic ;
         q_arr_0_1 : IN std_logic ;
         q_arr_0_0 : IN std_logic ;
         q_arr_1_31 : IN std_logic ;
         q_arr_1_30 : IN std_logic ;
         q_arr_1_29 : IN std_logic ;
         q_arr_1_28 : IN std_logic ;
         q_arr_1_27 : IN std_logic ;
         q_arr_1_26 : IN std_logic ;
         q_arr_1_25 : IN std_logic ;
         q_arr_1_24 : IN std_logic ;
         q_arr_1_23 : IN std_logic ;
         q_arr_1_22 : IN std_logic ;
         q_arr_1_21 : IN std_logic ;
         q_arr_1_20 : IN std_logic ;
         q_arr_1_19 : IN std_logic ;
         q_arr_1_18 : IN std_logic ;
         q_arr_1_17 : IN std_logic ;
         q_arr_1_16 : IN std_logic ;
         q_arr_1_15 : IN std_logic ;
         q_arr_1_14 : IN std_logic ;
         q_arr_1_13 : IN std_logic ;
         q_arr_1_12 : IN std_logic ;
         q_arr_1_11 : IN std_logic ;
         q_arr_1_10 : IN std_logic ;
         q_arr_1_9 : IN std_logic ;
         q_arr_1_8 : IN std_logic ;
         q_arr_1_7 : IN std_logic ;
         q_arr_1_6 : IN std_logic ;
         q_arr_1_5 : IN std_logic ;
         q_arr_1_4 : IN std_logic ;
         q_arr_1_3 : IN std_logic ;
         q_arr_1_2 : IN std_logic ;
         q_arr_1_1 : IN std_logic ;
         q_arr_1_0 : IN std_logic ;
         q_arr_2_31 : IN std_logic ;
         q_arr_2_30 : IN std_logic ;
         q_arr_2_29 : IN std_logic ;
         q_arr_2_28 : IN std_logic ;
         q_arr_2_27 : IN std_logic ;
         q_arr_2_26 : IN std_logic ;
         q_arr_2_25 : IN std_logic ;
         q_arr_2_24 : IN std_logic ;
         q_arr_2_23 : IN std_logic ;
         q_arr_2_22 : IN std_logic ;
         q_arr_2_21 : IN std_logic ;
         q_arr_2_20 : IN std_logic ;
         q_arr_2_19 : IN std_logic ;
         q_arr_2_18 : IN std_logic ;
         q_arr_2_17 : IN std_logic ;
         q_arr_2_16 : IN std_logic ;
         q_arr_2_15 : IN std_logic ;
         q_arr_2_14 : IN std_logic ;
         q_arr_2_13 : IN std_logic ;
         q_arr_2_12 : IN std_logic ;
         q_arr_2_11 : IN std_logic ;
         q_arr_2_10 : IN std_logic ;
         q_arr_2_9 : IN std_logic ;
         q_arr_2_8 : IN std_logic ;
         q_arr_2_7 : IN std_logic ;
         q_arr_2_6 : IN std_logic ;
         q_arr_2_5 : IN std_logic ;
         q_arr_2_4 : IN std_logic ;
         q_arr_2_3 : IN std_logic ;
         q_arr_2_2 : IN std_logic ;
         q_arr_2_1 : IN std_logic ;
         q_arr_2_0 : IN std_logic ;
         q_arr_3_31 : IN std_logic ;
         q_arr_3_30 : IN std_logic ;
         q_arr_3_29 : IN std_logic ;
         q_arr_3_28 : IN std_logic ;
         q_arr_3_27 : IN std_logic ;
         q_arr_3_26 : IN std_logic ;
         q_arr_3_25 : IN std_logic ;
         q_arr_3_24 : IN std_logic ;
         q_arr_3_23 : IN std_logic ;
         q_arr_3_22 : IN std_logic ;
         q_arr_3_21 : IN std_logic ;
         q_arr_3_20 : IN std_logic ;
         q_arr_3_19 : IN std_logic ;
         q_arr_3_18 : IN std_logic ;
         q_arr_3_17 : IN std_logic ;
         q_arr_3_16 : IN std_logic ;
         q_arr_3_15 : IN std_logic ;
         q_arr_3_14 : IN std_logic ;
         q_arr_3_13 : IN std_logic ;
         q_arr_3_12 : IN std_logic ;
         q_arr_3_11 : IN std_logic ;
         q_arr_3_10 : IN std_logic ;
         q_arr_3_9 : IN std_logic ;
         q_arr_3_8 : IN std_logic ;
         q_arr_3_7 : IN std_logic ;
         q_arr_3_6 : IN std_logic ;
         q_arr_3_5 : IN std_logic ;
         q_arr_3_4 : IN std_logic ;
         q_arr_3_3 : IN std_logic ;
         q_arr_3_2 : IN std_logic ;
         q_arr_3_1 : IN std_logic ;
         q_arr_3_0 : IN std_logic ;
         q_arr_4_31 : IN std_logic ;
         q_arr_4_30 : IN std_logic ;
         q_arr_4_29 : IN std_logic ;
         q_arr_4_28 : IN std_logic ;
         q_arr_4_27 : IN std_logic ;
         q_arr_4_26 : IN std_logic ;
         q_arr_4_25 : IN std_logic ;
         q_arr_4_24 : IN std_logic ;
         q_arr_4_23 : IN std_logic ;
         q_arr_4_22 : IN std_logic ;
         q_arr_4_21 : IN std_logic ;
         q_arr_4_20 : IN std_logic ;
         q_arr_4_19 : IN std_logic ;
         q_arr_4_18 : IN std_logic ;
         q_arr_4_17 : IN std_logic ;
         q_arr_4_16 : IN std_logic ;
         q_arr_4_15 : IN std_logic ;
         q_arr_4_14 : IN std_logic ;
         q_arr_4_13 : IN std_logic ;
         q_arr_4_12 : IN std_logic ;
         q_arr_4_11 : IN std_logic ;
         q_arr_4_10 : IN std_logic ;
         q_arr_4_9 : IN std_logic ;
         q_arr_4_8 : IN std_logic ;
         q_arr_4_7 : IN std_logic ;
         q_arr_4_6 : IN std_logic ;
         q_arr_4_5 : IN std_logic ;
         q_arr_4_4 : IN std_logic ;
         q_arr_4_3 : IN std_logic ;
         q_arr_4_2 : IN std_logic ;
         q_arr_4_1 : IN std_logic ;
         q_arr_4_0 : IN std_logic ;
         q_arr_5_31 : IN std_logic ;
         q_arr_5_30 : IN std_logic ;
         q_arr_5_29 : IN std_logic ;
         q_arr_5_28 : IN std_logic ;
         q_arr_5_27 : IN std_logic ;
         q_arr_5_26 : IN std_logic ;
         q_arr_5_25 : IN std_logic ;
         q_arr_5_24 : IN std_logic ;
         q_arr_5_23 : IN std_logic ;
         q_arr_5_22 : IN std_logic ;
         q_arr_5_21 : IN std_logic ;
         q_arr_5_20 : IN std_logic ;
         q_arr_5_19 : IN std_logic ;
         q_arr_5_18 : IN std_logic ;
         q_arr_5_17 : IN std_logic ;
         q_arr_5_16 : IN std_logic ;
         q_arr_5_15 : IN std_logic ;
         q_arr_5_14 : IN std_logic ;
         q_arr_5_13 : IN std_logic ;
         q_arr_5_12 : IN std_logic ;
         q_arr_5_11 : IN std_logic ;
         q_arr_5_10 : IN std_logic ;
         q_arr_5_9 : IN std_logic ;
         q_arr_5_8 : IN std_logic ;
         q_arr_5_7 : IN std_logic ;
         q_arr_5_6 : IN std_logic ;
         q_arr_5_5 : IN std_logic ;
         q_arr_5_4 : IN std_logic ;
         q_arr_5_3 : IN std_logic ;
         q_arr_5_2 : IN std_logic ;
         q_arr_5_1 : IN std_logic ;
         q_arr_5_0 : IN std_logic ;
         q_arr_6_31 : IN std_logic ;
         q_arr_6_30 : IN std_logic ;
         q_arr_6_29 : IN std_logic ;
         q_arr_6_28 : IN std_logic ;
         q_arr_6_27 : IN std_logic ;
         q_arr_6_26 : IN std_logic ;
         q_arr_6_25 : IN std_logic ;
         q_arr_6_24 : IN std_logic ;
         q_arr_6_23 : IN std_logic ;
         q_arr_6_22 : IN std_logic ;
         q_arr_6_21 : IN std_logic ;
         q_arr_6_20 : IN std_logic ;
         q_arr_6_19 : IN std_logic ;
         q_arr_6_18 : IN std_logic ;
         q_arr_6_17 : IN std_logic ;
         q_arr_6_16 : IN std_logic ;
         q_arr_6_15 : IN std_logic ;
         q_arr_6_14 : IN std_logic ;
         q_arr_6_13 : IN std_logic ;
         q_arr_6_12 : IN std_logic ;
         q_arr_6_11 : IN std_logic ;
         q_arr_6_10 : IN std_logic ;
         q_arr_6_9 : IN std_logic ;
         q_arr_6_8 : IN std_logic ;
         q_arr_6_7 : IN std_logic ;
         q_arr_6_6 : IN std_logic ;
         q_arr_6_5 : IN std_logic ;
         q_arr_6_4 : IN std_logic ;
         q_arr_6_3 : IN std_logic ;
         q_arr_6_2 : IN std_logic ;
         q_arr_6_1 : IN std_logic ;
         q_arr_6_0 : IN std_logic ;
         q_arr_7_31 : IN std_logic ;
         q_arr_7_30 : IN std_logic ;
         q_arr_7_29 : IN std_logic ;
         q_arr_7_28 : IN std_logic ;
         q_arr_7_27 : IN std_logic ;
         q_arr_7_26 : IN std_logic ;
         q_arr_7_25 : IN std_logic ;
         q_arr_7_24 : IN std_logic ;
         q_arr_7_23 : IN std_logic ;
         q_arr_7_22 : IN std_logic ;
         q_arr_7_21 : IN std_logic ;
         q_arr_7_20 : IN std_logic ;
         q_arr_7_19 : IN std_logic ;
         q_arr_7_18 : IN std_logic ;
         q_arr_7_17 : IN std_logic ;
         q_arr_7_16 : IN std_logic ;
         q_arr_7_15 : IN std_logic ;
         q_arr_7_14 : IN std_logic ;
         q_arr_7_13 : IN std_logic ;
         q_arr_7_12 : IN std_logic ;
         q_arr_7_11 : IN std_logic ;
         q_arr_7_10 : IN std_logic ;
         q_arr_7_9 : IN std_logic ;
         q_arr_7_8 : IN std_logic ;
         q_arr_7_7 : IN std_logic ;
         q_arr_7_6 : IN std_logic ;
         q_arr_7_5 : IN std_logic ;
         q_arr_7_4 : IN std_logic ;
         q_arr_7_3 : IN std_logic ;
         q_arr_7_2 : IN std_logic ;
         q_arr_7_1 : IN std_logic ;
         q_arr_7_0 : IN std_logic ;
         q_arr_8_31 : IN std_logic ;
         q_arr_8_30 : IN std_logic ;
         q_arr_8_29 : IN std_logic ;
         q_arr_8_28 : IN std_logic ;
         q_arr_8_27 : IN std_logic ;
         q_arr_8_26 : IN std_logic ;
         q_arr_8_25 : IN std_logic ;
         q_arr_8_24 : IN std_logic ;
         q_arr_8_23 : IN std_logic ;
         q_arr_8_22 : IN std_logic ;
         q_arr_8_21 : IN std_logic ;
         q_arr_8_20 : IN std_logic ;
         q_arr_8_19 : IN std_logic ;
         q_arr_8_18 : IN std_logic ;
         q_arr_8_17 : IN std_logic ;
         q_arr_8_16 : IN std_logic ;
         q_arr_8_15 : IN std_logic ;
         q_arr_8_14 : IN std_logic ;
         q_arr_8_13 : IN std_logic ;
         q_arr_8_12 : IN std_logic ;
         q_arr_8_11 : IN std_logic ;
         q_arr_8_10 : IN std_logic ;
         q_arr_8_9 : IN std_logic ;
         q_arr_8_8 : IN std_logic ;
         q_arr_8_7 : IN std_logic ;
         q_arr_8_6 : IN std_logic ;
         q_arr_8_5 : IN std_logic ;
         q_arr_8_4 : IN std_logic ;
         q_arr_8_3 : IN std_logic ;
         q_arr_8_2 : IN std_logic ;
         q_arr_8_1 : IN std_logic ;
         q_arr_8_0 : IN std_logic ;
         q_arr_9_31 : IN std_logic ;
         q_arr_9_30 : IN std_logic ;
         q_arr_9_29 : IN std_logic ;
         q_arr_9_28 : IN std_logic ;
         q_arr_9_27 : IN std_logic ;
         q_arr_9_26 : IN std_logic ;
         q_arr_9_25 : IN std_logic ;
         q_arr_9_24 : IN std_logic ;
         q_arr_9_23 : IN std_logic ;
         q_arr_9_22 : IN std_logic ;
         q_arr_9_21 : IN std_logic ;
         q_arr_9_20 : IN std_logic ;
         q_arr_9_19 : IN std_logic ;
         q_arr_9_18 : IN std_logic ;
         q_arr_9_17 : IN std_logic ;
         q_arr_9_16 : IN std_logic ;
         q_arr_9_15 : IN std_logic ;
         q_arr_9_14 : IN std_logic ;
         q_arr_9_13 : IN std_logic ;
         q_arr_9_12 : IN std_logic ;
         q_arr_9_11 : IN std_logic ;
         q_arr_9_10 : IN std_logic ;
         q_arr_9_9 : IN std_logic ;
         q_arr_9_8 : IN std_logic ;
         q_arr_9_7 : IN std_logic ;
         q_arr_9_6 : IN std_logic ;
         q_arr_9_5 : IN std_logic ;
         q_arr_9_4 : IN std_logic ;
         q_arr_9_3 : IN std_logic ;
         q_arr_9_2 : IN std_logic ;
         q_arr_9_1 : IN std_logic ;
         q_arr_9_0 : IN std_logic ;
         q_arr_10_31 : IN std_logic ;
         q_arr_10_30 : IN std_logic ;
         q_arr_10_29 : IN std_logic ;
         q_arr_10_28 : IN std_logic ;
         q_arr_10_27 : IN std_logic ;
         q_arr_10_26 : IN std_logic ;
         q_arr_10_25 : IN std_logic ;
         q_arr_10_24 : IN std_logic ;
         q_arr_10_23 : IN std_logic ;
         q_arr_10_22 : IN std_logic ;
         q_arr_10_21 : IN std_logic ;
         q_arr_10_20 : IN std_logic ;
         q_arr_10_19 : IN std_logic ;
         q_arr_10_18 : IN std_logic ;
         q_arr_10_17 : IN std_logic ;
         q_arr_10_16 : IN std_logic ;
         q_arr_10_15 : IN std_logic ;
         q_arr_10_14 : IN std_logic ;
         q_arr_10_13 : IN std_logic ;
         q_arr_10_12 : IN std_logic ;
         q_arr_10_11 : IN std_logic ;
         q_arr_10_10 : IN std_logic ;
         q_arr_10_9 : IN std_logic ;
         q_arr_10_8 : IN std_logic ;
         q_arr_10_7 : IN std_logic ;
         q_arr_10_6 : IN std_logic ;
         q_arr_10_5 : IN std_logic ;
         q_arr_10_4 : IN std_logic ;
         q_arr_10_3 : IN std_logic ;
         q_arr_10_2 : IN std_logic ;
         q_arr_10_1 : IN std_logic ;
         q_arr_10_0 : IN std_logic ;
         q_arr_11_31 : IN std_logic ;
         q_arr_11_30 : IN std_logic ;
         q_arr_11_29 : IN std_logic ;
         q_arr_11_28 : IN std_logic ;
         q_arr_11_27 : IN std_logic ;
         q_arr_11_26 : IN std_logic ;
         q_arr_11_25 : IN std_logic ;
         q_arr_11_24 : IN std_logic ;
         q_arr_11_23 : IN std_logic ;
         q_arr_11_22 : IN std_logic ;
         q_arr_11_21 : IN std_logic ;
         q_arr_11_20 : IN std_logic ;
         q_arr_11_19 : IN std_logic ;
         q_arr_11_18 : IN std_logic ;
         q_arr_11_17 : IN std_logic ;
         q_arr_11_16 : IN std_logic ;
         q_arr_11_15 : IN std_logic ;
         q_arr_11_14 : IN std_logic ;
         q_arr_11_13 : IN std_logic ;
         q_arr_11_12 : IN std_logic ;
         q_arr_11_11 : IN std_logic ;
         q_arr_11_10 : IN std_logic ;
         q_arr_11_9 : IN std_logic ;
         q_arr_11_8 : IN std_logic ;
         q_arr_11_7 : IN std_logic ;
         q_arr_11_6 : IN std_logic ;
         q_arr_11_5 : IN std_logic ;
         q_arr_11_4 : IN std_logic ;
         q_arr_11_3 : IN std_logic ;
         q_arr_11_2 : IN std_logic ;
         q_arr_11_1 : IN std_logic ;
         q_arr_11_0 : IN std_logic ;
         q_arr_12_31 : IN std_logic ;
         q_arr_12_30 : IN std_logic ;
         q_arr_12_29 : IN std_logic ;
         q_arr_12_28 : IN std_logic ;
         q_arr_12_27 : IN std_logic ;
         q_arr_12_26 : IN std_logic ;
         q_arr_12_25 : IN std_logic ;
         q_arr_12_24 : IN std_logic ;
         q_arr_12_23 : IN std_logic ;
         q_arr_12_22 : IN std_logic ;
         q_arr_12_21 : IN std_logic ;
         q_arr_12_20 : IN std_logic ;
         q_arr_12_19 : IN std_logic ;
         q_arr_12_18 : IN std_logic ;
         q_arr_12_17 : IN std_logic ;
         q_arr_12_16 : IN std_logic ;
         q_arr_12_15 : IN std_logic ;
         q_arr_12_14 : IN std_logic ;
         q_arr_12_13 : IN std_logic ;
         q_arr_12_12 : IN std_logic ;
         q_arr_12_11 : IN std_logic ;
         q_arr_12_10 : IN std_logic ;
         q_arr_12_9 : IN std_logic ;
         q_arr_12_8 : IN std_logic ;
         q_arr_12_7 : IN std_logic ;
         q_arr_12_6 : IN std_logic ;
         q_arr_12_5 : IN std_logic ;
         q_arr_12_4 : IN std_logic ;
         q_arr_12_3 : IN std_logic ;
         q_arr_12_2 : IN std_logic ;
         q_arr_12_1 : IN std_logic ;
         q_arr_12_0 : IN std_logic ;
         q_arr_13_31 : IN std_logic ;
         q_arr_13_30 : IN std_logic ;
         q_arr_13_29 : IN std_logic ;
         q_arr_13_28 : IN std_logic ;
         q_arr_13_27 : IN std_logic ;
         q_arr_13_26 : IN std_logic ;
         q_arr_13_25 : IN std_logic ;
         q_arr_13_24 : IN std_logic ;
         q_arr_13_23 : IN std_logic ;
         q_arr_13_22 : IN std_logic ;
         q_arr_13_21 : IN std_logic ;
         q_arr_13_20 : IN std_logic ;
         q_arr_13_19 : IN std_logic ;
         q_arr_13_18 : IN std_logic ;
         q_arr_13_17 : IN std_logic ;
         q_arr_13_16 : IN std_logic ;
         q_arr_13_15 : IN std_logic ;
         q_arr_13_14 : IN std_logic ;
         q_arr_13_13 : IN std_logic ;
         q_arr_13_12 : IN std_logic ;
         q_arr_13_11 : IN std_logic ;
         q_arr_13_10 : IN std_logic ;
         q_arr_13_9 : IN std_logic ;
         q_arr_13_8 : IN std_logic ;
         q_arr_13_7 : IN std_logic ;
         q_arr_13_6 : IN std_logic ;
         q_arr_13_5 : IN std_logic ;
         q_arr_13_4 : IN std_logic ;
         q_arr_13_3 : IN std_logic ;
         q_arr_13_2 : IN std_logic ;
         q_arr_13_1 : IN std_logic ;
         q_arr_13_0 : IN std_logic ;
         q_arr_14_31 : IN std_logic ;
         q_arr_14_30 : IN std_logic ;
         q_arr_14_29 : IN std_logic ;
         q_arr_14_28 : IN std_logic ;
         q_arr_14_27 : IN std_logic ;
         q_arr_14_26 : IN std_logic ;
         q_arr_14_25 : IN std_logic ;
         q_arr_14_24 : IN std_logic ;
         q_arr_14_23 : IN std_logic ;
         q_arr_14_22 : IN std_logic ;
         q_arr_14_21 : IN std_logic ;
         q_arr_14_20 : IN std_logic ;
         q_arr_14_19 : IN std_logic ;
         q_arr_14_18 : IN std_logic ;
         q_arr_14_17 : IN std_logic ;
         q_arr_14_16 : IN std_logic ;
         q_arr_14_15 : IN std_logic ;
         q_arr_14_14 : IN std_logic ;
         q_arr_14_13 : IN std_logic ;
         q_arr_14_12 : IN std_logic ;
         q_arr_14_11 : IN std_logic ;
         q_arr_14_10 : IN std_logic ;
         q_arr_14_9 : IN std_logic ;
         q_arr_14_8 : IN std_logic ;
         q_arr_14_7 : IN std_logic ;
         q_arr_14_6 : IN std_logic ;
         q_arr_14_5 : IN std_logic ;
         q_arr_14_4 : IN std_logic ;
         q_arr_14_3 : IN std_logic ;
         q_arr_14_2 : IN std_logic ;
         q_arr_14_1 : IN std_logic ;
         q_arr_14_0 : IN std_logic ;
         q_arr_15_31 : IN std_logic ;
         q_arr_15_30 : IN std_logic ;
         q_arr_15_29 : IN std_logic ;
         q_arr_15_28 : IN std_logic ;
         q_arr_15_27 : IN std_logic ;
         q_arr_15_26 : IN std_logic ;
         q_arr_15_25 : IN std_logic ;
         q_arr_15_24 : IN std_logic ;
         q_arr_15_23 : IN std_logic ;
         q_arr_15_22 : IN std_logic ;
         q_arr_15_21 : IN std_logic ;
         q_arr_15_20 : IN std_logic ;
         q_arr_15_19 : IN std_logic ;
         q_arr_15_18 : IN std_logic ;
         q_arr_15_17 : IN std_logic ;
         q_arr_15_16 : IN std_logic ;
         q_arr_15_15 : IN std_logic ;
         q_arr_15_14 : IN std_logic ;
         q_arr_15_13 : IN std_logic ;
         q_arr_15_12 : IN std_logic ;
         q_arr_15_11 : IN std_logic ;
         q_arr_15_10 : IN std_logic ;
         q_arr_15_9 : IN std_logic ;
         q_arr_15_8 : IN std_logic ;
         q_arr_15_7 : IN std_logic ;
         q_arr_15_6 : IN std_logic ;
         q_arr_15_5 : IN std_logic ;
         q_arr_15_4 : IN std_logic ;
         q_arr_15_3 : IN std_logic ;
         q_arr_15_2 : IN std_logic ;
         q_arr_15_1 : IN std_logic ;
         q_arr_15_0 : IN std_logic ;
         q_arr_16_31 : IN std_logic ;
         q_arr_16_30 : IN std_logic ;
         q_arr_16_29 : IN std_logic ;
         q_arr_16_28 : IN std_logic ;
         q_arr_16_27 : IN std_logic ;
         q_arr_16_26 : IN std_logic ;
         q_arr_16_25 : IN std_logic ;
         q_arr_16_24 : IN std_logic ;
         q_arr_16_23 : IN std_logic ;
         q_arr_16_22 : IN std_logic ;
         q_arr_16_21 : IN std_logic ;
         q_arr_16_20 : IN std_logic ;
         q_arr_16_19 : IN std_logic ;
         q_arr_16_18 : IN std_logic ;
         q_arr_16_17 : IN std_logic ;
         q_arr_16_16 : IN std_logic ;
         q_arr_16_15 : IN std_logic ;
         q_arr_16_14 : IN std_logic ;
         q_arr_16_13 : IN std_logic ;
         q_arr_16_12 : IN std_logic ;
         q_arr_16_11 : IN std_logic ;
         q_arr_16_10 : IN std_logic ;
         q_arr_16_9 : IN std_logic ;
         q_arr_16_8 : IN std_logic ;
         q_arr_16_7 : IN std_logic ;
         q_arr_16_6 : IN std_logic ;
         q_arr_16_5 : IN std_logic ;
         q_arr_16_4 : IN std_logic ;
         q_arr_16_3 : IN std_logic ;
         q_arr_16_2 : IN std_logic ;
         q_arr_16_1 : IN std_logic ;
         q_arr_16_0 : IN std_logic ;
         q_arr_17_31 : IN std_logic ;
         q_arr_17_30 : IN std_logic ;
         q_arr_17_29 : IN std_logic ;
         q_arr_17_28 : IN std_logic ;
         q_arr_17_27 : IN std_logic ;
         q_arr_17_26 : IN std_logic ;
         q_arr_17_25 : IN std_logic ;
         q_arr_17_24 : IN std_logic ;
         q_arr_17_23 : IN std_logic ;
         q_arr_17_22 : IN std_logic ;
         q_arr_17_21 : IN std_logic ;
         q_arr_17_20 : IN std_logic ;
         q_arr_17_19 : IN std_logic ;
         q_arr_17_18 : IN std_logic ;
         q_arr_17_17 : IN std_logic ;
         q_arr_17_16 : IN std_logic ;
         q_arr_17_15 : IN std_logic ;
         q_arr_17_14 : IN std_logic ;
         q_arr_17_13 : IN std_logic ;
         q_arr_17_12 : IN std_logic ;
         q_arr_17_11 : IN std_logic ;
         q_arr_17_10 : IN std_logic ;
         q_arr_17_9 : IN std_logic ;
         q_arr_17_8 : IN std_logic ;
         q_arr_17_7 : IN std_logic ;
         q_arr_17_6 : IN std_logic ;
         q_arr_17_5 : IN std_logic ;
         q_arr_17_4 : IN std_logic ;
         q_arr_17_3 : IN std_logic ;
         q_arr_17_2 : IN std_logic ;
         q_arr_17_1 : IN std_logic ;
         q_arr_17_0 : IN std_logic ;
         q_arr_18_31 : IN std_logic ;
         q_arr_18_30 : IN std_logic ;
         q_arr_18_29 : IN std_logic ;
         q_arr_18_28 : IN std_logic ;
         q_arr_18_27 : IN std_logic ;
         q_arr_18_26 : IN std_logic ;
         q_arr_18_25 : IN std_logic ;
         q_arr_18_24 : IN std_logic ;
         q_arr_18_23 : IN std_logic ;
         q_arr_18_22 : IN std_logic ;
         q_arr_18_21 : IN std_logic ;
         q_arr_18_20 : IN std_logic ;
         q_arr_18_19 : IN std_logic ;
         q_arr_18_18 : IN std_logic ;
         q_arr_18_17 : IN std_logic ;
         q_arr_18_16 : IN std_logic ;
         q_arr_18_15 : IN std_logic ;
         q_arr_18_14 : IN std_logic ;
         q_arr_18_13 : IN std_logic ;
         q_arr_18_12 : IN std_logic ;
         q_arr_18_11 : IN std_logic ;
         q_arr_18_10 : IN std_logic ;
         q_arr_18_9 : IN std_logic ;
         q_arr_18_8 : IN std_logic ;
         q_arr_18_7 : IN std_logic ;
         q_arr_18_6 : IN std_logic ;
         q_arr_18_5 : IN std_logic ;
         q_arr_18_4 : IN std_logic ;
         q_arr_18_3 : IN std_logic ;
         q_arr_18_2 : IN std_logic ;
         q_arr_18_1 : IN std_logic ;
         q_arr_18_0 : IN std_logic ;
         q_arr_19_31 : IN std_logic ;
         q_arr_19_30 : IN std_logic ;
         q_arr_19_29 : IN std_logic ;
         q_arr_19_28 : IN std_logic ;
         q_arr_19_27 : IN std_logic ;
         q_arr_19_26 : IN std_logic ;
         q_arr_19_25 : IN std_logic ;
         q_arr_19_24 : IN std_logic ;
         q_arr_19_23 : IN std_logic ;
         q_arr_19_22 : IN std_logic ;
         q_arr_19_21 : IN std_logic ;
         q_arr_19_20 : IN std_logic ;
         q_arr_19_19 : IN std_logic ;
         q_arr_19_18 : IN std_logic ;
         q_arr_19_17 : IN std_logic ;
         q_arr_19_16 : IN std_logic ;
         q_arr_19_15 : IN std_logic ;
         q_arr_19_14 : IN std_logic ;
         q_arr_19_13 : IN std_logic ;
         q_arr_19_12 : IN std_logic ;
         q_arr_19_11 : IN std_logic ;
         q_arr_19_10 : IN std_logic ;
         q_arr_19_9 : IN std_logic ;
         q_arr_19_8 : IN std_logic ;
         q_arr_19_7 : IN std_logic ;
         q_arr_19_6 : IN std_logic ;
         q_arr_19_5 : IN std_logic ;
         q_arr_19_4 : IN std_logic ;
         q_arr_19_3 : IN std_logic ;
         q_arr_19_2 : IN std_logic ;
         q_arr_19_1 : IN std_logic ;
         q_arr_19_0 : IN std_logic ;
         q_arr_20_31 : IN std_logic ;
         q_arr_20_30 : IN std_logic ;
         q_arr_20_29 : IN std_logic ;
         q_arr_20_28 : IN std_logic ;
         q_arr_20_27 : IN std_logic ;
         q_arr_20_26 : IN std_logic ;
         q_arr_20_25 : IN std_logic ;
         q_arr_20_24 : IN std_logic ;
         q_arr_20_23 : IN std_logic ;
         q_arr_20_22 : IN std_logic ;
         q_arr_20_21 : IN std_logic ;
         q_arr_20_20 : IN std_logic ;
         q_arr_20_19 : IN std_logic ;
         q_arr_20_18 : IN std_logic ;
         q_arr_20_17 : IN std_logic ;
         q_arr_20_16 : IN std_logic ;
         q_arr_20_15 : IN std_logic ;
         q_arr_20_14 : IN std_logic ;
         q_arr_20_13 : IN std_logic ;
         q_arr_20_12 : IN std_logic ;
         q_arr_20_11 : IN std_logic ;
         q_arr_20_10 : IN std_logic ;
         q_arr_20_9 : IN std_logic ;
         q_arr_20_8 : IN std_logic ;
         q_arr_20_7 : IN std_logic ;
         q_arr_20_6 : IN std_logic ;
         q_arr_20_5 : IN std_logic ;
         q_arr_20_4 : IN std_logic ;
         q_arr_20_3 : IN std_logic ;
         q_arr_20_2 : IN std_logic ;
         q_arr_20_1 : IN std_logic ;
         q_arr_20_0 : IN std_logic ;
         q_arr_21_31 : IN std_logic ;
         q_arr_21_30 : IN std_logic ;
         q_arr_21_29 : IN std_logic ;
         q_arr_21_28 : IN std_logic ;
         q_arr_21_27 : IN std_logic ;
         q_arr_21_26 : IN std_logic ;
         q_arr_21_25 : IN std_logic ;
         q_arr_21_24 : IN std_logic ;
         q_arr_21_23 : IN std_logic ;
         q_arr_21_22 : IN std_logic ;
         q_arr_21_21 : IN std_logic ;
         q_arr_21_20 : IN std_logic ;
         q_arr_21_19 : IN std_logic ;
         q_arr_21_18 : IN std_logic ;
         q_arr_21_17 : IN std_logic ;
         q_arr_21_16 : IN std_logic ;
         q_arr_21_15 : IN std_logic ;
         q_arr_21_14 : IN std_logic ;
         q_arr_21_13 : IN std_logic ;
         q_arr_21_12 : IN std_logic ;
         q_arr_21_11 : IN std_logic ;
         q_arr_21_10 : IN std_logic ;
         q_arr_21_9 : IN std_logic ;
         q_arr_21_8 : IN std_logic ;
         q_arr_21_7 : IN std_logic ;
         q_arr_21_6 : IN std_logic ;
         q_arr_21_5 : IN std_logic ;
         q_arr_21_4 : IN std_logic ;
         q_arr_21_3 : IN std_logic ;
         q_arr_21_2 : IN std_logic ;
         q_arr_21_1 : IN std_logic ;
         q_arr_21_0 : IN std_logic ;
         q_arr_22_31 : IN std_logic ;
         q_arr_22_30 : IN std_logic ;
         q_arr_22_29 : IN std_logic ;
         q_arr_22_28 : IN std_logic ;
         q_arr_22_27 : IN std_logic ;
         q_arr_22_26 : IN std_logic ;
         q_arr_22_25 : IN std_logic ;
         q_arr_22_24 : IN std_logic ;
         q_arr_22_23 : IN std_logic ;
         q_arr_22_22 : IN std_logic ;
         q_arr_22_21 : IN std_logic ;
         q_arr_22_20 : IN std_logic ;
         q_arr_22_19 : IN std_logic ;
         q_arr_22_18 : IN std_logic ;
         q_arr_22_17 : IN std_logic ;
         q_arr_22_16 : IN std_logic ;
         q_arr_22_15 : IN std_logic ;
         q_arr_22_14 : IN std_logic ;
         q_arr_22_13 : IN std_logic ;
         q_arr_22_12 : IN std_logic ;
         q_arr_22_11 : IN std_logic ;
         q_arr_22_10 : IN std_logic ;
         q_arr_22_9 : IN std_logic ;
         q_arr_22_8 : IN std_logic ;
         q_arr_22_7 : IN std_logic ;
         q_arr_22_6 : IN std_logic ;
         q_arr_22_5 : IN std_logic ;
         q_arr_22_4 : IN std_logic ;
         q_arr_22_3 : IN std_logic ;
         q_arr_22_2 : IN std_logic ;
         q_arr_22_1 : IN std_logic ;
         q_arr_22_0 : IN std_logic ;
         q_arr_23_31 : IN std_logic ;
         q_arr_23_30 : IN std_logic ;
         q_arr_23_29 : IN std_logic ;
         q_arr_23_28 : IN std_logic ;
         q_arr_23_27 : IN std_logic ;
         q_arr_23_26 : IN std_logic ;
         q_arr_23_25 : IN std_logic ;
         q_arr_23_24 : IN std_logic ;
         q_arr_23_23 : IN std_logic ;
         q_arr_23_22 : IN std_logic ;
         q_arr_23_21 : IN std_logic ;
         q_arr_23_20 : IN std_logic ;
         q_arr_23_19 : IN std_logic ;
         q_arr_23_18 : IN std_logic ;
         q_arr_23_17 : IN std_logic ;
         q_arr_23_16 : IN std_logic ;
         q_arr_23_15 : IN std_logic ;
         q_arr_23_14 : IN std_logic ;
         q_arr_23_13 : IN std_logic ;
         q_arr_23_12 : IN std_logic ;
         q_arr_23_11 : IN std_logic ;
         q_arr_23_10 : IN std_logic ;
         q_arr_23_9 : IN std_logic ;
         q_arr_23_8 : IN std_logic ;
         q_arr_23_7 : IN std_logic ;
         q_arr_23_6 : IN std_logic ;
         q_arr_23_5 : IN std_logic ;
         q_arr_23_4 : IN std_logic ;
         q_arr_23_3 : IN std_logic ;
         q_arr_23_2 : IN std_logic ;
         q_arr_23_1 : IN std_logic ;
         q_arr_23_0 : IN std_logic ;
         q_arr_24_31 : IN std_logic ;
         q_arr_24_30 : IN std_logic ;
         q_arr_24_29 : IN std_logic ;
         q_arr_24_28 : IN std_logic ;
         q_arr_24_27 : IN std_logic ;
         q_arr_24_26 : IN std_logic ;
         q_arr_24_25 : IN std_logic ;
         q_arr_24_24 : IN std_logic ;
         q_arr_24_23 : IN std_logic ;
         q_arr_24_22 : IN std_logic ;
         q_arr_24_21 : IN std_logic ;
         q_arr_24_20 : IN std_logic ;
         q_arr_24_19 : IN std_logic ;
         q_arr_24_18 : IN std_logic ;
         q_arr_24_17 : IN std_logic ;
         q_arr_24_16 : IN std_logic ;
         q_arr_24_15 : IN std_logic ;
         q_arr_24_14 : IN std_logic ;
         q_arr_24_13 : IN std_logic ;
         q_arr_24_12 : IN std_logic ;
         q_arr_24_11 : IN std_logic ;
         q_arr_24_10 : IN std_logic ;
         q_arr_24_9 : IN std_logic ;
         q_arr_24_8 : IN std_logic ;
         q_arr_24_7 : IN std_logic ;
         q_arr_24_6 : IN std_logic ;
         q_arr_24_5 : IN std_logic ;
         q_arr_24_4 : IN std_logic ;
         q_arr_24_3 : IN std_logic ;
         q_arr_24_2 : IN std_logic ;
         q_arr_24_1 : IN std_logic ;
         q_arr_24_0 : IN std_logic ;
         output1_init : IN std_logic_vector (15 DOWNTO 0) ;
         output2_init : IN std_logic_vector (15 DOWNTO 0) ;
         filter_size : IN std_logic ;
         operation : IN std_logic ;
         compute_relu : IN std_logic ;
         clk : IN std_logic ;
         en : IN std_logic ;
         reset : IN std_logic ;
         buffer_ready : OUT std_logic ;
         semi_ready : OUT std_logic ;
         ready : OUT std_logic) ;
   end component ;
   component Queue_5_unfolded0
      port (
         d : IN std_logic_vector (15 DOWNTO 0) ;
         q_0_15 : OUT std_logic ;
         q_0_14 : OUT std_logic ;
         q_0_13 : OUT std_logic ;
         q_0_12 : OUT std_logic ;
         q_0_11 : OUT std_logic ;
         q_0_10 : OUT std_logic ;
         q_0_9 : OUT std_logic ;
         q_0_8 : OUT std_logic ;
         q_0_7 : OUT std_logic ;
         q_0_6 : OUT std_logic ;
         q_0_5 : OUT std_logic ;
         q_0_4 : OUT std_logic ;
         q_0_3 : OUT std_logic ;
         q_0_2 : OUT std_logic ;
         q_0_1 : OUT std_logic ;
         q_0_0 : OUT std_logic ;
         q_1_15 : OUT std_logic ;
         q_1_14 : OUT std_logic ;
         q_1_13 : OUT std_logic ;
         q_1_12 : OUT std_logic ;
         q_1_11 : OUT std_logic ;
         q_1_10 : OUT std_logic ;
         q_1_9 : OUT std_logic ;
         q_1_8 : OUT std_logic ;
         q_1_7 : OUT std_logic ;
         q_1_6 : OUT std_logic ;
         q_1_5 : OUT std_logic ;
         q_1_4 : OUT std_logic ;
         q_1_3 : OUT std_logic ;
         q_1_2 : OUT std_logic ;
         q_1_1 : OUT std_logic ;
         q_1_0 : OUT std_logic ;
         q_2_15 : OUT std_logic ;
         q_2_14 : OUT std_logic ;
         q_2_13 : OUT std_logic ;
         q_2_12 : OUT std_logic ;
         q_2_11 : OUT std_logic ;
         q_2_10 : OUT std_logic ;
         q_2_9 : OUT std_logic ;
         q_2_8 : OUT std_logic ;
         q_2_7 : OUT std_logic ;
         q_2_6 : OUT std_logic ;
         q_2_5 : OUT std_logic ;
         q_2_4 : OUT std_logic ;
         q_2_3 : OUT std_logic ;
         q_2_2 : OUT std_logic ;
         q_2_1 : OUT std_logic ;
         q_2_0 : OUT std_logic ;
         q_3_15 : OUT std_logic ;
         q_3_14 : OUT std_logic ;
         q_3_13 : OUT std_logic ;
         q_3_12 : OUT std_logic ;
         q_3_11 : OUT std_logic ;
         q_3_10 : OUT std_logic ;
         q_3_9 : OUT std_logic ;
         q_3_8 : OUT std_logic ;
         q_3_7 : OUT std_logic ;
         q_3_6 : OUT std_logic ;
         q_3_5 : OUT std_logic ;
         q_3_4 : OUT std_logic ;
         q_3_3 : OUT std_logic ;
         q_3_2 : OUT std_logic ;
         q_3_1 : OUT std_logic ;
         q_3_0 : OUT std_logic ;
         q_4_15 : OUT std_logic ;
         q_4_14 : OUT std_logic ;
         q_4_13 : OUT std_logic ;
         q_4_12 : OUT std_logic ;
         q_4_11 : OUT std_logic ;
         q_4_10 : OUT std_logic ;
         q_4_9 : OUT std_logic ;
         q_4_8 : OUT std_logic ;
         q_4_7 : OUT std_logic ;
         q_4_6 : OUT std_logic ;
         q_4_5 : OUT std_logic ;
         q_4_4 : OUT std_logic ;
         q_4_3 : OUT std_logic ;
         q_4_2 : OUT std_logic ;
         q_4_1 : OUT std_logic ;
         q_4_0 : OUT std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         reset : IN std_logic) ;
   end component ;
   component Queue_25
      port (
         d : IN std_logic_vector (15 DOWNTO 0) ;
         q_0_15 : OUT std_logic ;
         q_0_14 : OUT std_logic ;
         q_0_13 : OUT std_logic ;
         q_0_12 : OUT std_logic ;
         q_0_11 : OUT std_logic ;
         q_0_10 : OUT std_logic ;
         q_0_9 : OUT std_logic ;
         q_0_8 : OUT std_logic ;
         q_0_7 : OUT std_logic ;
         q_0_6 : OUT std_logic ;
         q_0_5 : OUT std_logic ;
         q_0_4 : OUT std_logic ;
         q_0_3 : OUT std_logic ;
         q_0_2 : OUT std_logic ;
         q_0_1 : OUT std_logic ;
         q_0_0 : OUT std_logic ;
         q_1_15 : OUT std_logic ;
         q_1_14 : OUT std_logic ;
         q_1_13 : OUT std_logic ;
         q_1_12 : OUT std_logic ;
         q_1_11 : OUT std_logic ;
         q_1_10 : OUT std_logic ;
         q_1_9 : OUT std_logic ;
         q_1_8 : OUT std_logic ;
         q_1_7 : OUT std_logic ;
         q_1_6 : OUT std_logic ;
         q_1_5 : OUT std_logic ;
         q_1_4 : OUT std_logic ;
         q_1_3 : OUT std_logic ;
         q_1_2 : OUT std_logic ;
         q_1_1 : OUT std_logic ;
         q_1_0 : OUT std_logic ;
         q_2_15 : OUT std_logic ;
         q_2_14 : OUT std_logic ;
         q_2_13 : OUT std_logic ;
         q_2_12 : OUT std_logic ;
         q_2_11 : OUT std_logic ;
         q_2_10 : OUT std_logic ;
         q_2_9 : OUT std_logic ;
         q_2_8 : OUT std_logic ;
         q_2_7 : OUT std_logic ;
         q_2_6 : OUT std_logic ;
         q_2_5 : OUT std_logic ;
         q_2_4 : OUT std_logic ;
         q_2_3 : OUT std_logic ;
         q_2_2 : OUT std_logic ;
         q_2_1 : OUT std_logic ;
         q_2_0 : OUT std_logic ;
         q_3_15 : OUT std_logic ;
         q_3_14 : OUT std_logic ;
         q_3_13 : OUT std_logic ;
         q_3_12 : OUT std_logic ;
         q_3_11 : OUT std_logic ;
         q_3_10 : OUT std_logic ;
         q_3_9 : OUT std_logic ;
         q_3_8 : OUT std_logic ;
         q_3_7 : OUT std_logic ;
         q_3_6 : OUT std_logic ;
         q_3_5 : OUT std_logic ;
         q_3_4 : OUT std_logic ;
         q_3_3 : OUT std_logic ;
         q_3_2 : OUT std_logic ;
         q_3_1 : OUT std_logic ;
         q_3_0 : OUT std_logic ;
         q_4_15 : OUT std_logic ;
         q_4_14 : OUT std_logic ;
         q_4_13 : OUT std_logic ;
         q_4_12 : OUT std_logic ;
         q_4_11 : OUT std_logic ;
         q_4_10 : OUT std_logic ;
         q_4_9 : OUT std_logic ;
         q_4_8 : OUT std_logic ;
         q_4_7 : OUT std_logic ;
         q_4_6 : OUT std_logic ;
         q_4_5 : OUT std_logic ;
         q_4_4 : OUT std_logic ;
         q_4_3 : OUT std_logic ;
         q_4_2 : OUT std_logic ;
         q_4_1 : OUT std_logic ;
         q_4_0 : OUT std_logic ;
         q_5_15 : OUT std_logic ;
         q_5_14 : OUT std_logic ;
         q_5_13 : OUT std_logic ;
         q_5_12 : OUT std_logic ;
         q_5_11 : OUT std_logic ;
         q_5_10 : OUT std_logic ;
         q_5_9 : OUT std_logic ;
         q_5_8 : OUT std_logic ;
         q_5_7 : OUT std_logic ;
         q_5_6 : OUT std_logic ;
         q_5_5 : OUT std_logic ;
         q_5_4 : OUT std_logic ;
         q_5_3 : OUT std_logic ;
         q_5_2 : OUT std_logic ;
         q_5_1 : OUT std_logic ;
         q_5_0 : OUT std_logic ;
         q_6_15 : OUT std_logic ;
         q_6_14 : OUT std_logic ;
         q_6_13 : OUT std_logic ;
         q_6_12 : OUT std_logic ;
         q_6_11 : OUT std_logic ;
         q_6_10 : OUT std_logic ;
         q_6_9 : OUT std_logic ;
         q_6_8 : OUT std_logic ;
         q_6_7 : OUT std_logic ;
         q_6_6 : OUT std_logic ;
         q_6_5 : OUT std_logic ;
         q_6_4 : OUT std_logic ;
         q_6_3 : OUT std_logic ;
         q_6_2 : OUT std_logic ;
         q_6_1 : OUT std_logic ;
         q_6_0 : OUT std_logic ;
         q_7_15 : OUT std_logic ;
         q_7_14 : OUT std_logic ;
         q_7_13 : OUT std_logic ;
         q_7_12 : OUT std_logic ;
         q_7_11 : OUT std_logic ;
         q_7_10 : OUT std_logic ;
         q_7_9 : OUT std_logic ;
         q_7_8 : OUT std_logic ;
         q_7_7 : OUT std_logic ;
         q_7_6 : OUT std_logic ;
         q_7_5 : OUT std_logic ;
         q_7_4 : OUT std_logic ;
         q_7_3 : OUT std_logic ;
         q_7_2 : OUT std_logic ;
         q_7_1 : OUT std_logic ;
         q_7_0 : OUT std_logic ;
         q_8_15 : OUT std_logic ;
         q_8_14 : OUT std_logic ;
         q_8_13 : OUT std_logic ;
         q_8_12 : OUT std_logic ;
         q_8_11 : OUT std_logic ;
         q_8_10 : OUT std_logic ;
         q_8_9 : OUT std_logic ;
         q_8_8 : OUT std_logic ;
         q_8_7 : OUT std_logic ;
         q_8_6 : OUT std_logic ;
         q_8_5 : OUT std_logic ;
         q_8_4 : OUT std_logic ;
         q_8_3 : OUT std_logic ;
         q_8_2 : OUT std_logic ;
         q_8_1 : OUT std_logic ;
         q_8_0 : OUT std_logic ;
         q_9_15 : OUT std_logic ;
         q_9_14 : OUT std_logic ;
         q_9_13 : OUT std_logic ;
         q_9_12 : OUT std_logic ;
         q_9_11 : OUT std_logic ;
         q_9_10 : OUT std_logic ;
         q_9_9 : OUT std_logic ;
         q_9_8 : OUT std_logic ;
         q_9_7 : OUT std_logic ;
         q_9_6 : OUT std_logic ;
         q_9_5 : OUT std_logic ;
         q_9_4 : OUT std_logic ;
         q_9_3 : OUT std_logic ;
         q_9_2 : OUT std_logic ;
         q_9_1 : OUT std_logic ;
         q_9_0 : OUT std_logic ;
         q_10_15 : OUT std_logic ;
         q_10_14 : OUT std_logic ;
         q_10_13 : OUT std_logic ;
         q_10_12 : OUT std_logic ;
         q_10_11 : OUT std_logic ;
         q_10_10 : OUT std_logic ;
         q_10_9 : OUT std_logic ;
         q_10_8 : OUT std_logic ;
         q_10_7 : OUT std_logic ;
         q_10_6 : OUT std_logic ;
         q_10_5 : OUT std_logic ;
         q_10_4 : OUT std_logic ;
         q_10_3 : OUT std_logic ;
         q_10_2 : OUT std_logic ;
         q_10_1 : OUT std_logic ;
         q_10_0 : OUT std_logic ;
         q_11_15 : OUT std_logic ;
         q_11_14 : OUT std_logic ;
         q_11_13 : OUT std_logic ;
         q_11_12 : OUT std_logic ;
         q_11_11 : OUT std_logic ;
         q_11_10 : OUT std_logic ;
         q_11_9 : OUT std_logic ;
         q_11_8 : OUT std_logic ;
         q_11_7 : OUT std_logic ;
         q_11_6 : OUT std_logic ;
         q_11_5 : OUT std_logic ;
         q_11_4 : OUT std_logic ;
         q_11_3 : OUT std_logic ;
         q_11_2 : OUT std_logic ;
         q_11_1 : OUT std_logic ;
         q_11_0 : OUT std_logic ;
         q_12_15 : OUT std_logic ;
         q_12_14 : OUT std_logic ;
         q_12_13 : OUT std_logic ;
         q_12_12 : OUT std_logic ;
         q_12_11 : OUT std_logic ;
         q_12_10 : OUT std_logic ;
         q_12_9 : OUT std_logic ;
         q_12_8 : OUT std_logic ;
         q_12_7 : OUT std_logic ;
         q_12_6 : OUT std_logic ;
         q_12_5 : OUT std_logic ;
         q_12_4 : OUT std_logic ;
         q_12_3 : OUT std_logic ;
         q_12_2 : OUT std_logic ;
         q_12_1 : OUT std_logic ;
         q_12_0 : OUT std_logic ;
         q_13_15 : OUT std_logic ;
         q_13_14 : OUT std_logic ;
         q_13_13 : OUT std_logic ;
         q_13_12 : OUT std_logic ;
         q_13_11 : OUT std_logic ;
         q_13_10 : OUT std_logic ;
         q_13_9 : OUT std_logic ;
         q_13_8 : OUT std_logic ;
         q_13_7 : OUT std_logic ;
         q_13_6 : OUT std_logic ;
         q_13_5 : OUT std_logic ;
         q_13_4 : OUT std_logic ;
         q_13_3 : OUT std_logic ;
         q_13_2 : OUT std_logic ;
         q_13_1 : OUT std_logic ;
         q_13_0 : OUT std_logic ;
         q_14_15 : OUT std_logic ;
         q_14_14 : OUT std_logic ;
         q_14_13 : OUT std_logic ;
         q_14_12 : OUT std_logic ;
         q_14_11 : OUT std_logic ;
         q_14_10 : OUT std_logic ;
         q_14_9 : OUT std_logic ;
         q_14_8 : OUT std_logic ;
         q_14_7 : OUT std_logic ;
         q_14_6 : OUT std_logic ;
         q_14_5 : OUT std_logic ;
         q_14_4 : OUT std_logic ;
         q_14_3 : OUT std_logic ;
         q_14_2 : OUT std_logic ;
         q_14_1 : OUT std_logic ;
         q_14_0 : OUT std_logic ;
         q_15_15 : OUT std_logic ;
         q_15_14 : OUT std_logic ;
         q_15_13 : OUT std_logic ;
         q_15_12 : OUT std_logic ;
         q_15_11 : OUT std_logic ;
         q_15_10 : OUT std_logic ;
         q_15_9 : OUT std_logic ;
         q_15_8 : OUT std_logic ;
         q_15_7 : OUT std_logic ;
         q_15_6 : OUT std_logic ;
         q_15_5 : OUT std_logic ;
         q_15_4 : OUT std_logic ;
         q_15_3 : OUT std_logic ;
         q_15_2 : OUT std_logic ;
         q_15_1 : OUT std_logic ;
         q_15_0 : OUT std_logic ;
         q_16_15 : OUT std_logic ;
         q_16_14 : OUT std_logic ;
         q_16_13 : OUT std_logic ;
         q_16_12 : OUT std_logic ;
         q_16_11 : OUT std_logic ;
         q_16_10 : OUT std_logic ;
         q_16_9 : OUT std_logic ;
         q_16_8 : OUT std_logic ;
         q_16_7 : OUT std_logic ;
         q_16_6 : OUT std_logic ;
         q_16_5 : OUT std_logic ;
         q_16_4 : OUT std_logic ;
         q_16_3 : OUT std_logic ;
         q_16_2 : OUT std_logic ;
         q_16_1 : OUT std_logic ;
         q_16_0 : OUT std_logic ;
         q_17_15 : OUT std_logic ;
         q_17_14 : OUT std_logic ;
         q_17_13 : OUT std_logic ;
         q_17_12 : OUT std_logic ;
         q_17_11 : OUT std_logic ;
         q_17_10 : OUT std_logic ;
         q_17_9 : OUT std_logic ;
         q_17_8 : OUT std_logic ;
         q_17_7 : OUT std_logic ;
         q_17_6 : OUT std_logic ;
         q_17_5 : OUT std_logic ;
         q_17_4 : OUT std_logic ;
         q_17_3 : OUT std_logic ;
         q_17_2 : OUT std_logic ;
         q_17_1 : OUT std_logic ;
         q_17_0 : OUT std_logic ;
         q_18_15 : OUT std_logic ;
         q_18_14 : OUT std_logic ;
         q_18_13 : OUT std_logic ;
         q_18_12 : OUT std_logic ;
         q_18_11 : OUT std_logic ;
         q_18_10 : OUT std_logic ;
         q_18_9 : OUT std_logic ;
         q_18_8 : OUT std_logic ;
         q_18_7 : OUT std_logic ;
         q_18_6 : OUT std_logic ;
         q_18_5 : OUT std_logic ;
         q_18_4 : OUT std_logic ;
         q_18_3 : OUT std_logic ;
         q_18_2 : OUT std_logic ;
         q_18_1 : OUT std_logic ;
         q_18_0 : OUT std_logic ;
         q_19_15 : OUT std_logic ;
         q_19_14 : OUT std_logic ;
         q_19_13 : OUT std_logic ;
         q_19_12 : OUT std_logic ;
         q_19_11 : OUT std_logic ;
         q_19_10 : OUT std_logic ;
         q_19_9 : OUT std_logic ;
         q_19_8 : OUT std_logic ;
         q_19_7 : OUT std_logic ;
         q_19_6 : OUT std_logic ;
         q_19_5 : OUT std_logic ;
         q_19_4 : OUT std_logic ;
         q_19_3 : OUT std_logic ;
         q_19_2 : OUT std_logic ;
         q_19_1 : OUT std_logic ;
         q_19_0 : OUT std_logic ;
         q_20_15 : OUT std_logic ;
         q_20_14 : OUT std_logic ;
         q_20_13 : OUT std_logic ;
         q_20_12 : OUT std_logic ;
         q_20_11 : OUT std_logic ;
         q_20_10 : OUT std_logic ;
         q_20_9 : OUT std_logic ;
         q_20_8 : OUT std_logic ;
         q_20_7 : OUT std_logic ;
         q_20_6 : OUT std_logic ;
         q_20_5 : OUT std_logic ;
         q_20_4 : OUT std_logic ;
         q_20_3 : OUT std_logic ;
         q_20_2 : OUT std_logic ;
         q_20_1 : OUT std_logic ;
         q_20_0 : OUT std_logic ;
         q_21_15 : OUT std_logic ;
         q_21_14 : OUT std_logic ;
         q_21_13 : OUT std_logic ;
         q_21_12 : OUT std_logic ;
         q_21_11 : OUT std_logic ;
         q_21_10 : OUT std_logic ;
         q_21_9 : OUT std_logic ;
         q_21_8 : OUT std_logic ;
         q_21_7 : OUT std_logic ;
         q_21_6 : OUT std_logic ;
         q_21_5 : OUT std_logic ;
         q_21_4 : OUT std_logic ;
         q_21_3 : OUT std_logic ;
         q_21_2 : OUT std_logic ;
         q_21_1 : OUT std_logic ;
         q_21_0 : OUT std_logic ;
         q_22_15 : OUT std_logic ;
         q_22_14 : OUT std_logic ;
         q_22_13 : OUT std_logic ;
         q_22_12 : OUT std_logic ;
         q_22_11 : OUT std_logic ;
         q_22_10 : OUT std_logic ;
         q_22_9 : OUT std_logic ;
         q_22_8 : OUT std_logic ;
         q_22_7 : OUT std_logic ;
         q_22_6 : OUT std_logic ;
         q_22_5 : OUT std_logic ;
         q_22_4 : OUT std_logic ;
         q_22_3 : OUT std_logic ;
         q_22_2 : OUT std_logic ;
         q_22_1 : OUT std_logic ;
         q_22_0 : OUT std_logic ;
         q_23_15 : OUT std_logic ;
         q_23_14 : OUT std_logic ;
         q_23_13 : OUT std_logic ;
         q_23_12 : OUT std_logic ;
         q_23_11 : OUT std_logic ;
         q_23_10 : OUT std_logic ;
         q_23_9 : OUT std_logic ;
         q_23_8 : OUT std_logic ;
         q_23_7 : OUT std_logic ;
         q_23_6 : OUT std_logic ;
         q_23_5 : OUT std_logic ;
         q_23_4 : OUT std_logic ;
         q_23_3 : OUT std_logic ;
         q_23_2 : OUT std_logic ;
         q_23_1 : OUT std_logic ;
         q_23_0 : OUT std_logic ;
         q_24_15 : OUT std_logic ;
         q_24_14 : OUT std_logic ;
         q_24_13 : OUT std_logic ;
         q_24_12 : OUT std_logic ;
         q_24_11 : OUT std_logic ;
         q_24_10 : OUT std_logic ;
         q_24_9 : OUT std_logic ;
         q_24_8 : OUT std_logic ;
         q_24_7 : OUT std_logic ;
         q_24_6 : OUT std_logic ;
         q_24_5 : OUT std_logic ;
         q_24_4 : OUT std_logic ;
         q_24_3 : OUT std_logic ;
         q_24_2 : OUT std_logic ;
         q_24_1 : OUT std_logic ;
         q_24_0 : OUT std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         reset : IN std_logic) ;
   end component ;
   component Reg_32
      port (
         d : IN std_logic_vector (31 DOWNTO 0) ;
         q : OUT std_logic_vector (31 DOWNTO 0) ;
         rst_data : IN std_logic_vector (31 DOWNTO 0) ;
         clk : IN std_logic ;
         load : IN std_logic ;
         reset : IN std_logic) ;
   end component ;
   signal output1_15_EXMPLR, output1_14_EXMPLR, output1_13_EXMPLR, 
      output1_12_EXMPLR, output1_11_EXMPLR, output1_10_EXMPLR, 
      output1_9_EXMPLR, output1_8_EXMPLR, output1_7_EXMPLR, output1_6_EXMPLR, 
      output1_5_EXMPLR, output1_4_EXMPLR, output1_3_EXMPLR, output1_2_EXMPLR, 
      output1_1_EXMPLR, output1_0_EXMPLR, output2_15_EXMPLR, 
      output2_14_EXMPLR, output2_13_EXMPLR, output2_12_EXMPLR, 
      output2_11_EXMPLR, output2_10_EXMPLR, output2_9_EXMPLR, 
      output2_8_EXMPLR, output2_7_EXMPLR, output2_6_EXMPLR, output2_5_EXMPLR, 
      output2_4_EXMPLR, output2_3_EXMPLR, output2_2_EXMPLR, output2_1_EXMPLR, 
      output2_0_EXMPLR, ready_EXMPLR, img_data_0_15, img_data_0_14, 
      img_data_0_13, img_data_0_12, img_data_0_11, img_data_0_10, 
      img_data_0_9, img_data_0_8, img_data_0_7, img_data_0_6, img_data_0_5, 
      img_data_0_4, img_data_0_3, img_data_0_2, img_data_0_1, img_data_0_0, 
      img_data_1_15, img_data_1_14, img_data_1_13, img_data_1_12, 
      img_data_1_11, img_data_1_10, img_data_1_9, img_data_1_8, img_data_1_7, 
      img_data_1_6, img_data_1_5, img_data_1_4, img_data_1_3, img_data_1_2, 
      img_data_1_1, img_data_1_0, img_data_2_15, img_data_2_14, 
      img_data_2_13, img_data_2_12, img_data_2_11, img_data_2_10, 
      img_data_2_9, img_data_2_8, img_data_2_7, img_data_2_6, img_data_2_5, 
      img_data_2_4, img_data_2_3, img_data_2_2, img_data_2_1, img_data_2_0, 
      img_data_3_15, img_data_3_14, img_data_3_13, img_data_3_12, 
      img_data_3_11, img_data_3_10, img_data_3_9, img_data_3_8, img_data_3_7, 
      img_data_3_6, img_data_3_5, img_data_3_4, img_data_3_3, img_data_3_2, 
      img_data_3_1, img_data_3_0, img_data_4_15, img_data_4_14, 
      img_data_4_13, img_data_4_12, img_data_4_11, img_data_4_10, 
      img_data_4_9, img_data_4_8, img_data_4_7, img_data_4_6, img_data_4_5, 
      img_data_4_4, img_data_4_3, img_data_4_2, img_data_4_1, img_data_4_0, 
      img_data_5_15, img_data_5_14, img_data_5_13, img_data_5_12, 
      img_data_5_11, img_data_5_10, img_data_5_9, img_data_5_8, img_data_5_7, 
      img_data_5_6, img_data_5_5, img_data_5_4, img_data_5_3, img_data_5_2, 
      img_data_5_1, img_data_5_0, img_data_6_15, img_data_6_14, 
      img_data_6_13, img_data_6_12, img_data_6_11, img_data_6_10, 
      img_data_6_9, img_data_6_8, img_data_6_7, img_data_6_6, img_data_6_5, 
      img_data_6_4, img_data_6_3, img_data_6_2, img_data_6_1, img_data_6_0, 
      img_data_7_15, img_data_7_14, img_data_7_13, img_data_7_12, 
      img_data_7_11, img_data_7_10, img_data_7_9, img_data_7_8, img_data_7_7, 
      img_data_7_6, img_data_7_5, img_data_7_4, img_data_7_3, img_data_7_2, 
      img_data_7_1, img_data_7_0, img_data_8_15, img_data_8_14, 
      img_data_8_13, img_data_8_12, img_data_8_11, img_data_8_10, 
      img_data_8_9, img_data_8_8, img_data_8_7, img_data_8_6, img_data_8_5, 
      img_data_8_4, img_data_8_3, img_data_8_2, img_data_8_1, img_data_8_0, 
      img_data_9_15, img_data_9_14, img_data_9_13, img_data_9_12, 
      img_data_9_11, img_data_9_10, img_data_9_9, img_data_9_8, img_data_9_7, 
      img_data_9_6, img_data_9_5, img_data_9_4, img_data_9_3, img_data_9_2, 
      img_data_9_1, img_data_9_0, img_data_10_15, img_data_10_14, 
      img_data_10_13, img_data_10_12, img_data_10_11, img_data_10_10, 
      img_data_10_9, img_data_10_8, img_data_10_7, img_data_10_6, 
      img_data_10_5, img_data_10_4, img_data_10_3, img_data_10_2, 
      img_data_10_1, img_data_10_0, img_data_11_15, img_data_11_14, 
      img_data_11_13, img_data_11_12, img_data_11_11, img_data_11_10, 
      img_data_11_9, img_data_11_8, img_data_11_7, img_data_11_6, 
      img_data_11_5, img_data_11_4, img_data_11_3, img_data_11_2, 
      img_data_11_1, img_data_11_0, img_data_12_15, img_data_12_14, 
      img_data_12_13, img_data_12_12, img_data_12_11, img_data_12_10, 
      img_data_12_9, img_data_12_8, img_data_12_7, img_data_12_6, 
      img_data_12_5, img_data_12_4, img_data_12_3, img_data_12_2, 
      img_data_12_1, img_data_12_0, img_data_13_15, img_data_13_14, 
      img_data_13_13, img_data_13_12, img_data_13_11, img_data_13_10, 
      img_data_13_9, img_data_13_8, img_data_13_7, img_data_13_6, 
      img_data_13_5, img_data_13_4, img_data_13_3, img_data_13_2, 
      img_data_13_1, img_data_13_0, img_data_14_15, img_data_14_14, 
      img_data_14_13, img_data_14_12, img_data_14_11, img_data_14_10, 
      img_data_14_9, img_data_14_8, img_data_14_7, img_data_14_6, 
      img_data_14_5, img_data_14_4, img_data_14_3, img_data_14_2, 
      img_data_14_1, img_data_14_0, img_data_15_15, img_data_15_14, 
      img_data_15_13, img_data_15_12, img_data_15_11, img_data_15_10, 
      img_data_15_9, img_data_15_8, img_data_15_7, img_data_15_6, 
      img_data_15_5, img_data_15_4, img_data_15_3, img_data_15_2, 
      img_data_15_1, img_data_15_0, img_data_16_15, img_data_16_14, 
      img_data_16_13, img_data_16_12, img_data_16_11, img_data_16_10, 
      img_data_16_9, img_data_16_8, img_data_16_7, img_data_16_6, 
      img_data_16_5, img_data_16_4, img_data_16_3, img_data_16_2, 
      img_data_16_1, img_data_16_0, img_data_17_15, img_data_17_14, 
      img_data_17_13, img_data_17_12, img_data_17_11, img_data_17_10, 
      img_data_17_9, img_data_17_8, img_data_17_7, img_data_17_6, 
      img_data_17_5, img_data_17_4, img_data_17_3, img_data_17_2, 
      img_data_17_1, img_data_17_0, img_data_18_15, img_data_18_14, 
      img_data_18_13, img_data_18_12, img_data_18_11, img_data_18_10, 
      img_data_18_9, img_data_18_8, img_data_18_7, img_data_18_6, 
      img_data_18_5, img_data_18_4, img_data_18_3, img_data_18_2, 
      img_data_18_1, img_data_18_0, img_data_19_15, img_data_19_14, 
      img_data_19_13, img_data_19_12, img_data_19_11, img_data_19_10, 
      img_data_19_9, img_data_19_8, img_data_19_7, img_data_19_6, 
      img_data_19_5, img_data_19_4, img_data_19_3, img_data_19_2, 
      img_data_19_1, img_data_19_0, img_data_20_15, img_data_20_14, 
      img_data_20_13, img_data_20_12, img_data_20_11, img_data_20_10, 
      img_data_20_9, img_data_20_8, img_data_20_7, img_data_20_6, 
      img_data_20_5, img_data_20_4, img_data_20_3, img_data_20_2, 
      img_data_20_1, img_data_20_0, img_data_21_15, img_data_21_14, 
      img_data_21_13, img_data_21_12, img_data_21_11, img_data_21_10, 
      img_data_21_9, img_data_21_8, img_data_21_7, img_data_21_6, 
      img_data_21_5, img_data_21_4, img_data_21_3, img_data_21_2, 
      img_data_21_1, img_data_21_0, img_data_22_15, img_data_22_14, 
      img_data_22_13, img_data_22_12, img_data_22_11, img_data_22_10, 
      img_data_22_9, img_data_22_8, img_data_22_7, img_data_22_6, 
      img_data_22_5, img_data_22_4, img_data_22_3, img_data_22_2, 
      img_data_22_1, img_data_22_0, img_data_23_15, img_data_23_14, 
      img_data_23_13, img_data_23_12, img_data_23_11, img_data_23_10, 
      img_data_23_9, img_data_23_8, img_data_23_7, img_data_23_6, 
      img_data_23_5, img_data_23_4, img_data_23_3, img_data_23_2, 
      img_data_23_1, img_data_23_0, img_data_24_15, img_data_24_14, 
      img_data_24_13, img_data_24_12, img_data_24_11, img_data_24_10, 
      img_data_24_9, img_data_24_8, img_data_24_7, img_data_24_6, 
      img_data_24_5, img_data_24_4, img_data_24_3, img_data_24_2, 
      img_data_24_1, img_data_24_0, filter_data_0_15, filter_data_0_14, 
      filter_data_0_13, filter_data_0_12, filter_data_0_11, filter_data_0_10, 
      filter_data_0_9, filter_data_0_8, filter_data_0_7, filter_data_0_6, 
      filter_data_0_5, filter_data_0_4, filter_data_0_3, filter_data_0_2, 
      filter_data_0_1, filter_data_0_0, filter_data_1_15, filter_data_1_14, 
      filter_data_1_13, filter_data_1_12, filter_data_1_11, filter_data_1_10, 
      filter_data_1_9, filter_data_1_8, filter_data_1_7, filter_data_1_6, 
      filter_data_1_5, filter_data_1_4, filter_data_1_3, filter_data_1_2, 
      filter_data_1_1, filter_data_1_0, filter_data_2_15, filter_data_2_14, 
      filter_data_2_13, filter_data_2_12, filter_data_2_11, filter_data_2_10, 
      filter_data_2_9, filter_data_2_8, filter_data_2_7, filter_data_2_6, 
      filter_data_2_5, filter_data_2_4, filter_data_2_3, filter_data_2_2, 
      filter_data_2_1, filter_data_2_0, filter_data_3_15, filter_data_3_14, 
      filter_data_3_13, filter_data_3_12, filter_data_3_11, filter_data_3_10, 
      filter_data_3_9, filter_data_3_8, filter_data_3_7, filter_data_3_6, 
      filter_data_3_5, filter_data_3_4, filter_data_3_3, filter_data_3_2, 
      filter_data_3_1, filter_data_3_0, filter_data_4_15, filter_data_4_14, 
      filter_data_4_13, filter_data_4_12, filter_data_4_11, filter_data_4_10, 
      filter_data_4_9, filter_data_4_8, filter_data_4_7, filter_data_4_6, 
      filter_data_4_5, filter_data_4_4, filter_data_4_3, filter_data_4_2, 
      filter_data_4_1, filter_data_4_0, filter_data_5_15, filter_data_5_14, 
      filter_data_5_13, filter_data_5_12, filter_data_5_11, filter_data_5_10, 
      filter_data_5_9, filter_data_5_8, filter_data_5_7, filter_data_5_6, 
      filter_data_5_5, filter_data_5_4, filter_data_5_3, filter_data_5_2, 
      filter_data_5_1, filter_data_5_0, filter_data_6_15, filter_data_6_14, 
      filter_data_6_13, filter_data_6_12, filter_data_6_11, filter_data_6_10, 
      filter_data_6_9, filter_data_6_8, filter_data_6_7, filter_data_6_6, 
      filter_data_6_5, filter_data_6_4, filter_data_6_3, filter_data_6_2, 
      filter_data_6_1, filter_data_6_0, filter_data_7_15, filter_data_7_14, 
      filter_data_7_13, filter_data_7_12, filter_data_7_11, filter_data_7_10, 
      filter_data_7_9, filter_data_7_8, filter_data_7_7, filter_data_7_6, 
      filter_data_7_5, filter_data_7_4, filter_data_7_3, filter_data_7_2, 
      filter_data_7_1, filter_data_7_0, filter_data_8_15, filter_data_8_14, 
      filter_data_8_13, filter_data_8_12, filter_data_8_11, filter_data_8_10, 
      filter_data_8_9, filter_data_8_8, filter_data_8_7, filter_data_8_6, 
      filter_data_8_5, filter_data_8_4, filter_data_8_3, filter_data_8_2, 
      filter_data_8_1, filter_data_8_0, filter_data_9_15, filter_data_9_14, 
      filter_data_9_13, filter_data_9_12, filter_data_9_11, filter_data_9_10, 
      filter_data_9_9, filter_data_9_8, filter_data_9_7, filter_data_9_6, 
      filter_data_9_5, filter_data_9_4, filter_data_9_3, filter_data_9_2, 
      filter_data_9_1, filter_data_9_0, filter_data_10_15, filter_data_10_14, 
      filter_data_10_13, filter_data_10_12, filter_data_10_11, 
      filter_data_10_10, filter_data_10_9, filter_data_10_8, 
      filter_data_10_7, filter_data_10_6, filter_data_10_5, filter_data_10_4, 
      filter_data_10_3, filter_data_10_2, filter_data_10_1, filter_data_10_0, 
      filter_data_11_15, filter_data_11_14, filter_data_11_13, 
      filter_data_11_12, filter_data_11_11, filter_data_11_10, 
      filter_data_11_9, filter_data_11_8, filter_data_11_7, filter_data_11_6, 
      filter_data_11_5, filter_data_11_4, filter_data_11_3, filter_data_11_2, 
      filter_data_11_1, filter_data_11_0, filter_data_12_15, 
      filter_data_12_14, filter_data_12_13, filter_data_12_12, 
      filter_data_12_11, filter_data_12_10, filter_data_12_9, 
      filter_data_12_8, filter_data_12_7, filter_data_12_6, filter_data_12_5, 
      filter_data_12_4, filter_data_12_3, filter_data_12_2, filter_data_12_1, 
      filter_data_12_0, filter_data_13_15, filter_data_13_14, 
      filter_data_13_13, filter_data_13_12, filter_data_13_11, 
      filter_data_13_10, filter_data_13_9, filter_data_13_8, 
      filter_data_13_7, filter_data_13_6, filter_data_13_5, filter_data_13_4, 
      filter_data_13_3, filter_data_13_2, filter_data_13_1, filter_data_13_0, 
      filter_data_14_15, filter_data_14_14, filter_data_14_13, 
      filter_data_14_12, filter_data_14_11, filter_data_14_10, 
      filter_data_14_9, filter_data_14_8, filter_data_14_7, filter_data_14_6, 
      filter_data_14_5, filter_data_14_4, filter_data_14_3, filter_data_14_2, 
      filter_data_14_1, filter_data_14_0, filter_data_15_15, 
      filter_data_15_14, filter_data_15_13, filter_data_15_12, 
      filter_data_15_11, filter_data_15_10, filter_data_15_9, 
      filter_data_15_8, filter_data_15_7, filter_data_15_6, filter_data_15_5, 
      filter_data_15_4, filter_data_15_3, filter_data_15_2, filter_data_15_1, 
      filter_data_15_0, filter_data_16_15, filter_data_16_14, 
      filter_data_16_13, filter_data_16_12, filter_data_16_11, 
      filter_data_16_10, filter_data_16_9, filter_data_16_8, 
      filter_data_16_7, filter_data_16_6, filter_data_16_5, filter_data_16_4, 
      filter_data_16_3, filter_data_16_2, filter_data_16_1, filter_data_16_0, 
      filter_data_17_15, filter_data_17_14, filter_data_17_13, 
      filter_data_17_12, filter_data_17_11, filter_data_17_10, 
      filter_data_17_9, filter_data_17_8, filter_data_17_7, filter_data_17_6, 
      filter_data_17_5, filter_data_17_4, filter_data_17_3, filter_data_17_2, 
      filter_data_17_1, filter_data_17_0, filter_data_18_15, 
      filter_data_18_14, filter_data_18_13, filter_data_18_12, 
      filter_data_18_11, filter_data_18_10, filter_data_18_9, 
      filter_data_18_8, filter_data_18_7, filter_data_18_6, filter_data_18_5, 
      filter_data_18_4, filter_data_18_3, filter_data_18_2, filter_data_18_1, 
      filter_data_18_0, filter_data_19_15, filter_data_19_14, 
      filter_data_19_13, filter_data_19_12, filter_data_19_11, 
      filter_data_19_10, filter_data_19_9, filter_data_19_8, 
      filter_data_19_7, filter_data_19_6, filter_data_19_5, filter_data_19_4, 
      filter_data_19_3, filter_data_19_2, filter_data_19_1, filter_data_19_0, 
      filter_data_20_15, filter_data_20_14, filter_data_20_13, 
      filter_data_20_12, filter_data_20_11, filter_data_20_10, 
      filter_data_20_9, filter_data_20_8, filter_data_20_7, filter_data_20_6, 
      filter_data_20_5, filter_data_20_4, filter_data_20_3, filter_data_20_2, 
      filter_data_20_1, filter_data_20_0, filter_data_21_15, 
      filter_data_21_14, filter_data_21_13, filter_data_21_12, 
      filter_data_21_11, filter_data_21_10, filter_data_21_9, 
      filter_data_21_8, filter_data_21_7, filter_data_21_6, filter_data_21_5, 
      filter_data_21_4, filter_data_21_3, filter_data_21_2, filter_data_21_1, 
      filter_data_21_0, filter_data_22_15, filter_data_22_14, 
      filter_data_22_13, filter_data_22_12, filter_data_22_11, 
      filter_data_22_10, filter_data_22_9, filter_data_22_8, 
      filter_data_22_7, filter_data_22_6, filter_data_22_5, filter_data_22_4, 
      filter_data_22_3, filter_data_22_2, filter_data_22_1, filter_data_22_0, 
      filter_data_23_15, filter_data_23_14, filter_data_23_13, 
      filter_data_23_12, filter_data_23_11, filter_data_23_10, 
      filter_data_23_9, filter_data_23_8, filter_data_23_7, filter_data_23_6, 
      filter_data_23_5, filter_data_23_4, filter_data_23_3, filter_data_23_2, 
      filter_data_23_1, filter_data_23_0, filter_data_24_15, 
      filter_data_24_14, filter_data_24_13, filter_data_24_12, 
      filter_data_24_11, filter_data_24_10, filter_data_24_9, 
      filter_data_24_8, filter_data_24_7, filter_data_24_6, filter_data_24_5, 
      filter_data_24_4, filter_data_24_3, filter_data_24_2, filter_data_24_1, 
      filter_data_24_0, d_cache_arr_0_31, d_cache_arr_0_30, d_cache_arr_0_29, 
      d_cache_arr_0_28, d_cache_arr_0_27, d_cache_arr_0_26, d_cache_arr_0_25, 
      d_cache_arr_0_24, d_cache_arr_0_23, d_cache_arr_0_22, d_cache_arr_0_21, 
      d_cache_arr_0_20, d_cache_arr_0_19, d_cache_arr_0_18, d_cache_arr_0_17, 
      d_cache_arr_0_16, d_cache_arr_0_15, d_cache_arr_0_14, d_cache_arr_0_13, 
      d_cache_arr_0_12, d_cache_arr_0_11, d_cache_arr_0_10, d_cache_arr_0_9, 
      d_cache_arr_0_8, d_cache_arr_0_7, d_cache_arr_0_6, d_cache_arr_0_5, 
      d_cache_arr_0_4, d_cache_arr_0_3, d_cache_arr_0_2, d_cache_arr_0_1, 
      d_cache_arr_0_0, d_cache_arr_1_31, d_cache_arr_1_30, d_cache_arr_1_29, 
      d_cache_arr_1_28, d_cache_arr_1_27, d_cache_arr_1_26, d_cache_arr_1_25, 
      d_cache_arr_1_24, d_cache_arr_1_23, d_cache_arr_1_22, d_cache_arr_1_21, 
      d_cache_arr_1_20, d_cache_arr_1_19, d_cache_arr_1_18, d_cache_arr_1_17, 
      d_cache_arr_1_16, d_cache_arr_1_15, d_cache_arr_1_14, d_cache_arr_1_13, 
      d_cache_arr_1_12, d_cache_arr_1_11, d_cache_arr_1_10, d_cache_arr_1_9, 
      d_cache_arr_1_8, d_cache_arr_1_7, d_cache_arr_1_6, d_cache_arr_1_5, 
      d_cache_arr_1_4, d_cache_arr_1_3, d_cache_arr_1_2, d_cache_arr_1_1, 
      d_cache_arr_1_0, d_cache_arr_2_31, d_cache_arr_2_30, d_cache_arr_2_29, 
      d_cache_arr_2_28, d_cache_arr_2_27, d_cache_arr_2_26, d_cache_arr_2_25, 
      d_cache_arr_2_24, d_cache_arr_2_23, d_cache_arr_2_22, d_cache_arr_2_21, 
      d_cache_arr_2_20, d_cache_arr_2_19, d_cache_arr_2_18, d_cache_arr_2_17, 
      d_cache_arr_2_16, d_cache_arr_2_15, d_cache_arr_2_14, d_cache_arr_2_13, 
      d_cache_arr_2_12, d_cache_arr_2_11, d_cache_arr_2_10, d_cache_arr_2_9, 
      d_cache_arr_2_8, d_cache_arr_2_7, d_cache_arr_2_6, d_cache_arr_2_5, 
      d_cache_arr_2_4, d_cache_arr_2_3, d_cache_arr_2_2, d_cache_arr_2_1, 
      d_cache_arr_2_0, d_cache_arr_3_31, d_cache_arr_3_30, d_cache_arr_3_29, 
      d_cache_arr_3_28, d_cache_arr_3_27, d_cache_arr_3_26, d_cache_arr_3_25, 
      d_cache_arr_3_24, d_cache_arr_3_23, d_cache_arr_3_22, d_cache_arr_3_21, 
      d_cache_arr_3_20, d_cache_arr_3_19, d_cache_arr_3_18, d_cache_arr_3_17, 
      d_cache_arr_3_16, d_cache_arr_3_15, d_cache_arr_3_14, d_cache_arr_3_13, 
      d_cache_arr_3_12, d_cache_arr_3_11, d_cache_arr_3_10, d_cache_arr_3_9, 
      d_cache_arr_3_8, d_cache_arr_3_7, d_cache_arr_3_6, d_cache_arr_3_5, 
      d_cache_arr_3_4, d_cache_arr_3_3, d_cache_arr_3_2, d_cache_arr_3_1, 
      d_cache_arr_3_0, d_cache_arr_4_31, d_cache_arr_4_30, d_cache_arr_4_29, 
      d_cache_arr_4_28, d_cache_arr_4_27, d_cache_arr_4_26, d_cache_arr_4_25, 
      d_cache_arr_4_24, d_cache_arr_4_23, d_cache_arr_4_22, d_cache_arr_4_21, 
      d_cache_arr_4_20, d_cache_arr_4_19, d_cache_arr_4_18, d_cache_arr_4_17, 
      d_cache_arr_4_16, d_cache_arr_4_15, d_cache_arr_4_14, d_cache_arr_4_13, 
      d_cache_arr_4_12, d_cache_arr_4_11, d_cache_arr_4_10, d_cache_arr_4_9, 
      d_cache_arr_4_8, d_cache_arr_4_7, d_cache_arr_4_6, d_cache_arr_4_5, 
      d_cache_arr_4_4, d_cache_arr_4_3, d_cache_arr_4_2, d_cache_arr_4_1, 
      d_cache_arr_4_0, d_cache_arr_5_31, d_cache_arr_5_30, d_cache_arr_5_29, 
      d_cache_arr_5_28, d_cache_arr_5_27, d_cache_arr_5_26, d_cache_arr_5_25, 
      d_cache_arr_5_24, d_cache_arr_5_23, d_cache_arr_5_22, d_cache_arr_5_21, 
      d_cache_arr_5_20, d_cache_arr_5_19, d_cache_arr_5_18, d_cache_arr_5_17, 
      d_cache_arr_5_16, d_cache_arr_5_15, d_cache_arr_5_14, d_cache_arr_5_13, 
      d_cache_arr_5_12, d_cache_arr_5_11, d_cache_arr_5_10, d_cache_arr_5_9, 
      d_cache_arr_5_8, d_cache_arr_5_7, d_cache_arr_5_6, d_cache_arr_5_5, 
      d_cache_arr_5_4, d_cache_arr_5_3, d_cache_arr_5_2, d_cache_arr_5_1, 
      d_cache_arr_5_0, d_cache_arr_6_31, d_cache_arr_6_30, d_cache_arr_6_29, 
      d_cache_arr_6_28, d_cache_arr_6_27, d_cache_arr_6_26, d_cache_arr_6_25, 
      d_cache_arr_6_24, d_cache_arr_6_23, d_cache_arr_6_22, d_cache_arr_6_21, 
      d_cache_arr_6_20, d_cache_arr_6_19, d_cache_arr_6_18, d_cache_arr_6_17, 
      d_cache_arr_6_16, d_cache_arr_6_15, d_cache_arr_6_14, d_cache_arr_6_13, 
      d_cache_arr_6_12, d_cache_arr_6_11, d_cache_arr_6_10, d_cache_arr_6_9, 
      d_cache_arr_6_8, d_cache_arr_6_7, d_cache_arr_6_6, d_cache_arr_6_5, 
      d_cache_arr_6_4, d_cache_arr_6_3, d_cache_arr_6_2, d_cache_arr_6_1, 
      d_cache_arr_6_0, d_cache_arr_7_31, d_cache_arr_7_30, d_cache_arr_7_29, 
      d_cache_arr_7_28, d_cache_arr_7_27, d_cache_arr_7_26, d_cache_arr_7_25, 
      d_cache_arr_7_24, d_cache_arr_7_23, d_cache_arr_7_22, d_cache_arr_7_21, 
      d_cache_arr_7_20, d_cache_arr_7_19, d_cache_arr_7_18, d_cache_arr_7_17, 
      d_cache_arr_7_16, d_cache_arr_7_15, d_cache_arr_7_14, d_cache_arr_7_13, 
      d_cache_arr_7_12, d_cache_arr_7_11, d_cache_arr_7_10, d_cache_arr_7_9, 
      d_cache_arr_7_8, d_cache_arr_7_7, d_cache_arr_7_6, d_cache_arr_7_5, 
      d_cache_arr_7_4, d_cache_arr_7_3, d_cache_arr_7_2, d_cache_arr_7_1, 
      d_cache_arr_7_0, d_cache_arr_8_31, d_cache_arr_8_30, d_cache_arr_8_29, 
      d_cache_arr_8_28, d_cache_arr_8_27, d_cache_arr_8_26, d_cache_arr_8_25, 
      d_cache_arr_8_24, d_cache_arr_8_23, d_cache_arr_8_22, d_cache_arr_8_21, 
      d_cache_arr_8_20, d_cache_arr_8_19, d_cache_arr_8_18, d_cache_arr_8_17, 
      d_cache_arr_8_16, d_cache_arr_8_15, d_cache_arr_8_14, d_cache_arr_8_13, 
      d_cache_arr_8_12, d_cache_arr_8_11, d_cache_arr_8_10, d_cache_arr_8_9, 
      d_cache_arr_8_8, d_cache_arr_8_7, d_cache_arr_8_6, d_cache_arr_8_5, 
      d_cache_arr_8_4, d_cache_arr_8_3, d_cache_arr_8_2, d_cache_arr_8_1, 
      d_cache_arr_8_0, d_cache_arr_9_31, d_cache_arr_9_30, d_cache_arr_9_29, 
      d_cache_arr_9_28, d_cache_arr_9_27, d_cache_arr_9_26, d_cache_arr_9_25, 
      d_cache_arr_9_24, d_cache_arr_9_23, d_cache_arr_9_22, d_cache_arr_9_21, 
      d_cache_arr_9_20, d_cache_arr_9_19, d_cache_arr_9_18, d_cache_arr_9_17, 
      d_cache_arr_9_16, d_cache_arr_9_15, d_cache_arr_9_14, d_cache_arr_9_13, 
      d_cache_arr_9_12, d_cache_arr_9_11, d_cache_arr_9_10, d_cache_arr_9_9, 
      d_cache_arr_9_8, d_cache_arr_9_7, d_cache_arr_9_6, d_cache_arr_9_5, 
      d_cache_arr_9_4, d_cache_arr_9_3, d_cache_arr_9_2, d_cache_arr_9_1, 
      d_cache_arr_9_0, d_cache_arr_10_31, d_cache_arr_10_30, 
      d_cache_arr_10_29, d_cache_arr_10_28, d_cache_arr_10_27, 
      d_cache_arr_10_26, d_cache_arr_10_25, d_cache_arr_10_24, 
      d_cache_arr_10_23, d_cache_arr_10_22, d_cache_arr_10_21, 
      d_cache_arr_10_20, d_cache_arr_10_19, d_cache_arr_10_18, 
      d_cache_arr_10_17, d_cache_arr_10_16, d_cache_arr_10_15, 
      d_cache_arr_10_14, d_cache_arr_10_13, d_cache_arr_10_12, 
      d_cache_arr_10_11, d_cache_arr_10_10, d_cache_arr_10_9, 
      d_cache_arr_10_8, d_cache_arr_10_7, d_cache_arr_10_6, d_cache_arr_10_5, 
      d_cache_arr_10_4, d_cache_arr_10_3, d_cache_arr_10_2, d_cache_arr_10_1, 
      d_cache_arr_10_0, d_cache_arr_11_31, d_cache_arr_11_30, 
      d_cache_arr_11_29, d_cache_arr_11_28, d_cache_arr_11_27, 
      d_cache_arr_11_26, d_cache_arr_11_25, d_cache_arr_11_24, 
      d_cache_arr_11_23, d_cache_arr_11_22, d_cache_arr_11_21, 
      d_cache_arr_11_20, d_cache_arr_11_19, d_cache_arr_11_18, 
      d_cache_arr_11_17, d_cache_arr_11_16, d_cache_arr_11_15, 
      d_cache_arr_11_14, d_cache_arr_11_13, d_cache_arr_11_12, 
      d_cache_arr_11_11, d_cache_arr_11_10, d_cache_arr_11_9, 
      d_cache_arr_11_8, d_cache_arr_11_7, d_cache_arr_11_6, d_cache_arr_11_5, 
      d_cache_arr_11_4, d_cache_arr_11_3, d_cache_arr_11_2, d_cache_arr_11_1, 
      d_cache_arr_11_0, d_cache_arr_12_31, d_cache_arr_12_30, 
      d_cache_arr_12_29, d_cache_arr_12_28, d_cache_arr_12_27, 
      d_cache_arr_12_26, d_cache_arr_12_25, d_cache_arr_12_24, 
      d_cache_arr_12_23, d_cache_arr_12_22, d_cache_arr_12_21, 
      d_cache_arr_12_20, d_cache_arr_12_19, d_cache_arr_12_18, 
      d_cache_arr_12_17, d_cache_arr_12_16, d_cache_arr_12_15, 
      d_cache_arr_12_14, d_cache_arr_12_13, d_cache_arr_12_12, 
      d_cache_arr_12_11, d_cache_arr_12_10, d_cache_arr_12_9, 
      d_cache_arr_12_8, d_cache_arr_12_7, d_cache_arr_12_6, d_cache_arr_12_5, 
      d_cache_arr_12_4, d_cache_arr_12_3, d_cache_arr_12_2, d_cache_arr_12_1, 
      d_cache_arr_12_0, d_cache_arr_13_31, d_cache_arr_13_30, 
      d_cache_arr_13_29, d_cache_arr_13_28, d_cache_arr_13_27, 
      d_cache_arr_13_26, d_cache_arr_13_25, d_cache_arr_13_24, 
      d_cache_arr_13_23, d_cache_arr_13_22, d_cache_arr_13_21, 
      d_cache_arr_13_20, d_cache_arr_13_19, d_cache_arr_13_18, 
      d_cache_arr_13_17, d_cache_arr_13_16, d_cache_arr_13_15, 
      d_cache_arr_13_14, d_cache_arr_13_13, d_cache_arr_13_12, 
      d_cache_arr_13_11, d_cache_arr_13_10, d_cache_arr_13_9, 
      d_cache_arr_13_8, d_cache_arr_13_7, d_cache_arr_13_6, d_cache_arr_13_5, 
      d_cache_arr_13_4, d_cache_arr_13_3, d_cache_arr_13_2, d_cache_arr_13_1, 
      d_cache_arr_13_0, d_cache_arr_14_31, d_cache_arr_14_30, 
      d_cache_arr_14_29, d_cache_arr_14_28, d_cache_arr_14_27, 
      d_cache_arr_14_26, d_cache_arr_14_25, d_cache_arr_14_24, 
      d_cache_arr_14_23, d_cache_arr_14_22, d_cache_arr_14_21, 
      d_cache_arr_14_20, d_cache_arr_14_19, d_cache_arr_14_18, 
      d_cache_arr_14_17, d_cache_arr_14_16, d_cache_arr_14_15, 
      d_cache_arr_14_14, d_cache_arr_14_13, d_cache_arr_14_12, 
      d_cache_arr_14_11, d_cache_arr_14_10, d_cache_arr_14_9, 
      d_cache_arr_14_8, d_cache_arr_14_7, d_cache_arr_14_6, d_cache_arr_14_5, 
      d_cache_arr_14_4, d_cache_arr_14_3, d_cache_arr_14_2, d_cache_arr_14_1, 
      d_cache_arr_14_0, d_cache_arr_15_31, d_cache_arr_15_30, 
      d_cache_arr_15_29, d_cache_arr_15_28, d_cache_arr_15_27, 
      d_cache_arr_15_26, d_cache_arr_15_25, d_cache_arr_15_24, 
      d_cache_arr_15_23, d_cache_arr_15_22, d_cache_arr_15_21, 
      d_cache_arr_15_20, d_cache_arr_15_19, d_cache_arr_15_18, 
      d_cache_arr_15_17, d_cache_arr_15_16, d_cache_arr_15_15, 
      d_cache_arr_15_14, d_cache_arr_15_13, d_cache_arr_15_12, 
      d_cache_arr_15_11, d_cache_arr_15_10, d_cache_arr_15_9, 
      d_cache_arr_15_8, d_cache_arr_15_7, d_cache_arr_15_6, d_cache_arr_15_5, 
      d_cache_arr_15_4, d_cache_arr_15_3, d_cache_arr_15_2, d_cache_arr_15_1, 
      d_cache_arr_15_0, d_cache_arr_16_31, d_cache_arr_16_30, 
      d_cache_arr_16_29, d_cache_arr_16_28, d_cache_arr_16_27, 
      d_cache_arr_16_26, d_cache_arr_16_25, d_cache_arr_16_24, 
      d_cache_arr_16_23, d_cache_arr_16_22, d_cache_arr_16_21, 
      d_cache_arr_16_20, d_cache_arr_16_19, d_cache_arr_16_18, 
      d_cache_arr_16_17, d_cache_arr_16_16, d_cache_arr_16_15, 
      d_cache_arr_16_14, d_cache_arr_16_13, d_cache_arr_16_12, 
      d_cache_arr_16_11, d_cache_arr_16_10, d_cache_arr_16_9, 
      d_cache_arr_16_8, d_cache_arr_16_7, d_cache_arr_16_6, d_cache_arr_16_5, 
      d_cache_arr_16_4, d_cache_arr_16_3, d_cache_arr_16_2, d_cache_arr_16_1, 
      d_cache_arr_16_0, d_cache_arr_17_31, d_cache_arr_17_30, 
      d_cache_arr_17_29, d_cache_arr_17_28, d_cache_arr_17_27, 
      d_cache_arr_17_26, d_cache_arr_17_25, d_cache_arr_17_24, 
      d_cache_arr_17_23, d_cache_arr_17_22, d_cache_arr_17_21, 
      d_cache_arr_17_20, d_cache_arr_17_19, d_cache_arr_17_18, 
      d_cache_arr_17_17, d_cache_arr_17_16, d_cache_arr_17_15, 
      d_cache_arr_17_14, d_cache_arr_17_13, d_cache_arr_17_12, 
      d_cache_arr_17_11, d_cache_arr_17_10, d_cache_arr_17_9, 
      d_cache_arr_17_8, d_cache_arr_17_7, d_cache_arr_17_6, d_cache_arr_17_5, 
      d_cache_arr_17_4, d_cache_arr_17_3, d_cache_arr_17_2, d_cache_arr_17_1, 
      d_cache_arr_17_0, d_cache_arr_18_31, d_cache_arr_18_30, 
      d_cache_arr_18_29, d_cache_arr_18_28, d_cache_arr_18_27, 
      d_cache_arr_18_26, d_cache_arr_18_25, d_cache_arr_18_24, 
      d_cache_arr_18_23, d_cache_arr_18_22, d_cache_arr_18_21, 
      d_cache_arr_18_20, d_cache_arr_18_19, d_cache_arr_18_18, 
      d_cache_arr_18_17, d_cache_arr_18_16, d_cache_arr_18_15, 
      d_cache_arr_18_14, d_cache_arr_18_13, d_cache_arr_18_12, 
      d_cache_arr_18_11, d_cache_arr_18_10, d_cache_arr_18_9, 
      d_cache_arr_18_8, d_cache_arr_18_7, d_cache_arr_18_6, d_cache_arr_18_5, 
      d_cache_arr_18_4, d_cache_arr_18_3, d_cache_arr_18_2, d_cache_arr_18_1, 
      d_cache_arr_18_0, d_cache_arr_19_31, d_cache_arr_19_30, 
      d_cache_arr_19_29, d_cache_arr_19_28, d_cache_arr_19_27, 
      d_cache_arr_19_26, d_cache_arr_19_25, d_cache_arr_19_24, 
      d_cache_arr_19_23, d_cache_arr_19_22, d_cache_arr_19_21, 
      d_cache_arr_19_20, d_cache_arr_19_19, d_cache_arr_19_18, 
      d_cache_arr_19_17, d_cache_arr_19_16, d_cache_arr_19_15, 
      d_cache_arr_19_14, d_cache_arr_19_13, d_cache_arr_19_12, 
      d_cache_arr_19_11, d_cache_arr_19_10, d_cache_arr_19_9, 
      d_cache_arr_19_8, d_cache_arr_19_7, d_cache_arr_19_6, d_cache_arr_19_5, 
      d_cache_arr_19_4, d_cache_arr_19_3, d_cache_arr_19_2, d_cache_arr_19_1, 
      d_cache_arr_19_0, d_cache_arr_20_31, d_cache_arr_20_30, 
      d_cache_arr_20_29, d_cache_arr_20_28, d_cache_arr_20_27, 
      d_cache_arr_20_26, d_cache_arr_20_25, d_cache_arr_20_24, 
      d_cache_arr_20_23, d_cache_arr_20_22, d_cache_arr_20_21, 
      d_cache_arr_20_20, d_cache_arr_20_19, d_cache_arr_20_18, 
      d_cache_arr_20_17, d_cache_arr_20_16, d_cache_arr_20_15, 
      d_cache_arr_20_14, d_cache_arr_20_13, d_cache_arr_20_12, 
      d_cache_arr_20_11, d_cache_arr_20_10, d_cache_arr_20_9, 
      d_cache_arr_20_8, d_cache_arr_20_7, d_cache_arr_20_6, d_cache_arr_20_5, 
      d_cache_arr_20_4, d_cache_arr_20_3, d_cache_arr_20_2, d_cache_arr_20_1, 
      d_cache_arr_20_0, d_cache_arr_21_31, d_cache_arr_21_30, 
      d_cache_arr_21_29, d_cache_arr_21_28, d_cache_arr_21_27, 
      d_cache_arr_21_26, d_cache_arr_21_25, d_cache_arr_21_24, 
      d_cache_arr_21_23, d_cache_arr_21_22, d_cache_arr_21_21, 
      d_cache_arr_21_20, d_cache_arr_21_19, d_cache_arr_21_18, 
      d_cache_arr_21_17, d_cache_arr_21_16, d_cache_arr_21_15, 
      d_cache_arr_21_14, d_cache_arr_21_13, d_cache_arr_21_12, 
      d_cache_arr_21_11, d_cache_arr_21_10, d_cache_arr_21_9, 
      d_cache_arr_21_8, d_cache_arr_21_7, d_cache_arr_21_6, d_cache_arr_21_5, 
      d_cache_arr_21_4, d_cache_arr_21_3, d_cache_arr_21_2, d_cache_arr_21_1, 
      d_cache_arr_21_0, d_cache_arr_22_31, d_cache_arr_22_30, 
      d_cache_arr_22_29, d_cache_arr_22_28, d_cache_arr_22_27, 
      d_cache_arr_22_26, d_cache_arr_22_25, d_cache_arr_22_24, 
      d_cache_arr_22_23, d_cache_arr_22_22, d_cache_arr_22_21, 
      d_cache_arr_22_20, d_cache_arr_22_19, d_cache_arr_22_18, 
      d_cache_arr_22_17, d_cache_arr_22_16, d_cache_arr_22_15, 
      d_cache_arr_22_14, d_cache_arr_22_13, d_cache_arr_22_12, 
      d_cache_arr_22_11, d_cache_arr_22_10, d_cache_arr_22_9, 
      d_cache_arr_22_8, d_cache_arr_22_7, d_cache_arr_22_6, d_cache_arr_22_5, 
      d_cache_arr_22_4, d_cache_arr_22_3, d_cache_arr_22_2, d_cache_arr_22_1, 
      d_cache_arr_22_0, d_cache_arr_23_31, d_cache_arr_23_30, 
      d_cache_arr_23_29, d_cache_arr_23_28, d_cache_arr_23_27, 
      d_cache_arr_23_26, d_cache_arr_23_25, d_cache_arr_23_24, 
      d_cache_arr_23_23, d_cache_arr_23_22, d_cache_arr_23_21, 
      d_cache_arr_23_20, d_cache_arr_23_19, d_cache_arr_23_18, 
      d_cache_arr_23_17, d_cache_arr_23_16, d_cache_arr_23_15, 
      d_cache_arr_23_14, d_cache_arr_23_13, d_cache_arr_23_12, 
      d_cache_arr_23_11, d_cache_arr_23_10, d_cache_arr_23_9, 
      d_cache_arr_23_8, d_cache_arr_23_7, d_cache_arr_23_6, d_cache_arr_23_5, 
      d_cache_arr_23_4, d_cache_arr_23_3, d_cache_arr_23_2, d_cache_arr_23_1, 
      d_cache_arr_23_0, d_cache_arr_24_31, d_cache_arr_24_30, 
      d_cache_arr_24_29, d_cache_arr_24_28, d_cache_arr_24_27, 
      d_cache_arr_24_26, d_cache_arr_24_25, d_cache_arr_24_24, 
      d_cache_arr_24_23, d_cache_arr_24_22, d_cache_arr_24_21, 
      d_cache_arr_24_20, d_cache_arr_24_19, d_cache_arr_24_18, 
      d_cache_arr_24_17, d_cache_arr_24_16, d_cache_arr_24_15, 
      d_cache_arr_24_14, d_cache_arr_24_13, d_cache_arr_24_12, 
      d_cache_arr_24_11, d_cache_arr_24_10, d_cache_arr_24_9, 
      d_cache_arr_24_8, d_cache_arr_24_7, d_cache_arr_24_6, d_cache_arr_24_5, 
      d_cache_arr_24_4, d_cache_arr_24_3, d_cache_arr_24_2, d_cache_arr_24_1, 
      d_cache_arr_24_0, q_cache_arr_0_31, q_cache_arr_0_30, q_cache_arr_0_29, 
      q_cache_arr_0_28, q_cache_arr_0_27, q_cache_arr_0_26, q_cache_arr_0_25, 
      q_cache_arr_0_24, q_cache_arr_0_23, q_cache_arr_0_22, q_cache_arr_0_21, 
      q_cache_arr_0_20, q_cache_arr_0_19, q_cache_arr_0_18, q_cache_arr_0_17, 
      q_cache_arr_0_16, q_cache_arr_0_15, q_cache_arr_0_14, q_cache_arr_0_13, 
      q_cache_arr_0_12, q_cache_arr_0_11, q_cache_arr_0_10, q_cache_arr_0_9, 
      q_cache_arr_0_8, q_cache_arr_0_7, q_cache_arr_0_6, q_cache_arr_0_5, 
      q_cache_arr_0_4, q_cache_arr_0_3, q_cache_arr_0_2, q_cache_arr_0_1, 
      q_cache_arr_0_0, q_cache_arr_1_31, q_cache_arr_1_30, q_cache_arr_1_29, 
      q_cache_arr_1_28, q_cache_arr_1_27, q_cache_arr_1_26, q_cache_arr_1_25, 
      q_cache_arr_1_24, q_cache_arr_1_23, q_cache_arr_1_22, q_cache_arr_1_21, 
      q_cache_arr_1_20, q_cache_arr_1_19, q_cache_arr_1_18, q_cache_arr_1_17, 
      q_cache_arr_1_16, q_cache_arr_1_15, q_cache_arr_1_14, q_cache_arr_1_13, 
      q_cache_arr_1_12, q_cache_arr_1_11, q_cache_arr_1_10, q_cache_arr_1_9, 
      q_cache_arr_1_8, q_cache_arr_1_7, q_cache_arr_1_6, q_cache_arr_1_5, 
      q_cache_arr_1_4, q_cache_arr_1_3, q_cache_arr_1_2, q_cache_arr_1_1, 
      q_cache_arr_1_0, q_cache_arr_2_31, q_cache_arr_2_30, q_cache_arr_2_29, 
      q_cache_arr_2_28, q_cache_arr_2_27, q_cache_arr_2_26, q_cache_arr_2_25, 
      q_cache_arr_2_24, q_cache_arr_2_23, q_cache_arr_2_22, q_cache_arr_2_21, 
      q_cache_arr_2_20, q_cache_arr_2_19, q_cache_arr_2_18, q_cache_arr_2_17, 
      q_cache_arr_2_16, q_cache_arr_2_15, q_cache_arr_2_14, q_cache_arr_2_13, 
      q_cache_arr_2_12, q_cache_arr_2_11, q_cache_arr_2_10, q_cache_arr_2_9, 
      q_cache_arr_2_8, q_cache_arr_2_7, q_cache_arr_2_6, q_cache_arr_2_5, 
      q_cache_arr_2_4, q_cache_arr_2_3, q_cache_arr_2_2, q_cache_arr_2_1, 
      q_cache_arr_2_0, q_cache_arr_3_31, q_cache_arr_3_30, q_cache_arr_3_29, 
      q_cache_arr_3_28, q_cache_arr_3_27, q_cache_arr_3_26, q_cache_arr_3_25, 
      q_cache_arr_3_24, q_cache_arr_3_23, q_cache_arr_3_22, q_cache_arr_3_21, 
      q_cache_arr_3_20, q_cache_arr_3_19, q_cache_arr_3_18, q_cache_arr_3_17, 
      q_cache_arr_3_16, q_cache_arr_3_15, q_cache_arr_3_14, q_cache_arr_3_13, 
      q_cache_arr_3_12, q_cache_arr_3_11, q_cache_arr_3_10, q_cache_arr_3_9, 
      q_cache_arr_3_8, q_cache_arr_3_7, q_cache_arr_3_6, q_cache_arr_3_5, 
      q_cache_arr_3_4, q_cache_arr_3_3, q_cache_arr_3_2, q_cache_arr_3_1, 
      q_cache_arr_3_0, q_cache_arr_4_31, q_cache_arr_4_30, q_cache_arr_4_29, 
      q_cache_arr_4_28, q_cache_arr_4_27, q_cache_arr_4_26, q_cache_arr_4_25, 
      q_cache_arr_4_24, q_cache_arr_4_23, q_cache_arr_4_22, q_cache_arr_4_21, 
      q_cache_arr_4_20, q_cache_arr_4_19, q_cache_arr_4_18, q_cache_arr_4_17, 
      q_cache_arr_4_16, q_cache_arr_4_15, q_cache_arr_4_14, q_cache_arr_4_13, 
      q_cache_arr_4_12, q_cache_arr_4_11, q_cache_arr_4_10, q_cache_arr_4_9, 
      q_cache_arr_4_8, q_cache_arr_4_7, q_cache_arr_4_6, q_cache_arr_4_5, 
      q_cache_arr_4_4, q_cache_arr_4_3, q_cache_arr_4_2, q_cache_arr_4_1, 
      q_cache_arr_4_0, q_cache_arr_5_31, q_cache_arr_5_30, q_cache_arr_5_29, 
      q_cache_arr_5_28, q_cache_arr_5_27, q_cache_arr_5_26, q_cache_arr_5_25, 
      q_cache_arr_5_24, q_cache_arr_5_23, q_cache_arr_5_22, q_cache_arr_5_21, 
      q_cache_arr_5_20, q_cache_arr_5_19, q_cache_arr_5_18, q_cache_arr_5_17, 
      q_cache_arr_5_16, q_cache_arr_5_15, q_cache_arr_5_14, q_cache_arr_5_13, 
      q_cache_arr_5_12, q_cache_arr_5_11, q_cache_arr_5_10, q_cache_arr_5_9, 
      q_cache_arr_5_8, q_cache_arr_5_7, q_cache_arr_5_6, q_cache_arr_5_5, 
      q_cache_arr_5_4, q_cache_arr_5_3, q_cache_arr_5_2, q_cache_arr_5_1, 
      q_cache_arr_5_0, q_cache_arr_6_31, q_cache_arr_6_30, q_cache_arr_6_29, 
      q_cache_arr_6_28, q_cache_arr_6_27, q_cache_arr_6_26, q_cache_arr_6_25, 
      q_cache_arr_6_24, q_cache_arr_6_23, q_cache_arr_6_22, q_cache_arr_6_21, 
      q_cache_arr_6_20, q_cache_arr_6_19, q_cache_arr_6_18, q_cache_arr_6_17, 
      q_cache_arr_6_16, q_cache_arr_6_15, q_cache_arr_6_14, q_cache_arr_6_13, 
      q_cache_arr_6_12, q_cache_arr_6_11, q_cache_arr_6_10, q_cache_arr_6_9, 
      q_cache_arr_6_8, q_cache_arr_6_7, q_cache_arr_6_6, q_cache_arr_6_5, 
      q_cache_arr_6_4, q_cache_arr_6_3, q_cache_arr_6_2, q_cache_arr_6_1, 
      q_cache_arr_6_0, q_cache_arr_7_31, q_cache_arr_7_30, q_cache_arr_7_29, 
      q_cache_arr_7_28, q_cache_arr_7_27, q_cache_arr_7_26, q_cache_arr_7_25, 
      q_cache_arr_7_24, q_cache_arr_7_23, q_cache_arr_7_22, q_cache_arr_7_21, 
      q_cache_arr_7_20, q_cache_arr_7_19, q_cache_arr_7_18, q_cache_arr_7_17, 
      q_cache_arr_7_16, q_cache_arr_7_15, q_cache_arr_7_14, q_cache_arr_7_13, 
      q_cache_arr_7_12, q_cache_arr_7_11, q_cache_arr_7_10, q_cache_arr_7_9, 
      q_cache_arr_7_8, q_cache_arr_7_7, q_cache_arr_7_6, q_cache_arr_7_5, 
      q_cache_arr_7_4, q_cache_arr_7_3, q_cache_arr_7_2, q_cache_arr_7_1, 
      q_cache_arr_7_0, q_cache_arr_8_31, q_cache_arr_8_30, q_cache_arr_8_29, 
      q_cache_arr_8_28, q_cache_arr_8_27, q_cache_arr_8_26, q_cache_arr_8_25, 
      q_cache_arr_8_24, q_cache_arr_8_23, q_cache_arr_8_22, q_cache_arr_8_21, 
      q_cache_arr_8_20, q_cache_arr_8_19, q_cache_arr_8_18, q_cache_arr_8_17, 
      q_cache_arr_8_16, q_cache_arr_8_15, q_cache_arr_8_14, q_cache_arr_8_13, 
      q_cache_arr_8_12, q_cache_arr_8_11, q_cache_arr_8_10, q_cache_arr_8_9, 
      q_cache_arr_8_8, q_cache_arr_8_7, q_cache_arr_8_6, q_cache_arr_8_5, 
      q_cache_arr_8_4, q_cache_arr_8_3, q_cache_arr_8_2, q_cache_arr_8_1, 
      q_cache_arr_8_0, q_cache_arr_9_31, q_cache_arr_9_30, q_cache_arr_9_29, 
      q_cache_arr_9_28, q_cache_arr_9_27, q_cache_arr_9_26, q_cache_arr_9_25, 
      q_cache_arr_9_24, q_cache_arr_9_23, q_cache_arr_9_22, q_cache_arr_9_21, 
      q_cache_arr_9_20, q_cache_arr_9_19, q_cache_arr_9_18, q_cache_arr_9_17, 
      q_cache_arr_9_16, q_cache_arr_9_15, q_cache_arr_9_14, q_cache_arr_9_13, 
      q_cache_arr_9_12, q_cache_arr_9_11, q_cache_arr_9_10, q_cache_arr_9_9, 
      q_cache_arr_9_8, q_cache_arr_9_7, q_cache_arr_9_6, q_cache_arr_9_5, 
      q_cache_arr_9_4, q_cache_arr_9_3, q_cache_arr_9_2, q_cache_arr_9_1, 
      q_cache_arr_9_0, q_cache_arr_10_31, q_cache_arr_10_30, 
      q_cache_arr_10_29, q_cache_arr_10_28, q_cache_arr_10_27, 
      q_cache_arr_10_26, q_cache_arr_10_25, q_cache_arr_10_24, 
      q_cache_arr_10_23, q_cache_arr_10_22, q_cache_arr_10_21, 
      q_cache_arr_10_20, q_cache_arr_10_19, q_cache_arr_10_18, 
      q_cache_arr_10_17, q_cache_arr_10_16, q_cache_arr_10_15, 
      q_cache_arr_10_14, q_cache_arr_10_13, q_cache_arr_10_12, 
      q_cache_arr_10_11, q_cache_arr_10_10, q_cache_arr_10_9, 
      q_cache_arr_10_8, q_cache_arr_10_7, q_cache_arr_10_6, q_cache_arr_10_5, 
      q_cache_arr_10_4, q_cache_arr_10_3, q_cache_arr_10_2, q_cache_arr_10_1, 
      q_cache_arr_10_0, q_cache_arr_11_31, q_cache_arr_11_30, 
      q_cache_arr_11_29, q_cache_arr_11_28, q_cache_arr_11_27, 
      q_cache_arr_11_26, q_cache_arr_11_25, q_cache_arr_11_24, 
      q_cache_arr_11_23, q_cache_arr_11_22, q_cache_arr_11_21, 
      q_cache_arr_11_20, q_cache_arr_11_19, q_cache_arr_11_18, 
      q_cache_arr_11_17, q_cache_arr_11_16, q_cache_arr_11_15, 
      q_cache_arr_11_14, q_cache_arr_11_13, q_cache_arr_11_12, 
      q_cache_arr_11_11, q_cache_arr_11_10, q_cache_arr_11_9, 
      q_cache_arr_11_8, q_cache_arr_11_7, q_cache_arr_11_6, q_cache_arr_11_5, 
      q_cache_arr_11_4, q_cache_arr_11_3, q_cache_arr_11_2, q_cache_arr_11_1, 
      q_cache_arr_11_0, q_cache_arr_12_31, q_cache_arr_12_30, 
      q_cache_arr_12_29, q_cache_arr_12_28, q_cache_arr_12_27, 
      q_cache_arr_12_26, q_cache_arr_12_25, q_cache_arr_12_24, 
      q_cache_arr_12_23, q_cache_arr_12_22, q_cache_arr_12_21, 
      q_cache_arr_12_20, q_cache_arr_12_19, q_cache_arr_12_18, 
      q_cache_arr_12_17, q_cache_arr_12_16, q_cache_arr_12_15, 
      q_cache_arr_12_14, q_cache_arr_12_13, q_cache_arr_12_12, 
      q_cache_arr_12_11, q_cache_arr_12_10, q_cache_arr_12_9, 
      q_cache_arr_12_8, q_cache_arr_12_7, q_cache_arr_12_6, q_cache_arr_12_5, 
      q_cache_arr_12_4, q_cache_arr_12_3, q_cache_arr_12_2, q_cache_arr_12_1, 
      q_cache_arr_12_0, q_cache_arr_13_31, q_cache_arr_13_30, 
      q_cache_arr_13_29, q_cache_arr_13_28, q_cache_arr_13_27, 
      q_cache_arr_13_26, q_cache_arr_13_25, q_cache_arr_13_24, 
      q_cache_arr_13_23, q_cache_arr_13_22, q_cache_arr_13_21, 
      q_cache_arr_13_20, q_cache_arr_13_19, q_cache_arr_13_18, 
      q_cache_arr_13_17, q_cache_arr_13_16, q_cache_arr_13_15, 
      q_cache_arr_13_14, q_cache_arr_13_13, q_cache_arr_13_12, 
      q_cache_arr_13_11, q_cache_arr_13_10, q_cache_arr_13_9, 
      q_cache_arr_13_8, q_cache_arr_13_7, q_cache_arr_13_6, q_cache_arr_13_5, 
      q_cache_arr_13_4, q_cache_arr_13_3, q_cache_arr_13_2, q_cache_arr_13_1, 
      q_cache_arr_13_0, q_cache_arr_14_31, q_cache_arr_14_30, 
      q_cache_arr_14_29, q_cache_arr_14_28, q_cache_arr_14_27, 
      q_cache_arr_14_26, q_cache_arr_14_25, q_cache_arr_14_24, 
      q_cache_arr_14_23, q_cache_arr_14_22, q_cache_arr_14_21, 
      q_cache_arr_14_20, q_cache_arr_14_19, q_cache_arr_14_18, 
      q_cache_arr_14_17, q_cache_arr_14_16, q_cache_arr_14_15, 
      q_cache_arr_14_14, q_cache_arr_14_13, q_cache_arr_14_12, 
      q_cache_arr_14_11, q_cache_arr_14_10, q_cache_arr_14_9, 
      q_cache_arr_14_8, q_cache_arr_14_7, q_cache_arr_14_6, q_cache_arr_14_5, 
      q_cache_arr_14_4, q_cache_arr_14_3, q_cache_arr_14_2, q_cache_arr_14_1, 
      q_cache_arr_14_0, q_cache_arr_15_31, q_cache_arr_15_30, 
      q_cache_arr_15_29, q_cache_arr_15_28, q_cache_arr_15_27, 
      q_cache_arr_15_26, q_cache_arr_15_25, q_cache_arr_15_24, 
      q_cache_arr_15_23, q_cache_arr_15_22, q_cache_arr_15_21, 
      q_cache_arr_15_20, q_cache_arr_15_19, q_cache_arr_15_18, 
      q_cache_arr_15_17, q_cache_arr_15_16, q_cache_arr_15_15, 
      q_cache_arr_15_14, q_cache_arr_15_13, q_cache_arr_15_12, 
      q_cache_arr_15_11, q_cache_arr_15_10, q_cache_arr_15_9, 
      q_cache_arr_15_8, q_cache_arr_15_7, q_cache_arr_15_6, q_cache_arr_15_5, 
      q_cache_arr_15_4, q_cache_arr_15_3, q_cache_arr_15_2, q_cache_arr_15_1, 
      q_cache_arr_15_0, q_cache_arr_16_31, q_cache_arr_16_30, 
      q_cache_arr_16_29, q_cache_arr_16_28, q_cache_arr_16_27, 
      q_cache_arr_16_26, q_cache_arr_16_25, q_cache_arr_16_24, 
      q_cache_arr_16_23, q_cache_arr_16_22, q_cache_arr_16_21, 
      q_cache_arr_16_20, q_cache_arr_16_19, q_cache_arr_16_18, 
      q_cache_arr_16_17, q_cache_arr_16_16, q_cache_arr_16_15, 
      q_cache_arr_16_14, q_cache_arr_16_13, q_cache_arr_16_12, 
      q_cache_arr_16_11, q_cache_arr_16_10, q_cache_arr_16_9, 
      q_cache_arr_16_8, q_cache_arr_16_7, q_cache_arr_16_6, q_cache_arr_16_5, 
      q_cache_arr_16_4, q_cache_arr_16_3, q_cache_arr_16_2, q_cache_arr_16_1, 
      q_cache_arr_16_0, q_cache_arr_17_31, q_cache_arr_17_30, 
      q_cache_arr_17_29, q_cache_arr_17_28, q_cache_arr_17_27, 
      q_cache_arr_17_26, q_cache_arr_17_25, q_cache_arr_17_24, 
      q_cache_arr_17_23, q_cache_arr_17_22, q_cache_arr_17_21, 
      q_cache_arr_17_20, q_cache_arr_17_19, q_cache_arr_17_18, 
      q_cache_arr_17_17, q_cache_arr_17_16, q_cache_arr_17_15, 
      q_cache_arr_17_14, q_cache_arr_17_13, q_cache_arr_17_12, 
      q_cache_arr_17_11, q_cache_arr_17_10, q_cache_arr_17_9, 
      q_cache_arr_17_8, q_cache_arr_17_7, q_cache_arr_17_6, q_cache_arr_17_5, 
      q_cache_arr_17_4, q_cache_arr_17_3, q_cache_arr_17_2, q_cache_arr_17_1, 
      q_cache_arr_17_0, q_cache_arr_18_31, q_cache_arr_18_30, 
      q_cache_arr_18_29, q_cache_arr_18_28, q_cache_arr_18_27, 
      q_cache_arr_18_26, q_cache_arr_18_25, q_cache_arr_18_24, 
      q_cache_arr_18_23, q_cache_arr_18_22, q_cache_arr_18_21, 
      q_cache_arr_18_20, q_cache_arr_18_19, q_cache_arr_18_18, 
      q_cache_arr_18_17, q_cache_arr_18_16, q_cache_arr_18_15, 
      q_cache_arr_18_14, q_cache_arr_18_13, q_cache_arr_18_12, 
      q_cache_arr_18_11, q_cache_arr_18_10, q_cache_arr_18_9, 
      q_cache_arr_18_8, q_cache_arr_18_7, q_cache_arr_18_6, q_cache_arr_18_5, 
      q_cache_arr_18_4, q_cache_arr_18_3, q_cache_arr_18_2, q_cache_arr_18_1, 
      q_cache_arr_18_0, q_cache_arr_19_31, q_cache_arr_19_30, 
      q_cache_arr_19_29, q_cache_arr_19_28, q_cache_arr_19_27, 
      q_cache_arr_19_26, q_cache_arr_19_25, q_cache_arr_19_24, 
      q_cache_arr_19_23, q_cache_arr_19_22, q_cache_arr_19_21, 
      q_cache_arr_19_20, q_cache_arr_19_19, q_cache_arr_19_18, 
      q_cache_arr_19_17, q_cache_arr_19_16, q_cache_arr_19_15, 
      q_cache_arr_19_14, q_cache_arr_19_13, q_cache_arr_19_12, 
      q_cache_arr_19_11, q_cache_arr_19_10, q_cache_arr_19_9, 
      q_cache_arr_19_8, q_cache_arr_19_7, q_cache_arr_19_6, q_cache_arr_19_5, 
      q_cache_arr_19_4, q_cache_arr_19_3, q_cache_arr_19_2, q_cache_arr_19_1, 
      q_cache_arr_19_0, q_cache_arr_20_31, q_cache_arr_20_30, 
      q_cache_arr_20_29, q_cache_arr_20_28, q_cache_arr_20_27, 
      q_cache_arr_20_26, q_cache_arr_20_25, q_cache_arr_20_24, 
      q_cache_arr_20_23, q_cache_arr_20_22, q_cache_arr_20_21, 
      q_cache_arr_20_20, q_cache_arr_20_19, q_cache_arr_20_18, 
      q_cache_arr_20_17, q_cache_arr_20_16, q_cache_arr_20_15, 
      q_cache_arr_20_14, q_cache_arr_20_13, q_cache_arr_20_12, 
      q_cache_arr_20_11, q_cache_arr_20_10, q_cache_arr_20_9, 
      q_cache_arr_20_8, q_cache_arr_20_7, q_cache_arr_20_6, q_cache_arr_20_5, 
      q_cache_arr_20_4, q_cache_arr_20_3, q_cache_arr_20_2, q_cache_arr_20_1, 
      q_cache_arr_20_0, q_cache_arr_21_31, q_cache_arr_21_30, 
      q_cache_arr_21_29, q_cache_arr_21_28, q_cache_arr_21_27, 
      q_cache_arr_21_26, q_cache_arr_21_25, q_cache_arr_21_24, 
      q_cache_arr_21_23, q_cache_arr_21_22, q_cache_arr_21_21, 
      q_cache_arr_21_20, q_cache_arr_21_19, q_cache_arr_21_18, 
      q_cache_arr_21_17, q_cache_arr_21_16, q_cache_arr_21_15, 
      q_cache_arr_21_14, q_cache_arr_21_13, q_cache_arr_21_12, 
      q_cache_arr_21_11, q_cache_arr_21_10, q_cache_arr_21_9, 
      q_cache_arr_21_8, q_cache_arr_21_7, q_cache_arr_21_6, q_cache_arr_21_5, 
      q_cache_arr_21_4, q_cache_arr_21_3, q_cache_arr_21_2, q_cache_arr_21_1, 
      q_cache_arr_21_0, q_cache_arr_22_31, q_cache_arr_22_30, 
      q_cache_arr_22_29, q_cache_arr_22_28, q_cache_arr_22_27, 
      q_cache_arr_22_26, q_cache_arr_22_25, q_cache_arr_22_24, 
      q_cache_arr_22_23, q_cache_arr_22_22, q_cache_arr_22_21, 
      q_cache_arr_22_20, q_cache_arr_22_19, q_cache_arr_22_18, 
      q_cache_arr_22_17, q_cache_arr_22_16, q_cache_arr_22_15, 
      q_cache_arr_22_14, q_cache_arr_22_13, q_cache_arr_22_12, 
      q_cache_arr_22_11, q_cache_arr_22_10, q_cache_arr_22_9, 
      q_cache_arr_22_8, q_cache_arr_22_7, q_cache_arr_22_6, q_cache_arr_22_5, 
      q_cache_arr_22_4, q_cache_arr_22_3, q_cache_arr_22_2, q_cache_arr_22_1, 
      q_cache_arr_22_0, q_cache_arr_23_31, q_cache_arr_23_30, 
      q_cache_arr_23_29, q_cache_arr_23_28, q_cache_arr_23_27, 
      q_cache_arr_23_26, q_cache_arr_23_25, q_cache_arr_23_24, 
      q_cache_arr_23_23, q_cache_arr_23_22, q_cache_arr_23_21, 
      q_cache_arr_23_20, q_cache_arr_23_19, q_cache_arr_23_18, 
      q_cache_arr_23_17, q_cache_arr_23_16, q_cache_arr_23_15, 
      q_cache_arr_23_14, q_cache_arr_23_13, q_cache_arr_23_12, 
      q_cache_arr_23_11, q_cache_arr_23_10, q_cache_arr_23_9, 
      q_cache_arr_23_8, q_cache_arr_23_7, q_cache_arr_23_6, q_cache_arr_23_5, 
      q_cache_arr_23_4, q_cache_arr_23_3, q_cache_arr_23_2, q_cache_arr_23_1, 
      q_cache_arr_23_0, q_cache_arr_24_31, q_cache_arr_24_30, 
      q_cache_arr_24_29, q_cache_arr_24_28, q_cache_arr_24_27, 
      q_cache_arr_24_26, q_cache_arr_24_25, q_cache_arr_24_24, 
      q_cache_arr_24_23, q_cache_arr_24_22, q_cache_arr_24_21, 
      q_cache_arr_24_20, q_cache_arr_24_19, q_cache_arr_24_18, 
      q_cache_arr_24_17, q_cache_arr_24_16, q_cache_arr_24_15, 
      q_cache_arr_24_14, q_cache_arr_24_13, q_cache_arr_24_12, 
      q_cache_arr_24_11, q_cache_arr_24_10, q_cache_arr_24_9, 
      q_cache_arr_24_8, q_cache_arr_24_7, q_cache_arr_24_6, q_cache_arr_24_5, 
      q_cache_arr_24_4, q_cache_arr_24_3, q_cache_arr_24_2, q_cache_arr_24_1, 
      q_cache_arr_24_0, img_load_tmp, filter_load_tmp, ready_tmp, 
      buffer_ready_tmp, comp_pipe_rst, comp_pipe_en, output1_init_q_15, 
      output1_init_q_14, output1_init_q_13, output1_init_q_12, 
      output1_init_q_11, output1_init_q_10, output1_init_q_9, 
      output1_init_q_8, output1_init_q_7, output1_init_q_6, output1_init_q_5, 
      output1_init_q_4, output1_init_q_3, output1_init_q_2, output1_init_q_1, 
      output1_init_q_0, output2_init_q_15, output2_init_q_14, 
      output2_init_q_13, output2_init_q_12, output2_init_q_11, 
      output2_init_q_10, output2_init_q_9, output2_init_q_8, 
      output2_init_q_7, output2_init_q_6, output2_init_q_5, output2_init_q_4, 
      output2_init_q_3, output2_init_q_2, output2_init_q_1, output2_init_q_0, 
      filter_size_q, operation_q, compute_relu_q, semi_ready, 
      buffer_ready_EXMPLR, nx4, nx10, NOT_nx4, buffer_ready_dup0, nx302, 
      nx201, nx211, nx221, nx231, nx241, nx251, nx261, nx271, nx281, nx291, 
      nx301, nx311, nx321, nx331, nx341, nx351, nx361, nx371, nx381, nx391, 
      nx401, nx411, nx421, nx431, nx441, nx451, nx461, nx471, nx481, nx491, 
      nx501, nx511, nx521, nx531, nx541, nx551, nx561, nx571, nx581, nx591, 
      nx601, nx611, nx621, nx631, nx641, nx651, nx661, nx671, nx681, nx691, 
      nx701, nx711, nx721, nx731, nx741, nx751, nx761, nx771, nx781, nx791, 
      nx801, nx811, nx821, nx831, nx841, nx851, nx861, nx875, nx879, nx996, 
      nx1103, nx1105, nx1107, nx1109, nx1111, nx1113, nx1115, nx1117, nx1119, 
      nx1121, nx1131, nx1133, nx1137, nx1139, nx1141, nx1143, nx1145, nx1147, 
      nx1151, nx1161, nx1167, nx1169, nx1171, nx1173, nx1175, nx1177, nx1179, 
      nx1181, nx1183, nx1185, nx1187, nx1189, nx1191, nx1193, nx1195: 
   std_logic ;

begin
   output1(15) <= output1_15_EXMPLR ;
   output1(14) <= output1_14_EXMPLR ;
   output1(13) <= output1_13_EXMPLR ;
   output1(12) <= output1_12_EXMPLR ;
   output1(11) <= output1_11_EXMPLR ;
   output1(10) <= output1_10_EXMPLR ;
   output1(9) <= output1_9_EXMPLR ;
   output1(8) <= output1_8_EXMPLR ;
   output1(7) <= output1_7_EXMPLR ;
   output1(6) <= output1_6_EXMPLR ;
   output1(5) <= output1_5_EXMPLR ;
   output1(4) <= output1_4_EXMPLR ;
   output1(3) <= output1_3_EXMPLR ;
   output1(2) <= output1_2_EXMPLR ;
   output1(1) <= output1_1_EXMPLR ;
   output1(0) <= output1_0_EXMPLR ;
   output2(15) <= output2_15_EXMPLR ;
   output2(14) <= output2_14_EXMPLR ;
   output2(13) <= output2_13_EXMPLR ;
   output2(12) <= output2_12_EXMPLR ;
   output2(11) <= output2_11_EXMPLR ;
   output2(10) <= output2_10_EXMPLR ;
   output2(9) <= output2_9_EXMPLR ;
   output2(8) <= output2_8_EXMPLR ;
   output2(7) <= output2_7_EXMPLR ;
   output2(6) <= output2_6_EXMPLR ;
   output2(5) <= output2_5_EXMPLR ;
   output2(4) <= output2_4_EXMPLR ;
   output2(3) <= output2_3_EXMPLR ;
   output2(2) <= output2_2_EXMPLR ;
   output2(1) <= output2_1_EXMPLR ;
   output2(0) <= output2_0_EXMPLR ;
   buffer_ready <= buffer_ready_EXMPLR ;
   ready <= ready_EXMPLR ;
   gen_comp_pipeline : ComputationPipeline port map ( img_data_0_15=>
      img_data_0_15, img_data_0_14=>img_data_0_14, img_data_0_13=>
      img_data_0_13, img_data_0_12=>img_data_0_12, img_data_0_11=>
      img_data_0_11, img_data_0_10=>img_data_0_10, img_data_0_9=>
      img_data_0_9, img_data_0_8=>img_data_0_8, img_data_0_7=>img_data_0_7, 
      img_data_0_6=>img_data_0_6, img_data_0_5=>img_data_0_5, img_data_0_4=>
      img_data_0_4, img_data_0_3=>img_data_0_3, img_data_0_2=>img_data_0_2, 
      img_data_0_1=>img_data_0_1, img_data_0_0=>img_data_0_0, img_data_1_15
      =>nx1103, img_data_1_14=>img_data_1_14, img_data_1_13=>img_data_1_13, 
      img_data_1_12=>img_data_1_12, img_data_1_11=>img_data_1_11, 
      img_data_1_10=>img_data_1_10, img_data_1_9=>img_data_1_9, img_data_1_8
      =>img_data_1_8, img_data_1_7=>img_data_1_7, img_data_1_6=>img_data_1_6, 
      img_data_1_5=>img_data_1_5, img_data_1_4=>img_data_1_4, img_data_1_3=>
      img_data_1_3, img_data_1_2=>img_data_1_2, img_data_1_1=>img_data_1_1, 
      img_data_1_0=>img_data_1_0, img_data_2_15=>nx1105, img_data_2_14=>
      img_data_2_14, img_data_2_13=>img_data_2_13, img_data_2_12=>
      img_data_2_12, img_data_2_11=>img_data_2_11, img_data_2_10=>
      img_data_2_10, img_data_2_9=>img_data_2_9, img_data_2_8=>img_data_2_8, 
      img_data_2_7=>img_data_2_7, img_data_2_6=>img_data_2_6, img_data_2_5=>
      img_data_2_5, img_data_2_4=>img_data_2_4, img_data_2_3=>img_data_2_3, 
      img_data_2_2=>img_data_2_2, img_data_2_1=>img_data_2_1, img_data_2_0=>
      img_data_2_0, img_data_3_15=>img_data_3_15, img_data_3_14=>
      img_data_3_14, img_data_3_13=>img_data_3_13, img_data_3_12=>
      img_data_3_12, img_data_3_11=>img_data_3_11, img_data_3_10=>
      img_data_3_10, img_data_3_9=>img_data_3_9, img_data_3_8=>img_data_3_8, 
      img_data_3_7=>img_data_3_7, img_data_3_6=>img_data_3_6, img_data_3_5=>
      img_data_3_5, img_data_3_4=>img_data_3_4, img_data_3_3=>img_data_3_3, 
      img_data_3_2=>img_data_3_2, img_data_3_1=>img_data_3_1, img_data_3_0=>
      img_data_3_0, img_data_4_15=>img_data_4_15, img_data_4_14=>
      img_data_4_14, img_data_4_13=>img_data_4_13, img_data_4_12=>
      img_data_4_12, img_data_4_11=>img_data_4_11, img_data_4_10=>
      img_data_4_10, img_data_4_9=>img_data_4_9, img_data_4_8=>img_data_4_8, 
      img_data_4_7=>img_data_4_7, img_data_4_6=>img_data_4_6, img_data_4_5=>
      img_data_4_5, img_data_4_4=>img_data_4_4, img_data_4_3=>img_data_4_3, 
      img_data_4_2=>img_data_4_2, img_data_4_1=>img_data_4_1, img_data_4_0=>
      img_data_4_0, img_data_5_15=>img_data_5_15, img_data_5_14=>
      img_data_5_14, img_data_5_13=>img_data_5_13, img_data_5_12=>
      img_data_5_12, img_data_5_11=>img_data_5_11, img_data_5_10=>
      img_data_5_10, img_data_5_9=>img_data_5_9, img_data_5_8=>img_data_5_8, 
      img_data_5_7=>img_data_5_7, img_data_5_6=>img_data_5_6, img_data_5_5=>
      img_data_5_5, img_data_5_4=>img_data_5_4, img_data_5_3=>img_data_5_3, 
      img_data_5_2=>img_data_5_2, img_data_5_1=>img_data_5_1, img_data_5_0=>
      img_data_5_0, img_data_6_15=>nx1107, img_data_6_14=>img_data_6_14, 
      img_data_6_13=>img_data_6_13, img_data_6_12=>img_data_6_12, 
      img_data_6_11=>img_data_6_11, img_data_6_10=>img_data_6_10, 
      img_data_6_9=>img_data_6_9, img_data_6_8=>img_data_6_8, img_data_6_7=>
      img_data_6_7, img_data_6_6=>img_data_6_6, img_data_6_5=>img_data_6_5, 
      img_data_6_4=>img_data_6_4, img_data_6_3=>img_data_6_3, img_data_6_2=>
      img_data_6_2, img_data_6_1=>img_data_6_1, img_data_6_0=>img_data_6_0, 
      img_data_7_15=>img_data_7_15, img_data_7_14=>img_data_7_14, 
      img_data_7_13=>img_data_7_13, img_data_7_12=>img_data_7_12, 
      img_data_7_11=>img_data_7_11, img_data_7_10=>img_data_7_10, 
      img_data_7_9=>img_data_7_9, img_data_7_8=>img_data_7_8, img_data_7_7=>
      img_data_7_7, img_data_7_6=>img_data_7_6, img_data_7_5=>img_data_7_5, 
      img_data_7_4=>img_data_7_4, img_data_7_3=>img_data_7_3, img_data_7_2=>
      img_data_7_2, img_data_7_1=>img_data_7_1, img_data_7_0=>img_data_7_0, 
      img_data_8_15=>img_data_8_15, img_data_8_14=>img_data_8_14, 
      img_data_8_13=>img_data_8_13, img_data_8_12=>img_data_8_12, 
      img_data_8_11=>img_data_8_11, img_data_8_10=>img_data_8_10, 
      img_data_8_9=>img_data_8_9, img_data_8_8=>img_data_8_8, img_data_8_7=>
      img_data_8_7, img_data_8_6=>img_data_8_6, img_data_8_5=>img_data_8_5, 
      img_data_8_4=>img_data_8_4, img_data_8_3=>img_data_8_3, img_data_8_2=>
      img_data_8_2, img_data_8_1=>img_data_8_1, img_data_8_0=>img_data_8_0, 
      img_data_9_15=>img_data_9_15, img_data_9_14=>img_data_9_14, 
      img_data_9_13=>img_data_9_13, img_data_9_12=>img_data_9_12, 
      img_data_9_11=>img_data_9_11, img_data_9_10=>img_data_9_10, 
      img_data_9_9=>img_data_9_9, img_data_9_8=>img_data_9_8, img_data_9_7=>
      img_data_9_7, img_data_9_6=>img_data_9_6, img_data_9_5=>img_data_9_5, 
      img_data_9_4=>img_data_9_4, img_data_9_3=>img_data_9_3, img_data_9_2=>
      img_data_9_2, img_data_9_1=>img_data_9_1, img_data_9_0=>img_data_9_0, 
      img_data_10_15=>img_data_10_15, img_data_10_14=>img_data_10_14, 
      img_data_10_13=>img_data_10_13, img_data_10_12=>img_data_10_12, 
      img_data_10_11=>img_data_10_11, img_data_10_10=>img_data_10_10, 
      img_data_10_9=>img_data_10_9, img_data_10_8=>img_data_10_8, 
      img_data_10_7=>img_data_10_7, img_data_10_6=>img_data_10_6, 
      img_data_10_5=>img_data_10_5, img_data_10_4=>img_data_10_4, 
      img_data_10_3=>img_data_10_3, img_data_10_2=>img_data_10_2, 
      img_data_10_1=>img_data_10_1, img_data_10_0=>img_data_10_0, 
      img_data_11_15=>img_data_11_15, img_data_11_14=>img_data_11_14, 
      img_data_11_13=>img_data_11_13, img_data_11_12=>img_data_11_12, 
      img_data_11_11=>img_data_11_11, img_data_11_10=>img_data_11_10, 
      img_data_11_9=>img_data_11_9, img_data_11_8=>img_data_11_8, 
      img_data_11_7=>img_data_11_7, img_data_11_6=>img_data_11_6, 
      img_data_11_5=>img_data_11_5, img_data_11_4=>img_data_11_4, 
      img_data_11_3=>img_data_11_3, img_data_11_2=>img_data_11_2, 
      img_data_11_1=>img_data_11_1, img_data_11_0=>img_data_11_0, 
      img_data_12_15=>img_data_12_15, img_data_12_14=>img_data_12_14, 
      img_data_12_13=>img_data_12_13, img_data_12_12=>img_data_12_12, 
      img_data_12_11=>img_data_12_11, img_data_12_10=>img_data_12_10, 
      img_data_12_9=>img_data_12_9, img_data_12_8=>img_data_12_8, 
      img_data_12_7=>img_data_12_7, img_data_12_6=>img_data_12_6, 
      img_data_12_5=>img_data_12_5, img_data_12_4=>img_data_12_4, 
      img_data_12_3=>img_data_12_3, img_data_12_2=>img_data_12_2, 
      img_data_12_1=>img_data_12_1, img_data_12_0=>img_data_12_0, 
      img_data_13_15=>img_data_13_15, img_data_13_14=>img_data_13_14, 
      img_data_13_13=>img_data_13_13, img_data_13_12=>img_data_13_12, 
      img_data_13_11=>img_data_13_11, img_data_13_10=>img_data_13_10, 
      img_data_13_9=>img_data_13_9, img_data_13_8=>img_data_13_8, 
      img_data_13_7=>img_data_13_7, img_data_13_6=>img_data_13_6, 
      img_data_13_5=>img_data_13_5, img_data_13_4=>img_data_13_4, 
      img_data_13_3=>img_data_13_3, img_data_13_2=>img_data_13_2, 
      img_data_13_1=>img_data_13_1, img_data_13_0=>img_data_13_0, 
      img_data_14_15=>img_data_14_15, img_data_14_14=>img_data_14_14, 
      img_data_14_13=>img_data_14_13, img_data_14_12=>img_data_14_12, 
      img_data_14_11=>img_data_14_11, img_data_14_10=>img_data_14_10, 
      img_data_14_9=>img_data_14_9, img_data_14_8=>img_data_14_8, 
      img_data_14_7=>img_data_14_7, img_data_14_6=>img_data_14_6, 
      img_data_14_5=>img_data_14_5, img_data_14_4=>img_data_14_4, 
      img_data_14_3=>img_data_14_3, img_data_14_2=>img_data_14_2, 
      img_data_14_1=>img_data_14_1, img_data_14_0=>img_data_14_0, 
      img_data_15_15=>img_data_15_15, img_data_15_14=>img_data_15_14, 
      img_data_15_13=>img_data_15_13, img_data_15_12=>img_data_15_12, 
      img_data_15_11=>img_data_15_11, img_data_15_10=>img_data_15_10, 
      img_data_15_9=>img_data_15_9, img_data_15_8=>img_data_15_8, 
      img_data_15_7=>img_data_15_7, img_data_15_6=>img_data_15_6, 
      img_data_15_5=>img_data_15_5, img_data_15_4=>img_data_15_4, 
      img_data_15_3=>img_data_15_3, img_data_15_2=>img_data_15_2, 
      img_data_15_1=>img_data_15_1, img_data_15_0=>img_data_15_0, 
      img_data_16_15=>img_data_16_15, img_data_16_14=>img_data_16_14, 
      img_data_16_13=>img_data_16_13, img_data_16_12=>img_data_16_12, 
      img_data_16_11=>img_data_16_11, img_data_16_10=>img_data_16_10, 
      img_data_16_9=>img_data_16_9, img_data_16_8=>img_data_16_8, 
      img_data_16_7=>img_data_16_7, img_data_16_6=>img_data_16_6, 
      img_data_16_5=>img_data_16_5, img_data_16_4=>img_data_16_4, 
      img_data_16_3=>img_data_16_3, img_data_16_2=>img_data_16_2, 
      img_data_16_1=>img_data_16_1, img_data_16_0=>img_data_16_0, 
      img_data_17_15=>img_data_17_15, img_data_17_14=>img_data_17_14, 
      img_data_17_13=>img_data_17_13, img_data_17_12=>img_data_17_12, 
      img_data_17_11=>img_data_17_11, img_data_17_10=>img_data_17_10, 
      img_data_17_9=>img_data_17_9, img_data_17_8=>img_data_17_8, 
      img_data_17_7=>img_data_17_7, img_data_17_6=>img_data_17_6, 
      img_data_17_5=>img_data_17_5, img_data_17_4=>img_data_17_4, 
      img_data_17_3=>img_data_17_3, img_data_17_2=>img_data_17_2, 
      img_data_17_1=>img_data_17_1, img_data_17_0=>img_data_17_0, 
      img_data_18_15=>img_data_18_15, img_data_18_14=>img_data_18_14, 
      img_data_18_13=>img_data_18_13, img_data_18_12=>img_data_18_12, 
      img_data_18_11=>img_data_18_11, img_data_18_10=>img_data_18_10, 
      img_data_18_9=>img_data_18_9, img_data_18_8=>img_data_18_8, 
      img_data_18_7=>img_data_18_7, img_data_18_6=>img_data_18_6, 
      img_data_18_5=>img_data_18_5, img_data_18_4=>img_data_18_4, 
      img_data_18_3=>img_data_18_3, img_data_18_2=>img_data_18_2, 
      img_data_18_1=>img_data_18_1, img_data_18_0=>img_data_18_0, 
      img_data_19_15=>img_data_19_15, img_data_19_14=>img_data_19_14, 
      img_data_19_13=>img_data_19_13, img_data_19_12=>img_data_19_12, 
      img_data_19_11=>img_data_19_11, img_data_19_10=>img_data_19_10, 
      img_data_19_9=>img_data_19_9, img_data_19_8=>img_data_19_8, 
      img_data_19_7=>img_data_19_7, img_data_19_6=>img_data_19_6, 
      img_data_19_5=>img_data_19_5, img_data_19_4=>img_data_19_4, 
      img_data_19_3=>img_data_19_3, img_data_19_2=>img_data_19_2, 
      img_data_19_1=>img_data_19_1, img_data_19_0=>img_data_19_0, 
      img_data_20_15=>img_data_20_15, img_data_20_14=>img_data_20_14, 
      img_data_20_13=>img_data_20_13, img_data_20_12=>img_data_20_12, 
      img_data_20_11=>img_data_20_11, img_data_20_10=>img_data_20_10, 
      img_data_20_9=>img_data_20_9, img_data_20_8=>img_data_20_8, 
      img_data_20_7=>img_data_20_7, img_data_20_6=>img_data_20_6, 
      img_data_20_5=>img_data_20_5, img_data_20_4=>img_data_20_4, 
      img_data_20_3=>img_data_20_3, img_data_20_2=>img_data_20_2, 
      img_data_20_1=>img_data_20_1, img_data_20_0=>img_data_20_0, 
      img_data_21_15=>img_data_21_15, img_data_21_14=>img_data_21_14, 
      img_data_21_13=>img_data_21_13, img_data_21_12=>img_data_21_12, 
      img_data_21_11=>img_data_21_11, img_data_21_10=>img_data_21_10, 
      img_data_21_9=>img_data_21_9, img_data_21_8=>img_data_21_8, 
      img_data_21_7=>img_data_21_7, img_data_21_6=>img_data_21_6, 
      img_data_21_5=>img_data_21_5, img_data_21_4=>img_data_21_4, 
      img_data_21_3=>img_data_21_3, img_data_21_2=>img_data_21_2, 
      img_data_21_1=>img_data_21_1, img_data_21_0=>img_data_21_0, 
      img_data_22_15=>img_data_22_15, img_data_22_14=>img_data_22_14, 
      img_data_22_13=>img_data_22_13, img_data_22_12=>img_data_22_12, 
      img_data_22_11=>img_data_22_11, img_data_22_10=>img_data_22_10, 
      img_data_22_9=>img_data_22_9, img_data_22_8=>img_data_22_8, 
      img_data_22_7=>img_data_22_7, img_data_22_6=>img_data_22_6, 
      img_data_22_5=>img_data_22_5, img_data_22_4=>img_data_22_4, 
      img_data_22_3=>img_data_22_3, img_data_22_2=>img_data_22_2, 
      img_data_22_1=>img_data_22_1, img_data_22_0=>img_data_22_0, 
      img_data_23_15=>img_data_23_15, img_data_23_14=>img_data_23_14, 
      img_data_23_13=>img_data_23_13, img_data_23_12=>img_data_23_12, 
      img_data_23_11=>img_data_23_11, img_data_23_10=>img_data_23_10, 
      img_data_23_9=>img_data_23_9, img_data_23_8=>img_data_23_8, 
      img_data_23_7=>img_data_23_7, img_data_23_6=>img_data_23_6, 
      img_data_23_5=>img_data_23_5, img_data_23_4=>img_data_23_4, 
      img_data_23_3=>img_data_23_3, img_data_23_2=>img_data_23_2, 
      img_data_23_1=>img_data_23_1, img_data_23_0=>img_data_23_0, 
      img_data_24_15=>img_data_24_15, img_data_24_14=>img_data_24_14, 
      img_data_24_13=>img_data_24_13, img_data_24_12=>img_data_24_12, 
      img_data_24_11=>img_data_24_11, img_data_24_10=>img_data_24_10, 
      img_data_24_9=>img_data_24_9, img_data_24_8=>img_data_24_8, 
      img_data_24_7=>img_data_24_7, img_data_24_6=>img_data_24_6, 
      img_data_24_5=>img_data_24_5, img_data_24_4=>img_data_24_4, 
      img_data_24_3=>img_data_24_3, img_data_24_2=>img_data_24_2, 
      img_data_24_1=>img_data_24_1, img_data_24_0=>img_data_24_0, 
      filter_data_0_15=>filter_data_0_15, filter_data_0_14=>filter_data_0_14, 
      filter_data_0_13=>filter_data_0_13, filter_data_0_12=>filter_data_0_12, 
      filter_data_0_11=>filter_data_0_11, filter_data_0_10=>filter_data_0_10, 
      filter_data_0_9=>filter_data_0_9, filter_data_0_8=>filter_data_0_8, 
      filter_data_0_7=>filter_data_0_7, filter_data_0_6=>filter_data_0_6, 
      filter_data_0_5=>filter_data_0_5, filter_data_0_4=>filter_data_0_4, 
      filter_data_0_3=>filter_data_0_3, filter_data_0_2=>filter_data_0_2, 
      filter_data_0_1=>filter_data_0_1, filter_data_0_0=>filter_data_0_0, 
      filter_data_1_15=>filter_data_1_15, filter_data_1_14=>filter_data_1_14, 
      filter_data_1_13=>filter_data_1_13, filter_data_1_12=>filter_data_1_12, 
      filter_data_1_11=>filter_data_1_11, filter_data_1_10=>filter_data_1_10, 
      filter_data_1_9=>filter_data_1_9, filter_data_1_8=>filter_data_1_8, 
      filter_data_1_7=>filter_data_1_7, filter_data_1_6=>filter_data_1_6, 
      filter_data_1_5=>filter_data_1_5, filter_data_1_4=>filter_data_1_4, 
      filter_data_1_3=>filter_data_1_3, filter_data_1_2=>filter_data_1_2, 
      filter_data_1_1=>filter_data_1_1, filter_data_1_0=>filter_data_1_0, 
      filter_data_2_15=>filter_data_2_15, filter_data_2_14=>filter_data_2_14, 
      filter_data_2_13=>filter_data_2_13, filter_data_2_12=>filter_data_2_12, 
      filter_data_2_11=>filter_data_2_11, filter_data_2_10=>filter_data_2_10, 
      filter_data_2_9=>filter_data_2_9, filter_data_2_8=>filter_data_2_8, 
      filter_data_2_7=>filter_data_2_7, filter_data_2_6=>filter_data_2_6, 
      filter_data_2_5=>filter_data_2_5, filter_data_2_4=>filter_data_2_4, 
      filter_data_2_3=>filter_data_2_3, filter_data_2_2=>filter_data_2_2, 
      filter_data_2_1=>filter_data_2_1, filter_data_2_0=>filter_data_2_0, 
      filter_data_3_15=>filter_data_3_15, filter_data_3_14=>filter_data_3_14, 
      filter_data_3_13=>filter_data_3_13, filter_data_3_12=>filter_data_3_12, 
      filter_data_3_11=>filter_data_3_11, filter_data_3_10=>filter_data_3_10, 
      filter_data_3_9=>filter_data_3_9, filter_data_3_8=>filter_data_3_8, 
      filter_data_3_7=>filter_data_3_7, filter_data_3_6=>filter_data_3_6, 
      filter_data_3_5=>filter_data_3_5, filter_data_3_4=>filter_data_3_4, 
      filter_data_3_3=>filter_data_3_3, filter_data_3_2=>filter_data_3_2, 
      filter_data_3_1=>filter_data_3_1, filter_data_3_0=>filter_data_3_0, 
      filter_data_4_15=>filter_data_4_15, filter_data_4_14=>filter_data_4_14, 
      filter_data_4_13=>filter_data_4_13, filter_data_4_12=>filter_data_4_12, 
      filter_data_4_11=>filter_data_4_11, filter_data_4_10=>filter_data_4_10, 
      filter_data_4_9=>filter_data_4_9, filter_data_4_8=>filter_data_4_8, 
      filter_data_4_7=>filter_data_4_7, filter_data_4_6=>filter_data_4_6, 
      filter_data_4_5=>filter_data_4_5, filter_data_4_4=>filter_data_4_4, 
      filter_data_4_3=>filter_data_4_3, filter_data_4_2=>filter_data_4_2, 
      filter_data_4_1=>filter_data_4_1, filter_data_4_0=>filter_data_4_0, 
      filter_data_5_15=>filter_data_5_15, filter_data_5_14=>filter_data_5_14, 
      filter_data_5_13=>filter_data_5_13, filter_data_5_12=>filter_data_5_12, 
      filter_data_5_11=>filter_data_5_11, filter_data_5_10=>filter_data_5_10, 
      filter_data_5_9=>filter_data_5_9, filter_data_5_8=>filter_data_5_8, 
      filter_data_5_7=>filter_data_5_7, filter_data_5_6=>filter_data_5_6, 
      filter_data_5_5=>filter_data_5_5, filter_data_5_4=>filter_data_5_4, 
      filter_data_5_3=>filter_data_5_3, filter_data_5_2=>filter_data_5_2, 
      filter_data_5_1=>filter_data_5_1, filter_data_5_0=>filter_data_5_0, 
      filter_data_6_15=>filter_data_6_15, filter_data_6_14=>filter_data_6_14, 
      filter_data_6_13=>filter_data_6_13, filter_data_6_12=>filter_data_6_12, 
      filter_data_6_11=>filter_data_6_11, filter_data_6_10=>filter_data_6_10, 
      filter_data_6_9=>filter_data_6_9, filter_data_6_8=>filter_data_6_8, 
      filter_data_6_7=>filter_data_6_7, filter_data_6_6=>filter_data_6_6, 
      filter_data_6_5=>filter_data_6_5, filter_data_6_4=>filter_data_6_4, 
      filter_data_6_3=>filter_data_6_3, filter_data_6_2=>filter_data_6_2, 
      filter_data_6_1=>filter_data_6_1, filter_data_6_0=>filter_data_6_0, 
      filter_data_7_15=>filter_data_7_15, filter_data_7_14=>filter_data_7_14, 
      filter_data_7_13=>filter_data_7_13, filter_data_7_12=>filter_data_7_12, 
      filter_data_7_11=>filter_data_7_11, filter_data_7_10=>filter_data_7_10, 
      filter_data_7_9=>filter_data_7_9, filter_data_7_8=>filter_data_7_8, 
      filter_data_7_7=>filter_data_7_7, filter_data_7_6=>filter_data_7_6, 
      filter_data_7_5=>filter_data_7_5, filter_data_7_4=>filter_data_7_4, 
      filter_data_7_3=>filter_data_7_3, filter_data_7_2=>filter_data_7_2, 
      filter_data_7_1=>filter_data_7_1, filter_data_7_0=>filter_data_7_0, 
      filter_data_8_15=>filter_data_8_15, filter_data_8_14=>filter_data_8_14, 
      filter_data_8_13=>filter_data_8_13, filter_data_8_12=>filter_data_8_12, 
      filter_data_8_11=>filter_data_8_11, filter_data_8_10=>filter_data_8_10, 
      filter_data_8_9=>filter_data_8_9, filter_data_8_8=>filter_data_8_8, 
      filter_data_8_7=>filter_data_8_7, filter_data_8_6=>filter_data_8_6, 
      filter_data_8_5=>filter_data_8_5, filter_data_8_4=>filter_data_8_4, 
      filter_data_8_3=>filter_data_8_3, filter_data_8_2=>filter_data_8_2, 
      filter_data_8_1=>filter_data_8_1, filter_data_8_0=>filter_data_8_0, 
      filter_data_9_15=>filter_data_9_15, filter_data_9_14=>filter_data_9_14, 
      filter_data_9_13=>filter_data_9_13, filter_data_9_12=>filter_data_9_12, 
      filter_data_9_11=>filter_data_9_11, filter_data_9_10=>filter_data_9_10, 
      filter_data_9_9=>filter_data_9_9, filter_data_9_8=>filter_data_9_8, 
      filter_data_9_7=>filter_data_9_7, filter_data_9_6=>filter_data_9_6, 
      filter_data_9_5=>filter_data_9_5, filter_data_9_4=>filter_data_9_4, 
      filter_data_9_3=>filter_data_9_3, filter_data_9_2=>filter_data_9_2, 
      filter_data_9_1=>filter_data_9_1, filter_data_9_0=>filter_data_9_0, 
      filter_data_10_15=>filter_data_10_15, filter_data_10_14=>
      filter_data_10_14, filter_data_10_13=>filter_data_10_13, 
      filter_data_10_12=>filter_data_10_12, filter_data_10_11=>
      filter_data_10_11, filter_data_10_10=>filter_data_10_10, 
      filter_data_10_9=>filter_data_10_9, filter_data_10_8=>filter_data_10_8, 
      filter_data_10_7=>filter_data_10_7, filter_data_10_6=>filter_data_10_6, 
      filter_data_10_5=>filter_data_10_5, filter_data_10_4=>filter_data_10_4, 
      filter_data_10_3=>filter_data_10_3, filter_data_10_2=>filter_data_10_2, 
      filter_data_10_1=>filter_data_10_1, filter_data_10_0=>filter_data_10_0, 
      filter_data_11_15=>filter_data_11_15, filter_data_11_14=>
      filter_data_11_14, filter_data_11_13=>filter_data_11_13, 
      filter_data_11_12=>filter_data_11_12, filter_data_11_11=>
      filter_data_11_11, filter_data_11_10=>filter_data_11_10, 
      filter_data_11_9=>filter_data_11_9, filter_data_11_8=>filter_data_11_8, 
      filter_data_11_7=>filter_data_11_7, filter_data_11_6=>filter_data_11_6, 
      filter_data_11_5=>filter_data_11_5, filter_data_11_4=>filter_data_11_4, 
      filter_data_11_3=>filter_data_11_3, filter_data_11_2=>filter_data_11_2, 
      filter_data_11_1=>filter_data_11_1, filter_data_11_0=>filter_data_11_0, 
      filter_data_12_15=>filter_data_12_15, filter_data_12_14=>
      filter_data_12_14, filter_data_12_13=>filter_data_12_13, 
      filter_data_12_12=>filter_data_12_12, filter_data_12_11=>
      filter_data_12_11, filter_data_12_10=>filter_data_12_10, 
      filter_data_12_9=>filter_data_12_9, filter_data_12_8=>filter_data_12_8, 
      filter_data_12_7=>filter_data_12_7, filter_data_12_6=>filter_data_12_6, 
      filter_data_12_5=>filter_data_12_5, filter_data_12_4=>filter_data_12_4, 
      filter_data_12_3=>filter_data_12_3, filter_data_12_2=>filter_data_12_2, 
      filter_data_12_1=>filter_data_12_1, filter_data_12_0=>filter_data_12_0, 
      filter_data_13_15=>filter_data_13_15, filter_data_13_14=>
      filter_data_13_14, filter_data_13_13=>filter_data_13_13, 
      filter_data_13_12=>filter_data_13_12, filter_data_13_11=>
      filter_data_13_11, filter_data_13_10=>filter_data_13_10, 
      filter_data_13_9=>filter_data_13_9, filter_data_13_8=>filter_data_13_8, 
      filter_data_13_7=>filter_data_13_7, filter_data_13_6=>filter_data_13_6, 
      filter_data_13_5=>filter_data_13_5, filter_data_13_4=>filter_data_13_4, 
      filter_data_13_3=>filter_data_13_3, filter_data_13_2=>filter_data_13_2, 
      filter_data_13_1=>filter_data_13_1, filter_data_13_0=>filter_data_13_0, 
      filter_data_14_15=>filter_data_14_15, filter_data_14_14=>
      filter_data_14_14, filter_data_14_13=>filter_data_14_13, 
      filter_data_14_12=>filter_data_14_12, filter_data_14_11=>
      filter_data_14_11, filter_data_14_10=>filter_data_14_10, 
      filter_data_14_9=>filter_data_14_9, filter_data_14_8=>filter_data_14_8, 
      filter_data_14_7=>filter_data_14_7, filter_data_14_6=>filter_data_14_6, 
      filter_data_14_5=>filter_data_14_5, filter_data_14_4=>filter_data_14_4, 
      filter_data_14_3=>filter_data_14_3, filter_data_14_2=>filter_data_14_2, 
      filter_data_14_1=>filter_data_14_1, filter_data_14_0=>filter_data_14_0, 
      filter_data_15_15=>filter_data_15_15, filter_data_15_14=>
      filter_data_15_14, filter_data_15_13=>filter_data_15_13, 
      filter_data_15_12=>filter_data_15_12, filter_data_15_11=>
      filter_data_15_11, filter_data_15_10=>filter_data_15_10, 
      filter_data_15_9=>filter_data_15_9, filter_data_15_8=>filter_data_15_8, 
      filter_data_15_7=>filter_data_15_7, filter_data_15_6=>filter_data_15_6, 
      filter_data_15_5=>filter_data_15_5, filter_data_15_4=>filter_data_15_4, 
      filter_data_15_3=>filter_data_15_3, filter_data_15_2=>filter_data_15_2, 
      filter_data_15_1=>filter_data_15_1, filter_data_15_0=>filter_data_15_0, 
      filter_data_16_15=>filter_data_16_15, filter_data_16_14=>
      filter_data_16_14, filter_data_16_13=>filter_data_16_13, 
      filter_data_16_12=>filter_data_16_12, filter_data_16_11=>
      filter_data_16_11, filter_data_16_10=>filter_data_16_10, 
      filter_data_16_9=>filter_data_16_9, filter_data_16_8=>filter_data_16_8, 
      filter_data_16_7=>filter_data_16_7, filter_data_16_6=>filter_data_16_6, 
      filter_data_16_5=>filter_data_16_5, filter_data_16_4=>filter_data_16_4, 
      filter_data_16_3=>filter_data_16_3, filter_data_16_2=>filter_data_16_2, 
      filter_data_16_1=>filter_data_16_1, filter_data_16_0=>filter_data_16_0, 
      filter_data_17_15=>filter_data_17_15, filter_data_17_14=>
      filter_data_17_14, filter_data_17_13=>filter_data_17_13, 
      filter_data_17_12=>filter_data_17_12, filter_data_17_11=>
      filter_data_17_11, filter_data_17_10=>filter_data_17_10, 
      filter_data_17_9=>filter_data_17_9, filter_data_17_8=>filter_data_17_8, 
      filter_data_17_7=>filter_data_17_7, filter_data_17_6=>filter_data_17_6, 
      filter_data_17_5=>filter_data_17_5, filter_data_17_4=>filter_data_17_4, 
      filter_data_17_3=>filter_data_17_3, filter_data_17_2=>filter_data_17_2, 
      filter_data_17_1=>filter_data_17_1, filter_data_17_0=>filter_data_17_0, 
      filter_data_18_15=>filter_data_18_15, filter_data_18_14=>
      filter_data_18_14, filter_data_18_13=>filter_data_18_13, 
      filter_data_18_12=>filter_data_18_12, filter_data_18_11=>
      filter_data_18_11, filter_data_18_10=>filter_data_18_10, 
      filter_data_18_9=>filter_data_18_9, filter_data_18_8=>filter_data_18_8, 
      filter_data_18_7=>filter_data_18_7, filter_data_18_6=>filter_data_18_6, 
      filter_data_18_5=>filter_data_18_5, filter_data_18_4=>filter_data_18_4, 
      filter_data_18_3=>filter_data_18_3, filter_data_18_2=>filter_data_18_2, 
      filter_data_18_1=>filter_data_18_1, filter_data_18_0=>filter_data_18_0, 
      filter_data_19_15=>filter_data_19_15, filter_data_19_14=>
      filter_data_19_14, filter_data_19_13=>filter_data_19_13, 
      filter_data_19_12=>filter_data_19_12, filter_data_19_11=>
      filter_data_19_11, filter_data_19_10=>filter_data_19_10, 
      filter_data_19_9=>filter_data_19_9, filter_data_19_8=>filter_data_19_8, 
      filter_data_19_7=>filter_data_19_7, filter_data_19_6=>filter_data_19_6, 
      filter_data_19_5=>filter_data_19_5, filter_data_19_4=>filter_data_19_4, 
      filter_data_19_3=>filter_data_19_3, filter_data_19_2=>filter_data_19_2, 
      filter_data_19_1=>filter_data_19_1, filter_data_19_0=>filter_data_19_0, 
      filter_data_20_15=>filter_data_20_15, filter_data_20_14=>
      filter_data_20_14, filter_data_20_13=>filter_data_20_13, 
      filter_data_20_12=>filter_data_20_12, filter_data_20_11=>
      filter_data_20_11, filter_data_20_10=>filter_data_20_10, 
      filter_data_20_9=>filter_data_20_9, filter_data_20_8=>filter_data_20_8, 
      filter_data_20_7=>filter_data_20_7, filter_data_20_6=>filter_data_20_6, 
      filter_data_20_5=>filter_data_20_5, filter_data_20_4=>filter_data_20_4, 
      filter_data_20_3=>filter_data_20_3, filter_data_20_2=>filter_data_20_2, 
      filter_data_20_1=>filter_data_20_1, filter_data_20_0=>filter_data_20_0, 
      filter_data_21_15=>filter_data_21_15, filter_data_21_14=>
      filter_data_21_14, filter_data_21_13=>filter_data_21_13, 
      filter_data_21_12=>filter_data_21_12, filter_data_21_11=>
      filter_data_21_11, filter_data_21_10=>filter_data_21_10, 
      filter_data_21_9=>filter_data_21_9, filter_data_21_8=>filter_data_21_8, 
      filter_data_21_7=>filter_data_21_7, filter_data_21_6=>filter_data_21_6, 
      filter_data_21_5=>filter_data_21_5, filter_data_21_4=>filter_data_21_4, 
      filter_data_21_3=>filter_data_21_3, filter_data_21_2=>filter_data_21_2, 
      filter_data_21_1=>filter_data_21_1, filter_data_21_0=>filter_data_21_0, 
      filter_data_22_15=>filter_data_22_15, filter_data_22_14=>
      filter_data_22_14, filter_data_22_13=>filter_data_22_13, 
      filter_data_22_12=>filter_data_22_12, filter_data_22_11=>
      filter_data_22_11, filter_data_22_10=>filter_data_22_10, 
      filter_data_22_9=>filter_data_22_9, filter_data_22_8=>filter_data_22_8, 
      filter_data_22_7=>filter_data_22_7, filter_data_22_6=>filter_data_22_6, 
      filter_data_22_5=>filter_data_22_5, filter_data_22_4=>filter_data_22_4, 
      filter_data_22_3=>filter_data_22_3, filter_data_22_2=>filter_data_22_2, 
      filter_data_22_1=>filter_data_22_1, filter_data_22_0=>filter_data_22_0, 
      filter_data_23_15=>filter_data_23_15, filter_data_23_14=>
      filter_data_23_14, filter_data_23_13=>filter_data_23_13, 
      filter_data_23_12=>filter_data_23_12, filter_data_23_11=>
      filter_data_23_11, filter_data_23_10=>filter_data_23_10, 
      filter_data_23_9=>filter_data_23_9, filter_data_23_8=>filter_data_23_8, 
      filter_data_23_7=>filter_data_23_7, filter_data_23_6=>filter_data_23_6, 
      filter_data_23_5=>filter_data_23_5, filter_data_23_4=>filter_data_23_4, 
      filter_data_23_3=>filter_data_23_3, filter_data_23_2=>filter_data_23_2, 
      filter_data_23_1=>filter_data_23_1, filter_data_23_0=>filter_data_23_0, 
      filter_data_24_15=>filter_data_24_15, filter_data_24_14=>
      filter_data_24_14, filter_data_24_13=>filter_data_24_13, 
      filter_data_24_12=>filter_data_24_12, filter_data_24_11=>
      filter_data_24_11, filter_data_24_10=>filter_data_24_10, 
      filter_data_24_9=>filter_data_24_9, filter_data_24_8=>filter_data_24_8, 
      filter_data_24_7=>filter_data_24_7, filter_data_24_6=>filter_data_24_6, 
      filter_data_24_5=>filter_data_24_5, filter_data_24_4=>filter_data_24_4, 
      filter_data_24_3=>filter_data_24_3, filter_data_24_2=>filter_data_24_2, 
      filter_data_24_1=>filter_data_24_1, filter_data_24_0=>filter_data_24_0, 
      d_arr_0_31=>d_cache_arr_0_31, d_arr_0_30=>d_cache_arr_0_30, d_arr_0_29
      =>d_cache_arr_0_29, d_arr_0_28=>d_cache_arr_0_28, d_arr_0_27=>
      d_cache_arr_0_27, d_arr_0_26=>d_cache_arr_0_26, d_arr_0_25=>
      d_cache_arr_0_25, d_arr_0_24=>d_cache_arr_0_24, d_arr_0_23=>
      d_cache_arr_0_23, d_arr_0_22=>d_cache_arr_0_22, d_arr_0_21=>
      d_cache_arr_0_21, d_arr_0_20=>d_cache_arr_0_20, d_arr_0_19=>
      d_cache_arr_0_19, d_arr_0_18=>d_cache_arr_0_18, d_arr_0_17=>
      d_cache_arr_0_17, d_arr_0_16=>d_cache_arr_0_16, d_arr_0_15=>
      d_cache_arr_0_15, d_arr_0_14=>d_cache_arr_0_14, d_arr_0_13=>
      d_cache_arr_0_13, d_arr_0_12=>d_cache_arr_0_12, d_arr_0_11=>
      d_cache_arr_0_11, d_arr_0_10=>d_cache_arr_0_10, d_arr_0_9=>
      d_cache_arr_0_9, d_arr_0_8=>d_cache_arr_0_8, d_arr_0_7=>
      d_cache_arr_0_7, d_arr_0_6=>d_cache_arr_0_6, d_arr_0_5=>
      d_cache_arr_0_5, d_arr_0_4=>d_cache_arr_0_4, d_arr_0_3=>
      d_cache_arr_0_3, d_arr_0_2=>d_cache_arr_0_2, d_arr_0_1=>
      d_cache_arr_0_1, d_arr_0_0=>d_cache_arr_0_0, d_arr_1_31=>
      d_cache_arr_1_31, d_arr_1_30=>d_cache_arr_1_30, d_arr_1_29=>
      d_cache_arr_1_29, d_arr_1_28=>d_cache_arr_1_28, d_arr_1_27=>
      d_cache_arr_1_27, d_arr_1_26=>d_cache_arr_1_26, d_arr_1_25=>
      d_cache_arr_1_25, d_arr_1_24=>d_cache_arr_1_24, d_arr_1_23=>
      d_cache_arr_1_23, d_arr_1_22=>d_cache_arr_1_22, d_arr_1_21=>
      d_cache_arr_1_21, d_arr_1_20=>d_cache_arr_1_20, d_arr_1_19=>
      d_cache_arr_1_19, d_arr_1_18=>d_cache_arr_1_18, d_arr_1_17=>
      d_cache_arr_1_17, d_arr_1_16=>d_cache_arr_1_16, d_arr_1_15=>
      d_cache_arr_1_15, d_arr_1_14=>d_cache_arr_1_14, d_arr_1_13=>
      d_cache_arr_1_13, d_arr_1_12=>d_cache_arr_1_12, d_arr_1_11=>
      d_cache_arr_1_11, d_arr_1_10=>d_cache_arr_1_10, d_arr_1_9=>
      d_cache_arr_1_9, d_arr_1_8=>d_cache_arr_1_8, d_arr_1_7=>
      d_cache_arr_1_7, d_arr_1_6=>d_cache_arr_1_6, d_arr_1_5=>
      d_cache_arr_1_5, d_arr_1_4=>d_cache_arr_1_4, d_arr_1_3=>
      d_cache_arr_1_3, d_arr_1_2=>d_cache_arr_1_2, d_arr_1_1=>
      d_cache_arr_1_1, d_arr_1_0=>d_cache_arr_1_0, d_arr_2_31=>
      d_cache_arr_2_31, d_arr_2_30=>d_cache_arr_2_30, d_arr_2_29=>
      d_cache_arr_2_29, d_arr_2_28=>d_cache_arr_2_28, d_arr_2_27=>
      d_cache_arr_2_27, d_arr_2_26=>d_cache_arr_2_26, d_arr_2_25=>
      d_cache_arr_2_25, d_arr_2_24=>d_cache_arr_2_24, d_arr_2_23=>
      d_cache_arr_2_23, d_arr_2_22=>d_cache_arr_2_22, d_arr_2_21=>
      d_cache_arr_2_21, d_arr_2_20=>d_cache_arr_2_20, d_arr_2_19=>
      d_cache_arr_2_19, d_arr_2_18=>d_cache_arr_2_18, d_arr_2_17=>
      d_cache_arr_2_17, d_arr_2_16=>d_cache_arr_2_16, d_arr_2_15=>
      d_cache_arr_2_15, d_arr_2_14=>d_cache_arr_2_14, d_arr_2_13=>
      d_cache_arr_2_13, d_arr_2_12=>d_cache_arr_2_12, d_arr_2_11=>
      d_cache_arr_2_11, d_arr_2_10=>d_cache_arr_2_10, d_arr_2_9=>
      d_cache_arr_2_9, d_arr_2_8=>d_cache_arr_2_8, d_arr_2_7=>
      d_cache_arr_2_7, d_arr_2_6=>d_cache_arr_2_6, d_arr_2_5=>
      d_cache_arr_2_5, d_arr_2_4=>d_cache_arr_2_4, d_arr_2_3=>
      d_cache_arr_2_3, d_arr_2_2=>d_cache_arr_2_2, d_arr_2_1=>
      d_cache_arr_2_1, d_arr_2_0=>d_cache_arr_2_0, d_arr_3_31=>
      d_cache_arr_3_31, d_arr_3_30=>d_cache_arr_3_30, d_arr_3_29=>
      d_cache_arr_3_29, d_arr_3_28=>d_cache_arr_3_28, d_arr_3_27=>
      d_cache_arr_3_27, d_arr_3_26=>d_cache_arr_3_26, d_arr_3_25=>
      d_cache_arr_3_25, d_arr_3_24=>d_cache_arr_3_24, d_arr_3_23=>
      d_cache_arr_3_23, d_arr_3_22=>d_cache_arr_3_22, d_arr_3_21=>
      d_cache_arr_3_21, d_arr_3_20=>d_cache_arr_3_20, d_arr_3_19=>
      d_cache_arr_3_19, d_arr_3_18=>d_cache_arr_3_18, d_arr_3_17=>
      d_cache_arr_3_17, d_arr_3_16=>d_cache_arr_3_16, d_arr_3_15=>
      d_cache_arr_3_15, d_arr_3_14=>d_cache_arr_3_14, d_arr_3_13=>
      d_cache_arr_3_13, d_arr_3_12=>d_cache_arr_3_12, d_arr_3_11=>
      d_cache_arr_3_11, d_arr_3_10=>d_cache_arr_3_10, d_arr_3_9=>
      d_cache_arr_3_9, d_arr_3_8=>d_cache_arr_3_8, d_arr_3_7=>
      d_cache_arr_3_7, d_arr_3_6=>d_cache_arr_3_6, d_arr_3_5=>
      d_cache_arr_3_5, d_arr_3_4=>d_cache_arr_3_4, d_arr_3_3=>
      d_cache_arr_3_3, d_arr_3_2=>d_cache_arr_3_2, d_arr_3_1=>
      d_cache_arr_3_1, d_arr_3_0=>d_cache_arr_3_0, d_arr_4_31=>
      d_cache_arr_4_31, d_arr_4_30=>d_cache_arr_4_30, d_arr_4_29=>
      d_cache_arr_4_29, d_arr_4_28=>d_cache_arr_4_28, d_arr_4_27=>
      d_cache_arr_4_27, d_arr_4_26=>d_cache_arr_4_26, d_arr_4_25=>
      d_cache_arr_4_25, d_arr_4_24=>d_cache_arr_4_24, d_arr_4_23=>
      d_cache_arr_4_23, d_arr_4_22=>d_cache_arr_4_22, d_arr_4_21=>
      d_cache_arr_4_21, d_arr_4_20=>d_cache_arr_4_20, d_arr_4_19=>
      d_cache_arr_4_19, d_arr_4_18=>d_cache_arr_4_18, d_arr_4_17=>
      d_cache_arr_4_17, d_arr_4_16=>d_cache_arr_4_16, d_arr_4_15=>
      d_cache_arr_4_15, d_arr_4_14=>d_cache_arr_4_14, d_arr_4_13=>
      d_cache_arr_4_13, d_arr_4_12=>d_cache_arr_4_12, d_arr_4_11=>
      d_cache_arr_4_11, d_arr_4_10=>d_cache_arr_4_10, d_arr_4_9=>
      d_cache_arr_4_9, d_arr_4_8=>d_cache_arr_4_8, d_arr_4_7=>
      d_cache_arr_4_7, d_arr_4_6=>d_cache_arr_4_6, d_arr_4_5=>
      d_cache_arr_4_5, d_arr_4_4=>d_cache_arr_4_4, d_arr_4_3=>
      d_cache_arr_4_3, d_arr_4_2=>d_cache_arr_4_2, d_arr_4_1=>
      d_cache_arr_4_1, d_arr_4_0=>d_cache_arr_4_0, d_arr_5_31=>
      d_cache_arr_5_31, d_arr_5_30=>d_cache_arr_5_30, d_arr_5_29=>
      d_cache_arr_5_29, d_arr_5_28=>d_cache_arr_5_28, d_arr_5_27=>
      d_cache_arr_5_27, d_arr_5_26=>d_cache_arr_5_26, d_arr_5_25=>
      d_cache_arr_5_25, d_arr_5_24=>d_cache_arr_5_24, d_arr_5_23=>
      d_cache_arr_5_23, d_arr_5_22=>d_cache_arr_5_22, d_arr_5_21=>
      d_cache_arr_5_21, d_arr_5_20=>d_cache_arr_5_20, d_arr_5_19=>
      d_cache_arr_5_19, d_arr_5_18=>d_cache_arr_5_18, d_arr_5_17=>
      d_cache_arr_5_17, d_arr_5_16=>d_cache_arr_5_16, d_arr_5_15=>
      d_cache_arr_5_15, d_arr_5_14=>d_cache_arr_5_14, d_arr_5_13=>
      d_cache_arr_5_13, d_arr_5_12=>d_cache_arr_5_12, d_arr_5_11=>
      d_cache_arr_5_11, d_arr_5_10=>d_cache_arr_5_10, d_arr_5_9=>
      d_cache_arr_5_9, d_arr_5_8=>d_cache_arr_5_8, d_arr_5_7=>
      d_cache_arr_5_7, d_arr_5_6=>d_cache_arr_5_6, d_arr_5_5=>
      d_cache_arr_5_5, d_arr_5_4=>d_cache_arr_5_4, d_arr_5_3=>
      d_cache_arr_5_3, d_arr_5_2=>d_cache_arr_5_2, d_arr_5_1=>
      d_cache_arr_5_1, d_arr_5_0=>d_cache_arr_5_0, d_arr_6_31=>
      d_cache_arr_6_31, d_arr_6_30=>d_cache_arr_6_30, d_arr_6_29=>
      d_cache_arr_6_29, d_arr_6_28=>d_cache_arr_6_28, d_arr_6_27=>
      d_cache_arr_6_27, d_arr_6_26=>d_cache_arr_6_26, d_arr_6_25=>
      d_cache_arr_6_25, d_arr_6_24=>d_cache_arr_6_24, d_arr_6_23=>
      d_cache_arr_6_23, d_arr_6_22=>d_cache_arr_6_22, d_arr_6_21=>
      d_cache_arr_6_21, d_arr_6_20=>d_cache_arr_6_20, d_arr_6_19=>
      d_cache_arr_6_19, d_arr_6_18=>d_cache_arr_6_18, d_arr_6_17=>
      d_cache_arr_6_17, d_arr_6_16=>d_cache_arr_6_16, d_arr_6_15=>
      d_cache_arr_6_15, d_arr_6_14=>d_cache_arr_6_14, d_arr_6_13=>
      d_cache_arr_6_13, d_arr_6_12=>d_cache_arr_6_12, d_arr_6_11=>
      d_cache_arr_6_11, d_arr_6_10=>d_cache_arr_6_10, d_arr_6_9=>
      d_cache_arr_6_9, d_arr_6_8=>d_cache_arr_6_8, d_arr_6_7=>
      d_cache_arr_6_7, d_arr_6_6=>d_cache_arr_6_6, d_arr_6_5=>
      d_cache_arr_6_5, d_arr_6_4=>d_cache_arr_6_4, d_arr_6_3=>
      d_cache_arr_6_3, d_arr_6_2=>d_cache_arr_6_2, d_arr_6_1=>
      d_cache_arr_6_1, d_arr_6_0=>d_cache_arr_6_0, d_arr_7_31=>
      d_cache_arr_7_31, d_arr_7_30=>d_cache_arr_7_30, d_arr_7_29=>
      d_cache_arr_7_29, d_arr_7_28=>d_cache_arr_7_28, d_arr_7_27=>
      d_cache_arr_7_27, d_arr_7_26=>d_cache_arr_7_26, d_arr_7_25=>
      d_cache_arr_7_25, d_arr_7_24=>d_cache_arr_7_24, d_arr_7_23=>
      d_cache_arr_7_23, d_arr_7_22=>d_cache_arr_7_22, d_arr_7_21=>
      d_cache_arr_7_21, d_arr_7_20=>d_cache_arr_7_20, d_arr_7_19=>
      d_cache_arr_7_19, d_arr_7_18=>d_cache_arr_7_18, d_arr_7_17=>
      d_cache_arr_7_17, d_arr_7_16=>d_cache_arr_7_16, d_arr_7_15=>
      d_cache_arr_7_15, d_arr_7_14=>d_cache_arr_7_14, d_arr_7_13=>
      d_cache_arr_7_13, d_arr_7_12=>d_cache_arr_7_12, d_arr_7_11=>
      d_cache_arr_7_11, d_arr_7_10=>d_cache_arr_7_10, d_arr_7_9=>
      d_cache_arr_7_9, d_arr_7_8=>d_cache_arr_7_8, d_arr_7_7=>
      d_cache_arr_7_7, d_arr_7_6=>d_cache_arr_7_6, d_arr_7_5=>
      d_cache_arr_7_5, d_arr_7_4=>d_cache_arr_7_4, d_arr_7_3=>
      d_cache_arr_7_3, d_arr_7_2=>d_cache_arr_7_2, d_arr_7_1=>
      d_cache_arr_7_1, d_arr_7_0=>d_cache_arr_7_0, d_arr_8_31=>
      d_cache_arr_8_31, d_arr_8_30=>d_cache_arr_8_30, d_arr_8_29=>
      d_cache_arr_8_29, d_arr_8_28=>d_cache_arr_8_28, d_arr_8_27=>
      d_cache_arr_8_27, d_arr_8_26=>d_cache_arr_8_26, d_arr_8_25=>
      d_cache_arr_8_25, d_arr_8_24=>d_cache_arr_8_24, d_arr_8_23=>
      d_cache_arr_8_23, d_arr_8_22=>d_cache_arr_8_22, d_arr_8_21=>
      d_cache_arr_8_21, d_arr_8_20=>d_cache_arr_8_20, d_arr_8_19=>
      d_cache_arr_8_19, d_arr_8_18=>d_cache_arr_8_18, d_arr_8_17=>
      d_cache_arr_8_17, d_arr_8_16=>d_cache_arr_8_16, d_arr_8_15=>
      d_cache_arr_8_15, d_arr_8_14=>d_cache_arr_8_14, d_arr_8_13=>
      d_cache_arr_8_13, d_arr_8_12=>d_cache_arr_8_12, d_arr_8_11=>
      d_cache_arr_8_11, d_arr_8_10=>d_cache_arr_8_10, d_arr_8_9=>
      d_cache_arr_8_9, d_arr_8_8=>d_cache_arr_8_8, d_arr_8_7=>
      d_cache_arr_8_7, d_arr_8_6=>d_cache_arr_8_6, d_arr_8_5=>
      d_cache_arr_8_5, d_arr_8_4=>d_cache_arr_8_4, d_arr_8_3=>
      d_cache_arr_8_3, d_arr_8_2=>d_cache_arr_8_2, d_arr_8_1=>
      d_cache_arr_8_1, d_arr_8_0=>d_cache_arr_8_0, d_arr_9_31=>
      d_cache_arr_9_31, d_arr_9_30=>d_cache_arr_9_30, d_arr_9_29=>
      d_cache_arr_9_29, d_arr_9_28=>d_cache_arr_9_28, d_arr_9_27=>
      d_cache_arr_9_27, d_arr_9_26=>d_cache_arr_9_26, d_arr_9_25=>
      d_cache_arr_9_25, d_arr_9_24=>d_cache_arr_9_24, d_arr_9_23=>
      d_cache_arr_9_23, d_arr_9_22=>d_cache_arr_9_22, d_arr_9_21=>
      d_cache_arr_9_21, d_arr_9_20=>d_cache_arr_9_20, d_arr_9_19=>
      d_cache_arr_9_19, d_arr_9_18=>d_cache_arr_9_18, d_arr_9_17=>
      d_cache_arr_9_17, d_arr_9_16=>d_cache_arr_9_16, d_arr_9_15=>
      d_cache_arr_9_15, d_arr_9_14=>d_cache_arr_9_14, d_arr_9_13=>
      d_cache_arr_9_13, d_arr_9_12=>d_cache_arr_9_12, d_arr_9_11=>
      d_cache_arr_9_11, d_arr_9_10=>d_cache_arr_9_10, d_arr_9_9=>
      d_cache_arr_9_9, d_arr_9_8=>d_cache_arr_9_8, d_arr_9_7=>
      d_cache_arr_9_7, d_arr_9_6=>d_cache_arr_9_6, d_arr_9_5=>
      d_cache_arr_9_5, d_arr_9_4=>d_cache_arr_9_4, d_arr_9_3=>
      d_cache_arr_9_3, d_arr_9_2=>d_cache_arr_9_2, d_arr_9_1=>
      d_cache_arr_9_1, d_arr_9_0=>d_cache_arr_9_0, d_arr_10_31=>
      d_cache_arr_10_31, d_arr_10_30=>d_cache_arr_10_30, d_arr_10_29=>
      d_cache_arr_10_29, d_arr_10_28=>d_cache_arr_10_28, d_arr_10_27=>
      d_cache_arr_10_27, d_arr_10_26=>d_cache_arr_10_26, d_arr_10_25=>
      d_cache_arr_10_25, d_arr_10_24=>d_cache_arr_10_24, d_arr_10_23=>
      d_cache_arr_10_23, d_arr_10_22=>d_cache_arr_10_22, d_arr_10_21=>
      d_cache_arr_10_21, d_arr_10_20=>d_cache_arr_10_20, d_arr_10_19=>
      d_cache_arr_10_19, d_arr_10_18=>d_cache_arr_10_18, d_arr_10_17=>
      d_cache_arr_10_17, d_arr_10_16=>d_cache_arr_10_16, d_arr_10_15=>
      d_cache_arr_10_15, d_arr_10_14=>d_cache_arr_10_14, d_arr_10_13=>
      d_cache_arr_10_13, d_arr_10_12=>d_cache_arr_10_12, d_arr_10_11=>
      d_cache_arr_10_11, d_arr_10_10=>d_cache_arr_10_10, d_arr_10_9=>
      d_cache_arr_10_9, d_arr_10_8=>d_cache_arr_10_8, d_arr_10_7=>
      d_cache_arr_10_7, d_arr_10_6=>d_cache_arr_10_6, d_arr_10_5=>
      d_cache_arr_10_5, d_arr_10_4=>d_cache_arr_10_4, d_arr_10_3=>
      d_cache_arr_10_3, d_arr_10_2=>d_cache_arr_10_2, d_arr_10_1=>
      d_cache_arr_10_1, d_arr_10_0=>d_cache_arr_10_0, d_arr_11_31=>
      d_cache_arr_11_31, d_arr_11_30=>d_cache_arr_11_30, d_arr_11_29=>
      d_cache_arr_11_29, d_arr_11_28=>d_cache_arr_11_28, d_arr_11_27=>
      d_cache_arr_11_27, d_arr_11_26=>d_cache_arr_11_26, d_arr_11_25=>
      d_cache_arr_11_25, d_arr_11_24=>d_cache_arr_11_24, d_arr_11_23=>
      d_cache_arr_11_23, d_arr_11_22=>d_cache_arr_11_22, d_arr_11_21=>
      d_cache_arr_11_21, d_arr_11_20=>d_cache_arr_11_20, d_arr_11_19=>
      d_cache_arr_11_19, d_arr_11_18=>d_cache_arr_11_18, d_arr_11_17=>
      d_cache_arr_11_17, d_arr_11_16=>d_cache_arr_11_16, d_arr_11_15=>
      d_cache_arr_11_15, d_arr_11_14=>d_cache_arr_11_14, d_arr_11_13=>
      d_cache_arr_11_13, d_arr_11_12=>d_cache_arr_11_12, d_arr_11_11=>
      d_cache_arr_11_11, d_arr_11_10=>d_cache_arr_11_10, d_arr_11_9=>
      d_cache_arr_11_9, d_arr_11_8=>d_cache_arr_11_8, d_arr_11_7=>
      d_cache_arr_11_7, d_arr_11_6=>d_cache_arr_11_6, d_arr_11_5=>
      d_cache_arr_11_5, d_arr_11_4=>d_cache_arr_11_4, d_arr_11_3=>
      d_cache_arr_11_3, d_arr_11_2=>d_cache_arr_11_2, d_arr_11_1=>
      d_cache_arr_11_1, d_arr_11_0=>d_cache_arr_11_0, d_arr_12_31=>
      d_cache_arr_12_31, d_arr_12_30=>d_cache_arr_12_30, d_arr_12_29=>
      d_cache_arr_12_29, d_arr_12_28=>d_cache_arr_12_28, d_arr_12_27=>
      d_cache_arr_12_27, d_arr_12_26=>d_cache_arr_12_26, d_arr_12_25=>
      d_cache_arr_12_25, d_arr_12_24=>d_cache_arr_12_24, d_arr_12_23=>
      d_cache_arr_12_23, d_arr_12_22=>d_cache_arr_12_22, d_arr_12_21=>
      d_cache_arr_12_21, d_arr_12_20=>d_cache_arr_12_20, d_arr_12_19=>
      d_cache_arr_12_19, d_arr_12_18=>d_cache_arr_12_18, d_arr_12_17=>
      d_cache_arr_12_17, d_arr_12_16=>d_cache_arr_12_16, d_arr_12_15=>
      d_cache_arr_12_15, d_arr_12_14=>d_cache_arr_12_14, d_arr_12_13=>
      d_cache_arr_12_13, d_arr_12_12=>d_cache_arr_12_12, d_arr_12_11=>
      d_cache_arr_12_11, d_arr_12_10=>d_cache_arr_12_10, d_arr_12_9=>
      d_cache_arr_12_9, d_arr_12_8=>d_cache_arr_12_8, d_arr_12_7=>
      d_cache_arr_12_7, d_arr_12_6=>d_cache_arr_12_6, d_arr_12_5=>
      d_cache_arr_12_5, d_arr_12_4=>d_cache_arr_12_4, d_arr_12_3=>
      d_cache_arr_12_3, d_arr_12_2=>d_cache_arr_12_2, d_arr_12_1=>
      d_cache_arr_12_1, d_arr_12_0=>d_cache_arr_12_0, d_arr_13_31=>
      d_cache_arr_13_31, d_arr_13_30=>d_cache_arr_13_30, d_arr_13_29=>
      d_cache_arr_13_29, d_arr_13_28=>d_cache_arr_13_28, d_arr_13_27=>
      d_cache_arr_13_27, d_arr_13_26=>d_cache_arr_13_26, d_arr_13_25=>
      d_cache_arr_13_25, d_arr_13_24=>d_cache_arr_13_24, d_arr_13_23=>
      d_cache_arr_13_23, d_arr_13_22=>d_cache_arr_13_22, d_arr_13_21=>
      d_cache_arr_13_21, d_arr_13_20=>d_cache_arr_13_20, d_arr_13_19=>
      d_cache_arr_13_19, d_arr_13_18=>d_cache_arr_13_18, d_arr_13_17=>
      d_cache_arr_13_17, d_arr_13_16=>d_cache_arr_13_16, d_arr_13_15=>
      d_cache_arr_13_15, d_arr_13_14=>d_cache_arr_13_14, d_arr_13_13=>
      d_cache_arr_13_13, d_arr_13_12=>d_cache_arr_13_12, d_arr_13_11=>
      d_cache_arr_13_11, d_arr_13_10=>d_cache_arr_13_10, d_arr_13_9=>
      d_cache_arr_13_9, d_arr_13_8=>d_cache_arr_13_8, d_arr_13_7=>
      d_cache_arr_13_7, d_arr_13_6=>d_cache_arr_13_6, d_arr_13_5=>
      d_cache_arr_13_5, d_arr_13_4=>d_cache_arr_13_4, d_arr_13_3=>
      d_cache_arr_13_3, d_arr_13_2=>d_cache_arr_13_2, d_arr_13_1=>
      d_cache_arr_13_1, d_arr_13_0=>d_cache_arr_13_0, d_arr_14_31=>
      d_cache_arr_14_31, d_arr_14_30=>d_cache_arr_14_30, d_arr_14_29=>
      d_cache_arr_14_29, d_arr_14_28=>d_cache_arr_14_28, d_arr_14_27=>
      d_cache_arr_14_27, d_arr_14_26=>d_cache_arr_14_26, d_arr_14_25=>
      d_cache_arr_14_25, d_arr_14_24=>d_cache_arr_14_24, d_arr_14_23=>
      d_cache_arr_14_23, d_arr_14_22=>d_cache_arr_14_22, d_arr_14_21=>
      d_cache_arr_14_21, d_arr_14_20=>d_cache_arr_14_20, d_arr_14_19=>
      d_cache_arr_14_19, d_arr_14_18=>d_cache_arr_14_18, d_arr_14_17=>
      d_cache_arr_14_17, d_arr_14_16=>d_cache_arr_14_16, d_arr_14_15=>
      d_cache_arr_14_15, d_arr_14_14=>d_cache_arr_14_14, d_arr_14_13=>
      d_cache_arr_14_13, d_arr_14_12=>d_cache_arr_14_12, d_arr_14_11=>
      d_cache_arr_14_11, d_arr_14_10=>d_cache_arr_14_10, d_arr_14_9=>
      d_cache_arr_14_9, d_arr_14_8=>d_cache_arr_14_8, d_arr_14_7=>
      d_cache_arr_14_7, d_arr_14_6=>d_cache_arr_14_6, d_arr_14_5=>
      d_cache_arr_14_5, d_arr_14_4=>d_cache_arr_14_4, d_arr_14_3=>
      d_cache_arr_14_3, d_arr_14_2=>d_cache_arr_14_2, d_arr_14_1=>
      d_cache_arr_14_1, d_arr_14_0=>d_cache_arr_14_0, d_arr_15_31=>
      d_cache_arr_15_31, d_arr_15_30=>d_cache_arr_15_30, d_arr_15_29=>
      d_cache_arr_15_29, d_arr_15_28=>d_cache_arr_15_28, d_arr_15_27=>
      d_cache_arr_15_27, d_arr_15_26=>d_cache_arr_15_26, d_arr_15_25=>
      d_cache_arr_15_25, d_arr_15_24=>d_cache_arr_15_24, d_arr_15_23=>
      d_cache_arr_15_23, d_arr_15_22=>d_cache_arr_15_22, d_arr_15_21=>
      d_cache_arr_15_21, d_arr_15_20=>d_cache_arr_15_20, d_arr_15_19=>
      d_cache_arr_15_19, d_arr_15_18=>d_cache_arr_15_18, d_arr_15_17=>
      d_cache_arr_15_17, d_arr_15_16=>d_cache_arr_15_16, d_arr_15_15=>
      d_cache_arr_15_15, d_arr_15_14=>d_cache_arr_15_14, d_arr_15_13=>
      d_cache_arr_15_13, d_arr_15_12=>d_cache_arr_15_12, d_arr_15_11=>
      d_cache_arr_15_11, d_arr_15_10=>d_cache_arr_15_10, d_arr_15_9=>
      d_cache_arr_15_9, d_arr_15_8=>d_cache_arr_15_8, d_arr_15_7=>
      d_cache_arr_15_7, d_arr_15_6=>d_cache_arr_15_6, d_arr_15_5=>
      d_cache_arr_15_5, d_arr_15_4=>d_cache_arr_15_4, d_arr_15_3=>
      d_cache_arr_15_3, d_arr_15_2=>d_cache_arr_15_2, d_arr_15_1=>
      d_cache_arr_15_1, d_arr_15_0=>d_cache_arr_15_0, d_arr_16_31=>
      d_cache_arr_16_31, d_arr_16_30=>d_cache_arr_16_30, d_arr_16_29=>
      d_cache_arr_16_29, d_arr_16_28=>d_cache_arr_16_28, d_arr_16_27=>
      d_cache_arr_16_27, d_arr_16_26=>d_cache_arr_16_26, d_arr_16_25=>
      d_cache_arr_16_25, d_arr_16_24=>d_cache_arr_16_24, d_arr_16_23=>
      d_cache_arr_16_23, d_arr_16_22=>d_cache_arr_16_22, d_arr_16_21=>
      d_cache_arr_16_21, d_arr_16_20=>d_cache_arr_16_20, d_arr_16_19=>
      d_cache_arr_16_19, d_arr_16_18=>d_cache_arr_16_18, d_arr_16_17=>
      d_cache_arr_16_17, d_arr_16_16=>d_cache_arr_16_16, d_arr_16_15=>
      d_cache_arr_16_15, d_arr_16_14=>d_cache_arr_16_14, d_arr_16_13=>
      d_cache_arr_16_13, d_arr_16_12=>d_cache_arr_16_12, d_arr_16_11=>
      d_cache_arr_16_11, d_arr_16_10=>d_cache_arr_16_10, d_arr_16_9=>
      d_cache_arr_16_9, d_arr_16_8=>d_cache_arr_16_8, d_arr_16_7=>
      d_cache_arr_16_7, d_arr_16_6=>d_cache_arr_16_6, d_arr_16_5=>
      d_cache_arr_16_5, d_arr_16_4=>d_cache_arr_16_4, d_arr_16_3=>
      d_cache_arr_16_3, d_arr_16_2=>d_cache_arr_16_2, d_arr_16_1=>
      d_cache_arr_16_1, d_arr_16_0=>d_cache_arr_16_0, d_arr_17_31=>
      d_cache_arr_17_31, d_arr_17_30=>d_cache_arr_17_30, d_arr_17_29=>
      d_cache_arr_17_29, d_arr_17_28=>d_cache_arr_17_28, d_arr_17_27=>
      d_cache_arr_17_27, d_arr_17_26=>d_cache_arr_17_26, d_arr_17_25=>
      d_cache_arr_17_25, d_arr_17_24=>d_cache_arr_17_24, d_arr_17_23=>
      d_cache_arr_17_23, d_arr_17_22=>d_cache_arr_17_22, d_arr_17_21=>
      d_cache_arr_17_21, d_arr_17_20=>d_cache_arr_17_20, d_arr_17_19=>
      d_cache_arr_17_19, d_arr_17_18=>d_cache_arr_17_18, d_arr_17_17=>
      d_cache_arr_17_17, d_arr_17_16=>d_cache_arr_17_16, d_arr_17_15=>
      d_cache_arr_17_15, d_arr_17_14=>d_cache_arr_17_14, d_arr_17_13=>
      d_cache_arr_17_13, d_arr_17_12=>d_cache_arr_17_12, d_arr_17_11=>
      d_cache_arr_17_11, d_arr_17_10=>d_cache_arr_17_10, d_arr_17_9=>
      d_cache_arr_17_9, d_arr_17_8=>d_cache_arr_17_8, d_arr_17_7=>
      d_cache_arr_17_7, d_arr_17_6=>d_cache_arr_17_6, d_arr_17_5=>
      d_cache_arr_17_5, d_arr_17_4=>d_cache_arr_17_4, d_arr_17_3=>
      d_cache_arr_17_3, d_arr_17_2=>d_cache_arr_17_2, d_arr_17_1=>
      d_cache_arr_17_1, d_arr_17_0=>d_cache_arr_17_0, d_arr_18_31=>
      d_cache_arr_18_31, d_arr_18_30=>d_cache_arr_18_30, d_arr_18_29=>
      d_cache_arr_18_29, d_arr_18_28=>d_cache_arr_18_28, d_arr_18_27=>
      d_cache_arr_18_27, d_arr_18_26=>d_cache_arr_18_26, d_arr_18_25=>
      d_cache_arr_18_25, d_arr_18_24=>d_cache_arr_18_24, d_arr_18_23=>
      d_cache_arr_18_23, d_arr_18_22=>d_cache_arr_18_22, d_arr_18_21=>
      d_cache_arr_18_21, d_arr_18_20=>d_cache_arr_18_20, d_arr_18_19=>
      d_cache_arr_18_19, d_arr_18_18=>d_cache_arr_18_18, d_arr_18_17=>
      d_cache_arr_18_17, d_arr_18_16=>d_cache_arr_18_16, d_arr_18_15=>
      d_cache_arr_18_15, d_arr_18_14=>d_cache_arr_18_14, d_arr_18_13=>
      d_cache_arr_18_13, d_arr_18_12=>d_cache_arr_18_12, d_arr_18_11=>
      d_cache_arr_18_11, d_arr_18_10=>d_cache_arr_18_10, d_arr_18_9=>
      d_cache_arr_18_9, d_arr_18_8=>d_cache_arr_18_8, d_arr_18_7=>
      d_cache_arr_18_7, d_arr_18_6=>d_cache_arr_18_6, d_arr_18_5=>
      d_cache_arr_18_5, d_arr_18_4=>d_cache_arr_18_4, d_arr_18_3=>
      d_cache_arr_18_3, d_arr_18_2=>d_cache_arr_18_2, d_arr_18_1=>
      d_cache_arr_18_1, d_arr_18_0=>d_cache_arr_18_0, d_arr_19_31=>
      d_cache_arr_19_31, d_arr_19_30=>d_cache_arr_19_30, d_arr_19_29=>
      d_cache_arr_19_29, d_arr_19_28=>d_cache_arr_19_28, d_arr_19_27=>
      d_cache_arr_19_27, d_arr_19_26=>d_cache_arr_19_26, d_arr_19_25=>
      d_cache_arr_19_25, d_arr_19_24=>d_cache_arr_19_24, d_arr_19_23=>
      d_cache_arr_19_23, d_arr_19_22=>d_cache_arr_19_22, d_arr_19_21=>
      d_cache_arr_19_21, d_arr_19_20=>d_cache_arr_19_20, d_arr_19_19=>
      d_cache_arr_19_19, d_arr_19_18=>d_cache_arr_19_18, d_arr_19_17=>
      d_cache_arr_19_17, d_arr_19_16=>d_cache_arr_19_16, d_arr_19_15=>
      d_cache_arr_19_15, d_arr_19_14=>d_cache_arr_19_14, d_arr_19_13=>
      d_cache_arr_19_13, d_arr_19_12=>d_cache_arr_19_12, d_arr_19_11=>
      d_cache_arr_19_11, d_arr_19_10=>d_cache_arr_19_10, d_arr_19_9=>
      d_cache_arr_19_9, d_arr_19_8=>d_cache_arr_19_8, d_arr_19_7=>
      d_cache_arr_19_7, d_arr_19_6=>d_cache_arr_19_6, d_arr_19_5=>
      d_cache_arr_19_5, d_arr_19_4=>d_cache_arr_19_4, d_arr_19_3=>
      d_cache_arr_19_3, d_arr_19_2=>d_cache_arr_19_2, d_arr_19_1=>
      d_cache_arr_19_1, d_arr_19_0=>d_cache_arr_19_0, d_arr_20_31=>
      d_cache_arr_20_31, d_arr_20_30=>d_cache_arr_20_30, d_arr_20_29=>
      d_cache_arr_20_29, d_arr_20_28=>d_cache_arr_20_28, d_arr_20_27=>
      d_cache_arr_20_27, d_arr_20_26=>d_cache_arr_20_26, d_arr_20_25=>
      d_cache_arr_20_25, d_arr_20_24=>d_cache_arr_20_24, d_arr_20_23=>
      d_cache_arr_20_23, d_arr_20_22=>d_cache_arr_20_22, d_arr_20_21=>
      d_cache_arr_20_21, d_arr_20_20=>d_cache_arr_20_20, d_arr_20_19=>
      d_cache_arr_20_19, d_arr_20_18=>d_cache_arr_20_18, d_arr_20_17=>
      d_cache_arr_20_17, d_arr_20_16=>d_cache_arr_20_16, d_arr_20_15=>
      d_cache_arr_20_15, d_arr_20_14=>d_cache_arr_20_14, d_arr_20_13=>
      d_cache_arr_20_13, d_arr_20_12=>d_cache_arr_20_12, d_arr_20_11=>
      d_cache_arr_20_11, d_arr_20_10=>d_cache_arr_20_10, d_arr_20_9=>
      d_cache_arr_20_9, d_arr_20_8=>d_cache_arr_20_8, d_arr_20_7=>
      d_cache_arr_20_7, d_arr_20_6=>d_cache_arr_20_6, d_arr_20_5=>
      d_cache_arr_20_5, d_arr_20_4=>d_cache_arr_20_4, d_arr_20_3=>
      d_cache_arr_20_3, d_arr_20_2=>d_cache_arr_20_2, d_arr_20_1=>
      d_cache_arr_20_1, d_arr_20_0=>d_cache_arr_20_0, d_arr_21_31=>
      d_cache_arr_21_31, d_arr_21_30=>d_cache_arr_21_30, d_arr_21_29=>
      d_cache_arr_21_29, d_arr_21_28=>d_cache_arr_21_28, d_arr_21_27=>
      d_cache_arr_21_27, d_arr_21_26=>d_cache_arr_21_26, d_arr_21_25=>
      d_cache_arr_21_25, d_arr_21_24=>d_cache_arr_21_24, d_arr_21_23=>
      d_cache_arr_21_23, d_arr_21_22=>d_cache_arr_21_22, d_arr_21_21=>
      d_cache_arr_21_21, d_arr_21_20=>d_cache_arr_21_20, d_arr_21_19=>
      d_cache_arr_21_19, d_arr_21_18=>d_cache_arr_21_18, d_arr_21_17=>
      d_cache_arr_21_17, d_arr_21_16=>d_cache_arr_21_16, d_arr_21_15=>
      d_cache_arr_21_15, d_arr_21_14=>d_cache_arr_21_14, d_arr_21_13=>
      d_cache_arr_21_13, d_arr_21_12=>d_cache_arr_21_12, d_arr_21_11=>
      d_cache_arr_21_11, d_arr_21_10=>d_cache_arr_21_10, d_arr_21_9=>
      d_cache_arr_21_9, d_arr_21_8=>d_cache_arr_21_8, d_arr_21_7=>
      d_cache_arr_21_7, d_arr_21_6=>d_cache_arr_21_6, d_arr_21_5=>
      d_cache_arr_21_5, d_arr_21_4=>d_cache_arr_21_4, d_arr_21_3=>
      d_cache_arr_21_3, d_arr_21_2=>d_cache_arr_21_2, d_arr_21_1=>
      d_cache_arr_21_1, d_arr_21_0=>d_cache_arr_21_0, d_arr_22_31=>
      d_cache_arr_22_31, d_arr_22_30=>d_cache_arr_22_30, d_arr_22_29=>
      d_cache_arr_22_29, d_arr_22_28=>d_cache_arr_22_28, d_arr_22_27=>
      d_cache_arr_22_27, d_arr_22_26=>d_cache_arr_22_26, d_arr_22_25=>
      d_cache_arr_22_25, d_arr_22_24=>d_cache_arr_22_24, d_arr_22_23=>
      d_cache_arr_22_23, d_arr_22_22=>d_cache_arr_22_22, d_arr_22_21=>
      d_cache_arr_22_21, d_arr_22_20=>d_cache_arr_22_20, d_arr_22_19=>
      d_cache_arr_22_19, d_arr_22_18=>d_cache_arr_22_18, d_arr_22_17=>
      d_cache_arr_22_17, d_arr_22_16=>d_cache_arr_22_16, d_arr_22_15=>
      d_cache_arr_22_15, d_arr_22_14=>d_cache_arr_22_14, d_arr_22_13=>
      d_cache_arr_22_13, d_arr_22_12=>d_cache_arr_22_12, d_arr_22_11=>
      d_cache_arr_22_11, d_arr_22_10=>d_cache_arr_22_10, d_arr_22_9=>
      d_cache_arr_22_9, d_arr_22_8=>d_cache_arr_22_8, d_arr_22_7=>
      d_cache_arr_22_7, d_arr_22_6=>d_cache_arr_22_6, d_arr_22_5=>
      d_cache_arr_22_5, d_arr_22_4=>d_cache_arr_22_4, d_arr_22_3=>
      d_cache_arr_22_3, d_arr_22_2=>d_cache_arr_22_2, d_arr_22_1=>
      d_cache_arr_22_1, d_arr_22_0=>d_cache_arr_22_0, d_arr_23_31=>
      d_cache_arr_23_31, d_arr_23_30=>d_cache_arr_23_30, d_arr_23_29=>
      d_cache_arr_23_29, d_arr_23_28=>d_cache_arr_23_28, d_arr_23_27=>
      d_cache_arr_23_27, d_arr_23_26=>d_cache_arr_23_26, d_arr_23_25=>
      d_cache_arr_23_25, d_arr_23_24=>d_cache_arr_23_24, d_arr_23_23=>
      d_cache_arr_23_23, d_arr_23_22=>d_cache_arr_23_22, d_arr_23_21=>
      d_cache_arr_23_21, d_arr_23_20=>d_cache_arr_23_20, d_arr_23_19=>
      d_cache_arr_23_19, d_arr_23_18=>d_cache_arr_23_18, d_arr_23_17=>
      d_cache_arr_23_17, d_arr_23_16=>d_cache_arr_23_16, d_arr_23_15=>
      d_cache_arr_23_15, d_arr_23_14=>d_cache_arr_23_14, d_arr_23_13=>
      d_cache_arr_23_13, d_arr_23_12=>d_cache_arr_23_12, d_arr_23_11=>
      d_cache_arr_23_11, d_arr_23_10=>d_cache_arr_23_10, d_arr_23_9=>
      d_cache_arr_23_9, d_arr_23_8=>d_cache_arr_23_8, d_arr_23_7=>
      d_cache_arr_23_7, d_arr_23_6=>d_cache_arr_23_6, d_arr_23_5=>
      d_cache_arr_23_5, d_arr_23_4=>d_cache_arr_23_4, d_arr_23_3=>
      d_cache_arr_23_3, d_arr_23_2=>d_cache_arr_23_2, d_arr_23_1=>
      d_cache_arr_23_1, d_arr_23_0=>d_cache_arr_23_0, d_arr_24_31=>
      d_cache_arr_24_31, d_arr_24_30=>d_cache_arr_24_30, d_arr_24_29=>
      d_cache_arr_24_29, d_arr_24_28=>d_cache_arr_24_28, d_arr_24_27=>
      d_cache_arr_24_27, d_arr_24_26=>d_cache_arr_24_26, d_arr_24_25=>
      d_cache_arr_24_25, d_arr_24_24=>d_cache_arr_24_24, d_arr_24_23=>
      d_cache_arr_24_23, d_arr_24_22=>d_cache_arr_24_22, d_arr_24_21=>
      d_cache_arr_24_21, d_arr_24_20=>d_cache_arr_24_20, d_arr_24_19=>
      d_cache_arr_24_19, d_arr_24_18=>d_cache_arr_24_18, d_arr_24_17=>
      d_cache_arr_24_17, d_arr_24_16=>d_cache_arr_24_16, d_arr_24_15=>
      d_cache_arr_24_15, d_arr_24_14=>d_cache_arr_24_14, d_arr_24_13=>
      d_cache_arr_24_13, d_arr_24_12=>d_cache_arr_24_12, d_arr_24_11=>
      d_cache_arr_24_11, d_arr_24_10=>d_cache_arr_24_10, d_arr_24_9=>
      d_cache_arr_24_9, d_arr_24_8=>d_cache_arr_24_8, d_arr_24_7=>
      d_cache_arr_24_7, d_arr_24_6=>d_cache_arr_24_6, d_arr_24_5=>
      d_cache_arr_24_5, d_arr_24_4=>d_cache_arr_24_4, d_arr_24_3=>
      d_cache_arr_24_3, d_arr_24_2=>d_cache_arr_24_2, d_arr_24_1=>
      d_cache_arr_24_1, d_arr_24_0=>d_cache_arr_24_0, q_arr_0_31=>
      q_cache_arr_0_31, q_arr_0_30=>q_cache_arr_0_30, q_arr_0_29=>
      q_cache_arr_0_29, q_arr_0_28=>q_cache_arr_0_28, q_arr_0_27=>
      q_cache_arr_0_27, q_arr_0_26=>q_cache_arr_0_26, q_arr_0_25=>
      q_cache_arr_0_25, q_arr_0_24=>q_cache_arr_0_24, q_arr_0_23=>
      q_cache_arr_0_23, q_arr_0_22=>q_cache_arr_0_22, q_arr_0_21=>
      q_cache_arr_0_21, q_arr_0_20=>q_cache_arr_0_20, q_arr_0_19=>
      q_cache_arr_0_19, q_arr_0_18=>q_cache_arr_0_18, q_arr_0_17=>
      q_cache_arr_0_17, q_arr_0_16=>q_cache_arr_0_16, q_arr_0_15=>
      q_cache_arr_0_15, q_arr_0_14=>q_cache_arr_0_14, q_arr_0_13=>
      q_cache_arr_0_13, q_arr_0_12=>q_cache_arr_0_12, q_arr_0_11=>
      q_cache_arr_0_11, q_arr_0_10=>q_cache_arr_0_10, q_arr_0_9=>
      q_cache_arr_0_9, q_arr_0_8=>q_cache_arr_0_8, q_arr_0_7=>
      q_cache_arr_0_7, q_arr_0_6=>q_cache_arr_0_6, q_arr_0_5=>
      q_cache_arr_0_5, q_arr_0_4=>q_cache_arr_0_4, q_arr_0_3=>
      q_cache_arr_0_3, q_arr_0_2=>q_cache_arr_0_2, q_arr_0_1=>
      q_cache_arr_0_1, q_arr_0_0=>q_cache_arr_0_0, q_arr_1_31=>
      q_cache_arr_1_31, q_arr_1_30=>q_cache_arr_1_30, q_arr_1_29=>
      q_cache_arr_1_29, q_arr_1_28=>q_cache_arr_1_28, q_arr_1_27=>
      q_cache_arr_1_27, q_arr_1_26=>q_cache_arr_1_26, q_arr_1_25=>
      q_cache_arr_1_25, q_arr_1_24=>q_cache_arr_1_24, q_arr_1_23=>
      q_cache_arr_1_23, q_arr_1_22=>q_cache_arr_1_22, q_arr_1_21=>
      q_cache_arr_1_21, q_arr_1_20=>q_cache_arr_1_20, q_arr_1_19=>
      q_cache_arr_1_19, q_arr_1_18=>q_cache_arr_1_18, q_arr_1_17=>
      q_cache_arr_1_17, q_arr_1_16=>q_cache_arr_1_16, q_arr_1_15=>
      q_cache_arr_1_15, q_arr_1_14=>q_cache_arr_1_14, q_arr_1_13=>
      q_cache_arr_1_13, q_arr_1_12=>q_cache_arr_1_12, q_arr_1_11=>
      q_cache_arr_1_11, q_arr_1_10=>q_cache_arr_1_10, q_arr_1_9=>
      q_cache_arr_1_9, q_arr_1_8=>q_cache_arr_1_8, q_arr_1_7=>
      q_cache_arr_1_7, q_arr_1_6=>q_cache_arr_1_6, q_arr_1_5=>
      q_cache_arr_1_5, q_arr_1_4=>q_cache_arr_1_4, q_arr_1_3=>
      q_cache_arr_1_3, q_arr_1_2=>q_cache_arr_1_2, q_arr_1_1=>
      q_cache_arr_1_1, q_arr_1_0=>q_cache_arr_1_0, q_arr_2_31=>
      q_cache_arr_2_31, q_arr_2_30=>q_cache_arr_2_30, q_arr_2_29=>
      q_cache_arr_2_29, q_arr_2_28=>q_cache_arr_2_28, q_arr_2_27=>
      q_cache_arr_2_27, q_arr_2_26=>q_cache_arr_2_26, q_arr_2_25=>
      q_cache_arr_2_25, q_arr_2_24=>q_cache_arr_2_24, q_arr_2_23=>
      q_cache_arr_2_23, q_arr_2_22=>q_cache_arr_2_22, q_arr_2_21=>
      q_cache_arr_2_21, q_arr_2_20=>q_cache_arr_2_20, q_arr_2_19=>
      q_cache_arr_2_19, q_arr_2_18=>q_cache_arr_2_18, q_arr_2_17=>
      q_cache_arr_2_17, q_arr_2_16=>q_cache_arr_2_16, q_arr_2_15=>
      q_cache_arr_2_15, q_arr_2_14=>q_cache_arr_2_14, q_arr_2_13=>
      q_cache_arr_2_13, q_arr_2_12=>q_cache_arr_2_12, q_arr_2_11=>
      q_cache_arr_2_11, q_arr_2_10=>q_cache_arr_2_10, q_arr_2_9=>
      q_cache_arr_2_9, q_arr_2_8=>q_cache_arr_2_8, q_arr_2_7=>
      q_cache_arr_2_7, q_arr_2_6=>q_cache_arr_2_6, q_arr_2_5=>
      q_cache_arr_2_5, q_arr_2_4=>q_cache_arr_2_4, q_arr_2_3=>
      q_cache_arr_2_3, q_arr_2_2=>q_cache_arr_2_2, q_arr_2_1=>
      q_cache_arr_2_1, q_arr_2_0=>q_cache_arr_2_0, q_arr_3_31=>
      q_cache_arr_3_31, q_arr_3_30=>q_cache_arr_3_30, q_arr_3_29=>
      q_cache_arr_3_29, q_arr_3_28=>q_cache_arr_3_28, q_arr_3_27=>
      q_cache_arr_3_27, q_arr_3_26=>q_cache_arr_3_26, q_arr_3_25=>
      q_cache_arr_3_25, q_arr_3_24=>q_cache_arr_3_24, q_arr_3_23=>
      q_cache_arr_3_23, q_arr_3_22=>q_cache_arr_3_22, q_arr_3_21=>
      q_cache_arr_3_21, q_arr_3_20=>q_cache_arr_3_20, q_arr_3_19=>
      q_cache_arr_3_19, q_arr_3_18=>q_cache_arr_3_18, q_arr_3_17=>
      q_cache_arr_3_17, q_arr_3_16=>q_cache_arr_3_16, q_arr_3_15=>
      q_cache_arr_3_15, q_arr_3_14=>q_cache_arr_3_14, q_arr_3_13=>
      q_cache_arr_3_13, q_arr_3_12=>q_cache_arr_3_12, q_arr_3_11=>
      q_cache_arr_3_11, q_arr_3_10=>q_cache_arr_3_10, q_arr_3_9=>
      q_cache_arr_3_9, q_arr_3_8=>q_cache_arr_3_8, q_arr_3_7=>
      q_cache_arr_3_7, q_arr_3_6=>q_cache_arr_3_6, q_arr_3_5=>
      q_cache_arr_3_5, q_arr_3_4=>q_cache_arr_3_4, q_arr_3_3=>
      q_cache_arr_3_3, q_arr_3_2=>q_cache_arr_3_2, q_arr_3_1=>
      q_cache_arr_3_1, q_arr_3_0=>q_cache_arr_3_0, q_arr_4_31=>
      q_cache_arr_4_31, q_arr_4_30=>q_cache_arr_4_30, q_arr_4_29=>
      q_cache_arr_4_29, q_arr_4_28=>q_cache_arr_4_28, q_arr_4_27=>
      q_cache_arr_4_27, q_arr_4_26=>q_cache_arr_4_26, q_arr_4_25=>
      q_cache_arr_4_25, q_arr_4_24=>q_cache_arr_4_24, q_arr_4_23=>
      q_cache_arr_4_23, q_arr_4_22=>q_cache_arr_4_22, q_arr_4_21=>
      q_cache_arr_4_21, q_arr_4_20=>q_cache_arr_4_20, q_arr_4_19=>
      q_cache_arr_4_19, q_arr_4_18=>q_cache_arr_4_18, q_arr_4_17=>
      q_cache_arr_4_17, q_arr_4_16=>q_cache_arr_4_16, q_arr_4_15=>
      q_cache_arr_4_15, q_arr_4_14=>q_cache_arr_4_14, q_arr_4_13=>
      q_cache_arr_4_13, q_arr_4_12=>q_cache_arr_4_12, q_arr_4_11=>
      q_cache_arr_4_11, q_arr_4_10=>q_cache_arr_4_10, q_arr_4_9=>
      q_cache_arr_4_9, q_arr_4_8=>q_cache_arr_4_8, q_arr_4_7=>
      q_cache_arr_4_7, q_arr_4_6=>q_cache_arr_4_6, q_arr_4_5=>
      q_cache_arr_4_5, q_arr_4_4=>q_cache_arr_4_4, q_arr_4_3=>
      q_cache_arr_4_3, q_arr_4_2=>q_cache_arr_4_2, q_arr_4_1=>
      q_cache_arr_4_1, q_arr_4_0=>q_cache_arr_4_0, q_arr_5_31=>
      q_cache_arr_5_31, q_arr_5_30=>q_cache_arr_5_30, q_arr_5_29=>
      q_cache_arr_5_29, q_arr_5_28=>q_cache_arr_5_28, q_arr_5_27=>
      q_cache_arr_5_27, q_arr_5_26=>q_cache_arr_5_26, q_arr_5_25=>
      q_cache_arr_5_25, q_arr_5_24=>q_cache_arr_5_24, q_arr_5_23=>
      q_cache_arr_5_23, q_arr_5_22=>q_cache_arr_5_22, q_arr_5_21=>
      q_cache_arr_5_21, q_arr_5_20=>q_cache_arr_5_20, q_arr_5_19=>
      q_cache_arr_5_19, q_arr_5_18=>q_cache_arr_5_18, q_arr_5_17=>
      q_cache_arr_5_17, q_arr_5_16=>q_cache_arr_5_16, q_arr_5_15=>
      q_cache_arr_5_15, q_arr_5_14=>q_cache_arr_5_14, q_arr_5_13=>
      q_cache_arr_5_13, q_arr_5_12=>q_cache_arr_5_12, q_arr_5_11=>
      q_cache_arr_5_11, q_arr_5_10=>q_cache_arr_5_10, q_arr_5_9=>
      q_cache_arr_5_9, q_arr_5_8=>q_cache_arr_5_8, q_arr_5_7=>
      q_cache_arr_5_7, q_arr_5_6=>q_cache_arr_5_6, q_arr_5_5=>
      q_cache_arr_5_5, q_arr_5_4=>q_cache_arr_5_4, q_arr_5_3=>
      q_cache_arr_5_3, q_arr_5_2=>q_cache_arr_5_2, q_arr_5_1=>
      q_cache_arr_5_1, q_arr_5_0=>q_cache_arr_5_0, q_arr_6_31=>
      q_cache_arr_6_31, q_arr_6_30=>q_cache_arr_6_30, q_arr_6_29=>
      q_cache_arr_6_29, q_arr_6_28=>q_cache_arr_6_28, q_arr_6_27=>
      q_cache_arr_6_27, q_arr_6_26=>q_cache_arr_6_26, q_arr_6_25=>
      q_cache_arr_6_25, q_arr_6_24=>q_cache_arr_6_24, q_arr_6_23=>
      q_cache_arr_6_23, q_arr_6_22=>q_cache_arr_6_22, q_arr_6_21=>
      q_cache_arr_6_21, q_arr_6_20=>q_cache_arr_6_20, q_arr_6_19=>
      q_cache_arr_6_19, q_arr_6_18=>q_cache_arr_6_18, q_arr_6_17=>
      q_cache_arr_6_17, q_arr_6_16=>q_cache_arr_6_16, q_arr_6_15=>
      q_cache_arr_6_15, q_arr_6_14=>q_cache_arr_6_14, q_arr_6_13=>
      q_cache_arr_6_13, q_arr_6_12=>q_cache_arr_6_12, q_arr_6_11=>
      q_cache_arr_6_11, q_arr_6_10=>q_cache_arr_6_10, q_arr_6_9=>
      q_cache_arr_6_9, q_arr_6_8=>q_cache_arr_6_8, q_arr_6_7=>
      q_cache_arr_6_7, q_arr_6_6=>q_cache_arr_6_6, q_arr_6_5=>
      q_cache_arr_6_5, q_arr_6_4=>q_cache_arr_6_4, q_arr_6_3=>
      q_cache_arr_6_3, q_arr_6_2=>q_cache_arr_6_2, q_arr_6_1=>
      q_cache_arr_6_1, q_arr_6_0=>q_cache_arr_6_0, q_arr_7_31=>
      q_cache_arr_7_31, q_arr_7_30=>q_cache_arr_7_30, q_arr_7_29=>
      q_cache_arr_7_29, q_arr_7_28=>q_cache_arr_7_28, q_arr_7_27=>
      q_cache_arr_7_27, q_arr_7_26=>q_cache_arr_7_26, q_arr_7_25=>
      q_cache_arr_7_25, q_arr_7_24=>q_cache_arr_7_24, q_arr_7_23=>
      q_cache_arr_7_23, q_arr_7_22=>q_cache_arr_7_22, q_arr_7_21=>
      q_cache_arr_7_21, q_arr_7_20=>q_cache_arr_7_20, q_arr_7_19=>
      q_cache_arr_7_19, q_arr_7_18=>q_cache_arr_7_18, q_arr_7_17=>
      q_cache_arr_7_17, q_arr_7_16=>q_cache_arr_7_16, q_arr_7_15=>
      q_cache_arr_7_15, q_arr_7_14=>q_cache_arr_7_14, q_arr_7_13=>
      q_cache_arr_7_13, q_arr_7_12=>q_cache_arr_7_12, q_arr_7_11=>
      q_cache_arr_7_11, q_arr_7_10=>q_cache_arr_7_10, q_arr_7_9=>
      q_cache_arr_7_9, q_arr_7_8=>q_cache_arr_7_8, q_arr_7_7=>
      q_cache_arr_7_7, q_arr_7_6=>q_cache_arr_7_6, q_arr_7_5=>
      q_cache_arr_7_5, q_arr_7_4=>q_cache_arr_7_4, q_arr_7_3=>
      q_cache_arr_7_3, q_arr_7_2=>q_cache_arr_7_2, q_arr_7_1=>
      q_cache_arr_7_1, q_arr_7_0=>q_cache_arr_7_0, q_arr_8_31=>
      q_cache_arr_8_31, q_arr_8_30=>q_cache_arr_8_30, q_arr_8_29=>
      q_cache_arr_8_29, q_arr_8_28=>q_cache_arr_8_28, q_arr_8_27=>
      q_cache_arr_8_27, q_arr_8_26=>q_cache_arr_8_26, q_arr_8_25=>
      q_cache_arr_8_25, q_arr_8_24=>q_cache_arr_8_24, q_arr_8_23=>
      q_cache_arr_8_23, q_arr_8_22=>q_cache_arr_8_22, q_arr_8_21=>
      q_cache_arr_8_21, q_arr_8_20=>q_cache_arr_8_20, q_arr_8_19=>
      q_cache_arr_8_19, q_arr_8_18=>q_cache_arr_8_18, q_arr_8_17=>
      q_cache_arr_8_17, q_arr_8_16=>q_cache_arr_8_16, q_arr_8_15=>
      q_cache_arr_8_15, q_arr_8_14=>q_cache_arr_8_14, q_arr_8_13=>
      q_cache_arr_8_13, q_arr_8_12=>q_cache_arr_8_12, q_arr_8_11=>
      q_cache_arr_8_11, q_arr_8_10=>q_cache_arr_8_10, q_arr_8_9=>
      q_cache_arr_8_9, q_arr_8_8=>q_cache_arr_8_8, q_arr_8_7=>
      q_cache_arr_8_7, q_arr_8_6=>q_cache_arr_8_6, q_arr_8_5=>
      q_cache_arr_8_5, q_arr_8_4=>q_cache_arr_8_4, q_arr_8_3=>
      q_cache_arr_8_3, q_arr_8_2=>q_cache_arr_8_2, q_arr_8_1=>
      q_cache_arr_8_1, q_arr_8_0=>q_cache_arr_8_0, q_arr_9_31=>
      q_cache_arr_9_31, q_arr_9_30=>q_cache_arr_9_30, q_arr_9_29=>
      q_cache_arr_9_29, q_arr_9_28=>q_cache_arr_9_28, q_arr_9_27=>
      q_cache_arr_9_27, q_arr_9_26=>q_cache_arr_9_26, q_arr_9_25=>
      q_cache_arr_9_25, q_arr_9_24=>q_cache_arr_9_24, q_arr_9_23=>
      q_cache_arr_9_23, q_arr_9_22=>q_cache_arr_9_22, q_arr_9_21=>
      q_cache_arr_9_21, q_arr_9_20=>q_cache_arr_9_20, q_arr_9_19=>
      q_cache_arr_9_19, q_arr_9_18=>q_cache_arr_9_18, q_arr_9_17=>
      q_cache_arr_9_17, q_arr_9_16=>q_cache_arr_9_16, q_arr_9_15=>
      q_cache_arr_9_15, q_arr_9_14=>q_cache_arr_9_14, q_arr_9_13=>
      q_cache_arr_9_13, q_arr_9_12=>q_cache_arr_9_12, q_arr_9_11=>
      q_cache_arr_9_11, q_arr_9_10=>q_cache_arr_9_10, q_arr_9_9=>
      q_cache_arr_9_9, q_arr_9_8=>q_cache_arr_9_8, q_arr_9_7=>
      q_cache_arr_9_7, q_arr_9_6=>q_cache_arr_9_6, q_arr_9_5=>
      q_cache_arr_9_5, q_arr_9_4=>q_cache_arr_9_4, q_arr_9_3=>
      q_cache_arr_9_3, q_arr_9_2=>q_cache_arr_9_2, q_arr_9_1=>
      q_cache_arr_9_1, q_arr_9_0=>q_cache_arr_9_0, q_arr_10_31=>
      q_cache_arr_10_31, q_arr_10_30=>q_cache_arr_10_30, q_arr_10_29=>
      q_cache_arr_10_29, q_arr_10_28=>q_cache_arr_10_28, q_arr_10_27=>
      q_cache_arr_10_27, q_arr_10_26=>q_cache_arr_10_26, q_arr_10_25=>
      q_cache_arr_10_25, q_arr_10_24=>q_cache_arr_10_24, q_arr_10_23=>
      q_cache_arr_10_23, q_arr_10_22=>q_cache_arr_10_22, q_arr_10_21=>
      q_cache_arr_10_21, q_arr_10_20=>q_cache_arr_10_20, q_arr_10_19=>
      q_cache_arr_10_19, q_arr_10_18=>q_cache_arr_10_18, q_arr_10_17=>
      q_cache_arr_10_17, q_arr_10_16=>q_cache_arr_10_16, q_arr_10_15=>
      q_cache_arr_10_15, q_arr_10_14=>q_cache_arr_10_14, q_arr_10_13=>
      q_cache_arr_10_13, q_arr_10_12=>q_cache_arr_10_12, q_arr_10_11=>
      q_cache_arr_10_11, q_arr_10_10=>q_cache_arr_10_10, q_arr_10_9=>
      q_cache_arr_10_9, q_arr_10_8=>q_cache_arr_10_8, q_arr_10_7=>
      q_cache_arr_10_7, q_arr_10_6=>q_cache_arr_10_6, q_arr_10_5=>
      q_cache_arr_10_5, q_arr_10_4=>q_cache_arr_10_4, q_arr_10_3=>
      q_cache_arr_10_3, q_arr_10_2=>q_cache_arr_10_2, q_arr_10_1=>
      q_cache_arr_10_1, q_arr_10_0=>q_cache_arr_10_0, q_arr_11_31=>
      q_cache_arr_11_31, q_arr_11_30=>q_cache_arr_11_30, q_arr_11_29=>
      q_cache_arr_11_29, q_arr_11_28=>q_cache_arr_11_28, q_arr_11_27=>
      q_cache_arr_11_27, q_arr_11_26=>q_cache_arr_11_26, q_arr_11_25=>
      q_cache_arr_11_25, q_arr_11_24=>q_cache_arr_11_24, q_arr_11_23=>
      q_cache_arr_11_23, q_arr_11_22=>q_cache_arr_11_22, q_arr_11_21=>
      q_cache_arr_11_21, q_arr_11_20=>q_cache_arr_11_20, q_arr_11_19=>
      q_cache_arr_11_19, q_arr_11_18=>q_cache_arr_11_18, q_arr_11_17=>
      q_cache_arr_11_17, q_arr_11_16=>q_cache_arr_11_16, q_arr_11_15=>
      q_cache_arr_11_15, q_arr_11_14=>q_cache_arr_11_14, q_arr_11_13=>
      q_cache_arr_11_13, q_arr_11_12=>q_cache_arr_11_12, q_arr_11_11=>
      q_cache_arr_11_11, q_arr_11_10=>q_cache_arr_11_10, q_arr_11_9=>
      q_cache_arr_11_9, q_arr_11_8=>q_cache_arr_11_8, q_arr_11_7=>
      q_cache_arr_11_7, q_arr_11_6=>q_cache_arr_11_6, q_arr_11_5=>
      q_cache_arr_11_5, q_arr_11_4=>q_cache_arr_11_4, q_arr_11_3=>
      q_cache_arr_11_3, q_arr_11_2=>q_cache_arr_11_2, q_arr_11_1=>
      q_cache_arr_11_1, q_arr_11_0=>q_cache_arr_11_0, q_arr_12_31=>
      q_cache_arr_12_31, q_arr_12_30=>q_cache_arr_12_30, q_arr_12_29=>
      q_cache_arr_12_29, q_arr_12_28=>q_cache_arr_12_28, q_arr_12_27=>
      q_cache_arr_12_27, q_arr_12_26=>q_cache_arr_12_26, q_arr_12_25=>
      q_cache_arr_12_25, q_arr_12_24=>q_cache_arr_12_24, q_arr_12_23=>
      q_cache_arr_12_23, q_arr_12_22=>q_cache_arr_12_22, q_arr_12_21=>
      q_cache_arr_12_21, q_arr_12_20=>q_cache_arr_12_20, q_arr_12_19=>
      q_cache_arr_12_19, q_arr_12_18=>q_cache_arr_12_18, q_arr_12_17=>
      q_cache_arr_12_17, q_arr_12_16=>q_cache_arr_12_16, q_arr_12_15=>
      q_cache_arr_12_15, q_arr_12_14=>q_cache_arr_12_14, q_arr_12_13=>
      q_cache_arr_12_13, q_arr_12_12=>q_cache_arr_12_12, q_arr_12_11=>
      q_cache_arr_12_11, q_arr_12_10=>q_cache_arr_12_10, q_arr_12_9=>
      q_cache_arr_12_9, q_arr_12_8=>q_cache_arr_12_8, q_arr_12_7=>
      q_cache_arr_12_7, q_arr_12_6=>q_cache_arr_12_6, q_arr_12_5=>
      q_cache_arr_12_5, q_arr_12_4=>q_cache_arr_12_4, q_arr_12_3=>
      q_cache_arr_12_3, q_arr_12_2=>q_cache_arr_12_2, q_arr_12_1=>
      q_cache_arr_12_1, q_arr_12_0=>q_cache_arr_12_0, q_arr_13_31=>
      q_cache_arr_13_31, q_arr_13_30=>q_cache_arr_13_30, q_arr_13_29=>
      q_cache_arr_13_29, q_arr_13_28=>q_cache_arr_13_28, q_arr_13_27=>
      q_cache_arr_13_27, q_arr_13_26=>q_cache_arr_13_26, q_arr_13_25=>
      q_cache_arr_13_25, q_arr_13_24=>q_cache_arr_13_24, q_arr_13_23=>
      q_cache_arr_13_23, q_arr_13_22=>q_cache_arr_13_22, q_arr_13_21=>
      q_cache_arr_13_21, q_arr_13_20=>q_cache_arr_13_20, q_arr_13_19=>
      q_cache_arr_13_19, q_arr_13_18=>q_cache_arr_13_18, q_arr_13_17=>
      q_cache_arr_13_17, q_arr_13_16=>q_cache_arr_13_16, q_arr_13_15=>
      q_cache_arr_13_15, q_arr_13_14=>q_cache_arr_13_14, q_arr_13_13=>
      q_cache_arr_13_13, q_arr_13_12=>q_cache_arr_13_12, q_arr_13_11=>
      q_cache_arr_13_11, q_arr_13_10=>q_cache_arr_13_10, q_arr_13_9=>
      q_cache_arr_13_9, q_arr_13_8=>q_cache_arr_13_8, q_arr_13_7=>
      q_cache_arr_13_7, q_arr_13_6=>q_cache_arr_13_6, q_arr_13_5=>
      q_cache_arr_13_5, q_arr_13_4=>q_cache_arr_13_4, q_arr_13_3=>
      q_cache_arr_13_3, q_arr_13_2=>q_cache_arr_13_2, q_arr_13_1=>
      q_cache_arr_13_1, q_arr_13_0=>q_cache_arr_13_0, q_arr_14_31=>
      q_cache_arr_14_31, q_arr_14_30=>q_cache_arr_14_30, q_arr_14_29=>
      q_cache_arr_14_29, q_arr_14_28=>q_cache_arr_14_28, q_arr_14_27=>
      q_cache_arr_14_27, q_arr_14_26=>q_cache_arr_14_26, q_arr_14_25=>
      q_cache_arr_14_25, q_arr_14_24=>q_cache_arr_14_24, q_arr_14_23=>
      q_cache_arr_14_23, q_arr_14_22=>q_cache_arr_14_22, q_arr_14_21=>
      q_cache_arr_14_21, q_arr_14_20=>q_cache_arr_14_20, q_arr_14_19=>
      q_cache_arr_14_19, q_arr_14_18=>q_cache_arr_14_18, q_arr_14_17=>
      q_cache_arr_14_17, q_arr_14_16=>q_cache_arr_14_16, q_arr_14_15=>
      q_cache_arr_14_15, q_arr_14_14=>q_cache_arr_14_14, q_arr_14_13=>
      q_cache_arr_14_13, q_arr_14_12=>q_cache_arr_14_12, q_arr_14_11=>
      q_cache_arr_14_11, q_arr_14_10=>q_cache_arr_14_10, q_arr_14_9=>
      q_cache_arr_14_9, q_arr_14_8=>q_cache_arr_14_8, q_arr_14_7=>
      q_cache_arr_14_7, q_arr_14_6=>q_cache_arr_14_6, q_arr_14_5=>
      q_cache_arr_14_5, q_arr_14_4=>q_cache_arr_14_4, q_arr_14_3=>
      q_cache_arr_14_3, q_arr_14_2=>q_cache_arr_14_2, q_arr_14_1=>
      q_cache_arr_14_1, q_arr_14_0=>q_cache_arr_14_0, q_arr_15_31=>
      q_cache_arr_15_31, q_arr_15_30=>q_cache_arr_15_30, q_arr_15_29=>
      q_cache_arr_15_29, q_arr_15_28=>q_cache_arr_15_28, q_arr_15_27=>
      q_cache_arr_15_27, q_arr_15_26=>q_cache_arr_15_26, q_arr_15_25=>
      q_cache_arr_15_25, q_arr_15_24=>q_cache_arr_15_24, q_arr_15_23=>
      q_cache_arr_15_23, q_arr_15_22=>q_cache_arr_15_22, q_arr_15_21=>
      q_cache_arr_15_21, q_arr_15_20=>q_cache_arr_15_20, q_arr_15_19=>
      q_cache_arr_15_19, q_arr_15_18=>q_cache_arr_15_18, q_arr_15_17=>
      q_cache_arr_15_17, q_arr_15_16=>q_cache_arr_15_16, q_arr_15_15=>
      q_cache_arr_15_15, q_arr_15_14=>q_cache_arr_15_14, q_arr_15_13=>
      q_cache_arr_15_13, q_arr_15_12=>q_cache_arr_15_12, q_arr_15_11=>
      q_cache_arr_15_11, q_arr_15_10=>q_cache_arr_15_10, q_arr_15_9=>
      q_cache_arr_15_9, q_arr_15_8=>q_cache_arr_15_8, q_arr_15_7=>
      q_cache_arr_15_7, q_arr_15_6=>q_cache_arr_15_6, q_arr_15_5=>
      q_cache_arr_15_5, q_arr_15_4=>q_cache_arr_15_4, q_arr_15_3=>
      q_cache_arr_15_3, q_arr_15_2=>q_cache_arr_15_2, q_arr_15_1=>
      q_cache_arr_15_1, q_arr_15_0=>q_cache_arr_15_0, q_arr_16_31=>
      q_cache_arr_16_31, q_arr_16_30=>q_cache_arr_16_30, q_arr_16_29=>
      q_cache_arr_16_29, q_arr_16_28=>q_cache_arr_16_28, q_arr_16_27=>
      q_cache_arr_16_27, q_arr_16_26=>q_cache_arr_16_26, q_arr_16_25=>
      q_cache_arr_16_25, q_arr_16_24=>q_cache_arr_16_24, q_arr_16_23=>
      q_cache_arr_16_23, q_arr_16_22=>q_cache_arr_16_22, q_arr_16_21=>
      q_cache_arr_16_21, q_arr_16_20=>q_cache_arr_16_20, q_arr_16_19=>
      q_cache_arr_16_19, q_arr_16_18=>q_cache_arr_16_18, q_arr_16_17=>
      q_cache_arr_16_17, q_arr_16_16=>q_cache_arr_16_16, q_arr_16_15=>
      q_cache_arr_16_15, q_arr_16_14=>q_cache_arr_16_14, q_arr_16_13=>
      q_cache_arr_16_13, q_arr_16_12=>q_cache_arr_16_12, q_arr_16_11=>
      q_cache_arr_16_11, q_arr_16_10=>q_cache_arr_16_10, q_arr_16_9=>
      q_cache_arr_16_9, q_arr_16_8=>q_cache_arr_16_8, q_arr_16_7=>
      q_cache_arr_16_7, q_arr_16_6=>q_cache_arr_16_6, q_arr_16_5=>
      q_cache_arr_16_5, q_arr_16_4=>q_cache_arr_16_4, q_arr_16_3=>
      q_cache_arr_16_3, q_arr_16_2=>q_cache_arr_16_2, q_arr_16_1=>
      q_cache_arr_16_1, q_arr_16_0=>q_cache_arr_16_0, q_arr_17_31=>
      q_cache_arr_17_31, q_arr_17_30=>q_cache_arr_17_30, q_arr_17_29=>
      q_cache_arr_17_29, q_arr_17_28=>q_cache_arr_17_28, q_arr_17_27=>
      q_cache_arr_17_27, q_arr_17_26=>q_cache_arr_17_26, q_arr_17_25=>
      q_cache_arr_17_25, q_arr_17_24=>q_cache_arr_17_24, q_arr_17_23=>
      q_cache_arr_17_23, q_arr_17_22=>q_cache_arr_17_22, q_arr_17_21=>
      q_cache_arr_17_21, q_arr_17_20=>q_cache_arr_17_20, q_arr_17_19=>
      q_cache_arr_17_19, q_arr_17_18=>q_cache_arr_17_18, q_arr_17_17=>
      q_cache_arr_17_17, q_arr_17_16=>q_cache_arr_17_16, q_arr_17_15=>
      q_cache_arr_17_15, q_arr_17_14=>q_cache_arr_17_14, q_arr_17_13=>
      q_cache_arr_17_13, q_arr_17_12=>q_cache_arr_17_12, q_arr_17_11=>
      q_cache_arr_17_11, q_arr_17_10=>q_cache_arr_17_10, q_arr_17_9=>
      q_cache_arr_17_9, q_arr_17_8=>q_cache_arr_17_8, q_arr_17_7=>
      q_cache_arr_17_7, q_arr_17_6=>q_cache_arr_17_6, q_arr_17_5=>
      q_cache_arr_17_5, q_arr_17_4=>q_cache_arr_17_4, q_arr_17_3=>
      q_cache_arr_17_3, q_arr_17_2=>q_cache_arr_17_2, q_arr_17_1=>
      q_cache_arr_17_1, q_arr_17_0=>q_cache_arr_17_0, q_arr_18_31=>
      q_cache_arr_18_31, q_arr_18_30=>q_cache_arr_18_30, q_arr_18_29=>
      q_cache_arr_18_29, q_arr_18_28=>q_cache_arr_18_28, q_arr_18_27=>
      q_cache_arr_18_27, q_arr_18_26=>q_cache_arr_18_26, q_arr_18_25=>
      q_cache_arr_18_25, q_arr_18_24=>q_cache_arr_18_24, q_arr_18_23=>
      q_cache_arr_18_23, q_arr_18_22=>q_cache_arr_18_22, q_arr_18_21=>
      q_cache_arr_18_21, q_arr_18_20=>q_cache_arr_18_20, q_arr_18_19=>
      q_cache_arr_18_19, q_arr_18_18=>q_cache_arr_18_18, q_arr_18_17=>
      q_cache_arr_18_17, q_arr_18_16=>q_cache_arr_18_16, q_arr_18_15=>
      q_cache_arr_18_15, q_arr_18_14=>q_cache_arr_18_14, q_arr_18_13=>
      q_cache_arr_18_13, q_arr_18_12=>q_cache_arr_18_12, q_arr_18_11=>
      q_cache_arr_18_11, q_arr_18_10=>q_cache_arr_18_10, q_arr_18_9=>
      q_cache_arr_18_9, q_arr_18_8=>q_cache_arr_18_8, q_arr_18_7=>
      q_cache_arr_18_7, q_arr_18_6=>q_cache_arr_18_6, q_arr_18_5=>
      q_cache_arr_18_5, q_arr_18_4=>q_cache_arr_18_4, q_arr_18_3=>
      q_cache_arr_18_3, q_arr_18_2=>q_cache_arr_18_2, q_arr_18_1=>
      q_cache_arr_18_1, q_arr_18_0=>q_cache_arr_18_0, q_arr_19_31=>
      q_cache_arr_19_31, q_arr_19_30=>q_cache_arr_19_30, q_arr_19_29=>
      q_cache_arr_19_29, q_arr_19_28=>q_cache_arr_19_28, q_arr_19_27=>
      q_cache_arr_19_27, q_arr_19_26=>q_cache_arr_19_26, q_arr_19_25=>
      q_cache_arr_19_25, q_arr_19_24=>q_cache_arr_19_24, q_arr_19_23=>
      q_cache_arr_19_23, q_arr_19_22=>q_cache_arr_19_22, q_arr_19_21=>
      q_cache_arr_19_21, q_arr_19_20=>q_cache_arr_19_20, q_arr_19_19=>
      q_cache_arr_19_19, q_arr_19_18=>q_cache_arr_19_18, q_arr_19_17=>
      q_cache_arr_19_17, q_arr_19_16=>q_cache_arr_19_16, q_arr_19_15=>
      q_cache_arr_19_15, q_arr_19_14=>q_cache_arr_19_14, q_arr_19_13=>
      q_cache_arr_19_13, q_arr_19_12=>q_cache_arr_19_12, q_arr_19_11=>
      q_cache_arr_19_11, q_arr_19_10=>q_cache_arr_19_10, q_arr_19_9=>
      q_cache_arr_19_9, q_arr_19_8=>q_cache_arr_19_8, q_arr_19_7=>
      q_cache_arr_19_7, q_arr_19_6=>q_cache_arr_19_6, q_arr_19_5=>
      q_cache_arr_19_5, q_arr_19_4=>q_cache_arr_19_4, q_arr_19_3=>
      q_cache_arr_19_3, q_arr_19_2=>q_cache_arr_19_2, q_arr_19_1=>
      q_cache_arr_19_1, q_arr_19_0=>q_cache_arr_19_0, q_arr_20_31=>
      q_cache_arr_20_31, q_arr_20_30=>q_cache_arr_20_30, q_arr_20_29=>
      q_cache_arr_20_29, q_arr_20_28=>q_cache_arr_20_28, q_arr_20_27=>
      q_cache_arr_20_27, q_arr_20_26=>q_cache_arr_20_26, q_arr_20_25=>
      q_cache_arr_20_25, q_arr_20_24=>q_cache_arr_20_24, q_arr_20_23=>
      q_cache_arr_20_23, q_arr_20_22=>q_cache_arr_20_22, q_arr_20_21=>
      q_cache_arr_20_21, q_arr_20_20=>q_cache_arr_20_20, q_arr_20_19=>
      q_cache_arr_20_19, q_arr_20_18=>q_cache_arr_20_18, q_arr_20_17=>
      q_cache_arr_20_17, q_arr_20_16=>q_cache_arr_20_16, q_arr_20_15=>
      q_cache_arr_20_15, q_arr_20_14=>q_cache_arr_20_14, q_arr_20_13=>
      q_cache_arr_20_13, q_arr_20_12=>q_cache_arr_20_12, q_arr_20_11=>
      q_cache_arr_20_11, q_arr_20_10=>q_cache_arr_20_10, q_arr_20_9=>
      q_cache_arr_20_9, q_arr_20_8=>q_cache_arr_20_8, q_arr_20_7=>
      q_cache_arr_20_7, q_arr_20_6=>q_cache_arr_20_6, q_arr_20_5=>
      q_cache_arr_20_5, q_arr_20_4=>q_cache_arr_20_4, q_arr_20_3=>
      q_cache_arr_20_3, q_arr_20_2=>q_cache_arr_20_2, q_arr_20_1=>
      q_cache_arr_20_1, q_arr_20_0=>q_cache_arr_20_0, q_arr_21_31=>
      q_cache_arr_21_31, q_arr_21_30=>q_cache_arr_21_30, q_arr_21_29=>
      q_cache_arr_21_29, q_arr_21_28=>q_cache_arr_21_28, q_arr_21_27=>
      q_cache_arr_21_27, q_arr_21_26=>q_cache_arr_21_26, q_arr_21_25=>
      q_cache_arr_21_25, q_arr_21_24=>q_cache_arr_21_24, q_arr_21_23=>
      q_cache_arr_21_23, q_arr_21_22=>q_cache_arr_21_22, q_arr_21_21=>
      q_cache_arr_21_21, q_arr_21_20=>q_cache_arr_21_20, q_arr_21_19=>
      q_cache_arr_21_19, q_arr_21_18=>q_cache_arr_21_18, q_arr_21_17=>
      q_cache_arr_21_17, q_arr_21_16=>q_cache_arr_21_16, q_arr_21_15=>
      q_cache_arr_21_15, q_arr_21_14=>q_cache_arr_21_14, q_arr_21_13=>
      q_cache_arr_21_13, q_arr_21_12=>q_cache_arr_21_12, q_arr_21_11=>
      q_cache_arr_21_11, q_arr_21_10=>q_cache_arr_21_10, q_arr_21_9=>
      q_cache_arr_21_9, q_arr_21_8=>q_cache_arr_21_8, q_arr_21_7=>
      q_cache_arr_21_7, q_arr_21_6=>q_cache_arr_21_6, q_arr_21_5=>
      q_cache_arr_21_5, q_arr_21_4=>q_cache_arr_21_4, q_arr_21_3=>
      q_cache_arr_21_3, q_arr_21_2=>q_cache_arr_21_2, q_arr_21_1=>
      q_cache_arr_21_1, q_arr_21_0=>q_cache_arr_21_0, q_arr_22_31=>
      q_cache_arr_22_31, q_arr_22_30=>q_cache_arr_22_30, q_arr_22_29=>
      q_cache_arr_22_29, q_arr_22_28=>q_cache_arr_22_28, q_arr_22_27=>
      q_cache_arr_22_27, q_arr_22_26=>q_cache_arr_22_26, q_arr_22_25=>
      q_cache_arr_22_25, q_arr_22_24=>q_cache_arr_22_24, q_arr_22_23=>
      q_cache_arr_22_23, q_arr_22_22=>q_cache_arr_22_22, q_arr_22_21=>
      q_cache_arr_22_21, q_arr_22_20=>q_cache_arr_22_20, q_arr_22_19=>
      q_cache_arr_22_19, q_arr_22_18=>q_cache_arr_22_18, q_arr_22_17=>
      q_cache_arr_22_17, q_arr_22_16=>q_cache_arr_22_16, q_arr_22_15=>
      q_cache_arr_22_15, q_arr_22_14=>q_cache_arr_22_14, q_arr_22_13=>
      q_cache_arr_22_13, q_arr_22_12=>q_cache_arr_22_12, q_arr_22_11=>
      q_cache_arr_22_11, q_arr_22_10=>q_cache_arr_22_10, q_arr_22_9=>
      q_cache_arr_22_9, q_arr_22_8=>q_cache_arr_22_8, q_arr_22_7=>
      q_cache_arr_22_7, q_arr_22_6=>q_cache_arr_22_6, q_arr_22_5=>
      q_cache_arr_22_5, q_arr_22_4=>q_cache_arr_22_4, q_arr_22_3=>
      q_cache_arr_22_3, q_arr_22_2=>q_cache_arr_22_2, q_arr_22_1=>
      q_cache_arr_22_1, q_arr_22_0=>q_cache_arr_22_0, q_arr_23_31=>
      q_cache_arr_23_31, q_arr_23_30=>q_cache_arr_23_30, q_arr_23_29=>
      q_cache_arr_23_29, q_arr_23_28=>q_cache_arr_23_28, q_arr_23_27=>
      q_cache_arr_23_27, q_arr_23_26=>q_cache_arr_23_26, q_arr_23_25=>
      q_cache_arr_23_25, q_arr_23_24=>q_cache_arr_23_24, q_arr_23_23=>
      q_cache_arr_23_23, q_arr_23_22=>q_cache_arr_23_22, q_arr_23_21=>
      q_cache_arr_23_21, q_arr_23_20=>q_cache_arr_23_20, q_arr_23_19=>
      q_cache_arr_23_19, q_arr_23_18=>q_cache_arr_23_18, q_arr_23_17=>
      q_cache_arr_23_17, q_arr_23_16=>q_cache_arr_23_16, q_arr_23_15=>
      q_cache_arr_23_15, q_arr_23_14=>q_cache_arr_23_14, q_arr_23_13=>
      q_cache_arr_23_13, q_arr_23_12=>q_cache_arr_23_12, q_arr_23_11=>
      q_cache_arr_23_11, q_arr_23_10=>q_cache_arr_23_10, q_arr_23_9=>
      q_cache_arr_23_9, q_arr_23_8=>q_cache_arr_23_8, q_arr_23_7=>
      q_cache_arr_23_7, q_arr_23_6=>q_cache_arr_23_6, q_arr_23_5=>
      q_cache_arr_23_5, q_arr_23_4=>q_cache_arr_23_4, q_arr_23_3=>
      q_cache_arr_23_3, q_arr_23_2=>q_cache_arr_23_2, q_arr_23_1=>
      q_cache_arr_23_1, q_arr_23_0=>q_cache_arr_23_0, q_arr_24_31=>
      q_cache_arr_24_31, q_arr_24_30=>q_cache_arr_24_30, q_arr_24_29=>
      q_cache_arr_24_29, q_arr_24_28=>q_cache_arr_24_28, q_arr_24_27=>
      q_cache_arr_24_27, q_arr_24_26=>q_cache_arr_24_26, q_arr_24_25=>
      q_cache_arr_24_25, q_arr_24_24=>q_cache_arr_24_24, q_arr_24_23=>
      q_cache_arr_24_23, q_arr_24_22=>q_cache_arr_24_22, q_arr_24_21=>
      q_cache_arr_24_21, q_arr_24_20=>q_cache_arr_24_20, q_arr_24_19=>
      q_cache_arr_24_19, q_arr_24_18=>q_cache_arr_24_18, q_arr_24_17=>
      q_cache_arr_24_17, q_arr_24_16=>q_cache_arr_24_16, q_arr_24_15=>
      q_cache_arr_24_15, q_arr_24_14=>q_cache_arr_24_14, q_arr_24_13=>
      q_cache_arr_24_13, q_arr_24_12=>q_cache_arr_24_12, q_arr_24_11=>
      q_cache_arr_24_11, q_arr_24_10=>q_cache_arr_24_10, q_arr_24_9=>
      q_cache_arr_24_9, q_arr_24_8=>q_cache_arr_24_8, q_arr_24_7=>
      q_cache_arr_24_7, q_arr_24_6=>q_cache_arr_24_6, q_arr_24_5=>
      q_cache_arr_24_5, q_arr_24_4=>q_cache_arr_24_4, q_arr_24_3=>
      q_cache_arr_24_3, q_arr_24_2=>q_cache_arr_24_2, q_arr_24_1=>
      q_cache_arr_24_1, q_arr_24_0=>q_cache_arr_24_0, output1_init(15)=>
      output1_init_q_15, output1_init(14)=>output1_init_q_14, 
      output1_init(13)=>output1_init_q_13, output1_init(12)=>
      output1_init_q_12, output1_init(11)=>output1_init_q_11, 
      output1_init(10)=>output1_init_q_10, output1_init(9)=>output1_init_q_9, 
      output1_init(8)=>output1_init_q_8, output1_init(7)=>output1_init_q_7, 
      output1_init(6)=>output1_init_q_6, output1_init(5)=>output1_init_q_5, 
      output1_init(4)=>output1_init_q_4, output1_init(3)=>output1_init_q_3, 
      output1_init(2)=>output1_init_q_2, output1_init(1)=>output1_init_q_1, 
      output1_init(0)=>output1_init_q_0, output2_init(15)=>output2_init_q_15, 
      output2_init(14)=>output2_init_q_14, output2_init(13)=>
      output2_init_q_13, output2_init(12)=>output2_init_q_12, 
      output2_init(11)=>output2_init_q_11, output2_init(10)=>
      output2_init_q_10, output2_init(9)=>output2_init_q_9, output2_init(8)
      =>output2_init_q_8, output2_init(7)=>output2_init_q_7, output2_init(6)
      =>output2_init_q_6, output2_init(5)=>output2_init_q_5, output2_init(4)
      =>output2_init_q_4, output2_init(3)=>output2_init_q_3, output2_init(2)
      =>output2_init_q_2, output2_init(1)=>output2_init_q_1, output2_init(0)
      =>output2_init_q_0, filter_size=>nx1119, operation=>operation_q, 
      compute_relu=>compute_relu_q, clk=>clk, en=>comp_pipe_en, reset=>
      comp_pipe_rst, buffer_ready=>buffer_ready_tmp, semi_ready=>semi_ready, 
      ready=>ready_tmp);
   gen_img_window_gen_queues_0_queuei : Queue_5_unfolded0 port map ( d(15)=>
      img_data_col_0(15), d(14)=>img_data_col_0(14), d(13)=>
      img_data_col_0(13), d(12)=>img_data_col_0(12), d(11)=>
      img_data_col_0(11), d(10)=>img_data_col_0(10), d(9)=>img_data_col_0(9), 
      d(8)=>img_data_col_0(8), d(7)=>img_data_col_0(7), d(6)=>
      img_data_col_0(6), d(5)=>img_data_col_0(5), d(4)=>img_data_col_0(4), 
      d(3)=>img_data_col_0(3), d(2)=>img_data_col_0(2), d(1)=>
      img_data_col_0(1), d(0)=>img_data_col_0(0), q_0_15=>img_data_0_15, 
      q_0_14=>img_data_0_14, q_0_13=>img_data_0_13, q_0_12=>img_data_0_12, 
      q_0_11=>img_data_0_11, q_0_10=>img_data_0_10, q_0_9=>img_data_0_9, 
      q_0_8=>img_data_0_8, q_0_7=>img_data_0_7, q_0_6=>img_data_0_6, q_0_5=>
      img_data_0_5, q_0_4=>img_data_0_4, q_0_3=>img_data_0_3, q_0_2=>
      img_data_0_2, q_0_1=>img_data_0_1, q_0_0=>img_data_0_0, q_1_15=>
      img_data_1_15, q_1_14=>img_data_1_14, q_1_13=>img_data_1_13, q_1_12=>
      img_data_1_12, q_1_11=>img_data_1_11, q_1_10=>img_data_1_10, q_1_9=>
      img_data_1_9, q_1_8=>img_data_1_8, q_1_7=>img_data_1_7, q_1_6=>
      img_data_1_6, q_1_5=>img_data_1_5, q_1_4=>img_data_1_4, q_1_3=>
      img_data_1_3, q_1_2=>img_data_1_2, q_1_1=>img_data_1_1, q_1_0=>
      img_data_1_0, q_2_15=>img_data_2_15, q_2_14=>img_data_2_14, q_2_13=>
      img_data_2_13, q_2_12=>img_data_2_12, q_2_11=>img_data_2_11, q_2_10=>
      img_data_2_10, q_2_9=>img_data_2_9, q_2_8=>img_data_2_8, q_2_7=>
      img_data_2_7, q_2_6=>img_data_2_6, q_2_5=>img_data_2_5, q_2_4=>
      img_data_2_4, q_2_3=>img_data_2_3, q_2_2=>img_data_2_2, q_2_1=>
      img_data_2_1, q_2_0=>img_data_2_0, q_3_15=>img_data_3_15, q_3_14=>
      img_data_3_14, q_3_13=>img_data_3_13, q_3_12=>img_data_3_12, q_3_11=>
      img_data_3_11, q_3_10=>img_data_3_10, q_3_9=>img_data_3_9, q_3_8=>
      img_data_3_8, q_3_7=>img_data_3_7, q_3_6=>img_data_3_6, q_3_5=>
      img_data_3_5, q_3_4=>img_data_3_4, q_3_3=>img_data_3_3, q_3_2=>
      img_data_3_2, q_3_1=>img_data_3_1, q_3_0=>img_data_3_0, q_4_15=>
      img_data_4_15, q_4_14=>img_data_4_14, q_4_13=>img_data_4_13, q_4_12=>
      img_data_4_12, q_4_11=>img_data_4_11, q_4_10=>img_data_4_10, q_4_9=>
      img_data_4_9, q_4_8=>img_data_4_8, q_4_7=>img_data_4_7, q_4_6=>
      img_data_4_6, q_4_5=>img_data_4_5, q_4_4=>img_data_4_4, q_4_3=>
      img_data_4_3, q_4_2=>img_data_4_2, q_4_1=>img_data_4_1, q_4_0=>
      img_data_4_0, clk=>nx1181, load=>nx1177, reset=>buffer_ready_EXMPLR);
   gen_img_window_gen_queues_1_queuei : Queue_5_unfolded0 port map ( d(15)=>
      img_data_col_1(15), d(14)=>img_data_col_1(14), d(13)=>
      img_data_col_1(13), d(12)=>img_data_col_1(12), d(11)=>
      img_data_col_1(11), d(10)=>img_data_col_1(10), d(9)=>img_data_col_1(9), 
      d(8)=>img_data_col_1(8), d(7)=>img_data_col_1(7), d(6)=>
      img_data_col_1(6), d(5)=>img_data_col_1(5), d(4)=>img_data_col_1(4), 
      d(3)=>img_data_col_1(3), d(2)=>img_data_col_1(2), d(1)=>
      img_data_col_1(1), d(0)=>img_data_col_1(0), q_0_15=>img_data_5_15, 
      q_0_14=>img_data_5_14, q_0_13=>img_data_5_13, q_0_12=>img_data_5_12, 
      q_0_11=>img_data_5_11, q_0_10=>img_data_5_10, q_0_9=>img_data_5_9, 
      q_0_8=>img_data_5_8, q_0_7=>img_data_5_7, q_0_6=>img_data_5_6, q_0_5=>
      img_data_5_5, q_0_4=>img_data_5_4, q_0_3=>img_data_5_3, q_0_2=>
      img_data_5_2, q_0_1=>img_data_5_1, q_0_0=>img_data_5_0, q_1_15=>
      img_data_6_15, q_1_14=>img_data_6_14, q_1_13=>img_data_6_13, q_1_12=>
      img_data_6_12, q_1_11=>img_data_6_11, q_1_10=>img_data_6_10, q_1_9=>
      img_data_6_9, q_1_8=>img_data_6_8, q_1_7=>img_data_6_7, q_1_6=>
      img_data_6_6, q_1_5=>img_data_6_5, q_1_4=>img_data_6_4, q_1_3=>
      img_data_6_3, q_1_2=>img_data_6_2, q_1_1=>img_data_6_1, q_1_0=>
      img_data_6_0, q_2_15=>img_data_7_15, q_2_14=>img_data_7_14, q_2_13=>
      img_data_7_13, q_2_12=>img_data_7_12, q_2_11=>img_data_7_11, q_2_10=>
      img_data_7_10, q_2_9=>img_data_7_9, q_2_8=>img_data_7_8, q_2_7=>
      img_data_7_7, q_2_6=>img_data_7_6, q_2_5=>img_data_7_5, q_2_4=>
      img_data_7_4, q_2_3=>img_data_7_3, q_2_2=>img_data_7_2, q_2_1=>
      img_data_7_1, q_2_0=>img_data_7_0, q_3_15=>img_data_8_15, q_3_14=>
      img_data_8_14, q_3_13=>img_data_8_13, q_3_12=>img_data_8_12, q_3_11=>
      img_data_8_11, q_3_10=>img_data_8_10, q_3_9=>img_data_8_9, q_3_8=>
      img_data_8_8, q_3_7=>img_data_8_7, q_3_6=>img_data_8_6, q_3_5=>
      img_data_8_5, q_3_4=>img_data_8_4, q_3_3=>img_data_8_3, q_3_2=>
      img_data_8_2, q_3_1=>img_data_8_1, q_3_0=>img_data_8_0, q_4_15=>
      img_data_9_15, q_4_14=>img_data_9_14, q_4_13=>img_data_9_13, q_4_12=>
      img_data_9_12, q_4_11=>img_data_9_11, q_4_10=>img_data_9_10, q_4_9=>
      img_data_9_9, q_4_8=>img_data_9_8, q_4_7=>img_data_9_7, q_4_6=>
      img_data_9_6, q_4_5=>img_data_9_5, q_4_4=>img_data_9_4, q_4_3=>
      img_data_9_3, q_4_2=>img_data_9_2, q_4_1=>img_data_9_1, q_4_0=>
      img_data_9_0, clk=>nx1181, load=>nx1177, reset=>buffer_ready_EXMPLR);
   gen_img_window_gen_queues_2_queuei : Queue_5_unfolded0 port map ( d(15)=>
      img_data_col_2(15), d(14)=>img_data_col_2(14), d(13)=>
      img_data_col_2(13), d(12)=>img_data_col_2(12), d(11)=>
      img_data_col_2(11), d(10)=>img_data_col_2(10), d(9)=>img_data_col_2(9), 
      d(8)=>img_data_col_2(8), d(7)=>img_data_col_2(7), d(6)=>
      img_data_col_2(6), d(5)=>img_data_col_2(5), d(4)=>img_data_col_2(4), 
      d(3)=>img_data_col_2(3), d(2)=>img_data_col_2(2), d(1)=>
      img_data_col_2(1), d(0)=>img_data_col_2(0), q_0_15=>img_data_10_15, 
      q_0_14=>img_data_10_14, q_0_13=>img_data_10_13, q_0_12=>img_data_10_12, 
      q_0_11=>img_data_10_11, q_0_10=>img_data_10_10, q_0_9=>img_data_10_9, 
      q_0_8=>img_data_10_8, q_0_7=>img_data_10_7, q_0_6=>img_data_10_6, 
      q_0_5=>img_data_10_5, q_0_4=>img_data_10_4, q_0_3=>img_data_10_3, 
      q_0_2=>img_data_10_2, q_0_1=>img_data_10_1, q_0_0=>img_data_10_0, 
      q_1_15=>img_data_11_15, q_1_14=>img_data_11_14, q_1_13=>img_data_11_13, 
      q_1_12=>img_data_11_12, q_1_11=>img_data_11_11, q_1_10=>img_data_11_10, 
      q_1_9=>img_data_11_9, q_1_8=>img_data_11_8, q_1_7=>img_data_11_7, 
      q_1_6=>img_data_11_6, q_1_5=>img_data_11_5, q_1_4=>img_data_11_4, 
      q_1_3=>img_data_11_3, q_1_2=>img_data_11_2, q_1_1=>img_data_11_1, 
      q_1_0=>img_data_11_0, q_2_15=>img_data_12_15, q_2_14=>img_data_12_14, 
      q_2_13=>img_data_12_13, q_2_12=>img_data_12_12, q_2_11=>img_data_12_11, 
      q_2_10=>img_data_12_10, q_2_9=>img_data_12_9, q_2_8=>img_data_12_8, 
      q_2_7=>img_data_12_7, q_2_6=>img_data_12_6, q_2_5=>img_data_12_5, 
      q_2_4=>img_data_12_4, q_2_3=>img_data_12_3, q_2_2=>img_data_12_2, 
      q_2_1=>img_data_12_1, q_2_0=>img_data_12_0, q_3_15=>img_data_13_15, 
      q_3_14=>img_data_13_14, q_3_13=>img_data_13_13, q_3_12=>img_data_13_12, 
      q_3_11=>img_data_13_11, q_3_10=>img_data_13_10, q_3_9=>img_data_13_9, 
      q_3_8=>img_data_13_8, q_3_7=>img_data_13_7, q_3_6=>img_data_13_6, 
      q_3_5=>img_data_13_5, q_3_4=>img_data_13_4, q_3_3=>img_data_13_3, 
      q_3_2=>img_data_13_2, q_3_1=>img_data_13_1, q_3_0=>img_data_13_0, 
      q_4_15=>img_data_14_15, q_4_14=>img_data_14_14, q_4_13=>img_data_14_13, 
      q_4_12=>img_data_14_12, q_4_11=>img_data_14_11, q_4_10=>img_data_14_10, 
      q_4_9=>img_data_14_9, q_4_8=>img_data_14_8, q_4_7=>img_data_14_7, 
      q_4_6=>img_data_14_6, q_4_5=>img_data_14_5, q_4_4=>img_data_14_4, 
      q_4_3=>img_data_14_3, q_4_2=>img_data_14_2, q_4_1=>img_data_14_1, 
      q_4_0=>img_data_14_0, clk=>nx1181, load=>nx1177, reset=>
      buffer_ready_EXMPLR);
   gen_img_window_gen_queues_3_queuei : Queue_5_unfolded0 port map ( d(15)=>
      img_data_col_3(15), d(14)=>img_data_col_3(14), d(13)=>
      img_data_col_3(13), d(12)=>img_data_col_3(12), d(11)=>
      img_data_col_3(11), d(10)=>img_data_col_3(10), d(9)=>img_data_col_3(9), 
      d(8)=>img_data_col_3(8), d(7)=>img_data_col_3(7), d(6)=>
      img_data_col_3(6), d(5)=>img_data_col_3(5), d(4)=>img_data_col_3(4), 
      d(3)=>img_data_col_3(3), d(2)=>img_data_col_3(2), d(1)=>
      img_data_col_3(1), d(0)=>img_data_col_3(0), q_0_15=>img_data_15_15, 
      q_0_14=>img_data_15_14, q_0_13=>img_data_15_13, q_0_12=>img_data_15_12, 
      q_0_11=>img_data_15_11, q_0_10=>img_data_15_10, q_0_9=>img_data_15_9, 
      q_0_8=>img_data_15_8, q_0_7=>img_data_15_7, q_0_6=>img_data_15_6, 
      q_0_5=>img_data_15_5, q_0_4=>img_data_15_4, q_0_3=>img_data_15_3, 
      q_0_2=>img_data_15_2, q_0_1=>img_data_15_1, q_0_0=>img_data_15_0, 
      q_1_15=>img_data_16_15, q_1_14=>img_data_16_14, q_1_13=>img_data_16_13, 
      q_1_12=>img_data_16_12, q_1_11=>img_data_16_11, q_1_10=>img_data_16_10, 
      q_1_9=>img_data_16_9, q_1_8=>img_data_16_8, q_1_7=>img_data_16_7, 
      q_1_6=>img_data_16_6, q_1_5=>img_data_16_5, q_1_4=>img_data_16_4, 
      q_1_3=>img_data_16_3, q_1_2=>img_data_16_2, q_1_1=>img_data_16_1, 
      q_1_0=>img_data_16_0, q_2_15=>img_data_17_15, q_2_14=>img_data_17_14, 
      q_2_13=>img_data_17_13, q_2_12=>img_data_17_12, q_2_11=>img_data_17_11, 
      q_2_10=>img_data_17_10, q_2_9=>img_data_17_9, q_2_8=>img_data_17_8, 
      q_2_7=>img_data_17_7, q_2_6=>img_data_17_6, q_2_5=>img_data_17_5, 
      q_2_4=>img_data_17_4, q_2_3=>img_data_17_3, q_2_2=>img_data_17_2, 
      q_2_1=>img_data_17_1, q_2_0=>img_data_17_0, q_3_15=>img_data_18_15, 
      q_3_14=>img_data_18_14, q_3_13=>img_data_18_13, q_3_12=>img_data_18_12, 
      q_3_11=>img_data_18_11, q_3_10=>img_data_18_10, q_3_9=>img_data_18_9, 
      q_3_8=>img_data_18_8, q_3_7=>img_data_18_7, q_3_6=>img_data_18_6, 
      q_3_5=>img_data_18_5, q_3_4=>img_data_18_4, q_3_3=>img_data_18_3, 
      q_3_2=>img_data_18_2, q_3_1=>img_data_18_1, q_3_0=>img_data_18_0, 
      q_4_15=>img_data_19_15, q_4_14=>img_data_19_14, q_4_13=>img_data_19_13, 
      q_4_12=>img_data_19_12, q_4_11=>img_data_19_11, q_4_10=>img_data_19_10, 
      q_4_9=>img_data_19_9, q_4_8=>img_data_19_8, q_4_7=>img_data_19_7, 
      q_4_6=>img_data_19_6, q_4_5=>img_data_19_5, q_4_4=>img_data_19_4, 
      q_4_3=>img_data_19_3, q_4_2=>img_data_19_2, q_4_1=>img_data_19_1, 
      q_4_0=>img_data_19_0, clk=>nx1183, load=>nx1179, reset=>
      buffer_ready_EXMPLR);
   gen_img_window_gen_queues_4_queuei : Queue_5_unfolded0 port map ( d(15)=>
      img_data_col_4(15), d(14)=>img_data_col_4(14), d(13)=>
      img_data_col_4(13), d(12)=>img_data_col_4(12), d(11)=>
      img_data_col_4(11), d(10)=>img_data_col_4(10), d(9)=>img_data_col_4(9), 
      d(8)=>img_data_col_4(8), d(7)=>img_data_col_4(7), d(6)=>
      img_data_col_4(6), d(5)=>img_data_col_4(5), d(4)=>img_data_col_4(4), 
      d(3)=>img_data_col_4(3), d(2)=>img_data_col_4(2), d(1)=>
      img_data_col_4(1), d(0)=>img_data_col_4(0), q_0_15=>img_data_20_15, 
      q_0_14=>img_data_20_14, q_0_13=>img_data_20_13, q_0_12=>img_data_20_12, 
      q_0_11=>img_data_20_11, q_0_10=>img_data_20_10, q_0_9=>img_data_20_9, 
      q_0_8=>img_data_20_8, q_0_7=>img_data_20_7, q_0_6=>img_data_20_6, 
      q_0_5=>img_data_20_5, q_0_4=>img_data_20_4, q_0_3=>img_data_20_3, 
      q_0_2=>img_data_20_2, q_0_1=>img_data_20_1, q_0_0=>img_data_20_0, 
      q_1_15=>img_data_21_15, q_1_14=>img_data_21_14, q_1_13=>img_data_21_13, 
      q_1_12=>img_data_21_12, q_1_11=>img_data_21_11, q_1_10=>img_data_21_10, 
      q_1_9=>img_data_21_9, q_1_8=>img_data_21_8, q_1_7=>img_data_21_7, 
      q_1_6=>img_data_21_6, q_1_5=>img_data_21_5, q_1_4=>img_data_21_4, 
      q_1_3=>img_data_21_3, q_1_2=>img_data_21_2, q_1_1=>img_data_21_1, 
      q_1_0=>img_data_21_0, q_2_15=>img_data_22_15, q_2_14=>img_data_22_14, 
      q_2_13=>img_data_22_13, q_2_12=>img_data_22_12, q_2_11=>img_data_22_11, 
      q_2_10=>img_data_22_10, q_2_9=>img_data_22_9, q_2_8=>img_data_22_8, 
      q_2_7=>img_data_22_7, q_2_6=>img_data_22_6, q_2_5=>img_data_22_5, 
      q_2_4=>img_data_22_4, q_2_3=>img_data_22_3, q_2_2=>img_data_22_2, 
      q_2_1=>img_data_22_1, q_2_0=>img_data_22_0, q_3_15=>img_data_23_15, 
      q_3_14=>img_data_23_14, q_3_13=>img_data_23_13, q_3_12=>img_data_23_12, 
      q_3_11=>img_data_23_11, q_3_10=>img_data_23_10, q_3_9=>img_data_23_9, 
      q_3_8=>img_data_23_8, q_3_7=>img_data_23_7, q_3_6=>img_data_23_6, 
      q_3_5=>img_data_23_5, q_3_4=>img_data_23_4, q_3_3=>img_data_23_3, 
      q_3_2=>img_data_23_2, q_3_1=>img_data_23_1, q_3_0=>img_data_23_0, 
      q_4_15=>img_data_24_15, q_4_14=>img_data_24_14, q_4_13=>img_data_24_13, 
      q_4_12=>img_data_24_12, q_4_11=>img_data_24_11, q_4_10=>img_data_24_10, 
      q_4_9=>img_data_24_9, q_4_8=>img_data_24_8, q_4_7=>img_data_24_7, 
      q_4_6=>img_data_24_6, q_4_5=>img_data_24_5, q_4_4=>img_data_24_4, 
      q_4_3=>img_data_24_3, q_4_2=>img_data_24_2, q_4_1=>img_data_24_1, 
      q_4_0=>img_data_24_0, clk=>nx1183, load=>nx1179, reset=>
      buffer_ready_EXMPLR);
   gen_filter_window_queuei : Queue_25 port map ( d(15)=>
      filter_data_word(15), d(14)=>filter_data_word(14), d(13)=>
      filter_data_word(13), d(12)=>filter_data_word(12), d(11)=>
      filter_data_word(11), d(10)=>filter_data_word(10), d(9)=>
      filter_data_word(9), d(8)=>filter_data_word(8), d(7)=>
      filter_data_word(7), d(6)=>filter_data_word(6), d(5)=>
      filter_data_word(5), d(4)=>filter_data_word(4), d(3)=>
      filter_data_word(3), d(2)=>filter_data_word(2), d(1)=>
      filter_data_word(1), d(0)=>filter_data_word(0), q_0_15=>
      filter_data_0_15, q_0_14=>filter_data_0_14, q_0_13=>filter_data_0_13, 
      q_0_12=>filter_data_0_12, q_0_11=>filter_data_0_11, q_0_10=>
      filter_data_0_10, q_0_9=>filter_data_0_9, q_0_8=>filter_data_0_8, 
      q_0_7=>filter_data_0_7, q_0_6=>filter_data_0_6, q_0_5=>filter_data_0_5, 
      q_0_4=>filter_data_0_4, q_0_3=>filter_data_0_3, q_0_2=>filter_data_0_2, 
      q_0_1=>filter_data_0_1, q_0_0=>filter_data_0_0, q_1_15=>
      filter_data_1_15, q_1_14=>filter_data_1_14, q_1_13=>filter_data_1_13, 
      q_1_12=>filter_data_1_12, q_1_11=>filter_data_1_11, q_1_10=>
      filter_data_1_10, q_1_9=>filter_data_1_9, q_1_8=>filter_data_1_8, 
      q_1_7=>filter_data_1_7, q_1_6=>filter_data_1_6, q_1_5=>filter_data_1_5, 
      q_1_4=>filter_data_1_4, q_1_3=>filter_data_1_3, q_1_2=>filter_data_1_2, 
      q_1_1=>filter_data_1_1, q_1_0=>filter_data_1_0, q_2_15=>
      filter_data_2_15, q_2_14=>filter_data_2_14, q_2_13=>filter_data_2_13, 
      q_2_12=>filter_data_2_12, q_2_11=>filter_data_2_11, q_2_10=>
      filter_data_2_10, q_2_9=>filter_data_2_9, q_2_8=>filter_data_2_8, 
      q_2_7=>filter_data_2_7, q_2_6=>filter_data_2_6, q_2_5=>filter_data_2_5, 
      q_2_4=>filter_data_2_4, q_2_3=>filter_data_2_3, q_2_2=>filter_data_2_2, 
      q_2_1=>filter_data_2_1, q_2_0=>filter_data_2_0, q_3_15=>
      filter_data_3_15, q_3_14=>filter_data_3_14, q_3_13=>filter_data_3_13, 
      q_3_12=>filter_data_3_12, q_3_11=>filter_data_3_11, q_3_10=>
      filter_data_3_10, q_3_9=>filter_data_3_9, q_3_8=>filter_data_3_8, 
      q_3_7=>filter_data_3_7, q_3_6=>filter_data_3_6, q_3_5=>filter_data_3_5, 
      q_3_4=>filter_data_3_4, q_3_3=>filter_data_3_3, q_3_2=>filter_data_3_2, 
      q_3_1=>filter_data_3_1, q_3_0=>filter_data_3_0, q_4_15=>
      filter_data_4_15, q_4_14=>filter_data_4_14, q_4_13=>filter_data_4_13, 
      q_4_12=>filter_data_4_12, q_4_11=>filter_data_4_11, q_4_10=>
      filter_data_4_10, q_4_9=>filter_data_4_9, q_4_8=>filter_data_4_8, 
      q_4_7=>filter_data_4_7, q_4_6=>filter_data_4_6, q_4_5=>filter_data_4_5, 
      q_4_4=>filter_data_4_4, q_4_3=>filter_data_4_3, q_4_2=>filter_data_4_2, 
      q_4_1=>filter_data_4_1, q_4_0=>filter_data_4_0, q_5_15=>
      filter_data_5_15, q_5_14=>filter_data_5_14, q_5_13=>filter_data_5_13, 
      q_5_12=>filter_data_5_12, q_5_11=>filter_data_5_11, q_5_10=>
      filter_data_5_10, q_5_9=>filter_data_5_9, q_5_8=>filter_data_5_8, 
      q_5_7=>filter_data_5_7, q_5_6=>filter_data_5_6, q_5_5=>filter_data_5_5, 
      q_5_4=>filter_data_5_4, q_5_3=>filter_data_5_3, q_5_2=>filter_data_5_2, 
      q_5_1=>filter_data_5_1, q_5_0=>filter_data_5_0, q_6_15=>
      filter_data_6_15, q_6_14=>filter_data_6_14, q_6_13=>filter_data_6_13, 
      q_6_12=>filter_data_6_12, q_6_11=>filter_data_6_11, q_6_10=>
      filter_data_6_10, q_6_9=>filter_data_6_9, q_6_8=>filter_data_6_8, 
      q_6_7=>filter_data_6_7, q_6_6=>filter_data_6_6, q_6_5=>filter_data_6_5, 
      q_6_4=>filter_data_6_4, q_6_3=>filter_data_6_3, q_6_2=>filter_data_6_2, 
      q_6_1=>filter_data_6_1, q_6_0=>filter_data_6_0, q_7_15=>
      filter_data_7_15, q_7_14=>filter_data_7_14, q_7_13=>filter_data_7_13, 
      q_7_12=>filter_data_7_12, q_7_11=>filter_data_7_11, q_7_10=>
      filter_data_7_10, q_7_9=>filter_data_7_9, q_7_8=>filter_data_7_8, 
      q_7_7=>filter_data_7_7, q_7_6=>filter_data_7_6, q_7_5=>filter_data_7_5, 
      q_7_4=>filter_data_7_4, q_7_3=>filter_data_7_3, q_7_2=>filter_data_7_2, 
      q_7_1=>filter_data_7_1, q_7_0=>filter_data_7_0, q_8_15=>
      filter_data_8_15, q_8_14=>filter_data_8_14, q_8_13=>filter_data_8_13, 
      q_8_12=>filter_data_8_12, q_8_11=>filter_data_8_11, q_8_10=>
      filter_data_8_10, q_8_9=>filter_data_8_9, q_8_8=>filter_data_8_8, 
      q_8_7=>filter_data_8_7, q_8_6=>filter_data_8_6, q_8_5=>filter_data_8_5, 
      q_8_4=>filter_data_8_4, q_8_3=>filter_data_8_3, q_8_2=>filter_data_8_2, 
      q_8_1=>filter_data_8_1, q_8_0=>filter_data_8_0, q_9_15=>
      filter_data_9_15, q_9_14=>filter_data_9_14, q_9_13=>filter_data_9_13, 
      q_9_12=>filter_data_9_12, q_9_11=>filter_data_9_11, q_9_10=>
      filter_data_9_10, q_9_9=>filter_data_9_9, q_9_8=>filter_data_9_8, 
      q_9_7=>filter_data_9_7, q_9_6=>filter_data_9_6, q_9_5=>filter_data_9_5, 
      q_9_4=>filter_data_9_4, q_9_3=>filter_data_9_3, q_9_2=>filter_data_9_2, 
      q_9_1=>filter_data_9_1, q_9_0=>filter_data_9_0, q_10_15=>
      filter_data_10_15, q_10_14=>filter_data_10_14, q_10_13=>
      filter_data_10_13, q_10_12=>filter_data_10_12, q_10_11=>
      filter_data_10_11, q_10_10=>filter_data_10_10, q_10_9=>
      filter_data_10_9, q_10_8=>filter_data_10_8, q_10_7=>filter_data_10_7, 
      q_10_6=>filter_data_10_6, q_10_5=>filter_data_10_5, q_10_4=>
      filter_data_10_4, q_10_3=>filter_data_10_3, q_10_2=>filter_data_10_2, 
      q_10_1=>filter_data_10_1, q_10_0=>filter_data_10_0, q_11_15=>
      filter_data_11_15, q_11_14=>filter_data_11_14, q_11_13=>
      filter_data_11_13, q_11_12=>filter_data_11_12, q_11_11=>
      filter_data_11_11, q_11_10=>filter_data_11_10, q_11_9=>
      filter_data_11_9, q_11_8=>filter_data_11_8, q_11_7=>filter_data_11_7, 
      q_11_6=>filter_data_11_6, q_11_5=>filter_data_11_5, q_11_4=>
      filter_data_11_4, q_11_3=>filter_data_11_3, q_11_2=>filter_data_11_2, 
      q_11_1=>filter_data_11_1, q_11_0=>filter_data_11_0, q_12_15=>
      filter_data_12_15, q_12_14=>filter_data_12_14, q_12_13=>
      filter_data_12_13, q_12_12=>filter_data_12_12, q_12_11=>
      filter_data_12_11, q_12_10=>filter_data_12_10, q_12_9=>
      filter_data_12_9, q_12_8=>filter_data_12_8, q_12_7=>filter_data_12_7, 
      q_12_6=>filter_data_12_6, q_12_5=>filter_data_12_5, q_12_4=>
      filter_data_12_4, q_12_3=>filter_data_12_3, q_12_2=>filter_data_12_2, 
      q_12_1=>filter_data_12_1, q_12_0=>filter_data_12_0, q_13_15=>
      filter_data_13_15, q_13_14=>filter_data_13_14, q_13_13=>
      filter_data_13_13, q_13_12=>filter_data_13_12, q_13_11=>
      filter_data_13_11, q_13_10=>filter_data_13_10, q_13_9=>
      filter_data_13_9, q_13_8=>filter_data_13_8, q_13_7=>filter_data_13_7, 
      q_13_6=>filter_data_13_6, q_13_5=>filter_data_13_5, q_13_4=>
      filter_data_13_4, q_13_3=>filter_data_13_3, q_13_2=>filter_data_13_2, 
      q_13_1=>filter_data_13_1, q_13_0=>filter_data_13_0, q_14_15=>
      filter_data_14_15, q_14_14=>filter_data_14_14, q_14_13=>
      filter_data_14_13, q_14_12=>filter_data_14_12, q_14_11=>
      filter_data_14_11, q_14_10=>filter_data_14_10, q_14_9=>
      filter_data_14_9, q_14_8=>filter_data_14_8, q_14_7=>filter_data_14_7, 
      q_14_6=>filter_data_14_6, q_14_5=>filter_data_14_5, q_14_4=>
      filter_data_14_4, q_14_3=>filter_data_14_3, q_14_2=>filter_data_14_2, 
      q_14_1=>filter_data_14_1, q_14_0=>filter_data_14_0, q_15_15=>
      filter_data_15_15, q_15_14=>filter_data_15_14, q_15_13=>
      filter_data_15_13, q_15_12=>filter_data_15_12, q_15_11=>
      filter_data_15_11, q_15_10=>filter_data_15_10, q_15_9=>
      filter_data_15_9, q_15_8=>filter_data_15_8, q_15_7=>filter_data_15_7, 
      q_15_6=>filter_data_15_6, q_15_5=>filter_data_15_5, q_15_4=>
      filter_data_15_4, q_15_3=>filter_data_15_3, q_15_2=>filter_data_15_2, 
      q_15_1=>filter_data_15_1, q_15_0=>filter_data_15_0, q_16_15=>
      filter_data_16_15, q_16_14=>filter_data_16_14, q_16_13=>
      filter_data_16_13, q_16_12=>filter_data_16_12, q_16_11=>
      filter_data_16_11, q_16_10=>filter_data_16_10, q_16_9=>
      filter_data_16_9, q_16_8=>filter_data_16_8, q_16_7=>filter_data_16_7, 
      q_16_6=>filter_data_16_6, q_16_5=>filter_data_16_5, q_16_4=>
      filter_data_16_4, q_16_3=>filter_data_16_3, q_16_2=>filter_data_16_2, 
      q_16_1=>filter_data_16_1, q_16_0=>filter_data_16_0, q_17_15=>
      filter_data_17_15, q_17_14=>filter_data_17_14, q_17_13=>
      filter_data_17_13, q_17_12=>filter_data_17_12, q_17_11=>
      filter_data_17_11, q_17_10=>filter_data_17_10, q_17_9=>
      filter_data_17_9, q_17_8=>filter_data_17_8, q_17_7=>filter_data_17_7, 
      q_17_6=>filter_data_17_6, q_17_5=>filter_data_17_5, q_17_4=>
      filter_data_17_4, q_17_3=>filter_data_17_3, q_17_2=>filter_data_17_2, 
      q_17_1=>filter_data_17_1, q_17_0=>filter_data_17_0, q_18_15=>
      filter_data_18_15, q_18_14=>filter_data_18_14, q_18_13=>
      filter_data_18_13, q_18_12=>filter_data_18_12, q_18_11=>
      filter_data_18_11, q_18_10=>filter_data_18_10, q_18_9=>
      filter_data_18_9, q_18_8=>filter_data_18_8, q_18_7=>filter_data_18_7, 
      q_18_6=>filter_data_18_6, q_18_5=>filter_data_18_5, q_18_4=>
      filter_data_18_4, q_18_3=>filter_data_18_3, q_18_2=>filter_data_18_2, 
      q_18_1=>filter_data_18_1, q_18_0=>filter_data_18_0, q_19_15=>
      filter_data_19_15, q_19_14=>filter_data_19_14, q_19_13=>
      filter_data_19_13, q_19_12=>filter_data_19_12, q_19_11=>
      filter_data_19_11, q_19_10=>filter_data_19_10, q_19_9=>
      filter_data_19_9, q_19_8=>filter_data_19_8, q_19_7=>filter_data_19_7, 
      q_19_6=>filter_data_19_6, q_19_5=>filter_data_19_5, q_19_4=>
      filter_data_19_4, q_19_3=>filter_data_19_3, q_19_2=>filter_data_19_2, 
      q_19_1=>filter_data_19_1, q_19_0=>filter_data_19_0, q_20_15=>
      filter_data_20_15, q_20_14=>filter_data_20_14, q_20_13=>
      filter_data_20_13, q_20_12=>filter_data_20_12, q_20_11=>
      filter_data_20_11, q_20_10=>filter_data_20_10, q_20_9=>
      filter_data_20_9, q_20_8=>filter_data_20_8, q_20_7=>filter_data_20_7, 
      q_20_6=>filter_data_20_6, q_20_5=>filter_data_20_5, q_20_4=>
      filter_data_20_4, q_20_3=>filter_data_20_3, q_20_2=>filter_data_20_2, 
      q_20_1=>filter_data_20_1, q_20_0=>filter_data_20_0, q_21_15=>
      filter_data_21_15, q_21_14=>filter_data_21_14, q_21_13=>
      filter_data_21_13, q_21_12=>filter_data_21_12, q_21_11=>
      filter_data_21_11, q_21_10=>filter_data_21_10, q_21_9=>
      filter_data_21_9, q_21_8=>filter_data_21_8, q_21_7=>filter_data_21_7, 
      q_21_6=>filter_data_21_6, q_21_5=>filter_data_21_5, q_21_4=>
      filter_data_21_4, q_21_3=>filter_data_21_3, q_21_2=>filter_data_21_2, 
      q_21_1=>filter_data_21_1, q_21_0=>filter_data_21_0, q_22_15=>
      filter_data_22_15, q_22_14=>filter_data_22_14, q_22_13=>
      filter_data_22_13, q_22_12=>filter_data_22_12, q_22_11=>
      filter_data_22_11, q_22_10=>filter_data_22_10, q_22_9=>
      filter_data_22_9, q_22_8=>filter_data_22_8, q_22_7=>filter_data_22_7, 
      q_22_6=>filter_data_22_6, q_22_5=>filter_data_22_5, q_22_4=>
      filter_data_22_4, q_22_3=>filter_data_22_3, q_22_2=>filter_data_22_2, 
      q_22_1=>filter_data_22_1, q_22_0=>filter_data_22_0, q_23_15=>
      filter_data_23_15, q_23_14=>filter_data_23_14, q_23_13=>
      filter_data_23_13, q_23_12=>filter_data_23_12, q_23_11=>
      filter_data_23_11, q_23_10=>filter_data_23_10, q_23_9=>
      filter_data_23_9, q_23_8=>filter_data_23_8, q_23_7=>filter_data_23_7, 
      q_23_6=>filter_data_23_6, q_23_5=>filter_data_23_5, q_23_4=>
      filter_data_23_4, q_23_3=>filter_data_23_3, q_23_2=>filter_data_23_2, 
      q_23_1=>filter_data_23_1, q_23_0=>filter_data_23_0, q_24_15=>
      filter_data_24_15, q_24_14=>filter_data_24_14, q_24_13=>
      filter_data_24_13, q_24_12=>filter_data_24_12, q_24_11=>
      filter_data_24_11, q_24_10=>filter_data_24_10, q_24_9=>
      filter_data_24_9, q_24_8=>filter_data_24_8, q_24_7=>filter_data_24_7, 
      q_24_6=>filter_data_24_6, q_24_5=>filter_data_24_5, q_24_4=>
      filter_data_24_4, q_24_3=>filter_data_24_3, q_24_2=>filter_data_24_2, 
      q_24_1=>filter_data_24_1, q_24_0=>filter_data_24_0, clk=>nx1181, load
      =>filter_load_tmp, reset=>filter_reset);
   gen_comp_cache_gen_regs_0_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_0_31, d(30)=>d_cache_arr_0_30, d(29)=>d_cache_arr_0_29, 
      d(28)=>d_cache_arr_0_28, d(27)=>d_cache_arr_0_27, d(26)=>
      d_cache_arr_0_26, d(25)=>d_cache_arr_0_25, d(24)=>d_cache_arr_0_24, 
      d(23)=>d_cache_arr_0_23, d(22)=>d_cache_arr_0_22, d(21)=>
      d_cache_arr_0_21, d(20)=>d_cache_arr_0_20, d(19)=>d_cache_arr_0_19, 
      d(18)=>d_cache_arr_0_18, d(17)=>d_cache_arr_0_17, d(16)=>
      d_cache_arr_0_16, d(15)=>d_cache_arr_0_15, d(14)=>d_cache_arr_0_14, 
      d(13)=>d_cache_arr_0_13, d(12)=>d_cache_arr_0_12, d(11)=>
      d_cache_arr_0_11, d(10)=>d_cache_arr_0_10, d(9)=>d_cache_arr_0_9, d(8)
      =>d_cache_arr_0_8, d(7)=>d_cache_arr_0_7, d(6)=>d_cache_arr_0_6, d(5)
      =>d_cache_arr_0_5, d(4)=>d_cache_arr_0_4, d(3)=>d_cache_arr_0_3, d(2)
      =>d_cache_arr_0_2, d(1)=>d_cache_arr_0_1, d(0)=>d_cache_arr_0_0, q(31)
      =>q_cache_arr_0_31, q(30)=>q_cache_arr_0_30, q(29)=>q_cache_arr_0_29, 
      q(28)=>q_cache_arr_0_28, q(27)=>q_cache_arr_0_27, q(26)=>
      q_cache_arr_0_26, q(25)=>q_cache_arr_0_25, q(24)=>q_cache_arr_0_24, 
      q(23)=>q_cache_arr_0_23, q(22)=>q_cache_arr_0_22, q(21)=>
      q_cache_arr_0_21, q(20)=>q_cache_arr_0_20, q(19)=>q_cache_arr_0_19, 
      q(18)=>q_cache_arr_0_18, q(17)=>q_cache_arr_0_17, q(16)=>
      q_cache_arr_0_16, q(15)=>q_cache_arr_0_15, q(14)=>q_cache_arr_0_14, 
      q(13)=>q_cache_arr_0_13, q(12)=>q_cache_arr_0_12, q(11)=>
      q_cache_arr_0_11, q(10)=>q_cache_arr_0_10, q(9)=>q_cache_arr_0_9, q(8)
      =>q_cache_arr_0_8, q(7)=>q_cache_arr_0_7, q(6)=>q_cache_arr_0_6, q(5)
      =>q_cache_arr_0_5, q(4)=>q_cache_arr_0_4, q(3)=>q_cache_arr_0_3, q(2)
      =>q_cache_arr_0_2, q(1)=>q_cache_arr_0_1, q(0)=>q_cache_arr_0_0, 
      rst_data(31)=>buffer_ready_EXMPLR, rst_data(30)=>buffer_ready_EXMPLR, 
      rst_data(29)=>buffer_ready_EXMPLR, rst_data(28)=>buffer_ready_EXMPLR, 
      rst_data(27)=>buffer_ready_EXMPLR, rst_data(26)=>buffer_ready_EXMPLR, 
      rst_data(25)=>buffer_ready_EXMPLR, rst_data(24)=>buffer_ready_EXMPLR, 
      rst_data(23)=>buffer_ready_EXMPLR, rst_data(22)=>buffer_ready_EXMPLR, 
      rst_data(21)=>buffer_ready_EXMPLR, rst_data(20)=>buffer_ready_EXMPLR, 
      rst_data(19)=>buffer_ready_EXMPLR, rst_data(18)=>buffer_ready_EXMPLR, 
      rst_data(17)=>buffer_ready_EXMPLR, rst_data(16)=>buffer_ready_EXMPLR, 
      rst_data(15)=>buffer_ready_EXMPLR, rst_data(14)=>buffer_ready_EXMPLR, 
      rst_data(13)=>buffer_ready_EXMPLR, rst_data(12)=>buffer_ready_EXMPLR, 
      rst_data(11)=>buffer_ready_EXMPLR, rst_data(10)=>buffer_ready_EXMPLR, 
      rst_data(9)=>buffer_ready_EXMPLR, rst_data(8)=>buffer_ready_EXMPLR, 
      rst_data(7)=>buffer_ready_EXMPLR, rst_data(6)=>buffer_ready_EXMPLR, 
      rst_data(5)=>buffer_ready_EXMPLR, rst_data(4)=>buffer_ready_EXMPLR, 
      rst_data(3)=>buffer_ready_EXMPLR, rst_data(2)=>buffer_ready_EXMPLR, 
      rst_data(1)=>buffer_ready_EXMPLR, rst_data(0)=>buffer_ready_EXMPLR, 
      clk=>clk, load=>nx1109, reset=>filter_reset);
   gen_comp_cache_gen_regs_1_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_1_31, d(30)=>d_cache_arr_1_30, d(29)=>d_cache_arr_1_29, 
      d(28)=>d_cache_arr_1_28, d(27)=>d_cache_arr_1_27, d(26)=>
      d_cache_arr_1_26, d(25)=>d_cache_arr_1_25, d(24)=>d_cache_arr_1_24, 
      d(23)=>d_cache_arr_1_23, d(22)=>d_cache_arr_1_22, d(21)=>
      d_cache_arr_1_21, d(20)=>d_cache_arr_1_20, d(19)=>d_cache_arr_1_19, 
      d(18)=>d_cache_arr_1_18, d(17)=>d_cache_arr_1_17, d(16)=>
      d_cache_arr_1_16, d(15)=>d_cache_arr_1_15, d(14)=>d_cache_arr_1_14, 
      d(13)=>d_cache_arr_1_13, d(12)=>d_cache_arr_1_12, d(11)=>
      d_cache_arr_1_11, d(10)=>d_cache_arr_1_10, d(9)=>d_cache_arr_1_9, d(8)
      =>d_cache_arr_1_8, d(7)=>d_cache_arr_1_7, d(6)=>d_cache_arr_1_6, d(5)
      =>d_cache_arr_1_5, d(4)=>d_cache_arr_1_4, d(3)=>d_cache_arr_1_3, d(2)
      =>d_cache_arr_1_2, d(1)=>d_cache_arr_1_1, d(0)=>d_cache_arr_1_0, q(31)
      =>q_cache_arr_1_31, q(30)=>q_cache_arr_1_30, q(29)=>q_cache_arr_1_29, 
      q(28)=>q_cache_arr_1_28, q(27)=>q_cache_arr_1_27, q(26)=>
      q_cache_arr_1_26, q(25)=>q_cache_arr_1_25, q(24)=>q_cache_arr_1_24, 
      q(23)=>q_cache_arr_1_23, q(22)=>q_cache_arr_1_22, q(21)=>
      q_cache_arr_1_21, q(20)=>q_cache_arr_1_20, q(19)=>q_cache_arr_1_19, 
      q(18)=>q_cache_arr_1_18, q(17)=>q_cache_arr_1_17, q(16)=>
      q_cache_arr_1_16, q(15)=>q_cache_arr_1_15, q(14)=>q_cache_arr_1_14, 
      q(13)=>q_cache_arr_1_13, q(12)=>q_cache_arr_1_12, q(11)=>
      q_cache_arr_1_11, q(10)=>q_cache_arr_1_10, q(9)=>q_cache_arr_1_9, q(8)
      =>q_cache_arr_1_8, q(7)=>q_cache_arr_1_7, q(6)=>q_cache_arr_1_6, q(5)
      =>q_cache_arr_1_5, q(4)=>q_cache_arr_1_4, q(3)=>q_cache_arr_1_3, q(2)
      =>q_cache_arr_1_2, q(1)=>q_cache_arr_1_1, q(0)=>q_cache_arr_1_0, 
      rst_data(31)=>buffer_ready_EXMPLR, rst_data(30)=>buffer_ready_EXMPLR, 
      rst_data(29)=>buffer_ready_EXMPLR, rst_data(28)=>buffer_ready_EXMPLR, 
      rst_data(27)=>buffer_ready_EXMPLR, rst_data(26)=>buffer_ready_EXMPLR, 
      rst_data(25)=>buffer_ready_EXMPLR, rst_data(24)=>buffer_ready_EXMPLR, 
      rst_data(23)=>buffer_ready_EXMPLR, rst_data(22)=>buffer_ready_EXMPLR, 
      rst_data(21)=>buffer_ready_EXMPLR, rst_data(20)=>buffer_ready_EXMPLR, 
      rst_data(19)=>buffer_ready_EXMPLR, rst_data(18)=>buffer_ready_EXMPLR, 
      rst_data(17)=>buffer_ready_EXMPLR, rst_data(16)=>buffer_ready_EXMPLR, 
      rst_data(15)=>buffer_ready_EXMPLR, rst_data(14)=>buffer_ready_EXMPLR, 
      rst_data(13)=>buffer_ready_EXMPLR, rst_data(12)=>buffer_ready_EXMPLR, 
      rst_data(11)=>buffer_ready_EXMPLR, rst_data(10)=>buffer_ready_EXMPLR, 
      rst_data(9)=>buffer_ready_EXMPLR, rst_data(8)=>buffer_ready_EXMPLR, 
      rst_data(7)=>buffer_ready_EXMPLR, rst_data(6)=>buffer_ready_EXMPLR, 
      rst_data(5)=>buffer_ready_EXMPLR, rst_data(4)=>buffer_ready_EXMPLR, 
      rst_data(3)=>buffer_ready_EXMPLR, rst_data(2)=>buffer_ready_EXMPLR, 
      rst_data(1)=>buffer_ready_EXMPLR, rst_data(0)=>buffer_ready_EXMPLR, 
      clk=>clk, load=>nx1109, reset=>filter_reset);
   gen_comp_cache_gen_regs_2_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_2_31, d(30)=>d_cache_arr_2_30, d(29)=>d_cache_arr_2_29, 
      d(28)=>d_cache_arr_2_28, d(27)=>d_cache_arr_2_27, d(26)=>
      d_cache_arr_2_26, d(25)=>d_cache_arr_2_25, d(24)=>d_cache_arr_2_24, 
      d(23)=>d_cache_arr_2_23, d(22)=>d_cache_arr_2_22, d(21)=>
      d_cache_arr_2_21, d(20)=>d_cache_arr_2_20, d(19)=>d_cache_arr_2_19, 
      d(18)=>d_cache_arr_2_18, d(17)=>d_cache_arr_2_17, d(16)=>
      d_cache_arr_2_16, d(15)=>d_cache_arr_2_15, d(14)=>d_cache_arr_2_14, 
      d(13)=>d_cache_arr_2_13, d(12)=>d_cache_arr_2_12, d(11)=>
      d_cache_arr_2_11, d(10)=>d_cache_arr_2_10, d(9)=>d_cache_arr_2_9, d(8)
      =>d_cache_arr_2_8, d(7)=>d_cache_arr_2_7, d(6)=>d_cache_arr_2_6, d(5)
      =>d_cache_arr_2_5, d(4)=>d_cache_arr_2_4, d(3)=>d_cache_arr_2_3, d(2)
      =>d_cache_arr_2_2, d(1)=>d_cache_arr_2_1, d(0)=>d_cache_arr_2_0, q(31)
      =>q_cache_arr_2_31, q(30)=>q_cache_arr_2_30, q(29)=>q_cache_arr_2_29, 
      q(28)=>q_cache_arr_2_28, q(27)=>q_cache_arr_2_27, q(26)=>
      q_cache_arr_2_26, q(25)=>q_cache_arr_2_25, q(24)=>q_cache_arr_2_24, 
      q(23)=>q_cache_arr_2_23, q(22)=>q_cache_arr_2_22, q(21)=>
      q_cache_arr_2_21, q(20)=>q_cache_arr_2_20, q(19)=>q_cache_arr_2_19, 
      q(18)=>q_cache_arr_2_18, q(17)=>q_cache_arr_2_17, q(16)=>
      q_cache_arr_2_16, q(15)=>q_cache_arr_2_15, q(14)=>q_cache_arr_2_14, 
      q(13)=>q_cache_arr_2_13, q(12)=>q_cache_arr_2_12, q(11)=>
      q_cache_arr_2_11, q(10)=>q_cache_arr_2_10, q(9)=>q_cache_arr_2_9, q(8)
      =>q_cache_arr_2_8, q(7)=>q_cache_arr_2_7, q(6)=>q_cache_arr_2_6, q(5)
      =>q_cache_arr_2_5, q(4)=>q_cache_arr_2_4, q(3)=>q_cache_arr_2_3, q(2)
      =>q_cache_arr_2_2, q(1)=>q_cache_arr_2_1, q(0)=>q_cache_arr_2_0, 
      rst_data(31)=>buffer_ready_EXMPLR, rst_data(30)=>buffer_ready_EXMPLR, 
      rst_data(29)=>buffer_ready_EXMPLR, rst_data(28)=>buffer_ready_EXMPLR, 
      rst_data(27)=>buffer_ready_EXMPLR, rst_data(26)=>buffer_ready_EXMPLR, 
      rst_data(25)=>buffer_ready_EXMPLR, rst_data(24)=>buffer_ready_EXMPLR, 
      rst_data(23)=>buffer_ready_EXMPLR, rst_data(22)=>buffer_ready_EXMPLR, 
      rst_data(21)=>buffer_ready_EXMPLR, rst_data(20)=>buffer_ready_EXMPLR, 
      rst_data(19)=>buffer_ready_EXMPLR, rst_data(18)=>buffer_ready_EXMPLR, 
      rst_data(17)=>buffer_ready_EXMPLR, rst_data(16)=>buffer_ready_EXMPLR, 
      rst_data(15)=>buffer_ready_EXMPLR, rst_data(14)=>buffer_ready_EXMPLR, 
      rst_data(13)=>buffer_ready_EXMPLR, rst_data(12)=>buffer_ready_EXMPLR, 
      rst_data(11)=>buffer_ready_EXMPLR, rst_data(10)=>buffer_ready_EXMPLR, 
      rst_data(9)=>buffer_ready_EXMPLR, rst_data(8)=>buffer_ready_EXMPLR, 
      rst_data(7)=>buffer_ready_EXMPLR, rst_data(6)=>buffer_ready_EXMPLR, 
      rst_data(5)=>buffer_ready_EXMPLR, rst_data(4)=>buffer_ready_EXMPLR, 
      rst_data(3)=>buffer_ready_EXMPLR, rst_data(2)=>buffer_ready_EXMPLR, 
      rst_data(1)=>buffer_ready_EXMPLR, rst_data(0)=>buffer_ready_EXMPLR, 
      clk=>clk, load=>nx1109, reset=>filter_reset);
   gen_comp_cache_gen_regs_3_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_3_31, d(30)=>d_cache_arr_3_30, d(29)=>d_cache_arr_3_29, 
      d(28)=>d_cache_arr_3_28, d(27)=>d_cache_arr_3_27, d(26)=>
      d_cache_arr_3_26, d(25)=>d_cache_arr_3_25, d(24)=>d_cache_arr_3_24, 
      d(23)=>d_cache_arr_3_23, d(22)=>d_cache_arr_3_22, d(21)=>
      d_cache_arr_3_21, d(20)=>d_cache_arr_3_20, d(19)=>d_cache_arr_3_19, 
      d(18)=>d_cache_arr_3_18, d(17)=>d_cache_arr_3_17, d(16)=>
      d_cache_arr_3_16, d(15)=>d_cache_arr_3_15, d(14)=>d_cache_arr_3_14, 
      d(13)=>d_cache_arr_3_13, d(12)=>d_cache_arr_3_12, d(11)=>
      d_cache_arr_3_11, d(10)=>d_cache_arr_3_10, d(9)=>d_cache_arr_3_9, d(8)
      =>d_cache_arr_3_8, d(7)=>d_cache_arr_3_7, d(6)=>d_cache_arr_3_6, d(5)
      =>d_cache_arr_3_5, d(4)=>d_cache_arr_3_4, d(3)=>d_cache_arr_3_3, d(2)
      =>d_cache_arr_3_2, d(1)=>d_cache_arr_3_1, d(0)=>d_cache_arr_3_0, q(31)
      =>q_cache_arr_3_31, q(30)=>q_cache_arr_3_30, q(29)=>q_cache_arr_3_29, 
      q(28)=>q_cache_arr_3_28, q(27)=>q_cache_arr_3_27, q(26)=>
      q_cache_arr_3_26, q(25)=>q_cache_arr_3_25, q(24)=>q_cache_arr_3_24, 
      q(23)=>q_cache_arr_3_23, q(22)=>q_cache_arr_3_22, q(21)=>
      q_cache_arr_3_21, q(20)=>q_cache_arr_3_20, q(19)=>q_cache_arr_3_19, 
      q(18)=>q_cache_arr_3_18, q(17)=>q_cache_arr_3_17, q(16)=>
      q_cache_arr_3_16, q(15)=>q_cache_arr_3_15, q(14)=>q_cache_arr_3_14, 
      q(13)=>q_cache_arr_3_13, q(12)=>q_cache_arr_3_12, q(11)=>
      q_cache_arr_3_11, q(10)=>q_cache_arr_3_10, q(9)=>q_cache_arr_3_9, q(8)
      =>q_cache_arr_3_8, q(7)=>q_cache_arr_3_7, q(6)=>q_cache_arr_3_6, q(5)
      =>q_cache_arr_3_5, q(4)=>q_cache_arr_3_4, q(3)=>q_cache_arr_3_3, q(2)
      =>q_cache_arr_3_2, q(1)=>q_cache_arr_3_1, q(0)=>q_cache_arr_3_0, 
      rst_data(31)=>buffer_ready_EXMPLR, rst_data(30)=>buffer_ready_EXMPLR, 
      rst_data(29)=>buffer_ready_EXMPLR, rst_data(28)=>buffer_ready_EXMPLR, 
      rst_data(27)=>buffer_ready_EXMPLR, rst_data(26)=>buffer_ready_EXMPLR, 
      rst_data(25)=>buffer_ready_EXMPLR, rst_data(24)=>buffer_ready_EXMPLR, 
      rst_data(23)=>buffer_ready_EXMPLR, rst_data(22)=>buffer_ready_EXMPLR, 
      rst_data(21)=>buffer_ready_EXMPLR, rst_data(20)=>buffer_ready_EXMPLR, 
      rst_data(19)=>buffer_ready_EXMPLR, rst_data(18)=>buffer_ready_EXMPLR, 
      rst_data(17)=>buffer_ready_EXMPLR, rst_data(16)=>buffer_ready_EXMPLR, 
      rst_data(15)=>buffer_ready_EXMPLR, rst_data(14)=>buffer_ready_EXMPLR, 
      rst_data(13)=>buffer_ready_EXMPLR, rst_data(12)=>buffer_ready_EXMPLR, 
      rst_data(11)=>buffer_ready_EXMPLR, rst_data(10)=>buffer_ready_EXMPLR, 
      rst_data(9)=>buffer_ready_EXMPLR, rst_data(8)=>buffer_ready_EXMPLR, 
      rst_data(7)=>buffer_ready_EXMPLR, rst_data(6)=>buffer_ready_EXMPLR, 
      rst_data(5)=>buffer_ready_EXMPLR, rst_data(4)=>buffer_ready_EXMPLR, 
      rst_data(3)=>buffer_ready_EXMPLR, rst_data(2)=>buffer_ready_EXMPLR, 
      rst_data(1)=>buffer_ready_EXMPLR, rst_data(0)=>buffer_ready_EXMPLR, 
      clk=>clk, load=>nx1109, reset=>filter_reset);
   gen_comp_cache_gen_regs_4_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_4_31, d(30)=>d_cache_arr_4_30, d(29)=>d_cache_arr_4_29, 
      d(28)=>d_cache_arr_4_28, d(27)=>d_cache_arr_4_27, d(26)=>
      d_cache_arr_4_26, d(25)=>d_cache_arr_4_25, d(24)=>d_cache_arr_4_24, 
      d(23)=>d_cache_arr_4_23, d(22)=>d_cache_arr_4_22, d(21)=>
      d_cache_arr_4_21, d(20)=>d_cache_arr_4_20, d(19)=>d_cache_arr_4_19, 
      d(18)=>d_cache_arr_4_18, d(17)=>d_cache_arr_4_17, d(16)=>
      d_cache_arr_4_16, d(15)=>d_cache_arr_4_15, d(14)=>d_cache_arr_4_14, 
      d(13)=>d_cache_arr_4_13, d(12)=>d_cache_arr_4_12, d(11)=>
      d_cache_arr_4_11, d(10)=>d_cache_arr_4_10, d(9)=>d_cache_arr_4_9, d(8)
      =>d_cache_arr_4_8, d(7)=>d_cache_arr_4_7, d(6)=>d_cache_arr_4_6, d(5)
      =>d_cache_arr_4_5, d(4)=>d_cache_arr_4_4, d(3)=>d_cache_arr_4_3, d(2)
      =>d_cache_arr_4_2, d(1)=>d_cache_arr_4_1, d(0)=>d_cache_arr_4_0, q(31)
      =>q_cache_arr_4_31, q(30)=>q_cache_arr_4_30, q(29)=>q_cache_arr_4_29, 
      q(28)=>q_cache_arr_4_28, q(27)=>q_cache_arr_4_27, q(26)=>
      q_cache_arr_4_26, q(25)=>q_cache_arr_4_25, q(24)=>q_cache_arr_4_24, 
      q(23)=>q_cache_arr_4_23, q(22)=>q_cache_arr_4_22, q(21)=>
      q_cache_arr_4_21, q(20)=>q_cache_arr_4_20, q(19)=>q_cache_arr_4_19, 
      q(18)=>q_cache_arr_4_18, q(17)=>q_cache_arr_4_17, q(16)=>
      q_cache_arr_4_16, q(15)=>q_cache_arr_4_15, q(14)=>q_cache_arr_4_14, 
      q(13)=>q_cache_arr_4_13, q(12)=>q_cache_arr_4_12, q(11)=>
      q_cache_arr_4_11, q(10)=>q_cache_arr_4_10, q(9)=>q_cache_arr_4_9, q(8)
      =>q_cache_arr_4_8, q(7)=>q_cache_arr_4_7, q(6)=>q_cache_arr_4_6, q(5)
      =>q_cache_arr_4_5, q(4)=>q_cache_arr_4_4, q(3)=>q_cache_arr_4_3, q(2)
      =>q_cache_arr_4_2, q(1)=>q_cache_arr_4_1, q(0)=>q_cache_arr_4_0, 
      rst_data(31)=>buffer_ready_EXMPLR, rst_data(30)=>buffer_ready_EXMPLR, 
      rst_data(29)=>buffer_ready_EXMPLR, rst_data(28)=>buffer_ready_EXMPLR, 
      rst_data(27)=>buffer_ready_EXMPLR, rst_data(26)=>buffer_ready_EXMPLR, 
      rst_data(25)=>buffer_ready_EXMPLR, rst_data(24)=>buffer_ready_EXMPLR, 
      rst_data(23)=>buffer_ready_EXMPLR, rst_data(22)=>buffer_ready_EXMPLR, 
      rst_data(21)=>buffer_ready_EXMPLR, rst_data(20)=>buffer_ready_EXMPLR, 
      rst_data(19)=>buffer_ready_EXMPLR, rst_data(18)=>buffer_ready_EXMPLR, 
      rst_data(17)=>buffer_ready_EXMPLR, rst_data(16)=>buffer_ready_EXMPLR, 
      rst_data(15)=>buffer_ready_EXMPLR, rst_data(14)=>buffer_ready_EXMPLR, 
      rst_data(13)=>buffer_ready_EXMPLR, rst_data(12)=>buffer_ready_EXMPLR, 
      rst_data(11)=>buffer_ready_EXMPLR, rst_data(10)=>buffer_ready_EXMPLR, 
      rst_data(9)=>buffer_ready_EXMPLR, rst_data(8)=>buffer_ready_EXMPLR, 
      rst_data(7)=>buffer_ready_EXMPLR, rst_data(6)=>buffer_ready_EXMPLR, 
      rst_data(5)=>buffer_ready_EXMPLR, rst_data(4)=>buffer_ready_EXMPLR, 
      rst_data(3)=>buffer_ready_EXMPLR, rst_data(2)=>buffer_ready_EXMPLR, 
      rst_data(1)=>buffer_ready_EXMPLR, rst_data(0)=>buffer_ready_EXMPLR, 
      clk=>clk, load=>nx1109, reset=>filter_reset);
   gen_comp_cache_gen_regs_5_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_5_31, d(30)=>d_cache_arr_5_30, d(29)=>d_cache_arr_5_29, 
      d(28)=>d_cache_arr_5_28, d(27)=>d_cache_arr_5_27, d(26)=>
      d_cache_arr_5_26, d(25)=>d_cache_arr_5_25, d(24)=>d_cache_arr_5_24, 
      d(23)=>d_cache_arr_5_23, d(22)=>d_cache_arr_5_22, d(21)=>
      d_cache_arr_5_21, d(20)=>d_cache_arr_5_20, d(19)=>d_cache_arr_5_19, 
      d(18)=>d_cache_arr_5_18, d(17)=>d_cache_arr_5_17, d(16)=>
      d_cache_arr_5_16, d(15)=>d_cache_arr_5_15, d(14)=>d_cache_arr_5_14, 
      d(13)=>d_cache_arr_5_13, d(12)=>d_cache_arr_5_12, d(11)=>
      d_cache_arr_5_11, d(10)=>d_cache_arr_5_10, d(9)=>d_cache_arr_5_9, d(8)
      =>d_cache_arr_5_8, d(7)=>d_cache_arr_5_7, d(6)=>d_cache_arr_5_6, d(5)
      =>d_cache_arr_5_5, d(4)=>d_cache_arr_5_4, d(3)=>d_cache_arr_5_3, d(2)
      =>d_cache_arr_5_2, d(1)=>d_cache_arr_5_1, d(0)=>d_cache_arr_5_0, q(31)
      =>q_cache_arr_5_31, q(30)=>q_cache_arr_5_30, q(29)=>q_cache_arr_5_29, 
      q(28)=>q_cache_arr_5_28, q(27)=>q_cache_arr_5_27, q(26)=>
      q_cache_arr_5_26, q(25)=>q_cache_arr_5_25, q(24)=>q_cache_arr_5_24, 
      q(23)=>q_cache_arr_5_23, q(22)=>q_cache_arr_5_22, q(21)=>
      q_cache_arr_5_21, q(20)=>q_cache_arr_5_20, q(19)=>q_cache_arr_5_19, 
      q(18)=>q_cache_arr_5_18, q(17)=>q_cache_arr_5_17, q(16)=>
      q_cache_arr_5_16, q(15)=>q_cache_arr_5_15, q(14)=>q_cache_arr_5_14, 
      q(13)=>q_cache_arr_5_13, q(12)=>q_cache_arr_5_12, q(11)=>
      q_cache_arr_5_11, q(10)=>q_cache_arr_5_10, q(9)=>q_cache_arr_5_9, q(8)
      =>q_cache_arr_5_8, q(7)=>q_cache_arr_5_7, q(6)=>q_cache_arr_5_6, q(5)
      =>q_cache_arr_5_5, q(4)=>q_cache_arr_5_4, q(3)=>q_cache_arr_5_3, q(2)
      =>q_cache_arr_5_2, q(1)=>q_cache_arr_5_1, q(0)=>q_cache_arr_5_0, 
      rst_data(31)=>buffer_ready_EXMPLR, rst_data(30)=>buffer_ready_EXMPLR, 
      rst_data(29)=>buffer_ready_EXMPLR, rst_data(28)=>buffer_ready_EXMPLR, 
      rst_data(27)=>buffer_ready_EXMPLR, rst_data(26)=>buffer_ready_EXMPLR, 
      rst_data(25)=>buffer_ready_EXMPLR, rst_data(24)=>buffer_ready_EXMPLR, 
      rst_data(23)=>buffer_ready_EXMPLR, rst_data(22)=>buffer_ready_EXMPLR, 
      rst_data(21)=>buffer_ready_EXMPLR, rst_data(20)=>buffer_ready_EXMPLR, 
      rst_data(19)=>buffer_ready_EXMPLR, rst_data(18)=>buffer_ready_EXMPLR, 
      rst_data(17)=>buffer_ready_EXMPLR, rst_data(16)=>buffer_ready_EXMPLR, 
      rst_data(15)=>buffer_ready_EXMPLR, rst_data(14)=>buffer_ready_EXMPLR, 
      rst_data(13)=>buffer_ready_EXMPLR, rst_data(12)=>buffer_ready_EXMPLR, 
      rst_data(11)=>buffer_ready_EXMPLR, rst_data(10)=>buffer_ready_EXMPLR, 
      rst_data(9)=>buffer_ready_EXMPLR, rst_data(8)=>buffer_ready_EXMPLR, 
      rst_data(7)=>buffer_ready_EXMPLR, rst_data(6)=>buffer_ready_EXMPLR, 
      rst_data(5)=>buffer_ready_EXMPLR, rst_data(4)=>buffer_ready_EXMPLR, 
      rst_data(3)=>buffer_ready_EXMPLR, rst_data(2)=>buffer_ready_EXMPLR, 
      rst_data(1)=>buffer_ready_EXMPLR, rst_data(0)=>buffer_ready_EXMPLR, 
      clk=>clk, load=>nx1109, reset=>filter_reset);
   gen_comp_cache_gen_regs_6_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_6_31, d(30)=>d_cache_arr_6_30, d(29)=>d_cache_arr_6_29, 
      d(28)=>d_cache_arr_6_28, d(27)=>d_cache_arr_6_27, d(26)=>
      d_cache_arr_6_26, d(25)=>d_cache_arr_6_25, d(24)=>d_cache_arr_6_24, 
      d(23)=>d_cache_arr_6_23, d(22)=>d_cache_arr_6_22, d(21)=>
      d_cache_arr_6_21, d(20)=>d_cache_arr_6_20, d(19)=>d_cache_arr_6_19, 
      d(18)=>d_cache_arr_6_18, d(17)=>d_cache_arr_6_17, d(16)=>
      d_cache_arr_6_16, d(15)=>d_cache_arr_6_15, d(14)=>d_cache_arr_6_14, 
      d(13)=>d_cache_arr_6_13, d(12)=>d_cache_arr_6_12, d(11)=>
      d_cache_arr_6_11, d(10)=>d_cache_arr_6_10, d(9)=>d_cache_arr_6_9, d(8)
      =>d_cache_arr_6_8, d(7)=>d_cache_arr_6_7, d(6)=>d_cache_arr_6_6, d(5)
      =>d_cache_arr_6_5, d(4)=>d_cache_arr_6_4, d(3)=>d_cache_arr_6_3, d(2)
      =>d_cache_arr_6_2, d(1)=>d_cache_arr_6_1, d(0)=>d_cache_arr_6_0, q(31)
      =>q_cache_arr_6_31, q(30)=>q_cache_arr_6_30, q(29)=>q_cache_arr_6_29, 
      q(28)=>q_cache_arr_6_28, q(27)=>q_cache_arr_6_27, q(26)=>
      q_cache_arr_6_26, q(25)=>q_cache_arr_6_25, q(24)=>q_cache_arr_6_24, 
      q(23)=>q_cache_arr_6_23, q(22)=>q_cache_arr_6_22, q(21)=>
      q_cache_arr_6_21, q(20)=>q_cache_arr_6_20, q(19)=>q_cache_arr_6_19, 
      q(18)=>q_cache_arr_6_18, q(17)=>q_cache_arr_6_17, q(16)=>
      q_cache_arr_6_16, q(15)=>q_cache_arr_6_15, q(14)=>q_cache_arr_6_14, 
      q(13)=>q_cache_arr_6_13, q(12)=>q_cache_arr_6_12, q(11)=>
      q_cache_arr_6_11, q(10)=>q_cache_arr_6_10, q(9)=>q_cache_arr_6_9, q(8)
      =>q_cache_arr_6_8, q(7)=>q_cache_arr_6_7, q(6)=>q_cache_arr_6_6, q(5)
      =>q_cache_arr_6_5, q(4)=>q_cache_arr_6_4, q(3)=>q_cache_arr_6_3, q(2)
      =>q_cache_arr_6_2, q(1)=>q_cache_arr_6_1, q(0)=>q_cache_arr_6_0, 
      rst_data(31)=>buffer_ready_EXMPLR, rst_data(30)=>buffer_ready_EXMPLR, 
      rst_data(29)=>buffer_ready_EXMPLR, rst_data(28)=>buffer_ready_EXMPLR, 
      rst_data(27)=>buffer_ready_EXMPLR, rst_data(26)=>buffer_ready_EXMPLR, 
      rst_data(25)=>buffer_ready_EXMPLR, rst_data(24)=>buffer_ready_EXMPLR, 
      rst_data(23)=>buffer_ready_EXMPLR, rst_data(22)=>buffer_ready_EXMPLR, 
      rst_data(21)=>buffer_ready_EXMPLR, rst_data(20)=>buffer_ready_EXMPLR, 
      rst_data(19)=>buffer_ready_EXMPLR, rst_data(18)=>buffer_ready_EXMPLR, 
      rst_data(17)=>buffer_ready_EXMPLR, rst_data(16)=>buffer_ready_EXMPLR, 
      rst_data(15)=>buffer_ready_EXMPLR, rst_data(14)=>buffer_ready_EXMPLR, 
      rst_data(13)=>buffer_ready_EXMPLR, rst_data(12)=>buffer_ready_EXMPLR, 
      rst_data(11)=>buffer_ready_EXMPLR, rst_data(10)=>buffer_ready_EXMPLR, 
      rst_data(9)=>buffer_ready_EXMPLR, rst_data(8)=>buffer_ready_EXMPLR, 
      rst_data(7)=>buffer_ready_EXMPLR, rst_data(6)=>buffer_ready_EXMPLR, 
      rst_data(5)=>buffer_ready_EXMPLR, rst_data(4)=>buffer_ready_EXMPLR, 
      rst_data(3)=>buffer_ready_EXMPLR, rst_data(2)=>buffer_ready_EXMPLR, 
      rst_data(1)=>buffer_ready_EXMPLR, rst_data(0)=>buffer_ready_EXMPLR, 
      clk=>clk, load=>nx1109, reset=>filter_reset);
   gen_comp_cache_gen_regs_7_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_7_31, d(30)=>d_cache_arr_7_30, d(29)=>d_cache_arr_7_29, 
      d(28)=>d_cache_arr_7_28, d(27)=>d_cache_arr_7_27, d(26)=>
      d_cache_arr_7_26, d(25)=>d_cache_arr_7_25, d(24)=>d_cache_arr_7_24, 
      d(23)=>d_cache_arr_7_23, d(22)=>d_cache_arr_7_22, d(21)=>
      d_cache_arr_7_21, d(20)=>d_cache_arr_7_20, d(19)=>d_cache_arr_7_19, 
      d(18)=>d_cache_arr_7_18, d(17)=>d_cache_arr_7_17, d(16)=>
      d_cache_arr_7_16, d(15)=>d_cache_arr_7_15, d(14)=>d_cache_arr_7_14, 
      d(13)=>d_cache_arr_7_13, d(12)=>d_cache_arr_7_12, d(11)=>
      d_cache_arr_7_11, d(10)=>d_cache_arr_7_10, d(9)=>d_cache_arr_7_9, d(8)
      =>d_cache_arr_7_8, d(7)=>d_cache_arr_7_7, d(6)=>d_cache_arr_7_6, d(5)
      =>d_cache_arr_7_5, d(4)=>d_cache_arr_7_4, d(3)=>d_cache_arr_7_3, d(2)
      =>d_cache_arr_7_2, d(1)=>d_cache_arr_7_1, d(0)=>d_cache_arr_7_0, q(31)
      =>q_cache_arr_7_31, q(30)=>q_cache_arr_7_30, q(29)=>q_cache_arr_7_29, 
      q(28)=>q_cache_arr_7_28, q(27)=>q_cache_arr_7_27, q(26)=>
      q_cache_arr_7_26, q(25)=>q_cache_arr_7_25, q(24)=>q_cache_arr_7_24, 
      q(23)=>q_cache_arr_7_23, q(22)=>q_cache_arr_7_22, q(21)=>
      q_cache_arr_7_21, q(20)=>q_cache_arr_7_20, q(19)=>q_cache_arr_7_19, 
      q(18)=>q_cache_arr_7_18, q(17)=>q_cache_arr_7_17, q(16)=>
      q_cache_arr_7_16, q(15)=>q_cache_arr_7_15, q(14)=>q_cache_arr_7_14, 
      q(13)=>q_cache_arr_7_13, q(12)=>q_cache_arr_7_12, q(11)=>
      q_cache_arr_7_11, q(10)=>q_cache_arr_7_10, q(9)=>q_cache_arr_7_9, q(8)
      =>q_cache_arr_7_8, q(7)=>q_cache_arr_7_7, q(6)=>q_cache_arr_7_6, q(5)
      =>q_cache_arr_7_5, q(4)=>q_cache_arr_7_4, q(3)=>q_cache_arr_7_3, q(2)
      =>q_cache_arr_7_2, q(1)=>q_cache_arr_7_1, q(0)=>q_cache_arr_7_0, 
      rst_data(31)=>buffer_ready_EXMPLR, rst_data(30)=>buffer_ready_EXMPLR, 
      rst_data(29)=>buffer_ready_EXMPLR, rst_data(28)=>buffer_ready_EXMPLR, 
      rst_data(27)=>buffer_ready_EXMPLR, rst_data(26)=>buffer_ready_EXMPLR, 
      rst_data(25)=>buffer_ready_EXMPLR, rst_data(24)=>buffer_ready_EXMPLR, 
      rst_data(23)=>buffer_ready_EXMPLR, rst_data(22)=>buffer_ready_EXMPLR, 
      rst_data(21)=>buffer_ready_EXMPLR, rst_data(20)=>buffer_ready_EXMPLR, 
      rst_data(19)=>buffer_ready_EXMPLR, rst_data(18)=>buffer_ready_EXMPLR, 
      rst_data(17)=>buffer_ready_EXMPLR, rst_data(16)=>buffer_ready_EXMPLR, 
      rst_data(15)=>buffer_ready_EXMPLR, rst_data(14)=>buffer_ready_EXMPLR, 
      rst_data(13)=>buffer_ready_EXMPLR, rst_data(12)=>buffer_ready_EXMPLR, 
      rst_data(11)=>buffer_ready_EXMPLR, rst_data(10)=>buffer_ready_EXMPLR, 
      rst_data(9)=>buffer_ready_EXMPLR, rst_data(8)=>buffer_ready_EXMPLR, 
      rst_data(7)=>buffer_ready_EXMPLR, rst_data(6)=>buffer_ready_EXMPLR, 
      rst_data(5)=>buffer_ready_EXMPLR, rst_data(4)=>buffer_ready_EXMPLR, 
      rst_data(3)=>buffer_ready_EXMPLR, rst_data(2)=>buffer_ready_EXMPLR, 
      rst_data(1)=>buffer_ready_EXMPLR, rst_data(0)=>buffer_ready_EXMPLR, 
      clk=>clk, load=>nx1111, reset=>filter_reset);
   gen_comp_cache_gen_regs_8_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_8_31, d(30)=>d_cache_arr_8_30, d(29)=>d_cache_arr_8_29, 
      d(28)=>d_cache_arr_8_28, d(27)=>d_cache_arr_8_27, d(26)=>
      d_cache_arr_8_26, d(25)=>d_cache_arr_8_25, d(24)=>d_cache_arr_8_24, 
      d(23)=>d_cache_arr_8_23, d(22)=>d_cache_arr_8_22, d(21)=>
      d_cache_arr_8_21, d(20)=>d_cache_arr_8_20, d(19)=>d_cache_arr_8_19, 
      d(18)=>d_cache_arr_8_18, d(17)=>d_cache_arr_8_17, d(16)=>
      d_cache_arr_8_16, d(15)=>d_cache_arr_8_15, d(14)=>d_cache_arr_8_14, 
      d(13)=>d_cache_arr_8_13, d(12)=>d_cache_arr_8_12, d(11)=>
      d_cache_arr_8_11, d(10)=>d_cache_arr_8_10, d(9)=>d_cache_arr_8_9, d(8)
      =>d_cache_arr_8_8, d(7)=>d_cache_arr_8_7, d(6)=>d_cache_arr_8_6, d(5)
      =>d_cache_arr_8_5, d(4)=>d_cache_arr_8_4, d(3)=>d_cache_arr_8_3, d(2)
      =>d_cache_arr_8_2, d(1)=>d_cache_arr_8_1, d(0)=>d_cache_arr_8_0, q(31)
      =>q_cache_arr_8_31, q(30)=>q_cache_arr_8_30, q(29)=>q_cache_arr_8_29, 
      q(28)=>q_cache_arr_8_28, q(27)=>q_cache_arr_8_27, q(26)=>
      q_cache_arr_8_26, q(25)=>q_cache_arr_8_25, q(24)=>q_cache_arr_8_24, 
      q(23)=>q_cache_arr_8_23, q(22)=>q_cache_arr_8_22, q(21)=>
      q_cache_arr_8_21, q(20)=>q_cache_arr_8_20, q(19)=>q_cache_arr_8_19, 
      q(18)=>q_cache_arr_8_18, q(17)=>q_cache_arr_8_17, q(16)=>
      q_cache_arr_8_16, q(15)=>q_cache_arr_8_15, q(14)=>q_cache_arr_8_14, 
      q(13)=>q_cache_arr_8_13, q(12)=>q_cache_arr_8_12, q(11)=>
      q_cache_arr_8_11, q(10)=>q_cache_arr_8_10, q(9)=>q_cache_arr_8_9, q(8)
      =>q_cache_arr_8_8, q(7)=>q_cache_arr_8_7, q(6)=>q_cache_arr_8_6, q(5)
      =>q_cache_arr_8_5, q(4)=>q_cache_arr_8_4, q(3)=>q_cache_arr_8_3, q(2)
      =>q_cache_arr_8_2, q(1)=>q_cache_arr_8_1, q(0)=>q_cache_arr_8_0, 
      rst_data(31)=>buffer_ready_EXMPLR, rst_data(30)=>buffer_ready_EXMPLR, 
      rst_data(29)=>buffer_ready_EXMPLR, rst_data(28)=>buffer_ready_EXMPLR, 
      rst_data(27)=>buffer_ready_EXMPLR, rst_data(26)=>buffer_ready_EXMPLR, 
      rst_data(25)=>buffer_ready_EXMPLR, rst_data(24)=>buffer_ready_EXMPLR, 
      rst_data(23)=>buffer_ready_EXMPLR, rst_data(22)=>buffer_ready_EXMPLR, 
      rst_data(21)=>buffer_ready_EXMPLR, rst_data(20)=>buffer_ready_EXMPLR, 
      rst_data(19)=>buffer_ready_EXMPLR, rst_data(18)=>buffer_ready_EXMPLR, 
      rst_data(17)=>buffer_ready_EXMPLR, rst_data(16)=>buffer_ready_EXMPLR, 
      rst_data(15)=>buffer_ready_EXMPLR, rst_data(14)=>buffer_ready_EXMPLR, 
      rst_data(13)=>buffer_ready_EXMPLR, rst_data(12)=>buffer_ready_EXMPLR, 
      rst_data(11)=>buffer_ready_EXMPLR, rst_data(10)=>buffer_ready_EXMPLR, 
      rst_data(9)=>buffer_ready_EXMPLR, rst_data(8)=>buffer_ready_EXMPLR, 
      rst_data(7)=>buffer_ready_EXMPLR, rst_data(6)=>buffer_ready_EXMPLR, 
      rst_data(5)=>buffer_ready_EXMPLR, rst_data(4)=>buffer_ready_EXMPLR, 
      rst_data(3)=>buffer_ready_EXMPLR, rst_data(2)=>buffer_ready_EXMPLR, 
      rst_data(1)=>buffer_ready_EXMPLR, rst_data(0)=>buffer_ready_EXMPLR, 
      clk=>clk, load=>nx1111, reset=>filter_reset);
   gen_comp_cache_gen_regs_9_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_9_31, d(30)=>d_cache_arr_9_30, d(29)=>d_cache_arr_9_29, 
      d(28)=>d_cache_arr_9_28, d(27)=>d_cache_arr_9_27, d(26)=>
      d_cache_arr_9_26, d(25)=>d_cache_arr_9_25, d(24)=>d_cache_arr_9_24, 
      d(23)=>d_cache_arr_9_23, d(22)=>d_cache_arr_9_22, d(21)=>
      d_cache_arr_9_21, d(20)=>d_cache_arr_9_20, d(19)=>d_cache_arr_9_19, 
      d(18)=>d_cache_arr_9_18, d(17)=>d_cache_arr_9_17, d(16)=>
      d_cache_arr_9_16, d(15)=>d_cache_arr_9_15, d(14)=>d_cache_arr_9_14, 
      d(13)=>d_cache_arr_9_13, d(12)=>d_cache_arr_9_12, d(11)=>
      d_cache_arr_9_11, d(10)=>d_cache_arr_9_10, d(9)=>d_cache_arr_9_9, d(8)
      =>d_cache_arr_9_8, d(7)=>d_cache_arr_9_7, d(6)=>d_cache_arr_9_6, d(5)
      =>d_cache_arr_9_5, d(4)=>d_cache_arr_9_4, d(3)=>d_cache_arr_9_3, d(2)
      =>d_cache_arr_9_2, d(1)=>d_cache_arr_9_1, d(0)=>d_cache_arr_9_0, q(31)
      =>q_cache_arr_9_31, q(30)=>q_cache_arr_9_30, q(29)=>q_cache_arr_9_29, 
      q(28)=>q_cache_arr_9_28, q(27)=>q_cache_arr_9_27, q(26)=>
      q_cache_arr_9_26, q(25)=>q_cache_arr_9_25, q(24)=>q_cache_arr_9_24, 
      q(23)=>q_cache_arr_9_23, q(22)=>q_cache_arr_9_22, q(21)=>
      q_cache_arr_9_21, q(20)=>q_cache_arr_9_20, q(19)=>q_cache_arr_9_19, 
      q(18)=>q_cache_arr_9_18, q(17)=>q_cache_arr_9_17, q(16)=>
      q_cache_arr_9_16, q(15)=>q_cache_arr_9_15, q(14)=>q_cache_arr_9_14, 
      q(13)=>q_cache_arr_9_13, q(12)=>q_cache_arr_9_12, q(11)=>
      q_cache_arr_9_11, q(10)=>q_cache_arr_9_10, q(9)=>q_cache_arr_9_9, q(8)
      =>q_cache_arr_9_8, q(7)=>q_cache_arr_9_7, q(6)=>q_cache_arr_9_6, q(5)
      =>q_cache_arr_9_5, q(4)=>q_cache_arr_9_4, q(3)=>q_cache_arr_9_3, q(2)
      =>q_cache_arr_9_2, q(1)=>q_cache_arr_9_1, q(0)=>q_cache_arr_9_0, 
      rst_data(31)=>buffer_ready_EXMPLR, rst_data(30)=>buffer_ready_EXMPLR, 
      rst_data(29)=>buffer_ready_EXMPLR, rst_data(28)=>buffer_ready_EXMPLR, 
      rst_data(27)=>buffer_ready_EXMPLR, rst_data(26)=>buffer_ready_EXMPLR, 
      rst_data(25)=>buffer_ready_EXMPLR, rst_data(24)=>buffer_ready_EXMPLR, 
      rst_data(23)=>buffer_ready_EXMPLR, rst_data(22)=>buffer_ready_EXMPLR, 
      rst_data(21)=>buffer_ready_EXMPLR, rst_data(20)=>buffer_ready_EXMPLR, 
      rst_data(19)=>buffer_ready_EXMPLR, rst_data(18)=>buffer_ready_EXMPLR, 
      rst_data(17)=>buffer_ready_EXMPLR, rst_data(16)=>buffer_ready_EXMPLR, 
      rst_data(15)=>buffer_ready_EXMPLR, rst_data(14)=>buffer_ready_EXMPLR, 
      rst_data(13)=>buffer_ready_EXMPLR, rst_data(12)=>buffer_ready_EXMPLR, 
      rst_data(11)=>buffer_ready_EXMPLR, rst_data(10)=>buffer_ready_EXMPLR, 
      rst_data(9)=>buffer_ready_EXMPLR, rst_data(8)=>buffer_ready_EXMPLR, 
      rst_data(7)=>buffer_ready_EXMPLR, rst_data(6)=>buffer_ready_EXMPLR, 
      rst_data(5)=>buffer_ready_EXMPLR, rst_data(4)=>buffer_ready_EXMPLR, 
      rst_data(3)=>buffer_ready_EXMPLR, rst_data(2)=>buffer_ready_EXMPLR, 
      rst_data(1)=>buffer_ready_EXMPLR, rst_data(0)=>buffer_ready_EXMPLR, 
      clk=>clk, load=>nx1111, reset=>filter_reset);
   gen_comp_cache_gen_regs_10_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_10_31, d(30)=>d_cache_arr_10_30, d(29)=>d_cache_arr_10_29, 
      d(28)=>d_cache_arr_10_28, d(27)=>d_cache_arr_10_27, d(26)=>
      d_cache_arr_10_26, d(25)=>d_cache_arr_10_25, d(24)=>d_cache_arr_10_24, 
      d(23)=>d_cache_arr_10_23, d(22)=>d_cache_arr_10_22, d(21)=>
      d_cache_arr_10_21, d(20)=>d_cache_arr_10_20, d(19)=>d_cache_arr_10_19, 
      d(18)=>d_cache_arr_10_18, d(17)=>d_cache_arr_10_17, d(16)=>
      d_cache_arr_10_16, d(15)=>d_cache_arr_10_15, d(14)=>d_cache_arr_10_14, 
      d(13)=>d_cache_arr_10_13, d(12)=>d_cache_arr_10_12, d(11)=>
      d_cache_arr_10_11, d(10)=>d_cache_arr_10_10, d(9)=>d_cache_arr_10_9, 
      d(8)=>d_cache_arr_10_8, d(7)=>d_cache_arr_10_7, d(6)=>d_cache_arr_10_6, 
      d(5)=>d_cache_arr_10_5, d(4)=>d_cache_arr_10_4, d(3)=>d_cache_arr_10_3, 
      d(2)=>d_cache_arr_10_2, d(1)=>d_cache_arr_10_1, d(0)=>d_cache_arr_10_0, 
      q(31)=>q_cache_arr_10_31, q(30)=>q_cache_arr_10_30, q(29)=>
      q_cache_arr_10_29, q(28)=>q_cache_arr_10_28, q(27)=>q_cache_arr_10_27, 
      q(26)=>q_cache_arr_10_26, q(25)=>q_cache_arr_10_25, q(24)=>
      q_cache_arr_10_24, q(23)=>q_cache_arr_10_23, q(22)=>q_cache_arr_10_22, 
      q(21)=>q_cache_arr_10_21, q(20)=>q_cache_arr_10_20, q(19)=>
      q_cache_arr_10_19, q(18)=>q_cache_arr_10_18, q(17)=>q_cache_arr_10_17, 
      q(16)=>q_cache_arr_10_16, q(15)=>q_cache_arr_10_15, q(14)=>
      q_cache_arr_10_14, q(13)=>q_cache_arr_10_13, q(12)=>q_cache_arr_10_12, 
      q(11)=>q_cache_arr_10_11, q(10)=>q_cache_arr_10_10, q(9)=>
      q_cache_arr_10_9, q(8)=>q_cache_arr_10_8, q(7)=>q_cache_arr_10_7, q(6)
      =>q_cache_arr_10_6, q(5)=>q_cache_arr_10_5, q(4)=>q_cache_arr_10_4, 
      q(3)=>q_cache_arr_10_3, q(2)=>q_cache_arr_10_2, q(1)=>q_cache_arr_10_1, 
      q(0)=>q_cache_arr_10_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1111, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_11_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_11_31, d(30)=>d_cache_arr_11_30, d(29)=>d_cache_arr_11_29, 
      d(28)=>d_cache_arr_11_28, d(27)=>d_cache_arr_11_27, d(26)=>
      d_cache_arr_11_26, d(25)=>d_cache_arr_11_25, d(24)=>d_cache_arr_11_24, 
      d(23)=>d_cache_arr_11_23, d(22)=>d_cache_arr_11_22, d(21)=>
      d_cache_arr_11_21, d(20)=>d_cache_arr_11_20, d(19)=>d_cache_arr_11_19, 
      d(18)=>d_cache_arr_11_18, d(17)=>d_cache_arr_11_17, d(16)=>
      d_cache_arr_11_16, d(15)=>d_cache_arr_11_15, d(14)=>d_cache_arr_11_14, 
      d(13)=>d_cache_arr_11_13, d(12)=>d_cache_arr_11_12, d(11)=>
      d_cache_arr_11_11, d(10)=>d_cache_arr_11_10, d(9)=>d_cache_arr_11_9, 
      d(8)=>d_cache_arr_11_8, d(7)=>d_cache_arr_11_7, d(6)=>d_cache_arr_11_6, 
      d(5)=>d_cache_arr_11_5, d(4)=>d_cache_arr_11_4, d(3)=>d_cache_arr_11_3, 
      d(2)=>d_cache_arr_11_2, d(1)=>d_cache_arr_11_1, d(0)=>d_cache_arr_11_0, 
      q(31)=>q_cache_arr_11_31, q(30)=>q_cache_arr_11_30, q(29)=>
      q_cache_arr_11_29, q(28)=>q_cache_arr_11_28, q(27)=>q_cache_arr_11_27, 
      q(26)=>q_cache_arr_11_26, q(25)=>q_cache_arr_11_25, q(24)=>
      q_cache_arr_11_24, q(23)=>q_cache_arr_11_23, q(22)=>q_cache_arr_11_22, 
      q(21)=>q_cache_arr_11_21, q(20)=>q_cache_arr_11_20, q(19)=>
      q_cache_arr_11_19, q(18)=>q_cache_arr_11_18, q(17)=>q_cache_arr_11_17, 
      q(16)=>q_cache_arr_11_16, q(15)=>q_cache_arr_11_15, q(14)=>
      q_cache_arr_11_14, q(13)=>q_cache_arr_11_13, q(12)=>q_cache_arr_11_12, 
      q(11)=>q_cache_arr_11_11, q(10)=>q_cache_arr_11_10, q(9)=>
      q_cache_arr_11_9, q(8)=>q_cache_arr_11_8, q(7)=>q_cache_arr_11_7, q(6)
      =>q_cache_arr_11_6, q(5)=>q_cache_arr_11_5, q(4)=>q_cache_arr_11_4, 
      q(3)=>q_cache_arr_11_3, q(2)=>q_cache_arr_11_2, q(1)=>q_cache_arr_11_1, 
      q(0)=>q_cache_arr_11_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1111, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_12_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_12_31, d(30)=>d_cache_arr_12_30, d(29)=>d_cache_arr_12_29, 
      d(28)=>d_cache_arr_12_28, d(27)=>d_cache_arr_12_27, d(26)=>
      d_cache_arr_12_26, d(25)=>d_cache_arr_12_25, d(24)=>d_cache_arr_12_24, 
      d(23)=>d_cache_arr_12_23, d(22)=>d_cache_arr_12_22, d(21)=>
      d_cache_arr_12_21, d(20)=>d_cache_arr_12_20, d(19)=>d_cache_arr_12_19, 
      d(18)=>d_cache_arr_12_18, d(17)=>d_cache_arr_12_17, d(16)=>
      d_cache_arr_12_16, d(15)=>d_cache_arr_12_15, d(14)=>d_cache_arr_12_14, 
      d(13)=>d_cache_arr_12_13, d(12)=>d_cache_arr_12_12, d(11)=>
      d_cache_arr_12_11, d(10)=>d_cache_arr_12_10, d(9)=>d_cache_arr_12_9, 
      d(8)=>d_cache_arr_12_8, d(7)=>d_cache_arr_12_7, d(6)=>d_cache_arr_12_6, 
      d(5)=>d_cache_arr_12_5, d(4)=>d_cache_arr_12_4, d(3)=>d_cache_arr_12_3, 
      d(2)=>d_cache_arr_12_2, d(1)=>d_cache_arr_12_1, d(0)=>d_cache_arr_12_0, 
      q(31)=>q_cache_arr_12_31, q(30)=>q_cache_arr_12_30, q(29)=>
      q_cache_arr_12_29, q(28)=>q_cache_arr_12_28, q(27)=>q_cache_arr_12_27, 
      q(26)=>q_cache_arr_12_26, q(25)=>q_cache_arr_12_25, q(24)=>
      q_cache_arr_12_24, q(23)=>q_cache_arr_12_23, q(22)=>q_cache_arr_12_22, 
      q(21)=>q_cache_arr_12_21, q(20)=>q_cache_arr_12_20, q(19)=>
      q_cache_arr_12_19, q(18)=>q_cache_arr_12_18, q(17)=>q_cache_arr_12_17, 
      q(16)=>q_cache_arr_12_16, q(15)=>q_cache_arr_12_15, q(14)=>
      q_cache_arr_12_14, q(13)=>q_cache_arr_12_13, q(12)=>q_cache_arr_12_12, 
      q(11)=>q_cache_arr_12_11, q(10)=>q_cache_arr_12_10, q(9)=>
      q_cache_arr_12_9, q(8)=>q_cache_arr_12_8, q(7)=>q_cache_arr_12_7, q(6)
      =>q_cache_arr_12_6, q(5)=>q_cache_arr_12_5, q(4)=>q_cache_arr_12_4, 
      q(3)=>q_cache_arr_12_3, q(2)=>q_cache_arr_12_2, q(1)=>q_cache_arr_12_1, 
      q(0)=>q_cache_arr_12_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1111, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_13_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_13_31, d(30)=>d_cache_arr_13_30, d(29)=>d_cache_arr_13_29, 
      d(28)=>d_cache_arr_13_28, d(27)=>d_cache_arr_13_27, d(26)=>
      d_cache_arr_13_26, d(25)=>d_cache_arr_13_25, d(24)=>d_cache_arr_13_24, 
      d(23)=>d_cache_arr_13_23, d(22)=>d_cache_arr_13_22, d(21)=>
      d_cache_arr_13_21, d(20)=>d_cache_arr_13_20, d(19)=>d_cache_arr_13_19, 
      d(18)=>d_cache_arr_13_18, d(17)=>d_cache_arr_13_17, d(16)=>
      d_cache_arr_13_16, d(15)=>d_cache_arr_13_15, d(14)=>d_cache_arr_13_14, 
      d(13)=>d_cache_arr_13_13, d(12)=>d_cache_arr_13_12, d(11)=>
      d_cache_arr_13_11, d(10)=>d_cache_arr_13_10, d(9)=>d_cache_arr_13_9, 
      d(8)=>d_cache_arr_13_8, d(7)=>d_cache_arr_13_7, d(6)=>d_cache_arr_13_6, 
      d(5)=>d_cache_arr_13_5, d(4)=>d_cache_arr_13_4, d(3)=>d_cache_arr_13_3, 
      d(2)=>d_cache_arr_13_2, d(1)=>d_cache_arr_13_1, d(0)=>d_cache_arr_13_0, 
      q(31)=>q_cache_arr_13_31, q(30)=>q_cache_arr_13_30, q(29)=>
      q_cache_arr_13_29, q(28)=>q_cache_arr_13_28, q(27)=>q_cache_arr_13_27, 
      q(26)=>q_cache_arr_13_26, q(25)=>q_cache_arr_13_25, q(24)=>
      q_cache_arr_13_24, q(23)=>q_cache_arr_13_23, q(22)=>q_cache_arr_13_22, 
      q(21)=>q_cache_arr_13_21, q(20)=>q_cache_arr_13_20, q(19)=>
      q_cache_arr_13_19, q(18)=>q_cache_arr_13_18, q(17)=>q_cache_arr_13_17, 
      q(16)=>q_cache_arr_13_16, q(15)=>q_cache_arr_13_15, q(14)=>
      q_cache_arr_13_14, q(13)=>q_cache_arr_13_13, q(12)=>q_cache_arr_13_12, 
      q(11)=>q_cache_arr_13_11, q(10)=>q_cache_arr_13_10, q(9)=>
      q_cache_arr_13_9, q(8)=>q_cache_arr_13_8, q(7)=>q_cache_arr_13_7, q(6)
      =>q_cache_arr_13_6, q(5)=>q_cache_arr_13_5, q(4)=>q_cache_arr_13_4, 
      q(3)=>q_cache_arr_13_3, q(2)=>q_cache_arr_13_2, q(1)=>q_cache_arr_13_1, 
      q(0)=>q_cache_arr_13_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1111, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_14_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_14_31, d(30)=>d_cache_arr_14_30, d(29)=>d_cache_arr_14_29, 
      d(28)=>d_cache_arr_14_28, d(27)=>d_cache_arr_14_27, d(26)=>
      d_cache_arr_14_26, d(25)=>d_cache_arr_14_25, d(24)=>d_cache_arr_14_24, 
      d(23)=>d_cache_arr_14_23, d(22)=>d_cache_arr_14_22, d(21)=>
      d_cache_arr_14_21, d(20)=>d_cache_arr_14_20, d(19)=>d_cache_arr_14_19, 
      d(18)=>d_cache_arr_14_18, d(17)=>d_cache_arr_14_17, d(16)=>
      d_cache_arr_14_16, d(15)=>d_cache_arr_14_15, d(14)=>d_cache_arr_14_14, 
      d(13)=>d_cache_arr_14_13, d(12)=>d_cache_arr_14_12, d(11)=>
      d_cache_arr_14_11, d(10)=>d_cache_arr_14_10, d(9)=>d_cache_arr_14_9, 
      d(8)=>d_cache_arr_14_8, d(7)=>d_cache_arr_14_7, d(6)=>d_cache_arr_14_6, 
      d(5)=>d_cache_arr_14_5, d(4)=>d_cache_arr_14_4, d(3)=>d_cache_arr_14_3, 
      d(2)=>d_cache_arr_14_2, d(1)=>d_cache_arr_14_1, d(0)=>d_cache_arr_14_0, 
      q(31)=>q_cache_arr_14_31, q(30)=>q_cache_arr_14_30, q(29)=>
      q_cache_arr_14_29, q(28)=>q_cache_arr_14_28, q(27)=>q_cache_arr_14_27, 
      q(26)=>q_cache_arr_14_26, q(25)=>q_cache_arr_14_25, q(24)=>
      q_cache_arr_14_24, q(23)=>q_cache_arr_14_23, q(22)=>q_cache_arr_14_22, 
      q(21)=>q_cache_arr_14_21, q(20)=>q_cache_arr_14_20, q(19)=>
      q_cache_arr_14_19, q(18)=>q_cache_arr_14_18, q(17)=>q_cache_arr_14_17, 
      q(16)=>q_cache_arr_14_16, q(15)=>q_cache_arr_14_15, q(14)=>
      q_cache_arr_14_14, q(13)=>q_cache_arr_14_13, q(12)=>q_cache_arr_14_12, 
      q(11)=>q_cache_arr_14_11, q(10)=>q_cache_arr_14_10, q(9)=>
      q_cache_arr_14_9, q(8)=>q_cache_arr_14_8, q(7)=>q_cache_arr_14_7, q(6)
      =>q_cache_arr_14_6, q(5)=>q_cache_arr_14_5, q(4)=>q_cache_arr_14_4, 
      q(3)=>q_cache_arr_14_3, q(2)=>q_cache_arr_14_2, q(1)=>q_cache_arr_14_1, 
      q(0)=>q_cache_arr_14_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1113, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_15_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_15_31, d(30)=>d_cache_arr_15_30, d(29)=>d_cache_arr_15_29, 
      d(28)=>d_cache_arr_15_28, d(27)=>d_cache_arr_15_27, d(26)=>
      d_cache_arr_15_26, d(25)=>d_cache_arr_15_25, d(24)=>d_cache_arr_15_24, 
      d(23)=>d_cache_arr_15_23, d(22)=>d_cache_arr_15_22, d(21)=>
      d_cache_arr_15_21, d(20)=>d_cache_arr_15_20, d(19)=>d_cache_arr_15_19, 
      d(18)=>d_cache_arr_15_18, d(17)=>d_cache_arr_15_17, d(16)=>
      d_cache_arr_15_16, d(15)=>d_cache_arr_15_15, d(14)=>d_cache_arr_15_14, 
      d(13)=>d_cache_arr_15_13, d(12)=>d_cache_arr_15_12, d(11)=>
      d_cache_arr_15_11, d(10)=>d_cache_arr_15_10, d(9)=>d_cache_arr_15_9, 
      d(8)=>d_cache_arr_15_8, d(7)=>d_cache_arr_15_7, d(6)=>d_cache_arr_15_6, 
      d(5)=>d_cache_arr_15_5, d(4)=>d_cache_arr_15_4, d(3)=>d_cache_arr_15_3, 
      d(2)=>d_cache_arr_15_2, d(1)=>d_cache_arr_15_1, d(0)=>d_cache_arr_15_0, 
      q(31)=>q_cache_arr_15_31, q(30)=>q_cache_arr_15_30, q(29)=>
      q_cache_arr_15_29, q(28)=>q_cache_arr_15_28, q(27)=>q_cache_arr_15_27, 
      q(26)=>q_cache_arr_15_26, q(25)=>q_cache_arr_15_25, q(24)=>
      q_cache_arr_15_24, q(23)=>q_cache_arr_15_23, q(22)=>q_cache_arr_15_22, 
      q(21)=>q_cache_arr_15_21, q(20)=>q_cache_arr_15_20, q(19)=>
      q_cache_arr_15_19, q(18)=>q_cache_arr_15_18, q(17)=>q_cache_arr_15_17, 
      q(16)=>q_cache_arr_15_16, q(15)=>q_cache_arr_15_15, q(14)=>
      q_cache_arr_15_14, q(13)=>q_cache_arr_15_13, q(12)=>q_cache_arr_15_12, 
      q(11)=>q_cache_arr_15_11, q(10)=>q_cache_arr_15_10, q(9)=>
      q_cache_arr_15_9, q(8)=>q_cache_arr_15_8, q(7)=>q_cache_arr_15_7, q(6)
      =>q_cache_arr_15_6, q(5)=>q_cache_arr_15_5, q(4)=>q_cache_arr_15_4, 
      q(3)=>q_cache_arr_15_3, q(2)=>q_cache_arr_15_2, q(1)=>q_cache_arr_15_1, 
      q(0)=>q_cache_arr_15_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1113, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_16_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_16_31, d(30)=>d_cache_arr_16_30, d(29)=>d_cache_arr_16_29, 
      d(28)=>d_cache_arr_16_28, d(27)=>d_cache_arr_16_27, d(26)=>
      d_cache_arr_16_26, d(25)=>d_cache_arr_16_25, d(24)=>d_cache_arr_16_24, 
      d(23)=>d_cache_arr_16_23, d(22)=>d_cache_arr_16_22, d(21)=>
      d_cache_arr_16_21, d(20)=>d_cache_arr_16_20, d(19)=>d_cache_arr_16_19, 
      d(18)=>d_cache_arr_16_18, d(17)=>d_cache_arr_16_17, d(16)=>
      d_cache_arr_16_16, d(15)=>d_cache_arr_16_15, d(14)=>d_cache_arr_16_14, 
      d(13)=>d_cache_arr_16_13, d(12)=>d_cache_arr_16_12, d(11)=>
      d_cache_arr_16_11, d(10)=>d_cache_arr_16_10, d(9)=>d_cache_arr_16_9, 
      d(8)=>d_cache_arr_16_8, d(7)=>d_cache_arr_16_7, d(6)=>d_cache_arr_16_6, 
      d(5)=>d_cache_arr_16_5, d(4)=>d_cache_arr_16_4, d(3)=>d_cache_arr_16_3, 
      d(2)=>d_cache_arr_16_2, d(1)=>d_cache_arr_16_1, d(0)=>d_cache_arr_16_0, 
      q(31)=>q_cache_arr_16_31, q(30)=>q_cache_arr_16_30, q(29)=>
      q_cache_arr_16_29, q(28)=>q_cache_arr_16_28, q(27)=>q_cache_arr_16_27, 
      q(26)=>q_cache_arr_16_26, q(25)=>q_cache_arr_16_25, q(24)=>
      q_cache_arr_16_24, q(23)=>q_cache_arr_16_23, q(22)=>q_cache_arr_16_22, 
      q(21)=>q_cache_arr_16_21, q(20)=>q_cache_arr_16_20, q(19)=>
      q_cache_arr_16_19, q(18)=>q_cache_arr_16_18, q(17)=>q_cache_arr_16_17, 
      q(16)=>q_cache_arr_16_16, q(15)=>q_cache_arr_16_15, q(14)=>
      q_cache_arr_16_14, q(13)=>q_cache_arr_16_13, q(12)=>q_cache_arr_16_12, 
      q(11)=>q_cache_arr_16_11, q(10)=>q_cache_arr_16_10, q(9)=>
      q_cache_arr_16_9, q(8)=>q_cache_arr_16_8, q(7)=>q_cache_arr_16_7, q(6)
      =>q_cache_arr_16_6, q(5)=>q_cache_arr_16_5, q(4)=>q_cache_arr_16_4, 
      q(3)=>q_cache_arr_16_3, q(2)=>q_cache_arr_16_2, q(1)=>q_cache_arr_16_1, 
      q(0)=>q_cache_arr_16_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1113, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_17_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_17_31, d(30)=>d_cache_arr_17_30, d(29)=>d_cache_arr_17_29, 
      d(28)=>d_cache_arr_17_28, d(27)=>d_cache_arr_17_27, d(26)=>
      d_cache_arr_17_26, d(25)=>d_cache_arr_17_25, d(24)=>d_cache_arr_17_24, 
      d(23)=>d_cache_arr_17_23, d(22)=>d_cache_arr_17_22, d(21)=>
      d_cache_arr_17_21, d(20)=>d_cache_arr_17_20, d(19)=>d_cache_arr_17_19, 
      d(18)=>d_cache_arr_17_18, d(17)=>d_cache_arr_17_17, d(16)=>
      d_cache_arr_17_16, d(15)=>d_cache_arr_17_15, d(14)=>d_cache_arr_17_14, 
      d(13)=>d_cache_arr_17_13, d(12)=>d_cache_arr_17_12, d(11)=>
      d_cache_arr_17_11, d(10)=>d_cache_arr_17_10, d(9)=>d_cache_arr_17_9, 
      d(8)=>d_cache_arr_17_8, d(7)=>d_cache_arr_17_7, d(6)=>d_cache_arr_17_6, 
      d(5)=>d_cache_arr_17_5, d(4)=>d_cache_arr_17_4, d(3)=>d_cache_arr_17_3, 
      d(2)=>d_cache_arr_17_2, d(1)=>d_cache_arr_17_1, d(0)=>d_cache_arr_17_0, 
      q(31)=>q_cache_arr_17_31, q(30)=>q_cache_arr_17_30, q(29)=>
      q_cache_arr_17_29, q(28)=>q_cache_arr_17_28, q(27)=>q_cache_arr_17_27, 
      q(26)=>q_cache_arr_17_26, q(25)=>q_cache_arr_17_25, q(24)=>
      q_cache_arr_17_24, q(23)=>q_cache_arr_17_23, q(22)=>q_cache_arr_17_22, 
      q(21)=>q_cache_arr_17_21, q(20)=>q_cache_arr_17_20, q(19)=>
      q_cache_arr_17_19, q(18)=>q_cache_arr_17_18, q(17)=>q_cache_arr_17_17, 
      q(16)=>q_cache_arr_17_16, q(15)=>q_cache_arr_17_15, q(14)=>
      q_cache_arr_17_14, q(13)=>q_cache_arr_17_13, q(12)=>q_cache_arr_17_12, 
      q(11)=>q_cache_arr_17_11, q(10)=>q_cache_arr_17_10, q(9)=>
      q_cache_arr_17_9, q(8)=>q_cache_arr_17_8, q(7)=>q_cache_arr_17_7, q(6)
      =>q_cache_arr_17_6, q(5)=>q_cache_arr_17_5, q(4)=>q_cache_arr_17_4, 
      q(3)=>q_cache_arr_17_3, q(2)=>q_cache_arr_17_2, q(1)=>q_cache_arr_17_1, 
      q(0)=>q_cache_arr_17_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1113, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_18_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_18_31, d(30)=>d_cache_arr_18_30, d(29)=>d_cache_arr_18_29, 
      d(28)=>d_cache_arr_18_28, d(27)=>d_cache_arr_18_27, d(26)=>
      d_cache_arr_18_26, d(25)=>d_cache_arr_18_25, d(24)=>d_cache_arr_18_24, 
      d(23)=>d_cache_arr_18_23, d(22)=>d_cache_arr_18_22, d(21)=>
      d_cache_arr_18_21, d(20)=>d_cache_arr_18_20, d(19)=>d_cache_arr_18_19, 
      d(18)=>d_cache_arr_18_18, d(17)=>d_cache_arr_18_17, d(16)=>
      d_cache_arr_18_16, d(15)=>d_cache_arr_18_15, d(14)=>d_cache_arr_18_14, 
      d(13)=>d_cache_arr_18_13, d(12)=>d_cache_arr_18_12, d(11)=>
      d_cache_arr_18_11, d(10)=>d_cache_arr_18_10, d(9)=>d_cache_arr_18_9, 
      d(8)=>d_cache_arr_18_8, d(7)=>d_cache_arr_18_7, d(6)=>d_cache_arr_18_6, 
      d(5)=>d_cache_arr_18_5, d(4)=>d_cache_arr_18_4, d(3)=>d_cache_arr_18_3, 
      d(2)=>d_cache_arr_18_2, d(1)=>d_cache_arr_18_1, d(0)=>d_cache_arr_18_0, 
      q(31)=>q_cache_arr_18_31, q(30)=>q_cache_arr_18_30, q(29)=>
      q_cache_arr_18_29, q(28)=>q_cache_arr_18_28, q(27)=>q_cache_arr_18_27, 
      q(26)=>q_cache_arr_18_26, q(25)=>q_cache_arr_18_25, q(24)=>
      q_cache_arr_18_24, q(23)=>q_cache_arr_18_23, q(22)=>q_cache_arr_18_22, 
      q(21)=>q_cache_arr_18_21, q(20)=>q_cache_arr_18_20, q(19)=>
      q_cache_arr_18_19, q(18)=>q_cache_arr_18_18, q(17)=>q_cache_arr_18_17, 
      q(16)=>q_cache_arr_18_16, q(15)=>q_cache_arr_18_15, q(14)=>
      q_cache_arr_18_14, q(13)=>q_cache_arr_18_13, q(12)=>q_cache_arr_18_12, 
      q(11)=>q_cache_arr_18_11, q(10)=>q_cache_arr_18_10, q(9)=>
      q_cache_arr_18_9, q(8)=>q_cache_arr_18_8, q(7)=>q_cache_arr_18_7, q(6)
      =>q_cache_arr_18_6, q(5)=>q_cache_arr_18_5, q(4)=>q_cache_arr_18_4, 
      q(3)=>q_cache_arr_18_3, q(2)=>q_cache_arr_18_2, q(1)=>q_cache_arr_18_1, 
      q(0)=>q_cache_arr_18_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1113, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_19_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_19_31, d(30)=>d_cache_arr_19_30, d(29)=>d_cache_arr_19_29, 
      d(28)=>d_cache_arr_19_28, d(27)=>d_cache_arr_19_27, d(26)=>
      d_cache_arr_19_26, d(25)=>d_cache_arr_19_25, d(24)=>d_cache_arr_19_24, 
      d(23)=>d_cache_arr_19_23, d(22)=>d_cache_arr_19_22, d(21)=>
      d_cache_arr_19_21, d(20)=>d_cache_arr_19_20, d(19)=>d_cache_arr_19_19, 
      d(18)=>d_cache_arr_19_18, d(17)=>d_cache_arr_19_17, d(16)=>
      d_cache_arr_19_16, d(15)=>d_cache_arr_19_15, d(14)=>d_cache_arr_19_14, 
      d(13)=>d_cache_arr_19_13, d(12)=>d_cache_arr_19_12, d(11)=>
      d_cache_arr_19_11, d(10)=>d_cache_arr_19_10, d(9)=>d_cache_arr_19_9, 
      d(8)=>d_cache_arr_19_8, d(7)=>d_cache_arr_19_7, d(6)=>d_cache_arr_19_6, 
      d(5)=>d_cache_arr_19_5, d(4)=>d_cache_arr_19_4, d(3)=>d_cache_arr_19_3, 
      d(2)=>d_cache_arr_19_2, d(1)=>d_cache_arr_19_1, d(0)=>d_cache_arr_19_0, 
      q(31)=>q_cache_arr_19_31, q(30)=>q_cache_arr_19_30, q(29)=>
      q_cache_arr_19_29, q(28)=>q_cache_arr_19_28, q(27)=>q_cache_arr_19_27, 
      q(26)=>q_cache_arr_19_26, q(25)=>q_cache_arr_19_25, q(24)=>
      q_cache_arr_19_24, q(23)=>q_cache_arr_19_23, q(22)=>q_cache_arr_19_22, 
      q(21)=>q_cache_arr_19_21, q(20)=>q_cache_arr_19_20, q(19)=>
      q_cache_arr_19_19, q(18)=>q_cache_arr_19_18, q(17)=>q_cache_arr_19_17, 
      q(16)=>q_cache_arr_19_16, q(15)=>q_cache_arr_19_15, q(14)=>
      q_cache_arr_19_14, q(13)=>q_cache_arr_19_13, q(12)=>q_cache_arr_19_12, 
      q(11)=>q_cache_arr_19_11, q(10)=>q_cache_arr_19_10, q(9)=>
      q_cache_arr_19_9, q(8)=>q_cache_arr_19_8, q(7)=>q_cache_arr_19_7, q(6)
      =>q_cache_arr_19_6, q(5)=>q_cache_arr_19_5, q(4)=>q_cache_arr_19_4, 
      q(3)=>q_cache_arr_19_3, q(2)=>q_cache_arr_19_2, q(1)=>q_cache_arr_19_1, 
      q(0)=>q_cache_arr_19_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1113, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_20_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_20_31, d(30)=>d_cache_arr_20_30, d(29)=>d_cache_arr_20_29, 
      d(28)=>d_cache_arr_20_28, d(27)=>d_cache_arr_20_27, d(26)=>
      d_cache_arr_20_26, d(25)=>d_cache_arr_20_25, d(24)=>d_cache_arr_20_24, 
      d(23)=>d_cache_arr_20_23, d(22)=>d_cache_arr_20_22, d(21)=>
      d_cache_arr_20_21, d(20)=>d_cache_arr_20_20, d(19)=>d_cache_arr_20_19, 
      d(18)=>d_cache_arr_20_18, d(17)=>d_cache_arr_20_17, d(16)=>
      d_cache_arr_20_16, d(15)=>d_cache_arr_20_15, d(14)=>d_cache_arr_20_14, 
      d(13)=>d_cache_arr_20_13, d(12)=>d_cache_arr_20_12, d(11)=>
      d_cache_arr_20_11, d(10)=>d_cache_arr_20_10, d(9)=>d_cache_arr_20_9, 
      d(8)=>d_cache_arr_20_8, d(7)=>d_cache_arr_20_7, d(6)=>d_cache_arr_20_6, 
      d(5)=>d_cache_arr_20_5, d(4)=>d_cache_arr_20_4, d(3)=>d_cache_arr_20_3, 
      d(2)=>d_cache_arr_20_2, d(1)=>d_cache_arr_20_1, d(0)=>d_cache_arr_20_0, 
      q(31)=>q_cache_arr_20_31, q(30)=>q_cache_arr_20_30, q(29)=>
      q_cache_arr_20_29, q(28)=>q_cache_arr_20_28, q(27)=>q_cache_arr_20_27, 
      q(26)=>q_cache_arr_20_26, q(25)=>q_cache_arr_20_25, q(24)=>
      q_cache_arr_20_24, q(23)=>q_cache_arr_20_23, q(22)=>q_cache_arr_20_22, 
      q(21)=>q_cache_arr_20_21, q(20)=>q_cache_arr_20_20, q(19)=>
      q_cache_arr_20_19, q(18)=>q_cache_arr_20_18, q(17)=>q_cache_arr_20_17, 
      q(16)=>q_cache_arr_20_16, q(15)=>q_cache_arr_20_15, q(14)=>
      q_cache_arr_20_14, q(13)=>q_cache_arr_20_13, q(12)=>q_cache_arr_20_12, 
      q(11)=>q_cache_arr_20_11, q(10)=>q_cache_arr_20_10, q(9)=>
      q_cache_arr_20_9, q(8)=>q_cache_arr_20_8, q(7)=>q_cache_arr_20_7, q(6)
      =>q_cache_arr_20_6, q(5)=>q_cache_arr_20_5, q(4)=>q_cache_arr_20_4, 
      q(3)=>q_cache_arr_20_3, q(2)=>q_cache_arr_20_2, q(1)=>q_cache_arr_20_1, 
      q(0)=>q_cache_arr_20_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1113, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_21_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_21_31, d(30)=>d_cache_arr_21_30, d(29)=>d_cache_arr_21_29, 
      d(28)=>d_cache_arr_21_28, d(27)=>d_cache_arr_21_27, d(26)=>
      d_cache_arr_21_26, d(25)=>d_cache_arr_21_25, d(24)=>d_cache_arr_21_24, 
      d(23)=>d_cache_arr_21_23, d(22)=>d_cache_arr_21_22, d(21)=>
      d_cache_arr_21_21, d(20)=>d_cache_arr_21_20, d(19)=>d_cache_arr_21_19, 
      d(18)=>d_cache_arr_21_18, d(17)=>d_cache_arr_21_17, d(16)=>
      d_cache_arr_21_16, d(15)=>d_cache_arr_21_15, d(14)=>d_cache_arr_21_14, 
      d(13)=>d_cache_arr_21_13, d(12)=>d_cache_arr_21_12, d(11)=>
      d_cache_arr_21_11, d(10)=>d_cache_arr_21_10, d(9)=>d_cache_arr_21_9, 
      d(8)=>d_cache_arr_21_8, d(7)=>d_cache_arr_21_7, d(6)=>d_cache_arr_21_6, 
      d(5)=>d_cache_arr_21_5, d(4)=>d_cache_arr_21_4, d(3)=>d_cache_arr_21_3, 
      d(2)=>d_cache_arr_21_2, d(1)=>d_cache_arr_21_1, d(0)=>d_cache_arr_21_0, 
      q(31)=>q_cache_arr_21_31, q(30)=>q_cache_arr_21_30, q(29)=>
      q_cache_arr_21_29, q(28)=>q_cache_arr_21_28, q(27)=>q_cache_arr_21_27, 
      q(26)=>q_cache_arr_21_26, q(25)=>q_cache_arr_21_25, q(24)=>
      q_cache_arr_21_24, q(23)=>q_cache_arr_21_23, q(22)=>q_cache_arr_21_22, 
      q(21)=>q_cache_arr_21_21, q(20)=>q_cache_arr_21_20, q(19)=>
      q_cache_arr_21_19, q(18)=>q_cache_arr_21_18, q(17)=>q_cache_arr_21_17, 
      q(16)=>q_cache_arr_21_16, q(15)=>q_cache_arr_21_15, q(14)=>
      q_cache_arr_21_14, q(13)=>q_cache_arr_21_13, q(12)=>q_cache_arr_21_12, 
      q(11)=>q_cache_arr_21_11, q(10)=>q_cache_arr_21_10, q(9)=>
      q_cache_arr_21_9, q(8)=>q_cache_arr_21_8, q(7)=>q_cache_arr_21_7, q(6)
      =>q_cache_arr_21_6, q(5)=>q_cache_arr_21_5, q(4)=>q_cache_arr_21_4, 
      q(3)=>q_cache_arr_21_3, q(2)=>q_cache_arr_21_2, q(1)=>q_cache_arr_21_1, 
      q(0)=>q_cache_arr_21_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1115, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_22_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_22_31, d(30)=>d_cache_arr_22_30, d(29)=>d_cache_arr_22_29, 
      d(28)=>d_cache_arr_22_28, d(27)=>d_cache_arr_22_27, d(26)=>
      d_cache_arr_22_26, d(25)=>d_cache_arr_22_25, d(24)=>d_cache_arr_22_24, 
      d(23)=>d_cache_arr_22_23, d(22)=>d_cache_arr_22_22, d(21)=>
      d_cache_arr_22_21, d(20)=>d_cache_arr_22_20, d(19)=>d_cache_arr_22_19, 
      d(18)=>d_cache_arr_22_18, d(17)=>d_cache_arr_22_17, d(16)=>
      d_cache_arr_22_16, d(15)=>d_cache_arr_22_15, d(14)=>d_cache_arr_22_14, 
      d(13)=>d_cache_arr_22_13, d(12)=>d_cache_arr_22_12, d(11)=>
      d_cache_arr_22_11, d(10)=>d_cache_arr_22_10, d(9)=>d_cache_arr_22_9, 
      d(8)=>d_cache_arr_22_8, d(7)=>d_cache_arr_22_7, d(6)=>d_cache_arr_22_6, 
      d(5)=>d_cache_arr_22_5, d(4)=>d_cache_arr_22_4, d(3)=>d_cache_arr_22_3, 
      d(2)=>d_cache_arr_22_2, d(1)=>d_cache_arr_22_1, d(0)=>d_cache_arr_22_0, 
      q(31)=>q_cache_arr_22_31, q(30)=>q_cache_arr_22_30, q(29)=>
      q_cache_arr_22_29, q(28)=>q_cache_arr_22_28, q(27)=>q_cache_arr_22_27, 
      q(26)=>q_cache_arr_22_26, q(25)=>q_cache_arr_22_25, q(24)=>
      q_cache_arr_22_24, q(23)=>q_cache_arr_22_23, q(22)=>q_cache_arr_22_22, 
      q(21)=>q_cache_arr_22_21, q(20)=>q_cache_arr_22_20, q(19)=>
      q_cache_arr_22_19, q(18)=>q_cache_arr_22_18, q(17)=>q_cache_arr_22_17, 
      q(16)=>q_cache_arr_22_16, q(15)=>q_cache_arr_22_15, q(14)=>
      q_cache_arr_22_14, q(13)=>q_cache_arr_22_13, q(12)=>q_cache_arr_22_12, 
      q(11)=>q_cache_arr_22_11, q(10)=>q_cache_arr_22_10, q(9)=>
      q_cache_arr_22_9, q(8)=>q_cache_arr_22_8, q(7)=>q_cache_arr_22_7, q(6)
      =>q_cache_arr_22_6, q(5)=>q_cache_arr_22_5, q(4)=>q_cache_arr_22_4, 
      q(3)=>q_cache_arr_22_3, q(2)=>q_cache_arr_22_2, q(1)=>q_cache_arr_22_1, 
      q(0)=>q_cache_arr_22_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1115, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_23_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_23_31, d(30)=>d_cache_arr_23_30, d(29)=>d_cache_arr_23_29, 
      d(28)=>d_cache_arr_23_28, d(27)=>d_cache_arr_23_27, d(26)=>
      d_cache_arr_23_26, d(25)=>d_cache_arr_23_25, d(24)=>d_cache_arr_23_24, 
      d(23)=>d_cache_arr_23_23, d(22)=>d_cache_arr_23_22, d(21)=>
      d_cache_arr_23_21, d(20)=>d_cache_arr_23_20, d(19)=>d_cache_arr_23_19, 
      d(18)=>d_cache_arr_23_18, d(17)=>d_cache_arr_23_17, d(16)=>
      d_cache_arr_23_16, d(15)=>d_cache_arr_23_15, d(14)=>d_cache_arr_23_14, 
      d(13)=>d_cache_arr_23_13, d(12)=>d_cache_arr_23_12, d(11)=>
      d_cache_arr_23_11, d(10)=>d_cache_arr_23_10, d(9)=>d_cache_arr_23_9, 
      d(8)=>d_cache_arr_23_8, d(7)=>d_cache_arr_23_7, d(6)=>d_cache_arr_23_6, 
      d(5)=>d_cache_arr_23_5, d(4)=>d_cache_arr_23_4, d(3)=>d_cache_arr_23_3, 
      d(2)=>d_cache_arr_23_2, d(1)=>d_cache_arr_23_1, d(0)=>d_cache_arr_23_0, 
      q(31)=>q_cache_arr_23_31, q(30)=>q_cache_arr_23_30, q(29)=>
      q_cache_arr_23_29, q(28)=>q_cache_arr_23_28, q(27)=>q_cache_arr_23_27, 
      q(26)=>q_cache_arr_23_26, q(25)=>q_cache_arr_23_25, q(24)=>
      q_cache_arr_23_24, q(23)=>q_cache_arr_23_23, q(22)=>q_cache_arr_23_22, 
      q(21)=>q_cache_arr_23_21, q(20)=>q_cache_arr_23_20, q(19)=>
      q_cache_arr_23_19, q(18)=>q_cache_arr_23_18, q(17)=>q_cache_arr_23_17, 
      q(16)=>q_cache_arr_23_16, q(15)=>q_cache_arr_23_15, q(14)=>
      q_cache_arr_23_14, q(13)=>q_cache_arr_23_13, q(12)=>q_cache_arr_23_12, 
      q(11)=>q_cache_arr_23_11, q(10)=>q_cache_arr_23_10, q(9)=>
      q_cache_arr_23_9, q(8)=>q_cache_arr_23_8, q(7)=>q_cache_arr_23_7, q(6)
      =>q_cache_arr_23_6, q(5)=>q_cache_arr_23_5, q(4)=>q_cache_arr_23_4, 
      q(3)=>q_cache_arr_23_3, q(2)=>q_cache_arr_23_2, q(1)=>q_cache_arr_23_1, 
      q(0)=>q_cache_arr_23_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1115, reset=>
      filter_reset);
   gen_comp_cache_gen_regs_24_gen_regi : Reg_32 port map ( d(31)=>
      d_cache_arr_24_31, d(30)=>d_cache_arr_24_30, d(29)=>d_cache_arr_24_29, 
      d(28)=>d_cache_arr_24_28, d(27)=>d_cache_arr_24_27, d(26)=>
      d_cache_arr_24_26, d(25)=>d_cache_arr_24_25, d(24)=>d_cache_arr_24_24, 
      d(23)=>d_cache_arr_24_23, d(22)=>d_cache_arr_24_22, d(21)=>
      d_cache_arr_24_21, d(20)=>d_cache_arr_24_20, d(19)=>d_cache_arr_24_19, 
      d(18)=>d_cache_arr_24_18, d(17)=>d_cache_arr_24_17, d(16)=>
      d_cache_arr_24_16, d(15)=>d_cache_arr_24_15, d(14)=>d_cache_arr_24_14, 
      d(13)=>d_cache_arr_24_13, d(12)=>d_cache_arr_24_12, d(11)=>
      d_cache_arr_24_11, d(10)=>d_cache_arr_24_10, d(9)=>d_cache_arr_24_9, 
      d(8)=>d_cache_arr_24_8, d(7)=>d_cache_arr_24_7, d(6)=>d_cache_arr_24_6, 
      d(5)=>d_cache_arr_24_5, d(4)=>d_cache_arr_24_4, d(3)=>d_cache_arr_24_3, 
      d(2)=>d_cache_arr_24_2, d(1)=>d_cache_arr_24_1, d(0)=>d_cache_arr_24_0, 
      q(31)=>q_cache_arr_24_31, q(30)=>q_cache_arr_24_30, q(29)=>
      q_cache_arr_24_29, q(28)=>q_cache_arr_24_28, q(27)=>q_cache_arr_24_27, 
      q(26)=>q_cache_arr_24_26, q(25)=>q_cache_arr_24_25, q(24)=>
      q_cache_arr_24_24, q(23)=>q_cache_arr_24_23, q(22)=>q_cache_arr_24_22, 
      q(21)=>q_cache_arr_24_21, q(20)=>q_cache_arr_24_20, q(19)=>
      q_cache_arr_24_19, q(18)=>q_cache_arr_24_18, q(17)=>q_cache_arr_24_17, 
      q(16)=>q_cache_arr_24_16, q(15)=>q_cache_arr_24_15, q(14)=>
      q_cache_arr_24_14, q(13)=>q_cache_arr_24_13, q(12)=>q_cache_arr_24_12, 
      q(11)=>q_cache_arr_24_11, q(10)=>q_cache_arr_24_10, q(9)=>
      q_cache_arr_24_9, q(8)=>q_cache_arr_24_8, q(7)=>q_cache_arr_24_7, q(6)
      =>q_cache_arr_24_6, q(5)=>q_cache_arr_24_5, q(4)=>q_cache_arr_24_4, 
      q(3)=>q_cache_arr_24_3, q(2)=>q_cache_arr_24_2, q(1)=>q_cache_arr_24_1, 
      q(0)=>q_cache_arr_24_0, rst_data(31)=>buffer_ready_EXMPLR, 
      rst_data(30)=>buffer_ready_EXMPLR, rst_data(29)=>buffer_ready_EXMPLR, 
      rst_data(28)=>buffer_ready_EXMPLR, rst_data(27)=>buffer_ready_EXMPLR, 
      rst_data(26)=>buffer_ready_EXMPLR, rst_data(25)=>buffer_ready_EXMPLR, 
      rst_data(24)=>buffer_ready_EXMPLR, rst_data(23)=>buffer_ready_EXMPLR, 
      rst_data(22)=>buffer_ready_EXMPLR, rst_data(21)=>buffer_ready_EXMPLR, 
      rst_data(20)=>buffer_ready_EXMPLR, rst_data(19)=>buffer_ready_EXMPLR, 
      rst_data(18)=>buffer_ready_EXMPLR, rst_data(17)=>buffer_ready_EXMPLR, 
      rst_data(16)=>buffer_ready_EXMPLR, rst_data(15)=>buffer_ready_EXMPLR, 
      rst_data(14)=>buffer_ready_EXMPLR, rst_data(13)=>buffer_ready_EXMPLR, 
      rst_data(12)=>buffer_ready_EXMPLR, rst_data(11)=>buffer_ready_EXMPLR, 
      rst_data(10)=>buffer_ready_EXMPLR, rst_data(9)=>buffer_ready_EXMPLR, 
      rst_data(8)=>buffer_ready_EXMPLR, rst_data(7)=>buffer_ready_EXMPLR, 
      rst_data(6)=>buffer_ready_EXMPLR, rst_data(5)=>buffer_ready_EXMPLR, 
      rst_data(4)=>buffer_ready_EXMPLR, rst_data(3)=>buffer_ready_EXMPLR, 
      rst_data(2)=>buffer_ready_EXMPLR, rst_data(1)=>buffer_ready_EXMPLR, 
      rst_data(0)=>buffer_ready_EXMPLR, clk=>clk, load=>nx1115, reset=>
      filter_reset);
   ix48 : fake_gnd port map ( Y=>buffer_ready_EXMPLR);
   reg_compute_relu_q : dffs_ni port map ( Q=>compute_relu_q, QB=>OPEN, D=>
      nx541, CLK=>nx1137, S=>filter_reset);
   ix876 : nand02 port map ( Y=>nx875, A0=>start, A1=>ready_EXMPLR);
   reg_ready_q : dffs_ni port map ( Q=>ready_EXMPLR, QB=>OPEN, D=>nx10, CLK
      =>nx1183, S=>filter_reset);
   ix11 : inv01 port map ( Y=>nx10, A=>nx879);
   ix880 : oai21 port map ( Y=>nx879, A0=>ready_EXMPLR, A1=>ready_tmp, B0=>
      nx1151);
   reg_operation_q : dffr port map ( Q=>operation_q, QB=>OPEN, D=>nx531, CLK
      =>nx1137, R=>filter_reset);
   reg_filter_size_q : dffr port map ( Q=>filter_size_q, QB=>OPEN, D=>nx521, 
      CLK=>nx1137, R=>filter_reset);
   reg_output2_init_q_0 : dffr port map ( Q=>output2_init_q_0, QB=>OPEN, D=>
      nx361, CLK=>nx1137, R=>filter_reset);
   reg_output2_init_q_1 : dffr port map ( Q=>output2_init_q_1, QB=>OPEN, D=>
      nx371, CLK=>nx1137, R=>filter_reset);
   reg_output2_init_q_2 : dffr port map ( Q=>output2_init_q_2, QB=>OPEN, D=>
      nx381, CLK=>nx1137, R=>filter_reset);
   reg_output2_init_q_3 : dffr port map ( Q=>output2_init_q_3, QB=>OPEN, D=>
      nx391, CLK=>nx1137, R=>filter_reset);
   reg_output2_init_q_4 : dffr port map ( Q=>output2_init_q_4, QB=>OPEN, D=>
      nx401, CLK=>nx1139, R=>filter_reset);
   reg_output2_init_q_5 : dffr port map ( Q=>output2_init_q_5, QB=>OPEN, D=>
      nx411, CLK=>nx1139, R=>filter_reset);
   reg_output2_init_q_6 : dffr port map ( Q=>output2_init_q_6, QB=>OPEN, D=>
      nx421, CLK=>nx1139, R=>filter_reset);
   reg_output2_init_q_7 : dffr port map ( Q=>output2_init_q_7, QB=>OPEN, D=>
      nx431, CLK=>nx1139, R=>filter_reset);
   reg_output2_init_q_8 : dffr port map ( Q=>output2_init_q_8, QB=>OPEN, D=>
      nx441, CLK=>nx1139, R=>filter_reset);
   reg_output2_init_q_9 : dffr port map ( Q=>output2_init_q_9, QB=>OPEN, D=>
      nx451, CLK=>nx1139, R=>filter_reset);
   reg_output2_init_q_10 : dffr port map ( Q=>output2_init_q_10, QB=>OPEN, D
      =>nx461, CLK=>nx1139, R=>filter_reset);
   reg_output2_init_q_11 : dffr port map ( Q=>output2_init_q_11, QB=>OPEN, D
      =>nx471, CLK=>nx1141, R=>filter_reset);
   reg_output2_init_q_12 : dffr port map ( Q=>output2_init_q_12, QB=>OPEN, D
      =>nx481, CLK=>nx1141, R=>filter_reset);
   reg_output2_init_q_13 : dffr port map ( Q=>output2_init_q_13, QB=>OPEN, D
      =>nx491, CLK=>nx1141, R=>filter_reset);
   reg_output2_init_q_14 : dffr port map ( Q=>output2_init_q_14, QB=>OPEN, D
      =>nx501, CLK=>nx1141, R=>filter_reset);
   reg_output2_init_q_15 : dffr port map ( Q=>output2_init_q_15, QB=>OPEN, D
      =>nx511, CLK=>nx1141, R=>filter_reset);
   reg_output1_init_q_0 : dffr port map ( Q=>output1_init_q_0, QB=>OPEN, D=>
      nx201, CLK=>nx1141, R=>filter_reset);
   reg_output1_init_q_1 : dffr port map ( Q=>output1_init_q_1, QB=>OPEN, D=>
      nx211, CLK=>nx1141, R=>filter_reset);
   reg_output1_init_q_2 : dffr port map ( Q=>output1_init_q_2, QB=>OPEN, D=>
      nx221, CLK=>nx1143, R=>filter_reset);
   reg_output1_init_q_3 : dffr port map ( Q=>output1_init_q_3, QB=>OPEN, D=>
      nx231, CLK=>nx1143, R=>filter_reset);
   reg_output1_init_q_4 : dffr port map ( Q=>output1_init_q_4, QB=>OPEN, D=>
      nx241, CLK=>nx1143, R=>filter_reset);
   reg_output1_init_q_5 : dffr port map ( Q=>output1_init_q_5, QB=>OPEN, D=>
      nx251, CLK=>nx1143, R=>filter_reset);
   reg_output1_init_q_6 : dffr port map ( Q=>output1_init_q_6, QB=>OPEN, D=>
      nx261, CLK=>nx1143, R=>filter_reset);
   reg_output1_init_q_7 : dffr port map ( Q=>output1_init_q_7, QB=>OPEN, D=>
      nx271, CLK=>nx1143, R=>filter_reset);
   reg_output1_init_q_8 : dffr port map ( Q=>output1_init_q_8, QB=>OPEN, D=>
      nx281, CLK=>nx1143, R=>filter_reset);
   reg_output1_init_q_9 : dffr port map ( Q=>output1_init_q_9, QB=>OPEN, D=>
      nx291, CLK=>nx1145, R=>filter_reset);
   reg_output1_init_q_10 : dffr port map ( Q=>output1_init_q_10, QB=>OPEN, D
      =>nx301, CLK=>nx1145, R=>filter_reset);
   reg_output1_init_q_11 : dffr port map ( Q=>output1_init_q_11, QB=>OPEN, D
      =>nx311, CLK=>nx1145, R=>filter_reset);
   reg_output1_init_q_12 : dffr port map ( Q=>output1_init_q_12, QB=>OPEN, D
      =>nx321, CLK=>nx1145, R=>filter_reset);
   reg_output1_init_q_13 : dffr port map ( Q=>output1_init_q_13, QB=>OPEN, D
      =>nx331, CLK=>nx1145, R=>filter_reset);
   reg_output1_init_q_14 : dffr port map ( Q=>output1_init_q_14, QB=>OPEN, D
      =>nx341, CLK=>nx1145, R=>filter_reset);
   reg_output1_init_q_15 : dffr port map ( Q=>output1_init_q_15, QB=>OPEN, D
      =>nx351, CLK=>nx1145, R=>filter_reset);
   reg_comp_pipe_en : dffr port map ( Q=>comp_pipe_en, QB=>OPEN, D=>NOT_nx4, 
      CLK=>nx1147, R=>filter_reset);
   ix987 : nand02 port map ( Y=>NOT_nx4, A0=>ready_tmp, A1=>nx1161);
   reg_comp_pipe_rst : dffs_ni port map ( Q=>comp_pipe_rst, QB=>OPEN, D=>nx4, 
      CLK=>nx1147, S=>filter_reset);
   ix309 : and02 port map ( Y=>filter_load_tmp, A0=>filter_load, A1=>
      buffer_ready_dup0);
   reg_buffer_ready_q : dffs_ni port map ( Q=>buffer_ready_dup0, QB=>OPEN, D
      =>nx302, CLK=>nx1147, S=>filter_reset);
   ix303 : inv01 port map ( Y=>nx302, A=>nx996);
   ix997 : oai21 port map ( Y=>nx996, A0=>buffer_ready_dup0, A1=>
      buffer_ready_tmp, B0=>nx1161);
   ix311 : and02 port map ( Y=>img_load_tmp, A0=>img_load, A1=>
      buffer_ready_dup0);
   reg_output2_q_0 : dffr port map ( Q=>output2_0_EXMPLR, QB=>OPEN, D=>nx711, 
      CLK=>clk, R=>filter_reset);
   reg_output2_q_1 : dffr port map ( Q=>output2_1_EXMPLR, QB=>OPEN, D=>nx721, 
      CLK=>clk, R=>filter_reset);
   reg_output2_q_2 : dffr port map ( Q=>output2_2_EXMPLR, QB=>OPEN, D=>nx731, 
      CLK=>clk, R=>filter_reset);
   reg_output2_q_3 : dffr port map ( Q=>output2_3_EXMPLR, QB=>OPEN, D=>nx741, 
      CLK=>clk, R=>filter_reset);
   reg_output2_q_4 : dffr port map ( Q=>output2_4_EXMPLR, QB=>OPEN, D=>nx751, 
      CLK=>clk, R=>filter_reset);
   reg_output2_q_5 : dffr port map ( Q=>output2_5_EXMPLR, QB=>OPEN, D=>nx761, 
      CLK=>clk, R=>filter_reset);
   reg_output2_q_6 : dffr port map ( Q=>output2_6_EXMPLR, QB=>OPEN, D=>nx771, 
      CLK=>clk, R=>filter_reset);
   reg_output2_q_7 : dffr port map ( Q=>output2_7_EXMPLR, QB=>OPEN, D=>nx781, 
      CLK=>clk, R=>filter_reset);
   reg_output2_q_8 : dffr port map ( Q=>output2_8_EXMPLR, QB=>OPEN, D=>nx791, 
      CLK=>clk, R=>filter_reset);
   reg_output2_q_9 : dffr port map ( Q=>output2_9_EXMPLR, QB=>OPEN, D=>nx801, 
      CLK=>clk, R=>filter_reset);
   reg_output2_q_10 : dffr port map ( Q=>output2_10_EXMPLR, QB=>OPEN, D=>
      nx811, CLK=>clk, R=>filter_reset);
   reg_output2_q_11 : dffr port map ( Q=>output2_11_EXMPLR, QB=>OPEN, D=>
      nx821, CLK=>clk, R=>filter_reset);
   reg_output2_q_12 : dffr port map ( Q=>output2_12_EXMPLR, QB=>OPEN, D=>
      nx831, CLK=>clk, R=>filter_reset);
   reg_output2_q_13 : dffr port map ( Q=>output2_13_EXMPLR, QB=>OPEN, D=>
      nx841, CLK=>clk, R=>filter_reset);
   reg_output2_q_14 : dffr port map ( Q=>output2_14_EXMPLR, QB=>OPEN, D=>
      nx851, CLK=>clk, R=>filter_reset);
   reg_output2_q_15 : dffr port map ( Q=>output2_15_EXMPLR, QB=>OPEN, D=>
      nx861, CLK=>clk, R=>filter_reset);
   reg_output1_q_0 : dffr port map ( Q=>output1_0_EXMPLR, QB=>OPEN, D=>nx551, 
      CLK=>clk, R=>filter_reset);
   reg_output1_q_1 : dffr port map ( Q=>output1_1_EXMPLR, QB=>OPEN, D=>nx561, 
      CLK=>clk, R=>filter_reset);
   reg_output1_q_2 : dffr port map ( Q=>output1_2_EXMPLR, QB=>OPEN, D=>nx571, 
      CLK=>clk, R=>filter_reset);
   reg_output1_q_3 : dffr port map ( Q=>output1_3_EXMPLR, QB=>OPEN, D=>nx581, 
      CLK=>clk, R=>filter_reset);
   reg_output1_q_4 : dffr port map ( Q=>output1_4_EXMPLR, QB=>OPEN, D=>nx591, 
      CLK=>clk, R=>filter_reset);
   reg_output1_q_5 : dffr port map ( Q=>output1_5_EXMPLR, QB=>OPEN, D=>nx601, 
      CLK=>clk, R=>filter_reset);
   reg_output1_q_6 : dffr port map ( Q=>output1_6_EXMPLR, QB=>OPEN, D=>nx611, 
      CLK=>clk, R=>filter_reset);
   reg_output1_q_7 : dffr port map ( Q=>output1_7_EXMPLR, QB=>OPEN, D=>nx621, 
      CLK=>clk, R=>filter_reset);
   reg_output1_q_8 : dffr port map ( Q=>output1_8_EXMPLR, QB=>OPEN, D=>nx631, 
      CLK=>clk, R=>filter_reset);
   reg_output1_q_9 : dffr port map ( Q=>output1_9_EXMPLR, QB=>OPEN, D=>nx641, 
      CLK=>clk, R=>filter_reset);
   reg_output1_q_10 : dffr port map ( Q=>output1_10_EXMPLR, QB=>OPEN, D=>
      nx651, CLK=>clk, R=>filter_reset);
   reg_output1_q_11 : dffr port map ( Q=>output1_11_EXMPLR, QB=>OPEN, D=>
      nx661, CLK=>clk, R=>filter_reset);
   reg_output1_q_12 : dffr port map ( Q=>output1_12_EXMPLR, QB=>OPEN, D=>
      nx671, CLK=>clk, R=>filter_reset);
   reg_output1_q_13 : dffr port map ( Q=>output1_13_EXMPLR, QB=>OPEN, D=>
      nx681, CLK=>clk, R=>filter_reset);
   reg_output1_q_14 : dffr port map ( Q=>output1_14_EXMPLR, QB=>OPEN, D=>
      nx691, CLK=>clk, R=>filter_reset);
   reg_output1_q_15 : dffr port map ( Q=>output1_15_EXMPLR, QB=>OPEN, D=>
      nx701, CLK=>clk, R=>filter_reset);
   ix5 : inv01 port map ( Y=>nx4, A=>NOT_nx4);
   ix1102 : buf02 port map ( Y=>nx1103, A=>img_data_1_15);
   ix1104 : buf02 port map ( Y=>nx1105, A=>img_data_2_15);
   ix1106 : buf02 port map ( Y=>nx1107, A=>img_data_6_15);
   ix1108 : inv01 port map ( Y=>nx1109, A=>nx1131);
   ix1110 : inv01 port map ( Y=>nx1111, A=>nx1131);
   ix1112 : inv01 port map ( Y=>nx1113, A=>nx1131);
   ix1114 : inv01 port map ( Y=>nx1115, A=>nx1133);
   ix1116 : inv01 port map ( Y=>nx1117, A=>filter_size_q);
   ix1118 : inv01 port map ( Y=>nx1119, A=>nx1117);
   ix1120 : inv01 port map ( Y=>nx1121, A=>nx1117);
   ix1130 : inv02 port map ( Y=>nx1131, A=>nx1167);
   ix1132 : inv02 port map ( Y=>nx1133, A=>nx1167);
   ix1136 : inv02 port map ( Y=>nx1137, A=>clk);
   ix1138 : inv02 port map ( Y=>nx1139, A=>clk);
   ix1140 : inv02 port map ( Y=>nx1141, A=>clk);
   ix1142 : inv02 port map ( Y=>nx1143, A=>clk);
   ix1144 : inv02 port map ( Y=>nx1145, A=>clk);
   ix1146 : inv02 port map ( Y=>nx1147, A=>clk);
   ix1150 : inv02 port map ( Y=>nx1151, A=>nx1185);
   ix1160 : inv02 port map ( Y=>nx1161, A=>nx1185);
   ix542 : mux21_ni port map ( Y=>nx541, A0=>compute_relu_q, A1=>
      compute_relu, S0=>nx1185);
   ix532 : mux21_ni port map ( Y=>nx531, A0=>operation_q, A1=>operation, S0
      =>nx1185);
   ix522 : mux21_ni port map ( Y=>nx521, A0=>nx1121, A1=>filter_size, S0=>
      nx1185);
   ix362 : mux21_ni port map ( Y=>nx361, A0=>output2_init_q_0, A1=>
      output2_init(0), S0=>nx1185);
   ix372 : mux21_ni port map ( Y=>nx371, A0=>output2_init_q_1, A1=>
      output2_init(1), S0=>nx1185);
   ix382 : mux21_ni port map ( Y=>nx381, A0=>output2_init_q_2, A1=>
      output2_init(2), S0=>nx1187);
   ix392 : mux21_ni port map ( Y=>nx391, A0=>output2_init_q_3, A1=>
      output2_init(3), S0=>nx1187);
   ix402 : mux21_ni port map ( Y=>nx401, A0=>output2_init_q_4, A1=>
      output2_init(4), S0=>nx1187);
   ix412 : mux21_ni port map ( Y=>nx411, A0=>output2_init_q_5, A1=>
      output2_init(5), S0=>nx1187);
   ix422 : mux21_ni port map ( Y=>nx421, A0=>output2_init_q_6, A1=>
      output2_init(6), S0=>nx1187);
   ix432 : mux21_ni port map ( Y=>nx431, A0=>output2_init_q_7, A1=>
      output2_init(7), S0=>nx1187);
   ix442 : mux21_ni port map ( Y=>nx441, A0=>output2_init_q_8, A1=>
      output2_init(8), S0=>nx1187);
   ix452 : mux21_ni port map ( Y=>nx451, A0=>output2_init_q_9, A1=>
      output2_init(9), S0=>nx1189);
   ix462 : mux21_ni port map ( Y=>nx461, A0=>output2_init_q_10, A1=>
      output2_init(10), S0=>nx1189);
   ix472 : mux21_ni port map ( Y=>nx471, A0=>output2_init_q_11, A1=>
      output2_init(11), S0=>nx1189);
   ix482 : mux21_ni port map ( Y=>nx481, A0=>output2_init_q_12, A1=>
      output2_init(12), S0=>nx1189);
   ix492 : mux21_ni port map ( Y=>nx491, A0=>output2_init_q_13, A1=>
      output2_init(13), S0=>nx1189);
   ix502 : mux21_ni port map ( Y=>nx501, A0=>output2_init_q_14, A1=>
      output2_init(14), S0=>nx1189);
   ix512 : mux21_ni port map ( Y=>nx511, A0=>output2_init_q_15, A1=>
      output2_init(15), S0=>nx1189);
   ix202 : mux21_ni port map ( Y=>nx201, A0=>output1_init_q_0, A1=>
      output1_init(0), S0=>nx1191);
   ix212 : mux21_ni port map ( Y=>nx211, A0=>output1_init_q_1, A1=>
      output1_init(1), S0=>nx1191);
   ix222 : mux21_ni port map ( Y=>nx221, A0=>output1_init_q_2, A1=>
      output1_init(2), S0=>nx1191);
   ix232 : mux21_ni port map ( Y=>nx231, A0=>output1_init_q_3, A1=>
      output1_init(3), S0=>nx1191);
   ix242 : mux21_ni port map ( Y=>nx241, A0=>output1_init_q_4, A1=>
      output1_init(4), S0=>nx1191);
   ix252 : mux21_ni port map ( Y=>nx251, A0=>output1_init_q_5, A1=>
      output1_init(5), S0=>nx1191);
   ix262 : mux21_ni port map ( Y=>nx261, A0=>output1_init_q_6, A1=>
      output1_init(6), S0=>nx1191);
   ix272 : mux21_ni port map ( Y=>nx271, A0=>output1_init_q_7, A1=>
      output1_init(7), S0=>nx1193);
   ix282 : mux21_ni port map ( Y=>nx281, A0=>output1_init_q_8, A1=>
      output1_init(8), S0=>nx1193);
   ix292 : mux21_ni port map ( Y=>nx291, A0=>output1_init_q_9, A1=>
      output1_init(9), S0=>nx1193);
   ix302 : mux21_ni port map ( Y=>nx301, A0=>output1_init_q_10, A1=>
      output1_init(10), S0=>nx1193);
   ix312 : mux21_ni port map ( Y=>nx311, A0=>output1_init_q_11, A1=>
      output1_init(11), S0=>nx1193);
   ix322 : mux21_ni port map ( Y=>nx321, A0=>output1_init_q_12, A1=>
      output1_init(12), S0=>nx1193);
   ix332 : mux21_ni port map ( Y=>nx331, A0=>output1_init_q_13, A1=>
      output1_init(13), S0=>nx1193);
   ix342 : mux21_ni port map ( Y=>nx341, A0=>output1_init_q_14, A1=>
      output1_init(14), S0=>nx1195);
   ix352 : mux21_ni port map ( Y=>nx351, A0=>output1_init_q_15, A1=>
      output1_init(15), S0=>nx1195);
   ix712 : mux21_ni port map ( Y=>nx711, A0=>q_cache_arr_1_0, A1=>
      output2_0_EXMPLR, S0=>nx1167);
   ix722 : mux21_ni port map ( Y=>nx721, A0=>q_cache_arr_1_1, A1=>
      output2_1_EXMPLR, S0=>nx1167);
   ix732 : mux21_ni port map ( Y=>nx731, A0=>q_cache_arr_1_2, A1=>
      output2_2_EXMPLR, S0=>nx1167);
   ix742 : mux21_ni port map ( Y=>nx741, A0=>q_cache_arr_1_3, A1=>
      output2_3_EXMPLR, S0=>nx1167);
   ix752 : mux21_ni port map ( Y=>nx751, A0=>q_cache_arr_1_4, A1=>
      output2_4_EXMPLR, S0=>nx1167);
   ix762 : mux21_ni port map ( Y=>nx761, A0=>q_cache_arr_1_5, A1=>
      output2_5_EXMPLR, S0=>nx1169);
   ix772 : mux21_ni port map ( Y=>nx771, A0=>q_cache_arr_1_6, A1=>
      output2_6_EXMPLR, S0=>nx1169);
   ix782 : mux21_ni port map ( Y=>nx781, A0=>q_cache_arr_1_7, A1=>
      output2_7_EXMPLR, S0=>nx1169);
   ix792 : mux21_ni port map ( Y=>nx791, A0=>q_cache_arr_1_8, A1=>
      output2_8_EXMPLR, S0=>nx1169);
   ix802 : mux21_ni port map ( Y=>nx801, A0=>q_cache_arr_1_9, A1=>
      output2_9_EXMPLR, S0=>nx1169);
   ix812 : mux21_ni port map ( Y=>nx811, A0=>q_cache_arr_1_10, A1=>
      output2_10_EXMPLR, S0=>nx1169);
   ix822 : mux21_ni port map ( Y=>nx821, A0=>q_cache_arr_1_11, A1=>
      output2_11_EXMPLR, S0=>nx1169);
   ix832 : mux21_ni port map ( Y=>nx831, A0=>q_cache_arr_1_12, A1=>
      output2_12_EXMPLR, S0=>nx1171);
   ix842 : mux21_ni port map ( Y=>nx841, A0=>q_cache_arr_1_13, A1=>
      output2_13_EXMPLR, S0=>nx1171);
   ix852 : mux21_ni port map ( Y=>nx851, A0=>q_cache_arr_1_14, A1=>
      output2_14_EXMPLR, S0=>nx1171);
   ix862 : mux21_ni port map ( Y=>nx861, A0=>q_cache_arr_1_15, A1=>
      output2_15_EXMPLR, S0=>nx1171);
   ix552 : mux21_ni port map ( Y=>nx551, A0=>q_cache_arr_0_0, A1=>
      output1_0_EXMPLR, S0=>nx1171);
   ix562 : mux21_ni port map ( Y=>nx561, A0=>q_cache_arr_0_1, A1=>
      output1_1_EXMPLR, S0=>nx1171);
   ix572 : mux21_ni port map ( Y=>nx571, A0=>q_cache_arr_0_2, A1=>
      output1_2_EXMPLR, S0=>nx1171);
   ix582 : mux21_ni port map ( Y=>nx581, A0=>q_cache_arr_0_3, A1=>
      output1_3_EXMPLR, S0=>nx1173);
   ix592 : mux21_ni port map ( Y=>nx591, A0=>q_cache_arr_0_4, A1=>
      output1_4_EXMPLR, S0=>nx1173);
   ix602 : mux21_ni port map ( Y=>nx601, A0=>q_cache_arr_0_5, A1=>
      output1_5_EXMPLR, S0=>nx1173);
   ix612 : mux21_ni port map ( Y=>nx611, A0=>q_cache_arr_0_6, A1=>
      output1_6_EXMPLR, S0=>nx1173);
   ix622 : mux21_ni port map ( Y=>nx621, A0=>q_cache_arr_0_7, A1=>
      output1_7_EXMPLR, S0=>nx1173);
   ix632 : mux21_ni port map ( Y=>nx631, A0=>q_cache_arr_0_8, A1=>
      output1_8_EXMPLR, S0=>nx1173);
   ix642 : mux21_ni port map ( Y=>nx641, A0=>q_cache_arr_0_9, A1=>
      output1_9_EXMPLR, S0=>nx1173);
   ix652 : mux21_ni port map ( Y=>nx651, A0=>q_cache_arr_0_10, A1=>
      output1_10_EXMPLR, S0=>nx1175);
   ix662 : mux21_ni port map ( Y=>nx661, A0=>q_cache_arr_0_11, A1=>
      output1_11_EXMPLR, S0=>nx1175);
   ix672 : mux21_ni port map ( Y=>nx671, A0=>q_cache_arr_0_12, A1=>
      output1_12_EXMPLR, S0=>nx1175);
   ix682 : mux21_ni port map ( Y=>nx681, A0=>q_cache_arr_0_13, A1=>
      output1_13_EXMPLR, S0=>nx1175);
   ix692 : mux21_ni port map ( Y=>nx691, A0=>q_cache_arr_0_14, A1=>
      output1_14_EXMPLR, S0=>nx1175);
   ix702 : mux21_ni port map ( Y=>nx701, A0=>q_cache_arr_0_15, A1=>
      output1_15_EXMPLR, S0=>nx1175);
   ix1166 : inv02 port map ( Y=>nx1167, A=>semi_ready);
   ix1168 : inv02 port map ( Y=>nx1169, A=>semi_ready);
   ix1170 : inv02 port map ( Y=>nx1171, A=>semi_ready);
   ix1172 : inv02 port map ( Y=>nx1173, A=>semi_ready);
   ix1174 : inv02 port map ( Y=>nx1175, A=>semi_ready);
   ix1176 : buf02 port map ( Y=>nx1177, A=>img_load_tmp);
   ix1178 : buf02 port map ( Y=>nx1179, A=>img_load_tmp);
   ix1180 : inv02 port map ( Y=>nx1181, A=>clk);
   ix1182 : inv02 port map ( Y=>nx1183, A=>clk);
   ix1184 : inv02 port map ( Y=>nx1185, A=>nx875);
   ix1186 : inv02 port map ( Y=>nx1187, A=>nx875);
   ix1188 : inv02 port map ( Y=>nx1189, A=>nx875);
   ix1190 : inv02 port map ( Y=>nx1191, A=>nx875);
   ix1192 : inv02 port map ( Y=>nx1193, A=>nx875);
   ix1194 : inv02 port map ( Y=>nx1195, A=>nx875);
end Structural_unfold_2968_0 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity NAdder_16 is
   port (
      a : IN std_logic_vector (15 DOWNTO 0) ;
      b : IN std_logic_vector (15 DOWNTO 0) ;
      cin : IN std_logic ;
      s : OUT std_logic_vector (15 DOWNTO 0) ;
      cout : OUT std_logic) ;
end NAdder_16 ;

architecture DataFlow_unfold_2313 of NAdder_16 is
   signal cout_EXMPLR, nx12, nx16, nx61, nx103, nx105, nx125, nx127, nx129, 
      nx135, nx152, nx153, nx154, nx155, nx156, nx157, nx158, nx159, nx160, 
      nx161, nx162, nx163, nx164, nx165, nx166, nx167, nx168, nx169, nx170, 
      nx38, nx171, nx172, nx173, nx174, nx175, nx176, nx177, nx62, nx178, 
      nx179, nx180, nx97, nx181, nx182, nx183, nx184, nx185, nx186, nx98, 
      nx223, nx225: std_logic ;

begin
   s(14) <= cout_EXMPLR ;
   s(13) <= cout_EXMPLR ;
   s(12) <= cout_EXMPLR ;
   s(11) <= cout_EXMPLR ;
   s(10) <= cout_EXMPLR ;
   s(9) <= cout_EXMPLR ;
   s(8) <= cout_EXMPLR ;
   s(7) <= cout_EXMPLR ;
   s(6) <= cout_EXMPLR ;
   s(5) <= cout_EXMPLR ;
   s(4) <= cout_EXMPLR ;
   s(3) <= cout_EXMPLR ;
   s(2) <= cout_EXMPLR ;
   s(1) <= cout_EXMPLR ;
   s(0) <= cout_EXMPLR ;
   cout <= cout_EXMPLR ;
   ix25 : fake_gnd port map ( Y=>cout_EXMPLR);
   ix13 : xor2 port map ( Y=>nx12, A0=>a(8), A1=>b(8));
   ix104 : xnor2 port map ( Y=>nx103, A0=>a(7), A1=>b(7));
   ix106 : aoi22 port map ( Y=>nx105, A0=>b(6), A1=>a(6), B0=>nx16, B1=>
      nx225);
   ix17 : xor2 port map ( Y=>nx16, A0=>a(6), A1=>b(6));
   ix27 : xor2 port map ( Y=>nx61, A0=>a(2), A1=>b(2));
   ix126 : xnor2 port map ( Y=>nx125, A0=>a(1), A1=>b(1));
   ix128 : nor02_2x port map ( Y=>nx127, A0=>b(0), A1=>a(0));
   ix130 : nand02 port map ( Y=>nx129, A0=>b(1), A1=>a(1));
   ix136 : nand02 port map ( Y=>nx135, A0=>b(7), A1=>a(7));
   ix187 : or02 port map ( Y=>nx152, A0=>a(13), A1=>b(13));
   ix188 : nor02_2x port map ( Y=>nx153, A0=>a(11), A1=>b(11));
   ix189 : nand02_2x port map ( Y=>nx154, A0=>a(11), A1=>b(11));
   ix190 : inv02 port map ( Y=>nx155, A=>a(12));
   ix191 : inv02 port map ( Y=>nx156, A=>b(12));
   ix192 : aoi22 port map ( Y=>nx157, A0=>b(12), A1=>nx155, B0=>a(12), B1=>
      nx156);
   ix193 : nor02_2x port map ( Y=>nx158, A0=>a(13), A1=>b(13));
   ix194 : nor02_2x port map ( Y=>nx159, A0=>nx157, A1=>nx158);
   ix195 : aoi322 port map ( Y=>nx160, A0=>nx152, A1=>b(12), A2=>a(12), B0=>
      a(13), B1=>b(13), C0=>nx98, C1=>nx159);
   ix196 : inv02 port map ( Y=>nx161, A=>a(15));
   ix197 : inv02 port map ( Y=>nx162, A=>b(15));
   ix198 : aoi22 port map ( Y=>nx163, A0=>b(15), A1=>nx161, B0=>a(15), B1=>
      nx162);
   ix199 : and02 port map ( Y=>nx164, A0=>b(14), A1=>a(14));
   ix200 : nor02_2x port map ( Y=>nx165, A0=>nx223, A1=>nx164);
   ix201 : oai21 port map ( Y=>nx166, A0=>b(14), A1=>a(14), B0=>nx223);
   ix202 : nor03_2x port map ( Y=>nx167, A0=>nx223, A1=>b(14), A2=>a(14));
   ix203 : aoi21 port map ( Y=>nx168, A0=>nx223, A1=>nx164, B0=>nx167);
   ix204 : oai21 port map ( Y=>nx169, A0=>nx160, A1=>nx166, B0=>nx168);
   reg_s_15 : ao21 port map ( Y=>s(15), A0=>nx160, A1=>nx165, B0=>nx169);
   ix205 : or02 port map ( Y=>nx170, A0=>a(3), A1=>b(3));
   reg_nx38 : oai21 port map ( Y=>nx38, A0=>nx125, A1=>nx127, B0=>nx129);
   ix206 : aoi332 port map ( Y=>nx171, A0=>nx170, A1=>b(2), A2=>a(2), B0=>
      nx38, B1=>nx61, B2=>nx170, C0=>a(3), C1=>b(3));
   ix207 : inv02 port map ( Y=>nx172, A=>a(4));
   ix208 : inv02 port map ( Y=>nx173, A=>b(4));
   ix209 : aoi22 port map ( Y=>nx174, A0=>b(4), A1=>nx172, B0=>a(4), B1=>
      nx173);
   ix210 : nor02_2x port map ( Y=>nx175, A0=>a(5), A1=>b(5));
   ix211 : inv02 port map ( Y=>nx176, A=>a(5));
   ix212 : inv02 port map ( Y=>nx177, A=>b(5));
   reg_nx62 : oai332 port map ( Y=>nx62, A0=>nx171, A1=>nx174, A2=>nx175, B0
      =>nx175, B1=>nx173, B2=>nx172, C0=>nx176, C1=>nx177);
   ix213 : nor02_2x port map ( Y=>nx178, A0=>nx103, A1=>nx105);
   ix214 : inv02 port map ( Y=>nx179, A=>nx135);
   ix215 : and02 port map ( Y=>nx180, A0=>b(8), A1=>a(8));
   reg_nx97 : oai32 port map ( Y=>nx97, A0=>nx178, A1=>nx179, A2=>nx180, B0
      =>nx180, B1=>nx12);
   ix216 : nor02_2x port map ( Y=>nx181, A0=>a(9), A1=>b(9));
   ix217 : and02 port map ( Y=>nx182, A0=>a(9), A1=>b(9));
   ix218 : nor02_2x port map ( Y=>nx183, A0=>b(10), A1=>a(10));
   ix219 : or04 port map ( Y=>nx184, A0=>nx181, A1=>nx182, A2=>nx183, A3=>
      nx153);
   ix220 : or02 port map ( Y=>nx185, A0=>b(10), A1=>a(10));
   ix221 : aoi22 port map ( Y=>nx186, A0=>nx185, A1=>nx182, B0=>b(10), B1=>
      a(10));
   reg_nx98 : oai221 port map ( Y=>nx98, A0=>nx97, A1=>nx184, B0=>nx186, B1
      =>nx153, C0=>nx154);
   ix222 : buf02 port map ( Y=>nx223, A=>nx163);
   ix224 : buf02 port map ( Y=>nx225, A=>nx62);
end DataFlow_unfold_2313 ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity ArgMax is
   port (
      inp : IN std_logic_vector (15 DOWNTO 0) ;
      en : IN std_logic ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      ans : OUT std_logic_vector (3 DOWNTO 0)) ;
end ArgMax ;

architecture DataFlow of ArgMax is
   component NAdder_16
      port (
         a : IN std_logic_vector (15 DOWNTO 0) ;
         b : IN std_logic_vector (15 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (15 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal ans_3_EXMPLR, ans_2_EXMPLR, ans_1_EXMPLR, ans_0_EXMPLR, 
      reg_val_out_15, reg_val_out_14, reg_val_out_13, reg_val_out_12, 
      reg_val_out_11, reg_val_out_10, reg_val_out_9, reg_val_out_8, 
      reg_val_out_7, reg_val_out_6, reg_val_out_5, reg_val_out_4, 
      reg_val_out_3, reg_val_out_2, reg_val_out_1, reg_val_out_0, 
      compare_in1_inverted_15, compare_in1_inverted_14, 
      compare_in1_inverted_13, compare_in1_inverted_12, 
      compare_in1_inverted_11, compare_in1_inverted_10, 
      compare_in1_inverted_9, compare_in1_inverted_8, compare_in1_inverted_7, 
      compare_in1_inverted_6, compare_in1_inverted_5, compare_in1_inverted_4, 
      compare_in1_inverted_3, compare_in1_inverted_2, compare_in1_inverted_1, 
      compare_in1_inverted_0, compare_sub_res_15, tmp_15, curr_idx_0, nx54, 
      reg_idx_out_0, curr_idx_1, reg_idx_out_1, curr_idx_2, nx98, 
      reg_idx_out_2, curr_idx_3, nx157, reg_idx_out_3, nx140, nx152, nx164, 
      nx176, nx188, nx200, nx212, nx224, nx236, nx248, nx260, nx272, nx284, 
      nx296, nx308, nx165, nx175, nx185, nx195, nx205, nx215, nx225, nx235, 
      nx245, nx255, nx265, nx275, nx285, nx295, nx305, nx315, nx325, nx335, 
      nx345, nx355, nx365, nx375, nx385, nx395, nx405, nx411, nx482, nx484, 
      nx486, nx503, nx556, nx558, nx560, nx562, nx564, nx566, nx568, nx570: 
   std_logic ;
   
   signal DANGLING : std_logic_vector (15 downto 0 );

begin
   ans(3) <= ans_3_EXMPLR ;
   ans(2) <= ans_2_EXMPLR ;
   ans(1) <= ans_1_EXMPLR ;
   ans(0) <= ans_0_EXMPLR ;
   compare_DoSubtraction : NAdder_16 port map ( a(15)=>reg_val_out_15, a(14)
      =>reg_val_out_14, a(13)=>reg_val_out_13, a(12)=>reg_val_out_12, a(11)
      =>reg_val_out_11, a(10)=>reg_val_out_10, a(9)=>reg_val_out_9, a(8)=>
      reg_val_out_8, a(7)=>reg_val_out_7, a(6)=>reg_val_out_6, a(5)=>
      reg_val_out_5, a(4)=>reg_val_out_4, a(3)=>reg_val_out_3, a(2)=>
      reg_val_out_2, a(1)=>reg_val_out_1, a(0)=>reg_val_out_0, b(15)=>
      compare_in1_inverted_15, b(14)=>compare_in1_inverted_14, b(13)=>
      compare_in1_inverted_13, b(12)=>compare_in1_inverted_12, b(11)=>
      compare_in1_inverted_11, b(10)=>compare_in1_inverted_10, b(9)=>
      compare_in1_inverted_9, b(8)=>compare_in1_inverted_8, b(7)=>
      compare_in1_inverted_7, b(6)=>compare_in1_inverted_6, b(5)=>
      compare_in1_inverted_5, b(4)=>compare_in1_inverted_4, b(3)=>
      compare_in1_inverted_3, b(2)=>compare_in1_inverted_2, b(1)=>
      compare_in1_inverted_1, b(0)=>compare_in1_inverted_0, cin=>tmp_15, 
      s(15)=>compare_sub_res_15, s(14)=>DANGLING(0), s(13)=>DANGLING(1), 
      s(12)=>DANGLING(2), s(11)=>DANGLING(3), s(10)=>DANGLING(4), s(9)=>
      DANGLING(5), s(8)=>DANGLING(6), s(7)=>DANGLING(7), s(6)=>DANGLING(8), 
      s(5)=>DANGLING(9), s(4)=>DANGLING(10), s(3)=>DANGLING(11), s(2)=>
      DANGLING(12), s(1)=>DANGLING(13), s(0)=>DANGLING(14), cout=>DANGLING(
      15));
   ix115 : fake_vcc port map ( Y=>tmp_15);
   valReg_reg_q_0 : dffr port map ( Q=>reg_val_out_0, QB=>OPEN, D=>nx255, 
      CLK=>clk, R=>rst);
   ix256 : mux21_ni port map ( Y=>nx255, A0=>reg_val_out_0, A1=>nx140, S0=>
      nx558);
   ix55 : oai22 port map ( Y=>nx54, A0=>compare_sub_res_15, A1=>nx405, B0=>
      compare_in1_inverted_15, B1=>reg_val_out_15);
   ix176 : aoi21 port map ( Y=>nx175, A0=>nx558, A1=>compare_in1_inverted_15, 
      B0=>nx411);
   ix410 : inv01 port map ( Y=>compare_in1_inverted_15, A=>inp(15));
   valReg_reg_q_15 : dffs_ni port map ( Q=>reg_val_out_15, QB=>nx411, D=>
      nx175, CLK=>clk, S=>rst);
   valReg_reg_q_1 : dffr port map ( Q=>reg_val_out_1, QB=>OPEN, D=>nx265, 
      CLK=>clk, R=>rst);
   ix266 : mux21_ni port map ( Y=>nx265, A0=>reg_val_out_1, A1=>nx152, S0=>
      nx558);
   valReg_reg_q_2 : dffr port map ( Q=>reg_val_out_2, QB=>OPEN, D=>nx275, 
      CLK=>clk, R=>rst);
   ix276 : mux21_ni port map ( Y=>nx275, A0=>reg_val_out_2, A1=>nx164, S0=>
      nx558);
   valReg_reg_q_3 : dffr port map ( Q=>reg_val_out_3, QB=>OPEN, D=>nx285, 
      CLK=>clk, R=>rst);
   ix286 : mux21_ni port map ( Y=>nx285, A0=>reg_val_out_3, A1=>nx176, S0=>
      nx558);
   valReg_reg_q_4 : dffr port map ( Q=>reg_val_out_4, QB=>OPEN, D=>nx295, 
      CLK=>clk, R=>rst);
   ix296 : mux21_ni port map ( Y=>nx295, A0=>reg_val_out_4, A1=>nx188, S0=>
      nx558);
   valReg_reg_q_5 : dffr port map ( Q=>reg_val_out_5, QB=>OPEN, D=>nx305, 
      CLK=>clk, R=>rst);
   ix306 : mux21_ni port map ( Y=>nx305, A0=>reg_val_out_5, A1=>nx200, S0=>
      nx558);
   valReg_reg_q_6 : dffr port map ( Q=>reg_val_out_6, QB=>OPEN, D=>nx315, 
      CLK=>clk, R=>rst);
   ix316 : mux21_ni port map ( Y=>nx315, A0=>reg_val_out_6, A1=>nx212, S0=>
      nx560);
   valReg_reg_q_7 : dffr port map ( Q=>reg_val_out_7, QB=>OPEN, D=>nx325, 
      CLK=>clk, R=>rst);
   ix326 : mux21_ni port map ( Y=>nx325, A0=>reg_val_out_7, A1=>nx224, S0=>
      nx560);
   valReg_reg_q_8 : dffr port map ( Q=>reg_val_out_8, QB=>OPEN, D=>nx335, 
      CLK=>clk, R=>rst);
   ix336 : mux21_ni port map ( Y=>nx335, A0=>reg_val_out_8, A1=>nx236, S0=>
      nx560);
   valReg_reg_q_9 : dffr port map ( Q=>reg_val_out_9, QB=>OPEN, D=>nx345, 
      CLK=>clk, R=>rst);
   ix346 : mux21_ni port map ( Y=>nx345, A0=>reg_val_out_9, A1=>nx248, S0=>
      nx560);
   valReg_reg_q_10 : dffr port map ( Q=>reg_val_out_10, QB=>OPEN, D=>nx355, 
      CLK=>clk, R=>rst);
   ix356 : mux21_ni port map ( Y=>nx355, A0=>reg_val_out_10, A1=>nx260, S0=>
      nx560);
   valReg_reg_q_11 : dffr port map ( Q=>reg_val_out_11, QB=>OPEN, D=>nx365, 
      CLK=>clk, R=>rst);
   ix366 : mux21_ni port map ( Y=>nx365, A0=>reg_val_out_11, A1=>nx272, S0=>
      nx560);
   valReg_reg_q_12 : dffr port map ( Q=>reg_val_out_12, QB=>OPEN, D=>nx375, 
      CLK=>clk, R=>rst);
   ix376 : mux21_ni port map ( Y=>nx375, A0=>reg_val_out_12, A1=>nx284, S0=>
      nx560);
   valReg_reg_q_13 : dffr port map ( Q=>reg_val_out_13, QB=>OPEN, D=>nx385, 
      CLK=>clk, R=>rst);
   ix386 : mux21_ni port map ( Y=>nx385, A0=>reg_val_out_13, A1=>nx296, S0=>
      nx562);
   valReg_reg_q_14 : dffr port map ( Q=>reg_val_out_14, QB=>OPEN, D=>nx395, 
      CLK=>clk, R=>rst);
   ix396 : mux21_ni port map ( Y=>nx395, A0=>reg_val_out_14, A1=>nx308, S0=>
      nx562);
   reg_curr_idx_0 : dffr port map ( Q=>curr_idx_0, QB=>OPEN, D=>nx165, CLK=>
      clk, R=>rst);
   idxReg_reg_q_0 : dffr port map ( Q=>reg_idx_out_0, QB=>OPEN, D=>nx185, 
      CLK=>clk, R=>rst);
   ix186 : mux21_ni port map ( Y=>nx185, A0=>reg_idx_out_0, A1=>ans_0_EXMPLR, 
      S0=>nx562);
   ix196 : mux21 port map ( Y=>nx195, A0=>nx482, A1=>nx484, S0=>nx562);
   reg_curr_idx_1 : dffr port map ( Q=>curr_idx_1, QB=>nx482, D=>nx195, CLK
      =>clk, R=>rst);
   ix485 : oai21 port map ( Y=>nx484, A0=>curr_idx_0, A1=>curr_idx_1, B0=>
      nx486);
   ix487 : nand02 port map ( Y=>nx486, A0=>curr_idx_1, A1=>curr_idx_0);
   idxReg_reg_q_1 : dffr port map ( Q=>reg_idx_out_1, QB=>OPEN, D=>nx205, 
      CLK=>clk, R=>rst);
   ix206 : mux21_ni port map ( Y=>nx205, A0=>reg_idx_out_1, A1=>ans_1_EXMPLR, 
      S0=>nx562);
   reg_curr_idx_2 : dffr port map ( Q=>curr_idx_2, QB=>OPEN, D=>nx215, CLK=>
      clk, R=>rst);
   ix216 : mux21_ni port map ( Y=>nx215, A0=>curr_idx_2, A1=>nx98, S0=>nx562
   );
   ix99 : xnor2 port map ( Y=>nx98, A0=>curr_idx_2, A1=>nx486);
   idxReg_reg_q_2 : dffr port map ( Q=>reg_idx_out_2, QB=>OPEN, D=>nx225, 
      CLK=>clk, R=>rst);
   ix226 : mux21_ni port map ( Y=>nx225, A0=>reg_idx_out_2, A1=>ans_2_EXMPLR, 
      S0=>nx562);
   reg_curr_idx_3 : dffr port map ( Q=>curr_idx_3, QB=>OPEN, D=>nx235, CLK=>
      clk, R=>rst);
   ix236 : mux21_ni port map ( Y=>nx235, A0=>curr_idx_3, A1=>nx157, S0=>
      nx564);
   ix120 : xnor2 port map ( Y=>nx157, A0=>curr_idx_3, A1=>nx503);
   ix504 : nand03 port map ( Y=>nx503, A0=>curr_idx_2, A1=>curr_idx_1, A2=>
      curr_idx_0);
   idxReg_reg_q_3 : dffr port map ( Q=>reg_idx_out_3, QB=>OPEN, D=>nx245, 
      CLK=>clk, R=>rst);
   ix246 : mux21_ni port map ( Y=>nx245, A0=>reg_idx_out_3, A1=>ans_3_EXMPLR, 
      S0=>nx564);
   ix510 : inv01 port map ( Y=>compare_in1_inverted_0, A=>inp(0));
   ix512 : inv01 port map ( Y=>compare_in1_inverted_1, A=>inp(1));
   ix514 : inv01 port map ( Y=>compare_in1_inverted_2, A=>inp(2));
   ix516 : inv01 port map ( Y=>compare_in1_inverted_3, A=>inp(3));
   ix518 : inv01 port map ( Y=>compare_in1_inverted_4, A=>inp(4));
   ix520 : inv01 port map ( Y=>compare_in1_inverted_5, A=>inp(5));
   ix522 : inv01 port map ( Y=>compare_in1_inverted_6, A=>inp(6));
   ix524 : inv01 port map ( Y=>compare_in1_inverted_7, A=>inp(7));
   ix526 : inv01 port map ( Y=>compare_in1_inverted_8, A=>inp(8));
   ix528 : inv01 port map ( Y=>compare_in1_inverted_9, A=>inp(9));
   ix530 : inv01 port map ( Y=>compare_in1_inverted_10, A=>inp(10));
   ix532 : inv01 port map ( Y=>compare_in1_inverted_11, A=>inp(11));
   ix534 : inv01 port map ( Y=>compare_in1_inverted_12, A=>inp(12));
   ix536 : inv01 port map ( Y=>compare_in1_inverted_13, A=>inp(13));
   ix538 : inv01 port map ( Y=>compare_in1_inverted_14, A=>inp(14));
   ix141 : mux21_ni port map ( Y=>nx140, A0=>reg_val_out_0, A1=>inp(0), S0=>
      nx566);
   ix406 : xnor2 port map ( Y=>nx405, A0=>inp(15), A1=>nx411);
   ix153 : mux21_ni port map ( Y=>nx152, A0=>reg_val_out_1, A1=>inp(1), S0=>
      nx566);
   ix165 : mux21_ni port map ( Y=>nx164, A0=>reg_val_out_2, A1=>inp(2), S0=>
      nx566);
   ix177 : mux21_ni port map ( Y=>nx176, A0=>reg_val_out_3, A1=>inp(3), S0=>
      nx566);
   ix189 : mux21_ni port map ( Y=>nx188, A0=>reg_val_out_4, A1=>inp(4), S0=>
      nx566);
   ix201 : mux21_ni port map ( Y=>nx200, A0=>reg_val_out_5, A1=>inp(5), S0=>
      nx566);
   ix213 : mux21_ni port map ( Y=>nx212, A0=>reg_val_out_6, A1=>inp(6), S0=>
      nx566);
   ix225 : mux21_ni port map ( Y=>nx224, A0=>reg_val_out_7, A1=>inp(7), S0=>
      nx568);
   ix237 : mux21_ni port map ( Y=>nx236, A0=>reg_val_out_8, A1=>inp(8), S0=>
      nx568);
   ix249 : mux21_ni port map ( Y=>nx248, A0=>reg_val_out_9, A1=>inp(9), S0=>
      nx568);
   ix261 : mux21_ni port map ( Y=>nx260, A0=>reg_val_out_10, A1=>inp(10), S0
      =>nx568);
   ix273 : mux21_ni port map ( Y=>nx272, A0=>reg_val_out_11, A1=>inp(11), S0
      =>nx568);
   ix285 : mux21_ni port map ( Y=>nx284, A0=>reg_val_out_12, A1=>inp(12), S0
      =>nx568);
   ix297 : mux21_ni port map ( Y=>nx296, A0=>reg_val_out_13, A1=>inp(13), S0
      =>nx568);
   ix309 : mux21_ni port map ( Y=>nx308, A0=>reg_val_out_14, A1=>inp(14), S0
      =>nx570);
   ix67 : mux21_ni port map ( Y=>ans_0_EXMPLR, A0=>reg_idx_out_0, A1=>
      curr_idx_0, S0=>nx570);
   ix166 : xor2 port map ( Y=>nx165, A0=>curr_idx_0, A1=>nx564);
   ix91 : mux21_ni port map ( Y=>ans_1_EXMPLR, A0=>reg_idx_out_1, A1=>
      curr_idx_1, S0=>nx570);
   ix119 : mux21_ni port map ( Y=>ans_2_EXMPLR, A0=>reg_idx_out_2, A1=>
      curr_idx_2, S0=>nx570);
   ix133 : mux21_ni port map ( Y=>ans_3_EXMPLR, A0=>reg_idx_out_3, A1=>
      curr_idx_3, S0=>nx570);
   ix555 : inv01 port map ( Y=>nx556, A=>en);
   ix557 : inv02 port map ( Y=>nx558, A=>nx556);
   ix559 : inv02 port map ( Y=>nx560, A=>nx556);
   ix561 : inv02 port map ( Y=>nx562, A=>nx556);
   ix563 : inv02 port map ( Y=>nx564, A=>nx556);
   ix565 : inv02 port map ( Y=>nx566, A=>nx54);
   ix567 : inv02 port map ( Y=>nx568, A=>nx54);
   ix569 : inv02 port map ( Y=>nx570, A=>nx54);
end DataFlow ;

library adk; use adk.adk_components.all; library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity DCNNChip is
   port (
      clk : IN std_logic ;
      reset : IN std_logic ;
      io_ready_in : IN std_logic ;
      io_done_out : OUT std_logic ;
      mem_read_out : OUT std_logic ;
      mem_write_out : OUT std_logic ;
      mem_addr_out : OUT std_logic_vector (15 DOWNTO 0) ;
      mem_data_in : IN std_logic_vector (15 DOWNTO 0) ;
      mem_data_out : OUT std_logic_vector (15 DOWNTO 0)) ;
end DCNNChip ;

architecture Structural of DCNNChip is
   component Controller_16_16_5_16
      port (
         clk : IN std_logic ;
         reset : IN std_logic ;
         io_ready_in : IN std_logic ;
         io_done_out : OUT std_logic ;
         mem_data_in : IN std_logic_vector (15 DOWNTO 0) ;
         mem_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
         mem_addr_out : OUT std_logic_vector (15 DOWNTO 0) ;
         mem_write_out : OUT std_logic ;
         mem_read_out : OUT std_logic ;
         wind_en : OUT std_logic ;
         wind_rst : OUT std_logic ;
         wind_col_in_4_15 : OUT std_logic ;
         wind_col_in_4_14 : OUT std_logic ;
         wind_col_in_4_13 : OUT std_logic ;
         wind_col_in_4_12 : OUT std_logic ;
         wind_col_in_4_11 : OUT std_logic ;
         wind_col_in_4_10 : OUT std_logic ;
         wind_col_in_4_9 : OUT std_logic ;
         wind_col_in_4_8 : OUT std_logic ;
         wind_col_in_4_7 : OUT std_logic ;
         wind_col_in_4_6 : OUT std_logic ;
         wind_col_in_4_5 : OUT std_logic ;
         wind_col_in_4_4 : OUT std_logic ;
         wind_col_in_4_3 : OUT std_logic ;
         wind_col_in_4_2 : OUT std_logic ;
         wind_col_in_4_1 : OUT std_logic ;
         wind_col_in_4_0 : OUT std_logic ;
         wind_col_in_3_15 : OUT std_logic ;
         wind_col_in_3_14 : OUT std_logic ;
         wind_col_in_3_13 : OUT std_logic ;
         wind_col_in_3_12 : OUT std_logic ;
         wind_col_in_3_11 : OUT std_logic ;
         wind_col_in_3_10 : OUT std_logic ;
         wind_col_in_3_9 : OUT std_logic ;
         wind_col_in_3_8 : OUT std_logic ;
         wind_col_in_3_7 : OUT std_logic ;
         wind_col_in_3_6 : OUT std_logic ;
         wind_col_in_3_5 : OUT std_logic ;
         wind_col_in_3_4 : OUT std_logic ;
         wind_col_in_3_3 : OUT std_logic ;
         wind_col_in_3_2 : OUT std_logic ;
         wind_col_in_3_1 : OUT std_logic ;
         wind_col_in_3_0 : OUT std_logic ;
         wind_col_in_2_15 : OUT std_logic ;
         wind_col_in_2_14 : OUT std_logic ;
         wind_col_in_2_13 : OUT std_logic ;
         wind_col_in_2_12 : OUT std_logic ;
         wind_col_in_2_11 : OUT std_logic ;
         wind_col_in_2_10 : OUT std_logic ;
         wind_col_in_2_9 : OUT std_logic ;
         wind_col_in_2_8 : OUT std_logic ;
         wind_col_in_2_7 : OUT std_logic ;
         wind_col_in_2_6 : OUT std_logic ;
         wind_col_in_2_5 : OUT std_logic ;
         wind_col_in_2_4 : OUT std_logic ;
         wind_col_in_2_3 : OUT std_logic ;
         wind_col_in_2_2 : OUT std_logic ;
         wind_col_in_2_1 : OUT std_logic ;
         wind_col_in_2_0 : OUT std_logic ;
         wind_col_in_1_15 : OUT std_logic ;
         wind_col_in_1_14 : OUT std_logic ;
         wind_col_in_1_13 : OUT std_logic ;
         wind_col_in_1_12 : OUT std_logic ;
         wind_col_in_1_11 : OUT std_logic ;
         wind_col_in_1_10 : OUT std_logic ;
         wind_col_in_1_9 : OUT std_logic ;
         wind_col_in_1_8 : OUT std_logic ;
         wind_col_in_1_7 : OUT std_logic ;
         wind_col_in_1_6 : OUT std_logic ;
         wind_col_in_1_5 : OUT std_logic ;
         wind_col_in_1_4 : OUT std_logic ;
         wind_col_in_1_3 : OUT std_logic ;
         wind_col_in_1_2 : OUT std_logic ;
         wind_col_in_1_1 : OUT std_logic ;
         wind_col_in_1_0 : OUT std_logic ;
         wind_col_in_0_15 : OUT std_logic ;
         wind_col_in_0_14 : OUT std_logic ;
         wind_col_in_0_13 : OUT std_logic ;
         wind_col_in_0_12 : OUT std_logic ;
         wind_col_in_0_11 : OUT std_logic ;
         wind_col_in_0_10 : OUT std_logic ;
         wind_col_in_0_9 : OUT std_logic ;
         wind_col_in_0_8 : OUT std_logic ;
         wind_col_in_0_7 : OUT std_logic ;
         wind_col_in_0_6 : OUT std_logic ;
         wind_col_in_0_5 : OUT std_logic ;
         wind_col_in_0_4 : OUT std_logic ;
         wind_col_in_0_3 : OUT std_logic ;
         wind_col_in_0_2 : OUT std_logic ;
         wind_col_in_0_1 : OUT std_logic ;
         wind_col_in_0_0 : OUT std_logic ;
         filter_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
         filter_ready_out : OUT std_logic ;
         filter_reset : OUT std_logic ;
         comp_unit_ready : OUT std_logic ;
         comp_unit_operation : OUT std_logic ;
         comp_unit_flt_size : OUT std_logic ;
         comp_unit_relu : OUT std_logic ;
         comp_unit_data1_out : OUT std_logic_vector (15 DOWNTO 0) ;
         comp_unit_data2_out : OUT std_logic_vector (15 DOWNTO 0) ;
         comp_unit_buffer_finished : IN std_logic ;
         comp_unit_finished : IN std_logic ;
         comp_unit_data1_in : IN std_logic_vector (15 DOWNTO 0) ;
         comp_unit_data2_in : IN std_logic_vector (15 DOWNTO 0) ;
         argmax_ready : OUT std_logic ;
         argmax_data_out : OUT std_logic_vector (15 DOWNTO 0) ;
         argmax_data_in : IN std_logic_vector (15 DOWNTO 0)) ;
   
   end component ;
   component ComputationBlock
      port (
         img_data_col_0 : IN std_logic_vector (15 DOWNTO 0) ;
         img_data_col_1 : IN std_logic_vector (15 DOWNTO 0) ;
         img_data_col_2 : IN std_logic_vector (15 DOWNTO 0) ;
         img_data_col_3 : IN std_logic_vector (15 DOWNTO 0) ;
         img_data_col_4 : IN std_logic_vector (15 DOWNTO 0) ;
         img_load : IN std_logic ;
         img_reset : IN std_logic ;
         filter_data_word : IN std_logic_vector (15 DOWNTO 0) ;
         filter_load : IN std_logic ;
         filter_reset : IN std_logic ;
         start : IN std_logic ;
         operation : IN std_logic ;
         compute_relu : IN std_logic ;
         filter_size : IN std_logic ;
         output1_init : IN std_logic_vector (15 DOWNTO 0) ;
         output2_init : IN std_logic_vector (15 DOWNTO 0) ;
         output1 : OUT std_logic_vector (15 DOWNTO 0) ;
         output2 : OUT std_logic_vector (15 DOWNTO 0) ;
         buffer_ready : OUT std_logic ;
         ready : OUT std_logic ;
         clk : IN std_logic ;
         en : IN std_logic ;
         reset : IN std_logic) ;
   end component ;
   component ArgMax
      port (
         inp : IN std_logic_vector (15 DOWNTO 0) ;
         en : IN std_logic ;
         clk : IN std_logic ;
         rst : IN std_logic ;
         ans : OUT std_logic_vector (3 DOWNTO 0)) ;
   end component ;
   signal image_wind_en, image_wind_col_4_15, image_wind_col_4_14, 
      image_wind_col_4_13, image_wind_col_4_12, image_wind_col_4_11, 
      image_wind_col_4_10, image_wind_col_4_9, image_wind_col_4_8, 
      image_wind_col_4_7, image_wind_col_4_6, image_wind_col_4_5, 
      image_wind_col_4_4, image_wind_col_4_3, image_wind_col_4_2, 
      image_wind_col_4_1, image_wind_col_4_0, image_wind_col_3_15, 
      image_wind_col_3_14, image_wind_col_3_13, image_wind_col_3_12, 
      image_wind_col_3_11, image_wind_col_3_10, image_wind_col_3_9, 
      image_wind_col_3_8, image_wind_col_3_7, image_wind_col_3_6, 
      image_wind_col_3_5, image_wind_col_3_4, image_wind_col_3_3, 
      image_wind_col_3_2, image_wind_col_3_1, image_wind_col_3_0, 
      image_wind_col_2_15, image_wind_col_2_14, image_wind_col_2_13, 
      image_wind_col_2_12, image_wind_col_2_11, image_wind_col_2_10, 
      image_wind_col_2_9, image_wind_col_2_8, image_wind_col_2_7, 
      image_wind_col_2_6, image_wind_col_2_5, image_wind_col_2_4, 
      image_wind_col_2_3, image_wind_col_2_2, image_wind_col_2_1, 
      image_wind_col_2_0, image_wind_col_1_15, image_wind_col_1_14, 
      image_wind_col_1_13, image_wind_col_1_12, image_wind_col_1_11, 
      image_wind_col_1_10, image_wind_col_1_9, image_wind_col_1_8, 
      image_wind_col_1_7, image_wind_col_1_6, image_wind_col_1_5, 
      image_wind_col_1_4, image_wind_col_1_3, image_wind_col_1_2, 
      image_wind_col_1_1, image_wind_col_1_0, image_wind_col_0_15, 
      image_wind_col_0_14, image_wind_col_0_13, image_wind_col_0_12, 
      image_wind_col_0_11, image_wind_col_0_10, image_wind_col_0_9, 
      image_wind_col_0_8, image_wind_col_0_7, image_wind_col_0_6, 
      image_wind_col_0_5, image_wind_col_0_4, image_wind_col_0_3, 
      image_wind_col_0_2, image_wind_col_0_1, image_wind_col_0_0, 
      filter_window_ready, filter_window_data_15, filter_window_data_14, 
      filter_window_data_13, filter_window_data_12, filter_window_data_11, 
      filter_window_data_10, filter_window_data_9, filter_window_data_8, 
      filter_window_data_7, filter_window_data_6, filter_window_data_5, 
      filter_window_data_4, filter_window_data_3, filter_window_data_2, 
      filter_window_data_1, filter_window_data_0, comp_unit_ready, 
      comp_unit_operation, comp_unit_relu, comp_unit_flt_size, 
      comp_unit_finished, comp_unit_bias_1_15, comp_unit_bias_1_14, 
      comp_unit_bias_1_13, comp_unit_bias_1_12, comp_unit_bias_1_11, 
      comp_unit_bias_1_10, comp_unit_bias_1_9, comp_unit_bias_1_8, 
      comp_unit_bias_1_7, comp_unit_bias_1_6, comp_unit_bias_1_5, 
      comp_unit_bias_1_4, comp_unit_bias_1_3, comp_unit_bias_1_2, 
      comp_unit_bias_1_1, comp_unit_bias_1_0, comp_unit_bias_2_15, 
      comp_unit_bias_2_14, comp_unit_bias_2_13, comp_unit_bias_2_12, 
      comp_unit_bias_2_11, comp_unit_bias_2_10, comp_unit_bias_2_9, 
      comp_unit_bias_2_8, comp_unit_bias_2_7, comp_unit_bias_2_6, 
      comp_unit_bias_2_5, comp_unit_bias_2_4, comp_unit_bias_2_3, 
      comp_unit_bias_2_2, comp_unit_bias_2_1, comp_unit_bias_2_0, 
      comp_unit_result_1_15, comp_unit_result_1_14, comp_unit_result_1_13, 
      comp_unit_result_1_12, comp_unit_result_1_11, comp_unit_result_1_10, 
      comp_unit_result_1_9, comp_unit_result_1_8, comp_unit_result_1_7, 
      comp_unit_result_1_6, comp_unit_result_1_5, comp_unit_result_1_4, 
      comp_unit_result_1_3, comp_unit_result_1_2, comp_unit_result_1_1, 
      comp_unit_result_1_0, comp_unit_result_2_15, comp_unit_result_2_14, 
      comp_unit_result_2_13, comp_unit_result_2_12, comp_unit_result_2_11, 
      comp_unit_result_2_10, comp_unit_result_2_9, comp_unit_result_2_8, 
      comp_unit_result_2_7, comp_unit_result_2_6, comp_unit_result_2_5, 
      comp_unit_result_2_4, comp_unit_result_2_3, comp_unit_result_2_2, 
      comp_unit_result_2_1, comp_unit_result_2_0, controller_bias_1_15, 
      controller_bias_1_14, controller_bias_1_13, controller_bias_1_12, 
      controller_bias_1_11, controller_bias_1_10, controller_bias_1_9, 
      controller_bias_1_8, controller_bias_1_7, controller_bias_1_6, 
      controller_bias_1_5, controller_bias_1_4, controller_bias_1_3, 
      controller_bias_1_2, controller_bias_1_1, controller_bias_1_0, 
      controller_bias_2_15, controller_bias_2_14, controller_bias_2_13, 
      controller_bias_2_12, controller_bias_2_11, controller_bias_2_10, 
      controller_bias_2_9, controller_bias_2_8, controller_bias_2_7, 
      controller_bias_2_6, controller_bias_2_5, controller_bias_2_4, 
      controller_bias_2_3, controller_bias_2_2, controller_bias_2_1, 
      controller_bias_2_0, controller_result_1_15, controller_result_1_14, 
      controller_result_1_13, controller_result_1_12, controller_result_1_11, 
      controller_result_1_10, controller_result_1_9, controller_result_1_8, 
      controller_result_1_7, controller_result_1_6, controller_result_1_5, 
      controller_result_1_4, controller_result_1_3, controller_result_1_2, 
      controller_result_1_1, controller_result_1_0, controller_result_2_15, 
      controller_result_2_14, controller_result_2_13, controller_result_2_12, 
      controller_result_2_11, controller_result_2_10, controller_result_2_9, 
      controller_result_2_8, controller_result_2_7, controller_result_2_6, 
      controller_result_2_5, controller_result_2_4, controller_result_2_3, 
      controller_result_2_2, controller_result_2_1, controller_result_2_0, 
      argmax_ready, argmax_data_outof_controller_15, 
      argmax_data_outof_controller_14, argmax_data_outof_controller_13, 
      argmax_data_outof_controller_12, argmax_data_outof_controller_11, 
      argmax_data_outof_controller_10, argmax_data_outof_controller_9, 
      argmax_data_outof_controller_8, argmax_data_outof_controller_7, 
      argmax_data_outof_controller_6, argmax_data_outof_controller_5, 
      argmax_data_outof_controller_4, argmax_data_outof_controller_3, 
      argmax_data_outof_controller_2, argmax_data_outof_controller_1, 
      argmax_data_outof_controller_0, argmax_data_out_3, argmax_data_out_2, 
      argmax_data_out_1, argmax_data_out_0, io_done_out_EXMPLR, PWR, 
      flt_size_out_0, nx495, nx584, nx594, nx610, nx612, nx614, nx616, nx618, 
      nx620, nx622, nx624, nx626, nx628, nx630, nx632: std_logic ;
   
   signal DANGLING : std_logic_vector (3 downto 0 );

begin
   io_done_out <= io_done_out_EXMPLR ;
   controller_inst : Controller_16_16_5_16 port map ( clk=>clk, reset=>reset, 
      io_ready_in=>io_ready_in, io_done_out=>DANGLING(0), mem_data_in(15)=>
      mem_data_in(15), mem_data_in(14)=>mem_data_in(14), mem_data_in(13)=>
      mem_data_in(13), mem_data_in(12)=>mem_data_in(12), mem_data_in(11)=>
      mem_data_in(11), mem_data_in(10)=>mem_data_in(10), mem_data_in(9)=>
      mem_data_in(9), mem_data_in(8)=>mem_data_in(8), mem_data_in(7)=>
      mem_data_in(7), mem_data_in(6)=>mem_data_in(6), mem_data_in(5)=>
      mem_data_in(5), mem_data_in(4)=>mem_data_in(4), mem_data_in(3)=>
      mem_data_in(3), mem_data_in(2)=>mem_data_in(2), mem_data_in(1)=>
      mem_data_in(1), mem_data_in(0)=>mem_data_in(0), mem_data_out(15)=>
      mem_data_out(15), mem_data_out(14)=>mem_data_out(14), mem_data_out(13)
      =>mem_data_out(13), mem_data_out(12)=>mem_data_out(12), 
      mem_data_out(11)=>mem_data_out(11), mem_data_out(10)=>mem_data_out(10), 
      mem_data_out(9)=>mem_data_out(9), mem_data_out(8)=>mem_data_out(8), 
      mem_data_out(7)=>mem_data_out(7), mem_data_out(6)=>mem_data_out(6), 
      mem_data_out(5)=>mem_data_out(5), mem_data_out(4)=>mem_data_out(4), 
      mem_data_out(3)=>mem_data_out(3), mem_data_out(2)=>mem_data_out(2), 
      mem_data_out(1)=>mem_data_out(1), mem_data_out(0)=>mem_data_out(0), 
      mem_addr_out(15)=>mem_addr_out(15), mem_addr_out(14)=>mem_addr_out(14), 
      mem_addr_out(13)=>mem_addr_out(13), mem_addr_out(12)=>mem_addr_out(12), 
      mem_addr_out(11)=>mem_addr_out(11), mem_addr_out(10)=>mem_addr_out(10), 
      mem_addr_out(9)=>mem_addr_out(9), mem_addr_out(8)=>mem_addr_out(8), 
      mem_addr_out(7)=>mem_addr_out(7), mem_addr_out(6)=>mem_addr_out(6), 
      mem_addr_out(5)=>mem_addr_out(5), mem_addr_out(4)=>mem_addr_out(4), 
      mem_addr_out(3)=>mem_addr_out(3), mem_addr_out(2)=>mem_addr_out(2), 
      mem_addr_out(1)=>mem_addr_out(1), mem_addr_out(0)=>mem_addr_out(0), 
      mem_write_out=>mem_write_out, mem_read_out=>mem_read_out, wind_en=>
      image_wind_en, wind_rst=>DANGLING(1), wind_col_in_4_15=>
      image_wind_col_4_15, wind_col_in_4_14=>image_wind_col_4_14, 
      wind_col_in_4_13=>image_wind_col_4_13, wind_col_in_4_12=>
      image_wind_col_4_12, wind_col_in_4_11=>image_wind_col_4_11, 
      wind_col_in_4_10=>image_wind_col_4_10, wind_col_in_4_9=>
      image_wind_col_4_9, wind_col_in_4_8=>image_wind_col_4_8, 
      wind_col_in_4_7=>image_wind_col_4_7, wind_col_in_4_6=>
      image_wind_col_4_6, wind_col_in_4_5=>image_wind_col_4_5, 
      wind_col_in_4_4=>image_wind_col_4_4, wind_col_in_4_3=>
      image_wind_col_4_3, wind_col_in_4_2=>image_wind_col_4_2, 
      wind_col_in_4_1=>image_wind_col_4_1, wind_col_in_4_0=>
      image_wind_col_4_0, wind_col_in_3_15=>image_wind_col_3_15, 
      wind_col_in_3_14=>image_wind_col_3_14, wind_col_in_3_13=>
      image_wind_col_3_13, wind_col_in_3_12=>image_wind_col_3_12, 
      wind_col_in_3_11=>image_wind_col_3_11, wind_col_in_3_10=>
      image_wind_col_3_10, wind_col_in_3_9=>image_wind_col_3_9, 
      wind_col_in_3_8=>image_wind_col_3_8, wind_col_in_3_7=>
      image_wind_col_3_7, wind_col_in_3_6=>image_wind_col_3_6, 
      wind_col_in_3_5=>image_wind_col_3_5, wind_col_in_3_4=>
      image_wind_col_3_4, wind_col_in_3_3=>image_wind_col_3_3, 
      wind_col_in_3_2=>image_wind_col_3_2, wind_col_in_3_1=>
      image_wind_col_3_1, wind_col_in_3_0=>image_wind_col_3_0, 
      wind_col_in_2_15=>image_wind_col_2_15, wind_col_in_2_14=>
      image_wind_col_2_14, wind_col_in_2_13=>image_wind_col_2_13, 
      wind_col_in_2_12=>image_wind_col_2_12, wind_col_in_2_11=>
      image_wind_col_2_11, wind_col_in_2_10=>image_wind_col_2_10, 
      wind_col_in_2_9=>image_wind_col_2_9, wind_col_in_2_8=>
      image_wind_col_2_8, wind_col_in_2_7=>image_wind_col_2_7, 
      wind_col_in_2_6=>image_wind_col_2_6, wind_col_in_2_5=>
      image_wind_col_2_5, wind_col_in_2_4=>image_wind_col_2_4, 
      wind_col_in_2_3=>image_wind_col_2_3, wind_col_in_2_2=>
      image_wind_col_2_2, wind_col_in_2_1=>image_wind_col_2_1, 
      wind_col_in_2_0=>image_wind_col_2_0, wind_col_in_1_15=>
      image_wind_col_1_15, wind_col_in_1_14=>image_wind_col_1_14, 
      wind_col_in_1_13=>image_wind_col_1_13, wind_col_in_1_12=>
      image_wind_col_1_12, wind_col_in_1_11=>image_wind_col_1_11, 
      wind_col_in_1_10=>image_wind_col_1_10, wind_col_in_1_9=>
      image_wind_col_1_9, wind_col_in_1_8=>image_wind_col_1_8, 
      wind_col_in_1_7=>image_wind_col_1_7, wind_col_in_1_6=>
      image_wind_col_1_6, wind_col_in_1_5=>image_wind_col_1_5, 
      wind_col_in_1_4=>image_wind_col_1_4, wind_col_in_1_3=>
      image_wind_col_1_3, wind_col_in_1_2=>image_wind_col_1_2, 
      wind_col_in_1_1=>image_wind_col_1_1, wind_col_in_1_0=>
      image_wind_col_1_0, wind_col_in_0_15=>image_wind_col_0_15, 
      wind_col_in_0_14=>image_wind_col_0_14, wind_col_in_0_13=>
      image_wind_col_0_13, wind_col_in_0_12=>image_wind_col_0_12, 
      wind_col_in_0_11=>image_wind_col_0_11, wind_col_in_0_10=>
      image_wind_col_0_10, wind_col_in_0_9=>image_wind_col_0_9, 
      wind_col_in_0_8=>image_wind_col_0_8, wind_col_in_0_7=>
      image_wind_col_0_7, wind_col_in_0_6=>image_wind_col_0_6, 
      wind_col_in_0_5=>image_wind_col_0_5, wind_col_in_0_4=>
      image_wind_col_0_4, wind_col_in_0_3=>image_wind_col_0_3, 
      wind_col_in_0_2=>image_wind_col_0_2, wind_col_in_0_1=>
      image_wind_col_0_1, wind_col_in_0_0=>image_wind_col_0_0, 
      filter_data_out(15)=>filter_window_data_15, filter_data_out(14)=>
      filter_window_data_14, filter_data_out(13)=>filter_window_data_13, 
      filter_data_out(12)=>filter_window_data_12, filter_data_out(11)=>
      filter_window_data_11, filter_data_out(10)=>filter_window_data_10, 
      filter_data_out(9)=>filter_window_data_9, filter_data_out(8)=>
      filter_window_data_8, filter_data_out(7)=>filter_window_data_7, 
      filter_data_out(6)=>filter_window_data_6, filter_data_out(5)=>
      filter_window_data_5, filter_data_out(4)=>filter_window_data_4, 
      filter_data_out(3)=>filter_window_data_3, filter_data_out(2)=>
      filter_window_data_2, filter_data_out(1)=>filter_window_data_1, 
      filter_data_out(0)=>filter_window_data_0, filter_ready_out=>
      filter_window_ready, filter_reset=>DANGLING(2), comp_unit_ready=>
      comp_unit_ready, comp_unit_operation=>comp_unit_operation, 
      comp_unit_flt_size=>comp_unit_flt_size, comp_unit_relu=>comp_unit_relu, 
      comp_unit_data1_out(15)=>controller_bias_1_15, comp_unit_data1_out(14)
      =>controller_bias_1_14, comp_unit_data1_out(13)=>controller_bias_1_13, 
      comp_unit_data1_out(12)=>controller_bias_1_12, comp_unit_data1_out(11)
      =>controller_bias_1_11, comp_unit_data1_out(10)=>controller_bias_1_10, 
      comp_unit_data1_out(9)=>controller_bias_1_9, comp_unit_data1_out(8)=>
      controller_bias_1_8, comp_unit_data1_out(7)=>controller_bias_1_7, 
      comp_unit_data1_out(6)=>controller_bias_1_6, comp_unit_data1_out(5)=>
      controller_bias_1_5, comp_unit_data1_out(4)=>controller_bias_1_4, 
      comp_unit_data1_out(3)=>controller_bias_1_3, comp_unit_data1_out(2)=>
      controller_bias_1_2, comp_unit_data1_out(1)=>controller_bias_1_1, 
      comp_unit_data1_out(0)=>controller_bias_1_0, comp_unit_data2_out(15)=>
      controller_bias_2_15, comp_unit_data2_out(14)=>controller_bias_2_14, 
      comp_unit_data2_out(13)=>controller_bias_2_13, comp_unit_data2_out(12)
      =>controller_bias_2_12, comp_unit_data2_out(11)=>controller_bias_2_11, 
      comp_unit_data2_out(10)=>controller_bias_2_10, comp_unit_data2_out(9)
      =>controller_bias_2_9, comp_unit_data2_out(8)=>controller_bias_2_8, 
      comp_unit_data2_out(7)=>controller_bias_2_7, comp_unit_data2_out(6)=>
      controller_bias_2_6, comp_unit_data2_out(5)=>controller_bias_2_5, 
      comp_unit_data2_out(4)=>controller_bias_2_4, comp_unit_data2_out(3)=>
      controller_bias_2_3, comp_unit_data2_out(2)=>controller_bias_2_2, 
      comp_unit_data2_out(1)=>controller_bias_2_1, comp_unit_data2_out(0)=>
      controller_bias_2_0, comp_unit_buffer_finished=>io_done_out_EXMPLR, 
      comp_unit_finished=>comp_unit_finished, comp_unit_data1_in(15)=>
      controller_result_1_15, comp_unit_data1_in(14)=>controller_result_1_14, 
      comp_unit_data1_in(13)=>controller_result_1_13, comp_unit_data1_in(12)
      =>controller_result_1_12, comp_unit_data1_in(11)=>
      controller_result_1_11, comp_unit_data1_in(10)=>controller_result_1_10, 
      comp_unit_data1_in(9)=>controller_result_1_9, comp_unit_data1_in(8)=>
      controller_result_1_8, comp_unit_data1_in(7)=>controller_result_1_7, 
      comp_unit_data1_in(6)=>controller_result_1_6, comp_unit_data1_in(5)=>
      controller_result_1_5, comp_unit_data1_in(4)=>controller_result_1_4, 
      comp_unit_data1_in(3)=>controller_result_1_3, comp_unit_data1_in(2)=>
      controller_result_1_2, comp_unit_data1_in(1)=>controller_result_1_1, 
      comp_unit_data1_in(0)=>controller_result_1_0, comp_unit_data2_in(15)=>
      controller_result_2_15, comp_unit_data2_in(14)=>controller_result_2_14, 
      comp_unit_data2_in(13)=>controller_result_2_13, comp_unit_data2_in(12)
      =>controller_result_2_12, comp_unit_data2_in(11)=>
      controller_result_2_11, comp_unit_data2_in(10)=>controller_result_2_10, 
      comp_unit_data2_in(9)=>controller_result_2_9, comp_unit_data2_in(8)=>
      controller_result_2_8, comp_unit_data2_in(7)=>controller_result_2_7, 
      comp_unit_data2_in(6)=>controller_result_2_6, comp_unit_data2_in(5)=>
      controller_result_2_5, comp_unit_data2_in(4)=>controller_result_2_4, 
      comp_unit_data2_in(3)=>controller_result_2_3, comp_unit_data2_in(2)=>
      controller_result_2_2, comp_unit_data2_in(1)=>controller_result_2_1, 
      comp_unit_data2_in(0)=>controller_result_2_0, argmax_ready=>
      argmax_ready, argmax_data_out(15)=>argmax_data_outof_controller_15, 
      argmax_data_out(14)=>argmax_data_outof_controller_14, 
      argmax_data_out(13)=>argmax_data_outof_controller_13, 
      argmax_data_out(12)=>argmax_data_outof_controller_12, 
      argmax_data_out(11)=>argmax_data_outof_controller_11, 
      argmax_data_out(10)=>argmax_data_outof_controller_10, 
      argmax_data_out(9)=>argmax_data_outof_controller_9, argmax_data_out(8)
      =>argmax_data_outof_controller_8, argmax_data_out(7)=>
      argmax_data_outof_controller_7, argmax_data_out(6)=>
      argmax_data_outof_controller_6, argmax_data_out(5)=>
      argmax_data_outof_controller_5, argmax_data_out(4)=>
      argmax_data_outof_controller_4, argmax_data_out(3)=>
      argmax_data_outof_controller_3, argmax_data_out(2)=>
      argmax_data_outof_controller_2, argmax_data_out(1)=>
      argmax_data_outof_controller_1, argmax_data_out(0)=>
      argmax_data_outof_controller_0, argmax_data_in(15)=>io_done_out_EXMPLR, 
      argmax_data_in(14)=>io_done_out_EXMPLR, argmax_data_in(13)=>
      io_done_out_EXMPLR, argmax_data_in(12)=>io_done_out_EXMPLR, 
      argmax_data_in(11)=>io_done_out_EXMPLR, argmax_data_in(10)=>
      io_done_out_EXMPLR, argmax_data_in(9)=>io_done_out_EXMPLR, 
      argmax_data_in(8)=>io_done_out_EXMPLR, argmax_data_in(7)=>
      io_done_out_EXMPLR, argmax_data_in(6)=>io_done_out_EXMPLR, 
      argmax_data_in(5)=>io_done_out_EXMPLR, argmax_data_in(4)=>
      io_done_out_EXMPLR, argmax_data_in(3)=>argmax_data_out_3, 
      argmax_data_in(2)=>argmax_data_out_2, argmax_data_in(1)=>
      argmax_data_out_1, argmax_data_in(0)=>argmax_data_out_0);
   computation_block_inst : ComputationBlock port map ( img_data_col_0(15)=>
      image_wind_col_0_15, img_data_col_0(14)=>image_wind_col_0_14, 
      img_data_col_0(13)=>image_wind_col_0_13, img_data_col_0(12)=>
      image_wind_col_0_12, img_data_col_0(11)=>image_wind_col_0_11, 
      img_data_col_0(10)=>image_wind_col_0_10, img_data_col_0(9)=>
      image_wind_col_0_9, img_data_col_0(8)=>image_wind_col_0_8, 
      img_data_col_0(7)=>image_wind_col_0_7, img_data_col_0(6)=>
      image_wind_col_0_6, img_data_col_0(5)=>image_wind_col_0_5, 
      img_data_col_0(4)=>image_wind_col_0_4, img_data_col_0(3)=>
      image_wind_col_0_3, img_data_col_0(2)=>image_wind_col_0_2, 
      img_data_col_0(1)=>image_wind_col_0_1, img_data_col_0(0)=>
      image_wind_col_0_0, img_data_col_1(15)=>image_wind_col_1_15, 
      img_data_col_1(14)=>image_wind_col_1_14, img_data_col_1(13)=>
      image_wind_col_1_13, img_data_col_1(12)=>image_wind_col_1_12, 
      img_data_col_1(11)=>image_wind_col_1_11, img_data_col_1(10)=>
      image_wind_col_1_10, img_data_col_1(9)=>image_wind_col_1_9, 
      img_data_col_1(8)=>image_wind_col_1_8, img_data_col_1(7)=>
      image_wind_col_1_7, img_data_col_1(6)=>image_wind_col_1_6, 
      img_data_col_1(5)=>image_wind_col_1_5, img_data_col_1(4)=>
      image_wind_col_1_4, img_data_col_1(3)=>image_wind_col_1_3, 
      img_data_col_1(2)=>image_wind_col_1_2, img_data_col_1(1)=>
      image_wind_col_1_1, img_data_col_1(0)=>image_wind_col_1_0, 
      img_data_col_2(15)=>image_wind_col_2_15, img_data_col_2(14)=>
      image_wind_col_2_14, img_data_col_2(13)=>image_wind_col_2_13, 
      img_data_col_2(12)=>image_wind_col_2_12, img_data_col_2(11)=>
      image_wind_col_2_11, img_data_col_2(10)=>image_wind_col_2_10, 
      img_data_col_2(9)=>image_wind_col_2_9, img_data_col_2(8)=>
      image_wind_col_2_8, img_data_col_2(7)=>image_wind_col_2_7, 
      img_data_col_2(6)=>image_wind_col_2_6, img_data_col_2(5)=>
      image_wind_col_2_5, img_data_col_2(4)=>image_wind_col_2_4, 
      img_data_col_2(3)=>image_wind_col_2_3, img_data_col_2(2)=>
      image_wind_col_2_2, img_data_col_2(1)=>image_wind_col_2_1, 
      img_data_col_2(0)=>image_wind_col_2_0, img_data_col_3(15)=>
      image_wind_col_3_15, img_data_col_3(14)=>image_wind_col_3_14, 
      img_data_col_3(13)=>image_wind_col_3_13, img_data_col_3(12)=>
      image_wind_col_3_12, img_data_col_3(11)=>image_wind_col_3_11, 
      img_data_col_3(10)=>image_wind_col_3_10, img_data_col_3(9)=>
      image_wind_col_3_9, img_data_col_3(8)=>image_wind_col_3_8, 
      img_data_col_3(7)=>image_wind_col_3_7, img_data_col_3(6)=>
      image_wind_col_3_6, img_data_col_3(5)=>image_wind_col_3_5, 
      img_data_col_3(4)=>image_wind_col_3_4, img_data_col_3(3)=>
      image_wind_col_3_3, img_data_col_3(2)=>image_wind_col_3_2, 
      img_data_col_3(1)=>image_wind_col_3_1, img_data_col_3(0)=>
      image_wind_col_3_0, img_data_col_4(15)=>image_wind_col_4_15, 
      img_data_col_4(14)=>image_wind_col_4_14, img_data_col_4(13)=>
      image_wind_col_4_13, img_data_col_4(12)=>image_wind_col_4_12, 
      img_data_col_4(11)=>image_wind_col_4_11, img_data_col_4(10)=>
      image_wind_col_4_10, img_data_col_4(9)=>image_wind_col_4_9, 
      img_data_col_4(8)=>image_wind_col_4_8, img_data_col_4(7)=>
      image_wind_col_4_7, img_data_col_4(6)=>image_wind_col_4_6, 
      img_data_col_4(5)=>image_wind_col_4_5, img_data_col_4(4)=>
      image_wind_col_4_4, img_data_col_4(3)=>image_wind_col_4_3, 
      img_data_col_4(2)=>image_wind_col_4_2, img_data_col_4(1)=>
      image_wind_col_4_1, img_data_col_4(0)=>image_wind_col_4_0, img_load=>
      image_wind_en, img_reset=>io_done_out_EXMPLR, filter_data_word(15)=>
      filter_window_data_15, filter_data_word(14)=>filter_window_data_14, 
      filter_data_word(13)=>filter_window_data_13, filter_data_word(12)=>
      filter_window_data_12, filter_data_word(11)=>filter_window_data_11, 
      filter_data_word(10)=>filter_window_data_10, filter_data_word(9)=>
      filter_window_data_9, filter_data_word(8)=>filter_window_data_8, 
      filter_data_word(7)=>filter_window_data_7, filter_data_word(6)=>
      filter_window_data_6, filter_data_word(5)=>filter_window_data_5, 
      filter_data_word(4)=>filter_window_data_4, filter_data_word(3)=>
      filter_window_data_3, filter_data_word(2)=>filter_window_data_2, 
      filter_data_word(1)=>filter_window_data_1, filter_data_word(0)=>
      filter_window_data_0, filter_load=>filter_window_ready, filter_reset=>
      reset, start=>comp_unit_ready, operation=>comp_unit_operation, 
      compute_relu=>comp_unit_relu, filter_size=>comp_unit_flt_size, 
      output1_init(15)=>comp_unit_bias_1_15, output1_init(14)=>
      comp_unit_bias_1_14, output1_init(13)=>comp_unit_bias_1_13, 
      output1_init(12)=>comp_unit_bias_1_12, output1_init(11)=>
      comp_unit_bias_1_11, output1_init(10)=>comp_unit_bias_1_10, 
      output1_init(9)=>comp_unit_bias_1_9, output1_init(8)=>
      comp_unit_bias_1_8, output1_init(7)=>comp_unit_bias_1_7, 
      output1_init(6)=>comp_unit_bias_1_6, output1_init(5)=>
      comp_unit_bias_1_5, output1_init(4)=>comp_unit_bias_1_4, 
      output1_init(3)=>comp_unit_bias_1_3, output1_init(2)=>
      comp_unit_bias_1_2, output1_init(1)=>comp_unit_bias_1_1, 
      output1_init(0)=>comp_unit_bias_1_0, output2_init(15)=>
      comp_unit_bias_2_15, output2_init(14)=>comp_unit_bias_2_14, 
      output2_init(13)=>comp_unit_bias_2_13, output2_init(12)=>
      comp_unit_bias_2_12, output2_init(11)=>comp_unit_bias_2_11, 
      output2_init(10)=>comp_unit_bias_2_10, output2_init(9)=>
      comp_unit_bias_2_9, output2_init(8)=>comp_unit_bias_2_8, 
      output2_init(7)=>comp_unit_bias_2_7, output2_init(6)=>
      comp_unit_bias_2_6, output2_init(5)=>comp_unit_bias_2_5, 
      output2_init(4)=>comp_unit_bias_2_4, output2_init(3)=>
      comp_unit_bias_2_3, output2_init(2)=>comp_unit_bias_2_2, 
      output2_init(1)=>comp_unit_bias_2_1, output2_init(0)=>
      comp_unit_bias_2_0, output1(15)=>comp_unit_result_1_15, output1(14)=>
      comp_unit_result_1_14, output1(13)=>comp_unit_result_1_13, output1(12)
      =>comp_unit_result_1_12, output1(11)=>comp_unit_result_1_11, 
      output1(10)=>comp_unit_result_1_10, output1(9)=>comp_unit_result_1_9, 
      output1(8)=>comp_unit_result_1_8, output1(7)=>comp_unit_result_1_7, 
      output1(6)=>comp_unit_result_1_6, output1(5)=>comp_unit_result_1_5, 
      output1(4)=>comp_unit_result_1_4, output1(3)=>comp_unit_result_1_3, 
      output1(2)=>comp_unit_result_1_2, output1(1)=>comp_unit_result_1_1, 
      output1(0)=>comp_unit_result_1_0, output2(15)=>comp_unit_result_2_15, 
      output2(14)=>comp_unit_result_2_14, output2(13)=>comp_unit_result_2_13, 
      output2(12)=>comp_unit_result_2_12, output2(11)=>comp_unit_result_2_11, 
      output2(10)=>comp_unit_result_2_10, output2(9)=>comp_unit_result_2_9, 
      output2(8)=>comp_unit_result_2_8, output2(7)=>comp_unit_result_2_7, 
      output2(6)=>comp_unit_result_2_6, output2(5)=>comp_unit_result_2_5, 
      output2(4)=>comp_unit_result_2_4, output2(3)=>comp_unit_result_2_3, 
      output2(2)=>comp_unit_result_2_2, output2(1)=>comp_unit_result_2_1, 
      output2(0)=>comp_unit_result_2_0, buffer_ready=>DANGLING(3), ready=>
      comp_unit_finished, clk=>clk, en=>PWR, reset=>io_done_out_EXMPLR);
   argmax_inst : ArgMax port map ( inp(15)=>argmax_data_outof_controller_15, 
      inp(14)=>argmax_data_outof_controller_14, inp(13)=>
      argmax_data_outof_controller_13, inp(12)=>
      argmax_data_outof_controller_12, inp(11)=>
      argmax_data_outof_controller_11, inp(10)=>
      argmax_data_outof_controller_10, inp(9)=>
      argmax_data_outof_controller_9, inp(8)=>argmax_data_outof_controller_8, 
      inp(7)=>argmax_data_outof_controller_7, inp(6)=>
      argmax_data_outof_controller_6, inp(5)=>argmax_data_outof_controller_5, 
      inp(4)=>argmax_data_outof_controller_4, inp(3)=>
      argmax_data_outof_controller_3, inp(2)=>argmax_data_outof_controller_2, 
      inp(1)=>argmax_data_outof_controller_1, inp(0)=>
      argmax_data_outof_controller_0, en=>argmax_ready, clk=>clk, rst=>reset, 
      ans(3)=>argmax_data_out_3, ans(2)=>argmax_data_out_2, ans(1)=>
      argmax_data_out_1, ans(0)=>argmax_data_out_0);
   ix415 : fake_vcc port map ( Y=>PWR);
   ix413 : fake_gnd port map ( Y=>io_done_out_EXMPLR);
   flt_size_reg_reg_q_0 : dffr port map ( Q=>flt_size_out_0, QB=>OPEN, D=>
      nx495, CLK=>clk, R=>reset);
   ix496 : mux21_ni port map ( Y=>nx495, A0=>nx584, A1=>comp_unit_flt_size, 
      S0=>comp_unit_ready);
   ix583 : inv02 port map ( Y=>nx584, A=>nx612);
   ix11 : mux21_ni port map ( Y=>controller_result_2_0, A0=>
      comp_unit_result_1_0, A1=>comp_unit_result_2_0, S0=>nx612);
   ix19 : mux21_ni port map ( Y=>controller_result_2_1, A0=>
      comp_unit_result_1_1, A1=>comp_unit_result_2_1, S0=>nx612);
   ix27 : mux21_ni port map ( Y=>controller_result_2_2, A0=>
      comp_unit_result_1_2, A1=>comp_unit_result_2_2, S0=>nx612);
   ix35 : mux21_ni port map ( Y=>controller_result_2_3, A0=>
      comp_unit_result_1_3, A1=>comp_unit_result_2_3, S0=>nx612);
   ix43 : mux21_ni port map ( Y=>controller_result_2_4, A0=>
      comp_unit_result_1_4, A1=>comp_unit_result_2_4, S0=>nx612);
   ix51 : mux21_ni port map ( Y=>controller_result_2_5, A0=>
      comp_unit_result_1_5, A1=>comp_unit_result_2_5, S0=>nx612);
   ix59 : mux21_ni port map ( Y=>controller_result_2_6, A0=>
      comp_unit_result_1_6, A1=>comp_unit_result_2_6, S0=>nx614);
   ix67 : mux21_ni port map ( Y=>controller_result_2_7, A0=>
      comp_unit_result_1_7, A1=>comp_unit_result_2_7, S0=>nx614);
   ix75 : mux21_ni port map ( Y=>controller_result_2_8, A0=>
      comp_unit_result_1_8, A1=>comp_unit_result_2_8, S0=>nx614);
   ix83 : mux21_ni port map ( Y=>controller_result_2_9, A0=>
      comp_unit_result_1_9, A1=>comp_unit_result_2_9, S0=>nx614);
   ix91 : mux21_ni port map ( Y=>controller_result_2_10, A0=>
      comp_unit_result_1_10, A1=>comp_unit_result_2_10, S0=>nx614);
   ix99 : mux21_ni port map ( Y=>controller_result_2_11, A0=>
      comp_unit_result_1_11, A1=>comp_unit_result_2_11, S0=>nx614);
   ix107 : mux21_ni port map ( Y=>controller_result_2_12, A0=>
      comp_unit_result_1_12, A1=>comp_unit_result_2_12, S0=>nx614);
   ix115 : mux21_ni port map ( Y=>controller_result_2_13, A0=>
      comp_unit_result_1_13, A1=>comp_unit_result_2_13, S0=>nx616);
   ix123 : mux21_ni port map ( Y=>controller_result_2_14, A0=>
      comp_unit_result_1_14, A1=>comp_unit_result_2_14, S0=>nx616);
   ix131 : mux21_ni port map ( Y=>controller_result_2_15, A0=>
      comp_unit_result_1_15, A1=>comp_unit_result_2_15, S0=>nx616);
   ix139 : mux21_ni port map ( Y=>controller_result_1_0, A0=>
      comp_unit_result_2_0, A1=>comp_unit_result_1_0, S0=>nx616);
   ix147 : mux21_ni port map ( Y=>controller_result_1_1, A0=>
      comp_unit_result_2_1, A1=>comp_unit_result_1_1, S0=>nx616);
   ix155 : mux21_ni port map ( Y=>controller_result_1_2, A0=>
      comp_unit_result_2_2, A1=>comp_unit_result_1_2, S0=>nx616);
   ix163 : mux21_ni port map ( Y=>controller_result_1_3, A0=>
      comp_unit_result_2_3, A1=>comp_unit_result_1_3, S0=>nx616);
   ix171 : mux21_ni port map ( Y=>controller_result_1_4, A0=>
      comp_unit_result_2_4, A1=>comp_unit_result_1_4, S0=>nx618);
   ix179 : mux21_ni port map ( Y=>controller_result_1_5, A0=>
      comp_unit_result_2_5, A1=>comp_unit_result_1_5, S0=>nx618);
   ix187 : mux21_ni port map ( Y=>controller_result_1_6, A0=>
      comp_unit_result_2_6, A1=>comp_unit_result_1_6, S0=>nx618);
   ix195 : mux21_ni port map ( Y=>controller_result_1_7, A0=>
      comp_unit_result_2_7, A1=>comp_unit_result_1_7, S0=>nx618);
   ix203 : mux21_ni port map ( Y=>controller_result_1_8, A0=>
      comp_unit_result_2_8, A1=>comp_unit_result_1_8, S0=>nx618);
   ix211 : mux21_ni port map ( Y=>controller_result_1_9, A0=>
      comp_unit_result_2_9, A1=>comp_unit_result_1_9, S0=>nx618);
   ix219 : mux21_ni port map ( Y=>controller_result_1_10, A0=>
      comp_unit_result_2_10, A1=>comp_unit_result_1_10, S0=>nx618);
   ix227 : mux21_ni port map ( Y=>controller_result_1_11, A0=>
      comp_unit_result_2_11, A1=>comp_unit_result_1_11, S0=>nx620);
   ix235 : mux21_ni port map ( Y=>controller_result_1_12, A0=>
      comp_unit_result_2_12, A1=>comp_unit_result_1_12, S0=>nx620);
   ix243 : mux21_ni port map ( Y=>controller_result_1_13, A0=>
      comp_unit_result_2_13, A1=>comp_unit_result_1_13, S0=>nx620);
   ix251 : mux21_ni port map ( Y=>controller_result_1_14, A0=>
      comp_unit_result_2_14, A1=>comp_unit_result_1_14, S0=>nx620);
   ix259 : mux21_ni port map ( Y=>controller_result_1_15, A0=>
      comp_unit_result_2_15, A1=>comp_unit_result_1_15, S0=>nx620);
   ix269 : mux21_ni port map ( Y=>comp_unit_bias_2_0, A0=>
      controller_bias_2_0, A1=>controller_bias_1_0, S0=>nx624);
   ix545 : nand02 port map ( Y=>nx594, A0=>nx620, A1=>nx610);
   ix609 : inv01 port map ( Y=>nx610, A=>comp_unit_flt_size);
   ix277 : mux21_ni port map ( Y=>comp_unit_bias_2_1, A0=>
      controller_bias_2_1, A1=>controller_bias_1_1, S0=>nx624);
   ix285 : mux21_ni port map ( Y=>comp_unit_bias_2_2, A0=>
      controller_bias_2_2, A1=>controller_bias_1_2, S0=>nx624);
   ix293 : mux21_ni port map ( Y=>comp_unit_bias_2_3, A0=>
      controller_bias_2_3, A1=>controller_bias_1_3, S0=>nx624);
   ix301 : mux21_ni port map ( Y=>comp_unit_bias_2_4, A0=>
      controller_bias_2_4, A1=>controller_bias_1_4, S0=>nx624);
   ix309 : mux21_ni port map ( Y=>comp_unit_bias_2_5, A0=>
      controller_bias_2_5, A1=>controller_bias_1_5, S0=>nx624);
   ix317 : mux21_ni port map ( Y=>comp_unit_bias_2_6, A0=>
      controller_bias_2_6, A1=>controller_bias_1_6, S0=>nx624);
   ix325 : mux21_ni port map ( Y=>comp_unit_bias_2_7, A0=>
      controller_bias_2_7, A1=>controller_bias_1_7, S0=>nx626);
   ix333 : mux21_ni port map ( Y=>comp_unit_bias_2_8, A0=>
      controller_bias_2_8, A1=>controller_bias_1_8, S0=>nx626);
   ix341 : mux21_ni port map ( Y=>comp_unit_bias_2_9, A0=>
      controller_bias_2_9, A1=>controller_bias_1_9, S0=>nx626);
   ix349 : mux21_ni port map ( Y=>comp_unit_bias_2_10, A0=>
      controller_bias_2_10, A1=>controller_bias_1_10, S0=>nx626);
   ix357 : mux21_ni port map ( Y=>comp_unit_bias_2_11, A0=>
      controller_bias_2_11, A1=>controller_bias_1_11, S0=>nx626);
   ix365 : mux21_ni port map ( Y=>comp_unit_bias_2_12, A0=>
      controller_bias_2_12, A1=>controller_bias_1_12, S0=>nx626);
   ix373 : mux21_ni port map ( Y=>comp_unit_bias_2_13, A0=>
      controller_bias_2_13, A1=>controller_bias_1_13, S0=>nx626);
   ix381 : mux21_ni port map ( Y=>comp_unit_bias_2_14, A0=>
      controller_bias_2_14, A1=>controller_bias_1_14, S0=>nx628);
   ix389 : mux21_ni port map ( Y=>comp_unit_bias_2_15, A0=>
      controller_bias_2_15, A1=>controller_bias_1_15, S0=>nx628);
   ix397 : mux21_ni port map ( Y=>comp_unit_bias_1_0, A0=>
      controller_bias_1_0, A1=>controller_bias_2_0, S0=>nx628);
   ix405 : mux21_ni port map ( Y=>comp_unit_bias_1_1, A0=>
      controller_bias_1_1, A1=>controller_bias_2_1, S0=>nx628);
   ix417 : mux21_ni port map ( Y=>comp_unit_bias_1_2, A0=>
      controller_bias_1_2, A1=>controller_bias_2_2, S0=>nx628);
   ix421 : mux21_ni port map ( Y=>comp_unit_bias_1_3, A0=>
      controller_bias_1_3, A1=>controller_bias_2_3, S0=>nx628);
   ix429 : mux21_ni port map ( Y=>comp_unit_bias_1_4, A0=>
      controller_bias_1_4, A1=>controller_bias_2_4, S0=>nx628);
   ix437 : mux21_ni port map ( Y=>comp_unit_bias_1_5, A0=>
      controller_bias_1_5, A1=>controller_bias_2_5, S0=>nx630);
   ix445 : mux21_ni port map ( Y=>comp_unit_bias_1_6, A0=>
      controller_bias_1_6, A1=>controller_bias_2_6, S0=>nx630);
   ix453 : mux21_ni port map ( Y=>comp_unit_bias_1_7, A0=>
      controller_bias_1_7, A1=>controller_bias_2_7, S0=>nx630);
   ix461 : mux21_ni port map ( Y=>comp_unit_bias_1_8, A0=>
      controller_bias_1_8, A1=>controller_bias_2_8, S0=>nx630);
   ix469 : mux21_ni port map ( Y=>comp_unit_bias_1_9, A0=>
      controller_bias_1_9, A1=>controller_bias_2_9, S0=>nx630);
   ix477 : mux21_ni port map ( Y=>comp_unit_bias_1_10, A0=>
      controller_bias_1_10, A1=>controller_bias_2_10, S0=>nx630);
   ix485 : mux21_ni port map ( Y=>comp_unit_bias_1_11, A0=>
      controller_bias_1_11, A1=>controller_bias_2_11, S0=>nx630);
   ix493 : mux21_ni port map ( Y=>comp_unit_bias_1_12, A0=>
      controller_bias_1_12, A1=>controller_bias_2_12, S0=>nx632);
   ix501 : mux21_ni port map ( Y=>comp_unit_bias_1_13, A0=>
      controller_bias_1_13, A1=>controller_bias_2_13, S0=>nx632);
   ix509 : mux21_ni port map ( Y=>comp_unit_bias_1_14, A0=>
      controller_bias_1_14, A1=>controller_bias_2_14, S0=>nx632);
   ix517 : mux21_ni port map ( Y=>comp_unit_bias_1_15, A0=>
      controller_bias_1_15, A1=>controller_bias_2_15, S0=>nx632);
   ix611 : inv02 port map ( Y=>nx612, A=>flt_size_out_0);
   ix613 : inv02 port map ( Y=>nx614, A=>flt_size_out_0);
   ix615 : inv02 port map ( Y=>nx616, A=>flt_size_out_0);
   ix617 : inv02 port map ( Y=>nx618, A=>flt_size_out_0);
   ix619 : inv02 port map ( Y=>nx620, A=>flt_size_out_0);
   ix621 : inv01 port map ( Y=>nx622, A=>nx594);
   ix623 : inv02 port map ( Y=>nx624, A=>nx622);
   ix625 : inv02 port map ( Y=>nx626, A=>nx622);
   ix627 : inv02 port map ( Y=>nx628, A=>nx622);
   ix629 : inv02 port map ( Y=>nx630, A=>nx622);
   ix631 : inv02 port map ( Y=>nx632, A=>nx622);
end Structural ;

