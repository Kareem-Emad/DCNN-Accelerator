//
// Verilog description for cell Controller, 
// Sat May 11 13:08:18 2019
//
// LeonardoSpectrum Level 3, 2018a.2 
//


module Controller ( clk, reset, io_ready_in, io_done_out, mem_data_in, 
                    mem_data_out, mem_addr_out, mem_write_out, mem_read_out, 
                    wind_en, wind_rst, wind_col_in_4__15, wind_col_in_4__14, 
                    wind_col_in_4__13, wind_col_in_4__12, wind_col_in_4__11, 
                    wind_col_in_4__10, wind_col_in_4__9, wind_col_in_4__8, 
                    wind_col_in_4__7, wind_col_in_4__6, wind_col_in_4__5, 
                    wind_col_in_4__4, wind_col_in_4__3, wind_col_in_4__2, 
                    wind_col_in_4__1, wind_col_in_4__0, wind_col_in_3__15, 
                    wind_col_in_3__14, wind_col_in_3__13, wind_col_in_3__12, 
                    wind_col_in_3__11, wind_col_in_3__10, wind_col_in_3__9, 
                    wind_col_in_3__8, wind_col_in_3__7, wind_col_in_3__6, 
                    wind_col_in_3__5, wind_col_in_3__4, wind_col_in_3__3, 
                    wind_col_in_3__2, wind_col_in_3__1, wind_col_in_3__0, 
                    wind_col_in_2__15, wind_col_in_2__14, wind_col_in_2__13, 
                    wind_col_in_2__12, wind_col_in_2__11, wind_col_in_2__10, 
                    wind_col_in_2__9, wind_col_in_2__8, wind_col_in_2__7, 
                    wind_col_in_2__6, wind_col_in_2__5, wind_col_in_2__4, 
                    wind_col_in_2__3, wind_col_in_2__2, wind_col_in_2__1, 
                    wind_col_in_2__0, wind_col_in_1__15, wind_col_in_1__14, 
                    wind_col_in_1__13, wind_col_in_1__12, wind_col_in_1__11, 
                    wind_col_in_1__10, wind_col_in_1__9, wind_col_in_1__8, 
                    wind_col_in_1__7, wind_col_in_1__6, wind_col_in_1__5, 
                    wind_col_in_1__4, wind_col_in_1__3, wind_col_in_1__2, 
                    wind_col_in_1__1, wind_col_in_1__0, wind_col_in_0__15, 
                    wind_col_in_0__14, wind_col_in_0__13, wind_col_in_0__12, 
                    wind_col_in_0__11, wind_col_in_0__10, wind_col_in_0__9, 
                    wind_col_in_0__8, wind_col_in_0__7, wind_col_in_0__6, 
                    wind_col_in_0__5, wind_col_in_0__4, wind_col_in_0__3, 
                    wind_col_in_0__2, wind_col_in_0__1, wind_col_in_0__0, 
                    filter_data_out, filter_ready_out, filter_reset, 
                    comp_unit_ready, comp_unit_operation, comp_unit_flt_size, 
                    comp_unit_relu, comp_unit_data1_out, comp_unit_data2_out, 
                    comp_unit_buffer_finished, comp_unit_finished, 
                    comp_unit_data1_in, comp_unit_data2_in, argmax_ready, 
                    argmax_data_out, argmax_data_in ) ;

    input clk ;
    input reset ;
    input io_ready_in ;
    output io_done_out ;
    input [15:0]mem_data_in ;
    output [15:0]mem_data_out ;
    output [15:0]mem_addr_out ;
    output mem_write_out ;
    output mem_read_out ;
    output wind_en ;
    output wind_rst ;
    output wind_col_in_4__15 ;
    output wind_col_in_4__14 ;
    output wind_col_in_4__13 ;
    output wind_col_in_4__12 ;
    output wind_col_in_4__11 ;
    output wind_col_in_4__10 ;
    output wind_col_in_4__9 ;
    output wind_col_in_4__8 ;
    output wind_col_in_4__7 ;
    output wind_col_in_4__6 ;
    output wind_col_in_4__5 ;
    output wind_col_in_4__4 ;
    output wind_col_in_4__3 ;
    output wind_col_in_4__2 ;
    output wind_col_in_4__1 ;
    output wind_col_in_4__0 ;
    output wind_col_in_3__15 ;
    output wind_col_in_3__14 ;
    output wind_col_in_3__13 ;
    output wind_col_in_3__12 ;
    output wind_col_in_3__11 ;
    output wind_col_in_3__10 ;
    output wind_col_in_3__9 ;
    output wind_col_in_3__8 ;
    output wind_col_in_3__7 ;
    output wind_col_in_3__6 ;
    output wind_col_in_3__5 ;
    output wind_col_in_3__4 ;
    output wind_col_in_3__3 ;
    output wind_col_in_3__2 ;
    output wind_col_in_3__1 ;
    output wind_col_in_3__0 ;
    output wind_col_in_2__15 ;
    output wind_col_in_2__14 ;
    output wind_col_in_2__13 ;
    output wind_col_in_2__12 ;
    output wind_col_in_2__11 ;
    output wind_col_in_2__10 ;
    output wind_col_in_2__9 ;
    output wind_col_in_2__8 ;
    output wind_col_in_2__7 ;
    output wind_col_in_2__6 ;
    output wind_col_in_2__5 ;
    output wind_col_in_2__4 ;
    output wind_col_in_2__3 ;
    output wind_col_in_2__2 ;
    output wind_col_in_2__1 ;
    output wind_col_in_2__0 ;
    output wind_col_in_1__15 ;
    output wind_col_in_1__14 ;
    output wind_col_in_1__13 ;
    output wind_col_in_1__12 ;
    output wind_col_in_1__11 ;
    output wind_col_in_1__10 ;
    output wind_col_in_1__9 ;
    output wind_col_in_1__8 ;
    output wind_col_in_1__7 ;
    output wind_col_in_1__6 ;
    output wind_col_in_1__5 ;
    output wind_col_in_1__4 ;
    output wind_col_in_1__3 ;
    output wind_col_in_1__2 ;
    output wind_col_in_1__1 ;
    output wind_col_in_1__0 ;
    output wind_col_in_0__15 ;
    output wind_col_in_0__14 ;
    output wind_col_in_0__13 ;
    output wind_col_in_0__12 ;
    output wind_col_in_0__11 ;
    output wind_col_in_0__10 ;
    output wind_col_in_0__9 ;
    output wind_col_in_0__8 ;
    output wind_col_in_0__7 ;
    output wind_col_in_0__6 ;
    output wind_col_in_0__5 ;
    output wind_col_in_0__4 ;
    output wind_col_in_0__3 ;
    output wind_col_in_0__2 ;
    output wind_col_in_0__1 ;
    output wind_col_in_0__0 ;
    output [15:0]filter_data_out ;
    output filter_ready_out ;
    output filter_reset ;
    output comp_unit_ready ;
    output comp_unit_operation ;
    output comp_unit_flt_size ;
    output comp_unit_relu ;
    output [15:0]comp_unit_data1_out ;
    output [15:0]comp_unit_data2_out ;
    input comp_unit_buffer_finished ;
    input comp_unit_finished ;
    input [15:0]comp_unit_data1_in ;
    input [15:0]comp_unit_data2_in ;
    output argmax_ready ;
    output [15:0]argmax_data_out ;
    input [15:0]argmax_data_in ;

    wire current_state_13, wind_width_count_4, wind_width_count_3, 
         wind_width_count_2, wind_width_count_1, wind_width_count_0, 
         cache_height_count_en, cache_height_ended, max_height_2, max_height_0, 
         cache_width_count_4, cache_width_count_3, cache_width_count_2, 
         cache_width_count_1, cache_width_count_0, cache_data_in_15, 
         cache_data_in_14, cache_data_in_13, cache_data_in_12, cache_data_in_11, 
         cache_data_in_10, cache_data_in_9, cache_data_in_8, cache_data_in_7, 
         cache_data_in_6, cache_data_in_5, cache_data_in_4, cache_data_in_3, 
         cache_data_in_2, cache_data_in_1, cache_data_in_0, cache_data_out_4__15, 
         cache_data_out_4__14, cache_data_out_4__13, cache_data_out_4__12, 
         cache_data_out_4__11, cache_data_out_4__10, cache_data_out_4__9, 
         cache_data_out_4__8, cache_data_out_4__7, cache_data_out_4__6, 
         cache_data_out_4__5, cache_data_out_4__4, cache_data_out_4__3, 
         cache_data_out_4__2, cache_data_out_4__1, cache_data_out_4__0, 
         cache_data_out_3__15, cache_data_out_3__14, cache_data_out_3__13, 
         cache_data_out_3__12, cache_data_out_3__11, cache_data_out_3__10, 
         cache_data_out_3__9, cache_data_out_3__8, cache_data_out_3__7, 
         cache_data_out_3__6, cache_data_out_3__5, cache_data_out_3__4, 
         cache_data_out_3__3, cache_data_out_3__2, cache_data_out_3__1, 
         cache_data_out_3__0, cache_data_out_2__15, cache_data_out_2__14, 
         cache_data_out_2__13, cache_data_out_2__12, cache_data_out_2__11, 
         cache_data_out_2__10, cache_data_out_2__9, cache_data_out_2__8, 
         cache_data_out_2__7, cache_data_out_2__6, cache_data_out_2__5, 
         cache_data_out_2__4, cache_data_out_2__3, cache_data_out_2__2, 
         cache_data_out_2__1, cache_data_out_2__0, cache_data_out_1__15, 
         cache_data_out_1__14, cache_data_out_1__13, cache_data_out_1__12, 
         cache_data_out_1__11, cache_data_out_1__10, cache_data_out_1__9, 
         cache_data_out_1__8, cache_data_out_1__7, cache_data_out_1__6, 
         cache_data_out_1__5, cache_data_out_1__4, cache_data_out_1__3, 
         cache_data_out_1__2, cache_data_out_1__1, cache_data_out_1__0, 
         cache_data_out_0__15, cache_data_out_0__14, cache_data_out_0__13, 
         cache_data_out_0__12, cache_data_out_0__11, cache_data_out_0__10, 
         cache_data_out_0__9, cache_data_out_0__8, cache_data_out_0__7, 
         cache_data_out_0__6, cache_data_out_0__5, cache_data_out_0__4, 
         cache_data_out_0__3, cache_data_out_0__2, cache_data_out_0__1, 
         cache_data_out_0__0, cache_load, cache_rst_actual, max_height_4, 
         max_height_3, max_height_1, current_state_21, layer_type_out_1, 
         current_state_3, current_state_26, nflt_layer_out_3, current_state_4, 
         nflt_layer_out_1, nflt_layer_out_0, nx78, nx12873, nx92, 
         current_state_8, current_state_7, current_state_6, current_state_5, 
         nx118, current_state_2, nx134, nx140, nx148, nx12875, current_state_24, 
         ftc_cntrl_reg_out_12, current_state_16, ftc_cntrl_reg_out_8, nx12877, 
         nx158, ftc_cntrl_reg_out_14, current_state_10, nx174, nx182, nx196, 
         cntr1_inst_counter_out_1, cntr1_inst_counter_out_0, nx206, 
         cntr1_inst_counter_out_3, cntr1_inst_counter_out_2, nx230, nx244, 
         cntr1_inst_counter_out_4, nx12882, nx262, nx276, nx278, flt_size_out_0, 
         flt_size_out_2, flt_size_out_1, nx308, nx310, nx316, nx330, nx12883, 
         nx336, ftc_cntrl_reg_out_13, nx362, ftc_cntrl_reg_out_11, nx12884, 
         window_width_cntr_counter_out_14, nx12885, 
         window_width_cntr_counter_out_13, window_width_cntr_counter_out_12, 
         nx12887, window_width_cntr_counter_out_11, 
         window_width_cntr_counter_out_10, nx12889, 
         window_width_cntr_counter_out_9, window_width_cntr_counter_out_8, 
         nx12891, window_width_cntr_counter_out_7, 
         window_width_cntr_counter_out_6, nx12893, 
         window_width_cntr_counter_out_5, nx378, nx384, nx392, nx400, nx408, 
         nx428, nx452, nx476, nx500, nx524, nx550, nx564, nx576, img_width_out_0, 
         nx582, new_width_out_0, nx602, nx604, nx612, img_width_out_1, 
         new_width_out_1, nx630, nx636, nx640, img_width_out_2, new_width_out_2, 
         nx674, img_width_out_3, new_width_out_3, nx704, img_width_out_4, 
         new_width_out_4, nx722, nx732, current_state_15, 
         write_offset_data_out_0, nx760, new_size_squared_out_0, 
         write_offset_data_out_1, nx780, new_size_squared_out_1, 
         write_offset_data_out_2, new_size_squared_out_2, 
         write_offset_data_out_3, nx832, new_size_squared_out_3, nx850, 
         write_offset_data_out_4, nx852, nx858, new_size_squared_out_4, 
         write_offset_data_out_5, new_size_squared_out_5, 
         write_offset_data_out_6, nx898, nx904, new_size_squared_out_6, 
         write_offset_data_out_7, new_size_squared_out_7, nx944, 
         write_offset_data_out_8, nx948, nx954, new_size_squared_out_8, 
         write_offset_data_out_9, new_size_squared_out_9, 
         write_offset_data_out_10, nx994, nx1000, new_size_squared_out_10, 
         write_offset_data_out_11, new_size_squared_out_11, nx1040, 
         write_offset_data_out_12, nx1042, nx1048, new_size_squared_out_12, 
         write_offset_data_out_13, new_size_squared_out_13, 
         write_offset_data_out_14, nx1088, nx1094, new_size_squared_out_14, 
         write_offset_data_out_15, new_size_squared_out_15, nx1128, nx1138, 
         ftc_cntrl_reg_out_9, nx1146, nx1154, nx1168, ftc_cntrl_reg_out_10, 
         nx1182, nx1206, nx1212, cache_width_cntr_counter_out_14, nx12896, 
         cache_width_cntr_counter_out_13, cache_width_cntr_counter_out_12, 
         nx12898, cache_width_cntr_counter_out_11, 
         cache_width_cntr_counter_out_10, nx12900, 
         cache_width_cntr_counter_out_9, cache_width_cntr_counter_out_8, nx12902, 
         cache_width_cntr_counter_out_7, cache_width_cntr_counter_out_6, nx12904, 
         nx1224, nx1230, nx1238, nx1246, nx1254, cache_width_cntr_counter_out_5, 
         nx1260, nx1280, nx1304, nx1328, nx1352, nx1376, nx1402, nx1416, nx1434, 
         nx1436, nx1438, nx1446, nx1448, nx1456, nx1460, current_state_19, 
         current_state_18, nx1478, nx1484, nx1500, nx12906, nx1518, nx1524, 
         nx1534, nx1546, num_channels_counter_out_3, nflt_layer_temp_3, 
         num_channels_counter_out_2, nflt_layer_temp_2, nx12908, 
         num_channels_counter_out_1, nflt_layer_temp_1, 
         num_channels_counter_out_0, nflt_layer_temp_0, 
         max_num_channels_data_out_0, nx1608, nx1618, nx1642, nx1648, nx1660, 
         max_num_channels_data_out_2, nx1674, nx1686, 
         max_num_channels_data_out_3, nx1700, nx1712, 
         max_num_channels_data_out_4, nlayers_counter_out_0, nx12910, 
         nlayers_counter_out_2, nlayers_counter_out_1, nx1764, nx1780, nx1796, 
         nx12912, nx1838, nx1876, current_state_27, class_cntr_counter_out_3, 
         class_cntr_counter_out_2, class_cntr_counter_out_1, 
         class_cntr_counter_out_0, nx1904, nx1912, nx1926, nx1938, nx1946, 
         flt_bias_out_0, nx2128, nx2140, nx2142, flt_bias_out_1, nx2168, 
         flt_bias_out_2, nx2194, flt_bias_out_3, nx2220, flt_bias_out_4, nx2246, 
         flt_bias_out_5, nx2272, flt_bias_out_6, nx2298, flt_bias_out_7, nx2324, 
         flt_bias_out_8, nx2350, flt_bias_out_9, nx2376, flt_bias_out_10, nx2402, 
         flt_bias_out_11, nx2428, flt_bias_out_12, nx2454, flt_bias_out_13, 
         nx2480, flt_bias_out_14, nx2506, flt_bias_out_15, nx2532, nx2546, 
         ftc_cntrl_reg_out_15, nx2566, nx2580, nx2622, nx2642, 
         bias_offset_data_out_0, nx2664, nx2668, img_base_addr_0, 
         write_base_prev_data_out_0, nx2674, nx2678, img_addr_offset_0, nx2712, 
         nx2724, nx2738, nx2740, addr1_data_0, nx2754, nx2766, 
         write_base_data_out_1, addr1_data_1, nx2822, img_base_addr_1, 
         write_base_prev_data_out_1, img_addr_offset_1, bias_offset_data_out_1, 
         nx2874, nx2882, nx2892, write_base_data_out_2, nx2914, nx2924, nx2926, 
         nx2928, nx2932, addr1_data_2, nx2942, img_base_addr_2, 
         write_base_prev_data_out_2, nx2968, nx2974, img_addr_offset_2, nx2988, 
         nx2996, bias_offset_data_out_2, nx3016, write_base_data_out_3, nx3048, 
         nx3050, nx3060, nx3074, nx3076, nx3078, addr1_data_3, nx3092, 
         bias_offset_data_out_3, nx3122, img_base_addr_3, 
         write_base_prev_data_out_3, nx3146, img_addr_offset_3, nx3160, nx3168, 
         write_base_data_out_4, nx3206, addr1_data_4, nx3232, nx3238, nx3246, 
         img_base_addr_4, nx3264, nx3270, img_addr_offset_4, nx3278, nx3284, 
         nx3292, bias_offset_data_out_4, nx3312, write_base_data_out_5, nx3346, 
         nx3356, nx3360, nx3370, addr1_data_5, img_base_addr_5, 
         write_base_prev_data_out_5, nx3412, img_addr_offset_5, nx3434, 
         bias_offset_data_out_5, nx3454, nx3458, write_base_data_out_6, 
         addr1_data_6, nx3516, nx3522, nx3532, img_base_addr_6, nx3548, nx3554, 
         img_addr_offset_6, nx3562, nx3568, bias_offset_data_out_6, nx3608, 
         write_base_data_out_7, nx3630, nx3640, nx3654, addr1_data_7, 
         img_base_addr_7, write_base_prev_data_out_7, nx3696, img_addr_offset_7, 
         nx3718, bias_offset_data_out_7, nx3738, nx3742, write_base_data_out_8, 
         nx3780, addr1_data_8, nx3800, nx3806, nx3816, img_base_addr_8, nx3832, 
         nx3838, img_addr_offset_8, nx3846, nx3852, bias_offset_data_out_8, 
         nx3892, write_base_data_out_9, nx3914, nx3924, nx3938, addr1_data_9, 
         img_base_addr_9, write_base_prev_data_out_9, nx3980, img_addr_offset_9, 
         nx4002, bias_offset_data_out_9, nx4022, nx4026, nx4044, 
         write_base_data_out_10, addr1_data_10, nx4084, nx4090, nx4100, 
         img_base_addr_10, nx4116, nx4122, img_addr_offset_10, nx4130, nx4136, 
         bias_offset_data_out_10, nx4176, write_base_data_out_11, nx4198, nx4208, 
         nx4222, addr1_data_11, img_base_addr_11, write_base_prev_data_out_11, 
         nx4264, img_addr_offset_11, nx4286, bias_offset_data_out_11, nx4306, 
         write_base_data_out_12, addr1_data_12, nx4368, nx4374, img_base_addr_12, 
         nx4400, nx4406, img_addr_offset_12, nx4414, nx4420, 
         bias_offset_data_out_12, write_base_data_out_13, nx4492, nx4506, 
         addr1_data_13, nx4534, img_base_addr_13, write_base_prev_data_out_13, 
         nx4548, img_addr_offset_13, nx4568, nx4570, bias_offset_data_out_13, 
         nx4590, nx4594, write_base_data_out_14, addr1_data_14, nx4652, nx4658, 
         nx4668, img_base_addr_14, nx4684, nx4690, img_addr_offset_14, nx4698, 
         nx4704, bias_offset_data_out_14, nx4744, nx4754, 
         bias_offset_data_out_15, write_base_data_out_15, nx4782, addr1_data_15, 
         nx4802, nx4804, nx4812, nx4816, nx4826, img_base_addr_15, 
         write_base_prev_data_out_15, nx4834, nx4850, nx12921, nx12931, nx12941, 
         nx12951, nx12961, nx12971, nx12981, nx12991, nx13001, nx13011, nx13021, 
         nx13031, nx13041, nx13051, nx13061, nx13071, nx13081, nx13091, nx13101, 
         nx13111, nx13121, nx13131, nx13141, nx13151, nx13161, nx13171, nx13181, 
         nx13191, nx13201, nx13211, nx13221, nx13231, nx13241, nx13251, nx13261, 
         nx13271, nx13281, nx13291, nx13301, nx13311, nx13321, nx13331, nx13341, 
         nx13351, nx13361, nx13371, nx13381, nx13391, nx13401, nx13411, nx13421, 
         nx13431, nx13441, nx13451, nx13461, nx13471, nx13481, nx13491, nx13501, 
         nx13511, nx13521, nx13531, nx13541, nx13551, nx13561, nx13571, nx13581, 
         nx13591, nx13601, nx13611, nx13621, nx13631, nx13641, nx13651, nx13661, 
         nx13671, nx13681, nx13691, nx13701, nx13711, nx13721, nx13731, nx13741, 
         nx13751, nx13761, nx13771, nx13781, nx13791, nx13801, nx13811, nx13821, 
         nx13831, nx13841, nx13851, nx13861, nx13871, nx13881, nx13891, nx13901, 
         nx13911, nx13921, nx13931, nx13941, nx13951, nx13961, nx13971, nx13981, 
         nx13991, nx14001, nx14011, nx14021, nx14031, nx14041, nx14051, nx14061, 
         nx14071, nx14081, nx14091, nx14101, nx14111, nx14121, nx14131, nx14141, 
         nx14151, nx14161, nx14171, nx14181, nx14191, nx14201, nx14211, nx14221, 
         nx14231, nx14241, nx14251, nx14261, nx14271, nx14281, nx14291, nx14301, 
         nx14311, nx14321, nx14331, nx14341, nx14351, nx14361, nx14371, nx14381, 
         nx14391, nx14401, nx14411, nx14421, nx14431, nx14441, nx14451, nx14461, 
         nx14471, nx14481, nx14491, nx14501, nx14511, nx14521, nx14531, nx14541, 
         nx14551, nx14561, nx14571, nx14581, nx14591, nx14601, nx14611, nx14621, 
         nx14631, nx14641, nx14651, nx14661, nx14671, nx14681, nx14691, nx14701, 
         nx14711, nx14721, nx14731, nx14741, nx14751, nx14761, nx14771, nx14781, 
         nx14791, nx14801, nx14811, nx14821, nx14831, nx14841, nx14851, nx14861, 
         nx14871, nx14881, nx14891, nx14901, nx14911, nx14921, nx14931, nx14941, 
         nx14951, nx14961, nx14971, nx14981, nx14991, nx15001, nx15011, nx15021, 
         nx15031, nx15041, nx15051, nx15061, nx15071, nx15081, nx15091, nx15101, 
         nx15111, nx15121, nx15131, nx15141, nx15161, nx15171, nx15181, nx15191, 
         nx15201, nx15221, nx15231, nx15241, nx15251, nx15261, nx15281, nx15291, 
         nx15301, nx15311, nx15321, nx15331, nx15351, nx15361, nx15371, nx15381, 
         nx15392, nx15396, nx15402, nx15407, nx15412, nx15416, nx15422, nx15426, 
         nx15428, nx15432, nx15435, nx15445, nx15450, nx15452, nx15460, nx15466, 
         nx15470, nx15474, nx15479, nx15486, nx15488, nx15491, nx15496, nx15500, 
         nx15502, nx15504, nx15506, nx15508, nx15512, nx15514, nx15516, nx15518, 
         nx15523, nx15525, nx15527, nx15530, nx15531, nx15533, nx15537, nx15541, 
         nx15544, nx15546, nx15548, nx15554, nx15559, nx15561, nx15563, nx15567, 
         nx15571, nx15573, nx15575, nx15580, nx15586, nx15588, nx15591, nx15596, 
         nx15598, nx15602, nx15605, nx15609, nx15614, nx15617, nx15619, nx15621, 
         nx15626, nx15630, nx15635, nx15637, nx15640, nx15644, nx15647, nx15653, 
         nx15657, nx15660, nx15666, nx15670, nx15673, nx15679, nx15683, nx15686, 
         nx15692, nx15696, nx15711, nx15716, nx15717, nx15720, nx15726, nx15730, 
         nx15732, nx15735, nx15741, nx15745, nx15750, nx15753, nx15756, nx15759, 
         nx15763, nx15765, nx15768, nx15770, nx15772, nx15774, nx15776, nx15781, 
         nx15785, nx15786, nx15791, nx15795, nx15797, nx15802, nx15806, nx15807, 
         nx15812, nx15816, nx15818, nx15823, nx15827, nx15828, nx15833, nx15837, 
         nx15839, nx15844, nx15848, nx15849, nx15854, nx15859, nx15861, nx15865, 
         nx15868, nx15873, nx15876, nx15878, nx15883, nx15885, nx15888, nx15890, 
         nx15893, nx15898, nx15902, nx15904, nx15907, nx15912, nx15916, nx15918, 
         nx15921, nx15926, nx15930, nx15932, nx15935, nx15940, nx15944, nx15946, 
         nx15949, nx15954, nx15959, nx15970, nx15974, nx15983, nx15989, nx15995, 
         nx15997, nx16005, nx16013, nx16019, nx16025, nx16028, nx16037, nx16039, 
         nx16042, nx16046, nx16052, nx16055, nx16063, nx16065, nx16067, nx16070, 
         nx16075, nx16079, nx16081, nx16084, nx16089, nx16093, nx16095, nx16098, 
         nx16103, nx16107, nx16109, nx16112, nx16117, nx16121, nx16123, nx16126, 
         nx16131, nx16136, nx16148, nx16150, nx16153, nx16155, nx16166, nx16172, 
         nx16178, nx16180, nx16189, nx16191, nx16196, nx16198, nx16202, nx16204, 
         nx16213, nx16216, nx16222, nx16224, nx16226, nx16228, nx16234, nx16239, 
         nx16243, nx16247, nx16253, nx16258, nx16262, nx16265, nx16269, nx16274, 
         nx16278, nx16280, nx16282, nx16284, nx16290, nx16299, nx16302, nx16305, 
         nx16307, nx16313, nx16318, nx16324, nx16327, nx16332, nx16334, nx16336, 
         nx16338, nx16346, nx16348, nx16373, nx16455, nx16459, nx16463, nx16507, 
         nx16511, nx16514, nx16518, nx16521, nx16524, nx16527, nx16530, nx16533, 
         nx16536, nx16539, nx16542, nx16545, nx16548, nx16551, nx16554, nx16557, 
         nx16560, nx16563, nx16566, nx16569, nx16572, nx16575, nx16578, nx16581, 
         nx16584, nx16587, nx16590, nx16593, nx16596, nx16599, nx16602, nx16605, 
         nx16608, nx16610, nx16629, nx16715, nx16721, nx16727, nx16729, nx16732, 
         nx16736, nx16738, nx16742, nx16745, nx16747, nx16756, nx16764, nx16768, 
         nx16770, nx16774, nx16776, nx16780, nx16786, nx16788, nx16791, nx16796, 
         nx16798, nx16802, nx16804, nx16806, nx16810, nx16812, nx16818, nx16820, 
         nx16825, nx16829, nx16831, nx16833, nx16835, nx16837, nx16839, nx16843, 
         nx16846, nx16849, nx16852, nx16857, nx16861, nx16863, nx16868, nx16870, 
         nx16874, nx16878, nx16880, nx16895, nx16906, nx16911, nx16915, nx16916, 
         nx16924, nx16927, nx16931, nx16934, nx16943, nx16945, nx16948, nx16956, 
         nx16962, nx16967, nx16973, nx16976, nx16978, nx16983, nx16993, nx17002, 
         nx17004, nx17021, nx17031, nx17035, nx17038, nx17042, nx17044, nx17047, 
         nx17051, nx17054, nx17056, nx17060, nx17065, nx17074, nx17076, nx17077, 
         nx17081, nx17085, nx17089, nx17100, nx17102, nx17104, nx17106, nx17110, 
         nx17112, nx17114, nx17125, nx17135, nx17138, nx17140, nx17147, nx17157, 
         nx17161, nx17164, nx17168, nx17175, nx17178, nx17183, nx17186, nx17188, 
         nx17194, nx17199, nx17204, nx17210, nx17214, nx17218, nx17229, nx17231, 
         nx17233, nx17235, nx17239, nx17242, nx17244, nx17255, nx17265, nx17268, 
         nx17270, nx17277, nx17287, nx17291, nx17294, nx17298, nx17307, nx17310, 
         nx17312, nx17315, nx17321, nx17326, nx17331, nx17337, nx17341, nx17345, 
         nx17356, nx17358, nx17360, nx17362, nx17366, nx17369, nx17371, nx17374, 
         nx17377, nx17382, nx17392, nx17395, nx17397, nx17404, nx17414, nx17418, 
         nx17421, nx17425, nx17434, nx17437, nx17439, nx17442, nx17448, nx17453, 
         nx17458, nx17464, nx17468, nx17472, nx17483, nx17485, nx17487, nx17489, 
         nx17493, nx17496, nx17498, nx17509, nx17519, nx17522, nx17541, nx17545, 
         nx17548, nx17552, nx17561, nx17564, nx17566, nx17575, nx17580, nx17591, 
         nx17595, nx17599, nx17610, nx17612, nx17614, nx17616, nx17620, nx17623, 
         nx17625, nx17636, nx17641, nx17646, nx17649, nx17658, nx17660, nx17663, 
         nx17670, nx17671, nx17673, nx17677, nx17679, nx17682, nx17685, nx17687, 
         nx17692, nx17696, nx17700, nx17711, nx17723, nx17726, nx17728, nx17737, 
         nx17740, nx17744, nx17748, nx17751, nx17754, nx17757, nx17760, nx17763, 
         nx17766, nx17769, nx17772, nx17775, nx17778, nx17781, nx17784, nx17787, 
         nx17790, nx17793, nx17796, nx17803, nx17805, nx17807, nx17809, nx17811, 
         nx17813, nx17815, nx17817, nx17819, nx17821, nx17823, nx17825, nx17827, 
         nx17829, nx17831, nx17833, nx17835, nx17837, nx17839, nx17841, nx17843, 
         nx17845, nx17847, nx17855, nx17857, nx17859, nx17863, nx17865, nx17869, 
         nx17871, nx17873, nx17875, nx17877, nx17879, nx17887, nx17893, nx17895, 
         nx17897, nx17899, nx17907, nx17909, nx17911, nx17913, nx17915, nx17917, 
         nx17919, nx17921, nx17923, nx17927, nx17929, nx17937, nx17939, nx17941, 
         nx17943, nx17945, nx17947, nx17949, nx17951, nx17959, nx17961, nx17963, 
         nx17965, nx17971, nx17973, nx17975, nx17979, nx17981, nx17983, nx17993, 
         nx17995, nx17997, nx17999, nx18001, nx18003, nx18005, nx18007, nx18011, 
         nx18017, nx18021, nx18023, nx18027, nx18029, nx18031, nx18033, nx18035, 
         nx18037, nx18039, nx18041, nx18045, nx18047, nx18049, nx18051, nx18053, 
         nx18055, nx18059, nx18063, nx18065, nx18067, nx18069, nx18077, nx18081, 
         nx18085, nx18087, nx18089, nx18091, nx18117, nx18119, nx18121, nx18137, 
         nx18139, nx18141, nx18143, nx18151, nx18153, nx18155, nx18157, nx18163, 
         nx18165, nx18167, nx18169, nx18171, nx18173, nx18175, nx18177, nx18179, 
         nx18181, nx18183, nx18185, nx18187, nx18189, nx18191, nx18193, nx18195, 
         nx18197, nx18199, nx18201, nx18203, nx18205, nx18207, nx18211, nx18217, 
         nx18219, nx18225, nx18227, nx18229, nx18231, nx18233, nx18235, nx18237, 
         nx18239, nx18241, nx18243, nx18245, nx18247, nx18249, nx18251, nx18253, 
         nx18255, nx18257, nx18259, nx18261, nx18263, nx18265, nx18269, nx18271, 
         nx18273, nx18275, nx18277, nx18279, nx18281, nx18283, nx18285, nx18287, 
         nx18289, nx18291, nx18293, nx18295, nx18297, nx18299, nx18301, nx18303, 
         nx18305, nx18307, nx18309, nx18311, nx18313, nx18315, nx18317, nx18319, 
         nx18321, nx18323, nx18325, nx18327, nx18329, nx18331, nx18333, nx18335, 
         nx18339, nx18341, nx18343, nx18345, nx18347, nx18349, nx18351, nx18353, 
         nx18355, nx18357, nx18359, nx18361, nx18363, nx18365, nx18367, nx18369, 
         nx18371, nx18373, nx18375, nx18381, nx18383, nx18385, nx17067, nx3366, 
         nx16995, nx18543, nx18544, nx18545, nx18546, nx18547, nx18548, nx18549, 
         nx18550, nx18551, nx18552, nx18553, nx15341, nx18554, nx18555, nx18556, 
         nx18557, nx18558, nx18559, nx18560, nx18561, nx18562, nx18009, nx18563, 
         nx18564, nx18565, nx18566, nx18567, nx18568, nx3046, nx16882, nx16885, 
         nx16808, nx18569, nx18570, nx18571, nx18572, nx18573, nx18574, nx18575, 
         NOT_nx4768, nx18576, nx18577, nx18578, nx18579, nx16888, nx18580, 
         nx18581, nx18582, nx18583, nx18584, nx18585, nx3444, nx18586, nx18587, 
         nx17013, nx18588, nx17016, nx3112, nx16891, nx18589, nx18590, nx16987, 
         nx18591, nx18592, nx18593, nx18594, nx18595, nx18596, nx18597, nx18598, 
         nx18599, nx17118, nx18600, nx18601, nx17121, nx3184, nx18602, nx18603, 
         nx16990, nx18604, nx17656, nx18605, nx18223, nx18606, nx18607, nx18608, 
         nx18609, nx18610, nx18043, nx18611, nx18612, nx18613, nx18614, nx18615, 
         nx15271, nx18616, nx18617, nx18618, nx18619, nx18620, nx18621, nx18622, 
         nx18623, nx18624, nx18625, nx4612, nx18626, nx17731, nx18627, nx18628, 
         nx18629, nx17629, nx18630, nx18631, nx17632, nx4328, nx18632, nx17502, 
         nx17505, nx17529, nx18633, nx18634, nx18635, nx18636, nx15151, nx18267, 
         nx18337, nx18637, nx18638, nx18639, nx18640, nx18641, nx18642, nx18643, 
         nx18644, nx18645, nx18646, nx17023, nx18647, nx3132, nx18648, nx16898, 
         nx18649, nx16901, nx16814, nx18650, nx18651, nx18652, nx18653, nx18654, 
         nx18655, nx18656, nx18657, nx18658, nx17127, nx18659, nx18660, nx18661, 
         nx18662, nx18663, nx18664, nx18665, nx18666, nx18667, nx18668, nx18669, 
         nx18670, nx18671, nx18672, nx18673, nx15211, nx17585, nx18674, nx18675, 
         nx18676, nx18677, nx18678, nx17526, nx18679, nx18680, nx17402, nx18681, 
         nx18682, nx18683, nx18684, nx18685, nx18686, nx18687, nx18688, nx4194, 
         nx18689, nx18690, nx18691, nx18692, nx17399, nx18693, nx18694, nx18695, 
         nx18696, nx17272, nx18697, nx18698, nx17275, nx3626, nx18699, nx18700, 
         nx17145, nx18701, nx18702, nx18703, nx18704, nx18705, nx18706, nx18707, 
         nx18708, nx18709, nx18710, nx18711, nx4502, nx18712, nx18713, nx18714, 
         nx18715, nx18716, nx17556, nx4218, nx17429, nx4168, nx18717, nx18718, 
         nx18719, nx18720, nx18721, nx18722, nx18723, nx18724, nx17638, nx18725, 
         nx18726, nx18727, nx18728, nx18729, nx18730, nx17511, nx18731, nx17514, 
         nx4296, nx18732, nx18733, nx17384, nx17387, nx18734, nx18735, nx18736, 
         nx18737, nx18738, nx18739, nx18740, nx18741, nx18742, NOT_nx3476, 
         nx18743, nx18744, nx18745, nx18746, nx18747, nx18748, nx18749, nx18750, 
         nx3682, nx18751, nx18752, nx18753, nx18754, nx18755, nx18756, nx3966, 
         nx18757, nx18758, nx17279, nx18759, nx17282, nx18760, nx18761, nx18762, 
         nx17149, nx18763, nx17152, nx3398, nx17026, nx18764, nx18765, nx18766, 
         nx18767, nx18768, nx18769, nx3342, nx18770, nx18771, nx17006, nx18772, 
         nx18773, nx17009, nx18774, nx18775, nx18776, nx18777, nx18778, nx18779, 
         nx18780, nx4496, nx18781, nx17431, nx18782, nx18783, nx18784, nx18785, 
         nx18786, nx18787, nx18788, nx17323, nx18789, nx18790, nx3934, nx18791, 
         nx18792, nx3644, nx18793, nx18794, nx18795, nx17196, nx3884, nx3928, 
         nx17302, nx3650, nx17172, nx3600, nx18796, nx18797, nx18798, nx18799, 
         nx18800, nx18801, nx18802, nx18803, nx18804, nx18805, nx18806, nx18807, 
         NOT_nx3910, nx18808, nx18809, nx18810, nx18811, nx18812, nx18813, 
         nx18814, nx18815, nx18816, nx17531, nx18817, nx17571, nx18818, nx18819, 
         nx18820, nx18135, nx18821, nx18822, nx18075, nx17536, nx18823, nx18824, 
         nx18213, nx17977, nx4250, nx17450, nx18825, nx17409, nx18826, nx18827, 
         nx18828, nx18829, nx18830, nx18831, nx18832, nx17247, nx17250, nx18833, 
         nx18834, nx18835, nx18836, nx18837, nx18838, nx17533, nx18839, nx17406, 
         nx18840, nx18841, nx18842, nx18843, nx3760, nx17577, nx4736, nx18844, 
         nx18845, nx18846, nx18847, nx17257, nx3728, nx17130, nx18848, nx18849, 
         nx18850, nx18851, nx18852, nx18853, nx18854, nx18855, nx4012, nx18856, 
         nx18857, nx18858, nx17260, nx18859, nx18860, nx18861, nx18862, nx18863, 
         nx18864, nx18865, nx18866, nx16998, nx18867, nx18868, nx3216, nx16937, 
         nx18869, nx18870, nx18871, nx18872, nx18873, nx18874, nx4580, nx18875, 
         nx18876, nx18877, nx18878, nx18879, nx18880, nx17142, nx18881, nx18882, 
         nx18883, nx18884, nx18885, nx18886, nx18887, nx18888, nx18889, nx18890, 
         nx18891, nx18892, nx18893, nx18894, nx18895, nx18896, nx18897, nx18898, 
         nx18899, nx18900, nx18901, nx18902, nx18903, nx18904, nx18905, nx18906, 
         nx18907, nx18908, nx18909, nx18910, nx18911, nx18912, nx18913, nx18914, 
         nx18915, nx18916, nx19292, nx19294, nx19296, nx19298, nx19300, nx19302, 
         nx19308;
    wire [148:0] \$dummy ;




    assign wind_rst = io_done_out ;
    assign filter_reset = reset ;
    assign comp_unit_relu = io_done_out ;
    Cache_5_16_28_5 img_cache (.in_word ({cache_data_in_15,cache_data_in_14,
                    cache_data_in_13,cache_data_in_12,cache_data_in_11,
                    cache_data_in_10,cache_data_in_9,cache_data_in_8,
                    cache_data_in_7,cache_data_in_6,cache_data_in_5,
                    cache_data_in_4,cache_data_in_3,cache_data_in_2,
                    cache_data_in_1,cache_data_in_0}), .cache_in_sel ({nx17815,
                    cache_width_count_3,nx17819,cache_width_count_1,
                    cache_width_count_0}), .cache_out_sel ({wind_width_count_4,
                    wind_width_count_3,wind_width_count_2,wind_width_count_1,
                    nx17811}), .decoder_enable (cache_load), .out_column_0__15 (
                    cache_data_out_4__15), .out_column_0__14 (
                    cache_data_out_4__14), .out_column_0__13 (
                    cache_data_out_4__13), .out_column_0__12 (
                    cache_data_out_4__12), .out_column_0__11 (
                    cache_data_out_4__11), .out_column_0__10 (
                    cache_data_out_4__10), .out_column_0__9 (cache_data_out_4__9
                    ), .out_column_0__8 (cache_data_out_4__8), .out_column_0__7 (
                    cache_data_out_4__7), .out_column_0__6 (cache_data_out_4__6)
                    , .out_column_0__5 (cache_data_out_4__5), .out_column_0__4 (
                    cache_data_out_4__4), .out_column_0__3 (cache_data_out_4__3)
                    , .out_column_0__2 (cache_data_out_4__2), .out_column_0__1 (
                    cache_data_out_4__1), .out_column_0__0 (cache_data_out_4__0)
                    , .out_column_1__15 (cache_data_out_3__15), .out_column_1__14 (
                    cache_data_out_3__14), .out_column_1__13 (
                    cache_data_out_3__13), .out_column_1__12 (
                    cache_data_out_3__12), .out_column_1__11 (
                    cache_data_out_3__11), .out_column_1__10 (
                    cache_data_out_3__10), .out_column_1__9 (cache_data_out_3__9
                    ), .out_column_1__8 (cache_data_out_3__8), .out_column_1__7 (
                    cache_data_out_3__7), .out_column_1__6 (cache_data_out_3__6)
                    , .out_column_1__5 (cache_data_out_3__5), .out_column_1__4 (
                    cache_data_out_3__4), .out_column_1__3 (cache_data_out_3__3)
                    , .out_column_1__2 (cache_data_out_3__2), .out_column_1__1 (
                    cache_data_out_3__1), .out_column_1__0 (cache_data_out_3__0)
                    , .out_column_2__15 (cache_data_out_2__15), .out_column_2__14 (
                    cache_data_out_2__14), .out_column_2__13 (
                    cache_data_out_2__13), .out_column_2__12 (
                    cache_data_out_2__12), .out_column_2__11 (
                    cache_data_out_2__11), .out_column_2__10 (
                    cache_data_out_2__10), .out_column_2__9 (cache_data_out_2__9
                    ), .out_column_2__8 (cache_data_out_2__8), .out_column_2__7 (
                    cache_data_out_2__7), .out_column_2__6 (cache_data_out_2__6)
                    , .out_column_2__5 (cache_data_out_2__5), .out_column_2__4 (
                    cache_data_out_2__4), .out_column_2__3 (cache_data_out_2__3)
                    , .out_column_2__2 (cache_data_out_2__2), .out_column_2__1 (
                    cache_data_out_2__1), .out_column_2__0 (cache_data_out_2__0)
                    , .out_column_3__15 (cache_data_out_1__15), .out_column_3__14 (
                    cache_data_out_1__14), .out_column_3__13 (
                    cache_data_out_1__13), .out_column_3__12 (
                    cache_data_out_1__12), .out_column_3__11 (
                    cache_data_out_1__11), .out_column_3__10 (
                    cache_data_out_1__10), .out_column_3__9 (cache_data_out_1__9
                    ), .out_column_3__8 (cache_data_out_1__8), .out_column_3__7 (
                    cache_data_out_1__7), .out_column_3__6 (cache_data_out_1__6)
                    , .out_column_3__5 (cache_data_out_1__5), .out_column_3__4 (
                    cache_data_out_1__4), .out_column_3__3 (cache_data_out_1__3)
                    , .out_column_3__2 (cache_data_out_1__2), .out_column_3__1 (
                    cache_data_out_1__1), .out_column_3__0 (cache_data_out_1__0)
                    , .out_column_4__15 (cache_data_out_0__15), .out_column_4__14 (
                    cache_data_out_0__14), .out_column_4__13 (
                    cache_data_out_0__13), .out_column_4__12 (
                    cache_data_out_0__12), .out_column_4__11 (
                    cache_data_out_0__11), .out_column_4__10 (
                    cache_data_out_0__10), .out_column_4__9 (cache_data_out_0__9
                    ), .out_column_4__8 (cache_data_out_0__8), .out_column_4__7 (
                    cache_data_out_0__7), .out_column_4__6 (cache_data_out_0__6)
                    , .out_column_4__5 (cache_data_out_0__5), .out_column_4__4 (
                    cache_data_out_0__4), .out_column_4__3 (cache_data_out_0__3)
                    , .out_column_4__2 (cache_data_out_0__2), .out_column_4__1 (
                    cache_data_out_0__1), .out_column_4__0 (cache_data_out_0__0)
                    , .clk (nx17823), .reset (cache_rst_actual)) ;
    AdvancedCounter_16 cache_height_cntr (.clk (clk), .reset (nx17805), .enable (
                       cache_height_count_en), .mode_in ({io_done_out,
                       io_done_out}), .max_val_in ({io_done_out,io_done_out,
                       io_done_out,io_done_out,io_done_out,io_done_out,
                       io_done_out,io_done_out,io_done_out,io_done_out,
                       io_done_out,max_height_4,max_height_3,max_height_2,
                       max_height_1,max_height_0}), .max_reached_out (
                       cache_height_ended), .counter_out ({\$dummy [0],
                       \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],
                       \$dummy [5],\$dummy [6],\$dummy [7],\$dummy [8],
                       \$dummy [9],\$dummy [10],\$dummy [11],\$dummy [12],
                       \$dummy [13],\$dummy [14],\$dummy [15]})) ;
    fake_gnd ix12710 (.Y (io_done_out)) ;
    oai21 ix321 (.Y (filter_ready_out), .A0 (nx18255), .A1 (nx15396), .B0 (
          nx16313)) ;
    dffr reg_current_state_11 (.Q (\$dummy [16]), .QB (nx15392), .D (nx17865), .CLK (
         nx17823), .R (reset)) ;
    nand04 ix15403 (.Y (nx15402), .A0 (cntr1_inst_counter_out_3), .A1 (
           cntr1_inst_counter_out_2), .A2 (cntr1_inst_counter_out_1), .A3 (
           cntr1_inst_counter_out_0)) ;
    dffr reg_cntr1_inst_counter_out_3 (.Q (cntr1_inst_counter_out_3), .QB (
         \$dummy [17]), .D (nx13001), .CLK (clk), .R (nx17929)) ;
    xnor2 ix245 (.Y (nx244), .A0 (cntr1_inst_counter_out_3), .A1 (nx15407)) ;
    nand03 ix15408 (.Y (nx15407), .A0 (cntr1_inst_counter_out_2), .A1 (
           cntr1_inst_counter_out_1), .A2 (cntr1_inst_counter_out_0)) ;
    dffr reg_cntr1_inst_counter_out_2 (.Q (cntr1_inst_counter_out_2), .QB (
         \$dummy [18]), .D (nx12991), .CLK (clk), .R (nx17929)) ;
    xnor2 ix231 (.Y (nx230), .A0 (cntr1_inst_counter_out_2), .A1 (nx15412)) ;
    nand02 ix15413 (.Y (nx15412), .A0 (cntr1_inst_counter_out_1), .A1 (
           cntr1_inst_counter_out_0)) ;
    dffr reg_cntr1_inst_counter_out_1 (.Q (cntr1_inst_counter_out_1), .QB (
         nx15416), .D (nx12981), .CLK (clk), .R (nx17929)) ;
    oai21 ix183 (.Y (nx182), .A0 (nx15422), .A1 (nx15537), .B0 (nx16302)) ;
    mux21 ix13992 (.Y (nx13991), .A0 (nx15426), .A1 (nx15428), .S0 (nx17973)) ;
    dffr num_channels_counter_out_4 (.Q (\$dummy [19]), .QB (nx15426), .D (
         nx13991), .CLK (clk), .R (reset)) ;
    aoi222 ix15429 (.Y (nx15428), .A0 (max_num_channels_data_out_4), .A1 (nx1642
           ), .B0 (mem_data_in[4]), .B1 (nx17899), .C0 (nx18271), .C1 (nx1712)
           ) ;
    oai22 ix13982 (.Y (nx13981), .A0 (nx15432), .A1 (nx582), .B0 (nx16299), .B1 (
          nx15435)) ;
    dffr max_num_channels_inst_reg_q_4 (.Q (max_num_channels_data_out_4), .QB (
         nx15432), .D (nx13981), .CLK (clk), .R (reset)) ;
    and02 ix119 (.Y (nx118), .A0 (current_state_8), .A1 (nx15546)) ;
    dffr reg_current_state_8 (.Q (current_state_8), .QB (\$dummy [20]), .D (
         nx17907), .CLK (nx17837), .R (reset)) ;
    dffr reg_current_state_7 (.Q (current_state_7), .QB (\$dummy [21]), .D (
         current_state_6), .CLK (nx17835), .R (reset)) ;
    dffr reg_current_state_6 (.Q (current_state_6), .QB (\$dummy [22]), .D (
         current_state_5), .CLK (nx17835), .R (reset)) ;
    dffr reg_current_state_5 (.Q (current_state_5), .QB (\$dummy [23]), .D (
         nx17895), .CLK (nx17835), .R (reset)) ;
    dffr reg_current_state_4 (.Q (current_state_4), .QB (\$dummy [24]), .D (
         current_state_3), .CLK (nx17835), .R (reset)) ;
    dffr reg_current_state_3 (.Q (current_state_3), .QB (\$dummy [25]), .D (
         nx12910), .CLK (nx17835), .R (reset)) ;
    dffr reg_current_state_2 (.Q (current_state_2), .QB (nx15445), .D (nx140), .CLK (
         nx17823), .R (reset)) ;
    oai21 ix135 (.Y (nx134), .A0 (io_ready_in), .A1 (nx15450), .B0 (nx15452)) ;
    dffr reg_current_state_1 (.Q (\$dummy [26]), .QB (nx15450), .D (nx134), .CLK (
         nx17823), .R (reset)) ;
    dffs_ni reg_current_state_0 (.Q (\$dummy [27]), .QB (nx15452), .D (
            io_done_out), .CLK (nx17823), .S (reset)) ;
    nand02 ix1733 (.Y (nx12875), .A0 (nx15460), .A1 (nx15426)) ;
    nor04 ix15461 (.Y (nx15460), .A0 (num_channels_counter_out_0), .A1 (
          num_channels_counter_out_1), .A2 (num_channels_counter_out_2), .A3 (
          num_channels_counter_out_3)) ;
    mux21_ni ix13912 (.Y (nx13911), .A0 (num_channels_counter_out_0), .A1 (
             nx1618), .S0 (nx17973)) ;
    mux21_ni ix1619 (.Y (nx1618), .A0 (nx1608), .A1 (nx15531), .S0 (nx18269)) ;
    nand03 ix1609 (.Y (nx1608), .A0 (nx15466), .A1 (nx15474), .A2 (nx15445)) ;
    oai21 ix15467 (.Y (nx15466), .A0 (max_num_channels_data_out_0), .A1 (nx18151
          ), .B0 (nx17887)) ;
    oai32 ix13902 (.Y (nx13901), .A0 (nx15470), .A1 (nx17897), .A2 (nx17875), .B0 (
          nx15474), .B1 (nx18259)) ;
    dffr max_num_channels_inst_reg_q_0 (.Q (max_num_channels_data_out_0), .QB (
         nx15470), .D (nx13901), .CLK (clk), .R (reset)) ;
    dffr reg_current_state_9 (.Q (\$dummy [28]), .QB (nx15435), .D (nx118), .CLK (
         nx17823), .R (reset)) ;
    dffr reg_current_state_26 (.Q (current_state_26), .QB (\$dummy [29]), .D (
         nx1796), .CLK (nx17823), .R (reset)) ;
    aoi22 ix15475 (.Y (nx15474), .A0 (mem_data_in[0]), .A1 (nx17897), .B0 (
          nx17875), .B1 (nflt_layer_temp_0)) ;
    dffr nflt_layer_total_reg_q_0 (.Q (nflt_layer_temp_0), .QB (\$dummy [30]), .D (
         nx13891), .CLK (clk), .R (reset)) ;
    mux21_ni ix13892 (.Y (nx13891), .A0 (nflt_layer_temp_0), .A1 (mem_data_in[0]
             ), .S0 (nx17893)) ;
    dffr layer_type_reg_q_0 (.Q (comp_unit_operation), .QB (\$dummy [31]), .D (
         nx12961), .CLK (clk), .R (reset)) ;
    mux21_ni ix12962 (.Y (nx12961), .A0 (nx18151), .A1 (mem_data_in[0]), .S0 (
             current_state_3)) ;
    dffr reg_current_state_25 (.Q (\$dummy [32]), .QB (nx15530), .D (nx92), .CLK (
         nx17825), .R (reset)) ;
    oai32 ix12922 (.Y (nx12921), .A0 (nx15488), .A1 (nx17893), .A2 (nx17887), .B0 (
          nx15491), .B1 (nx18263)) ;
    dffr reg_nflt_layer_out_0 (.Q (nflt_layer_out_0), .QB (nx15488), .D (nx12921
         ), .CLK (clk), .R (reset)) ;
    oai32 ix12932 (.Y (nx12931), .A0 (nx15500), .A1 (nx17893), .A2 (nx17887), .B0 (
          nx15502), .B1 (nx18263)) ;
    dffr reg_nflt_layer_out_1 (.Q (nflt_layer_out_1), .QB (nx15500), .D (nx12931
         ), .CLK (clk), .R (reset)) ;
    mux21_ni ix15503 (.Y (nx15502), .A0 (nx15504), .A1 (nx15508), .S0 (nx17893)
             ) ;
    aoi21 ix15505 (.Y (nx15504), .A0 (nflt_layer_out_1), .A1 (nflt_layer_out_0)
          , .B0 (nx15506)) ;
    inv01 ix15509 (.Y (nx15508), .A (mem_data_in[1])) ;
    oai32 ix12942 (.Y (nx12941), .A0 (nx15512), .A1 (nx17893), .A2 (nx17887), .B0 (
          nx15514), .B1 (nx18263)) ;
    dffr nflt_layer_out_2 (.Q (\$dummy [33]), .QB (nx15512), .D (nx12941), .CLK (
         clk), .R (reset)) ;
    mux21_ni ix15515 (.Y (nx15514), .A0 (nx15516), .A1 (nx15518), .S0 (nx17895)
             ) ;
    inv01 ix15519 (.Y (nx15518), .A (mem_data_in[2])) ;
    dffr reg_nflt_layer_out_3 (.Q (nflt_layer_out_3), .QB (\$dummy [34]), .D (
         nx12951), .CLK (clk), .R (reset)) ;
    mux21_ni ix12952 (.Y (nx12951), .A0 (nx78), .A1 (nflt_layer_out_3), .S0 (
             nx18263)) ;
    mux21 ix79 (.Y (nx78), .A0 (nx15523), .A1 (nx15527), .S0 (nx17895)) ;
    xnor2 ix15524 (.Y (nx15523), .A0 (nflt_layer_out_3), .A1 (nx15525)) ;
    inv01 ix15528 (.Y (nx15527), .A (mem_data_in[3])) ;
    dffr reg_num_channels_counter_out_0 (.Q (num_channels_counter_out_0), .QB (
         nx15531), .D (nx13911), .CLK (clk), .R (reset)) ;
    oai21 ix1547 (.Y (nx1546), .A0 (nx15422), .A1 (nx15537), .B0 (nx18269)) ;
    nand02 ix15538 (.Y (nx15537), .A0 (current_state_24), .A1 (nx15637)) ;
    oai21 ix1535 (.Y (nx1534), .A0 (nx15541), .A1 (nx17847), .B0 (nx15716)) ;
    nand02 ix1519 (.Y (nx1518), .A0 (nx15544), .A1 (nx16065)) ;
    aoi32 ix15545 (.Y (nx15544), .A0 (nx15546), .A1 (comp_unit_finished), .A2 (
          current_state_19), .B0 (nx15561), .B1 (nx12906)) ;
    mux21_ni ix14032 (.Y (nx14031), .A0 (layer_type_out_1), .A1 (mem_data_in[1])
             , .S0 (current_state_3)) ;
    dffr layer_type_reg_q_1 (.Q (layer_type_out_1), .QB (nx15548), .D (nx14031)
         , .CLK (clk), .R (reset)) ;
    oai221 ix1501 (.Y (nx1500), .A0 (nx18273), .A1 (nx17847), .B0 (
           comp_unit_finished), .B1 (nx15573), .C0 (nx18059)) ;
    dffr reg_current_state_17 (.Q (\$dummy [35]), .QB (nx15554), .D (nx1478), .CLK (
         nx17835), .R (reset)) ;
    mux21 ix13342 (.Y (nx13341), .A0 (nx15559), .A1 (nx15575), .S0 (nx18045)) ;
    aoi32 ix15560 (.Y (nx15559), .A0 (nx15561), .A1 (ftc_cntrl_reg_out_11), .A2 (
          current_state_21), .B0 (ftc_cntrl_reg_out_8), .B1 (nx158)) ;
    mux21_ni ix13072 (.Y (nx13071), .A0 (nx362), .A1 (ftc_cntrl_reg_out_14), .S0 (
             nx18045)) ;
    oai22 ix363 (.Y (nx362), .A0 (nx15561), .A1 (nx15567), .B0 (nx15563), .B1 (
          nx16198)) ;
    aoi21 ix15568 (.Y (nx15567), .A0 (nx17873), .A1 (nx15621), .B0 (
          current_state_21)) ;
    oai321 ix1839 (.Y (nx1838), .A0 (nx15546), .A1 (nx15571), .A2 (nx15573), .B0 (
           nx15575), .B1 (nx15602), .C0 (nx16196)) ;
    inv01 ix15572 (.Y (nx15571), .A (comp_unit_finished)) ;
    dffr reg_current_state_19 (.Q (current_state_19), .QB (nx15573), .D (nx1500)
         , .CLK (nx17825), .R (reset)) ;
    dffr ftc_cntrl_reg_reg_q_8 (.Q (ftc_cntrl_reg_out_8), .QB (nx15575), .D (
         nx13341), .CLK (nx17825), .R (nx17805)) ;
    dffr reg_current_state_13 (.Q (current_state_13), .QB (\$dummy [36]), .D (
         nx330), .CLK (nx17825), .R (reset)) ;
    oai22 ix331 (.Y (nx330), .A0 (nx18255), .A1 (nx316), .B0 (nx15598), .B1 (
          nx196)) ;
    nand04 ix317 (.Y (nx316), .A0 (nx15580), .A1 (cntr1_inst_counter_out_0), .A2 (
           cntr1_inst_counter_out_3), .A3 (nx15596)) ;
    nor03_2x ix15581 (.Y (nx15580), .A0 (nx310), .A1 (nx278), .A2 (nx276)) ;
    dffr cntr1_inst_counter_out_5 (.Q (\$dummy [37]), .QB (nx15586), .D (nx13021
         ), .CLK (clk), .R (nx17929)) ;
    dffr reg_cntr1_inst_counter_out_4 (.Q (cntr1_inst_counter_out_4), .QB (
         nx15591), .D (nx13011), .CLK (clk), .R (nx17929)) ;
    dffr reg_cntr1_inst_counter_out_0 (.Q (cntr1_inst_counter_out_0), .QB (
         \$dummy [38]), .D (nx12971), .CLK (clk), .R (nx17929)) ;
    xnor2 ix12972 (.Y (nx12971), .A0 (cntr1_inst_counter_out_0), .A1 (nx18255)
          ) ;
    dffr reg_current_state_10 (.Q (current_state_10), .QB (nx15598), .D (nx182)
         , .CLK (nx17825), .R (reset)) ;
    nand02 ix197 (.Y (nx196), .A0 (nx18151), .A1 (nx15548)) ;
    dffr reg_current_state_20 (.Q (\$dummy [39]), .QB (nx15605), .D (nx1838), .CLK (
         nx17825), .R (reset)) ;
    mux21 ix13852 (.Y (nx13851), .A0 (nx15609), .A1 (nx15621), .S0 (nx18045)) ;
    nand04 ix15610 (.Y (nx15609), .A0 (nx1402), .A1 (nx1416), .A2 (nx1434), .A3 (
           nx1456)) ;
    dffr cache_width_cntr_counter_out_15 (.Q (\$dummy [40]), .QB (nx15614), .D (
         nx13841), .CLK (clk), .R (nx17961)) ;
    nand02 ix1225 (.Y (nx1224), .A0 (nx15617), .A1 (nx16065)) ;
    aoi21 ix15618 (.Y (nx15617), .A0 (nx15619), .A1 (nx17921), .B0 (nx17807)) ;
    dffr ftc_cntrl_reg_reg_q_12 (.Q (ftc_cntrl_reg_out_12), .QB (nx15621), .D (
         nx13851), .CLK (nx17825), .R (nx17805)) ;
    or02 ix337 (.Y (nx336), .A0 (nx12883), .A1 (nx17805)) ;
    dffr reg_current_state_14 (.Q (\$dummy [41]), .QB (nx15626), .D (nx336), .CLK (
         nx17827), .R (reset)) ;
    mux21_ni ix13062 (.Y (nx13061), .A0 (cache_height_ended), .A1 (
             ftc_cntrl_reg_out_13), .S0 (nx18045)) ;
    dffr reg_current_state_15 (.Q (current_state_15), .QB (nx15861), .D (nx1138)
         , .CLK (nx17833), .R (reset)) ;
    oai22 ix1139 (.Y (nx1138), .A0 (nx15635), .A1 (nx15637), .B0 (nx18279), .B1 (
          nx15859)) ;
    dffr reg_current_state_24 (.Q (current_state_24), .QB (nx15635), .D (nx1534)
         , .CLK (nx17827), .R (reset)) ;
    nor04 ix15638 (.Y (nx15637), .A0 (nx1128), .A1 (nx1040), .A2 (nx944), .A3 (
          nx850)) ;
    nand04 ix1129 (.Y (nx1128), .A0 (nx15640), .A1 (nx15781), .A2 (nx15786), .A3 (
           nx15791)) ;
    oai22 ix13652 (.Y (nx13651), .A0 (nx15644), .A1 (nx18053), .B0 (nx15776), .B1 (
          nx17951)) ;
    dffr reg_write_offset_reg_q_14 (.Q (write_offset_data_out_14), .QB (nx15647)
         , .D (nx13631), .CLK (nx17827), .R (reset)) ;
    nand02 ix15654 (.Y (nx15653), .A0 (write_offset_data_out_13), .A1 (nx1042)
           ) ;
    oai22 ix13612 (.Y (nx13611), .A0 (nx15657), .A1 (nx18053), .B0 (nx15774), .B1 (
          nx17949)) ;
    oai21 ix15658 (.Y (nx15657), .A0 (nx1042), .A1 (write_offset_data_out_13), .B0 (
          nx15653)) ;
    dffr reg_write_offset_reg_q_12 (.Q (write_offset_data_out_12), .QB (nx15660)
         , .D (nx13591), .CLK (nx17827), .R (reset)) ;
    nand02 ix15667 (.Y (nx15666), .A0 (write_offset_data_out_11), .A1 (nx994)) ;
    oai22 ix13572 (.Y (nx13571), .A0 (nx15670), .A1 (nx18051), .B0 (nx15772), .B1 (
          nx17949)) ;
    oai21 ix15671 (.Y (nx15670), .A0 (nx994), .A1 (write_offset_data_out_11), .B0 (
          nx15666)) ;
    dffr reg_write_offset_reg_q_10 (.Q (write_offset_data_out_10), .QB (nx15673)
         , .D (nx13551), .CLK (nx17827), .R (reset)) ;
    nand02 ix15680 (.Y (nx15679), .A0 (write_offset_data_out_9), .A1 (nx948)) ;
    oai22 ix13532 (.Y (nx13531), .A0 (nx15683), .A1 (nx18051), .B0 (nx15770), .B1 (
          nx17949)) ;
    oai21 ix15684 (.Y (nx15683), .A0 (nx948), .A1 (write_offset_data_out_9), .B0 (
          nx15679)) ;
    dffr reg_write_offset_reg_q_8 (.Q (write_offset_data_out_8), .QB (nx15686), 
         .D (nx13511), .CLK (nx17827), .R (reset)) ;
    nand02 ix15693 (.Y (nx15692), .A0 (write_offset_data_out_7), .A1 (nx898)) ;
    oai22 ix13492 (.Y (nx13491), .A0 (nx15696), .A1 (nx17947), .B0 (nx15717), .B1 (
          nx18051)) ;
    dffr reg_write_offset_reg_q_7 (.Q (write_offset_data_out_7), .QB (nx15696), 
         .D (nx13491), .CLK (nx17827), .R (reset)) ;
    dffr reg_current_state_22 (.Q (\$dummy [42]), .QB (nx15541), .D (nx1518), .CLK (
         nx17829), .R (reset)) ;
    dffr reg_current_state_23 (.Q (\$dummy [43]), .QB (nx15716), .D (nx1524), .CLK (
         nx17829), .R (reset)) ;
    mux21_ni ix13032 (.Y (nx13031), .A0 (flt_size_out_0), .A1 (mem_data_in[0]), 
             .S0 (current_state_5)) ;
    dffr flt_size_reg_q_0 (.Q (flt_size_out_0), .QB (\$dummy [44]), .D (nx13031)
         , .CLK (clk), .R (reset)) ;
    dffr flt_size_reg_q_2 (.Q (flt_size_out_2), .QB (nx15711), .D (nx13041), .CLK (
         clk), .R (reset)) ;
    mux21_ni ix13042 (.Y (nx13041), .A0 (flt_size_out_2), .A1 (mem_data_in[2]), 
             .S0 (current_state_5)) ;
    mux21_ni ix13052 (.Y (nx13051), .A0 (flt_size_out_1), .A1 (mem_data_in[1]), 
             .S0 (current_state_5)) ;
    dffr flt_size_reg_q_1 (.Q (flt_size_out_1), .QB (\$dummy [45]), .D (nx13051)
         , .CLK (clk), .R (reset)) ;
    oai21 ix15718 (.Y (nx15717), .A0 (nx898), .A1 (write_offset_data_out_7), .B0 (
          nx15692)) ;
    dffr reg_write_offset_reg_q_6 (.Q (write_offset_data_out_6), .QB (nx15720), 
         .D (nx13471), .CLK (nx17829), .R (reset)) ;
    nand02 ix15727 (.Y (nx15726), .A0 (write_offset_data_out_5), .A1 (nx852)) ;
    oai22 ix13452 (.Y (nx13451), .A0 (nx15730), .A1 (nx17947), .B0 (nx15732), .B1 (
          nx18049)) ;
    dffr reg_write_offset_reg_q_5 (.Q (write_offset_data_out_5), .QB (nx15730), 
         .D (nx13451), .CLK (nx17829), .R (reset)) ;
    oai21 ix15733 (.Y (nx15732), .A0 (nx852), .A1 (write_offset_data_out_5), .B0 (
          nx15726)) ;
    dffr reg_write_offset_reg_q_4 (.Q (write_offset_data_out_4), .QB (nx15735), 
         .D (nx13431), .CLK (nx17829), .R (reset)) ;
    dffr reg_write_offset_reg_q_3 (.Q (write_offset_data_out_3), .QB (nx15745), 
         .D (nx13411), .CLK (nx17829), .R (reset)) ;
    oai22 ix13392 (.Y (nx13391), .A0 (nx15750), .A1 (nx17947), .B0 (nx15753), .B1 (
          nx18049)) ;
    oai21 ix15754 (.Y (nx15753), .A0 (nx780), .A1 (write_offset_data_out_2), .B0 (
          nx15768)) ;
    oai22 ix13372 (.Y (nx13371), .A0 (nx15756), .A1 (nx17947), .B0 (nx15759), .B1 (
          nx18049)) ;
    oai21 ix15760 (.Y (nx15759), .A0 (write_offset_data_out_0), .A1 (
          write_offset_data_out_1), .B0 (nx15765)) ;
    dffr reg_write_offset_reg_q_0 (.Q (write_offset_data_out_0), .QB (nx15763), 
         .D (nx13351), .CLK (nx17829), .R (reset)) ;
    dffr reg_write_offset_reg_q_1 (.Q (write_offset_data_out_1), .QB (nx15756), 
         .D (nx13371), .CLK (nx17831), .R (reset)) ;
    dffr reg_write_offset_reg_q_2 (.Q (write_offset_data_out_2), .QB (nx15750), 
         .D (nx13391), .CLK (nx17831), .R (reset)) ;
    dffr reg_write_offset_reg_q_9 (.Q (write_offset_data_out_9), .QB (nx15770), 
         .D (nx13531), .CLK (nx17831), .R (reset)) ;
    dffr reg_write_offset_reg_q_11 (.Q (write_offset_data_out_11), .QB (nx15772)
         , .D (nx13571), .CLK (nx17831), .R (reset)) ;
    dffr reg_write_offset_reg_q_13 (.Q (write_offset_data_out_13), .QB (nx15774)
         , .D (nx13611), .CLK (nx17831), .R (reset)) ;
    dffr reg_write_offset_reg_q_15 (.Q (write_offset_data_out_15), .QB (nx15776)
         , .D (nx13651), .CLK (nx17831), .R (reset)) ;
    dffr new_size_squared_reg_q_15 (.Q (new_size_squared_out_15), .QB (
         \$dummy [46]), .D (nx13661), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_14 (.Q (new_size_squared_out_14), .QB (nx15785)
         , .D (nx13641), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_13 (.Q (new_size_squared_out_13), .QB (
         \$dummy [47]), .D (nx13621), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_12 (.Q (new_size_squared_out_12), .QB (nx15795)
         , .D (nx13601), .CLK (clk), .R (reset)) ;
    nand04 ix1041 (.Y (nx1040), .A0 (nx15797), .A1 (nx15802), .A2 (nx15807), .A3 (
           nx15812)) ;
    dffr new_size_squared_reg_q_11 (.Q (new_size_squared_out_11), .QB (
         \$dummy [48]), .D (nx13581), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_10 (.Q (new_size_squared_out_10), .QB (nx15806)
         , .D (nx13561), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_9 (.Q (new_size_squared_out_9), .QB (
         \$dummy [49]), .D (nx13541), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_8 (.Q (new_size_squared_out_8), .QB (nx15816), .D (
         nx13521), .CLK (clk), .R (reset)) ;
    nand04 ix945 (.Y (nx944), .A0 (nx15818), .A1 (nx15823), .A2 (nx15828), .A3 (
           nx15833)) ;
    dffr new_size_squared_reg_q_7 (.Q (new_size_squared_out_7), .QB (
         \$dummy [50]), .D (nx13501), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_6 (.Q (new_size_squared_out_6), .QB (nx15827), .D (
         nx13481), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_5 (.Q (new_size_squared_out_5), .QB (
         \$dummy [51]), .D (nx13461), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_4 (.Q (new_size_squared_out_4), .QB (nx15837), .D (
         nx13441), .CLK (clk), .R (reset)) ;
    nand04 ix851 (.Y (nx850), .A0 (nx15839), .A1 (nx15844), .A2 (nx15849), .A3 (
           nx15854)) ;
    dffr new_size_squared_reg_q_3 (.Q (new_size_squared_out_3), .QB (
         \$dummy [52]), .D (nx13421), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_2 (.Q (new_size_squared_out_2), .QB (nx15848), .D (
         nx13401), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_1 (.Q (new_size_squared_out_1), .QB (
         \$dummy [53]), .D (nx13381), .CLK (clk), .R (reset)) ;
    dffr new_size_squared_reg_q_0 (.Q (new_size_squared_out_0), .QB (
         \$dummy [54]), .D (nx13361), .CLK (clk), .R (reset)) ;
    dffr ftc_cntrl_reg_reg_q_13 (.Q (ftc_cntrl_reg_out_13), .QB (nx15859), .D (
         nx13061), .CLK (nx17831), .R (nx17805)) ;
    nand02 ix1169 (.Y (nx1168), .A0 (nx18225), .A1 (nx15878)) ;
    mux21 ix13332 (.Y (nx13331), .A0 (nx15868), .A1 (nx15865), .S0 (nx18045)) ;
    nand04 ix15869 (.Y (nx15868), .A0 (nx550), .A1 (nx564), .A2 (nx612), .A3 (
           nx732)) ;
    dffr window_width_cntr_counter_out_15 (.Q (\$dummy [55]), .QB (nx15873), .D (
         nx13221), .CLK (clk), .R (nx17939)) ;
    nand02 ix379 (.Y (nx378), .A0 (nx15876), .A1 (nx15878)) ;
    aoi22 ix15877 (.Y (nx15876), .A0 (nx17921), .A1 (ftc_cntrl_reg_out_13), .B0 (
          nx17871), .B1 (ftc_cntrl_reg_out_12)) ;
    mux21_ni ix13672 (.Y (nx13671), .A0 (nx1154), .A1 (ftc_cntrl_reg_out_9), .S0 (
             nx18045)) ;
    oai21 ix1155 (.Y (nx1154), .A0 (nx15883), .A1 (nx15885), .B0 (nx15876)) ;
    dffr ftc_cntrl_reg_reg_q_9 (.Q (ftc_cntrl_reg_out_9), .QB (nx15883), .D (
         nx13671), .CLK (nx17833), .R (nx17805)) ;
    aoi21 ix15886 (.Y (nx15885), .A0 (nx18225), .A1 (nx1146), .B0 (nx17921)) ;
    dffr reg_current_state_16 (.Q (current_state_16), .QB (nx15888), .D (nx1168)
         , .CLK (nx17833), .R (reset)) ;
    dffr reg_window_width_cntr_counter_out_14 (.Q (
         window_width_cntr_counter_out_14), .QB (nx15893), .D (nx13211), .CLK (
         clk), .R (nx17939)) ;
    nand02 ix15899 (.Y (nx15898), .A0 (window_width_cntr_counter_out_13), .A1 (
           nx12887)) ;
    dffr reg_window_width_cntr_counter_out_13 (.Q (
         window_width_cntr_counter_out_13), .QB (nx15902), .D (nx13201), .CLK (
         clk), .R (nx17939)) ;
    oai21 ix15905 (.Y (nx15904), .A0 (nx12887), .A1 (
          window_width_cntr_counter_out_13), .B0 (nx15898)) ;
    dffr reg_window_width_cntr_counter_out_12 (.Q (
         window_width_cntr_counter_out_12), .QB (nx15907), .D (nx13191), .CLK (
         clk), .R (nx17939)) ;
    nand02 ix15913 (.Y (nx15912), .A0 (window_width_cntr_counter_out_11), .A1 (
           nx12889)) ;
    dffr reg_window_width_cntr_counter_out_11 (.Q (
         window_width_cntr_counter_out_11), .QB (nx15916), .D (nx13181), .CLK (
         clk), .R (nx17939)) ;
    oai21 ix15919 (.Y (nx15918), .A0 (nx12889), .A1 (
          window_width_cntr_counter_out_11), .B0 (nx15912)) ;
    dffr reg_window_width_cntr_counter_out_10 (.Q (
         window_width_cntr_counter_out_10), .QB (nx15921), .D (nx13171), .CLK (
         clk), .R (nx17939)) ;
    nand02 ix15927 (.Y (nx15926), .A0 (window_width_cntr_counter_out_9), .A1 (
           nx12891)) ;
    dffr reg_window_width_cntr_counter_out_9 (.Q (
         window_width_cntr_counter_out_9), .QB (nx15930), .D (nx13161), .CLK (
         clk), .R (nx17939)) ;
    oai21 ix15933 (.Y (nx15932), .A0 (nx12891), .A1 (
          window_width_cntr_counter_out_9), .B0 (nx15926)) ;
    dffr reg_window_width_cntr_counter_out_8 (.Q (
         window_width_cntr_counter_out_8), .QB (nx15935), .D (nx13151), .CLK (
         clk), .R (nx17941)) ;
    nand02 ix15941 (.Y (nx15940), .A0 (window_width_cntr_counter_out_7), .A1 (
           nx12893)) ;
    dffr reg_window_width_cntr_counter_out_7 (.Q (
         window_width_cntr_counter_out_7), .QB (nx15944), .D (nx13141), .CLK (
         clk), .R (nx17941)) ;
    oai21 ix15947 (.Y (nx15946), .A0 (nx12893), .A1 (
          window_width_cntr_counter_out_7), .B0 (nx15940)) ;
    dffr reg_window_width_cntr_counter_out_6 (.Q (
         window_width_cntr_counter_out_6), .QB (nx15949), .D (nx13131), .CLK (
         clk), .R (nx17941)) ;
    dffr reg_wind_width_count_4 (.Q (wind_width_count_4), .QB (\$dummy [56]), .D (
         nx14041), .CLK (clk), .R (nx17943)) ;
    xnor2 ix1877 (.Y (nx1876), .A0 (wind_width_count_4), .A1 (nx15959)) ;
    nand04 ix15960 (.Y (nx15959), .A0 (wind_width_count_1), .A1 (nx17811), .A2 (
           wind_width_count_2), .A3 (wind_width_count_3)) ;
    dffr reg_wind_width_count_1 (.Q (wind_width_count_1), .QB (\$dummy [57]), .D (
         nx13091), .CLK (clk), .R (nx17941)) ;
    xor2 ix385 (.Y (nx384), .A0 (wind_width_count_1), .A1 (nx17811)) ;
    dffr reg_wind_width_count_0 (.Q (wind_width_count_0), .QB (\$dummy [58]), .D (
         nx13081), .CLK (clk), .R (nx17941)) ;
    dffr reg_current_state_21 (.Q (current_state_21), .QB (nx15970), .D (nx12877
         ), .CLK (nx17833), .R (reset)) ;
    dffr ftc_cntrl_reg_reg_q_11 (.Q (ftc_cntrl_reg_out_11), .QB (nx15865), .D (
         nx13331), .CLK (nx17833), .R (nx17805)) ;
    oai22 ix1875 (.Y (nx12884), .A0 (ftc_cntrl_reg_out_9), .A1 (nx18225), .B0 (
          nx15970), .B1 (ftc_cntrl_reg_out_11)) ;
    dffr reg_wind_width_count_2 (.Q (wind_width_count_2), .QB (\$dummy [59]), .D (
         nx13101), .CLK (clk), .R (nx17941)) ;
    xnor2 ix393 (.Y (nx392), .A0 (wind_width_count_2), .A1 (nx15983)) ;
    nand02 ix15984 (.Y (nx15983), .A0 (wind_width_count_1), .A1 (nx17813)) ;
    dffr reg_wind_width_count_3 (.Q (wind_width_count_3), .QB (\$dummy [60]), .D (
         nx13111), .CLK (clk), .R (nx17941)) ;
    xnor2 ix401 (.Y (nx400), .A0 (wind_width_count_3), .A1 (nx15989)) ;
    nand03 ix15990 (.Y (nx15989), .A0 (wind_width_count_1), .A1 (nx17813), .A2 (
           wind_width_count_2)) ;
    dffr reg_window_width_cntr_counter_out_5 (.Q (
         window_width_cntr_counter_out_5), .QB (nx15995), .D (nx13121), .CLK (
         clk), .R (nx17943)) ;
    oai21 ix15998 (.Y (nx15997), .A0 (nx408), .A1 (
          window_width_cntr_counter_out_5), .B0 (nx15954)) ;
    nor02ii ix409 (.Y (nx408), .A0 (nx15959), .A1 (wind_width_count_4)) ;
    xor2 ix605 (.Y (nx604), .A0 (nx602), .A1 (nx17813)) ;
    dffr img_width_reg_q_0 (.Q (img_width_out_0), .QB (nx16005), .D (nx13241), .CLK (
         clk), .R (reset)) ;
    mux21_ni ix13232 (.Y (nx13231), .A0 (new_width_out_0), .A1 (mem_data_in[0])
             , .S0 (current_state_6)) ;
    dffr new_width_reg_q_0 (.Q (new_width_out_0), .QB (\$dummy [61]), .D (
         nx13231), .CLK (clk), .R (reset)) ;
    and04 ix733 (.Y (nx732), .A0 (nx16013), .A1 (nx16025), .A2 (nx16039), .A3 (
          nx16052)) ;
    xnor2 ix16014 (.Y (nx16013), .A0 (wind_width_count_1), .A1 (nx640)) ;
    dffr img_width_reg_q_1 (.Q (img_width_out_1), .QB (nx16019), .D (nx13261), .CLK (
         clk), .R (reset)) ;
    mux21_ni ix13252 (.Y (nx13251), .A0 (new_width_out_1), .A1 (mem_data_in[1])
             , .S0 (current_state_6)) ;
    dffr new_width_reg_q_1 (.Q (new_width_out_1), .QB (\$dummy [62]), .D (
         nx13251), .CLK (clk), .R (reset)) ;
    xnor2 ix16026 (.Y (nx16025), .A0 (wind_width_count_2), .A1 (nx674)) ;
    mux21 ix675 (.Y (nx674), .A0 (nx17845), .A1 (nx18055), .S0 (nx18225)) ;
    aoi21 ix16029 (.Y (nx16028), .A0 (img_width_out_2), .A1 (nx630), .B0 (
          nx16037)) ;
    dffs_ni img_width_reg_q_2 (.Q (img_width_out_2), .QB (\$dummy [63]), .D (
            nx13281), .CLK (clk), .S (reset)) ;
    ao221 ix13282 (.Y (nx13281), .A0 (nx17875), .A1 (new_width_out_2), .B0 (
          img_width_out_2), .B1 (nx18259), .C0 (nx17897)) ;
    dffr new_width_reg_q_2 (.Q (new_width_out_2), .QB (\$dummy [64]), .D (
         nx13271), .CLK (clk), .R (reset)) ;
    mux21_ni ix13272 (.Y (nx13271), .A0 (new_width_out_2), .A1 (mem_data_in[2])
             , .S0 (current_state_6)) ;
    nor03_2x ix16038 (.Y (nx16037), .A0 (img_width_out_0), .A1 (img_width_out_1)
             , .A2 (img_width_out_2)) ;
    xnor2 ix16040 (.Y (nx16039), .A0 (wind_width_count_3), .A1 (nx704)) ;
    dffs_ni img_width_reg_q_3 (.Q (img_width_out_3), .QB (nx16046), .D (nx13301)
            , .CLK (clk), .S (reset)) ;
    mux21_ni ix13292 (.Y (nx13291), .A0 (new_width_out_3), .A1 (mem_data_in[3])
             , .S0 (current_state_6)) ;
    dffr new_width_reg_q_3 (.Q (new_width_out_3), .QB (\$dummy [65]), .D (
         nx13291), .CLK (clk), .R (reset)) ;
    xnor2 ix16053 (.Y (nx16052), .A0 (wind_width_count_4), .A1 (nx722)) ;
    xnor2 ix16056 (.Y (nx16055), .A0 (img_width_out_4), .A1 (nx16063)) ;
    dffs_ni img_width_reg_q_4 (.Q (img_width_out_4), .QB (\$dummy [66]), .D (
            nx13321), .CLK (clk), .S (reset)) ;
    ao22 ix13322 (.Y (nx13321), .A0 (nx17875), .A1 (new_width_out_4), .B0 (
         img_width_out_4), .B1 (nx18259)) ;
    dffr new_width_reg_q_4 (.Q (new_width_out_4), .QB (\$dummy [67]), .D (
         nx13311), .CLK (clk), .R (reset)) ;
    mux21_ni ix13312 (.Y (nx13311), .A0 (new_width_out_4), .A1 (mem_data_in[4])
             , .S0 (current_state_6)) ;
    dffr reg_cache_width_cntr_counter_out_14 (.Q (
         cache_width_cntr_counter_out_14), .QB (nx16070), .D (nx13831), .CLK (
         clk), .R (nx17961)) ;
    nand02 ix16076 (.Y (nx16075), .A0 (cache_width_cntr_counter_out_13), .A1 (
           nx12898)) ;
    dffr reg_cache_width_cntr_counter_out_13 (.Q (
         cache_width_cntr_counter_out_13), .QB (nx16079), .D (nx13821), .CLK (
         clk), .R (nx17961)) ;
    oai21 ix16082 (.Y (nx16081), .A0 (nx12898), .A1 (
          cache_width_cntr_counter_out_13), .B0 (nx16075)) ;
    dffr reg_cache_width_cntr_counter_out_12 (.Q (
         cache_width_cntr_counter_out_12), .QB (nx16084), .D (nx13811), .CLK (
         clk), .R (nx17961)) ;
    nand02 ix16090 (.Y (nx16089), .A0 (cache_width_cntr_counter_out_11), .A1 (
           nx12900)) ;
    dffr reg_cache_width_cntr_counter_out_11 (.Q (
         cache_width_cntr_counter_out_11), .QB (nx16093), .D (nx13801), .CLK (
         clk), .R (nx17961)) ;
    oai21 ix16096 (.Y (nx16095), .A0 (nx12900), .A1 (
          cache_width_cntr_counter_out_11), .B0 (nx16089)) ;
    dffr reg_cache_width_cntr_counter_out_10 (.Q (
         cache_width_cntr_counter_out_10), .QB (nx16098), .D (nx13791), .CLK (
         clk), .R (nx17961)) ;
    nand02 ix16104 (.Y (nx16103), .A0 (cache_width_cntr_counter_out_9), .A1 (
           nx12902)) ;
    dffr reg_cache_width_cntr_counter_out_9 (.Q (cache_width_cntr_counter_out_9)
         , .QB (nx16107), .D (nx13781), .CLK (clk), .R (nx17961)) ;
    oai21 ix16110 (.Y (nx16109), .A0 (nx12902), .A1 (
          cache_width_cntr_counter_out_9), .B0 (nx16103)) ;
    dffr reg_cache_width_cntr_counter_out_8 (.Q (cache_width_cntr_counter_out_8)
         , .QB (nx16112), .D (nx13771), .CLK (clk), .R (nx17963)) ;
    nand02 ix16118 (.Y (nx16117), .A0 (cache_width_cntr_counter_out_7), .A1 (
           nx12904)) ;
    dffr reg_cache_width_cntr_counter_out_7 (.Q (cache_width_cntr_counter_out_7)
         , .QB (nx16121), .D (nx13761), .CLK (clk), .R (nx17963)) ;
    oai21 ix16124 (.Y (nx16123), .A0 (nx12904), .A1 (
          cache_width_cntr_counter_out_7), .B0 (nx16117)) ;
    dffr reg_cache_width_cntr_counter_out_6 (.Q (cache_width_cntr_counter_out_6)
         , .QB (nx16126), .D (nx13751), .CLK (clk), .R (nx17963)) ;
    dffr reg_cache_width_count_4 (.Q (cache_width_count_4), .QB (\$dummy [68]), 
         .D (nx13731), .CLK (clk), .R (nx17965)) ;
    xnor2 ix1255 (.Y (nx1254), .A0 (nx17815), .A1 (nx16136)) ;
    nand04 ix16137 (.Y (nx16136), .A0 (cache_width_count_1), .A1 (
           cache_width_count_0), .A2 (nx17819), .A3 (cache_width_count_3)) ;
    dffr reg_cache_width_count_1 (.Q (cache_width_count_1), .QB (\$dummy [69]), 
         .D (nx13701), .CLK (clk), .R (nx17963)) ;
    xor2 ix1231 (.Y (nx1230), .A0 (cache_width_count_1), .A1 (
         cache_width_count_0)) ;
    dffr reg_cache_width_count_0 (.Q (cache_width_count_0), .QB (\$dummy [70]), 
         .D (nx13691), .CLK (clk), .R (nx17963)) ;
    mux21_ni ix13682 (.Y (nx13681), .A0 (nx1206), .A1 (ftc_cntrl_reg_out_10), .S0 (
             nx18045)) ;
    oai21 ix1207 (.Y (nx1206), .A0 (nx16148), .A1 (nx16150), .B0 (nx16155)) ;
    dffr ftc_cntrl_reg_reg_q_10 (.Q (ftc_cntrl_reg_out_10), .QB (nx16148), .D (
         nx13681), .CLK (nx17833), .R (nx17807)) ;
    nor03_2x ix1195 (.Y (cache_height_count_en), .A0 (nx16153), .A1 (
             ftc_cntrl_reg_out_13), .A2 (nx15621)) ;
    oai21 ix16156 (.Y (nx16155), .A0 (nx17871), .A1 (nx12883), .B0 (nx15621)) ;
    dffr reg_cache_width_count_2 (.Q (cache_width_count_2), .QB (\$dummy [71]), 
         .D (nx13711), .CLK (clk), .R (nx17963)) ;
    xnor2 ix1239 (.Y (nx1238), .A0 (nx17819), .A1 (nx16166)) ;
    nand02 ix16167 (.Y (nx16166), .A0 (cache_width_count_1), .A1 (
           cache_width_count_0)) ;
    dffr reg_cache_width_count_3 (.Q (cache_width_count_3), .QB (\$dummy [72]), 
         .D (nx13721), .CLK (clk), .R (nx17963)) ;
    xnor2 ix1247 (.Y (nx1246), .A0 (cache_width_count_3), .A1 (nx16172)) ;
    nand03 ix16173 (.Y (nx16172), .A0 (cache_width_count_1), .A1 (
           cache_width_count_0), .A2 (nx17821)) ;
    dffr reg_cache_width_cntr_counter_out_5 (.Q (cache_width_cntr_counter_out_5)
         , .QB (nx16178), .D (nx13741), .CLK (clk), .R (nx17965)) ;
    oai21 ix16181 (.Y (nx16180), .A0 (nx1260), .A1 (
          cache_width_cntr_counter_out_5), .B0 (nx16131)) ;
    nor02ii ix1261 (.Y (nx1260), .A0 (nx16136), .A1 (nx17817)) ;
    nor04 ix1457 (.Y (nx1456), .A0 (nx1436), .A1 (nx1438), .A2 (nx1446), .A3 (
          nx1448)) ;
    aoi21 ix16190 (.Y (nx16189), .A0 (img_width_out_1), .A1 (img_width_out_0), .B0 (
          nx16191)) ;
    xnor2 ix1439 (.Y (nx1438), .A0 (nx17821), .A1 (nx18055)) ;
    xnor2 ix1447 (.Y (nx1446), .A0 (cache_width_count_3), .A1 (nx16042)) ;
    xnor2 ix1449 (.Y (nx1448), .A0 (nx17817), .A1 (nx16055)) ;
    aoi43 ix16197 (.Y (nx16196), .A0 (nx15563), .A1 (nx17845), .A2 (nx17871), .A3 (
          nx15621), .B0 (nx15561), .B1 (ftc_cntrl_reg_out_11), .B2 (
          current_state_21)) ;
    aoi22 ix16199 (.Y (nx16198), .A0 (nx17921), .A1 (nx15859), .B0 (nx15970), .B1 (
          nx16153)) ;
    dffr ftc_cntrl_reg_reg_q_14 (.Q (ftc_cntrl_reg_out_14), .QB (nx15563), .D (
         nx13071), .CLK (nx17833), .R (nx17807)) ;
    nand02 ix159 (.Y (nx158), .A0 (nx16202), .A1 (nx16204)) ;
    oai21 ix16203 (.Y (nx16202), .A0 (nx17873), .A1 (nx15970), .B0 (nx16065)) ;
    aoi43 ix16205 (.Y (nx16204), .A0 (nx17873), .A1 (nx15621), .A2 (nx15575), .A3 (
          nx15561), .B0 (current_state_21), .B1 (nx15563), .B2 (nx17845)) ;
    dffr reg_current_state_18 (.Q (current_state_18), .QB (\$dummy [73]), .D (
         nx1484), .CLK (nx17835), .R (reset)) ;
    dffr reg_num_channels_counter_out_1 (.Q (num_channels_counter_out_1), .QB (
         \$dummy [74]), .D (nx13931), .CLK (clk), .R (reset)) ;
    mux21_ni ix13932 (.Y (nx13931), .A0 (num_channels_counter_out_1), .A1 (
             nx1648), .S0 (nx17973)) ;
    oai321 ix1649 (.Y (nx1648), .A0 (nx16213), .A1 (nx18265), .A2 (nx18151), .B0 (
           nx148), .B1 (nx16224), .C0 (nx16228)) ;
    dffr max_num_channels_inst_reg_q_1 (.Q (\$dummy [75]), .QB (nx16213), .D (
         nx13921), .CLK (clk), .R (reset)) ;
    oai32 ix13922 (.Y (nx13921), .A0 (nx16213), .A1 (nx17897), .A2 (nx17875), .B0 (
          nx16216), .B1 (nx18259)) ;
    aoi22 ix16217 (.Y (nx16216), .A0 (mem_data_in[1]), .A1 (nx17897), .B0 (
          nx17875), .B1 (nflt_layer_temp_1)) ;
    dffr nflt_layer_total_reg_q_1 (.Q (nflt_layer_temp_1), .QB (\$dummy [76]), .D (
         nx13881), .CLK (clk), .R (reset)) ;
    mux21_ni ix13882 (.Y (nx13881), .A0 (nflt_layer_temp_1), .A1 (mem_data_in[1]
             ), .S0 (nx17895)) ;
    aoi21 ix16225 (.Y (nx16224), .A0 (num_channels_counter_out_1), .A1 (
          num_channels_counter_out_0), .B0 (nx16226)) ;
    aoi22 ix16229 (.Y (nx16228), .A0 (mem_data_in[1]), .A1 (nx17899), .B0 (
          nx17877), .B1 (nflt_layer_temp_1)) ;
    mux21_ni ix13952 (.Y (nx13951), .A0 (num_channels_counter_out_2), .A1 (
             nx1674), .S0 (nx17973)) ;
    oai21 ix1675 (.Y (nx1674), .A0 (nx16234), .A1 (nx18269), .B0 (nx16239)) ;
    aoi22 ix16235 (.Y (nx16234), .A0 (mem_data_in[2]), .A1 (nx17899), .B0 (
          nx17877), .B1 (nflt_layer_temp_2)) ;
    dffr nflt_layer_total_reg_q_2 (.Q (nflt_layer_temp_2), .QB (\$dummy [77]), .D (
         nx13871), .CLK (clk), .R (reset)) ;
    mux21_ni ix13872 (.Y (nx13871), .A0 (nflt_layer_temp_2), .A1 (mem_data_in[2]
             ), .S0 (nx17895)) ;
    aoi22 ix16240 (.Y (nx16239), .A0 (max_num_channels_data_out_2), .A1 (nx1642)
          , .B0 (nx18269), .B1 (nx1660)) ;
    oai32 ix13942 (.Y (nx13941), .A0 (nx16243), .A1 (nx17899), .A2 (nx17877), .B0 (
          nx16234), .B1 (nx18259)) ;
    dffr max_num_channels_inst_reg_q_2 (.Q (max_num_channels_data_out_2), .QB (
         nx16243), .D (nx13941), .CLK (clk), .R (reset)) ;
    nor02_2x ix1643 (.Y (nx1642), .A0 (nx18265), .A1 (nx18151)) ;
    oai21 ix1661 (.Y (nx1660), .A0 (nx16247), .A1 (nx16226), .B0 (nx12908)) ;
    dffr reg_num_channels_counter_out_2 (.Q (num_channels_counter_out_2), .QB (
         nx16247), .D (nx13951), .CLK (clk), .R (reset)) ;
    dffr reg_num_channels_counter_out_3 (.Q (num_channels_counter_out_3), .QB (
         \$dummy [78]), .D (nx13971), .CLK (clk), .R (reset)) ;
    mux21_ni ix13972 (.Y (nx13971), .A0 (num_channels_counter_out_3), .A1 (
             nx1700), .S0 (nx17973)) ;
    oai21 ix1701 (.Y (nx1700), .A0 (nx16253), .A1 (nx18269), .B0 (nx16258)) ;
    aoi22 ix16254 (.Y (nx16253), .A0 (mem_data_in[3]), .A1 (nx17899), .B0 (
          nx17877), .B1 (nflt_layer_temp_3)) ;
    dffr nflt_layer_total_reg_q_3 (.Q (nflt_layer_temp_3), .QB (\$dummy [79]), .D (
         nx13861), .CLK (clk), .R (reset)) ;
    mux21_ni ix13862 (.Y (nx13861), .A0 (nflt_layer_temp_3), .A1 (mem_data_in[3]
             ), .S0 (nx17895)) ;
    aoi22 ix16259 (.Y (nx16258), .A0 (max_num_channels_data_out_3), .A1 (nx1642)
          , .B0 (nx18269), .B1 (nx1686)) ;
    oai32 ix13962 (.Y (nx13961), .A0 (nx16262), .A1 (nx17899), .A2 (nx17877), .B0 (
          nx16253), .B1 (nx18259)) ;
    dffr max_num_channels_inst_reg_q_3 (.Q (max_num_channels_data_out_3), .QB (
         nx16262), .D (nx13961), .CLK (clk), .R (reset)) ;
    xor2 ix1687 (.Y (nx1686), .A0 (num_channels_counter_out_3), .A1 (nx16265)) ;
    nor03_2x ix16266 (.Y (nx16265), .A0 (num_channels_counter_out_0), .A1 (
             num_channels_counter_out_1), .A2 (num_channels_counter_out_2)) ;
    nor03_2x ix16270 (.Y (nx16269), .A0 (nlayers_counter_out_1), .A1 (
             nlayers_counter_out_2), .A2 (nx16278)) ;
    dffr reg_nlayers_counter_out_1 (.Q (nlayers_counter_out_1), .QB (
         \$dummy [80]), .D (nx14011), .CLK (clk), .R (reset)) ;
    mux21_ni ix14012 (.Y (nx14011), .A0 (nx1764), .A1 (nlayers_counter_out_1), .S0 (
             nx16282)) ;
    aoi21 ix16275 (.Y (nx16274), .A0 (nlayers_counter_out_1), .A1 (
          nlayers_counter_out_0), .B0 (nx16284)) ;
    oai32 ix14002 (.Y (nx14001), .A0 (nx16278), .A1 (current_state_2), .A2 (
          nx17877), .B0 (nx16280), .B1 (nx16282)) ;
    dffr reg_nlayers_counter_out_0 (.Q (nlayers_counter_out_0), .QB (nx16278), .D (
         nx14001), .CLK (clk), .R (reset)) ;
    dffr reg_nlayers_counter_out_2 (.Q (nlayers_counter_out_2), .QB (
         \$dummy [81]), .D (nx14021), .CLK (clk), .R (reset)) ;
    mux21_ni ix14022 (.Y (nx14021), .A0 (nx1780), .A1 (nlayers_counter_out_2), .S0 (
             nx16282)) ;
    xnor2 ix16291 (.Y (nx16290), .A0 (nlayers_counter_out_2), .A1 (nx16284)) ;
    inv01 ix16300 (.Y (nx16299), .A (mem_data_in[4])) ;
    oai21 ix1713 (.Y (nx1712), .A0 (nx15426), .A1 (nx15460), .B0 (nx12875)) ;
    dffr reg_current_state_12 (.Q (\$dummy [82]), .QB (nx16302), .D (nx174), .CLK (
         nx17837), .R (reset)) ;
    nand03 ix175 (.Y (nx174), .A0 (nx16305), .A1 (nx15435), .A2 (nx18265)) ;
    oai21 ix16306 (.Y (nx16305), .A0 (nx18151), .A1 (nx15548), .B0 (
          current_state_8)) ;
    oai21 ix16308 (.Y (nx16307), .A0 (cntr1_inst_counter_out_0), .A1 (
          cntr1_inst_counter_out_1), .B0 (nx15412)) ;
    nand02 ix16314 (.Y (nx16313), .A0 (current_state_10), .A1 (nx196)) ;
    nand02 ix1939 (.Y (nx1938), .A0 (nx16318), .A1 (nx18075)) ;
    nand03 ix16319 (.Y (nx16318), .A0 (nx12873), .A1 (nx15486), .A2 (nx16269)) ;
    nor02_2x ix1737 (.Y (nx12873), .A0 (nx12875), .A1 (nx15537)) ;
    dffr reg_current_state_27 (.Q (current_state_27), .QB (nx16327), .D (nx1938)
         , .CLK (nx17837), .R (reset)) ;
    dffr reg_class_cntr_counter_out_0 (.Q (class_cntr_counter_out_0), .QB (
         nx16324), .D (nx14051), .CLK (nx17837), .R (reset)) ;
    dffr reg_class_cntr_counter_out_1 (.Q (class_cntr_counter_out_1), .QB (
         nx16332), .D (nx14061), .CLK (nx17837), .R (reset)) ;
    oai21 ix16335 (.Y (nx16334), .A0 (class_cntr_counter_out_0), .A1 (
          class_cntr_counter_out_1), .B0 (nx16336)) ;
    dffr reg_class_cntr_counter_out_2 (.Q (class_cntr_counter_out_2), .QB (
         nx16338), .D (nx14071), .CLK (nx17837), .R (reset)) ;
    dffr reg_class_cntr_counter_out_3 (.Q (class_cntr_counter_out_3), .QB (
         nx16348), .D (nx14081), .CLK (nx17837), .R (reset)) ;
    dff reg_flt_bias1_reg_q_0 (.Q (flt_bias_out_0), .QB (\$dummy [83]), .D (
        nx14101), .CLK (clk)) ;
    mux21_ni ix14102 (.Y (nx14101), .A0 (flt_bias_out_0), .A1 (mem_data_in[0]), 
             .S0 (nx17993)) ;
    nor02_2x ix2129 (.Y (nx2128), .A0 (nx16302), .A1 (nx18153)) ;
    oai21 ix14092 (.Y (nx14091), .A0 (nx18297), .A1 (nx182), .B0 (nx16302)) ;
    dffr channel_zero_reg_q_0 (.Q (\$dummy [84]), .QB (nx16373), .D (nx14091), .CLK (
         clk), .R (reset)) ;
    dff reg_flt_bias1_reg_q_1 (.Q (flt_bias_out_1), .QB (\$dummy [85]), .D (
        nx14121), .CLK (clk)) ;
    mux21_ni ix14122 (.Y (nx14121), .A0 (flt_bias_out_1), .A1 (mem_data_in[1]), 
             .S0 (nx17993)) ;
    dff reg_flt_bias1_reg_q_2 (.Q (flt_bias_out_2), .QB (\$dummy [86]), .D (
        nx14141), .CLK (clk)) ;
    mux21_ni ix14142 (.Y (nx14141), .A0 (flt_bias_out_2), .A1 (mem_data_in[2]), 
             .S0 (nx17993)) ;
    dff reg_flt_bias1_reg_q_3 (.Q (flt_bias_out_3), .QB (\$dummy [87]), .D (
        nx14161), .CLK (clk)) ;
    mux21_ni ix14162 (.Y (nx14161), .A0 (flt_bias_out_3), .A1 (mem_data_in[3]), 
             .S0 (nx17993)) ;
    dff reg_flt_bias1_reg_q_4 (.Q (flt_bias_out_4), .QB (\$dummy [88]), .D (
        nx14181), .CLK (clk)) ;
    mux21_ni ix14182 (.Y (nx14181), .A0 (flt_bias_out_4), .A1 (mem_data_in[4]), 
             .S0 (nx17993)) ;
    dff reg_flt_bias1_reg_q_5 (.Q (flt_bias_out_5), .QB (\$dummy [89]), .D (
        nx14201), .CLK (clk)) ;
    mux21_ni ix14202 (.Y (nx14201), .A0 (flt_bias_out_5), .A1 (mem_data_in[5]), 
             .S0 (nx17993)) ;
    dff reg_flt_bias1_reg_q_6 (.Q (flt_bias_out_6), .QB (\$dummy [90]), .D (
        nx14221), .CLK (clk)) ;
    mux21_ni ix14222 (.Y (nx14221), .A0 (flt_bias_out_6), .A1 (mem_data_in[6]), 
             .S0 (nx17995)) ;
    dff reg_flt_bias1_reg_q_7 (.Q (flt_bias_out_7), .QB (\$dummy [91]), .D (
        nx14241), .CLK (clk)) ;
    mux21_ni ix14242 (.Y (nx14241), .A0 (flt_bias_out_7), .A1 (mem_data_in[7]), 
             .S0 (nx17995)) ;
    dff reg_flt_bias1_reg_q_8 (.Q (flt_bias_out_8), .QB (\$dummy [92]), .D (
        nx14261), .CLK (clk)) ;
    mux21_ni ix14262 (.Y (nx14261), .A0 (flt_bias_out_8), .A1 (mem_data_in[8]), 
             .S0 (nx17995)) ;
    dff reg_flt_bias1_reg_q_9 (.Q (flt_bias_out_9), .QB (\$dummy [93]), .D (
        nx14281), .CLK (clk)) ;
    mux21_ni ix14282 (.Y (nx14281), .A0 (flt_bias_out_9), .A1 (mem_data_in[9]), 
             .S0 (nx17995)) ;
    dff reg_flt_bias1_reg_q_10 (.Q (flt_bias_out_10), .QB (\$dummy [94]), .D (
        nx14301), .CLK (clk)) ;
    mux21_ni ix14302 (.Y (nx14301), .A0 (flt_bias_out_10), .A1 (mem_data_in[10])
             , .S0 (nx17995)) ;
    dff reg_flt_bias1_reg_q_11 (.Q (flt_bias_out_11), .QB (\$dummy [95]), .D (
        nx14321), .CLK (clk)) ;
    mux21_ni ix14322 (.Y (nx14321), .A0 (flt_bias_out_11), .A1 (mem_data_in[11])
             , .S0 (nx17995)) ;
    dff reg_flt_bias1_reg_q_12 (.Q (flt_bias_out_12), .QB (\$dummy [96]), .D (
        nx14341), .CLK (clk)) ;
    mux21_ni ix14342 (.Y (nx14341), .A0 (flt_bias_out_12), .A1 (mem_data_in[12])
             , .S0 (nx2128)) ;
    dff reg_flt_bias1_reg_q_13 (.Q (flt_bias_out_13), .QB (\$dummy [97]), .D (
        nx14361), .CLK (clk)) ;
    mux21_ni ix14362 (.Y (nx14361), .A0 (flt_bias_out_13), .A1 (mem_data_in[13])
             , .S0 (nx2128)) ;
    dff reg_flt_bias1_reg_q_14 (.Q (flt_bias_out_14), .QB (\$dummy [98]), .D (
        nx14381), .CLK (clk)) ;
    mux21_ni ix14382 (.Y (nx14381), .A0 (flt_bias_out_14), .A1 (mem_data_in[14])
             , .S0 (nx2128)) ;
    dff reg_flt_bias1_reg_q_15 (.Q (flt_bias_out_15), .QB (\$dummy [99]), .D (
        nx14401), .CLK (clk)) ;
    mux21_ni ix14402 (.Y (nx14401), .A0 (flt_bias_out_15), .A1 (mem_data_in[15])
             , .S0 (nx2128)) ;
    nor03_2x ix5153 (.Y (max_height_3), .A0 (nx16042), .A1 (nx17807), .A2 (
             nx17923)) ;
    nor03_2x ix5157 (.Y (max_height_4), .A0 (nx16055), .A1 (nx17807), .A2 (
             nx17923)) ;
    or02 ix4861 (.Y (cache_rst_actual), .A0 (nx17809), .A1 (reset)) ;
    nand02 ix2619 (.Y (cache_load), .A0 (nx16455), .A1 (nx18081)) ;
    mux21 ix14422 (.Y (nx14421), .A0 (nx16459), .A1 (nx16463), .S0 (nx18047)) ;
    aoi32 ix16460 (.Y (nx16459), .A0 (nx1460), .A1 (cache_height_ended), .A2 (
          nx17873), .B0 (ftc_cntrl_reg_out_15), .B1 (nx2566)) ;
    nand03 ix2567 (.Y (nx2566), .A0 (ftc_cntrl_reg_out_13), .A1 (nx15605), .A2 (
           nx17923)) ;
    dffr ftc_cntrl_reg_reg_q_15 (.Q (ftc_cntrl_reg_out_15), .QB (nx16463), .D (
         nx14421), .CLK (nx17839), .R (nx17809)) ;
    nor03_2x ix1183 (.Y (nx1182), .A0 (ftc_cntrl_reg_out_12), .A1 (nx18279), .A2 (
             ftc_cntrl_reg_out_13)) ;
    nand02 ix5143 (.Y (max_height_0), .A0 (nx16507), .A1 (img_width_out_0)) ;
    nand02 ix5149 (.Y (max_height_2), .A0 (nx16507), .A1 (nx18055)) ;
    oai21 ix2153 (.Y (comp_unit_data1_out[0]), .A0 (nx18063), .A1 (nx16511), .B0 (
          nx16514)) ;
    dffr bias1_reg_reg_q_0 (.Q (\$dummy [100]), .QB (nx16511), .D (nx14111), .CLK (
         clk), .R (reset)) ;
    nand02 ix16515 (.Y (nx16514), .A0 (nx2140), .A1 (nx17997)) ;
    oai21 ix2179 (.Y (comp_unit_data1_out[1]), .A0 (nx18063), .A1 (nx16518), .B0 (
          nx16521)) ;
    dffr bias1_reg_reg_q_1 (.Q (\$dummy [101]), .QB (nx16518), .D (nx14131), .CLK (
         clk), .R (reset)) ;
    nand02 ix16522 (.Y (nx16521), .A0 (nx2168), .A1 (nx17997)) ;
    oai21 ix2205 (.Y (comp_unit_data1_out[2]), .A0 (nx18063), .A1 (nx16524), .B0 (
          nx16527)) ;
    dffr bias1_reg_reg_q_2 (.Q (\$dummy [102]), .QB (nx16524), .D (nx14151), .CLK (
         clk), .R (reset)) ;
    nand02 ix16528 (.Y (nx16527), .A0 (nx2194), .A1 (nx17997)) ;
    oai21 ix2231 (.Y (comp_unit_data1_out[3]), .A0 (nx18063), .A1 (nx16530), .B0 (
          nx16533)) ;
    dffr bias1_reg_reg_q_3 (.Q (\$dummy [103]), .QB (nx16530), .D (nx14171), .CLK (
         clk), .R (reset)) ;
    nand02 ix16534 (.Y (nx16533), .A0 (nx2220), .A1 (nx17997)) ;
    oai21 ix2257 (.Y (comp_unit_data1_out[4]), .A0 (nx18065), .A1 (nx16536), .B0 (
          nx16539)) ;
    dffr bias1_reg_reg_q_4 (.Q (\$dummy [104]), .QB (nx16536), .D (nx14191), .CLK (
         clk), .R (reset)) ;
    nand02 ix16540 (.Y (nx16539), .A0 (nx2246), .A1 (nx17997)) ;
    oai21 ix2283 (.Y (comp_unit_data1_out[5]), .A0 (nx18065), .A1 (nx16542), .B0 (
          nx16545)) ;
    dffr bias1_reg_reg_q_5 (.Q (\$dummy [105]), .QB (nx16542), .D (nx14211), .CLK (
         clk), .R (reset)) ;
    nand02 ix16546 (.Y (nx16545), .A0 (nx2272), .A1 (nx17997)) ;
    oai21 ix2309 (.Y (comp_unit_data1_out[6]), .A0 (nx18065), .A1 (nx16548), .B0 (
          nx16551)) ;
    dffr bias1_reg_reg_q_6 (.Q (\$dummy [106]), .QB (nx16548), .D (nx14231), .CLK (
         clk), .R (reset)) ;
    nand02 ix16552 (.Y (nx16551), .A0 (nx2298), .A1 (nx17997)) ;
    oai21 ix2335 (.Y (comp_unit_data1_out[7]), .A0 (nx18065), .A1 (nx16554), .B0 (
          nx16557)) ;
    dffr bias1_reg_reg_q_7 (.Q (\$dummy [107]), .QB (nx16554), .D (nx14251), .CLK (
         clk), .R (reset)) ;
    nand02 ix16558 (.Y (nx16557), .A0 (nx2324), .A1 (nx17999)) ;
    oai21 ix2361 (.Y (comp_unit_data1_out[8]), .A0 (nx18065), .A1 (nx16560), .B0 (
          nx16563)) ;
    dffr bias1_reg_reg_q_8 (.Q (\$dummy [108]), .QB (nx16560), .D (nx14271), .CLK (
         clk), .R (reset)) ;
    nand02 ix16564 (.Y (nx16563), .A0 (nx2350), .A1 (nx17999)) ;
    oai21 ix2387 (.Y (comp_unit_data1_out[9]), .A0 (nx18065), .A1 (nx16566), .B0 (
          nx16569)) ;
    dffr bias1_reg_reg_q_9 (.Q (\$dummy [109]), .QB (nx16566), .D (nx14291), .CLK (
         clk), .R (reset)) ;
    nand02 ix16570 (.Y (nx16569), .A0 (nx2376), .A1 (nx17999)) ;
    oai21 ix2413 (.Y (comp_unit_data1_out[10]), .A0 (nx18067), .A1 (nx16572), .B0 (
          nx16575)) ;
    dffr bias1_reg_reg_q_10 (.Q (\$dummy [110]), .QB (nx16572), .D (nx14311), .CLK (
         clk), .R (reset)) ;
    nand02 ix16576 (.Y (nx16575), .A0 (nx2402), .A1 (nx17999)) ;
    oai21 ix2439 (.Y (comp_unit_data1_out[11]), .A0 (nx18067), .A1 (nx16578), .B0 (
          nx16581)) ;
    dffr bias1_reg_reg_q_11 (.Q (\$dummy [111]), .QB (nx16578), .D (nx14331), .CLK (
         clk), .R (reset)) ;
    nand02 ix16582 (.Y (nx16581), .A0 (nx2428), .A1 (nx17999)) ;
    oai21 ix2465 (.Y (comp_unit_data1_out[12]), .A0 (nx18067), .A1 (nx16584), .B0 (
          nx16587)) ;
    dffr bias1_reg_reg_q_12 (.Q (\$dummy [112]), .QB (nx16584), .D (nx14351), .CLK (
         clk), .R (reset)) ;
    nand02 ix16588 (.Y (nx16587), .A0 (nx2454), .A1 (nx17999)) ;
    oai21 ix2491 (.Y (comp_unit_data1_out[13]), .A0 (nx18067), .A1 (nx16590), .B0 (
          nx16593)) ;
    dffr bias1_reg_reg_q_13 (.Q (\$dummy [113]), .QB (nx16590), .D (nx14371), .CLK (
         clk), .R (reset)) ;
    nand02 ix16594 (.Y (nx16593), .A0 (nx2480), .A1 (nx17999)) ;
    oai21 ix2517 (.Y (comp_unit_data1_out[14]), .A0 (nx18067), .A1 (nx16596), .B0 (
          nx16599)) ;
    dffr bias1_reg_reg_q_14 (.Q (\$dummy [114]), .QB (nx16596), .D (nx14391), .CLK (
         clk), .R (reset)) ;
    nand02 ix16600 (.Y (nx16599), .A0 (nx2506), .A1 (nx18001)) ;
    oai21 ix2543 (.Y (comp_unit_data1_out[15]), .A0 (nx18067), .A1 (nx16602), .B0 (
          nx16605)) ;
    dffr bias1_reg_reg_q_15 (.Q (\$dummy [115]), .QB (nx16602), .D (nx14411), .CLK (
         clk), .R (reset)) ;
    nand02 ix16606 (.Y (nx16605), .A0 (nx2532), .A1 (nx18001)) ;
    oai21 ix2117 (.Y (comp_unit_ready), .A0 (nx18273), .A1 (nx196), .B0 (nx16608
          )) ;
    aoi21 ix16609 (.Y (nx16608), .A0 (nx17971), .A1 (nx18305), .B0 (nx18233)) ;
    nand03 ix16611 (.Y (nx16610), .A0 (flt_size_out_0), .A1 (nx15711), .A2 (
           flt_size_out_1)) ;
    aoi21 ix4883 (.Y (mem_read_out), .A0 (nx16715), .A1 (nx16721), .B0 (reset)
          ) ;
    nor04 ix16722 (.Y (nx16721), .A0 (nx18003), .A1 (nx17869), .A2 (nx2754), .A3 (
          nx2128)) ;
    nand02 ix2755 (.Y (nx2754), .A0 (nx16727), .A1 (nx16729)) ;
    nor04 ix16728 (.Y (nx16727), .A0 (current_state_2), .A1 (current_state_3), .A2 (
          nx17895), .A3 (current_state_5)) ;
    nor04 ix16730 (.Y (nx16729), .A0 (current_state_6), .A1 (nx17907), .A2 (
          current_state_8), .A3 (nx17899)) ;
    aoi21 ix4867 (.Y (mem_write_out), .A0 (nx18053), .A1 (nx18883), .B0 (reset)
          ) ;
    dffr reg_current_state_28 (.Q (\$dummy [116]), .QB (nx16732), .D (nx1946), .CLK (
         nx17839), .R (reset)) ;
    nand04 ix2779 (.Y (mem_addr_out[0]), .A0 (nx16736), .A1 (nx16756), .A2 (
           nx16780), .A3 (nx16788)) ;
    aoi221 ix16737 (.Y (nx16736), .A0 (nx16738), .A1 (nx17855), .B0 (
           addr1_data_0), .B1 (nx18037), .C0 (nx2740)) ;
    oai21 ix16739 (.Y (nx16738), .A0 (class_cntr_counter_out_0), .A1 (nx18007), 
          .B0 (nx16747)) ;
    oai33 ix14432 (.Y (nx14431), .A0 (nx16742), .A1 (nx2622), .A2 (nx18069), .B0 (
          nx16745), .B1 (nx17887), .B2 (nx17879)) ;
    dffr reg_write_base_reg_q_0 (.Q (\$dummy [117]), .QB (nx16745), .D (nx14431)
         , .CLK (nx17839), .R (reset)) ;
    dffr reg_addr1_data_0 (.Q (addr1_data_0), .QB (\$dummy [118]), .D (nx14481)
         , .CLK (clk), .R (reset)) ;
    nand02 ix2767 (.Y (nx2766), .A0 (nx16313), .A1 (nx18121)) ;
    nor02_2x ix2741 (.Y (nx2740), .A0 (nx18883), .A1 (nx16738)) ;
    oai21 ix16757 (.Y (nx16756), .A0 (img_addr_offset_0), .A1 (img_base_addr_0)
          , .B0 (nx2724)) ;
    dffr reg_img_addr_offset_0 (.Q (img_addr_offset_0), .QB (\$dummy [119]), .D (
         nx14471), .CLK (clk), .R (nx18031)) ;
    or02 ix2713 (.Y (nx2712), .A0 (nx12873), .A1 (reset)) ;
    dffs_ni img_base_addr_inst_reg_q_0 (.Q (img_base_addr_0), .QB (\$dummy [120]
            ), .D (nx14461), .CLK (clk), .S (reset)) ;
    dffr reg_write_base_prev_reg_q_0 (.Q (write_base_prev_data_out_0), .QB (
         nx16764), .D (nx14451), .CLK (clk), .R (reset)) ;
    nand04 ix16769 (.Y (nx16768), .A0 (nx16770), .A1 (nx2678), .A2 (nx16774), .A3 (
           nx16776)) ;
    nor02_2x ix2679 (.Y (nx2678), .A0 (nx16302), .A1 (nx2674)) ;
    xnor2 ix16777 (.Y (nx16776), .A0 (nflt_layer_temp_3), .A1 (nflt_layer_out_3)
          ) ;
    aoi21 ix2725 (.Y (nx2724), .A0 (img_base_addr_0), .A1 (img_addr_offset_0), .B0 (
          nx18085)) ;
    oai21 ix16781 (.Y (nx16780), .A0 (nx18007), .A1 (bias_offset_data_out_0), .B0 (
          nx2668)) ;
    dffr reg_bias_offset_reg_q_0 (.Q (bias_offset_data_out_0), .QB (
         \$dummy [121]), .D (nx14441), .CLK (clk), .R (reset)) ;
    aoi21 ix2669 (.Y (nx2668), .A0 (bias_offset_data_out_0), .A1 (nx18007), .B0 (
          nx18135)) ;
    nand02 ix16787 (.Y (nx16786), .A0 (nx18233), .A1 (nx18297)) ;
    oai221 ix16789 (.Y (nx16788), .A0 (nx18011), .A1 (nx18229), .B0 (
           write_offset_data_out_0), .B1 (nx18007), .C0 (nx16791)) ;
    or02 ix2885 (.Y (mem_addr_out[1]), .A0 (nx2882), .A1 (nx2822)) ;
    oai222 ix2883 (.Y (nx2882), .A0 (nx2874), .A1 (nx18075), .B0 (nx16810), .B1 (
           nx18085), .C0 (nx16835), .C1 (nx18135)) ;
    nand02 ix2875 (.Y (nx2874), .A0 (nx16796), .A1 (nx16738)) ;
    xnor2 ix16797 (.Y (nx16796), .A0 (nx16747), .A1 (nx16798)) ;
    dffr reg_write_base_reg_q_1 (.Q (write_base_data_out_1), .QB (nx16802), .D (
         nx14491), .CLK (nx17839), .R (reset)) ;
    xnor2 ix16805 (.Y (nx16804), .A0 (nx16806), .A1 (nx16808)) ;
    nand02 ix16807 (.Y (nx16806), .A0 (new_size_squared_out_0), .A1 (nx18009)) ;
    xnor2 ix16811 (.Y (nx16810), .A0 (nx16812), .A1 (nx16814)) ;
    nand02 ix16813 (.Y (nx16812), .A0 (img_base_addr_0), .A1 (img_addr_offset_0)
           ) ;
    dffs_ni img_base_addr_inst_reg_q_1 (.Q (img_base_addr_1), .QB (nx16818), .D (
            nx14521), .CLK (clk), .S (reset)) ;
    aoi21 ix16821 (.Y (nx16820), .A0 (write_base_prev_data_out_1), .A1 (
          write_base_prev_data_out_0), .B0 (nx16825)) ;
    dffr reg_write_base_prev_reg_q_1 (.Q (write_base_prev_data_out_1), .QB (
         \$dummy [122]), .D (nx14511), .CLK (clk), .R (reset)) ;
    oai21 ix16830 (.Y (nx16829), .A0 (img_addr_offset_0), .A1 (img_addr_offset_1
          ), .B0 (nx16831)) ;
    nand02 ix16832 (.Y (nx16831), .A0 (img_addr_offset_1), .A1 (
           img_addr_offset_0)) ;
    dffr reg_img_addr_offset_1 (.Q (img_addr_offset_1), .QB (nx16833), .D (
         nx14531), .CLK (clk), .R (nx18031)) ;
    xnor2 ix16836 (.Y (nx16835), .A0 (nx16837), .A1 (nx16839)) ;
    nand02 ix16838 (.Y (nx16837), .A0 (bias_offset_data_out_0), .A1 (nx18009)) ;
    dffr reg_bias_offset_reg_q_1 (.Q (bias_offset_data_out_1), .QB (nx16843), .D (
         nx14541), .CLK (clk), .R (reset)) ;
    oai222 ix2823 (.Y (nx2822), .A0 (nx16846), .A1 (nx18139), .B0 (nx16796), .B1 (
           nx16857), .C0 (nx16861), .C1 (nx18143)) ;
    oai21 ix16850 (.Y (nx16849), .A0 (addr1_data_0), .A1 (addr1_data_1), .B0 (
          nx16852)) ;
    dffr reg_addr1_data_1 (.Q (addr1_data_1), .QB (nx16846), .D (nx14501), .CLK (
         clk), .R (reset)) ;
    nand02 ix16853 (.Y (nx16852), .A0 (addr1_data_1), .A1 (addr1_data_0)) ;
    aoi21 ix16858 (.Y (nx16857), .A0 (nx2738), .A1 (nx17855), .B0 (nx17975)) ;
    xnor2 ix16862 (.Y (nx16861), .A0 (nx16791), .A1 (nx16863)) ;
    nand02 ix3031 (.Y (mem_addr_out[2]), .A0 (nx16868), .A1 (nx16916)) ;
    aoi222 ix16869 (.Y (nx16868), .A0 (nx16870), .A1 (nx17855), .B0 (nx3016), .B1 (
           nx18021), .C0 (nx2996), .C1 (nx18003)) ;
    nor02_2x ix16871 (.Y (nx16870), .A0 (nx2928), .A1 (nx2874)) ;
    xnor2 ix2929 (.Y (nx2928), .A0 (nx2924), .A1 (nx16874)) ;
    oai22 ix2925 (.Y (nx2924), .A0 (nx16747), .A1 (nx16798), .B0 (nx16332), .B1 (
          nx16802)) ;
    dffr reg_write_base_reg_q_2 (.Q (write_base_data_out_2), .QB (nx16878), .D (
         nx14551), .CLK (nx17839), .R (reset)) ;
    xnor2 ix16881 (.Y (nx16880), .A0 (nx16882), .A1 (nx16885)) ;
    xor2 ix3017 (.Y (nx3016), .A0 (nx16888), .A1 (nx16891)) ;
    dffr reg_bias_offset_reg_q_2 (.Q (bias_offset_data_out_2), .QB (nx16895), .D (
         nx14601), .CLK (clk), .R (reset)) ;
    xor2 ix2997 (.Y (nx2996), .A0 (nx16898), .A1 (nx16901)) ;
    dffs_ni img_base_addr_inst_reg_q_2 (.Q (img_base_addr_2), .QB (nx16911), .D (
            nx14581), .CLK (clk), .S (reset)) ;
    oai21 ix2975 (.Y (nx2974), .A0 (nx16906), .A1 (nx16825), .B0 (nx2968)) ;
    dffr reg_write_base_prev_reg_q_2 (.Q (write_base_prev_data_out_2), .QB (
         nx16906), .D (nx14571), .CLK (clk), .R (reset)) ;
    dffr reg_img_addr_offset_2 (.Q (img_addr_offset_2), .QB (nx16915), .D (
         nx14591), .CLK (clk), .R (nx18031)) ;
    aoi222 ix16917 (.Y (nx16916), .A0 (addr1_data_2), .A1 (nx18037), .B0 (nx2914
           ), .B1 (nx18017), .C0 (nx2928), .C1 (nx2932)) ;
    dffr reg_addr1_data_2 (.Q (addr1_data_2), .QB (\$dummy [123]), .D (nx14561)
         , .CLK (clk), .R (reset)) ;
    xnor2 ix2943 (.Y (nx2942), .A0 (addr1_data_2), .A1 (nx16852)) ;
    xnor2 ix2915 (.Y (nx2914), .A0 (nx2892), .A1 (nx16924)) ;
    oai22 ix2893 (.Y (nx2892), .A0 (nx16791), .A1 (nx16863), .B0 (nx15756), .B1 (
          nx16802)) ;
    nand02 ix2643 (.Y (nx2642), .A0 (nx18313), .A1 (nx18053)) ;
    nand02 ix3177 (.Y (mem_addr_out[3]), .A0 (nx16931), .A1 (nx16973)) ;
    aoi222 ix16932 (.Y (nx16931), .A0 (nx17975), .A1 (nx3074), .B0 (nx3168), .B1 (
           nx18003), .C0 (nx3122), .C1 (nx18021)) ;
    aoi22 ix16935 (.Y (nx16934), .A0 (class_cntr_counter_out_2), .A1 (
          write_base_data_out_2), .B0 (nx2924), .B1 (nx2926)) ;
    dffs_ni reg_write_base_reg_q_3 (.Q (write_base_data_out_3), .QB (nx16945), .D (
            nx14611), .CLK (nx17839), .S (reset)) ;
    xnor2 ix3051 (.Y (nx3050), .A0 (nx3046), .A1 (nx16943)) ;
    xnor2 ix3169 (.Y (nx3168), .A0 (nx3132), .A1 (nx16948)) ;
    xnor2 ix16949 (.Y (nx16948), .A0 (img_base_addr_3), .A1 (img_addr_offset_3)
          ) ;
    dffr img_base_addr_inst_reg_q_3 (.Q (img_base_addr_3), .QB (\$dummy [124]), 
         .D (nx14651), .CLK (clk), .R (reset)) ;
    xor2 ix3147 (.Y (nx3146), .A0 (write_base_prev_data_out_3), .A1 (nx16956)) ;
    dffr reg_write_base_prev_reg_q_3 (.Q (write_base_prev_data_out_3), .QB (
         \$dummy [125]), .D (nx14641), .CLK (clk), .R (reset)) ;
    nor03_2x ix16957 (.Y (nx16956), .A0 (write_base_prev_data_out_0), .A1 (
             write_base_prev_data_out_1), .A2 (write_base_prev_data_out_2)) ;
    dffr reg_img_addr_offset_3 (.Q (img_addr_offset_3), .QB (\$dummy [126]), .D (
         nx14661), .CLK (clk), .R (nx18031)) ;
    xnor2 ix3161 (.Y (nx3160), .A0 (img_addr_offset_3), .A1 (nx16962)) ;
    nand03 ix16963 (.Y (nx16962), .A0 (img_addr_offset_2), .A1 (
           img_addr_offset_1), .A2 (nx18027)) ;
    xnor2 ix3123 (.Y (nx3122), .A0 (nx3112), .A1 (nx16967)) ;
    dffr reg_bias_offset_reg_q_3 (.Q (bias_offset_data_out_3), .QB (
         \$dummy [127]), .D (nx14631), .CLK (clk), .R (reset)) ;
    aoi322 ix16974 (.Y (nx16973), .A0 (nx3076), .A1 (nx16978), .A2 (nx17855), .B0 (
           addr1_data_3), .B1 (nx18037), .C0 (nx3060), .C1 (nx18017)) ;
    nand02 ix3077 (.Y (nx3076), .A0 (nx16976), .A1 (nx16870)) ;
    xnor2 ix16977 (.Y (nx16976), .A0 (nx16934), .A1 (nx16937)) ;
    dffr reg_addr1_data_3 (.Q (addr1_data_3), .QB (\$dummy [128]), .D (nx14621)
         , .CLK (clk), .R (reset)) ;
    xnor2 ix3093 (.Y (nx3092), .A0 (addr1_data_3), .A1 (nx16983)) ;
    nand03 ix16984 (.Y (nx16983), .A0 (addr1_data_2), .A1 (addr1_data_1), .A2 (
           addr1_data_0)) ;
    xor2 ix3061 (.Y (nx3060), .A0 (nx16987), .A1 (nx16990)) ;
    nand02 ix3327 (.Y (mem_addr_out[4]), .A0 (nx16993), .A1 (nx17047)) ;
    aoi222 ix16994 (.Y (nx16993), .A0 (nx16995), .A1 (nx17855), .B0 (nx3312), .B1 (
           nx18021), .C0 (nx3292), .C1 (nx18003)) ;
    nor02_2x ix3079 (.Y (nx3078), .A0 (nx16870), .A1 (nx16976)) ;
    dffr reg_write_base_reg_q_4 (.Q (write_base_data_out_4), .QB (nx17002), .D (
         nx14671), .CLK (nx17839), .R (reset)) ;
    xnor2 ix17005 (.Y (nx17004), .A0 (nx17006), .A1 (nx17009)) ;
    xor2 ix3313 (.Y (nx3312), .A0 (nx17013), .A1 (nx17016)) ;
    dffr reg_bias_offset_reg_q_4 (.Q (bias_offset_data_out_4), .QB (nx17021), .D (
         nx14721), .CLK (clk), .R (reset)) ;
    aoi21 ix859 (.Y (nx858), .A0 (nx15741), .A1 (nx15735), .B0 (nx852)) ;
    xor2 ix3293 (.Y (nx3292), .A0 (nx17023), .A1 (nx17026)) ;
    dffs_ni img_base_addr_inst_reg_q_4 (.Q (img_base_addr_4), .QB (nx17038), .D (
            nx14701), .CLK (clk), .S (reset)) ;
    oai21 ix3271 (.Y (nx3270), .A0 (nx17031), .A1 (nx17035), .B0 (nx3264)) ;
    dffr reg_write_base_prev_reg_q_4 (.Q (\$dummy [129]), .QB (nx17031), .D (
         nx14691), .CLK (clk), .R (reset)) ;
    nor04 ix17036 (.Y (nx17035), .A0 (write_base_prev_data_out_0), .A1 (
          write_base_prev_data_out_1), .A2 (write_base_prev_data_out_2), .A3 (
          write_base_prev_data_out_3)) ;
    nand02 ix3265 (.Y (nx3264), .A0 (nx17035), .A1 (nx17031)) ;
    aoi21 ix3285 (.Y (nx3284), .A0 (nx17042), .A1 (nx17044), .B0 (nx3278)) ;
    nand04 ix17043 (.Y (nx17042), .A0 (img_addr_offset_3), .A1 (
           img_addr_offset_2), .A2 (img_addr_offset_1), .A3 (nx18027)) ;
    dffr reg_img_addr_offset_4 (.Q (img_addr_offset_4), .QB (nx17044), .D (
         nx14711), .CLK (clk), .R (nx18031)) ;
    aoi21 ix17048 (.Y (nx17047), .A0 (nx3206), .A1 (nx18017), .B0 (nx3246)) ;
    xnor2 ix3207 (.Y (nx3206), .A0 (nx3184), .A1 (nx17051)) ;
    oai22 ix3247 (.Y (nx3246), .A0 (nx16998), .A1 (nx17054), .B0 (nx17056), .B1 (
          nx18139)) ;
    aoi21 ix17055 (.Y (nx17054), .A0 (nx3078), .A1 (nx17855), .B0 (nx17975)) ;
    aoi21 ix3239 (.Y (nx3238), .A0 (nx17060), .A1 (nx17056), .B0 (nx3232)) ;
    nand04 ix17061 (.Y (nx17060), .A0 (addr1_data_3), .A1 (addr1_data_2), .A2 (
           addr1_data_1), .A3 (addr1_data_0)) ;
    dffr reg_addr1_data_4 (.Q (addr1_data_4), .QB (nx17056), .D (nx14681), .CLK (
         clk), .R (reset)) ;
    nand02 ix3469 (.Y (mem_addr_out[5]), .A0 (nx17065), .A1 (nx17106)) ;
    aoi222 ix17066 (.Y (nx17065), .A0 (nx18543), .A1 (nx17857), .B0 (nx3454), .B1 (
           nx18021), .C0 (nx3434), .C1 (nx18003)) ;
    dffs_ni reg_write_base_reg_q_5 (.Q (write_base_data_out_5), .QB (nx17076), .D (
            nx14731), .CLK (nx17841), .S (reset)) ;
    xnor2 ix3347 (.Y (nx3346), .A0 (nx3342), .A1 (nx17074)) ;
    nand02 ix17078 (.Y (nx17077), .A0 (write_base_data_out_4), .A1 (nx3216)) ;
    xnor2 ix3455 (.Y (nx3454), .A0 (nx3444), .A1 (nx17081)) ;
    dffr reg_bias_offset_reg_q_5 (.Q (bias_offset_data_out_5), .QB (nx17085), .D (
         nx14781), .CLK (clk), .R (reset)) ;
    xnor2 ix3435 (.Y (nx3434), .A0 (nx3398), .A1 (nx17089)) ;
    dffr img_base_addr_inst_reg_q_5 (.Q (img_base_addr_5), .QB (\$dummy [130]), 
         .D (nx14761), .CLK (clk), .R (reset)) ;
    xnor2 ix3413 (.Y (nx3412), .A0 (write_base_prev_data_out_5), .A1 (nx3264)) ;
    dffr reg_write_base_prev_reg_q_5 (.Q (write_base_prev_data_out_5), .QB (
         \$dummy [131]), .D (nx14751), .CLK (clk), .R (reset)) ;
    oai21 ix17101 (.Y (nx17100), .A0 (nx3278), .A1 (img_addr_offset_5), .B0 (
          nx17102)) ;
    nand02 ix17103 (.Y (nx17102), .A0 (img_addr_offset_5), .A1 (nx3278)) ;
    dffr reg_img_addr_offset_5 (.Q (img_addr_offset_5), .QB (nx17104), .D (
         nx14771), .CLK (clk), .R (nx18031)) ;
    aoi222 ix17107 (.Y (nx17106), .A0 (addr1_data_5), .A1 (nx18037), .B0 (nx3366
           ), .B1 (nx3370), .C0 (nx3356), .C1 (nx18017)) ;
    oai21 ix17111 (.Y (nx17110), .A0 (nx3232), .A1 (addr1_data_5), .B0 (nx17112)
          ) ;
    nand02 ix17113 (.Y (nx17112), .A0 (addr1_data_5), .A1 (nx3232)) ;
    dffr reg_addr1_data_5 (.Q (addr1_data_5), .QB (nx17114), .D (nx14741), .CLK (
         clk), .R (reset)) ;
    oai21 ix3371 (.Y (nx3370), .A0 (nx16995), .A1 (nx18075), .B0 (nx18883)) ;
    xor2 ix3357 (.Y (nx3356), .A0 (nx17118), .A1 (nx17121)) ;
    or02 ix3611 (.Y (mem_addr_out[6]), .A0 (nx3608), .A1 (nx3532)) ;
    oai222 ix3609 (.Y (nx3608), .A0 (nx17125), .A1 (nx18135), .B0 (nx17147), .B1 (
           nx18087), .C0 (nx3600), .C1 (nx18075)) ;
    xnor2 ix17126 (.Y (nx17125), .A0 (nx17127), .A1 (nx17130)) ;
    dffr reg_bias_offset_reg_q_6 (.Q (bias_offset_data_out_6), .QB (nx17135), .D (
         nx14841), .CLK (clk), .R (reset)) ;
    aoi21 ix905 (.Y (nx904), .A0 (nx15726), .A1 (nx15720), .B0 (nx898)) ;
    dffs_ni reg_write_base_reg_q_6 (.Q (write_base_data_out_6), .QB (nx17138), .D (
            nx14791), .CLK (nx17841), .S (reset)) ;
    xnor2 ix17141 (.Y (nx17140), .A0 (nx17142), .A1 (nx17145)) ;
    xnor2 ix17148 (.Y (nx17147), .A0 (nx17149), .A1 (nx17152)) ;
    dffs_ni img_base_addr_inst_reg_q_6 (.Q (img_base_addr_6), .QB (nx17164), .D (
            nx14821), .CLK (clk), .S (reset)) ;
    oai21 ix3555 (.Y (nx3554), .A0 (nx17157), .A1 (nx17161), .B0 (nx3548)) ;
    dffr reg_write_base_prev_reg_q_6 (.Q (\$dummy [132]), .QB (nx17157), .D (
         nx14811), .CLK (clk), .R (reset)) ;
    nor02_2x ix17162 (.Y (nx17161), .A0 (nx3264), .A1 (
             write_base_prev_data_out_5)) ;
    nand02 ix3549 (.Y (nx3548), .A0 (nx17161), .A1 (nx17157)) ;
    aoi21 ix3569 (.Y (nx3568), .A0 (nx17102), .A1 (nx17168), .B0 (nx3562)) ;
    dffr reg_img_addr_offset_6 (.Q (img_addr_offset_6), .QB (nx17168), .D (
         nx14831), .CLK (clk), .R (nx18031)) ;
    nand02 ix17176 (.Y (nx17175), .A0 (write_base_data_out_6), .A1 (nx3360)) ;
    oai222 ix3533 (.Y (nx3532), .A0 (nx17172), .A1 (nx17178), .B0 (nx17183), .B1 (
           nx18143), .C0 (nx17188), .C1 (nx18139)) ;
    aoi21 ix17179 (.Y (nx17178), .A0 (nx3458), .A1 (nx17857), .B0 (nx17975)) ;
    xor2 ix17184 (.Y (nx17183), .A0 (nx18597), .A1 (nx17186)) ;
    dffr reg_addr1_data_6 (.Q (addr1_data_6), .QB (nx17188), .D (nx14801), .CLK (
         clk), .R (reset)) ;
    nand02 ix3753 (.Y (mem_addr_out[7]), .A0 (nx17194), .A1 (nx17235)) ;
    aoi222 ix17195 (.Y (nx17194), .A0 (nx17196), .A1 (nx17857), .B0 (nx3738), .B1 (
           nx18021), .C0 (nx3718), .C1 (nx18003)) ;
    xnor2 ix3631 (.Y (nx3630), .A0 (nx3626), .A1 (nx17204)) ;
    dffr reg_write_base_reg_q_7 (.Q (write_base_data_out_7), .QB (nx17199), .D (
         nx14851), .CLK (nx17841), .R (reset)) ;
    xnor2 ix3739 (.Y (nx3738), .A0 (nx3728), .A1 (nx17210)) ;
    dffr reg_bias_offset_reg_q_7 (.Q (bias_offset_data_out_7), .QB (nx17214), .D (
         nx14901), .CLK (clk), .R (reset)) ;
    xnor2 ix3719 (.Y (nx3718), .A0 (nx18760), .A1 (nx17218)) ;
    dffr img_base_addr_inst_reg_q_7 (.Q (img_base_addr_7), .QB (\$dummy [133]), 
         .D (nx14881), .CLK (clk), .R (reset)) ;
    xnor2 ix3697 (.Y (nx3696), .A0 (write_base_prev_data_out_7), .A1 (nx3548)) ;
    dffr reg_write_base_prev_reg_q_7 (.Q (write_base_prev_data_out_7), .QB (
         \$dummy [134]), .D (nx14871), .CLK (clk), .R (reset)) ;
    oai21 ix17230 (.Y (nx17229), .A0 (nx3562), .A1 (img_addr_offset_7), .B0 (
          nx17231)) ;
    nand02 ix17232 (.Y (nx17231), .A0 (img_addr_offset_7), .A1 (nx3562)) ;
    dffr reg_img_addr_offset_7 (.Q (img_addr_offset_7), .QB (nx17233), .D (
         nx14891), .CLK (clk), .R (nx18033)) ;
    aoi222 ix17236 (.Y (nx17235), .A0 (addr1_data_7), .A1 (nx18037), .B0 (nx3640
           ), .B1 (nx18017), .C0 (nx3650), .C1 (nx3654)) ;
    oai21 ix17240 (.Y (nx17239), .A0 (nx3516), .A1 (addr1_data_7), .B0 (nx17242)
          ) ;
    nand02 ix17243 (.Y (nx17242), .A0 (addr1_data_7), .A1 (nx3516)) ;
    dffr reg_addr1_data_7 (.Q (addr1_data_7), .QB (nx17244), .D (nx14861), .CLK (
         clk), .R (reset)) ;
    xor2 ix3641 (.Y (nx3640), .A0 (nx17247), .A1 (nx17250)) ;
    or02 ix3895 (.Y (mem_addr_out[8]), .A0 (nx3892), .A1 (nx3816)) ;
    oai222 ix3893 (.Y (nx3892), .A0 (nx17255), .A1 (nx18135), .B0 (nx17277), .B1 (
           nx18089), .C0 (nx3884), .C1 (nx18075)) ;
    xnor2 ix17256 (.Y (nx17255), .A0 (nx17257), .A1 (nx17260)) ;
    dffr reg_bias_offset_reg_q_8 (.Q (bias_offset_data_out_8), .QB (nx17265), .D (
         nx14961), .CLK (clk), .R (reset)) ;
    aoi21 ix955 (.Y (nx954), .A0 (nx15692), .A1 (nx15686), .B0 (nx948)) ;
    dffs_ni reg_write_base_reg_q_8 (.Q (write_base_data_out_8), .QB (nx17268), .D (
            nx14911), .CLK (nx17841), .S (reset)) ;
    xnor2 ix17271 (.Y (nx17270), .A0 (nx17272), .A1 (nx17275)) ;
    xnor2 ix17278 (.Y (nx17277), .A0 (nx17279), .A1 (nx17282)) ;
    dffr img_base_addr_inst_reg_q_8 (.Q (img_base_addr_8), .QB (nx17294), .D (
         nx14941), .CLK (clk), .R (reset)) ;
    oai21 ix3839 (.Y (nx3838), .A0 (nx17287), .A1 (nx17291), .B0 (nx3832)) ;
    dffr reg_write_base_prev_reg_q_8 (.Q (\$dummy [135]), .QB (nx17287), .D (
         nx14931), .CLK (clk), .R (reset)) ;
    nor02_2x ix17292 (.Y (nx17291), .A0 (nx3548), .A1 (
             write_base_prev_data_out_7)) ;
    nand02 ix3833 (.Y (nx3832), .A0 (nx17291), .A1 (nx17287)) ;
    aoi21 ix3853 (.Y (nx3852), .A0 (nx17231), .A1 (nx17298), .B0 (nx3846)) ;
    dffr reg_img_addr_offset_8 (.Q (img_addr_offset_8), .QB (nx17298), .D (
         nx14951), .CLK (clk), .R (nx18033)) ;
    oai222 ix3817 (.Y (nx3816), .A0 (nx17307), .A1 (nx18143), .B0 (nx17302), .B1 (
           nx17312), .C0 (nx17315), .C1 (nx18139)) ;
    xor2 ix17308 (.Y (nx17307), .A0 (nx3760), .A1 (nx17310)) ;
    aoi21 ix17313 (.Y (nx17312), .A0 (nx3742), .A1 (nx17857), .B0 (nx17975)) ;
    dffr reg_addr1_data_8 (.Q (addr1_data_8), .QB (nx17315), .D (nx14921), .CLK (
         clk), .R (reset)) ;
    nand02 ix4037 (.Y (mem_addr_out[9]), .A0 (nx17321), .A1 (nx17362)) ;
    aoi222 ix17322 (.Y (nx17321), .A0 (nx17323), .A1 (nx17857), .B0 (nx4022), .B1 (
           nx18021), .C0 (nx4002), .C1 (nx18003)) ;
    xnor2 ix3915 (.Y (nx3914), .A0 (nx18694), .A1 (nx17331)) ;
    dffs_ni reg_write_base_reg_q_9 (.Q (write_base_data_out_9), .QB (nx17326), .D (
            nx14971), .CLK (nx17841), .S (reset)) ;
    xnor2 ix4023 (.Y (nx4022), .A0 (nx4012), .A1 (nx17337)) ;
    dffr reg_bias_offset_reg_q_9 (.Q (bias_offset_data_out_9), .QB (nx17341), .D (
         nx15021), .CLK (clk), .R (reset)) ;
    xnor2 ix4003 (.Y (nx4002), .A0 (nx3966), .A1 (nx17345)) ;
    dffr img_base_addr_inst_reg_q_9 (.Q (img_base_addr_9), .QB (\$dummy [136]), 
         .D (nx15001), .CLK (clk), .R (reset)) ;
    xnor2 ix3981 (.Y (nx3980), .A0 (write_base_prev_data_out_9), .A1 (nx3832)) ;
    dffr reg_write_base_prev_reg_q_9 (.Q (write_base_prev_data_out_9), .QB (
         \$dummy [137]), .D (nx14991), .CLK (clk), .R (reset)) ;
    oai21 ix17357 (.Y (nx17356), .A0 (nx3846), .A1 (img_addr_offset_9), .B0 (
          nx17358)) ;
    nand02 ix17359 (.Y (nx17358), .A0 (img_addr_offset_9), .A1 (nx3846)) ;
    dffr reg_img_addr_offset_9 (.Q (img_addr_offset_9), .QB (nx17360), .D (
         nx15011), .CLK (clk), .R (nx18033)) ;
    aoi222 ix17363 (.Y (nx17362), .A0 (addr1_data_9), .A1 (nx18037), .B0 (nx3924
           ), .B1 (nx18017), .C0 (nx3934), .C1 (nx3938)) ;
    oai21 ix17367 (.Y (nx17366), .A0 (nx3800), .A1 (addr1_data_9), .B0 (nx17369)
          ) ;
    nand02 ix17370 (.Y (nx17369), .A0 (addr1_data_9), .A1 (nx3800)) ;
    dffr reg_addr1_data_9 (.Q (addr1_data_9), .QB (nx17371), .D (nx14981), .CLK (
         clk), .R (reset)) ;
    xor2 ix3925 (.Y (nx3924), .A0 (nx17374), .A1 (nx17377)) ;
    aoi22 ix17375 (.Y (nx17374), .A0 (write_offset_data_out_8), .A1 (nx18897), .B0 (
          nx3760), .B1 (nx3780)) ;
    or02 ix4179 (.Y (mem_addr_out[10]), .A0 (nx4176), .A1 (nx4100)) ;
    oai222 ix4177 (.Y (nx4176), .A0 (nx17382), .A1 (nx18135), .B0 (nx17404), .B1 (
           nx18089), .C0 (nx4168), .C1 (nx18075)) ;
    xnor2 ix17383 (.Y (nx17382), .A0 (nx17384), .A1 (nx17387)) ;
    dffr reg_bias_offset_reg_q_10 (.Q (bias_offset_data_out_10), .QB (nx17392), 
         .D (nx15081), .CLK (clk), .R (reset)) ;
    aoi21 ix1001 (.Y (nx1000), .A0 (nx15679), .A1 (nx15673), .B0 (nx994)) ;
    dffr reg_write_base_reg_q_10 (.Q (write_base_data_out_10), .QB (nx17395), .D (
         nx15031), .CLK (nx17841), .R (reset)) ;
    xnor2 ix17398 (.Y (nx17397), .A0 (nx17399), .A1 (nx17402)) ;
    xnor2 ix17405 (.Y (nx17404), .A0 (nx17406), .A1 (nx17409)) ;
    dffr img_base_addr_inst_reg_q_10 (.Q (img_base_addr_10), .QB (nx17421), .D (
         nx15061), .CLK (clk), .R (reset)) ;
    oai21 ix4123 (.Y (nx4122), .A0 (nx17414), .A1 (nx17418), .B0 (nx4116)) ;
    dffr reg_write_base_prev_reg_q_10 (.Q (\$dummy [138]), .QB (nx17414), .D (
         nx15051), .CLK (clk), .R (reset)) ;
    nor02_2x ix17419 (.Y (nx17418), .A0 (nx3832), .A1 (
             write_base_prev_data_out_9)) ;
    nand02 ix4117 (.Y (nx4116), .A0 (nx17418), .A1 (nx17414)) ;
    aoi21 ix4137 (.Y (nx4136), .A0 (nx17358), .A1 (nx17425), .B0 (nx4130)) ;
    dffr reg_img_addr_offset_10 (.Q (img_addr_offset_10), .QB (nx17425), .D (
         nx15071), .CLK (clk), .R (nx18033)) ;
    oai222 ix4101 (.Y (nx4100), .A0 (nx17434), .A1 (nx18143), .B0 (nx17429), .B1 (
           nx17439), .C0 (nx17442), .C1 (nx18139)) ;
    xor2 ix17435 (.Y (nx17434), .A0 (nx4044), .A1 (nx17437)) ;
    oai22 ix4045 (.Y (nx4044), .A0 (nx17374), .A1 (nx17377), .B0 (nx15770), .B1 (
          nx17326)) ;
    aoi21 ix17440 (.Y (nx17439), .A0 (nx4026), .A1 (nx17859), .B0 (nx17977)) ;
    dffr reg_addr1_data_10 (.Q (addr1_data_10), .QB (nx17442), .D (nx15041), .CLK (
         clk), .R (reset)) ;
    nand02 ix4321 (.Y (mem_addr_out[11]), .A0 (nx17448), .A1 (nx17489)) ;
    aoi222 ix17449 (.Y (nx17448), .A0 (nx17450), .A1 (nx17859), .B0 (nx4306), .B1 (
           nx18023), .C0 (nx4286), .C1 (nx18005)) ;
    xnor2 ix4199 (.Y (nx4198), .A0 (nx4194), .A1 (nx17458)) ;
    dffs_ni reg_write_base_reg_q_11 (.Q (write_base_data_out_11), .QB (nx17453)
            , .D (nx15091), .CLK (nx17841), .S (reset)) ;
    xnor2 ix4307 (.Y (nx4306), .A0 (nx4296), .A1 (nx17464)) ;
    dffr reg_bias_offset_reg_q_11 (.Q (bias_offset_data_out_11), .QB (nx17468), 
         .D (nx15141), .CLK (clk), .R (reset)) ;
    xnor2 ix4287 (.Y (nx4286), .A0 (nx4250), .A1 (nx17472)) ;
    dffs_ni img_base_addr_inst_reg_q_11 (.Q (img_base_addr_11), .QB (
            \$dummy [139]), .D (nx15121), .CLK (clk), .S (reset)) ;
    xnor2 ix4265 (.Y (nx4264), .A0 (write_base_prev_data_out_11), .A1 (nx4116)
          ) ;
    dffr reg_write_base_prev_reg_q_11 (.Q (write_base_prev_data_out_11), .QB (
         \$dummy [140]), .D (nx15111), .CLK (clk), .R (reset)) ;
    oai21 ix17484 (.Y (nx17483), .A0 (nx4130), .A1 (img_addr_offset_11), .B0 (
          nx17485)) ;
    nand02 ix17486 (.Y (nx17485), .A0 (img_addr_offset_11), .A1 (nx4130)) ;
    dffr reg_img_addr_offset_11 (.Q (img_addr_offset_11), .QB (nx17487), .D (
         nx15131), .CLK (clk), .R (nx18033)) ;
    aoi222 ix17490 (.Y (nx17489), .A0 (addr1_data_11), .A1 (nx18037), .B0 (
           nx4218), .B1 (nx4222), .C0 (nx4208), .C1 (nx18017)) ;
    oai21 ix17494 (.Y (nx17493), .A0 (nx4084), .A1 (addr1_data_11), .B0 (nx17496
          )) ;
    nand02 ix17497 (.Y (nx17496), .A0 (addr1_data_11), .A1 (nx4084)) ;
    dffr reg_addr1_data_11 (.Q (addr1_data_11), .QB (nx17498), .D (nx15101), .CLK (
         clk), .R (reset)) ;
    xor2 ix4209 (.Y (nx4208), .A0 (nx17502), .A1 (nx17505)) ;
    xnor2 ix17510 (.Y (nx17509), .A0 (nx17511), .A1 (nx17514)) ;
    dffr reg_bias_offset_reg_q_12 (.Q (bias_offset_data_out_12), .QB (nx17519), 
         .D (nx15201), .CLK (clk), .R (reset)) ;
    aoi21 ix1049 (.Y (nx1048), .A0 (nx15666), .A1 (nx15660), .B0 (nx1042)) ;
    dffs_ni reg_write_base_reg_q_12 (.Q (write_base_data_out_12), .QB (nx17522)
            , .D (nx15151), .CLK (nx17843), .S (reset)) ;
    dffs_ni img_base_addr_inst_reg_q_12 (.Q (img_base_addr_12), .QB (nx17548), .D (
            nx15181), .CLK (clk), .S (reset)) ;
    oai21 ix4407 (.Y (nx4406), .A0 (nx17541), .A1 (nx17545), .B0 (nx4400)) ;
    dffr reg_write_base_prev_reg_q_12 (.Q (\$dummy [141]), .QB (nx17541), .D (
         nx15171), .CLK (clk), .R (reset)) ;
    nor02_2x ix17546 (.Y (nx17545), .A0 (nx4116), .A1 (
             write_base_prev_data_out_11)) ;
    nand02 ix4401 (.Y (nx4400), .A0 (nx17545), .A1 (nx17541)) ;
    aoi21 ix4421 (.Y (nx4420), .A0 (nx17485), .A1 (nx17552), .B0 (nx4414)) ;
    dffr reg_img_addr_offset_12 (.Q (img_addr_offset_12), .QB (nx17552), .D (
         nx15191), .CLK (clk), .R (nx18033)) ;
    xor2 ix17562 (.Y (nx17561), .A0 (nx4328), .A1 (nx17564)) ;
    dffr reg_addr1_data_12 (.Q (addr1_data_12), .QB (nx17566), .D (nx15161), .CLK (
         clk), .R (reset)) ;
    nand02 ix4605 (.Y (mem_addr_out[13]), .A0 (nx17575), .A1 (nx17616)) ;
    aoi222 ix17576 (.Y (nx17575), .A0 (nx17577), .A1 (nx17859), .B0 (nx4590), .B1 (
           nx18023), .C0 (nx4570), .C1 (nx18005)) ;
    dffr reg_write_base_reg_q_13 (.Q (write_base_data_out_13), .QB (nx17580), .D (
         nx15211), .CLK (nx17843), .R (reset)) ;
    xnor2 ix4591 (.Y (nx4590), .A0 (nx18726), .A1 (nx17591)) ;
    dffr reg_bias_offset_reg_q_13 (.Q (bias_offset_data_out_13), .QB (nx17595), 
         .D (nx15261), .CLK (clk), .R (reset)) ;
    xnor2 ix4571 (.Y (nx4570), .A0 (nx4534), .A1 (nx17599)) ;
    oai22 ix4535 (.Y (nx4534), .A0 (nx18838), .A1 (nx17536), .B0 (nx17552), .B1 (
          nx17548)) ;
    dffr img_base_addr_inst_reg_q_13 (.Q (img_base_addr_13), .QB (\$dummy [142])
         , .D (nx15241), .CLK (clk), .R (reset)) ;
    xnor2 ix4549 (.Y (nx4548), .A0 (write_base_prev_data_out_13), .A1 (nx4400)
          ) ;
    dffr reg_write_base_prev_reg_q_13 (.Q (write_base_prev_data_out_13), .QB (
         \$dummy [143]), .D (nx15231), .CLK (clk), .R (reset)) ;
    oai21 ix17611 (.Y (nx17610), .A0 (nx4414), .A1 (img_addr_offset_13), .B0 (
          nx17612)) ;
    nand02 ix17613 (.Y (nx17612), .A0 (img_addr_offset_13), .A1 (nx4414)) ;
    dffr reg_img_addr_offset_13 (.Q (img_addr_offset_13), .QB (nx17614), .D (
         nx15251), .CLK (clk), .R (nx18033)) ;
    aoi222 ix17617 (.Y (nx17616), .A0 (addr1_data_13), .A1 (nx18039), .B0 (
           nx4502), .B1 (nx4506), .C0 (nx4492), .C1 (nx2642)) ;
    oai21 ix17621 (.Y (nx17620), .A0 (nx4368), .A1 (addr1_data_13), .B0 (nx17623
          )) ;
    nand02 ix17624 (.Y (nx17623), .A0 (addr1_data_13), .A1 (nx4368)) ;
    dffr reg_addr1_data_13 (.Q (addr1_data_13), .QB (nx17625), .D (nx15221), .CLK (
         clk), .R (reset)) ;
    xor2 ix4493 (.Y (nx4492), .A0 (nx17629), .A1 (nx17632)) ;
    or02 ix4747 (.Y (mem_addr_out[14]), .A0 (nx4744), .A1 (nx4668)) ;
    oai222 ix4745 (.Y (nx4744), .A0 (nx17636), .A1 (nx18135), .B0 (nx17658), .B1 (
           nx18091), .C0 (nx4736), .C1 (nx18339)) ;
    xnor2 ix17637 (.Y (nx17636), .A0 (nx17638), .A1 (nx17641)) ;
    dffr reg_bias_offset_reg_q_14 (.Q (bias_offset_data_out_14), .QB (nx17646), 
         .D (nx15321), .CLK (clk), .R (reset)) ;
    dffr reg_write_base_reg_q_14 (.Q (write_base_data_out_14), .QB (nx17649), .D (
         nx15271), .CLK (nx17843), .R (reset)) ;
    xnor2 ix17659 (.Y (nx17658), .A0 (nx17660), .A1 (nx17663)) ;
    aoi22 ix17661 (.Y (nx17660), .A0 (img_addr_offset_13), .A1 (img_base_addr_13
          ), .B0 (nx4534), .B1 (nx4568)) ;
    dffr img_base_addr_inst_reg_q_14 (.Q (img_base_addr_14), .QB (nx17673), .D (
         nx15301), .CLK (clk), .R (reset)) ;
    dffr reg_write_base_prev_reg_q_14 (.Q (\$dummy [144]), .QB (nx17670), .D (
         nx15291), .CLK (clk), .R (reset)) ;
    nor02_2x ix17672 (.Y (nx17671), .A0 (nx4400), .A1 (
             write_base_prev_data_out_13)) ;
    dffr reg_img_addr_offset_14 (.Q (img_addr_offset_14), .QB (nx17677), .D (
         nx15311), .CLK (clk), .R (nx18035)) ;
    oai222 ix4669 (.Y (nx4668), .A0 (nx17682), .A1 (nx18143), .B0 (nx17687), .B1 (
           nx18139), .C0 (nx17679), .C1 (nx17692)) ;
    xor2 ix17683 (.Y (nx17682), .A0 (nx18627), .A1 (nx17685)) ;
    dffr reg_addr1_data_14 (.Q (addr1_data_14), .QB (nx17687), .D (nx15281), .CLK (
         clk), .R (reset)) ;
    aoi21 ix17693 (.Y (nx17692), .A0 (nx4594), .A1 (nx17859), .B0 (nx17977)) ;
    nand02 ix4859 (.Y (mem_addr_out[15]), .A0 (nx17696), .A1 (nx17728)) ;
    aoi222 ix17697 (.Y (nx17696), .A0 (nx4816), .A1 (nx18381), .B0 (nx17977), .B1 (
           nx4812), .C0 (nx4850), .C1 (nx18005)) ;
    xnor2 ix4817 (.Y (nx4816), .A0 (nx4736), .A1 (nx4812)) ;
    xnor2 ix4813 (.Y (nx4812), .A0 (nx17700), .A1 (write_base_data_out_15)) ;
    nand02 ix17701 (.Y (nx17700), .A0 (write_base_data_out_14), .A1 (nx4496)) ;
    dffs_ni reg_write_base_reg_q_15 (.Q (write_base_data_out_15), .QB (
            \$dummy [145]), .D (nx15341), .CLK (nx17843), .S (reset)) ;
    xnor2 ix4851 (.Y (nx4850), .A0 (nx4826), .A1 (nx17711)) ;
    oai22 ix4827 (.Y (nx4826), .A0 (nx17660), .A1 (nx17663), .B0 (nx17677), .B1 (
          nx17673)) ;
    dffs_ni img_base_addr_inst_reg_q_15 (.Q (img_base_addr_15), .QB (
            \$dummy [146]), .D (nx15371), .CLK (clk), .S (reset)) ;
    xnor2 ix4835 (.Y (nx4834), .A0 (write_base_prev_data_out_15), .A1 (nx4684)
          ) ;
    dffr reg_write_base_prev_reg_q_15 (.Q (write_base_prev_data_out_15), .QB (
         \$dummy [147]), .D (nx15361), .CLK (clk), .R (reset)) ;
    nand02 ix4685 (.Y (nx4684), .A0 (nx17671), .A1 (nx17670)) ;
    dffr img_addr_offset_15 (.Q (\$dummy [148]), .QB (nx17726), .D (nx15381), .CLK (
         clk), .R (nx18035)) ;
    aoi222 ix17729 (.Y (nx17728), .A0 (nx4804), .A1 (nx2642), .B0 (addr1_data_15
           ), .B1 (nx18039), .C0 (nx4782), .C1 (nx18023)) ;
    xnor2 ix4805 (.Y (nx4804), .A0 (nx17731), .A1 (nx4802)) ;
    dffr reg_addr1_data_15 (.Q (addr1_data_15), .QB (nx17740), .D (nx15351), .CLK (
         clk), .R (reset)) ;
    xnor2 ix4783 (.Y (nx4782), .A0 (nx4754), .A1 (nx17744)) ;
    oai22 ix4755 (.Y (nx4754), .A0 (nx18725), .A1 (nx17641), .B0 (nx18915), .B1 (
          nx17646)) ;
    dffr reg_bias_offset_reg_q_15 (.Q (bias_offset_data_out_15), .QB (nx17748), 
         .D (nx15331), .CLK (clk), .R (reset)) ;
    inv01 ix1961 (.Y (mem_data_out[0]), .A (nx17751)) ;
    aoi222 ix17752 (.Y (nx17751), .A0 (comp_unit_data2_in[0]), .A1 (nx17909), .B0 (
           comp_unit_data1_in[0]), .B1 (nx17915), .C0 (argmax_data_in[0]), .C1 (
           nx17979)) ;
    inv01 ix1971 (.Y (mem_data_out[1]), .A (nx17754)) ;
    aoi222 ix17755 (.Y (nx17754), .A0 (comp_unit_data2_in[1]), .A1 (nx17909), .B0 (
           comp_unit_data1_in[1]), .B1 (nx17915), .C0 (argmax_data_in[1]), .C1 (
           nx17979)) ;
    inv01 ix1981 (.Y (mem_data_out[2]), .A (nx17757)) ;
    aoi222 ix17758 (.Y (nx17757), .A0 (comp_unit_data2_in[2]), .A1 (nx17909), .B0 (
           comp_unit_data1_in[2]), .B1 (nx17915), .C0 (argmax_data_in[2]), .C1 (
           nx17979)) ;
    inv01 ix1991 (.Y (mem_data_out[3]), .A (nx17760)) ;
    aoi222 ix17761 (.Y (nx17760), .A0 (comp_unit_data2_in[3]), .A1 (nx17909), .B0 (
           comp_unit_data1_in[3]), .B1 (nx17915), .C0 (argmax_data_in[3]), .C1 (
           nx17979)) ;
    inv01 ix2001 (.Y (mem_data_out[4]), .A (nx17763)) ;
    aoi222 ix17764 (.Y (nx17763), .A0 (comp_unit_data2_in[4]), .A1 (nx17909), .B0 (
           comp_unit_data1_in[4]), .B1 (nx17915), .C0 (argmax_data_in[4]), .C1 (
           nx17979)) ;
    inv01 ix2011 (.Y (mem_data_out[5]), .A (nx17766)) ;
    aoi222 ix17767 (.Y (nx17766), .A0 (comp_unit_data2_in[5]), .A1 (nx17909), .B0 (
           comp_unit_data1_in[5]), .B1 (nx17917), .C0 (argmax_data_in[5]), .C1 (
           nx17979)) ;
    inv01 ix2021 (.Y (mem_data_out[6]), .A (nx17769)) ;
    aoi222 ix17770 (.Y (nx17769), .A0 (comp_unit_data2_in[6]), .A1 (nx17911), .B0 (
           comp_unit_data1_in[6]), .B1 (nx17917), .C0 (argmax_data_in[6]), .C1 (
           nx17979)) ;
    inv01 ix2031 (.Y (mem_data_out[7]), .A (nx17772)) ;
    aoi222 ix17773 (.Y (nx17772), .A0 (comp_unit_data2_in[7]), .A1 (nx17911), .B0 (
           comp_unit_data1_in[7]), .B1 (nx17917), .C0 (argmax_data_in[7]), .C1 (
           nx17981)) ;
    inv01 ix2041 (.Y (mem_data_out[8]), .A (nx17775)) ;
    aoi222 ix17776 (.Y (nx17775), .A0 (comp_unit_data2_in[8]), .A1 (nx17911), .B0 (
           comp_unit_data1_in[8]), .B1 (nx17917), .C0 (argmax_data_in[8]), .C1 (
           nx17981)) ;
    inv01 ix2051 (.Y (mem_data_out[9]), .A (nx17778)) ;
    aoi222 ix17779 (.Y (nx17778), .A0 (comp_unit_data2_in[9]), .A1 (nx17911), .B0 (
           comp_unit_data1_in[9]), .B1 (nx17917), .C0 (argmax_data_in[9]), .C1 (
           nx17981)) ;
    inv01 ix2061 (.Y (mem_data_out[10]), .A (nx17781)) ;
    aoi222 ix17782 (.Y (nx17781), .A0 (comp_unit_data2_in[10]), .A1 (nx17911), .B0 (
           comp_unit_data1_in[10]), .B1 (nx17917), .C0 (argmax_data_in[10]), .C1 (
           nx17981)) ;
    inv01 ix2071 (.Y (mem_data_out[11]), .A (nx17784)) ;
    aoi222 ix17785 (.Y (nx17784), .A0 (comp_unit_data2_in[11]), .A1 (nx17911), .B0 (
           comp_unit_data1_in[11]), .B1 (nx17917), .C0 (argmax_data_in[11]), .C1 (
           nx17981)) ;
    inv01 ix2081 (.Y (mem_data_out[12]), .A (nx17787)) ;
    aoi222 ix17788 (.Y (nx17787), .A0 (comp_unit_data2_in[12]), .A1 (nx17911), .B0 (
           comp_unit_data1_in[12]), .B1 (nx17919), .C0 (argmax_data_in[12]), .C1 (
           nx17981)) ;
    inv01 ix2091 (.Y (mem_data_out[13]), .A (nx17790)) ;
    aoi222 ix17791 (.Y (nx17790), .A0 (comp_unit_data2_in[13]), .A1 (nx17913), .B0 (
           comp_unit_data1_in[13]), .B1 (nx17919), .C0 (argmax_data_in[13]), .C1 (
           nx17981)) ;
    inv01 ix2101 (.Y (mem_data_out[14]), .A (nx17793)) ;
    aoi222 ix17794 (.Y (nx17793), .A0 (comp_unit_data2_in[14]), .A1 (nx17913), .B0 (
           comp_unit_data1_in[14]), .B1 (nx17919), .C0 (argmax_data_in[14]), .C1 (
           nx17983)) ;
    inv01 ix2111 (.Y (mem_data_out[15]), .A (nx17796)) ;
    aoi222 ix17797 (.Y (nx17796), .A0 (comp_unit_data2_in[15]), .A1 (nx17913), .B0 (
           comp_unit_data1_in[15]), .B1 (nx17919), .C0 (argmax_data_in[15]), .C1 (
           nx17983)) ;
    inv01 ix4595 (.Y (nx4594), .A (nx17577)) ;
    inv01 ix4569 (.Y (nx4568), .A (nx17599)) ;
    inv01 ix4027 (.Y (nx4026), .A (nx17323)) ;
    inv01 ix3781 (.Y (nx3780), .A (nx17310)) ;
    inv01 ix3743 (.Y (nx3742), .A (nx17196)) ;
    inv01 ix3459 (.Y (nx3458), .A (nx18543)) ;
    inv01 ix16979 (.Y (nx16978), .A (nx3078)) ;
    inv01 ix3075 (.Y (nx3074), .A (nx16976)) ;
    inv01 ix3049 (.Y (nx3048), .A (nx16943)) ;
    inv01 ix2969 (.Y (nx2968), .A (nx16956)) ;
    inv01 ix2927 (.Y (nx2926), .A (nx16874)) ;
    inv01 ix2739 (.Y (nx2738), .A (nx16738)) ;
    inv01 ix2665 (.Y (nx2664), .A (nx16786)) ;
    inv01 ix2623 (.Y (nx2622), .A (nx16806)) ;
    inv01 ix16630 (.Y (nx16629), .A (nx2546)) ;
    inv01 ix1803 (.Y (nx12910), .A (nx16282)) ;
    inv01 ix1681 (.Y (nx12908), .A (nx16265)) ;
    inv01 ix1461 (.Y (nx1460), .A (nx15609)) ;
    inv01 ix15620 (.Y (nx15619), .A (nx1182)) ;
    inv01 ix781 (.Y (nx780), .A (nx15765)) ;
    inv01 ix637 (.Y (nx636), .A (nx16189)) ;
    inv01 ix631 (.Y (nx630), .A (nx16191)) ;
    inv01 ix583 (.Y (nx582), .A (nx15479)) ;
    inv01 ix15975 (.Y (nx15974), .A (nx576)) ;
    inv01 ix15397 (.Y (nx15396), .A (nx316)) ;
    inv01 ix1859 (.Y (nx12877), .A (nx16204)) ;
    inv01 ix15423 (.Y (nx15422), .A (nx12875)) ;
    inv01 ix149 (.Y (nx148), .A (nx15533)) ;
    inv01 ix303 (.Y (comp_unit_flt_size), .A (nx16610)) ;
    inv01 ix17802 (.Y (nx17803), .A (current_state_13)) ;
    inv02 ix17804 (.Y (nx17805), .A (nx17803)) ;
    inv02 ix17806 (.Y (nx17807), .A (nx17803)) ;
    inv02 ix17808 (.Y (nx17809), .A (nx17803)) ;
    buf02 ix17810 (.Y (nx17811), .A (wind_width_count_0)) ;
    buf02 ix17812 (.Y (nx17813), .A (wind_width_count_0)) ;
    buf02 ix17814 (.Y (nx17815), .A (cache_width_count_4)) ;
    buf02 ix17816 (.Y (nx17817), .A (cache_width_count_4)) ;
    buf02 ix17818 (.Y (nx17819), .A (cache_width_count_2)) ;
    buf02 ix17820 (.Y (nx17821), .A (cache_width_count_2)) ;
    inv02 ix17822 (.Y (nx17823), .A (clk)) ;
    inv02 ix17824 (.Y (nx17825), .A (clk)) ;
    inv02 ix17826 (.Y (nx17827), .A (clk)) ;
    inv02 ix17828 (.Y (nx17829), .A (clk)) ;
    inv02 ix17830 (.Y (nx17831), .A (clk)) ;
    inv02 ix17832 (.Y (nx17833), .A (clk)) ;
    inv02 ix17834 (.Y (nx17835), .A (clk)) ;
    inv02 ix17836 (.Y (nx17837), .A (clk)) ;
    inv02 ix17838 (.Y (nx17839), .A (clk)) ;
    inv02 ix17840 (.Y (nx17841), .A (clk)) ;
    inv02 ix17842 (.Y (nx17843), .A (clk)) ;
    inv02 ix17844 (.Y (nx17845), .A (nx18305)) ;
    inv02 ix17846 (.Y (nx17847), .A (nx18305)) ;
    inv02 ix17854 (.Y (nx17855), .A (nx18339)) ;
    inv02 ix17856 (.Y (nx17857), .A (nx18339)) ;
    inv02 ix17858 (.Y (nx17859), .A (nx18339)) ;
    inv01 ix17862 (.Y (nx17863), .A (filter_ready_out)) ;
    inv02 ix17864 (.Y (nx17865), .A (nx18319)) ;
    inv02 ix17868 (.Y (nx17869), .A (nx18319)) ;
    inv02 ix17870 (.Y (nx17871), .A (nx15605)) ;
    inv02 ix17872 (.Y (nx17873), .A (nx15605)) ;
    inv02 ix17874 (.Y (nx17875), .A (nx18333)) ;
    inv02 ix17876 (.Y (nx17877), .A (nx18333)) ;
    inv02 ix17878 (.Y (nx17879), .A (nx18333)) ;
    inv02 ix17886 (.Y (nx17887), .A (nx15530)) ;
    buf02 ix17892 (.Y (nx17893), .A (current_state_4)) ;
    buf02 ix17894 (.Y (nx17895), .A (current_state_4)) ;
    inv02 ix17896 (.Y (nx17897), .A (nx15435)) ;
    inv02 ix17898 (.Y (nx17899), .A (nx15435)) ;
    inv02 ix17906 (.Y (nx17907), .A (nx18323)) ;
    inv02 ix17908 (.Y (nx17909), .A (nx15716)) ;
    inv02 ix17910 (.Y (nx17911), .A (nx15716)) ;
    inv02 ix17912 (.Y (nx17913), .A (nx15716)) ;
    inv02 ix17914 (.Y (nx17915), .A (nx15541)) ;
    inv02 ix17916 (.Y (nx17917), .A (nx15541)) ;
    inv02 ix17918 (.Y (nx17919), .A (nx15541)) ;
    inv02 ix17920 (.Y (nx17921), .A (nx15626)) ;
    inv02 ix17922 (.Y (nx17923), .A (nx18279)) ;
    inv02 ix17926 (.Y (nx17927), .A (nx15392)) ;
    buf02 ix17928 (.Y (nx17929), .A (nx206)) ;
    inv01 ix17936 (.Y (nx17937), .A (nx378)) ;
    inv02 ix17938 (.Y (nx17939), .A (nx17937)) ;
    inv02 ix17940 (.Y (nx17941), .A (nx17937)) ;
    inv02 ix17942 (.Y (nx17943), .A (nx17937)) ;
    inv02 ix17946 (.Y (nx17947), .A (nx17945)) ;
    inv02 ix17948 (.Y (nx17949), .A (nx18329)) ;
    inv02 ix17950 (.Y (nx17951), .A (nx18329)) ;
    inv01 ix17958 (.Y (nx17959), .A (nx1224)) ;
    inv02 ix17960 (.Y (nx17961), .A (nx17959)) ;
    inv02 ix17962 (.Y (nx17963), .A (nx17959)) ;
    inv02 ix17964 (.Y (nx17965), .A (nx17959)) ;
    inv02 ix17970 (.Y (nx17971), .A (nx15554)) ;
    buf02 ix17972 (.Y (nx17973), .A (nx1546)) ;
    inv02 ix17974 (.Y (nx17975), .A (nx16732)) ;
    inv02 ix17978 (.Y (nx17979), .A (nx18883)) ;
    inv02 ix17980 (.Y (nx17981), .A (nx18884)) ;
    inv02 ix17982 (.Y (nx17983), .A (nx18884)) ;
    nor02_2x ix17992 (.Y (nx17993), .A0 (nx16302), .A1 (nx18153)) ;
    nor02_2x ix17994 (.Y (nx17995), .A0 (nx16302), .A1 (nx18153)) ;
    inv02 ix17996 (.Y (nx17997), .A (nx18117)) ;
    inv02 ix17998 (.Y (nx17999), .A (nx18117)) ;
    inv02 ix18000 (.Y (nx18001), .A (nx18117)) ;
    inv02 ix18002 (.Y (nx18003), .A (nx18091)) ;
    inv02 ix18004 (.Y (nx18005), .A (nx18091)) ;
    inv02 ix18006 (.Y (nx18007), .A (nx16745)) ;
    inv02 ix18010 (.Y (nx18011), .A (nx16927)) ;
    inv02 ix18016 (.Y (nx18017), .A (nx18143)) ;
    inv02 ix18020 (.Y (nx18021), .A (nx18137)) ;
    inv02 ix18022 (.Y (nx18023), .A (nx18137)) ;
    buf02 ix18026 (.Y (nx18027), .A (img_addr_offset_0)) ;
    inv01 ix18028 (.Y (nx18029), .A (nx2712)) ;
    inv02 ix18030 (.Y (nx18031), .A (nx18029)) ;
    inv02 ix18032 (.Y (nx18033), .A (nx18029)) ;
    inv02 ix18034 (.Y (nx18035), .A (nx18029)) ;
    inv02 ix18036 (.Y (nx18037), .A (nx18141)) ;
    inv02 ix18038 (.Y (nx18039), .A (nx18141)) ;
    inv02 ix18040 (.Y (nx18041), .A (nx18911)) ;
    buf02 ix18044 (.Y (nx18045), .A (nx15630)) ;
    buf02 ix18046 (.Y (nx18047), .A (nx15630)) ;
    inv02 ix18048 (.Y (nx18049), .A (nx760)) ;
    inv02 ix18050 (.Y (nx18051), .A (nx18229)) ;
    inv02 ix18052 (.Y (nx18053), .A (nx18229)) ;
    buf02 ix18054 (.Y (nx18055), .A (nx16028)) ;
    inv01 ix18058 (.Y (nx18059), .A (current_state_18)) ;
    inv01 ix18062 (.Y (nx18063), .A (nx18233)) ;
    inv01 ix18064 (.Y (nx18065), .A (nx18233)) ;
    inv01 ix18066 (.Y (nx18067), .A (nx18233)) ;
    inv02 ix18068 (.Y (nx18069), .A (nx19308)) ;
    inv02 ix18076 (.Y (nx18077), .A (nx18381)) ;
    inv02 ix18080 (.Y (nx18081), .A (nx2580)) ;
    inv02 ix18084 (.Y (nx18085), .A (nx18243)) ;
    inv02 ix18086 (.Y (nx18087), .A (nx18243)) ;
    inv02 ix18088 (.Y (nx18089), .A (nx18243)) ;
    inv02 ix18090 (.Y (nx18091), .A (nx18243)) ;
    inv02 ix18116 (.Y (nx18117), .A (nx2142)) ;
    inv02 ix18120 (.Y (nx18121), .A (nx18119)) ;
    inv02 ix18136 (.Y (nx18137), .A (nx2664)) ;
    inv02 ix18138 (.Y (nx18139), .A (nx2766)) ;
    inv02 ix18140 (.Y (nx18141), .A (nx2766)) ;
    inv02 ix18142 (.Y (nx18143), .A (nx2642)) ;
    buf02 ix18150 (.Y (nx18151), .A (comp_unit_operation)) ;
    buf02 ix18152 (.Y (nx18153), .A (comp_unit_operation)) ;
    inv01 ix18154 (.Y (nx18155), .A (nx18385)) ;
    inv01 ix18156 (.Y (nx18157), .A (nx18385)) ;
    xnor2 ix311 (.Y (nx310), .A0 (nx15591), .A1 (nx308)) ;
    mux21_ni ix13012 (.Y (nx13011), .A0 (nx262), .A1 (cntr1_inst_counter_out_4)
             , .S0 (nx18255)) ;
    xor2 ix263 (.Y (nx262), .A0 (nx15591), .A1 (nx15402)) ;
    mux21_ni ix13002 (.Y (nx13001), .A0 (nx244), .A1 (cntr1_inst_counter_out_3)
             , .S0 (nx18255)) ;
    mux21_ni ix12992 (.Y (nx12991), .A0 (nx230), .A1 (cntr1_inst_counter_out_2)
             , .S0 (nx18255)) ;
    mux21 ix12982 (.Y (nx12981), .A0 (nx16307), .A1 (nx15416), .S0 (nx18255)) ;
    nand02 ix207 (.Y (nx206), .A0 (nx16313), .A1 (nx17803)) ;
    nor02ii ix141 (.Y (nx140), .A0 (nx15450), .A1 (io_ready_in)) ;
    and03 ix1797 (.Y (nx1796), .A0 (nx12873), .A1 (nx15486), .A2 (nx18163)) ;
    inv01 ix18162 (.Y (nx18163), .A (nx16269)) ;
    and02 ix15480 (.Y (nx15479), .A0 (nx15435), .A1 (nx18333)) ;
    nor02ii ix93 (.Y (nx92), .A0 (nx15486), .A1 (nx12873)) ;
    and04 ix15487 (.Y (nx15486), .A0 (nflt_layer_out_0), .A1 (nx15500), .A2 (
          nx15512), .A3 (nx18165)) ;
    inv01 ix18164 (.Y (nx18165), .A (nflt_layer_out_3)) ;
    mux21 ix15492 (.Y (nx15491), .A0 (nx15488), .A1 (mem_data_in[0]), .S0 (
          nx17893)) ;
    nor02ii ix15497 (.Y (nx15496), .A0 (nx17893), .A1 (nx18265)) ;
    and02 ix15507 (.Y (nx15506), .A0 (nx15488), .A1 (nx15500)) ;
    xor2 ix15517 (.Y (nx15516), .A0 (nx15512), .A1 (nx15506)) ;
    and03 ix15526 (.Y (nx15525), .A0 (nx15488), .A1 (nx15500), .A2 (nx15512)) ;
    and03 ix15534 (.Y (nx15533), .A0 (nx15445), .A1 (nx15435), .A2 (nx19302)) ;
    nor02ii ix15547 (.Y (nx15546), .A0 (nx18151), .A1 (layer_type_out_1)) ;
    ao32 ix1479 (.Y (nx1478), .A0 (nx15575), .A1 (current_state_15), .A2 (
         nx15883), .B0 (current_state_16), .B1 (ftc_cntrl_reg_out_11)) ;
    or02 ix15562 (.Y (nx15561), .A0 (ftc_cntrl_reg_out_14), .A1 (nx18305)) ;
    xor2 ix279 (.Y (nx278), .A0 (nx18257), .A1 (cntr1_inst_counter_out_2)) ;
    xnor2 ix277 (.Y (nx276), .A0 (nx18257), .A1 (nx15586)) ;
    mux21 ix13022 (.Y (nx13021), .A0 (nx15588), .A1 (nx15586), .S0 (nx18257)) ;
    xor2 ix15589 (.Y (nx15588), .A0 (nx15586), .A1 (nx12882)) ;
    nor02ii ix269 (.Y (nx12882), .A0 (nx15402), .A1 (cntr1_inst_counter_out_4)
            ) ;
    xnor2 ix15597 (.Y (nx15596), .A0 (nx18257), .A1 (cntr1_inst_counter_out_1)
          ) ;
    nor02ii ix15603 (.Y (nx15602), .A0 (nx12912), .A1 (nx15861)) ;
    nor02ii ix1847 (.Y (nx12912), .A0 (nx15605), .A1 (nx15621)) ;
    and04 ix1403 (.Y (nx1402), .A0 (nx15614), .A1 (nx16070), .A2 (nx16079), .A3 (
          nx16084)) ;
    mux21 ix13842 (.Y (nx13841), .A0 (nx16067), .A1 (nx15614), .S0 (nx18289)) ;
    nor02ii ix349 (.Y (nx12883), .A0 (nx18279), .A1 (nx15859)) ;
    and04 ix15631 (.Y (nx15630), .A0 (nx16153), .A1 (nx15861), .A2 (nx15888), .A3 (
          nx15970)) ;
    xor2 ix15641 (.Y (nx15640), .A0 (nx15776), .A1 (new_size_squared_out_15)) ;
    xor2 ix15645 (.Y (nx15644), .A0 (nx15776), .A1 (nx1088)) ;
    nor02ii ix1089 (.Y (nx1088), .A0 (nx15653), .A1 (write_offset_data_out_14)
            ) ;
    ao22 ix13632 (.Y (nx13631), .A0 (nx1094), .A1 (nx18229), .B0 (
         write_offset_data_out_14), .B1 (nx18329)) ;
    nor02ii ix1043 (.Y (nx1042), .A0 (nx15666), .A1 (write_offset_data_out_12)
            ) ;
    ao22 ix13592 (.Y (nx13591), .A0 (nx1048), .A1 (nx18229), .B0 (
         write_offset_data_out_12), .B1 (nx18329)) ;
    nor02ii ix995 (.Y (nx994), .A0 (nx15679), .A1 (write_offset_data_out_10)) ;
    ao22 ix13552 (.Y (nx13551), .A0 (nx1000), .A1 (nx18229), .B0 (
         write_offset_data_out_10), .B1 (nx18329)) ;
    nor02ii ix949 (.Y (nx948), .A0 (nx15692), .A1 (write_offset_data_out_8)) ;
    ao22 ix13512 (.Y (nx13511), .A0 (nx954), .A1 (nx18231), .B0 (
         write_offset_data_out_8), .B1 (nx18329)) ;
    nor02ii ix763 (.Y (nx17945), .A0 (nx18231), .A1 (nx15537)) ;
    nand02 ix15700 (.Y (nx760), .A0 (nx15541), .A1 (nx15716)) ;
    nor02_2x ix1525 (.Y (nx1524), .A0 (nx15541), .A1 (nx18305)) ;
    nor02ii ix899 (.Y (nx898), .A0 (nx15726), .A1 (write_offset_data_out_6)) ;
    ao22 ix13472 (.Y (nx13471), .A0 (nx904), .A1 (nx18231), .B0 (
         write_offset_data_out_6), .B1 (nx18329)) ;
    nor02ii ix853 (.Y (nx852), .A0 (nx15741), .A1 (write_offset_data_out_4)) ;
    ao22 ix13432 (.Y (nx13431), .A0 (write_offset_data_out_4), .A1 (nx18331), .B0 (
         nx858), .B1 (nx18231)) ;
    or04 ix15742 (.Y (nx15741), .A0 (nx15745), .A1 (nx15750), .A2 (nx15756), .A3 (
         nx15763)) ;
    ao22 ix13412 (.Y (nx13411), .A0 (write_offset_data_out_3), .A1 (nx18331), .B0 (
         nx832), .B1 (nx18231)) ;
    mux21_ni ix13352 (.Y (nx13351), .A0 (nx18331), .A1 (nx18231), .S0 (nx15763)
             ) ;
    or02 ix15766 (.Y (nx15765), .A0 (nx15756), .A1 (nx15763)) ;
    or03 ix15769 (.Y (nx15768), .A0 (nx15750), .A1 (nx15756), .A2 (nx15763)) ;
    mux21_ni ix13662 (.Y (nx13661), .A0 (mem_data_in[15]), .A1 (
             new_size_squared_out_15), .S0 (nx18323)) ;
    xnor2 ix15782 (.Y (nx15781), .A0 (nx15647), .A1 (nx15785)) ;
    mux21_ni ix13642 (.Y (nx13641), .A0 (mem_data_in[14]), .A1 (
             new_size_squared_out_14), .S0 (nx18323)) ;
    xor2 ix15787 (.Y (nx15786), .A0 (nx15774), .A1 (new_size_squared_out_13)) ;
    mux21_ni ix13622 (.Y (nx13621), .A0 (mem_data_in[13]), .A1 (
             new_size_squared_out_13), .S0 (nx18323)) ;
    xnor2 ix15792 (.Y (nx15791), .A0 (nx15660), .A1 (nx15795)) ;
    mux21_ni ix13602 (.Y (nx13601), .A0 (mem_data_in[12]), .A1 (
             new_size_squared_out_12), .S0 (nx18323)) ;
    xor2 ix15798 (.Y (nx15797), .A0 (nx15772), .A1 (new_size_squared_out_11)) ;
    mux21_ni ix13582 (.Y (nx13581), .A0 (mem_data_in[11]), .A1 (
             new_size_squared_out_11), .S0 (nx18323)) ;
    xnor2 ix15803 (.Y (nx15802), .A0 (nx15673), .A1 (nx15806)) ;
    mux21_ni ix13562 (.Y (nx13561), .A0 (mem_data_in[10]), .A1 (
             new_size_squared_out_10), .S0 (nx18323)) ;
    xor2 ix15808 (.Y (nx15807), .A0 (nx15770), .A1 (new_size_squared_out_9)) ;
    mux21_ni ix13542 (.Y (nx13541), .A0 (mem_data_in[9]), .A1 (
             new_size_squared_out_9), .S0 (nx18325)) ;
    xnor2 ix15813 (.Y (nx15812), .A0 (nx15686), .A1 (nx15816)) ;
    mux21_ni ix13522 (.Y (nx13521), .A0 (mem_data_in[8]), .A1 (
             new_size_squared_out_8), .S0 (nx18325)) ;
    xor2 ix15819 (.Y (nx15818), .A0 (nx15696), .A1 (new_size_squared_out_7)) ;
    mux21_ni ix13502 (.Y (nx13501), .A0 (mem_data_in[7]), .A1 (
             new_size_squared_out_7), .S0 (nx18325)) ;
    xnor2 ix15824 (.Y (nx15823), .A0 (nx15720), .A1 (nx15827)) ;
    mux21_ni ix13482 (.Y (nx13481), .A0 (mem_data_in[6]), .A1 (
             new_size_squared_out_6), .S0 (nx18325)) ;
    xor2 ix15829 (.Y (nx15828), .A0 (nx15730), .A1 (new_size_squared_out_5)) ;
    mux21_ni ix13462 (.Y (nx13461), .A0 (mem_data_in[5]), .A1 (
             new_size_squared_out_5), .S0 (nx18325)) ;
    xnor2 ix15834 (.Y (nx15833), .A0 (nx15735), .A1 (nx15837)) ;
    mux21_ni ix13442 (.Y (nx13441), .A0 (mem_data_in[4]), .A1 (
             new_size_squared_out_4), .S0 (nx18325)) ;
    xor2 ix15840 (.Y (nx15839), .A0 (nx15745), .A1 (new_size_squared_out_3)) ;
    mux21_ni ix13422 (.Y (nx13421), .A0 (mem_data_in[3]), .A1 (
             new_size_squared_out_3), .S0 (nx18325)) ;
    xnor2 ix15845 (.Y (nx15844), .A0 (nx15750), .A1 (nx15848)) ;
    mux21_ni ix13402 (.Y (nx13401), .A0 (mem_data_in[2]), .A1 (
             new_size_squared_out_2), .S0 (nx18327)) ;
    xor2 ix15850 (.Y (nx15849), .A0 (nx15756), .A1 (new_size_squared_out_1)) ;
    mux21_ni ix13382 (.Y (nx13381), .A0 (mem_data_in[1]), .A1 (
             new_size_squared_out_1), .S0 (nx18327)) ;
    xor2 ix15855 (.Y (nx15854), .A0 (nx15763), .A1 (new_size_squared_out_0)) ;
    mux21_ni ix13362 (.Y (nx13361), .A0 (mem_data_in[0]), .A1 (
             new_size_squared_out_0), .S0 (nx18327)) ;
    or02 ix577 (.Y (nx576), .A0 (ftc_cntrl_reg_out_11), .A1 (nx15888)) ;
    and04 ix551 (.Y (nx550), .A0 (nx15873), .A1 (nx15893), .A2 (nx15902), .A3 (
          nx15907)) ;
    mux21 ix13222 (.Y (nx13221), .A0 (nx15890), .A1 (nx15873), .S0 (nx18283)) ;
    or03 ix15879 (.Y (nx15878), .A0 (ftc_cntrl_reg_out_8), .A1 (nx15861), .A2 (
         nx15883)) ;
    ao21 ix1147 (.Y (nx1146), .A0 (nx18279), .A1 (nx15605), .B0 (
         current_state_16)) ;
    xor2 ix15891 (.Y (nx15890), .A0 (nx15873), .A1 (nx12885)) ;
    nor02ii ix531 (.Y (nx12885), .A0 (nx15898), .A1 (
            window_width_cntr_counter_out_14)) ;
    mux21_ni ix13212 (.Y (nx13211), .A0 (nx524), .A1 (
             window_width_cntr_counter_out_14), .S0 (nx18283)) ;
    xor2 ix525 (.Y (nx524), .A0 (nx15893), .A1 (nx15898)) ;
    mux21 ix13202 (.Y (nx13201), .A0 (nx15904), .A1 (nx15902), .S0 (nx18283)) ;
    nor02ii ix507 (.Y (nx12887), .A0 (nx15912), .A1 (
            window_width_cntr_counter_out_12)) ;
    mux21_ni ix13192 (.Y (nx13191), .A0 (nx500), .A1 (
             window_width_cntr_counter_out_12), .S0 (nx18283)) ;
    xor2 ix501 (.Y (nx500), .A0 (nx15907), .A1 (nx15912)) ;
    mux21 ix13182 (.Y (nx13181), .A0 (nx15918), .A1 (nx15916), .S0 (nx18283)) ;
    nor02ii ix483 (.Y (nx12889), .A0 (nx15926), .A1 (
            window_width_cntr_counter_out_10)) ;
    mux21_ni ix13172 (.Y (nx13171), .A0 (nx476), .A1 (
             window_width_cntr_counter_out_10), .S0 (nx18283)) ;
    xor2 ix477 (.Y (nx476), .A0 (nx15921), .A1 (nx15926)) ;
    mux21 ix13162 (.Y (nx13161), .A0 (nx15932), .A1 (nx15930), .S0 (nx18283)) ;
    nor02ii ix459 (.Y (nx12891), .A0 (nx15940), .A1 (
            window_width_cntr_counter_out_8)) ;
    mux21_ni ix13152 (.Y (nx13151), .A0 (nx452), .A1 (
             window_width_cntr_counter_out_8), .S0 (nx18285)) ;
    xor2 ix453 (.Y (nx452), .A0 (nx15935), .A1 (nx15940)) ;
    mux21 ix13142 (.Y (nx13141), .A0 (nx15946), .A1 (nx15944), .S0 (nx18285)) ;
    nor02ii ix435 (.Y (nx12893), .A0 (nx15954), .A1 (
            window_width_cntr_counter_out_6)) ;
    mux21_ni ix13132 (.Y (nx13131), .A0 (nx428), .A1 (
             window_width_cntr_counter_out_6), .S0 (nx18285)) ;
    xor2 ix429 (.Y (nx428), .A0 (nx15949), .A1 (nx15954)) ;
    or03 ix15955 (.Y (nx15954), .A0 (nx18167), .A1 (nx15995), .A2 (nx15959)) ;
    inv01 ix18166 (.Y (nx18167), .A (wind_width_count_4)) ;
    mux21_ni ix14042 (.Y (nx14041), .A0 (nx1876), .A1 (wind_width_count_4), .S0 (
             nx18285)) ;
    mux21_ni ix13092 (.Y (nx13091), .A0 (nx384), .A1 (wind_width_count_1), .S0 (
             nx18285)) ;
    xor2 ix13082 (.Y (nx13081), .A0 (nx17811), .A1 (nx12884)) ;
    mux21_ni ix13102 (.Y (nx13101), .A0 (nx392), .A1 (wind_width_count_2), .S0 (
             nx18285)) ;
    mux21_ni ix13112 (.Y (nx13111), .A0 (nx400), .A1 (wind_width_count_3), .S0 (
             nx18285)) ;
    mux21 ix13122 (.Y (nx13121), .A0 (nx15997), .A1 (nx15995), .S0 (nx18287)) ;
    and04 ix565 (.Y (nx564), .A0 (nx15916), .A1 (nx15921), .A2 (nx15930), .A3 (
          nx15935)) ;
    and04 ix613 (.Y (nx612), .A0 (nx15944), .A1 (nx15949), .A2 (nx15995), .A3 (
          nx18169)) ;
    inv01 ix18168 (.Y (nx18169), .A (nx604)) ;
    mux21 ix603 (.Y (nx602), .A0 (nx18305), .A1 (img_width_out_0), .S0 (nx18225)
          ) ;
    ao221 ix13242 (.Y (nx13241), .A0 (img_width_out_0), .A1 (nx18259), .B0 (
          nx18911), .B1 (new_width_out_0), .C0 (nx17897)) ;
    mux21 ix641 (.Y (nx640), .A0 (nx18305), .A1 (nx16189), .S0 (nx18225)) ;
    ao22 ix13262 (.Y (nx13261), .A0 (img_width_out_1), .A1 (nx18261), .B0 (
         nx18911), .B1 (new_width_out_1)) ;
    nor02ii ix705 (.Y (nx704), .A0 (nx16042), .A1 (nx18225)) ;
    xor2 ix16043 (.Y (nx16042), .A0 (nx16046), .A1 (nx16037)) ;
    ao22 ix13302 (.Y (nx13301), .A0 (img_width_out_3), .A1 (nx18261), .B0 (
         nx18911), .B1 (new_width_out_3)) ;
    nor02ii ix723 (.Y (nx722), .A0 (nx16055), .A1 (nx18227)) ;
    and04 ix16064 (.Y (nx16063), .A0 (nx16005), .A1 (nx16019), .A2 (nx18171), .A3 (
          nx16046)) ;
    inv01 ix18170 (.Y (nx18171), .A (img_width_out_2)) ;
    or02 ix16066 (.Y (nx16065), .A0 (nx15605), .A1 (nx15621)) ;
    xor2 ix16068 (.Y (nx16067), .A0 (nx15614), .A1 (nx12896)) ;
    nor02ii ix1383 (.Y (nx12896), .A0 (nx16075), .A1 (
            cache_width_cntr_counter_out_14)) ;
    mux21_ni ix13832 (.Y (nx13831), .A0 (nx1376), .A1 (
             cache_width_cntr_counter_out_14), .S0 (nx18289)) ;
    xor2 ix1377 (.Y (nx1376), .A0 (nx16070), .A1 (nx16075)) ;
    mux21 ix13822 (.Y (nx13821), .A0 (nx16081), .A1 (nx16079), .S0 (nx18289)) ;
    nor02ii ix1359 (.Y (nx12898), .A0 (nx16089), .A1 (
            cache_width_cntr_counter_out_12)) ;
    mux21_ni ix13812 (.Y (nx13811), .A0 (nx1352), .A1 (
             cache_width_cntr_counter_out_12), .S0 (nx18289)) ;
    xor2 ix1353 (.Y (nx1352), .A0 (nx16084), .A1 (nx16089)) ;
    mux21 ix13802 (.Y (nx13801), .A0 (nx16095), .A1 (nx16093), .S0 (nx18289)) ;
    nor02ii ix1335 (.Y (nx12900), .A0 (nx16103), .A1 (
            cache_width_cntr_counter_out_10)) ;
    mux21_ni ix13792 (.Y (nx13791), .A0 (nx1328), .A1 (
             cache_width_cntr_counter_out_10), .S0 (nx18289)) ;
    xor2 ix1329 (.Y (nx1328), .A0 (nx16098), .A1 (nx16103)) ;
    mux21 ix13782 (.Y (nx13781), .A0 (nx16109), .A1 (nx16107), .S0 (nx18289)) ;
    nor02ii ix1311 (.Y (nx12902), .A0 (nx16117), .A1 (
            cache_width_cntr_counter_out_8)) ;
    mux21_ni ix13772 (.Y (nx13771), .A0 (nx1304), .A1 (
             cache_width_cntr_counter_out_8), .S0 (nx18291)) ;
    xor2 ix1305 (.Y (nx1304), .A0 (nx16112), .A1 (nx16117)) ;
    mux21 ix13762 (.Y (nx13761), .A0 (nx16123), .A1 (nx16121), .S0 (nx18291)) ;
    nor02ii ix1287 (.Y (nx12904), .A0 (nx16131), .A1 (
            cache_width_cntr_counter_out_6)) ;
    mux21_ni ix13752 (.Y (nx13751), .A0 (nx1280), .A1 (
             cache_width_cntr_counter_out_6), .S0 (nx18291)) ;
    xor2 ix1281 (.Y (nx1280), .A0 (nx16126), .A1 (nx16131)) ;
    or03 ix16132 (.Y (nx16131), .A0 (nx18173), .A1 (nx16178), .A2 (nx16136)) ;
    inv01 ix18172 (.Y (nx18173), .A (nx17817)) ;
    mux21_ni ix13732 (.Y (nx13731), .A0 (nx1254), .A1 (nx17815), .S0 (nx18291)
             ) ;
    mux21_ni ix13702 (.Y (nx13701), .A0 (nx1230), .A1 (cache_width_count_1), .S0 (
             nx18291)) ;
    xor2 ix13692 (.Y (nx13691), .A0 (cache_width_count_0), .A1 (nx18383)) ;
    mux21_ni ix16151 (.Y (nx16150), .A0 (cache_height_count_en), .A1 (nx17871), 
             .S0 (nx18279)) ;
    and02 ix16154 (.Y (nx16153), .A0 (nx18279), .A1 (nx15605)) ;
    nor02ii ix1213 (.Y (nx1212), .A0 (nx16155), .A1 (ftc_cntrl_reg_out_10)) ;
    mux21_ni ix13712 (.Y (nx13711), .A0 (nx1238), .A1 (nx17819), .S0 (nx18291)
             ) ;
    mux21_ni ix13722 (.Y (nx13721), .A0 (nx1246), .A1 (cache_width_count_3), .S0 (
             nx18291)) ;
    mux21 ix13742 (.Y (nx13741), .A0 (nx16180), .A1 (nx16178), .S0 (nx18293)) ;
    and04 ix1417 (.Y (nx1416), .A0 (nx16093), .A1 (nx16098), .A2 (nx16107), .A3 (
          nx16112)) ;
    and04 ix1435 (.Y (nx1434), .A0 (nx16121), .A1 (nx16126), .A2 (nx16178), .A3 (
          nx18175)) ;
    xnor2 ix1427 (.Y (nx18175), .A0 (nx16005), .A1 (cache_width_count_0)) ;
    xor2 ix1437 (.Y (nx1436), .A0 (cache_width_count_1), .A1 (nx636)) ;
    and02 ix16192 (.Y (nx16191), .A0 (nx16005), .A1 (nx16019)) ;
    nor02_2x ix1485 (.Y (nx1484), .A0 (nx18273), .A1 (nx18307)) ;
    and02 ix1867 (.Y (nx12906), .A0 (current_state_21), .A1 (nx15865)) ;
    and02 ix16223 (.Y (nx16222), .A0 (nx18265), .A1 (nx18333)) ;
    nor02ii ix16227 (.Y (nx16226), .A0 (num_channels_counter_out_1), .A1 (
            nx15531)) ;
    mux21 ix1765 (.Y (nx1764), .A0 (nx15508), .A1 (nx16274), .S0 (nx15445)) ;
    mux21 ix16281 (.Y (nx16280), .A0 (mem_data_in[0]), .A1 (nx16278), .S0 (
          nx15445)) ;
    and02 ix16283 (.Y (nx16282), .A0 (nx15445), .A1 (nx18333)) ;
    nor02ii ix16285 (.Y (nx16284), .A0 (nlayers_counter_out_1), .A1 (nx16278)) ;
    mux21 ix1781 (.Y (nx1780), .A0 (nx15518), .A1 (nx16290), .S0 (nx15445)) ;
    or02 ix309 (.Y (nx308), .A0 (nx18307), .A1 (nx18257)) ;
    nor02ii ix16322 (.Y (argmax_ready), .A0 (nx16327), .A1 (nx1926)) ;
    or04 ix1927 (.Y (nx1926), .A0 (class_cntr_counter_out_0), .A1 (nx16332), .A2 (
         class_cntr_counter_out_2), .A3 (nx18887)) ;
    mux21 ix14052 (.Y (nx14051), .A0 (current_state_27), .A1 (nx18339), .S0 (
          nx16324)) ;
    mux21 ix14062 (.Y (nx14061), .A0 (nx16334), .A1 (nx16332), .S0 (nx18339)) ;
    or02 ix16337 (.Y (nx16336), .A0 (nx16332), .A1 (nx16324)) ;
    mux21_ni ix14072 (.Y (nx14071), .A0 (nx1904), .A1 (class_cntr_counter_out_2)
             , .S0 (nx18339)) ;
    xor2 ix1905 (.Y (nx1904), .A0 (nx16338), .A1 (nx16336)) ;
    mux21_ni ix14082 (.Y (nx14081), .A0 (nx1912), .A1 (class_cntr_counter_out_3)
             , .S0 (nx18341)) ;
    xor2 ix1913 (.Y (nx1912), .A0 (nx18887), .A1 (nx16346)) ;
    or03 ix16347 (.Y (nx16346), .A0 (nx16338), .A1 (nx16332), .A2 (nx16324)) ;
    nor02ii ix4917 (.Y (argmax_data_out[0]), .A0 (nx18341), .A1 (mem_data_in[0])
            ) ;
    nor02ii ix4919 (.Y (argmax_data_out[1]), .A0 (nx18341), .A1 (mem_data_in[1])
            ) ;
    nor02ii ix4921 (.Y (argmax_data_out[2]), .A0 (nx18341), .A1 (mem_data_in[2])
            ) ;
    nor02ii ix4923 (.Y (argmax_data_out[3]), .A0 (nx18341), .A1 (mem_data_in[3])
            ) ;
    nor02ii ix4925 (.Y (argmax_data_out[4]), .A0 (nx18341), .A1 (mem_data_in[4])
            ) ;
    nor02ii ix4927 (.Y (argmax_data_out[5]), .A0 (nx18341), .A1 (mem_data_in[5])
            ) ;
    nor02ii ix4929 (.Y (argmax_data_out[6]), .A0 (nx18343), .A1 (mem_data_in[6])
            ) ;
    nor02ii ix4931 (.Y (argmax_data_out[7]), .A0 (nx18343), .A1 (mem_data_in[7])
            ) ;
    nor02ii ix4933 (.Y (argmax_data_out[8]), .A0 (nx18343), .A1 (mem_data_in[8])
            ) ;
    nor02ii ix4935 (.Y (argmax_data_out[9]), .A0 (nx18343), .A1 (mem_data_in[9])
            ) ;
    nor02ii ix4937 (.Y (argmax_data_out[10]), .A0 (nx18343), .A1 (
            mem_data_in[10])) ;
    nor02ii ix4939 (.Y (argmax_data_out[11]), .A0 (nx18343), .A1 (
            mem_data_in[11])) ;
    nor02ii ix4941 (.Y (argmax_data_out[12]), .A0 (nx18343), .A1 (
            mem_data_in[12])) ;
    nor02ii ix4943 (.Y (argmax_data_out[13]), .A0 (nx18345), .A1 (
            mem_data_in[13])) ;
    nor02ii ix4945 (.Y (argmax_data_out[14]), .A0 (nx18345), .A1 (
            mem_data_in[14])) ;
    nor02ii ix4947 (.Y (argmax_data_out[15]), .A0 (nx18345), .A1 (
            mem_data_in[15])) ;
    and02 ix4949 (.Y (comp_unit_data2_out[0]), .A0 (nx18233), .A1 (nx2140)) ;
    mux21_ni ix2141 (.Y (nx2140), .A0 (flt_bias_out_0), .A1 (mem_data_in[0]), .S0 (
             nx18297)) ;
    and02 ix4951 (.Y (comp_unit_data2_out[1]), .A0 (nx18233), .A1 (nx2168)) ;
    mux21_ni ix2169 (.Y (nx2168), .A0 (flt_bias_out_1), .A1 (mem_data_in[1]), .S0 (
             nx18297)) ;
    and02 ix4953 (.Y (comp_unit_data2_out[2]), .A0 (nx18235), .A1 (nx2194)) ;
    mux21_ni ix2195 (.Y (nx2194), .A0 (flt_bias_out_2), .A1 (mem_data_in[2]), .S0 (
             nx18297)) ;
    and02 ix4955 (.Y (comp_unit_data2_out[3]), .A0 (nx18235), .A1 (nx2220)) ;
    mux21_ni ix2221 (.Y (nx2220), .A0 (flt_bias_out_3), .A1 (mem_data_in[3]), .S0 (
             nx18297)) ;
    and02 ix4957 (.Y (comp_unit_data2_out[4]), .A0 (nx18235), .A1 (nx2246)) ;
    mux21_ni ix2247 (.Y (nx2246), .A0 (flt_bias_out_4), .A1 (mem_data_in[4]), .S0 (
             nx18297)) ;
    and02 ix4959 (.Y (comp_unit_data2_out[5]), .A0 (nx18235), .A1 (nx2272)) ;
    mux21_ni ix2273 (.Y (nx2272), .A0 (flt_bias_out_5), .A1 (mem_data_in[5]), .S0 (
             nx18299)) ;
    and02 ix4961 (.Y (comp_unit_data2_out[6]), .A0 (nx18235), .A1 (nx2298)) ;
    mux21_ni ix2299 (.Y (nx2298), .A0 (flt_bias_out_6), .A1 (mem_data_in[6]), .S0 (
             nx18299)) ;
    and02 ix4963 (.Y (comp_unit_data2_out[7]), .A0 (nx18235), .A1 (nx2324)) ;
    mux21_ni ix2325 (.Y (nx2324), .A0 (flt_bias_out_7), .A1 (mem_data_in[7]), .S0 (
             nx18299)) ;
    and02 ix4965 (.Y (comp_unit_data2_out[8]), .A0 (nx18235), .A1 (nx2350)) ;
    mux21_ni ix2351 (.Y (nx2350), .A0 (flt_bias_out_8), .A1 (mem_data_in[8]), .S0 (
             nx18299)) ;
    and02 ix4967 (.Y (comp_unit_data2_out[9]), .A0 (nx18237), .A1 (nx2376)) ;
    mux21_ni ix2377 (.Y (nx2376), .A0 (flt_bias_out_9), .A1 (mem_data_in[9]), .S0 (
             nx18299)) ;
    and02 ix4969 (.Y (comp_unit_data2_out[10]), .A0 (nx18237), .A1 (nx2402)) ;
    mux21_ni ix2403 (.Y (nx2402), .A0 (flt_bias_out_10), .A1 (mem_data_in[10]), 
             .S0 (nx18299)) ;
    and02 ix4971 (.Y (comp_unit_data2_out[11]), .A0 (nx18237), .A1 (nx2428)) ;
    mux21_ni ix2429 (.Y (nx2428), .A0 (flt_bias_out_11), .A1 (mem_data_in[11]), 
             .S0 (nx18299)) ;
    and02 ix4973 (.Y (comp_unit_data2_out[12]), .A0 (nx18237), .A1 (nx2454)) ;
    mux21_ni ix2455 (.Y (nx2454), .A0 (flt_bias_out_12), .A1 (mem_data_in[12]), 
             .S0 (nx18301)) ;
    and02 ix4975 (.Y (comp_unit_data2_out[13]), .A0 (nx18237), .A1 (nx2480)) ;
    mux21_ni ix2481 (.Y (nx2480), .A0 (flt_bias_out_13), .A1 (mem_data_in[13]), 
             .S0 (nx18301)) ;
    and02 ix4977 (.Y (comp_unit_data2_out[14]), .A0 (nx18237), .A1 (nx2506)) ;
    mux21_ni ix2507 (.Y (nx2506), .A0 (flt_bias_out_14), .A1 (mem_data_in[14]), 
             .S0 (nx18301)) ;
    and02 ix4979 (.Y (comp_unit_data2_out[15]), .A0 (nx18237), .A1 (nx2532)) ;
    mux21_ni ix2533 (.Y (nx2532), .A0 (flt_bias_out_15), .A1 (mem_data_in[15]), 
             .S0 (nx18301)) ;
    and03 ix5147 (.Y (max_height_1), .A0 (nx636), .A1 (nx17803), .A2 (nx18281)
          ) ;
    or03 ix16456 (.Y (nx16455), .A0 (nx18307), .A1 (nx15605), .A2 (nx16463)) ;
    ao21 ix16466 (.Y (nx2580), .A0 (nx16463), .A1 (nx12912), .B0 (nx1182)) ;
    and02 ix2583 (.Y (cache_data_in_0), .A0 (mem_data_in[0]), .A1 (nx18243)) ;
    and02 ix2585 (.Y (cache_data_in_1), .A0 (mem_data_in[1]), .A1 (nx18243)) ;
    and02 ix2587 (.Y (cache_data_in_2), .A0 (mem_data_in[2]), .A1 (nx18243)) ;
    and02 ix2589 (.Y (cache_data_in_3), .A0 (mem_data_in[3]), .A1 (nx18245)) ;
    and02 ix2591 (.Y (cache_data_in_4), .A0 (mem_data_in[4]), .A1 (nx18245)) ;
    and02 ix2593 (.Y (cache_data_in_5), .A0 (mem_data_in[5]), .A1 (nx18245)) ;
    and02 ix2595 (.Y (cache_data_in_6), .A0 (mem_data_in[6]), .A1 (nx18245)) ;
    and02 ix2597 (.Y (cache_data_in_7), .A0 (mem_data_in[7]), .A1 (nx18245)) ;
    and02 ix2599 (.Y (cache_data_in_8), .A0 (mem_data_in[8]), .A1 (nx18245)) ;
    and02 ix2601 (.Y (cache_data_in_9), .A0 (mem_data_in[9]), .A1 (nx18245)) ;
    and02 ix2603 (.Y (cache_data_in_10), .A0 (mem_data_in[10]), .A1 (nx18247)) ;
    and02 ix2605 (.Y (cache_data_in_11), .A0 (mem_data_in[11]), .A1 (nx18247)) ;
    and02 ix2607 (.Y (cache_data_in_12), .A0 (mem_data_in[12]), .A1 (nx18247)) ;
    and02 ix2609 (.Y (cache_data_in_13), .A0 (mem_data_in[13]), .A1 (nx18247)) ;
    and02 ix2611 (.Y (cache_data_in_14), .A0 (mem_data_in[14]), .A1 (nx18247)) ;
    and02 ix2613 (.Y (cache_data_in_15), .A0 (mem_data_in[15]), .A1 (nx18247)) ;
    and02 ix16508 (.Y (nx16507), .A0 (nx17803), .A1 (nx18281)) ;
    mux21 ix14112 (.Y (nx14111), .A0 (nx16514), .A1 (nx16511), .S0 (nx18273)) ;
    mux21 ix14132 (.Y (nx14131), .A0 (nx16521), .A1 (nx16518), .S0 (nx18273)) ;
    mux21 ix14152 (.Y (nx14151), .A0 (nx16527), .A1 (nx16524), .S0 (nx18273)) ;
    mux21 ix14172 (.Y (nx14171), .A0 (nx16533), .A1 (nx16530), .S0 (nx18273)) ;
    mux21 ix14192 (.Y (nx14191), .A0 (nx16539), .A1 (nx16536), .S0 (nx18275)) ;
    mux21 ix14212 (.Y (nx14211), .A0 (nx16545), .A1 (nx16542), .S0 (nx18275)) ;
    mux21 ix14232 (.Y (nx14231), .A0 (nx16551), .A1 (nx16548), .S0 (nx18275)) ;
    mux21 ix14252 (.Y (nx14251), .A0 (nx16557), .A1 (nx16554), .S0 (nx18275)) ;
    mux21 ix14272 (.Y (nx14271), .A0 (nx16563), .A1 (nx16560), .S0 (nx18275)) ;
    mux21 ix14292 (.Y (nx14291), .A0 (nx16569), .A1 (nx16566), .S0 (nx18275)) ;
    mux21 ix14312 (.Y (nx14311), .A0 (nx16575), .A1 (nx16572), .S0 (nx18275)) ;
    mux21 ix14332 (.Y (nx14331), .A0 (nx16581), .A1 (nx16578), .S0 (nx18277)) ;
    mux21 ix14352 (.Y (nx14351), .A0 (nx16587), .A1 (nx16584), .S0 (nx18277)) ;
    mux21 ix14372 (.Y (nx14371), .A0 (nx16593), .A1 (nx16590), .S0 (nx18277)) ;
    mux21 ix14392 (.Y (nx14391), .A0 (nx16599), .A1 (nx16596), .S0 (nx18277)) ;
    mux21 ix14412 (.Y (nx14411), .A0 (nx16605), .A1 (nx16602), .S0 (nx18277)) ;
    nor02ii ix4885 (.Y (filter_data_out[0]), .A0 (nx18319), .A1 (mem_data_in[0])
            ) ;
    nor02ii ix4887 (.Y (filter_data_out[1]), .A0 (nx18319), .A1 (mem_data_in[1])
            ) ;
    nor02ii ix4889 (.Y (filter_data_out[2]), .A0 (nx18319), .A1 (mem_data_in[2])
            ) ;
    nor02ii ix4891 (.Y (filter_data_out[3]), .A0 (nx18319), .A1 (mem_data_in[3])
            ) ;
    nor02ii ix4893 (.Y (filter_data_out[4]), .A0 (nx18319), .A1 (mem_data_in[4])
            ) ;
    nor02ii ix4895 (.Y (filter_data_out[5]), .A0 (nx18321), .A1 (mem_data_in[5])
            ) ;
    nor02ii ix4897 (.Y (filter_data_out[6]), .A0 (nx18321), .A1 (mem_data_in[6])
            ) ;
    nor02ii ix4899 (.Y (filter_data_out[7]), .A0 (nx18321), .A1 (mem_data_in[7])
            ) ;
    nor02ii ix4901 (.Y (filter_data_out[8]), .A0 (nx18321), .A1 (mem_data_in[8])
            ) ;
    nor02ii ix4903 (.Y (filter_data_out[9]), .A0 (nx18321), .A1 (mem_data_in[9])
            ) ;
    nor02ii ix4905 (.Y (filter_data_out[10]), .A0 (nx18321), .A1 (
            mem_data_in[10])) ;
    nor02ii ix4907 (.Y (filter_data_out[11]), .A0 (nx18321), .A1 (
            mem_data_in[11])) ;
    nor02ii ix4909 (.Y (filter_data_out[12]), .A0 (nx17863), .A1 (
            mem_data_in[12])) ;
    nor02ii ix4911 (.Y (filter_data_out[13]), .A0 (nx17863), .A1 (
            mem_data_in[13])) ;
    nor02ii ix4913 (.Y (filter_data_out[14]), .A0 (nx17863), .A1 (
            mem_data_in[14])) ;
    nor02ii ix4915 (.Y (filter_data_out[15]), .A0 (nx17863), .A1 (
            mem_data_in[15])) ;
    and02 ix4981 (.Y (wind_col_in_0__0), .A0 (nx18359), .A1 (cache_data_out_0__0
          )) ;
    and02 ix4983 (.Y (wind_col_in_0__1), .A0 (nx18359), .A1 (cache_data_out_0__1
          )) ;
    and02 ix4985 (.Y (wind_col_in_0__2), .A0 (nx18359), .A1 (cache_data_out_0__2
          )) ;
    and02 ix4987 (.Y (wind_col_in_0__3), .A0 (nx18359), .A1 (cache_data_out_0__3
          )) ;
    and02 ix4989 (.Y (wind_col_in_0__4), .A0 (nx18359), .A1 (cache_data_out_0__4
          )) ;
    and02 ix4991 (.Y (wind_col_in_0__5), .A0 (nx18359), .A1 (cache_data_out_0__5
          )) ;
    and02 ix4993 (.Y (wind_col_in_0__6), .A0 (nx18359), .A1 (cache_data_out_0__6
          )) ;
    and02 ix4995 (.Y (wind_col_in_0__7), .A0 (nx18361), .A1 (cache_data_out_0__7
          )) ;
    and02 ix4997 (.Y (wind_col_in_0__8), .A0 (nx18361), .A1 (cache_data_out_0__8
          )) ;
    and02 ix4999 (.Y (wind_col_in_0__9), .A0 (nx18361), .A1 (cache_data_out_0__9
          )) ;
    and02 ix5001 (.Y (wind_col_in_0__10), .A0 (nx18361), .A1 (
          cache_data_out_0__10)) ;
    and02 ix5003 (.Y (wind_col_in_0__11), .A0 (nx18361), .A1 (
          cache_data_out_0__11)) ;
    and02 ix5005 (.Y (wind_col_in_0__12), .A0 (nx18361), .A1 (
          cache_data_out_0__12)) ;
    and02 ix5007 (.Y (wind_col_in_0__13), .A0 (nx18361), .A1 (
          cache_data_out_0__13)) ;
    and02 ix5009 (.Y (wind_col_in_0__14), .A0 (nx18363), .A1 (
          cache_data_out_0__14)) ;
    and02 ix5011 (.Y (wind_col_in_0__15), .A0 (nx18363), .A1 (
          cache_data_out_0__15)) ;
    and02 ix5013 (.Y (wind_col_in_1__0), .A0 (nx18363), .A1 (cache_data_out_1__0
          )) ;
    and02 ix5015 (.Y (wind_col_in_1__1), .A0 (nx18363), .A1 (cache_data_out_1__1
          )) ;
    and02 ix5017 (.Y (wind_col_in_1__2), .A0 (nx18363), .A1 (cache_data_out_1__2
          )) ;
    and02 ix5019 (.Y (wind_col_in_1__3), .A0 (nx18363), .A1 (cache_data_out_1__3
          )) ;
    and02 ix5021 (.Y (wind_col_in_1__4), .A0 (nx18363), .A1 (cache_data_out_1__4
          )) ;
    and02 ix5023 (.Y (wind_col_in_1__5), .A0 (nx18365), .A1 (cache_data_out_1__5
          )) ;
    and02 ix5025 (.Y (wind_col_in_1__6), .A0 (nx18365), .A1 (cache_data_out_1__6
          )) ;
    and02 ix5027 (.Y (wind_col_in_1__7), .A0 (nx18365), .A1 (cache_data_out_1__7
          )) ;
    and02 ix5029 (.Y (wind_col_in_1__8), .A0 (nx18365), .A1 (cache_data_out_1__8
          )) ;
    and02 ix5031 (.Y (wind_col_in_1__9), .A0 (nx18365), .A1 (cache_data_out_1__9
          )) ;
    and02 ix5033 (.Y (wind_col_in_1__10), .A0 (nx18365), .A1 (
          cache_data_out_1__10)) ;
    and02 ix5035 (.Y (wind_col_in_1__11), .A0 (nx18365), .A1 (
          cache_data_out_1__11)) ;
    and02 ix5037 (.Y (wind_col_in_1__12), .A0 (nx18367), .A1 (
          cache_data_out_1__12)) ;
    and02 ix5039 (.Y (wind_col_in_1__13), .A0 (nx18367), .A1 (
          cache_data_out_1__13)) ;
    and02 ix5041 (.Y (wind_col_in_1__14), .A0 (nx18367), .A1 (
          cache_data_out_1__14)) ;
    and02 ix5043 (.Y (wind_col_in_1__15), .A0 (nx18367), .A1 (
          cache_data_out_1__15)) ;
    and02 ix5045 (.Y (wind_col_in_2__0), .A0 (nx18367), .A1 (cache_data_out_2__0
          )) ;
    and02 ix5047 (.Y (wind_col_in_2__1), .A0 (nx18367), .A1 (cache_data_out_2__1
          )) ;
    and02 ix5049 (.Y (wind_col_in_2__2), .A0 (nx18367), .A1 (cache_data_out_2__2
          )) ;
    and02 ix5051 (.Y (wind_col_in_2__3), .A0 (nx18155), .A1 (cache_data_out_2__3
          )) ;
    and02 ix5053 (.Y (wind_col_in_2__4), .A0 (nx18155), .A1 (cache_data_out_2__4
          )) ;
    and02 ix5055 (.Y (wind_col_in_2__5), .A0 (nx18155), .A1 (cache_data_out_2__5
          )) ;
    and02 ix5057 (.Y (wind_col_in_2__6), .A0 (nx18155), .A1 (cache_data_out_2__6
          )) ;
    and02 ix5059 (.Y (wind_col_in_2__7), .A0 (nx18155), .A1 (cache_data_out_2__7
          )) ;
    and02 ix5061 (.Y (wind_col_in_2__8), .A0 (nx18155), .A1 (cache_data_out_2__8
          )) ;
    and02 ix5063 (.Y (wind_col_in_2__9), .A0 (nx18155), .A1 (cache_data_out_2__9
          )) ;
    and02 ix5065 (.Y (wind_col_in_2__10), .A0 (nx18369), .A1 (
          cache_data_out_2__10)) ;
    and02 ix5067 (.Y (wind_col_in_2__11), .A0 (nx18369), .A1 (
          cache_data_out_2__11)) ;
    and02 ix5069 (.Y (wind_col_in_2__12), .A0 (nx18369), .A1 (
          cache_data_out_2__12)) ;
    and02 ix5071 (.Y (wind_col_in_2__13), .A0 (nx18369), .A1 (
          cache_data_out_2__13)) ;
    and02 ix5073 (.Y (wind_col_in_2__14), .A0 (nx18369), .A1 (
          cache_data_out_2__14)) ;
    and02 ix5075 (.Y (wind_col_in_2__15), .A0 (nx18369), .A1 (
          cache_data_out_2__15)) ;
    and02 ix5077 (.Y (wind_col_in_3__0), .A0 (nx18369), .A1 (cache_data_out_3__0
          )) ;
    and02 ix5079 (.Y (wind_col_in_3__1), .A0 (nx18371), .A1 (cache_data_out_3__1
          )) ;
    and02 ix5081 (.Y (wind_col_in_3__2), .A0 (nx18371), .A1 (cache_data_out_3__2
          )) ;
    and02 ix5083 (.Y (wind_col_in_3__3), .A0 (nx18371), .A1 (cache_data_out_3__3
          )) ;
    and02 ix5085 (.Y (wind_col_in_3__4), .A0 (nx18371), .A1 (cache_data_out_3__4
          )) ;
    and02 ix5087 (.Y (wind_col_in_3__5), .A0 (nx18371), .A1 (cache_data_out_3__5
          )) ;
    and02 ix5089 (.Y (wind_col_in_3__6), .A0 (nx18371), .A1 (cache_data_out_3__6
          )) ;
    and02 ix5091 (.Y (wind_col_in_3__7), .A0 (nx18371), .A1 (cache_data_out_3__7
          )) ;
    and02 ix5093 (.Y (wind_col_in_3__8), .A0 (nx18373), .A1 (cache_data_out_3__8
          )) ;
    and02 ix5095 (.Y (wind_col_in_3__9), .A0 (nx18373), .A1 (cache_data_out_3__9
          )) ;
    and02 ix5097 (.Y (wind_col_in_3__10), .A0 (nx18373), .A1 (
          cache_data_out_3__10)) ;
    and02 ix5099 (.Y (wind_col_in_3__11), .A0 (nx18373), .A1 (
          cache_data_out_3__11)) ;
    and02 ix5101 (.Y (wind_col_in_3__12), .A0 (nx18373), .A1 (
          cache_data_out_3__12)) ;
    and02 ix5103 (.Y (wind_col_in_3__13), .A0 (nx18373), .A1 (
          cache_data_out_3__13)) ;
    and02 ix5105 (.Y (wind_col_in_3__14), .A0 (nx18373), .A1 (
          cache_data_out_3__14)) ;
    and02 ix5107 (.Y (wind_col_in_3__15), .A0 (nx18375), .A1 (
          cache_data_out_3__15)) ;
    and02 ix5109 (.Y (wind_col_in_4__0), .A0 (nx18375), .A1 (cache_data_out_4__0
          )) ;
    and02 ix5111 (.Y (wind_col_in_4__1), .A0 (nx18375), .A1 (cache_data_out_4__1
          )) ;
    and02 ix5113 (.Y (wind_col_in_4__2), .A0 (nx18375), .A1 (cache_data_out_4__2
          )) ;
    and02 ix5115 (.Y (wind_col_in_4__3), .A0 (nx18375), .A1 (cache_data_out_4__3
          )) ;
    and02 ix5117 (.Y (wind_col_in_4__4), .A0 (nx18375), .A1 (cache_data_out_4__4
          )) ;
    and02 ix5119 (.Y (wind_col_in_4__5), .A0 (nx18375), .A1 (cache_data_out_4__5
          )) ;
    and02 ix5121 (.Y (wind_col_in_4__6), .A0 (nx18157), .A1 (cache_data_out_4__6
          )) ;
    and02 ix5123 (.Y (wind_col_in_4__7), .A0 (nx18157), .A1 (cache_data_out_4__7
          )) ;
    and02 ix5125 (.Y (wind_col_in_4__8), .A0 (nx18157), .A1 (cache_data_out_4__8
          )) ;
    and02 ix5127 (.Y (wind_col_in_4__9), .A0 (nx18157), .A1 (cache_data_out_4__9
          )) ;
    and02 ix5129 (.Y (wind_col_in_4__10), .A0 (nx18157), .A1 (
          cache_data_out_4__10)) ;
    and02 ix5131 (.Y (wind_col_in_4__11), .A0 (nx18157), .A1 (
          cache_data_out_4__11)) ;
    and02 ix5133 (.Y (wind_col_in_4__12), .A0 (nx18157), .A1 (
          cache_data_out_4__12)) ;
    and02 ix5135 (.Y (wind_col_in_4__13), .A0 (nx2546), .A1 (
          cache_data_out_4__13)) ;
    and02 ix5137 (.Y (wind_col_in_4__14), .A0 (nx2546), .A1 (
          cache_data_out_4__14)) ;
    and02 ix5139 (.Y (wind_col_in_4__15), .A0 (nx2546), .A1 (
          cache_data_out_4__15)) ;
    or03 ix2555 (.Y (wind_en), .A0 (nx15974), .A1 (nx18385), .A2 (nx12906)) ;
    or03 ix2547 (.Y (nx2546), .A0 (nx15865), .A1 (nx15970), .A2 (nx18307)) ;
    and03 ix16716 (.Y (nx16715), .A0 (nx18137), .A1 (nx18345), .A2 (nx18313)) ;
    nand02 ix2641 (.Y (nx16927), .A0 (nx18301), .A1 (nx18239)) ;
    nor02ii ix16720 (.Y (nx2142), .A0 (nx18277), .A1 (nx196)) ;
    nor02_2x ix1947 (.Y (nx1946), .A0 (nx1926), .A1 (nx16327)) ;
    nor02ii ix16743 (.Y (nx16742), .A0 (new_size_squared_out_0), .A1 (nx16745)
            ) ;
    or02 ix16748 (.Y (nx16747), .A0 (nx16745), .A1 (nx16324)) ;
    xor2 ix14482 (.Y (nx14481), .A0 (addr1_data_0), .A1 (nx18347)) ;
    or03 ix16752 (.Y (nx18119), .A0 (nx2128), .A1 (nx17927), .A2 (nx2754)) ;
    xor2 ix14472 (.Y (nx14471), .A0 (img_addr_offset_0), .A1 (nx18247)) ;
    mux21_ni ix14462 (.Y (nx14461), .A0 (nx16764), .A1 (img_base_addr_0), .S0 (
             nx18333)) ;
    mux21 ix14452 (.Y (nx14451), .A0 (nx16764), .A1 (nx16745), .S0 (nx18353)) ;
    xor2 ix16771 (.Y (nx16770), .A0 (nflt_layer_temp_1), .A1 (nx15500)) ;
    xor2 ix2675 (.Y (nx2674), .A0 (nflt_layer_temp_0), .A1 (nflt_layer_out_0)) ;
    xor2 ix16775 (.Y (nx16774), .A0 (nflt_layer_temp_2), .A1 (nx15512)) ;
    mux21_ni ix14442 (.Y (nx14441), .A0 (nx15763), .A1 (bias_offset_data_out_0)
             , .S0 (nx18313)) ;
    or02 ix16792 (.Y (nx16791), .A0 (nx16745), .A1 (nx15763)) ;
    xnor2 ix16799 (.Y (nx16798), .A0 (nx16802), .A1 (nx16332)) ;
    ao32 ix14492 (.Y (nx14491), .A0 (write_base_data_out_1), .A1 (nx18265), .A2 (
         nx18335), .B0 (nx19308), .B1 (nx18177)) ;
    inv01 ix18176 (.Y (nx18177), .A (nx16804)) ;
    mux21 ix14522 (.Y (nx14521), .A0 (nx16820), .A1 (nx16818), .S0 (nx18335)) ;
    mux21_ni ix14512 (.Y (nx14511), .A0 (write_base_prev_data_out_1), .A1 (
             write_base_data_out_1), .S0 (nx18353)) ;
    nor02ii ix16826 (.Y (nx16825), .A0 (write_base_prev_data_out_1), .A1 (
            nx16764)) ;
    mux21 ix14532 (.Y (nx14531), .A0 (nx16833), .A1 (nx16829), .S0 (nx18249)) ;
    xnor2 ix16840 (.Y (nx16839), .A0 (nx16843), .A1 (nx16802)) ;
    ao32 ix14542 (.Y (nx14541), .A0 (nx18179), .A1 (nx18301), .A2 (nx18239), .B0 (
         bias_offset_data_out_1), .B1 (nx18313)) ;
    inv01 ix18178 (.Y (nx18179), .A (nx15759)) ;
    mux21 ix14502 (.Y (nx14501), .A0 (nx16846), .A1 (nx16849), .S0 (nx18347)) ;
    xnor2 ix16864 (.Y (nx16863), .A0 (nx16802), .A1 (nx15756)) ;
    xnor2 ix16875 (.Y (nx16874), .A0 (nx18885), .A1 (nx16338)) ;
    ao32 ix14552 (.Y (nx14551), .A0 (write_base_data_out_2), .A1 (nx18265), .A2 (
         nx18335), .B0 (nx19308), .B1 (nx18181)) ;
    inv01 ix18180 (.Y (nx18181), .A (nx16880)) ;
    ao32 ix14602 (.Y (nx14601), .A0 (nx18183), .A1 (nx18301), .A2 (nx18239), .B0 (
         bias_offset_data_out_2), .B1 (nx18313)) ;
    inv01 ix18182 (.Y (nx18183), .A (nx15753)) ;
    mux21_ni ix14582 (.Y (nx14581), .A0 (nx2974), .A1 (img_base_addr_2), .S0 (
             nx18335)) ;
    mux21 ix14572 (.Y (nx14571), .A0 (nx16906), .A1 (nx18885), .S0 (nx18353)) ;
    mux21_ni ix14592 (.Y (nx14591), .A0 (img_addr_offset_2), .A1 (nx2988), .S0 (
             nx18249)) ;
    xor2 ix2989 (.Y (nx2988), .A0 (nx16915), .A1 (nx16831)) ;
    mux21_ni ix14562 (.Y (nx14561), .A0 (addr1_data_2), .A1 (nx2942), .S0 (
             nx18347)) ;
    xnor2 ix16925 (.Y (nx16924), .A0 (nx18885), .A1 (nx15750)) ;
    oai21 ix2933 (.Y (nx2932), .A0 (nx18185), .A1 (nx18345), .B0 (nx18311)) ;
    inv01 ix18184 (.Y (nx18185), .A (nx2874)) ;
    mux21_ni ix14612 (.Y (nx14611), .A0 (write_base_data_out_3), .A1 (nx3050), .S0 (
             nx19308)) ;
    xor2 ix16944 (.Y (nx16943), .A0 (new_size_squared_out_3), .A1 (nx18889)) ;
    mux21_ni ix14652 (.Y (nx14651), .A0 (nx3146), .A1 (img_base_addr_3), .S0 (
             nx18335)) ;
    mux21_ni ix14642 (.Y (nx14641), .A0 (write_base_prev_data_out_3), .A1 (
             write_base_data_out_3), .S0 (nx18353)) ;
    mux21_ni ix14662 (.Y (nx14661), .A0 (img_addr_offset_3), .A1 (nx3160), .S0 (
             nx18249)) ;
    xor2 ix16968 (.Y (nx16967), .A0 (bias_offset_data_out_3), .A1 (nx18889)) ;
    mux21_ni ix14632 (.Y (nx14631), .A0 (nx832), .A1 (bias_offset_data_out_3), .S0 (
             nx18313)) ;
    xor2 ix833 (.Y (nx832), .A0 (nx15745), .A1 (nx15768)) ;
    mux21_ni ix14622 (.Y (nx14621), .A0 (addr1_data_3), .A1 (nx3092), .S0 (
             nx18347)) ;
    ao32 ix14672 (.Y (nx14671), .A0 (write_base_data_out_4), .A1 (nx18267), .A2 (
         nx18335), .B0 (nx19308), .B1 (nx18187)) ;
    inv01 ix18186 (.Y (nx18187), .A (nx17004)) ;
    mux21_ni ix14722 (.Y (nx14721), .A0 (nx858), .A1 (bias_offset_data_out_4), .S0 (
             nx18313)) ;
    mux21_ni ix14702 (.Y (nx14701), .A0 (nx3270), .A1 (img_base_addr_4), .S0 (
             nx18335)) ;
    mux21 ix14692 (.Y (nx14691), .A0 (nx17031), .A1 (nx18891), .S0 (nx18353)) ;
    mux21_ni ix14712 (.Y (nx14711), .A0 (img_addr_offset_4), .A1 (nx3284), .S0 (
             nx18249)) ;
    nor02ii ix3279 (.Y (nx3278), .A0 (nx17042), .A1 (img_addr_offset_4)) ;
    xnor2 ix17052 (.Y (nx17051), .A0 (nx18891), .A1 (nx15735)) ;
    mux21_ni ix14682 (.Y (nx14681), .A0 (addr1_data_4), .A1 (nx3238), .S0 (
             nx18347)) ;
    nor02ii ix3233 (.Y (nx3232), .A0 (nx17060), .A1 (addr1_data_4)) ;
    mux21_ni ix14732 (.Y (nx14731), .A0 (write_base_data_out_5), .A1 (nx3346), .S0 (
             nx19308)) ;
    xor2 ix17075 (.Y (nx17074), .A0 (new_size_squared_out_5), .A1 (nx17076)) ;
    xnor2 ix17082 (.Y (nx17081), .A0 (nx17085), .A1 (nx17076)) ;
    ao32 ix14782 (.Y (nx14781), .A0 (nx18189), .A1 (nx18303), .A2 (nx18239), .B0 (
         bias_offset_data_out_5), .B1 (nx18315)) ;
    inv01 ix18188 (.Y (nx18189), .A (nx15732)) ;
    xor2 ix17090 (.Y (nx17089), .A0 (img_base_addr_5), .A1 (nx17104)) ;
    mux21_ni ix14762 (.Y (nx14761), .A0 (nx3412), .A1 (img_base_addr_5), .S0 (
             nx18041)) ;
    mux21_ni ix14752 (.Y (nx14751), .A0 (write_base_prev_data_out_5), .A1 (
             write_base_data_out_5), .S0 (nx18353)) ;
    mux21 ix14772 (.Y (nx14771), .A0 (nx17104), .A1 (nx17100), .S0 (nx18249)) ;
    mux21 ix14742 (.Y (nx14741), .A0 (nx17114), .A1 (nx17110), .S0 (nx18347)) ;
    mux21_ni ix14842 (.Y (nx14841), .A0 (nx904), .A1 (bias_offset_data_out_6), .S0 (
             nx18315)) ;
    ao32 ix14792 (.Y (nx14791), .A0 (write_base_data_out_6), .A1 (nx18267), .A2 (
         nx18041), .B0 (nx19308), .B1 (nx18191)) ;
    inv01 ix18190 (.Y (nx18191), .A (nx17140)) ;
    mux21_ni ix14822 (.Y (nx14821), .A0 (nx3554), .A1 (img_base_addr_6), .S0 (
             nx18041)) ;
    mux21 ix14812 (.Y (nx14811), .A0 (nx17157), .A1 (nx18893), .S0 (nx18353)) ;
    mux21_ni ix14832 (.Y (nx14831), .A0 (img_addr_offset_6), .A1 (nx3568), .S0 (
             nx18249)) ;
    nor02ii ix3563 (.Y (nx3562), .A0 (nx17102), .A1 (img_addr_offset_6)) ;
    nor02ii ix3361 (.Y (nx3360), .A0 (nx17077), .A1 (write_base_data_out_5)) ;
    xnor2 ix17187 (.Y (nx17186), .A0 (nx18893), .A1 (nx15720)) ;
    mux21_ni ix14802 (.Y (nx14801), .A0 (addr1_data_6), .A1 (nx3522), .S0 (
             nx18347)) ;
    xor2 ix3523 (.Y (nx3522), .A0 (nx17188), .A1 (nx17112)) ;
    mux21_ni ix14852 (.Y (nx14851), .A0 (nx18895), .A1 (nx3630), .S0 (nx19294)
             ) ;
    xor2_2x ix17205 (.Y (nx17204), .A0 (new_size_squared_out_7), .A1 (nx17199)
            ) ;
    xnor2 ix17211 (.Y (nx17210), .A0 (nx17214), .A1 (nx17199)) ;
    ao32 ix14902 (.Y (nx14901), .A0 (nx18193), .A1 (nx18303), .A2 (nx18239), .B0 (
         bias_offset_data_out_7), .B1 (nx18315)) ;
    inv01 ix18192 (.Y (nx18193), .A (nx15717)) ;
    xor2 ix17219 (.Y (nx17218), .A0 (img_base_addr_7), .A1 (nx17233)) ;
    mux21_ni ix14882 (.Y (nx14881), .A0 (nx3696), .A1 (img_base_addr_7), .S0 (
             nx18041)) ;
    mux21_ni ix14872 (.Y (nx14871), .A0 (write_base_prev_data_out_7), .A1 (
             nx18895), .S0 (nx18355)) ;
    mux21 ix14892 (.Y (nx14891), .A0 (nx17233), .A1 (nx17229), .S0 (nx18249)) ;
    mux21 ix14862 (.Y (nx14861), .A0 (nx17244), .A1 (nx17239), .S0 (nx18349)) ;
    nor02ii ix3517 (.Y (nx3516), .A0 (nx17112), .A1 (addr1_data_6)) ;
    oai21 ix3655 (.Y (nx3654), .A0 (nx18195), .A1 (nx18345), .B0 (nx18311)) ;
    inv01 ix18194 (.Y (nx18195), .A (nx3600)) ;
    mux21_ni ix14962 (.Y (nx14961), .A0 (nx954), .A1 (bias_offset_data_out_8), .S0 (
             nx18315)) ;
    ao32 ix14912 (.Y (nx14911), .A0 (nx18897), .A1 (nx18267), .A2 (nx18337), .B0 (
         nx19294), .B1 (nx18197)) ;
    inv01 ix18196 (.Y (nx18197), .A (nx17270)) ;
    mux21_ni ix14942 (.Y (nx14941), .A0 (nx3838), .A1 (img_base_addr_8), .S0 (
             nx18337)) ;
    mux21 ix14932 (.Y (nx14931), .A0 (nx17287), .A1 (nx18899), .S0 (nx18355)) ;
    mux21_ni ix14952 (.Y (nx14951), .A0 (img_addr_offset_8), .A1 (nx3852), .S0 (
             nx18251)) ;
    nor02ii ix3847 (.Y (nx3846), .A0 (nx17231), .A1 (img_addr_offset_8)) ;
    xnor2 ix17311 (.Y (nx17310), .A0 (nx18899), .A1 (nx15686)) ;
    mux21_ni ix14922 (.Y (nx14921), .A0 (addr1_data_8), .A1 (nx3806), .S0 (
             nx18349)) ;
    xor2 ix3807 (.Y (nx3806), .A0 (nx17315), .A1 (nx17242)) ;
    mux21_ni ix14972 (.Y (nx14971), .A0 (nx18901), .A1 (nx3914), .S0 (nx19294)
             ) ;
    xor2 ix17332 (.Y (nx17331), .A0 (new_size_squared_out_9), .A1 (nx17326)) ;
    xnor2 ix17338 (.Y (nx17337), .A0 (nx17341), .A1 (nx17326)) ;
    ao32 ix15022 (.Y (nx15021), .A0 (nx18199), .A1 (nx18303), .A2 (nx18239), .B0 (
         bias_offset_data_out_9), .B1 (nx18315)) ;
    inv01 ix18198 (.Y (nx18199), .A (nx15683)) ;
    xor2 ix17346 (.Y (nx17345), .A0 (img_base_addr_9), .A1 (nx17360)) ;
    mux21_ni ix15002 (.Y (nx15001), .A0 (nx3980), .A1 (img_base_addr_9), .S0 (
             nx18337)) ;
    mux21_ni ix14992 (.Y (nx14991), .A0 (write_base_prev_data_out_9), .A1 (
             nx18901), .S0 (nx18355)) ;
    mux21 ix15012 (.Y (nx15011), .A0 (nx17360), .A1 (nx17356), .S0 (nx18251)) ;
    mux21 ix14982 (.Y (nx14981), .A0 (nx17371), .A1 (nx17366), .S0 (nx18349)) ;
    nor02ii ix3801 (.Y (nx3800), .A0 (nx17242), .A1 (addr1_data_8)) ;
    xnor2 ix17378 (.Y (nx17377), .A0 (nx17326), .A1 (nx15770)) ;
    oai21 ix3939 (.Y (nx3938), .A0 (nx18201), .A1 (nx18345), .B0 (nx18311)) ;
    inv01 ix18200 (.Y (nx18201), .A (nx3884)) ;
    mux21_ni ix15082 (.Y (nx15081), .A0 (nx1000), .A1 (bias_offset_data_out_10)
             , .S0 (nx18315)) ;
    ao32 ix15032 (.Y (nx15031), .A0 (write_base_data_out_10), .A1 (nx18267), .A2 (
         nx18337), .B0 (nx19294), .B1 (nx18203)) ;
    inv01 ix18202 (.Y (nx18203), .A (nx17397)) ;
    mux21_ni ix15062 (.Y (nx15061), .A0 (nx4122), .A1 (img_base_addr_10), .S0 (
             nx18337)) ;
    mux21 ix15052 (.Y (nx15051), .A0 (nx17414), .A1 (nx18903), .S0 (nx18355)) ;
    mux21_ni ix15072 (.Y (nx15071), .A0 (img_addr_offset_10), .A1 (nx4136), .S0 (
             nx18251)) ;
    nor02ii ix4131 (.Y (nx4130), .A0 (nx17358), .A1 (img_addr_offset_10)) ;
    xnor2 ix17438 (.Y (nx17437), .A0 (nx18903), .A1 (nx15673)) ;
    mux21_ni ix15042 (.Y (nx15041), .A0 (addr1_data_10), .A1 (nx4090), .S0 (
             nx18349)) ;
    xor2 ix4091 (.Y (nx4090), .A0 (nx17442), .A1 (nx17369)) ;
    mux21_ni ix15092 (.Y (nx15091), .A0 (nx18905), .A1 (nx4198), .S0 (nx19294)
             ) ;
    xor2 ix17459 (.Y (nx17458), .A0 (new_size_squared_out_11), .A1 (nx18907)) ;
    xnor2 ix17465 (.Y (nx17464), .A0 (nx17468), .A1 (nx18907)) ;
    ao32 ix15142 (.Y (nx15141), .A0 (nx18205), .A1 (nx18303), .A2 (nx18239), .B0 (
         bias_offset_data_out_11), .B1 (nx18315)) ;
    inv01 ix18204 (.Y (nx18205), .A (nx15670)) ;
    xor2 ix17473 (.Y (nx17472), .A0 (img_base_addr_11), .A1 (nx17487)) ;
    mux21_ni ix15122 (.Y (nx15121), .A0 (nx4264), .A1 (img_base_addr_11), .S0 (
             nx18337)) ;
    mux21_ni ix15112 (.Y (nx15111), .A0 (write_base_prev_data_out_11), .A1 (
             nx18905), .S0 (nx18355)) ;
    mux21 ix15132 (.Y (nx15131), .A0 (nx17487), .A1 (nx17483), .S0 (nx18251)) ;
    mux21 ix15102 (.Y (nx15101), .A0 (nx17498), .A1 (nx17493), .S0 (nx18349)) ;
    nor02ii ix4085 (.Y (nx4084), .A0 (nx17369), .A1 (addr1_data_10)) ;
    oai21 ix4223 (.Y (nx4222), .A0 (nx18207), .A1 (nx18077), .B0 (nx18311)) ;
    inv01 ix18206 (.Y (nx18207), .A (nx4168)) ;
    mux21_ni ix15202 (.Y (nx15201), .A0 (nx1048), .A1 (bias_offset_data_out_12)
             , .S0 (nx18317)) ;
    mux21_ni ix15182 (.Y (nx15181), .A0 (nx4406), .A1 (img_base_addr_12), .S0 (
             nx18043)) ;
    mux21 ix15172 (.Y (nx15171), .A0 (nx17541), .A1 (nx18909), .S0 (nx18355)) ;
    mux21_ni ix15192 (.Y (nx15191), .A0 (img_addr_offset_12), .A1 (nx4420), .S0 (
             nx18251)) ;
    nor02ii ix4415 (.Y (nx4414), .A0 (nx17485), .A1 (img_addr_offset_12)) ;
    xnor2 ix17565 (.Y (nx17564), .A0 (nx18909), .A1 (nx15660)) ;
    mux21_ni ix15162 (.Y (nx15161), .A0 (addr1_data_12), .A1 (nx4374), .S0 (
             nx18349)) ;
    xor2 ix4375 (.Y (nx4374), .A0 (nx17566), .A1 (nx17496)) ;
    xnor2 ix17592 (.Y (nx17591), .A0 (nx17595), .A1 (nx18913)) ;
    ao32 ix15262 (.Y (nx15261), .A0 (nx18211), .A1 (nx18303), .A2 (nx18241), .B0 (
         bias_offset_data_out_13), .B1 (nx18317)) ;
    inv01 ix18210 (.Y (nx18211), .A (nx15657)) ;
    xor2 ix17600 (.Y (nx17599), .A0 (img_base_addr_13), .A1 (nx17614)) ;
    mux21_ni ix15242 (.Y (nx15241), .A0 (nx4548), .A1 (img_base_addr_13), .S0 (
             nx18043)) ;
    mux21_ni ix15232 (.Y (nx15231), .A0 (write_base_prev_data_out_13), .A1 (
             write_base_data_out_13), .S0 (nx18355)) ;
    mux21 ix15252 (.Y (nx15251), .A0 (nx17614), .A1 (nx17610), .S0 (nx18251)) ;
    mux21 ix15222 (.Y (nx15221), .A0 (nx17625), .A1 (nx17620), .S0 (nx18349)) ;
    nor02ii ix4369 (.Y (nx4368), .A0 (nx17496), .A1 (addr1_data_12)) ;
    oai21 ix4507 (.Y (nx4506), .A0 (nx18213), .A1 (nx18077), .B0 (nx18311)) ;
    xnor2 ix17642 (.Y (nx17641), .A0 (nx17646), .A1 (nx18915)) ;
    mux21_ni ix15322 (.Y (nx15321), .A0 (nx1094), .A1 (bias_offset_data_out_14)
             , .S0 (nx18317)) ;
    xor2 ix1095 (.Y (nx1094), .A0 (nx15647), .A1 (nx15653)) ;
    xnor2 ix17664 (.Y (nx17663), .A0 (nx17673), .A1 (nx17677)) ;
    mux21_ni ix15302 (.Y (nx15301), .A0 (nx4690), .A1 (img_base_addr_14), .S0 (
             nx18043)) ;
    xnor2 ix4691 (.Y (nx4690), .A0 (nx17670), .A1 (nx17671)) ;
    mux21 ix15292 (.Y (nx15291), .A0 (nx17670), .A1 (nx18915), .S0 (nx18357)) ;
    mux21_ni ix15312 (.Y (nx15311), .A0 (img_addr_offset_14), .A1 (nx4704), .S0 (
             nx18251)) ;
    xor2 ix4705 (.Y (nx4704), .A0 (nx17677), .A1 (nx17612)) ;
    xor2 ix17680 (.Y (nx17679), .A0 (nx18915), .A1 (nx4496)) ;
    xnor2 ix17686 (.Y (nx17685), .A0 (nx18916), .A1 (nx15647)) ;
    mux21_ni ix15282 (.Y (nx15281), .A0 (addr1_data_14), .A1 (nx4658), .S0 (
             nx18351)) ;
    xor2 ix4659 (.Y (nx4658), .A0 (nx17687), .A1 (nx17623)) ;
    xor2 ix17712 (.Y (nx17711), .A0 (img_base_addr_15), .A1 (nx17726)) ;
    mux21_ni ix15372 (.Y (nx15371), .A0 (nx4834), .A1 (img_base_addr_15), .S0 (
             nx18043)) ;
    mux21_ni ix15362 (.Y (nx15361), .A0 (write_base_prev_data_out_15), .A1 (
             write_base_data_out_15), .S0 (nx18357)) ;
    mux21 ix15382 (.Y (nx15381), .A0 (nx17726), .A1 (nx17723), .S0 (nx18253)) ;
    xor2 ix17724 (.Y (nx17723), .A0 (nx17726), .A1 (nx4698)) ;
    nor02ii ix4699 (.Y (nx4698), .A0 (nx17612), .A1 (img_addr_offset_14)) ;
    xor2 ix4803 (.Y (nx4802), .A0 (write_base_data_out_15), .A1 (
         write_offset_data_out_15)) ;
    mux21 ix15352 (.Y (nx15351), .A0 (nx17740), .A1 (nx17737), .S0 (nx18351)) ;
    xor2 ix17738 (.Y (nx17737), .A0 (nx17740), .A1 (nx4652)) ;
    nor02ii ix4653 (.Y (nx4652), .A0 (nx17623), .A1 (addr1_data_14)) ;
    xor2 ix17745 (.Y (nx17744), .A0 (nx17748), .A1 (write_base_data_out_15)) ;
    ao32 ix15332 (.Y (nx15331), .A0 (nx18217), .A1 (nx18303), .A2 (nx18241), .B0 (
         bias_offset_data_out_15), .B1 (nx18317)) ;
    inv01 ix18216 (.Y (nx18217), .A (nx15644)) ;
    inv02 ix18218 (.Y (nx18219), .A (nx16222)) ;
    inv02 ix18224 (.Y (nx18225), .A (nx15974)) ;
    inv02 ix18226 (.Y (nx18227), .A (nx15974)) ;
    inv01 ix18228 (.Y (nx18229), .A (nx18049)) ;
    inv01 ix18230 (.Y (nx18231), .A (nx18049)) ;
    inv01 ix18232 (.Y (nx18233), .A (nx18059)) ;
    inv01 ix18234 (.Y (nx18235), .A (nx18059)) ;
    inv01 ix18236 (.Y (nx18237), .A (nx18059)) ;
    inv02 ix18238 (.Y (nx18239), .A (nx18117)) ;
    inv02 ix18240 (.Y (nx18241), .A (nx18117)) ;
    inv02 ix18242 (.Y (nx18243), .A (nx18081)) ;
    inv02 ix18244 (.Y (nx18245), .A (nx18081)) ;
    inv02 ix18246 (.Y (nx18247), .A (nx18081)) ;
    inv02 ix18248 (.Y (nx18249), .A (nx18081)) ;
    inv02 ix18250 (.Y (nx18251), .A (nx18081)) ;
    inv02 ix18252 (.Y (nx18253), .A (nx18081)) ;
    inv02 ix18254 (.Y (nx18255), .A (nx17927)) ;
    inv02 ix18256 (.Y (nx18257), .A (nx17927)) ;
    inv02 ix18258 (.Y (nx18259), .A (nx582)) ;
    inv02 ix18260 (.Y (nx18261), .A (nx582)) ;
    buf02 ix18262 (.Y (nx18263), .A (nx15496)) ;
    inv02 ix18264 (.Y (nx18265), .A (nx17887)) ;
    inv01 ix18268 (.Y (nx18269), .A (nx148)) ;
    inv01 ix18270 (.Y (nx18271), .A (nx148)) ;
    inv02 ix18272 (.Y (nx18273), .A (nx17971)) ;
    inv02 ix18274 (.Y (nx18275), .A (nx17971)) ;
    inv02 ix18276 (.Y (nx18277), .A (nx17971)) ;
    inv02 ix18278 (.Y (nx18279), .A (nx17921)) ;
    inv02 ix18280 (.Y (nx18281), .A (nx17921)) ;
    inv02 ix18282 (.Y (nx18283), .A (nx12884)) ;
    inv02 ix18284 (.Y (nx18285), .A (nx12884)) ;
    inv02 ix18286 (.Y (nx18287), .A (nx12884)) ;
    inv02 ix18288 (.Y (nx18289), .A (nx1212)) ;
    inv02 ix18290 (.Y (nx18291), .A (nx18383)) ;
    inv02 ix18292 (.Y (nx18293), .A (nx18383)) ;
    inv01 ix18294 (.Y (nx18295), .A (nx16373)) ;
    inv02 ix18296 (.Y (nx18297), .A (nx18295)) ;
    inv02 ix18298 (.Y (nx18299), .A (nx18295)) ;
    inv02 ix18300 (.Y (nx18301), .A (nx18295)) ;
    inv02 ix18302 (.Y (nx18303), .A (nx18295)) ;
    inv02 ix18304 (.Y (nx18305), .A (comp_unit_flt_size)) ;
    inv02 ix18306 (.Y (nx18307), .A (comp_unit_flt_size)) ;
    inv02 ix18308 (.Y (nx18309), .A (nx17975)) ;
    inv02 ix18310 (.Y (nx18311), .A (nx17975)) ;
    inv02 ix18312 (.Y (nx18313), .A (nx18011)) ;
    inv02 ix18314 (.Y (nx18315), .A (nx18011)) ;
    inv02 ix18316 (.Y (nx18317), .A (nx18011)) ;
    inv01 ix18318 (.Y (nx18319), .A (filter_ready_out)) ;
    inv01 ix18320 (.Y (nx18321), .A (filter_ready_out)) ;
    inv02 ix18322 (.Y (nx18323), .A (current_state_7)) ;
    inv02 ix18324 (.Y (nx18325), .A (current_state_7)) ;
    inv02 ix18326 (.Y (nx18327), .A (current_state_7)) ;
    inv02 ix18328 (.Y (nx18329), .A (nx17947)) ;
    inv02 ix18330 (.Y (nx18331), .A (nx17947)) ;
    inv02 ix18332 (.Y (nx18333), .A (nx18912)) ;
    inv02 ix18334 (.Y (nx18335), .A (nx18912)) ;
    inv02 ix18338 (.Y (nx18339), .A (nx18381)) ;
    inv02 ix18340 (.Y (nx18341), .A (nx18381)) ;
    inv02 ix18342 (.Y (nx18343), .A (nx18381)) ;
    inv02 ix18344 (.Y (nx18345), .A (nx18381)) ;
    inv02 ix18346 (.Y (nx18347), .A (nx18121)) ;
    inv02 ix18348 (.Y (nx18349), .A (nx18121)) ;
    inv02 ix18350 (.Y (nx18351), .A (nx18121)) ;
    inv02 ix18352 (.Y (nx18353), .A (nx16768)) ;
    inv02 ix18354 (.Y (nx18355), .A (nx16768)) ;
    inv02 ix18356 (.Y (nx18357), .A (nx16768)) ;
    inv01 ix18358 (.Y (nx18359), .A (nx18385)) ;
    inv01 ix18360 (.Y (nx18361), .A (nx18385)) ;
    inv01 ix18362 (.Y (nx18363), .A (nx18385)) ;
    inv01 ix18364 (.Y (nx18365), .A (nx18385)) ;
    inv01 ix18366 (.Y (nx18367), .A (nx16629)) ;
    inv01 ix18368 (.Y (nx18369), .A (nx16629)) ;
    inv01 ix18370 (.Y (nx18371), .A (nx16629)) ;
    inv01 ix18372 (.Y (nx18373), .A (nx16629)) ;
    inv01 ix18374 (.Y (nx18375), .A (nx16629)) ;
    inv02 ix18380 (.Y (nx18381), .A (nx18075)) ;
    inv01 ix18382 (.Y (nx18383), .A (nx18289)) ;
    inv01 ix18384 (.Y (nx18385), .A (nx2546)) ;
    nor02ii ix17068 (.Y (nx17067), .A0 (nx3366), .A1 (nx16995)) ;
    xor2 ix3367 (.Y (nx3366), .A0 (nx17076), .A1 (nx17077)) ;
    nor02ii ix16996 (.Y (nx16995), .A0 (nx3078), .A1 (nx18867)) ;
    buf04 ix18917 (.Y (nx18543), .A (nx17067)) ;
    inv02 ix18918 (.Y (nx18544), .A (new_size_squared_out_15)) ;
    inv02 ix18919 (.Y (nx18545), .A (write_base_data_out_15)) ;
    oai32 ix18920 (.Y (nx18546), .A0 (nx19302), .A1 (nx18544), .A2 (
          write_base_data_out_15), .B0 (nx18545), .B1 (new_size_squared_out_15)
          ) ;
    and02 ix18921 (.Y (nx18547), .A0 (nx18909), .A1 (nx15795)) ;
    nor02_2x ix18922 (.Y (nx18548), .A0 (nx18909), .A1 (nx15795)) ;
    and02 ix18923 (.Y (nx18549), .A0 (nx18916), .A1 (nx15785)) ;
    inv02 ix18924 (.Y (nx18550), .A (write_base_data_out_13)) ;
    inv02 ix18925 (.Y (nx18551), .A (new_size_squared_out_13)) ;
    aoi32 ix18926 (.Y (nx18552), .A0 (nx18223), .A1 (nx18545), .A2 (nx18544), .B0 (
          write_base_data_out_15), .B1 (new_size_squared_out_15)) ;
    nor02_2x ix18927 (.Y (nx18553), .A0 (NOT_nx4768), .A1 (nx18552)) ;
    ao221 reg_nx15341 (.Y (nx15341), .A0 (nx18546), .A1 (NOT_nx4768), .B0 (
          write_base_data_out_15), .B1 (nx19302), .C0 (nx18553)) ;
    and02 ix18928 (.Y (nx18554), .A0 (write_base_data_out_13), .A1 (
          new_size_squared_out_13)) ;
    inv02 ix18929 (.Y (nx18555), .A (nx17585)) ;
    inv01 ix18930 (.Y (nx18556), .A (nx18916)) ;
    inv02 ix18931 (.Y (nx18557), .A (nx15785)) ;
    inv02 ix18932 (.Y (nx18558), .A (nx18909)) ;
    inv02 ix18933 (.Y (nx18559), .A (nx15795)) ;
    inv01 ix18934 (.Y (nx18560), .A (nx18885)) ;
    inv02 ix18935 (.Y (nx18561), .A (nx15848)) ;
    nand02_2x ix18936 (.Y (nx18562), .A0 (nx18886), .A1 (nx15848)) ;
    inv02 reg_nx18009 (.Y (nx18009), .A (nx16745)) ;
    inv02 ix18937 (.Y (nx18563), .A (nx16802)) ;
    nand03_2x ix18938 (.Y (nx18564), .A0 (new_size_squared_out_0), .A1 (nx18009)
              , .A2 (nx18563)) ;
    inv02 ix18939 (.Y (nx18565), .A (new_size_squared_out_1)) ;
    nand02_2x ix18940 (.Y (nx18566), .A0 (new_size_squared_out_1), .A1 (nx18563)
              ) ;
    nand03_2x ix18941 (.Y (nx18567), .A0 (nx18566), .A1 (new_size_squared_out_0)
              , .A2 (nx18009)) ;
    inv02 ix18942 (.Y (nx18568), .A (write_base_data_out_1)) ;
    inv01 reg_nx3046 (.Y (nx3046), .A (nx18877)) ;
    inv01 reg_nx16882 (.Y (nx16882), .A (nx18774)) ;
    oai22 reg_nx16885 (.Y (nx16885), .A0 (nx18560), .A1 (nx18561), .B0 (nx18886)
          , .B1 (nx15848)) ;
    oai22 reg_nx16808 (.Y (nx16808), .A0 (nx18563), .A1 (new_size_squared_out_1)
          , .B0 (nx18565), .B1 (nx16802)) ;
    nor02_2x ix18943 (.Y (nx18569), .A0 (nx18549), .A1 (nx17585)) ;
    nor02_2x ix18944 (.Y (nx18570), .A0 (nx18547), .A1 (nx17458)) ;
    inv02 ix18945 (.Y (nx18571), .A (nx18905)) ;
    inv02 ix18946 (.Y (nx18572), .A (new_size_squared_out_11)) ;
    nor03_2x ix18947 (.Y (nx18573), .A0 (nx18547), .A1 (nx18571), .A2 (nx18572)
             ) ;
    or02 ix18948 (.Y (nx18574), .A0 (nx18573), .A1 (nx18548)) ;
    oai32 ix18949 (.Y (nx18575), .A0 (nx18549), .A1 (nx18550), .A2 (nx18551), .B0 (
          nx18916), .B1 (nx15785)) ;
    aoi321 reg_NOT_nx4768 (.Y (NOT_nx4768), .A0 (nx18689), .A1 (nx18569), .A2 (
           nx18570), .B0 (nx18574), .B1 (nx18569), .C0 (nx18575)) ;
    inv01 ix18950 (.Y (nx18576), .A (nx18547)) ;
    and02 ix18951 (.Y (nx18577), .A0 (nx18905), .A1 (new_size_squared_out_11)) ;
    inv02 ix18952 (.Y (nx18578), .A (nx17458)) ;
    inv02 ix18953 (.Y (nx18579), .A (nx16839)) ;
    aoi32 reg_nx16888 (.Y (nx16888), .A0 (nx18579), .A1 (bias_offset_data_out_0)
          , .A2 (nx18009), .B0 (write_base_data_out_1), .B1 (
          bias_offset_data_out_1)) ;
    and02 ix18954 (.Y (nx18580), .A0 (nx18886), .A1 (nx16895)) ;
    nor02_2x ix18955 (.Y (nx18581), .A0 (nx16888), .A1 (nx18580)) ;
    nor02_2x ix18956 (.Y (nx18582), .A0 (nx18886), .A1 (nx16895)) ;
    and02 ix18957 (.Y (nx18583), .A0 (nx18891), .A1 (nx17021)) ;
    inv02 ix18958 (.Y (nx18584), .A (write_base_data_out_3)) ;
    inv02 ix18959 (.Y (nx18585), .A (bias_offset_data_out_3)) ;
    inv01 reg_nx3444 (.Y (nx3444), .A (nx18657)) ;
    and02 ix18960 (.Y (nx18586), .A0 (write_base_data_out_3), .A1 (
          bias_offset_data_out_3)) ;
    inv02 ix18961 (.Y (nx18587), .A (nx16967)) ;
    oai32 reg_nx17013 (.Y (nx17013), .A0 (nx18586), .A1 (nx18581), .A2 (nx18582)
          , .B0 (nx18587), .B1 (nx18586)) ;
    nor02_2x ix18962 (.Y (nx18588), .A0 (nx18891), .A1 (nx17021)) ;
    ao21 reg_nx17016 (.Y (nx17016), .A0 (nx18891), .A1 (nx17021), .B0 (nx18588)
         ) ;
    inv02 reg_nx3112 (.Y (nx3112), .A (nx18660)) ;
    ao21 reg_nx16891 (.Y (nx16891), .A0 (nx18886), .A1 (nx16895), .B0 (nx18582)
         ) ;
    nand02_2x ix18963 (.Y (nx18589), .A0 (write_offset_data_out_6), .A1 (
              write_base_data_out_6)) ;
    inv02 ix18964 (.Y (nx18590), .A (nx16924)) ;
    aoi22 reg_nx16987 (.Y (nx16987), .A0 (write_offset_data_out_2), .A1 (
          write_base_data_out_2), .B0 (nx2892), .B1 (nx18590)) ;
    and02 ix18965 (.Y (nx18591), .A0 (nx15745), .A1 (nx18889)) ;
    nor02_2x ix18966 (.Y (nx18592), .A0 (nx16987), .A1 (nx18591)) ;
    nor02_2x ix18967 (.Y (nx18593), .A0 (nx15745), .A1 (nx18889)) ;
    and02 ix18968 (.Y (nx18594), .A0 (nx15730), .A1 (nx17076)) ;
    inv02 ix18969 (.Y (nx18595), .A (write_offset_data_out_4)) ;
    inv02 ix18970 (.Y (nx18596), .A (write_base_data_out_4)) ;
    inv01 ix18971 (.Y (nx18597), .A (NOT_nx3476)) ;
    and02 ix18972 (.Y (nx18598), .A0 (write_offset_data_out_4), .A1 (
          write_base_data_out_4)) ;
    inv02 ix18973 (.Y (nx18599), .A (nx17051)) ;
    oai32 reg_nx17118 (.Y (nx17118), .A0 (nx18598), .A1 (nx18592), .A2 (nx18593)
          , .B0 (nx18599), .B1 (nx18598)) ;
    inv02 ix18974 (.Y (nx18600), .A (nx15730)) ;
    inv02 ix18975 (.Y (nx18601), .A (nx17076)) ;
    oai22 reg_nx17121 (.Y (nx17121), .A0 (nx18600), .A1 (nx18601), .B0 (nx15730)
          , .B1 (nx17076)) ;
    inv01 reg_nx3184 (.Y (nx3184), .A (nx18743)) ;
    inv02 ix18976 (.Y (nx18602), .A (nx15745)) ;
    inv02 ix18977 (.Y (nx18603), .A (nx18889)) ;
    oai22 reg_nx16990 (.Y (nx16990), .A0 (nx18602), .A1 (nx18603), .B0 (nx15745)
          , .B1 (nx18890)) ;
    aoi22 ix18978 (.Y (nx18604), .A0 (nx18576), .A1 (nx18577), .B0 (nx18690), .B1 (
          nx18570)) ;
    oai22 reg_nx17656 (.Y (nx17656), .A0 (nx18556), .A1 (nx18557), .B0 (nx18916)
          , .B1 (nx15785)) ;
    inv02 ix18979 (.Y (nx18605), .A (nx17656)) ;
    inv01 reg_nx18223 (.Y (nx18223), .A (nx19302)) ;
    nand02_2x ix18980 (.Y (nx18606), .A0 (nx18223), .A1 (nx18555)) ;
    inv01 ix18981 (.Y (nx18607), .A (nx18604)) ;
    inv02 ix18982 (.Y (nx18608), .A (nx18554)) ;
    inv02 ix18983 (.Y (nx18609), .A (nx18548)) ;
    nand04_2x ix18984 (.Y (nx18610), .A0 (nx18605), .A1 (nx18223), .A2 (nx18608)
              , .A3 (nx18609)) ;
    inv02 reg_nx18043 (.Y (nx18043), .A (nx18912)) ;
    aoi21 ix18985 (.Y (nx18611), .A0 (nx18548), .A1 (nx18555), .B0 (nx18554)) ;
    inv02 ix18986 (.Y (nx18612), .A (nx18555)) ;
    nand03_2x ix18987 (.Y (nx18613), .A0 (nx18605), .A1 (nx18608), .A2 (nx18612)
              ) ;
    oai21 ix18988 (.Y (nx18614), .A0 (nx18605), .A1 (nx18611), .B0 (nx18613)) ;
    aoi32 ix18989 (.Y (nx18615), .A0 (write_base_data_out_14), .A1 (nx18267), .A2 (
          nx18043), .B0 (nx18223), .B1 (nx18614)) ;
    oai321 reg_nx15271 (.Y (nx15271), .A0 (nx18604), .A1 (nx18605), .A2 (nx18606
           ), .B0 (nx18607), .B1 (nx18610), .C0 (nx18615)) ;
    nand02_2x ix18990 (.Y (nx18616), .A0 (write_offset_data_out_14), .A1 (
              write_base_data_out_14)) ;
    inv02 ix18991 (.Y (nx18617), .A (nx15772)) ;
    inv02 ix18992 (.Y (nx18618), .A (nx18907)) ;
    nand02_2x ix18993 (.Y (nx18619), .A0 (nx15772), .A1 (nx18907)) ;
    and02 ix18994 (.Y (nx18620), .A0 (write_offset_data_out_10), .A1 (
          write_base_data_out_10)) ;
    aoi21 ix18995 (.Y (nx18621), .A0 (nx15772), .A1 (nx18908), .B0 (nx17437)) ;
    aoi222 ix18996 (.Y (nx18622), .A0 (nx18617), .A1 (nx18618), .B0 (nx18619), .B1 (
           nx18620), .C0 (nx4044), .C1 (nx18621)) ;
    and02 ix18997 (.Y (nx18623), .A0 (nx15774), .A1 (nx18913)) ;
    inv02 ix18998 (.Y (nx18624), .A (write_offset_data_out_12)) ;
    inv02 ix18999 (.Y (nx18625), .A (write_base_data_out_12)) ;
    oai332 reg_nx4612 (.Y (nx4612), .A0 (nx18622), .A1 (nx18623), .A2 (nx17564)
           , .B0 (nx18623), .B1 (nx18624), .B2 (nx18625), .C0 (nx15774), .C1 (
           nx18913)) ;
    inv02 ix19000 (.Y (nx18626), .A (nx4612)) ;
    ao22 reg_nx17731 (.Y (nx17731), .A0 (nx18616), .A1 (nx18626), .B0 (nx17685)
         , .B1 (nx18616)) ;
    inv01 ix19001 (.Y (nx18627), .A (nx18626)) ;
    oai21 ix19002 (.Y (nx18628), .A0 (nx18624), .A1 (nx18625), .B0 (nx17564)) ;
    oai21 ix19003 (.Y (nx18629), .A0 (nx18624), .A1 (nx18625), .B0 (nx18622)) ;
    nand02_2x reg_nx17629 (.Y (nx17629), .A0 (nx18628), .A1 (nx18629)) ;
    inv02 ix19004 (.Y (nx18630), .A (nx15774)) ;
    inv01 ix19005 (.Y (nx18631), .A (nx18913)) ;
    oai22 reg_nx17632 (.Y (nx17632), .A0 (nx18630), .A1 (nx18631), .B0 (nx15774)
          , .B1 (nx18913)) ;
    inv01 reg_nx4328 (.Y (nx4328), .A (nx18622)) ;
    inv02 ix19006 (.Y (nx18632), .A (nx17437)) ;
    oai22 reg_nx17502 (.Y (nx17502), .A0 (nx18620), .A1 (nx4044), .B0 (nx18632)
          , .B1 (nx18620)) ;
    oai22 reg_nx17505 (.Y (nx17505), .A0 (nx18617), .A1 (nx18618), .B0 (nx15772)
          , .B1 (nx18908)) ;
    oai22 reg_nx17529 (.Y (nx17529), .A0 (nx18558), .A1 (nx18559), .B0 (nx18910)
          , .B1 (nx15795)) ;
    inv02 ix19007 (.Y (nx18633), .A (nx17529)) ;
    inv02 ix19008 (.Y (nx18634), .A (write_base_data_out_12)) ;
    or02 ix19009 (.Y (nx18635), .A0 (nx17887), .A1 (nx18912)) ;
    nand03_2x ix19010 (.Y (nx18636), .A0 (nx17526), .A1 (nx19294), .A2 (nx18633)
              ) ;
    oai321 reg_nx15151 (.Y (nx15151), .A0 (nx18679), .A1 (nx19302), .A2 (nx18633
           ), .B0 (nx18634), .B1 (nx18635), .C0 (nx18636)) ;
    inv02 reg_nx18267 (.Y (nx18267), .A (nx17887)) ;
    inv02 reg_nx18337 (.Y (nx18337), .A (nx18912)) ;
    nand02_2x ix19011 (.Y (nx18637), .A0 (img_addr_offset_3), .A1 (
              img_base_addr_3)) ;
    nand02_2x ix19012 (.Y (nx18638), .A0 (nx16915), .A1 (nx16911)) ;
    inv02 ix19013 (.Y (nx18639), .A (nx16818)) ;
    inv02 ix19014 (.Y (nx18640), .A (nx16833)) ;
    aoi22 ix19015 (.Y (nx18641), .A0 (nx16818), .A1 (nx16833), .B0 (nx18639), .B1 (
          nx18640)) ;
    and02 ix19016 (.Y (nx18642), .A0 (img_base_addr_0), .A1 (img_addr_offset_0)
          ) ;
    inv02 ix19017 (.Y (nx18643), .A (nx16915)) ;
    inv02 ix19018 (.Y (nx18644), .A (nx16911)) ;
    aoi332 ix19019 (.Y (nx18645), .A0 (nx18638), .A1 (img_addr_offset_1), .A2 (
           img_base_addr_1), .B0 (nx18641), .B1 (nx18638), .B2 (nx18642), .C0 (
           nx18643), .C1 (nx18644)) ;
    aoi22 ix19020 (.Y (nx18646), .A0 (nx18637), .A1 (nx18645), .B0 (nx16948), .B1 (
          nx18637)) ;
    inv01 reg_nx17023 (.Y (nx17023), .A (nx18646)) ;
    inv01 ix19021 (.Y (nx18647), .A (nx18646)) ;
    inv02 reg_nx3132 (.Y (nx3132), .A (nx18645)) ;
    and02 ix19022 (.Y (nx18648), .A0 (img_addr_offset_1), .A1 (img_base_addr_1)
          ) ;
    oai22 reg_nx16898 (.Y (nx16898), .A0 (nx18641), .A1 (nx18648), .B0 (nx18648)
          , .B1 (nx18642)) ;
    nor02_2x ix19023 (.Y (nx18649), .A0 (nx16915), .A1 (nx16911)) ;
    ao21 reg_nx16901 (.Y (nx16901), .A0 (nx16915), .A1 (nx16911), .B0 (nx18649)
         ) ;
    oai22 reg_nx16814 (.Y (nx16814), .A0 (nx18639), .A1 (nx18640), .B0 (nx16818)
          , .B1 (nx16833)) ;
    nand02_2x ix19024 (.Y (nx18650), .A0 (write_base_data_out_5), .A1 (
              bias_offset_data_out_5)) ;
    inv01 ix19025 (.Y (nx18651), .A (nx18583)) ;
    inv02 ix19026 (.Y (nx18652), .A (nx16967)) ;
    inv01 ix19027 (.Y (nx18653), .A (nx18891)) ;
    inv02 ix19028 (.Y (nx18654), .A (nx17021)) ;
    inv02 ix19029 (.Y (nx18655), .A (nx18582)) ;
    oai22 ix19030 (.Y (nx18656), .A0 (nx18655), .A1 (nx16967), .B0 (nx18584), .B1 (
          nx18585)) ;
    aoi322 ix19031 (.Y (nx18657), .A0 (nx18651), .A1 (nx18581), .A2 (nx18652), .B0 (
           nx18653), .B1 (nx18654), .C0 (nx18656), .C1 (nx18651)) ;
    aoi22 ix19032 (.Y (nx18658), .A0 (nx17081), .A1 (nx18650), .B0 (nx18650), .B1 (
          nx18657)) ;
    inv02 reg_nx17127 (.Y (nx17127), .A (nx18658)) ;
    inv02 ix19033 (.Y (nx18659), .A (nx18658)) ;
    nor02_2x ix19034 (.Y (nx18660), .A0 (nx18581), .A1 (nx18582)) ;
    nand02_2x ix19035 (.Y (nx18661), .A0 (nx18903), .A1 (nx15806)) ;
    inv01 ix19036 (.Y (nx18662), .A (nx18547)) ;
    and02 ix19037 (.Y (nx18663), .A0 (nx18578), .A1 (nx18662)) ;
    nor02_2x ix19038 (.Y (nx18664), .A0 (nx18903), .A1 (nx15806)) ;
    inv02 ix19039 (.Y (nx18665), .A (nx18577)) ;
    oai22 ix19040 (.Y (nx18666), .A0 (nx18910), .A1 (nx15795), .B0 (nx18665), .B1 (
          nx18547)) ;
    aoi321 ix19041 (.Y (nx18667), .A0 (nx18692), .A1 (nx18661), .A2 (nx18663), .B0 (
           nx18663), .B1 (nx18664), .C0 (nx18666)) ;
    inv02 ix19042 (.Y (nx18668), .A (new_size_squared_out_13)) ;
    inv01 ix19043 (.Y (nx18669), .A (nx18913)) ;
    aoi22 ix19044 (.Y (nx18670), .A0 (nx18914), .A1 (nx18668), .B0 (
          new_size_squared_out_13), .B1 (nx18669)) ;
    inv02 ix19045 (.Y (nx18671), .A (write_base_data_out_13)) ;
    oai22 ix19046 (.Y (nx18672), .A0 (nx18668), .A1 (nx18669), .B0 (
          new_size_squared_out_13), .B1 (nx18914)) ;
    nand03_2x ix19047 (.Y (nx18673), .A0 (nx18667), .A1 (nx19294), .A2 (nx18672)
              ) ;
    oai321 reg_nx15211 (.Y (nx15211), .A0 (nx18667), .A1 (nx19302), .A2 (nx18670
           ), .B0 (nx18671), .B1 (nx19296), .C0 (nx18673)) ;
    oai22 reg_nx17585 (.Y (nx17585), .A0 (nx18669), .A1 (new_size_squared_out_13
          ), .B0 (nx18668), .B1 (nx18914)) ;
    inv01 ix19048 (.Y (nx18674), .A (nx18903)) ;
    inv02 ix19049 (.Y (nx18675), .A (nx15806)) ;
    oai21 ix19050 (.Y (nx18676), .A0 (nx18674), .A1 (nx18675), .B0 (nx18578)) ;
    nor02_2x ix19051 (.Y (nx18677), .A0 (nx18664), .A1 (nx18577)) ;
    aoi22 ix19052 (.Y (nx18678), .A0 (nx18676), .A1 (nx18665), .B0 (nx18693), .B1 (
          nx18677)) ;
    inv02 reg_nx17526 (.Y (nx17526), .A (nx18678)) ;
    inv02 ix19053 (.Y (nx18679), .A (nx18678)) ;
    and02 ix19054 (.Y (nx18680), .A0 (nx18903), .A1 (nx15806)) ;
    ao21 reg_nx17402 (.Y (nx17402), .A0 (nx18904), .A1 (nx15806), .B0 (nx18664)
         ) ;
    and02 ix19055 (.Y (nx18681), .A0 (nx18893), .A1 (nx15827)) ;
    nor02_2x ix19056 (.Y (nx18682), .A0 (nx18681), .A1 (nx18881)) ;
    nor02_2x ix19057 (.Y (nx18683), .A0 (nx18893), .A1 (nx15827)) ;
    and02 ix19058 (.Y (nx18684), .A0 (nx18899), .A1 (nx15816)) ;
    inv02 ix19059 (.Y (nx18685), .A (nx18895)) ;
    inv02 ix19060 (.Y (nx18686), .A (new_size_squared_out_7)) ;
    inv02 ix19061 (.Y (nx18687), .A (nx18901)) ;
    inv02 ix19062 (.Y (nx18688), .A (new_size_squared_out_9)) ;
    inv01 reg_nx4194 (.Y (nx4194), .A (nx18805)) ;
    inv01 ix19063 (.Y (nx18689), .A (nx18805)) ;
    inv01 ix19064 (.Y (nx18690), .A (nx18805)) ;
    nand02_2x ix19065 (.Y (nx18691), .A0 (nx18901), .A1 (new_size_squared_out_9)
              ) ;
    aoi22 ix19066 (.Y (nx18692), .A0 (nx18691), .A1 (NOT_nx3910), .B0 (nx17331)
          , .B1 (nx18691)) ;
    inv02 reg_nx17399 (.Y (nx17399), .A (nx18692)) ;
    inv02 ix19067 (.Y (nx18693), .A (nx18692)) ;
    inv01 ix19068 (.Y (nx18694), .A (NOT_nx3910)) ;
    and02 ix19069 (.Y (nx18695), .A0 (nx18895), .A1 (new_size_squared_out_7)) ;
    inv02 ix19070 (.Y (nx18696), .A (nx17204)) ;
    oai32 reg_nx17272 (.Y (nx17272), .A0 (nx18695), .A1 (nx18682), .A2 (nx18683)
          , .B0 (nx18696), .B1 (nx18695)) ;
    inv02 ix19071 (.Y (nx18697), .A (nx18899)) ;
    inv02 ix19072 (.Y (nx18698), .A (nx15816)) ;
    oai22 reg_nx17275 (.Y (nx17275), .A0 (nx18697), .A1 (nx18698), .B0 (nx18899)
          , .B1 (nx15816)) ;
    oai22 reg_nx3626 (.Y (nx3626), .A0 (nx18893), .A1 (nx15827), .B0 (nx18681), 
          .B1 (nx18882)) ;
    inv02 ix19073 (.Y (nx18699), .A (nx18894)) ;
    inv02 ix19074 (.Y (nx18700), .A (nx15827)) ;
    oai22 reg_nx17145 (.Y (nx17145), .A0 (nx18699), .A1 (nx18700), .B0 (nx18894)
          , .B1 (nx15827)) ;
    inv02 ix19075 (.Y (nx18701), .A (nx18905)) ;
    inv02 ix19076 (.Y (nx18702), .A (write_base_data_out_12)) ;
    inv02 ix19077 (.Y (nx18703), .A (write_base_data_out_13)) ;
    inv02 ix19078 (.Y (nx18704), .A (nx3928)) ;
    inv01 ix19079 (.Y (nx18705), .A (nx18914)) ;
    inv02 ix19080 (.Y (nx18706), .A (nx18908)) ;
    nor04_2x ix19081 (.Y (nx18707), .A0 (write_base_data_out_12), .A1 (
             write_base_data_out_10), .A2 (nx18705), .A3 (nx18706)) ;
    and03 ix19082 (.Y (nx18708), .A0 (nx17431), .A1 (nx18704), .A2 (nx18707)) ;
    oai21 ix19083 (.Y (nx18709), .A0 (nx4496), .A1 (nx18708), .B0 (nx17323)) ;
    and02 ix19084 (.Y (nx18710), .A0 (write_base_data_out_12), .A1 (nx18906)) ;
    inv01 ix19085 (.Y (nx18711), .A (nx17431)) ;
    oai422 reg_nx4502 (.Y (nx4502), .A0 (nx17431), .A1 (nx18701), .A2 (nx18702)
           , .A3 (write_base_data_out_13), .B0 (nx18710), .B1 (nx18914), .C0 (
           nx18711), .C1 (nx18914)) ;
    nor02_2x ix19086 (.Y (nx18712), .A0 (nx18701), .A1 (nx17431)) ;
    oai32 ix19087 (.Y (nx18713), .A0 (nx18717), .A1 (nx18701), .A2 (
          write_base_data_out_12), .B0 (nx18702), .B1 (nx18712)) ;
    inv02 ix19088 (.Y (nx18714), .A (write_base_data_out_10)) ;
    nand04_2x ix19089 (.Y (nx18715), .A0 (nx18717), .A1 (nx18704), .A2 (nx18908)
              , .A3 (nx18714)) ;
    oai21 ix19090 (.Y (nx18716), .A0 (nx18701), .A1 (nx18717), .B0 (nx18715)) ;
    oai322 reg_nx17556 (.Y (nx17556), .A0 (nx18717), .A1 (nx18702), .A2 (nx18701
           ), .B0 (nx18906), .B1 (write_base_data_out_12), .C0 (nx18711), .C1 (
           write_base_data_out_12)) ;
    oai22 reg_nx4218 (.Y (nx4218), .A0 (nx18717), .A1 (nx18906), .B0 (nx18711), 
          .B1 (nx18908)) ;
    oai21 reg_nx17429 (.Y (nx17429), .A0 (nx3928), .A1 (write_base_data_out_10)
          , .B0 (nx18717)) ;
    nand02_2x reg_nx4168 (.Y (nx4168), .A0 (nx17429), .A1 (nx17323)) ;
    buf02 ix19091 (.Y (nx18717), .A (nx17431)) ;
    nand02_2x ix19092 (.Y (nx18718), .A0 (write_base_data_out_13), .A1 (
              bias_offset_data_out_13)) ;
    nand02_2x ix19093 (.Y (nx18719), .A0 (nx18904), .A1 (nx17392)) ;
    aoi21 ix19094 (.Y (nx18720), .A0 (nx18904), .A1 (nx17392), .B0 (nx17337)) ;
    nor02_2x ix19095 (.Y (nx18721), .A0 (nx18904), .A1 (nx17392)) ;
    and02 ix19096 (.Y (nx18722), .A0 (nx18910), .A1 (nx17519)) ;
    inv02 ix19097 (.Y (nx18723), .A (nx18906)) ;
    inv02 ix19098 (.Y (nx18724), .A (bias_offset_data_out_11)) ;
    inv02 reg_nx17638 (.Y (nx17638), .A (nx18851)) ;
    inv02 ix19099 (.Y (nx18725), .A (nx18851)) ;
    inv02 ix19100 (.Y (nx18726), .A (nx18850)) ;
    nand02_2x ix19101 (.Y (nx18727), .A0 (nx18906), .A1 (bias_offset_data_out_11
              )) ;
    inv02 ix19102 (.Y (nx18728), .A (nx17464)) ;
    and02 ix19103 (.Y (nx18729), .A0 (nx18906), .A1 (bias_offset_data_out_11)) ;
    nor02_2x ix19104 (.Y (nx18730), .A0 (nx18728), .A1 (nx18729)) ;
    ao21 reg_nx17511 (.Y (nx17511), .A0 (nx18727), .A1 (nx18875), .B0 (nx18730)
         ) ;
    nor02_2x ix19105 (.Y (nx18731), .A0 (nx18910), .A1 (nx17519)) ;
    ao21 reg_nx17514 (.Y (nx17514), .A0 (nx18910), .A1 (nx17519), .B0 (nx18731)
         ) ;
    inv02 reg_nx4296 (.Y (nx4296), .A (nx18875)) ;
    and02 ix19106 (.Y (nx18732), .A0 (nx18901), .A1 (bias_offset_data_out_9)) ;
    inv02 ix19107 (.Y (nx18733), .A (nx17337)) ;
    oai22 reg_nx17384 (.Y (nx17384), .A0 (nx18732), .A1 (nx18857), .B0 (nx18733)
          , .B1 (nx18732)) ;
    ao21 reg_nx17387 (.Y (nx17387), .A0 (nx18904), .A1 (nx17392), .B0 (nx18721)
         ) ;
    nor02_2x ix19108 (.Y (nx18734), .A0 (nx17186), .A1 (nx18594)) ;
    inv02 ix19109 (.Y (nx18735), .A (nx17051)) ;
    inv02 ix19110 (.Y (nx18736), .A (nx18593)) ;
    oai22 ix19111 (.Y (nx18737), .A0 (nx18736), .A1 (nx17051), .B0 (nx18595), .B1 (
          nx18596)) ;
    or02 ix19112 (.Y (nx18738), .A0 (nx15730), .A1 (nx17076)) ;
    oai21 ix19113 (.Y (nx18739), .A0 (nx17186), .A1 (nx18738), .B0 (nx18589)) ;
    inv01 ix19114 (.Y (nx18740), .A (nx18594)) ;
    inv02 ix19115 (.Y (nx18741), .A (nx15730)) ;
    inv02 ix19116 (.Y (nx18742), .A (nx17076)) ;
    aoi322 reg_NOT_nx3476 (.Y (NOT_nx3476), .A0 (nx18740), .A1 (nx18592), .A2 (
           nx18735), .B0 (nx18741), .B1 (nx18742), .C0 (nx18737), .C1 (nx18740)
           ) ;
    nor02_2x ix19117 (.Y (nx18743), .A0 (nx18593), .A1 (nx18592)) ;
    and02 ix19118 (.Y (nx18744), .A0 (nx17044), .A1 (nx17038)) ;
    nor02_2x ix19119 (.Y (nx18745), .A0 (nx18744), .A1 (nx18647)) ;
    nor02_2x ix19120 (.Y (nx18746), .A0 (nx17044), .A1 (nx17038)) ;
    nor02_2x ix19121 (.Y (nx18747), .A0 (nx18745), .A1 (nx18746)) ;
    and02 ix19122 (.Y (nx18748), .A0 (nx17168), .A1 (nx17164)) ;
    inv02 ix19123 (.Y (nx18749), .A (img_addr_offset_5)) ;
    inv02 ix19124 (.Y (nx18750), .A (img_base_addr_5)) ;
    oai332 reg_nx3682 (.Y (nx3682), .A0 (nx18747), .A1 (nx18748), .A2 (nx17089)
           , .B0 (nx18748), .B1 (nx18749), .B2 (nx18750), .C0 (nx17168), .C1 (
           nx17164)) ;
    inv01 ix19125 (.Y (nx18751), .A (nx3682)) ;
    and02 ix19126 (.Y (nx18752), .A0 (nx17298), .A1 (nx17294)) ;
    inv02 ix19127 (.Y (nx18753), .A (img_addr_offset_7)) ;
    inv02 ix19128 (.Y (nx18754), .A (img_base_addr_7)) ;
    oai332 ix19129 (.Y (nx18755), .A0 (nx18751), .A1 (nx18752), .A2 (nx17218), .B0 (
           nx18752), .B1 (nx18753), .B2 (nx18754), .C0 (nx17298), .C1 (nx17294)
           ) ;
    inv02 ix19130 (.Y (nx18756), .A (nx18755)) ;
    inv02 reg_nx3966 (.Y (nx3966), .A (nx18756)) ;
    oai21 ix19131 (.Y (nx18757), .A0 (nx18753), .A1 (nx18754), .B0 (nx17218)) ;
    oai21 ix19132 (.Y (nx18758), .A0 (nx18753), .A1 (nx18754), .B0 (nx18751)) ;
    nand02_2x reg_nx17279 (.Y (nx17279), .A0 (nx18757), .A1 (nx18758)) ;
    nor02_2x ix19133 (.Y (nx18759), .A0 (nx17298), .A1 (nx17294)) ;
    ao21 reg_nx17282 (.Y (nx17282), .A0 (nx17298), .A1 (nx17294), .B0 (nx18759)
         ) ;
    inv02 ix19134 (.Y (nx18760), .A (nx18751)) ;
    and02 ix19135 (.Y (nx18761), .A0 (img_addr_offset_5), .A1 (img_base_addr_5)
          ) ;
    inv02 ix19136 (.Y (nx18762), .A (nx17089)) ;
    oai32 reg_nx17149 (.Y (nx17149), .A0 (nx18761), .A1 (nx18745), .A2 (nx18746)
          , .B0 (nx18762), .B1 (nx18761)) ;
    nor02_2x ix19137 (.Y (nx18763), .A0 (nx17168), .A1 (nx17164)) ;
    ao21 reg_nx17152 (.Y (nx17152), .A0 (nx17168), .A1 (nx17164), .B0 (nx18763)
         ) ;
    oai22 reg_nx3398 (.Y (nx3398), .A0 (nx17044), .A1 (nx17038), .B0 (nx18744), 
          .B1 (nx18647)) ;
    ao21 reg_nx17026 (.Y (nx17026), .A0 (nx17044), .A1 (nx17038), .B0 (nx18746)
         ) ;
    nand02_2x ix19138 (.Y (nx18764), .A0 (nx18567), .A1 (nx18568)) ;
    nand02_2x ix19139 (.Y (nx18765), .A0 (nx18564), .A1 (nx18565)) ;
    inv02 ix19140 (.Y (nx18766), .A (nx3048)) ;
    and02 ix19141 (.Y (nx18767), .A0 (nx18891), .A1 (nx15837)) ;
    inv02 ix19142 (.Y (nx18768), .A (write_base_data_out_3)) ;
    inv02 ix19143 (.Y (nx18769), .A (new_size_squared_out_3)) ;
    inv01 reg_nx3342 (.Y (nx3342), .A (nx18879)) ;
    ao21 ix19144 (.Y (nx18770), .A0 (write_base_data_out_3), .A1 (
         new_size_squared_out_3), .B0 (nx3048)) ;
    oai21 ix19145 (.Y (nx18771), .A0 (nx18768), .A1 (nx18769), .B0 (nx18877)) ;
    nand02_2x reg_nx17006 (.Y (nx17006), .A0 (nx18770), .A1 (nx18771)) ;
    inv01 ix19146 (.Y (nx18772), .A (nx18891)) ;
    inv02 ix19147 (.Y (nx18773), .A (nx15837)) ;
    oai22 reg_nx17009 (.Y (nx17009), .A0 (nx18772), .A1 (nx18773), .B0 (nx18892)
          , .B1 (nx15837)) ;
    aoi22 ix19148 (.Y (nx18774), .A0 (nx18564), .A1 (nx18565), .B0 (nx18567), .B1 (
          nx18568)) ;
    inv02 ix19149 (.Y (nx18775), .A (nx18902)) ;
    inv02 ix19150 (.Y (nx18776), .A (write_base_data_out_10)) ;
    inv02 ix19151 (.Y (nx18777), .A (nx18897)) ;
    nor04_2x ix19152 (.Y (nx18778), .A0 (nx18775), .A1 (nx18703), .A2 (nx18776)
             , .A3 (nx18777)) ;
    inv01 ix19153 (.Y (nx18779), .A (nx18701)) ;
    inv02 ix19154 (.Y (nx18780), .A (nx18702)) ;
    and04 reg_nx4496 (.Y (nx4496), .A0 (nx3644), .A1 (nx18778), .A2 (nx18779), .A3 (
          nx18780)) ;
    and02 ix19155 (.Y (nx18781), .A0 (write_base_data_out_10), .A1 (nx18897)) ;
    nand03_2x reg_nx17431 (.Y (nx17431), .A0 (nx3644), .A1 (nx18902), .A2 (
              nx18781)) ;
    inv02 ix19156 (.Y (nx18782), .A (nx17067)) ;
    inv02 ix19157 (.Y (nx18783), .A (nx3360)) ;
    nor02_2x ix19158 (.Y (nx18784), .A0 (nx18897), .A1 (write_base_data_out_6)
             ) ;
    and02 ix19159 (.Y (nx18785), .A0 (nx17326), .A1 (nx17199)) ;
    inv01 ix19160 (.Y (nx18786), .A (nx18796)) ;
    and02 ix19161 (.Y (nx18787), .A0 (nx18898), .A1 (nx18896)) ;
    aoi43 ix19162 (.Y (nx18788), .A0 (nx18796), .A1 (nx18783), .A2 (nx18784), .A3 (
          nx18785), .B0 (nx18786), .B1 (nx18902), .B2 (nx18787)) ;
    nor02_2x reg_nx17323 (.Y (nx17323), .A0 (nx18782), .A1 (nx18788)) ;
    inv02 ix19163 (.Y (nx18789), .A (nx18902)) ;
    nand02_2x ix19164 (.Y (nx18790), .A0 (nx18789), .A1 (nx18787)) ;
    oai222 reg_nx3934 (.Y (nx3934), .A0 (nx18786), .A1 (nx17326), .B0 (nx18787)
           , .B1 (nx17326), .C0 (nx18796), .C1 (nx18790)) ;
    inv02 ix19165 (.Y (nx18791), .A (nx18896)) ;
    inv02 ix19166 (.Y (nx18792), .A (nx18898)) ;
    nor02_2x reg_nx3644 (.Y (nx3644), .A0 (nx18791), .A1 (nx18796)) ;
    inv02 ix19167 (.Y (nx18793), .A (write_base_data_out_6)) ;
    and04 ix19168 (.Y (nx18794), .A0 (nx18796), .A1 (nx18783), .A2 (nx17199), .A3 (
          nx18793)) ;
    nor02_2x ix19169 (.Y (nx18795), .A0 (nx18794), .A1 (nx3644)) ;
    nor02_2x reg_nx17196 (.Y (nx17196), .A0 (nx18782), .A1 (nx18795)) ;
    oai321 reg_nx3884 (.Y (nx3884), .A0 (nx18797), .A1 (nx18791), .A2 (nx18898)
           , .B0 (nx18792), .B1 (nx3644), .C0 (nx17196)) ;
    nor04_2x reg_nx3928 (.Y (nx3928), .A0 (nx18797), .A1 (nx18789), .A2 (nx18792
             ), .A3 (nx18791)) ;
    oai322 reg_nx17302 (.Y (nx17302), .A0 (nx18797), .A1 (nx18792), .A2 (nx18791
           ), .B0 (nx18898), .B1 (nx18896), .C0 (nx18786), .C1 (nx18898)) ;
    oai22 reg_nx3650 (.Y (nx3650), .A0 (nx18797), .A1 (nx18896), .B0 (nx18786), 
          .B1 (nx17199)) ;
    oai21 reg_nx17172 (.Y (nx17172), .A0 (nx3360), .A1 (write_base_data_out_6), 
          .B0 (nx18797)) ;
    nand02_2x reg_nx3600 (.Y (nx3600), .A0 (nx17067), .A1 (nx17172)) ;
    buf04 ix19170 (.Y (nx18796), .A (nx17175)) ;
    buf04 ix19171 (.Y (nx18797), .A (nx17175)) ;
    inv02 ix19172 (.Y (nx18798), .A (nx18683)) ;
    oai332 ix19173 (.Y (nx18799), .A0 (nx18684), .A1 (nx18798), .A2 (nx17204), .B0 (
           nx18684), .B1 (nx18685), .B2 (nx18686), .C0 (nx18900), .C1 (nx15816)
           ) ;
    nor02_2x ix19174 (.Y (nx18800), .A0 (nx18680), .A1 (nx17331)) ;
    inv01 ix19175 (.Y (nx18801), .A (nx18684)) ;
    inv02 ix19176 (.Y (nx18802), .A (nx17204)) ;
    nand03_2x ix19177 (.Y (nx18803), .A0 (nx18682), .A1 (nx18801), .A2 (nx18802)
              ) ;
    oai332 ix19178 (.Y (nx18804), .A0 (nx18803), .A1 (nx18680), .A2 (nx17331), .B0 (
           nx18687), .B1 (nx18680), .B2 (nx18688), .C0 (nx18904), .C1 (nx15806)
           ) ;
    aoi21 ix19179 (.Y (nx18805), .A0 (nx19298), .A1 (nx18800), .B0 (nx19300)) ;
    oai22 ix19180 (.Y (nx18806), .A0 (nx18798), .A1 (nx17204), .B0 (nx18685), .B1 (
          nx18686)) ;
    nor02_2x ix19181 (.Y (nx18807), .A0 (nx18900), .A1 (nx15816)) ;
    aoi321 reg_NOT_nx3910 (.Y (NOT_nx3910), .A0 (nx18801), .A1 (nx18682), .A2 (
           nx18802), .B0 (nx18806), .B1 (nx18801), .C0 (nx18807)) ;
    inv02 ix19182 (.Y (nx18808), .A (img_addr_offset_11)) ;
    inv02 ix19183 (.Y (nx18809), .A (img_base_addr_11)) ;
    oai21 ix19184 (.Y (nx18810), .A0 (nx18808), .A1 (nx18809), .B0 (nx17472)) ;
    and02 ix19185 (.Y (nx18811), .A0 (nx17425), .A1 (nx17421)) ;
    inv02 ix19186 (.Y (nx18812), .A (nx17548)) ;
    inv02 ix19187 (.Y (nx18813), .A (nx17552)) ;
    aoi22 ix19188 (.Y (nx18814), .A0 (nx17548), .A1 (nx17552), .B0 (nx18812), .B1 (
          nx18813)) ;
    oai22 ix19189 (.Y (nx18815), .A0 (nx18813), .A1 (nx17548), .B0 (nx18812), .B1 (
          nx17552)) ;
    nand02_2x ix19190 (.Y (nx18816), .A0 (nx18815), .A1 (nx17533)) ;
    oai21 reg_nx17531 (.Y (nx17531), .A0 (nx18839), .A1 (nx18814), .B0 (nx18816)
          ) ;
    inv02 ix19191 (.Y (nx18817), .A (nx17859)) ;
    ao32 reg_nx17571 (.Y (nx17571), .A0 (nx18716), .A1 (nx18884), .A2 (nx17323)
         , .B0 (nx18884), .B1 (nx18817)) ;
    nor02ii ix19192 (.Y (nx18818), .A0 (nx18713), .A1 (nx18716)) ;
    inv01 ix19193 (.Y (nx18819), .A (nx17561)) ;
    inv02 ix19194 (.Y (nx18820), .A (nx18143)) ;
    inv02 reg_nx18135 (.Y (nx18135), .A (nx2664)) ;
    oai22 ix19195 (.Y (nx18821), .A0 (nx18135), .A1 (nx17509), .B0 (nx17566), .B1 (
          nx18139)) ;
    aoi321 ix19196 (.Y (nx18822), .A0 (nx18818), .A1 (argmax_ready), .A2 (
           nx17323), .B0 (nx18819), .B1 (nx18820), .C0 (nx18821)) ;
    oai221 reg_mem_addr_out_12 (.Y (mem_addr_out[12]), .A0 (nx18091), .A1 (
           nx17531), .B0 (nx17556), .B1 (nx17571), .C0 (nx18822)) ;
    inv02 reg_nx18075 (.Y (nx18075), .A (argmax_ready)) ;
    oai22 reg_nx17536 (.Y (nx17536), .A0 (nx18812), .A1 (nx18813), .B0 (nx17548)
          , .B1 (nx17552)) ;
    inv01 ix19197 (.Y (nx18823), .A (nx18716)) ;
    inv02 ix19198 (.Y (nx18824), .A (nx17323)) ;
    nor03_2x reg_nx18213 (.Y (nx18213), .A0 (nx18713), .A1 (nx18823), .A2 (
             nx18824)) ;
    inv02 reg_nx17977 (.Y (nx17977), .A (nx18884)) ;
    oai22 reg_nx4250 (.Y (nx4250), .A0 (nx17425), .A1 (nx17421), .B0 (nx18811), 
          .B1 (nx17406)) ;
    and02 reg_nx17450 (.Y (nx17450), .A0 (nx18716), .A1 (nx17323)) ;
    nor02_2x ix19199 (.Y (nx18825), .A0 (nx17425), .A1 (nx17421)) ;
    ao21 reg_nx17409 (.Y (nx17409), .A0 (nx17425), .A1 (nx17421), .B0 (nx18825)
         ) ;
    inv02 ix19200 (.Y (nx18826), .A (nx15696)) ;
    inv02 ix19201 (.Y (nx18827), .A (nx17199)) ;
    nand02_2x ix19202 (.Y (nx18828), .A0 (nx15696), .A1 (nx17199)) ;
    or02 ix19203 (.Y (nx18829), .A0 (nx18737), .A1 (nx18739)) ;
    aoi21 ix19204 (.Y (nx18830), .A0 (nx18592), .A1 (nx18735), .B0 (nx18829)) ;
    nor02_2x ix19205 (.Y (nx18831), .A0 (nx18739), .A1 (nx18734)) ;
    and02 ix19206 (.Y (nx18832), .A0 (nx18592), .A1 (nx18735)) ;
    oai32 reg_nx17247 (.Y (nx17247), .A0 (nx18832), .A1 (nx18737), .A2 (nx18739)
          , .B0 (nx18739), .B1 (nx18734)) ;
    oai22 reg_nx17250 (.Y (nx17250), .A0 (nx18826), .A1 (nx18827), .B0 (nx15696)
          , .B1 (nx17199)) ;
    inv02 ix19207 (.Y (nx18833), .A (nx18756)) ;
    inv02 ix19208 (.Y (nx18834), .A (nx17345)) ;
    nor02ii ix19209 (.Y (nx18835), .A0 (nx18811), .A1 (nx18810)) ;
    oai22 ix19210 (.Y (nx18836), .A0 (nx17425), .A1 (nx17421), .B0 (nx18808), .B1 (
          nx18809)) ;
    and02 ix19211 (.Y (nx18837), .A0 (img_addr_offset_9), .A1 (img_base_addr_9)
          ) ;
    aoi322 ix19212 (.Y (nx18838), .A0 (nx18833), .A1 (nx18834), .A2 (nx18835), .B0 (
           nx18810), .B1 (nx18836), .C0 (nx18835), .C1 (nx18837)) ;
    inv02 reg_nx17533 (.Y (nx17533), .A (nx18838)) ;
    inv02 ix19213 (.Y (nx18839), .A (nx18838)) ;
    oai22 reg_nx17406 (.Y (nx17406), .A0 (nx18833), .A1 (nx18837), .B0 (nx18834)
          , .B1 (nx18837)) ;
    nand02_2x ix19214 (.Y (nx18840), .A0 (nx18826), .A1 (nx18827)) ;
    nor02ii ix19215 (.Y (nx18841), .A0 (nx18831), .A1 (nx18828)) ;
    and02 ix19216 (.Y (nx18842), .A0 (nx18826), .A1 (nx18827)) ;
    nor02_2x ix19217 (.Y (nx18843), .A0 (nx18841), .A1 (nx18842)) ;
    aoi21 reg_nx3760 (.Y (nx3760), .A0 (nx18830), .A1 (nx18840), .B0 (nx18843)
          ) ;
    inv01 reg_nx17577 (.Y (nx17577), .A (nx18709)) ;
    nand02_2x reg_nx4736 (.Y (nx4736), .A0 (nx17679), .A1 (nx17577)) ;
    nand02_2x ix19218 (.Y (nx18844), .A0 (nx18896), .A1 (bias_offset_data_out_7)
              ) ;
    and02 ix19219 (.Y (nx18845), .A0 (nx18894), .A1 (nx17135)) ;
    nor02_2x ix19220 (.Y (nx18846), .A0 (nx18894), .A1 (nx17135)) ;
    aoi22 ix19221 (.Y (nx18847), .A0 (nx18844), .A1 (nx18849), .B0 (nx17210), .B1 (
          nx18844)) ;
    inv01 reg_nx17257 (.Y (nx17257), .A (nx18847)) ;
    oai22 reg_nx3728 (.Y (nx3728), .A0 (nx18894), .A1 (nx17135), .B0 (nx18845), 
          .B1 (nx18659)) ;
    ao21 reg_nx17130 (.Y (nx17130), .A0 (nx18894), .A1 (nx17135), .B0 (nx18846)
         ) ;
    inv02 ix19222 (.Y (nx18848), .A (nx18846)) ;
    ao22 ix19223 (.Y (nx18849), .A0 (nx18845), .A1 (nx18848), .B0 (nx18659), .B1 (
         nx18848)) ;
    inv02 ix19224 (.Y (nx18850), .A (nx4580)) ;
    oai21 ix19225 (.Y (nx18851), .A0 (nx18850), .A1 (nx17591), .B0 (nx18718)) ;
    inv02 ix19226 (.Y (nx18852), .A (nx18900)) ;
    inv02 ix19227 (.Y (nx18853), .A (nx17265)) ;
    nand02_2x ix19228 (.Y (nx18854), .A0 (nx18900), .A1 (nx17265)) ;
    aoi22 ix19229 (.Y (nx18855), .A0 (nx18852), .A1 (nx18853), .B0 (nx18847), .B1 (
          nx18854)) ;
    inv02 reg_nx4012 (.Y (nx4012), .A (nx18855)) ;
    inv02 ix19230 (.Y (nx18856), .A (nx18855)) ;
    inv02 ix19231 (.Y (nx18857), .A (nx18855)) ;
    nor02_2x ix19232 (.Y (nx18858), .A0 (nx18900), .A1 (nx17265)) ;
    ao21 reg_nx17260 (.Y (nx17260), .A0 (nx18900), .A1 (nx17265), .B0 (nx18858)
         ) ;
    oai22 ix19233 (.Y (nx18859), .A0 (nx18892), .A1 (nx18890), .B0 (nx18892), .B1 (
          nx18887)) ;
    inv01 ix19234 (.Y (nx18860), .A (nx16934)) ;
    ao22 ix19235 (.Y (nx18861), .A0 (nx18892), .A1 (nx18890), .B0 (nx18892), .B1 (
         nx18887)) ;
    inv01 ix19236 (.Y (nx18862), .A (nx18888)) ;
    inv01 ix19237 (.Y (nx18863), .A (nx18892)) ;
    inv02 ix19238 (.Y (nx18864), .A (nx18890)) ;
    oai33 ix19239 (.Y (nx18865), .A0 (nx18862), .A1 (nx18863), .A2 (nx18864), .B0 (
          nx18888), .B1 (nx18892), .B2 (nx18890)) ;
    aoi221 ix19240 (.Y (nx18866), .A0 (nx18859), .A1 (nx18860), .B0 (nx16934), .B1 (
           nx18861), .C0 (nx18865)) ;
    inv01 reg_nx16998 (.Y (nx16998), .A (nx18866)) ;
    inv01 ix19241 (.Y (nx18867), .A (nx18866)) ;
    and02 ix19242 (.Y (nx18868), .A0 (nx18888), .A1 (nx18890)) ;
    oai22 reg_nx3216 (.Y (nx3216), .A0 (nx18888), .A1 (nx18890), .B0 (nx18868), 
          .B1 (nx16934)) ;
    oai22 reg_nx16937 (.Y (nx16937), .A0 (nx18862), .A1 (nx18864), .B0 (nx18888)
          , .B1 (nx18890)) ;
    nor02_2x ix19243 (.Y (nx18869), .A0 (nx18722), .A1 (nx17464)) ;
    nand03_2x ix19244 (.Y (nx18870), .A0 (nx18869), .A1 (nx18856), .A2 (nx18720)
              ) ;
    and03 ix19245 (.Y (nx18871), .A0 (nx18719), .A1 (nx18902), .A2 (
          bias_offset_data_out_9)) ;
    nor02_2x ix19246 (.Y (nx18872), .A0 (nx18871), .A1 (nx18721)) ;
    oai332 ix19247 (.Y (nx18873), .A0 (nx18872), .A1 (nx18722), .A2 (nx17464), .B0 (
           nx18723), .B1 (nx18722), .B2 (nx18724), .C0 (nx18910), .C1 (nx17519)
           ) ;
    inv02 ix19248 (.Y (nx18874), .A (nx18873)) ;
    nand02_2x reg_nx4580 (.Y (nx4580), .A0 (nx18870), .A1 (nx18874)) ;
    aoi321 ix19249 (.Y (nx18875), .A0 (nx18719), .A1 (nx18902), .A2 (
           bias_offset_data_out_9), .B0 (nx18856), .B1 (nx18720), .C0 (nx18721)
           ) ;
    nand02_2x ix19250 (.Y (nx18876), .A0 (write_base_data_out_5), .A1 (
              new_size_squared_out_5)) ;
    aoi32 ix19251 (.Y (nx18877), .A0 (nx18764), .A1 (nx18562), .A2 (nx18765), .B0 (
          nx18560), .B1 (nx18561)) ;
    oai332 ix19252 (.Y (nx18878), .A0 (nx18877), .A1 (nx18767), .A2 (nx18766), .B0 (
           nx18767), .B1 (nx18768), .B2 (nx18769), .C0 (nx18892), .C1 (nx15837)
           ) ;
    inv02 ix19253 (.Y (nx18879), .A (nx18878)) ;
    aoi22 ix19254 (.Y (nx18880), .A0 (nx17074), .A1 (nx18876), .B0 (nx18876), .B1 (
          nx18879)) ;
    inv02 reg_nx17142 (.Y (nx17142), .A (nx18880)) ;
    inv02 ix19255 (.Y (nx18881), .A (nx18880)) ;
    inv02 ix19256 (.Y (nx18882), .A (nx18880)) ;
    buf16 ix19257 (.Y (nx18883), .A (nx18309)) ;
    buf16 ix19258 (.Y (nx18884), .A (nx18309)) ;
    buf16 ix19259 (.Y (nx18885), .A (nx16878)) ;
    buf16 ix19260 (.Y (nx18886), .A (nx16878)) ;
    buf16 ix19261 (.Y (nx18887), .A (nx16348)) ;
    buf16 ix19262 (.Y (nx18888), .A (nx16348)) ;
    buf16 ix19263 (.Y (nx18889), .A (nx16945)) ;
    buf16 ix19264 (.Y (nx18890), .A (nx16945)) ;
    buf16 ix19265 (.Y (nx18891), .A (nx17002)) ;
    buf16 ix19266 (.Y (nx18892), .A (nx17002)) ;
    buf16 ix19267 (.Y (nx18893), .A (nx17138)) ;
    buf16 ix19268 (.Y (nx18894), .A (nx17138)) ;
    buf16 ix19269 (.Y (nx18895), .A (write_base_data_out_7)) ;
    buf16 ix19270 (.Y (nx18896), .A (write_base_data_out_7)) ;
    buf16 ix19271 (.Y (nx18897), .A (write_base_data_out_8)) ;
    buf16 ix19272 (.Y (nx18898), .A (write_base_data_out_8)) ;
    buf16 ix19273 (.Y (nx18899), .A (nx17268)) ;
    buf16 ix19274 (.Y (nx18900), .A (nx17268)) ;
    buf16 ix19275 (.Y (nx18901), .A (write_base_data_out_9)) ;
    buf16 ix19276 (.Y (nx18902), .A (write_base_data_out_9)) ;
    buf16 ix19277 (.Y (nx18903), .A (nx17395)) ;
    buf16 ix19278 (.Y (nx18904), .A (nx17395)) ;
    buf16 ix19279 (.Y (nx18905), .A (write_base_data_out_11)) ;
    buf16 ix19280 (.Y (nx18906), .A (write_base_data_out_11)) ;
    buf16 ix19281 (.Y (nx18907), .A (nx17453)) ;
    buf16 ix19282 (.Y (nx18908), .A (nx17453)) ;
    buf16 ix19283 (.Y (nx18909), .A (nx17522)) ;
    buf16 ix19284 (.Y (nx18910), .A (nx17522)) ;
    buf16 ix19285 (.Y (nx18911), .A (current_state_26)) ;
    buf16 ix19286 (.Y (nx18912), .A (current_state_26)) ;
    buf16 ix19287 (.Y (nx18913), .A (nx17580)) ;
    buf16 ix19288 (.Y (nx18914), .A (nx17580)) ;
    buf16 ix19289 (.Y (nx18915), .A (nx17649)) ;
    buf16 ix19290 (.Y (nx18916), .A (nx17649)) ;
    inv02 ix19291 (.Y (nx19292), .A (nx18219)) ;
    inv02 ix19293 (.Y (nx19294), .A (nx19292)) ;
    inv02 ix19295 (.Y (nx19296), .A (nx19292)) ;
    buf02 ix19297 (.Y (nx19298), .A (nx18799)) ;
    buf02 ix19299 (.Y (nx19300), .A (nx18804)) ;
    inv02 ix19301 (.Y (nx19302), .A (nx18219)) ;
    inv02 ix19307 (.Y (nx19308), .A (nx16222)) ;
endmodule


module AdvancedCounter_16 ( clk, reset, enable, mode_in, max_val_in, 
                            max_reached_out, counter_out ) ;

    input clk ;
    input reset ;
    input enable ;
    input [1:0]mode_in ;
    input [15:0]max_val_in ;
    output max_reached_out ;
    output [15:0]counter_out ;

    wire counter_out_15_rename, counter_out_14_rename, nx149, 
         counter_out_13_rename, counter_out_12_rename, nx152, 
         counter_out_11_rename, counter_out_10_rename, nx155, 
         counter_out_9_rename, counter_out_8_rename, nx157, counter_out_7_rename, 
         counter_out_6_rename, nx159, counter_out_5_rename, counter_out_4_rename, 
         nx161, counter_out_3_rename, counter_out_2_rename, counter_out_1_rename, 
         counter_out_dup0_0, nx22, nx34, nx46, nx70, nx94, nx118, nx142, nx166, 
         nx174, nx192, nx206, nx224, nx246, nx173, nx183, nx193, nx203, nx213, 
         nx223, nx233, nx243, nx253, nx263, nx273, nx283, nx293, nx303, nx313, 
         nx323, nx339, nx344, nx348, nx350, nx353, nx358, nx362, nx364, nx367, 
         nx372, nx376, nx378, nx381, nx386, nx390, nx392, nx395, nx400, nx404, 
         nx406, nx409, nx414, nx419, nx424, nx428, nx430, nx436, nx439, nx445, 
         nx447, nx449, nx451, nx458, nx460, nx462, nx464, nx466, nx468, nx470, 
         nx472, nx474;
    wire [1:0] \$dummy ;




    assign counter_out[14] = counter_out[15] ;
    assign counter_out[13] = counter_out[15] ;
    assign counter_out[12] = counter_out[15] ;
    assign counter_out[11] = counter_out[15] ;
    assign counter_out[10] = counter_out[15] ;
    assign counter_out[9] = counter_out[15] ;
    assign counter_out[8] = counter_out[15] ;
    assign counter_out[7] = counter_out[15] ;
    assign counter_out[6] = counter_out[15] ;
    assign counter_out[5] = counter_out[15] ;
    assign counter_out[4] = counter_out[15] ;
    assign counter_out[3] = counter_out[15] ;
    assign counter_out[2] = counter_out[15] ;
    assign counter_out[1] = counter_out[15] ;
    assign counter_out[0] = counter_out[15] ;
    fake_gnd ix140 (.Y (counter_out[15])) ;
    and04 ix251 (.Y (max_reached_out), .A0 (nx192), .A1 (nx206), .A2 (nx224), .A3 (
          nx246)) ;
    mux21_ni ix324 (.Y (nx323), .A0 (counter_out_15_rename), .A1 (nx174), .S0 (
             nx474)) ;
    mux21_ni ix314 (.Y (nx313), .A0 (counter_out_14_rename), .A1 (nx166), .S0 (
             nx472)) ;
    dffr reg_counter_data_14 (.Q (counter_out_14_rename), .QB (nx339), .D (nx313
         ), .CLK (clk), .R (nx462)) ;
    nand02 ix345 (.Y (nx344), .A0 (counter_out_13_rename), .A1 (nx152)) ;
    mux21 ix304 (.Y (nx303), .A0 (nx348), .A1 (nx350), .S0 (nx472)) ;
    dffr reg_counter_data_13 (.Q (counter_out_13_rename), .QB (nx348), .D (nx303
         ), .CLK (clk), .R (nx462)) ;
    oai21 ix351 (.Y (nx350), .A0 (nx152), .A1 (counter_out_13_rename), .B0 (
          nx344)) ;
    mux21_ni ix294 (.Y (nx293), .A0 (counter_out_12_rename), .A1 (nx142), .S0 (
             nx472)) ;
    dffr reg_counter_data_12 (.Q (counter_out_12_rename), .QB (nx353), .D (nx293
         ), .CLK (clk), .R (nx462)) ;
    nand02 ix359 (.Y (nx358), .A0 (counter_out_11_rename), .A1 (nx155)) ;
    mux21 ix284 (.Y (nx283), .A0 (nx362), .A1 (nx364), .S0 (nx472)) ;
    dffr reg_counter_data_11 (.Q (counter_out_11_rename), .QB (nx362), .D (nx283
         ), .CLK (clk), .R (nx462)) ;
    oai21 ix365 (.Y (nx364), .A0 (nx155), .A1 (counter_out_11_rename), .B0 (
          nx358)) ;
    mux21_ni ix274 (.Y (nx273), .A0 (counter_out_10_rename), .A1 (nx118), .S0 (
             nx472)) ;
    dffr reg_counter_data_10 (.Q (counter_out_10_rename), .QB (nx367), .D (nx273
         ), .CLK (clk), .R (nx462)) ;
    nand02 ix373 (.Y (nx372), .A0 (counter_out_9_rename), .A1 (nx157)) ;
    mux21 ix264 (.Y (nx263), .A0 (nx376), .A1 (nx378), .S0 (nx472)) ;
    dffr reg_counter_data_9 (.Q (counter_out_9_rename), .QB (nx376), .D (nx263)
         , .CLK (clk), .R (nx462)) ;
    oai21 ix379 (.Y (nx378), .A0 (nx157), .A1 (counter_out_9_rename), .B0 (nx372
          )) ;
    mux21_ni ix254 (.Y (nx253), .A0 (counter_out_8_rename), .A1 (nx94), .S0 (
             nx472)) ;
    dffr reg_counter_data_8 (.Q (counter_out_8_rename), .QB (nx381), .D (nx253)
         , .CLK (clk), .R (nx462)) ;
    nand02 ix387 (.Y (nx386), .A0 (counter_out_7_rename), .A1 (nx159)) ;
    mux21 ix244 (.Y (nx243), .A0 (nx390), .A1 (nx392), .S0 (nx470)) ;
    dffr reg_counter_data_7 (.Q (counter_out_7_rename), .QB (nx390), .D (nx243)
         , .CLK (clk), .R (nx464)) ;
    oai21 ix393 (.Y (nx392), .A0 (nx159), .A1 (counter_out_7_rename), .B0 (nx386
          )) ;
    mux21_ni ix234 (.Y (nx233), .A0 (counter_out_6_rename), .A1 (nx70), .S0 (
             nx470)) ;
    dffr reg_counter_data_6 (.Q (counter_out_6_rename), .QB (nx395), .D (nx233)
         , .CLK (clk), .R (nx464)) ;
    nand02 ix401 (.Y (nx400), .A0 (counter_out_5_rename), .A1 (nx161)) ;
    mux21 ix224 (.Y (nx223), .A0 (nx404), .A1 (nx406), .S0 (nx470)) ;
    dffr reg_counter_data_5 (.Q (counter_out_5_rename), .QB (nx404), .D (nx223)
         , .CLK (clk), .R (nx464)) ;
    oai21 ix407 (.Y (nx406), .A0 (nx161), .A1 (counter_out_5_rename), .B0 (nx400
          )) ;
    mux21_ni ix214 (.Y (nx213), .A0 (counter_out_4_rename), .A1 (nx46), .S0 (
             nx470)) ;
    dffr reg_counter_data_4 (.Q (counter_out_4_rename), .QB (nx409), .D (nx213)
         , .CLK (clk), .R (nx464)) ;
    aoi21 ix47 (.Y (nx46), .A0 (nx414), .A1 (nx409), .B0 (nx161)) ;
    nand04 ix415 (.Y (nx414), .A0 (counter_out_3_rename), .A1 (
           counter_out_2_rename), .A2 (counter_out_1_rename), .A3 (
           counter_out_dup0_0)) ;
    dffr reg_counter_data_3 (.Q (counter_out_3_rename), .QB (\$dummy [0]), .D (
         nx203), .CLK (clk), .R (nx466)) ;
    mux21_ni ix204 (.Y (nx203), .A0 (counter_out_3_rename), .A1 (nx34), .S0 (
             nx470)) ;
    xnor2 ix35 (.Y (nx34), .A0 (counter_out_3_rename), .A1 (nx419)) ;
    nand03 ix420 (.Y (nx419), .A0 (counter_out_2_rename), .A1 (
           counter_out_1_rename), .A2 (counter_out_dup0_0)) ;
    dffr reg_counter_data_2 (.Q (counter_out_2_rename), .QB (\$dummy [1]), .D (
         nx193), .CLK (clk), .R (nx464)) ;
    mux21_ni ix194 (.Y (nx193), .A0 (counter_out_2_rename), .A1 (nx22), .S0 (
             nx470)) ;
    xnor2 ix23 (.Y (nx22), .A0 (counter_out_2_rename), .A1 (nx424)) ;
    mux21 ix184 (.Y (nx183), .A0 (nx428), .A1 (nx430), .S0 (nx470)) ;
    dffr reg_counter_data_1 (.Q (counter_out_1_rename), .QB (nx428), .D (nx183)
         , .CLK (clk), .R (nx464)) ;
    oai21 ix431 (.Y (nx430), .A0 (counter_out_dup0_0), .A1 (counter_out_1_rename
          ), .B0 (nx424)) ;
    dffr reg_counter_data_0 (.Q (counter_out_dup0_0), .QB (nx436), .D (nx173), .CLK (
         clk), .R (nx464)) ;
    dffr reg_counter_data_15 (.Q (counter_out_15_rename), .QB (nx439), .D (nx323
         ), .CLK (clk), .R (nx466)) ;
    and04 ix247 (.Y (nx246), .A0 (nx445), .A1 (nx447), .A2 (nx449), .A3 (nx451)
          ) ;
    xnor2 ix448 (.Y (nx447), .A0 (counter_out_2_rename), .A1 (max_val_in[2])) ;
    xnor2 ix450 (.Y (nx449), .A0 (counter_out_3_rename), .A1 (max_val_in[3])) ;
    and04 ix193 (.Y (nx192), .A0 (nx439), .A1 (nx339), .A2 (nx348), .A3 (nx353)
          ) ;
    xor2 ix175 (.Y (nx174), .A0 (nx149), .A1 (counter_out_15_rename)) ;
    nor02ii ix173 (.Y (nx149), .A0 (nx344), .A1 (counter_out_14_rename)) ;
    xor2 ix167 (.Y (nx166), .A0 (nx339), .A1 (nx344)) ;
    nor02ii ix149 (.Y (nx152), .A0 (nx358), .A1 (counter_out_12_rename)) ;
    xor2 ix143 (.Y (nx142), .A0 (nx353), .A1 (nx358)) ;
    nor02ii ix125 (.Y (nx155), .A0 (nx372), .A1 (counter_out_10_rename)) ;
    xor2 ix119 (.Y (nx118), .A0 (nx367), .A1 (nx372)) ;
    nor02ii ix101 (.Y (nx157), .A0 (nx386), .A1 (counter_out_8_rename)) ;
    xor2 ix95 (.Y (nx94), .A0 (nx381), .A1 (nx386)) ;
    nor02ii ix77 (.Y (nx159), .A0 (nx400), .A1 (counter_out_6_rename)) ;
    xor2 ix71 (.Y (nx70), .A0 (nx395), .A1 (nx400)) ;
    nor02ii ix53 (.Y (nx161), .A0 (nx414), .A1 (counter_out_4_rename)) ;
    or02 ix425 (.Y (nx424), .A0 (nx428), .A1 (nx436)) ;
    xnor2 ix174 (.Y (nx173), .A0 (nx436), .A1 (nx474)) ;
    and04 ix207 (.Y (nx206), .A0 (nx362), .A1 (nx367), .A2 (nx376), .A3 (nx381)
          ) ;
    and04 ix225 (.Y (nx224), .A0 (nx390), .A1 (nx395), .A2 (nx404), .A3 (nx458)
          ) ;
    xnor2 ix217 (.Y (nx458), .A0 (max_val_in[0]), .A1 (counter_out_dup0_0)) ;
    xor2 ix446 (.Y (nx445), .A0 (nx428), .A1 (max_val_in[1])) ;
    xor2 ix452 (.Y (nx451), .A0 (nx409), .A1 (max_val_in[4])) ;
    inv01 ix459 (.Y (nx460), .A (reset)) ;
    inv02 ix461 (.Y (nx462), .A (nx460)) ;
    inv02 ix463 (.Y (nx464), .A (nx460)) ;
    inv02 ix465 (.Y (nx466), .A (nx460)) ;
    inv01 ix467 (.Y (nx468), .A (enable)) ;
    inv02 ix469 (.Y (nx470), .A (nx468)) ;
    inv02 ix471 (.Y (nx472), .A (nx468)) ;
    inv02 ix473 (.Y (nx474), .A (nx468)) ;
endmodule


module Cache_5_16_28_5 ( in_word, cache_in_sel, cache_out_sel, decoder_enable, 
                         out_column_0__15, out_column_0__14, out_column_0__13, 
                         out_column_0__12, out_column_0__11, out_column_0__10, 
                         out_column_0__9, out_column_0__8, out_column_0__7, 
                         out_column_0__6, out_column_0__5, out_column_0__4, 
                         out_column_0__3, out_column_0__2, out_column_0__1, 
                         out_column_0__0, out_column_1__15, out_column_1__14, 
                         out_column_1__13, out_column_1__12, out_column_1__11, 
                         out_column_1__10, out_column_1__9, out_column_1__8, 
                         out_column_1__7, out_column_1__6, out_column_1__5, 
                         out_column_1__4, out_column_1__3, out_column_1__2, 
                         out_column_1__1, out_column_1__0, out_column_2__15, 
                         out_column_2__14, out_column_2__13, out_column_2__12, 
                         out_column_2__11, out_column_2__10, out_column_2__9, 
                         out_column_2__8, out_column_2__7, out_column_2__6, 
                         out_column_2__5, out_column_2__4, out_column_2__3, 
                         out_column_2__2, out_column_2__1, out_column_2__0, 
                         out_column_3__15, out_column_3__14, out_column_3__13, 
                         out_column_3__12, out_column_3__11, out_column_3__10, 
                         out_column_3__9, out_column_3__8, out_column_3__7, 
                         out_column_3__6, out_column_3__5, out_column_3__4, 
                         out_column_3__3, out_column_3__2, out_column_3__1, 
                         out_column_3__0, out_column_4__15, out_column_4__14, 
                         out_column_4__13, out_column_4__12, out_column_4__11, 
                         out_column_4__10, out_column_4__9, out_column_4__8, 
                         out_column_4__7, out_column_4__6, out_column_4__5, 
                         out_column_4__4, out_column_4__3, out_column_4__2, 
                         out_column_4__1, out_column_4__0, clk, reset ) ;

    input [15:0]in_word ;
    input [4:0]cache_in_sel ;
    input [4:0]cache_out_sel ;
    input decoder_enable ;
    output out_column_0__15 ;
    output out_column_0__14 ;
    output out_column_0__13 ;
    output out_column_0__12 ;
    output out_column_0__11 ;
    output out_column_0__10 ;
    output out_column_0__9 ;
    output out_column_0__8 ;
    output out_column_0__7 ;
    output out_column_0__6 ;
    output out_column_0__5 ;
    output out_column_0__4 ;
    output out_column_0__3 ;
    output out_column_0__2 ;
    output out_column_0__1 ;
    output out_column_0__0 ;
    output out_column_1__15 ;
    output out_column_1__14 ;
    output out_column_1__13 ;
    output out_column_1__12 ;
    output out_column_1__11 ;
    output out_column_1__10 ;
    output out_column_1__9 ;
    output out_column_1__8 ;
    output out_column_1__7 ;
    output out_column_1__6 ;
    output out_column_1__5 ;
    output out_column_1__4 ;
    output out_column_1__3 ;
    output out_column_1__2 ;
    output out_column_1__1 ;
    output out_column_1__0 ;
    output out_column_2__15 ;
    output out_column_2__14 ;
    output out_column_2__13 ;
    output out_column_2__12 ;
    output out_column_2__11 ;
    output out_column_2__10 ;
    output out_column_2__9 ;
    output out_column_2__8 ;
    output out_column_2__7 ;
    output out_column_2__6 ;
    output out_column_2__5 ;
    output out_column_2__4 ;
    output out_column_2__3 ;
    output out_column_2__2 ;
    output out_column_2__1 ;
    output out_column_2__0 ;
    output out_column_3__15 ;
    output out_column_3__14 ;
    output out_column_3__13 ;
    output out_column_3__12 ;
    output out_column_3__11 ;
    output out_column_3__10 ;
    output out_column_3__9 ;
    output out_column_3__8 ;
    output out_column_3__7 ;
    output out_column_3__6 ;
    output out_column_3__5 ;
    output out_column_3__4 ;
    output out_column_3__3 ;
    output out_column_3__2 ;
    output out_column_3__1 ;
    output out_column_3__0 ;
    output out_column_4__15 ;
    output out_column_4__14 ;
    output out_column_4__13 ;
    output out_column_4__12 ;
    output out_column_4__11 ;
    output out_column_4__10 ;
    output out_column_4__9 ;
    output out_column_4__8 ;
    output out_column_4__7 ;
    output out_column_4__6 ;
    output out_column_4__5 ;
    output out_column_4__4 ;
    output out_column_4__3 ;
    output out_column_4__2 ;
    output out_column_4__1 ;
    output out_column_4__0 ;
    input clk ;
    input reset ;

    wire que_out_0__0__15, que_out_0__0__14, que_out_0__0__13, que_out_0__0__12, 
         que_out_0__0__11, que_out_0__0__10, que_out_0__0__9, que_out_0__0__8, 
         que_out_0__0__7, que_out_0__0__6, que_out_0__0__5, que_out_0__0__4, 
         que_out_0__0__3, que_out_0__0__2, que_out_0__0__1, que_out_0__0__0, 
         que_out_0__1__15, que_out_0__1__14, que_out_0__1__13, que_out_0__1__12, 
         que_out_0__1__11, que_out_0__1__10, que_out_0__1__9, que_out_0__1__8, 
         que_out_0__1__7, que_out_0__1__6, que_out_0__1__5, que_out_0__1__4, 
         que_out_0__1__3, que_out_0__1__2, que_out_0__1__1, que_out_0__1__0, 
         que_out_0__2__15, que_out_0__2__14, que_out_0__2__13, que_out_0__2__12, 
         que_out_0__2__11, que_out_0__2__10, que_out_0__2__9, que_out_0__2__8, 
         que_out_0__2__7, que_out_0__2__6, que_out_0__2__5, que_out_0__2__4, 
         que_out_0__2__3, que_out_0__2__2, que_out_0__2__1, que_out_0__2__0, 
         que_out_0__3__15, que_out_0__3__14, que_out_0__3__13, que_out_0__3__12, 
         que_out_0__3__11, que_out_0__3__10, que_out_0__3__9, que_out_0__3__8, 
         que_out_0__3__7, que_out_0__3__6, que_out_0__3__5, que_out_0__3__4, 
         que_out_0__3__3, que_out_0__3__2, que_out_0__3__1, que_out_0__3__0, 
         que_out_0__4__15, que_out_0__4__14, que_out_0__4__13, que_out_0__4__12, 
         que_out_0__4__11, que_out_0__4__10, que_out_0__4__9, que_out_0__4__8, 
         que_out_0__4__7, que_out_0__4__6, que_out_0__4__5, que_out_0__4__4, 
         que_out_0__4__3, que_out_0__4__2, que_out_0__4__1, que_out_0__4__0, 
         que_out_1__0__15, que_out_1__0__14, que_out_1__0__13, que_out_1__0__12, 
         que_out_1__0__11, que_out_1__0__10, que_out_1__0__9, que_out_1__0__8, 
         que_out_1__0__7, que_out_1__0__6, que_out_1__0__5, que_out_1__0__4, 
         que_out_1__0__3, que_out_1__0__2, que_out_1__0__1, que_out_1__0__0, 
         que_out_1__1__15, que_out_1__1__14, que_out_1__1__13, que_out_1__1__12, 
         que_out_1__1__11, que_out_1__1__10, que_out_1__1__9, que_out_1__1__8, 
         que_out_1__1__7, que_out_1__1__6, que_out_1__1__5, que_out_1__1__4, 
         que_out_1__1__3, que_out_1__1__2, que_out_1__1__1, que_out_1__1__0, 
         que_out_1__2__15, que_out_1__2__14, que_out_1__2__13, que_out_1__2__12, 
         que_out_1__2__11, que_out_1__2__10, que_out_1__2__9, que_out_1__2__8, 
         que_out_1__2__7, que_out_1__2__6, que_out_1__2__5, que_out_1__2__4, 
         que_out_1__2__3, que_out_1__2__2, que_out_1__2__1, que_out_1__2__0, 
         que_out_1__3__15, que_out_1__3__14, que_out_1__3__13, que_out_1__3__12, 
         que_out_1__3__11, que_out_1__3__10, que_out_1__3__9, que_out_1__3__8, 
         que_out_1__3__7, que_out_1__3__6, que_out_1__3__5, que_out_1__3__4, 
         que_out_1__3__3, que_out_1__3__2, que_out_1__3__1, que_out_1__3__0, 
         que_out_1__4__15, que_out_1__4__14, que_out_1__4__13, que_out_1__4__12, 
         que_out_1__4__11, que_out_1__4__10, que_out_1__4__9, que_out_1__4__8, 
         que_out_1__4__7, que_out_1__4__6, que_out_1__4__5, que_out_1__4__4, 
         que_out_1__4__3, que_out_1__4__2, que_out_1__4__1, que_out_1__4__0, 
         que_out_2__0__15, que_out_2__0__14, que_out_2__0__13, que_out_2__0__12, 
         que_out_2__0__11, que_out_2__0__10, que_out_2__0__9, que_out_2__0__8, 
         que_out_2__0__7, que_out_2__0__6, que_out_2__0__5, que_out_2__0__4, 
         que_out_2__0__3, que_out_2__0__2, que_out_2__0__1, que_out_2__0__0, 
         que_out_2__1__15, que_out_2__1__14, que_out_2__1__13, que_out_2__1__12, 
         que_out_2__1__11, que_out_2__1__10, que_out_2__1__9, que_out_2__1__8, 
         que_out_2__1__7, que_out_2__1__6, que_out_2__1__5, que_out_2__1__4, 
         que_out_2__1__3, que_out_2__1__2, que_out_2__1__1, que_out_2__1__0, 
         que_out_2__2__15, que_out_2__2__14, que_out_2__2__13, que_out_2__2__12, 
         que_out_2__2__11, que_out_2__2__10, que_out_2__2__9, que_out_2__2__8, 
         que_out_2__2__7, que_out_2__2__6, que_out_2__2__5, que_out_2__2__4, 
         que_out_2__2__3, que_out_2__2__2, que_out_2__2__1, que_out_2__2__0, 
         que_out_2__3__15, que_out_2__3__14, que_out_2__3__13, que_out_2__3__12, 
         que_out_2__3__11, que_out_2__3__10, que_out_2__3__9, que_out_2__3__8, 
         que_out_2__3__7, que_out_2__3__6, que_out_2__3__5, que_out_2__3__4, 
         que_out_2__3__3, que_out_2__3__2, que_out_2__3__1, que_out_2__3__0, 
         que_out_2__4__15, que_out_2__4__14, que_out_2__4__13, que_out_2__4__12, 
         que_out_2__4__11, que_out_2__4__10, que_out_2__4__9, que_out_2__4__8, 
         que_out_2__4__7, que_out_2__4__6, que_out_2__4__5, que_out_2__4__4, 
         que_out_2__4__3, que_out_2__4__2, que_out_2__4__1, que_out_2__4__0, 
         que_out_3__0__15, que_out_3__0__14, que_out_3__0__13, que_out_3__0__12, 
         que_out_3__0__11, que_out_3__0__10, que_out_3__0__9, que_out_3__0__8, 
         que_out_3__0__7, que_out_3__0__6, que_out_3__0__5, que_out_3__0__4, 
         que_out_3__0__3, que_out_3__0__2, que_out_3__0__1, que_out_3__0__0, 
         que_out_3__1__15, que_out_3__1__14, que_out_3__1__13, que_out_3__1__12, 
         que_out_3__1__11, que_out_3__1__10, que_out_3__1__9, que_out_3__1__8, 
         que_out_3__1__7, que_out_3__1__6, que_out_3__1__5, que_out_3__1__4, 
         que_out_3__1__3, que_out_3__1__2, que_out_3__1__1, que_out_3__1__0, 
         que_out_3__2__15, que_out_3__2__14, que_out_3__2__13, que_out_3__2__12, 
         que_out_3__2__11, que_out_3__2__10, que_out_3__2__9, que_out_3__2__8, 
         que_out_3__2__7, que_out_3__2__6, que_out_3__2__5, que_out_3__2__4, 
         que_out_3__2__3, que_out_3__2__2, que_out_3__2__1, que_out_3__2__0, 
         que_out_3__3__15, que_out_3__3__14, que_out_3__3__13, que_out_3__3__12, 
         que_out_3__3__11, que_out_3__3__10, que_out_3__3__9, que_out_3__3__8, 
         que_out_3__3__7, que_out_3__3__6, que_out_3__3__5, que_out_3__3__4, 
         que_out_3__3__3, que_out_3__3__2, que_out_3__3__1, que_out_3__3__0, 
         que_out_3__4__15, que_out_3__4__14, que_out_3__4__13, que_out_3__4__12, 
         que_out_3__4__11, que_out_3__4__10, que_out_3__4__9, que_out_3__4__8, 
         que_out_3__4__7, que_out_3__4__6, que_out_3__4__5, que_out_3__4__4, 
         que_out_3__4__3, que_out_3__4__2, que_out_3__4__1, que_out_3__4__0, 
         que_out_4__0__15, que_out_4__0__14, que_out_4__0__13, que_out_4__0__12, 
         que_out_4__0__11, que_out_4__0__10, que_out_4__0__9, que_out_4__0__8, 
         que_out_4__0__7, que_out_4__0__6, que_out_4__0__5, que_out_4__0__4, 
         que_out_4__0__3, que_out_4__0__2, que_out_4__0__1, que_out_4__0__0, 
         que_out_4__1__15, que_out_4__1__14, que_out_4__1__13, que_out_4__1__12, 
         que_out_4__1__11, que_out_4__1__10, que_out_4__1__9, que_out_4__1__8, 
         que_out_4__1__7, que_out_4__1__6, que_out_4__1__5, que_out_4__1__4, 
         que_out_4__1__3, que_out_4__1__2, que_out_4__1__1, que_out_4__1__0, 
         que_out_4__2__15, que_out_4__2__14, que_out_4__2__13, que_out_4__2__12, 
         que_out_4__2__11, que_out_4__2__10, que_out_4__2__9, que_out_4__2__8, 
         que_out_4__2__7, que_out_4__2__6, que_out_4__2__5, que_out_4__2__4, 
         que_out_4__2__3, que_out_4__2__2, que_out_4__2__1, que_out_4__2__0, 
         que_out_4__3__15, que_out_4__3__14, que_out_4__3__13, que_out_4__3__12, 
         que_out_4__3__11, que_out_4__3__10, que_out_4__3__9, que_out_4__3__8, 
         que_out_4__3__7, que_out_4__3__6, que_out_4__3__5, que_out_4__3__4, 
         que_out_4__3__3, que_out_4__3__2, que_out_4__3__1, que_out_4__3__0, 
         que_out_4__4__15, que_out_4__4__14, que_out_4__4__13, que_out_4__4__12, 
         que_out_4__4__11, que_out_4__4__10, que_out_4__4__9, que_out_4__4__8, 
         que_out_4__4__7, que_out_4__4__6, que_out_4__4__5, que_out_4__4__4, 
         que_out_4__4__3, que_out_4__4__2, que_out_4__4__1, que_out_4__4__0, 
         que_out_5__0__15, que_out_5__0__14, que_out_5__0__13, que_out_5__0__12, 
         que_out_5__0__11, que_out_5__0__10, que_out_5__0__9, que_out_5__0__8, 
         que_out_5__0__7, que_out_5__0__6, que_out_5__0__5, que_out_5__0__4, 
         que_out_5__0__3, que_out_5__0__2, que_out_5__0__1, que_out_5__0__0, 
         que_out_5__1__15, que_out_5__1__14, que_out_5__1__13, que_out_5__1__12, 
         que_out_5__1__11, que_out_5__1__10, que_out_5__1__9, que_out_5__1__8, 
         que_out_5__1__7, que_out_5__1__6, que_out_5__1__5, que_out_5__1__4, 
         que_out_5__1__3, que_out_5__1__2, que_out_5__1__1, que_out_5__1__0, 
         que_out_5__2__15, que_out_5__2__14, que_out_5__2__13, que_out_5__2__12, 
         que_out_5__2__11, que_out_5__2__10, que_out_5__2__9, que_out_5__2__8, 
         que_out_5__2__7, que_out_5__2__6, que_out_5__2__5, que_out_5__2__4, 
         que_out_5__2__3, que_out_5__2__2, que_out_5__2__1, que_out_5__2__0, 
         que_out_5__3__15, que_out_5__3__14, que_out_5__3__13, que_out_5__3__12, 
         que_out_5__3__11, que_out_5__3__10, que_out_5__3__9, que_out_5__3__8, 
         que_out_5__3__7, que_out_5__3__6, que_out_5__3__5, que_out_5__3__4, 
         que_out_5__3__3, que_out_5__3__2, que_out_5__3__1, que_out_5__3__0, 
         que_out_5__4__15, que_out_5__4__14, que_out_5__4__13, que_out_5__4__12, 
         que_out_5__4__11, que_out_5__4__10, que_out_5__4__9, que_out_5__4__8, 
         que_out_5__4__7, que_out_5__4__6, que_out_5__4__5, que_out_5__4__4, 
         que_out_5__4__3, que_out_5__4__2, que_out_5__4__1, que_out_5__4__0, 
         que_out_6__0__15, que_out_6__0__14, que_out_6__0__13, que_out_6__0__12, 
         que_out_6__0__11, que_out_6__0__10, que_out_6__0__9, que_out_6__0__8, 
         que_out_6__0__7, que_out_6__0__6, que_out_6__0__5, que_out_6__0__4, 
         que_out_6__0__3, que_out_6__0__2, que_out_6__0__1, que_out_6__0__0, 
         que_out_6__1__15, que_out_6__1__14, que_out_6__1__13, que_out_6__1__12, 
         que_out_6__1__11, que_out_6__1__10, que_out_6__1__9, que_out_6__1__8, 
         que_out_6__1__7, que_out_6__1__6, que_out_6__1__5, que_out_6__1__4, 
         que_out_6__1__3, que_out_6__1__2, que_out_6__1__1, que_out_6__1__0, 
         que_out_6__2__15, que_out_6__2__14, que_out_6__2__13, que_out_6__2__12, 
         que_out_6__2__11, que_out_6__2__10, que_out_6__2__9, que_out_6__2__8, 
         que_out_6__2__7, que_out_6__2__6, que_out_6__2__5, que_out_6__2__4, 
         que_out_6__2__3, que_out_6__2__2, que_out_6__2__1, que_out_6__2__0, 
         que_out_6__3__15, que_out_6__3__14, que_out_6__3__13, que_out_6__3__12, 
         que_out_6__3__11, que_out_6__3__10, que_out_6__3__9, que_out_6__3__8, 
         que_out_6__3__7, que_out_6__3__6, que_out_6__3__5, que_out_6__3__4, 
         que_out_6__3__3, que_out_6__3__2, que_out_6__3__1, que_out_6__3__0, 
         que_out_6__4__15, que_out_6__4__14, que_out_6__4__13, que_out_6__4__12, 
         que_out_6__4__11, que_out_6__4__10, que_out_6__4__9, que_out_6__4__8, 
         que_out_6__4__7, que_out_6__4__6, que_out_6__4__5, que_out_6__4__4, 
         que_out_6__4__3, que_out_6__4__2, que_out_6__4__1, que_out_6__4__0, 
         que_out_7__0__15, que_out_7__0__14, que_out_7__0__13, que_out_7__0__12, 
         que_out_7__0__11, que_out_7__0__10, que_out_7__0__9, que_out_7__0__8, 
         que_out_7__0__7, que_out_7__0__6, que_out_7__0__5, que_out_7__0__4, 
         que_out_7__0__3, que_out_7__0__2, que_out_7__0__1, que_out_7__0__0, 
         que_out_7__1__15, que_out_7__1__14, que_out_7__1__13, que_out_7__1__12, 
         que_out_7__1__11, que_out_7__1__10, que_out_7__1__9, que_out_7__1__8, 
         que_out_7__1__7, que_out_7__1__6, que_out_7__1__5, que_out_7__1__4, 
         que_out_7__1__3, que_out_7__1__2, que_out_7__1__1, que_out_7__1__0, 
         que_out_7__2__15, que_out_7__2__14, que_out_7__2__13, que_out_7__2__12, 
         que_out_7__2__11, que_out_7__2__10, que_out_7__2__9, que_out_7__2__8, 
         que_out_7__2__7, que_out_7__2__6, que_out_7__2__5, que_out_7__2__4, 
         que_out_7__2__3, que_out_7__2__2, que_out_7__2__1, que_out_7__2__0, 
         que_out_7__3__15, que_out_7__3__14, que_out_7__3__13, que_out_7__3__12, 
         que_out_7__3__11, que_out_7__3__10, que_out_7__3__9, que_out_7__3__8, 
         que_out_7__3__7, que_out_7__3__6, que_out_7__3__5, que_out_7__3__4, 
         que_out_7__3__3, que_out_7__3__2, que_out_7__3__1, que_out_7__3__0, 
         que_out_7__4__15, que_out_7__4__14, que_out_7__4__13, que_out_7__4__12, 
         que_out_7__4__11, que_out_7__4__10, que_out_7__4__9, que_out_7__4__8, 
         que_out_7__4__7, que_out_7__4__6, que_out_7__4__5, que_out_7__4__4, 
         que_out_7__4__3, que_out_7__4__2, que_out_7__4__1, que_out_7__4__0, 
         que_out_8__0__15, que_out_8__0__14, que_out_8__0__13, que_out_8__0__12, 
         que_out_8__0__11, que_out_8__0__10, que_out_8__0__9, que_out_8__0__8, 
         que_out_8__0__7, que_out_8__0__6, que_out_8__0__5, que_out_8__0__4, 
         que_out_8__0__3, que_out_8__0__2, que_out_8__0__1, que_out_8__0__0, 
         que_out_8__1__15, que_out_8__1__14, que_out_8__1__13, que_out_8__1__12, 
         que_out_8__1__11, que_out_8__1__10, que_out_8__1__9, que_out_8__1__8, 
         que_out_8__1__7, que_out_8__1__6, que_out_8__1__5, que_out_8__1__4, 
         que_out_8__1__3, que_out_8__1__2, que_out_8__1__1, que_out_8__1__0, 
         que_out_8__2__15, que_out_8__2__14, que_out_8__2__13, que_out_8__2__12, 
         que_out_8__2__11, que_out_8__2__10, que_out_8__2__9, que_out_8__2__8, 
         que_out_8__2__7, que_out_8__2__6, que_out_8__2__5, que_out_8__2__4, 
         que_out_8__2__3, que_out_8__2__2, que_out_8__2__1, que_out_8__2__0, 
         que_out_8__3__15, que_out_8__3__14, que_out_8__3__13, que_out_8__3__12, 
         que_out_8__3__11, que_out_8__3__10, que_out_8__3__9, que_out_8__3__8, 
         que_out_8__3__7, que_out_8__3__6, que_out_8__3__5, que_out_8__3__4, 
         que_out_8__3__3, que_out_8__3__2, que_out_8__3__1, que_out_8__3__0, 
         que_out_8__4__15, que_out_8__4__14, que_out_8__4__13, que_out_8__4__12, 
         que_out_8__4__11, que_out_8__4__10, que_out_8__4__9, que_out_8__4__8, 
         que_out_8__4__7, que_out_8__4__6, que_out_8__4__5, que_out_8__4__4, 
         que_out_8__4__3, que_out_8__4__2, que_out_8__4__1, que_out_8__4__0, 
         que_out_9__0__15, que_out_9__0__14, que_out_9__0__13, que_out_9__0__12, 
         que_out_9__0__11, que_out_9__0__10, que_out_9__0__9, que_out_9__0__8, 
         que_out_9__0__7, que_out_9__0__6, que_out_9__0__5, que_out_9__0__4, 
         que_out_9__0__3, que_out_9__0__2, que_out_9__0__1, que_out_9__0__0, 
         que_out_9__1__15, que_out_9__1__14, que_out_9__1__13, que_out_9__1__12, 
         que_out_9__1__11, que_out_9__1__10, que_out_9__1__9, que_out_9__1__8, 
         que_out_9__1__7, que_out_9__1__6, que_out_9__1__5, que_out_9__1__4, 
         que_out_9__1__3, que_out_9__1__2, que_out_9__1__1, que_out_9__1__0, 
         que_out_9__2__15, que_out_9__2__14, que_out_9__2__13, que_out_9__2__12, 
         que_out_9__2__11, que_out_9__2__10, que_out_9__2__9, que_out_9__2__8, 
         que_out_9__2__7, que_out_9__2__6, que_out_9__2__5, que_out_9__2__4, 
         que_out_9__2__3, que_out_9__2__2, que_out_9__2__1, que_out_9__2__0, 
         que_out_9__3__15, que_out_9__3__14, que_out_9__3__13, que_out_9__3__12, 
         que_out_9__3__11, que_out_9__3__10, que_out_9__3__9, que_out_9__3__8, 
         que_out_9__3__7, que_out_9__3__6, que_out_9__3__5, que_out_9__3__4, 
         que_out_9__3__3, que_out_9__3__2, que_out_9__3__1, que_out_9__3__0, 
         que_out_9__4__15, que_out_9__4__14, que_out_9__4__13, que_out_9__4__12, 
         que_out_9__4__11, que_out_9__4__10, que_out_9__4__9, que_out_9__4__8, 
         que_out_9__4__7, que_out_9__4__6, que_out_9__4__5, que_out_9__4__4, 
         que_out_9__4__3, que_out_9__4__2, que_out_9__4__1, que_out_9__4__0, 
         que_out_10__0__15, que_out_10__0__14, que_out_10__0__13, 
         que_out_10__0__12, que_out_10__0__11, que_out_10__0__10, 
         que_out_10__0__9, que_out_10__0__8, que_out_10__0__7, que_out_10__0__6, 
         que_out_10__0__5, que_out_10__0__4, que_out_10__0__3, que_out_10__0__2, 
         que_out_10__0__1, que_out_10__0__0, que_out_10__1__15, 
         que_out_10__1__14, que_out_10__1__13, que_out_10__1__12, 
         que_out_10__1__11, que_out_10__1__10, que_out_10__1__9, 
         que_out_10__1__8, que_out_10__1__7, que_out_10__1__6, que_out_10__1__5, 
         que_out_10__1__4, que_out_10__1__3, que_out_10__1__2, que_out_10__1__1, 
         que_out_10__1__0, que_out_10__2__15, que_out_10__2__14, 
         que_out_10__2__13, que_out_10__2__12, que_out_10__2__11, 
         que_out_10__2__10, que_out_10__2__9, que_out_10__2__8, que_out_10__2__7, 
         que_out_10__2__6, que_out_10__2__5, que_out_10__2__4, que_out_10__2__3, 
         que_out_10__2__2, que_out_10__2__1, que_out_10__2__0, que_out_10__3__15, 
         que_out_10__3__14, que_out_10__3__13, que_out_10__3__12, 
         que_out_10__3__11, que_out_10__3__10, que_out_10__3__9, 
         que_out_10__3__8, que_out_10__3__7, que_out_10__3__6, que_out_10__3__5, 
         que_out_10__3__4, que_out_10__3__3, que_out_10__3__2, que_out_10__3__1, 
         que_out_10__3__0, que_out_10__4__15, que_out_10__4__14, 
         que_out_10__4__13, que_out_10__4__12, que_out_10__4__11, 
         que_out_10__4__10, que_out_10__4__9, que_out_10__4__8, que_out_10__4__7, 
         que_out_10__4__6, que_out_10__4__5, que_out_10__4__4, que_out_10__4__3, 
         que_out_10__4__2, que_out_10__4__1, que_out_10__4__0, que_out_11__0__15, 
         que_out_11__0__14, que_out_11__0__13, que_out_11__0__12, 
         que_out_11__0__11, que_out_11__0__10, que_out_11__0__9, 
         que_out_11__0__8, que_out_11__0__7, que_out_11__0__6, que_out_11__0__5, 
         que_out_11__0__4, que_out_11__0__3, que_out_11__0__2, que_out_11__0__1, 
         que_out_11__0__0, que_out_11__1__15, que_out_11__1__14, 
         que_out_11__1__13, que_out_11__1__12, que_out_11__1__11, 
         que_out_11__1__10, que_out_11__1__9, que_out_11__1__8, que_out_11__1__7, 
         que_out_11__1__6, que_out_11__1__5, que_out_11__1__4, que_out_11__1__3, 
         que_out_11__1__2, que_out_11__1__1, que_out_11__1__0, que_out_11__2__15, 
         que_out_11__2__14, que_out_11__2__13, que_out_11__2__12, 
         que_out_11__2__11, que_out_11__2__10, que_out_11__2__9, 
         que_out_11__2__8, que_out_11__2__7, que_out_11__2__6, que_out_11__2__5, 
         que_out_11__2__4, que_out_11__2__3, que_out_11__2__2, que_out_11__2__1, 
         que_out_11__2__0, que_out_11__3__15, que_out_11__3__14, 
         que_out_11__3__13, que_out_11__3__12, que_out_11__3__11, 
         que_out_11__3__10, que_out_11__3__9, que_out_11__3__8, que_out_11__3__7, 
         que_out_11__3__6, que_out_11__3__5, que_out_11__3__4, que_out_11__3__3, 
         que_out_11__3__2, que_out_11__3__1, que_out_11__3__0, que_out_11__4__15, 
         que_out_11__4__14, que_out_11__4__13, que_out_11__4__12, 
         que_out_11__4__11, que_out_11__4__10, que_out_11__4__9, 
         que_out_11__4__8, que_out_11__4__7, que_out_11__4__6, que_out_11__4__5, 
         que_out_11__4__4, que_out_11__4__3, que_out_11__4__2, que_out_11__4__1, 
         que_out_11__4__0, que_out_12__0__15, que_out_12__0__14, 
         que_out_12__0__13, que_out_12__0__12, que_out_12__0__11, 
         que_out_12__0__10, que_out_12__0__9, que_out_12__0__8, que_out_12__0__7, 
         que_out_12__0__6, que_out_12__0__5, que_out_12__0__4, que_out_12__0__3, 
         que_out_12__0__2, que_out_12__0__1, que_out_12__0__0, que_out_12__1__15, 
         que_out_12__1__14, que_out_12__1__13, que_out_12__1__12, 
         que_out_12__1__11, que_out_12__1__10, que_out_12__1__9, 
         que_out_12__1__8, que_out_12__1__7, que_out_12__1__6, que_out_12__1__5, 
         que_out_12__1__4, que_out_12__1__3, que_out_12__1__2, que_out_12__1__1, 
         que_out_12__1__0, que_out_12__2__15, que_out_12__2__14, 
         que_out_12__2__13, que_out_12__2__12, que_out_12__2__11, 
         que_out_12__2__10, que_out_12__2__9, que_out_12__2__8, que_out_12__2__7, 
         que_out_12__2__6, que_out_12__2__5, que_out_12__2__4, que_out_12__2__3, 
         que_out_12__2__2, que_out_12__2__1, que_out_12__2__0, que_out_12__3__15, 
         que_out_12__3__14, que_out_12__3__13, que_out_12__3__12, 
         que_out_12__3__11, que_out_12__3__10, que_out_12__3__9, 
         que_out_12__3__8, que_out_12__3__7, que_out_12__3__6, que_out_12__3__5, 
         que_out_12__3__4, que_out_12__3__3, que_out_12__3__2, que_out_12__3__1, 
         que_out_12__3__0, que_out_12__4__15, que_out_12__4__14, 
         que_out_12__4__13, que_out_12__4__12, que_out_12__4__11, 
         que_out_12__4__10, que_out_12__4__9, que_out_12__4__8, que_out_12__4__7, 
         que_out_12__4__6, que_out_12__4__5, que_out_12__4__4, que_out_12__4__3, 
         que_out_12__4__2, que_out_12__4__1, que_out_12__4__0, que_out_13__0__15, 
         que_out_13__0__14, que_out_13__0__13, que_out_13__0__12, 
         que_out_13__0__11, que_out_13__0__10, que_out_13__0__9, 
         que_out_13__0__8, que_out_13__0__7, que_out_13__0__6, que_out_13__0__5, 
         que_out_13__0__4, que_out_13__0__3, que_out_13__0__2, que_out_13__0__1, 
         que_out_13__0__0, que_out_13__1__15, que_out_13__1__14, 
         que_out_13__1__13, que_out_13__1__12, que_out_13__1__11, 
         que_out_13__1__10, que_out_13__1__9, que_out_13__1__8, que_out_13__1__7, 
         que_out_13__1__6, que_out_13__1__5, que_out_13__1__4, que_out_13__1__3, 
         que_out_13__1__2, que_out_13__1__1, que_out_13__1__0, que_out_13__2__15, 
         que_out_13__2__14, que_out_13__2__13, que_out_13__2__12, 
         que_out_13__2__11, que_out_13__2__10, que_out_13__2__9, 
         que_out_13__2__8, que_out_13__2__7, que_out_13__2__6, que_out_13__2__5, 
         que_out_13__2__4, que_out_13__2__3, que_out_13__2__2, que_out_13__2__1, 
         que_out_13__2__0, que_out_13__3__15, que_out_13__3__14, 
         que_out_13__3__13, que_out_13__3__12, que_out_13__3__11, 
         que_out_13__3__10, que_out_13__3__9, que_out_13__3__8, que_out_13__3__7, 
         que_out_13__3__6, que_out_13__3__5, que_out_13__3__4, que_out_13__3__3, 
         que_out_13__3__2, que_out_13__3__1, que_out_13__3__0, que_out_13__4__15, 
         que_out_13__4__14, que_out_13__4__13, que_out_13__4__12, 
         que_out_13__4__11, que_out_13__4__10, que_out_13__4__9, 
         que_out_13__4__8, que_out_13__4__7, que_out_13__4__6, que_out_13__4__5, 
         que_out_13__4__4, que_out_13__4__3, que_out_13__4__2, que_out_13__4__1, 
         que_out_13__4__0, que_out_14__0__15, que_out_14__0__14, 
         que_out_14__0__13, que_out_14__0__12, que_out_14__0__11, 
         que_out_14__0__10, que_out_14__0__9, que_out_14__0__8, que_out_14__0__7, 
         que_out_14__0__6, que_out_14__0__5, que_out_14__0__4, que_out_14__0__3, 
         que_out_14__0__2, que_out_14__0__1, que_out_14__0__0, que_out_14__1__15, 
         que_out_14__1__14, que_out_14__1__13, que_out_14__1__12, 
         que_out_14__1__11, que_out_14__1__10, que_out_14__1__9, 
         que_out_14__1__8, que_out_14__1__7, que_out_14__1__6, que_out_14__1__5, 
         que_out_14__1__4, que_out_14__1__3, que_out_14__1__2, que_out_14__1__1, 
         que_out_14__1__0, que_out_14__2__15, que_out_14__2__14, 
         que_out_14__2__13, que_out_14__2__12, que_out_14__2__11, 
         que_out_14__2__10, que_out_14__2__9, que_out_14__2__8, que_out_14__2__7, 
         que_out_14__2__6, que_out_14__2__5, que_out_14__2__4, que_out_14__2__3, 
         que_out_14__2__2, que_out_14__2__1, que_out_14__2__0, que_out_14__3__15, 
         que_out_14__3__14, que_out_14__3__13, que_out_14__3__12, 
         que_out_14__3__11, que_out_14__3__10, que_out_14__3__9, 
         que_out_14__3__8, que_out_14__3__7, que_out_14__3__6, que_out_14__3__5, 
         que_out_14__3__4, que_out_14__3__3, que_out_14__3__2, que_out_14__3__1, 
         que_out_14__3__0, que_out_14__4__15, que_out_14__4__14, 
         que_out_14__4__13, que_out_14__4__12, que_out_14__4__11, 
         que_out_14__4__10, que_out_14__4__9, que_out_14__4__8, que_out_14__4__7, 
         que_out_14__4__6, que_out_14__4__5, que_out_14__4__4, que_out_14__4__3, 
         que_out_14__4__2, que_out_14__4__1, que_out_14__4__0, que_out_15__0__15, 
         que_out_15__0__14, que_out_15__0__13, que_out_15__0__12, 
         que_out_15__0__11, que_out_15__0__10, que_out_15__0__9, 
         que_out_15__0__8, que_out_15__0__7, que_out_15__0__6, que_out_15__0__5, 
         que_out_15__0__4, que_out_15__0__3, que_out_15__0__2, que_out_15__0__1, 
         que_out_15__0__0, que_out_15__1__15, que_out_15__1__14, 
         que_out_15__1__13, que_out_15__1__12, que_out_15__1__11, 
         que_out_15__1__10, que_out_15__1__9, que_out_15__1__8, que_out_15__1__7, 
         que_out_15__1__6, que_out_15__1__5, que_out_15__1__4, que_out_15__1__3, 
         que_out_15__1__2, que_out_15__1__1, que_out_15__1__0, que_out_15__2__15, 
         que_out_15__2__14, que_out_15__2__13, que_out_15__2__12, 
         que_out_15__2__11, que_out_15__2__10, que_out_15__2__9, 
         que_out_15__2__8, que_out_15__2__7, que_out_15__2__6, que_out_15__2__5, 
         que_out_15__2__4, que_out_15__2__3, que_out_15__2__2, que_out_15__2__1, 
         que_out_15__2__0, que_out_15__3__15, que_out_15__3__14, 
         que_out_15__3__13, que_out_15__3__12, que_out_15__3__11, 
         que_out_15__3__10, que_out_15__3__9, que_out_15__3__8, que_out_15__3__7, 
         que_out_15__3__6, que_out_15__3__5, que_out_15__3__4, que_out_15__3__3, 
         que_out_15__3__2, que_out_15__3__1, que_out_15__3__0, que_out_15__4__15, 
         que_out_15__4__14, que_out_15__4__13, que_out_15__4__12, 
         que_out_15__4__11, que_out_15__4__10, que_out_15__4__9, 
         que_out_15__4__8, que_out_15__4__7, que_out_15__4__6, que_out_15__4__5, 
         que_out_15__4__4, que_out_15__4__3, que_out_15__4__2, que_out_15__4__1, 
         que_out_15__4__0, que_out_16__0__15, que_out_16__0__14, 
         que_out_16__0__13, que_out_16__0__12, que_out_16__0__11, 
         que_out_16__0__10, que_out_16__0__9, que_out_16__0__8, que_out_16__0__7, 
         que_out_16__0__6, que_out_16__0__5, que_out_16__0__4, que_out_16__0__3, 
         que_out_16__0__2, que_out_16__0__1, que_out_16__0__0, que_out_16__1__15, 
         que_out_16__1__14, que_out_16__1__13, que_out_16__1__12, 
         que_out_16__1__11, que_out_16__1__10, que_out_16__1__9, 
         que_out_16__1__8, que_out_16__1__7, que_out_16__1__6, que_out_16__1__5, 
         que_out_16__1__4, que_out_16__1__3, que_out_16__1__2, que_out_16__1__1, 
         que_out_16__1__0, que_out_16__2__15, que_out_16__2__14, 
         que_out_16__2__13, que_out_16__2__12, que_out_16__2__11, 
         que_out_16__2__10, que_out_16__2__9, que_out_16__2__8, que_out_16__2__7, 
         que_out_16__2__6, que_out_16__2__5, que_out_16__2__4, que_out_16__2__3, 
         que_out_16__2__2, que_out_16__2__1, que_out_16__2__0, que_out_16__3__15, 
         que_out_16__3__14, que_out_16__3__13, que_out_16__3__12, 
         que_out_16__3__11, que_out_16__3__10, que_out_16__3__9, 
         que_out_16__3__8, que_out_16__3__7, que_out_16__3__6, que_out_16__3__5, 
         que_out_16__3__4, que_out_16__3__3, que_out_16__3__2, que_out_16__3__1, 
         que_out_16__3__0, que_out_16__4__15, que_out_16__4__14, 
         que_out_16__4__13, que_out_16__4__12, que_out_16__4__11, 
         que_out_16__4__10, que_out_16__4__9, que_out_16__4__8, que_out_16__4__7, 
         que_out_16__4__6, que_out_16__4__5, que_out_16__4__4, que_out_16__4__3, 
         que_out_16__4__2, que_out_16__4__1, que_out_16__4__0, que_out_17__0__15, 
         que_out_17__0__14, que_out_17__0__13, que_out_17__0__12, 
         que_out_17__0__11, que_out_17__0__10, que_out_17__0__9, 
         que_out_17__0__8, que_out_17__0__7, que_out_17__0__6, que_out_17__0__5, 
         que_out_17__0__4, que_out_17__0__3, que_out_17__0__2, que_out_17__0__1, 
         que_out_17__0__0, que_out_17__1__15, que_out_17__1__14, 
         que_out_17__1__13, que_out_17__1__12, que_out_17__1__11, 
         que_out_17__1__10, que_out_17__1__9, que_out_17__1__8, que_out_17__1__7, 
         que_out_17__1__6, que_out_17__1__5, que_out_17__1__4, que_out_17__1__3, 
         que_out_17__1__2, que_out_17__1__1, que_out_17__1__0, que_out_17__2__15, 
         que_out_17__2__14, que_out_17__2__13, que_out_17__2__12, 
         que_out_17__2__11, que_out_17__2__10, que_out_17__2__9, 
         que_out_17__2__8, que_out_17__2__7, que_out_17__2__6, que_out_17__2__5, 
         que_out_17__2__4, que_out_17__2__3, que_out_17__2__2, que_out_17__2__1, 
         que_out_17__2__0, que_out_17__3__15, que_out_17__3__14, 
         que_out_17__3__13, que_out_17__3__12, que_out_17__3__11, 
         que_out_17__3__10, que_out_17__3__9, que_out_17__3__8, que_out_17__3__7, 
         que_out_17__3__6, que_out_17__3__5, que_out_17__3__4, que_out_17__3__3, 
         que_out_17__3__2, que_out_17__3__1, que_out_17__3__0, que_out_17__4__15, 
         que_out_17__4__14, que_out_17__4__13, que_out_17__4__12, 
         que_out_17__4__11, que_out_17__4__10, que_out_17__4__9, 
         que_out_17__4__8, que_out_17__4__7, que_out_17__4__6, que_out_17__4__5, 
         que_out_17__4__4, que_out_17__4__3, que_out_17__4__2, que_out_17__4__1, 
         que_out_17__4__0, que_out_18__0__15, que_out_18__0__14, 
         que_out_18__0__13, que_out_18__0__12, que_out_18__0__11, 
         que_out_18__0__10, que_out_18__0__9, que_out_18__0__8, que_out_18__0__7, 
         que_out_18__0__6, que_out_18__0__5, que_out_18__0__4, que_out_18__0__3, 
         que_out_18__0__2, que_out_18__0__1, que_out_18__0__0, que_out_18__1__15, 
         que_out_18__1__14, que_out_18__1__13, que_out_18__1__12, 
         que_out_18__1__11, que_out_18__1__10, que_out_18__1__9, 
         que_out_18__1__8, que_out_18__1__7, que_out_18__1__6, que_out_18__1__5, 
         que_out_18__1__4, que_out_18__1__3, que_out_18__1__2, que_out_18__1__1, 
         que_out_18__1__0, que_out_18__2__15, que_out_18__2__14, 
         que_out_18__2__13, que_out_18__2__12, que_out_18__2__11, 
         que_out_18__2__10, que_out_18__2__9, que_out_18__2__8, que_out_18__2__7, 
         que_out_18__2__6, que_out_18__2__5, que_out_18__2__4, que_out_18__2__3, 
         que_out_18__2__2, que_out_18__2__1, que_out_18__2__0, que_out_18__3__15, 
         que_out_18__3__14, que_out_18__3__13, que_out_18__3__12, 
         que_out_18__3__11, que_out_18__3__10, que_out_18__3__9, 
         que_out_18__3__8, que_out_18__3__7, que_out_18__3__6, que_out_18__3__5, 
         que_out_18__3__4, que_out_18__3__3, que_out_18__3__2, que_out_18__3__1, 
         que_out_18__3__0, que_out_18__4__15, que_out_18__4__14, 
         que_out_18__4__13, que_out_18__4__12, que_out_18__4__11, 
         que_out_18__4__10, que_out_18__4__9, que_out_18__4__8, que_out_18__4__7, 
         que_out_18__4__6, que_out_18__4__5, que_out_18__4__4, que_out_18__4__3, 
         que_out_18__4__2, que_out_18__4__1, que_out_18__4__0, que_out_19__0__15, 
         que_out_19__0__14, que_out_19__0__13, que_out_19__0__12, 
         que_out_19__0__11, que_out_19__0__10, que_out_19__0__9, 
         que_out_19__0__8, que_out_19__0__7, que_out_19__0__6, que_out_19__0__5, 
         que_out_19__0__4, que_out_19__0__3, que_out_19__0__2, que_out_19__0__1, 
         que_out_19__0__0, que_out_19__1__15, que_out_19__1__14, 
         que_out_19__1__13, que_out_19__1__12, que_out_19__1__11, 
         que_out_19__1__10, que_out_19__1__9, que_out_19__1__8, que_out_19__1__7, 
         que_out_19__1__6, que_out_19__1__5, que_out_19__1__4, que_out_19__1__3, 
         que_out_19__1__2, que_out_19__1__1, que_out_19__1__0, que_out_19__2__15, 
         que_out_19__2__14, que_out_19__2__13, que_out_19__2__12, 
         que_out_19__2__11, que_out_19__2__10, que_out_19__2__9, 
         que_out_19__2__8, que_out_19__2__7, que_out_19__2__6, que_out_19__2__5, 
         que_out_19__2__4, que_out_19__2__3, que_out_19__2__2, que_out_19__2__1, 
         que_out_19__2__0, que_out_19__3__15, que_out_19__3__14, 
         que_out_19__3__13, que_out_19__3__12, que_out_19__3__11, 
         que_out_19__3__10, que_out_19__3__9, que_out_19__3__8, que_out_19__3__7, 
         que_out_19__3__6, que_out_19__3__5, que_out_19__3__4, que_out_19__3__3, 
         que_out_19__3__2, que_out_19__3__1, que_out_19__3__0, que_out_19__4__15, 
         que_out_19__4__14, que_out_19__4__13, que_out_19__4__12, 
         que_out_19__4__11, que_out_19__4__10, que_out_19__4__9, 
         que_out_19__4__8, que_out_19__4__7, que_out_19__4__6, que_out_19__4__5, 
         que_out_19__4__4, que_out_19__4__3, que_out_19__4__2, que_out_19__4__1, 
         que_out_19__4__0, que_out_20__0__15, que_out_20__0__14, 
         que_out_20__0__13, que_out_20__0__12, que_out_20__0__11, 
         que_out_20__0__10, que_out_20__0__9, que_out_20__0__8, que_out_20__0__7, 
         que_out_20__0__6, que_out_20__0__5, que_out_20__0__4, que_out_20__0__3, 
         que_out_20__0__2, que_out_20__0__1, que_out_20__0__0, que_out_20__1__15, 
         que_out_20__1__14, que_out_20__1__13, que_out_20__1__12, 
         que_out_20__1__11, que_out_20__1__10, que_out_20__1__9, 
         que_out_20__1__8, que_out_20__1__7, que_out_20__1__6, que_out_20__1__5, 
         que_out_20__1__4, que_out_20__1__3, que_out_20__1__2, que_out_20__1__1, 
         que_out_20__1__0, que_out_20__2__15, que_out_20__2__14, 
         que_out_20__2__13, que_out_20__2__12, que_out_20__2__11, 
         que_out_20__2__10, que_out_20__2__9, que_out_20__2__8, que_out_20__2__7, 
         que_out_20__2__6, que_out_20__2__5, que_out_20__2__4, que_out_20__2__3, 
         que_out_20__2__2, que_out_20__2__1, que_out_20__2__0, que_out_20__3__15, 
         que_out_20__3__14, que_out_20__3__13, que_out_20__3__12, 
         que_out_20__3__11, que_out_20__3__10, que_out_20__3__9, 
         que_out_20__3__8, que_out_20__3__7, que_out_20__3__6, que_out_20__3__5, 
         que_out_20__3__4, que_out_20__3__3, que_out_20__3__2, que_out_20__3__1, 
         que_out_20__3__0, que_out_20__4__15, que_out_20__4__14, 
         que_out_20__4__13, que_out_20__4__12, que_out_20__4__11, 
         que_out_20__4__10, que_out_20__4__9, que_out_20__4__8, que_out_20__4__7, 
         que_out_20__4__6, que_out_20__4__5, que_out_20__4__4, que_out_20__4__3, 
         que_out_20__4__2, que_out_20__4__1, que_out_20__4__0, que_out_21__0__15, 
         que_out_21__0__14, que_out_21__0__13, que_out_21__0__12, 
         que_out_21__0__11, que_out_21__0__10, que_out_21__0__9, 
         que_out_21__0__8, que_out_21__0__7, que_out_21__0__6, que_out_21__0__5, 
         que_out_21__0__4, que_out_21__0__3, que_out_21__0__2, que_out_21__0__1, 
         que_out_21__0__0, que_out_21__1__15, que_out_21__1__14, 
         que_out_21__1__13, que_out_21__1__12, que_out_21__1__11, 
         que_out_21__1__10, que_out_21__1__9, que_out_21__1__8, que_out_21__1__7, 
         que_out_21__1__6, que_out_21__1__5, que_out_21__1__4, que_out_21__1__3, 
         que_out_21__1__2, que_out_21__1__1, que_out_21__1__0, que_out_21__2__15, 
         que_out_21__2__14, que_out_21__2__13, que_out_21__2__12, 
         que_out_21__2__11, que_out_21__2__10, que_out_21__2__9, 
         que_out_21__2__8, que_out_21__2__7, que_out_21__2__6, que_out_21__2__5, 
         que_out_21__2__4, que_out_21__2__3, que_out_21__2__2, que_out_21__2__1, 
         que_out_21__2__0, que_out_21__3__15, que_out_21__3__14, 
         que_out_21__3__13, que_out_21__3__12, que_out_21__3__11, 
         que_out_21__3__10, que_out_21__3__9, que_out_21__3__8, que_out_21__3__7, 
         que_out_21__3__6, que_out_21__3__5, que_out_21__3__4, que_out_21__3__3, 
         que_out_21__3__2, que_out_21__3__1, que_out_21__3__0, que_out_21__4__15, 
         que_out_21__4__14, que_out_21__4__13, que_out_21__4__12, 
         que_out_21__4__11, que_out_21__4__10, que_out_21__4__9, 
         que_out_21__4__8, que_out_21__4__7, que_out_21__4__6, que_out_21__4__5, 
         que_out_21__4__4, que_out_21__4__3, que_out_21__4__2, que_out_21__4__1, 
         que_out_21__4__0, que_out_22__0__15, que_out_22__0__14, 
         que_out_22__0__13, que_out_22__0__12, que_out_22__0__11, 
         que_out_22__0__10, que_out_22__0__9, que_out_22__0__8, que_out_22__0__7, 
         que_out_22__0__6, que_out_22__0__5, que_out_22__0__4, que_out_22__0__3, 
         que_out_22__0__2, que_out_22__0__1, que_out_22__0__0, que_out_22__1__15, 
         que_out_22__1__14, que_out_22__1__13, que_out_22__1__12, 
         que_out_22__1__11, que_out_22__1__10, que_out_22__1__9, 
         que_out_22__1__8, que_out_22__1__7, que_out_22__1__6, que_out_22__1__5, 
         que_out_22__1__4, que_out_22__1__3, que_out_22__1__2, que_out_22__1__1, 
         que_out_22__1__0, que_out_22__2__15, que_out_22__2__14, 
         que_out_22__2__13, que_out_22__2__12, que_out_22__2__11, 
         que_out_22__2__10, que_out_22__2__9, que_out_22__2__8, que_out_22__2__7, 
         que_out_22__2__6, que_out_22__2__5, que_out_22__2__4, que_out_22__2__3, 
         que_out_22__2__2, que_out_22__2__1, que_out_22__2__0, que_out_22__3__15, 
         que_out_22__3__14, que_out_22__3__13, que_out_22__3__12, 
         que_out_22__3__11, que_out_22__3__10, que_out_22__3__9, 
         que_out_22__3__8, que_out_22__3__7, que_out_22__3__6, que_out_22__3__5, 
         que_out_22__3__4, que_out_22__3__3, que_out_22__3__2, que_out_22__3__1, 
         que_out_22__3__0, que_out_22__4__15, que_out_22__4__14, 
         que_out_22__4__13, que_out_22__4__12, que_out_22__4__11, 
         que_out_22__4__10, que_out_22__4__9, que_out_22__4__8, que_out_22__4__7, 
         que_out_22__4__6, que_out_22__4__5, que_out_22__4__4, que_out_22__4__3, 
         que_out_22__4__2, que_out_22__4__1, que_out_22__4__0, que_out_23__0__15, 
         que_out_23__0__14, que_out_23__0__13, que_out_23__0__12, 
         que_out_23__0__11, que_out_23__0__10, que_out_23__0__9, 
         que_out_23__0__8, que_out_23__0__7, que_out_23__0__6, que_out_23__0__5, 
         que_out_23__0__4, que_out_23__0__3, que_out_23__0__2, que_out_23__0__1, 
         que_out_23__0__0, que_out_23__1__15, que_out_23__1__14, 
         que_out_23__1__13, que_out_23__1__12, que_out_23__1__11, 
         que_out_23__1__10, que_out_23__1__9, que_out_23__1__8, que_out_23__1__7, 
         que_out_23__1__6, que_out_23__1__5, que_out_23__1__4, que_out_23__1__3, 
         que_out_23__1__2, que_out_23__1__1, que_out_23__1__0, que_out_23__2__15, 
         que_out_23__2__14, que_out_23__2__13, que_out_23__2__12, 
         que_out_23__2__11, que_out_23__2__10, que_out_23__2__9, 
         que_out_23__2__8, que_out_23__2__7, que_out_23__2__6, que_out_23__2__5, 
         que_out_23__2__4, que_out_23__2__3, que_out_23__2__2, que_out_23__2__1, 
         que_out_23__2__0, que_out_23__3__15, que_out_23__3__14, 
         que_out_23__3__13, que_out_23__3__12, que_out_23__3__11, 
         que_out_23__3__10, que_out_23__3__9, que_out_23__3__8, que_out_23__3__7, 
         que_out_23__3__6, que_out_23__3__5, que_out_23__3__4, que_out_23__3__3, 
         que_out_23__3__2, que_out_23__3__1, que_out_23__3__0, que_out_23__4__15, 
         que_out_23__4__14, que_out_23__4__13, que_out_23__4__12, 
         que_out_23__4__11, que_out_23__4__10, que_out_23__4__9, 
         que_out_23__4__8, que_out_23__4__7, que_out_23__4__6, que_out_23__4__5, 
         que_out_23__4__4, que_out_23__4__3, que_out_23__4__2, que_out_23__4__1, 
         que_out_23__4__0, que_out_24__0__15, que_out_24__0__14, 
         que_out_24__0__13, que_out_24__0__12, que_out_24__0__11, 
         que_out_24__0__10, que_out_24__0__9, que_out_24__0__8, que_out_24__0__7, 
         que_out_24__0__6, que_out_24__0__5, que_out_24__0__4, que_out_24__0__3, 
         que_out_24__0__2, que_out_24__0__1, que_out_24__0__0, que_out_24__1__15, 
         que_out_24__1__14, que_out_24__1__13, que_out_24__1__12, 
         que_out_24__1__11, que_out_24__1__10, que_out_24__1__9, 
         que_out_24__1__8, que_out_24__1__7, que_out_24__1__6, que_out_24__1__5, 
         que_out_24__1__4, que_out_24__1__3, que_out_24__1__2, que_out_24__1__1, 
         que_out_24__1__0, que_out_24__2__15, que_out_24__2__14, 
         que_out_24__2__13, que_out_24__2__12, que_out_24__2__11, 
         que_out_24__2__10, que_out_24__2__9, que_out_24__2__8, que_out_24__2__7, 
         que_out_24__2__6, que_out_24__2__5, que_out_24__2__4, que_out_24__2__3, 
         que_out_24__2__2, que_out_24__2__1, que_out_24__2__0, que_out_24__3__15, 
         que_out_24__3__14, que_out_24__3__13, que_out_24__3__12, 
         que_out_24__3__11, que_out_24__3__10, que_out_24__3__9, 
         que_out_24__3__8, que_out_24__3__7, que_out_24__3__6, que_out_24__3__5, 
         que_out_24__3__4, que_out_24__3__3, que_out_24__3__2, que_out_24__3__1, 
         que_out_24__3__0, que_out_24__4__15, que_out_24__4__14, 
         que_out_24__4__13, que_out_24__4__12, que_out_24__4__11, 
         que_out_24__4__10, que_out_24__4__9, que_out_24__4__8, que_out_24__4__7, 
         que_out_24__4__6, que_out_24__4__5, que_out_24__4__4, que_out_24__4__3, 
         que_out_24__4__2, que_out_24__4__1, que_out_24__4__0, que_out_25__0__15, 
         que_out_25__0__14, que_out_25__0__13, que_out_25__0__12, 
         que_out_25__0__11, que_out_25__0__10, que_out_25__0__9, 
         que_out_25__0__8, que_out_25__0__7, que_out_25__0__6, que_out_25__0__5, 
         que_out_25__0__4, que_out_25__0__3, que_out_25__0__2, que_out_25__0__1, 
         que_out_25__0__0, que_out_25__1__15, que_out_25__1__14, 
         que_out_25__1__13, que_out_25__1__12, que_out_25__1__11, 
         que_out_25__1__10, que_out_25__1__9, que_out_25__1__8, que_out_25__1__7, 
         que_out_25__1__6, que_out_25__1__5, que_out_25__1__4, que_out_25__1__3, 
         que_out_25__1__2, que_out_25__1__1, que_out_25__1__0, que_out_25__2__15, 
         que_out_25__2__14, que_out_25__2__13, que_out_25__2__12, 
         que_out_25__2__11, que_out_25__2__10, que_out_25__2__9, 
         que_out_25__2__8, que_out_25__2__7, que_out_25__2__6, que_out_25__2__5, 
         que_out_25__2__4, que_out_25__2__3, que_out_25__2__2, que_out_25__2__1, 
         que_out_25__2__0, que_out_25__3__15, que_out_25__3__14, 
         que_out_25__3__13, que_out_25__3__12, que_out_25__3__11, 
         que_out_25__3__10, que_out_25__3__9, que_out_25__3__8, que_out_25__3__7, 
         que_out_25__3__6, que_out_25__3__5, que_out_25__3__4, que_out_25__3__3, 
         que_out_25__3__2, que_out_25__3__1, que_out_25__3__0, que_out_25__4__15, 
         que_out_25__4__14, que_out_25__4__13, que_out_25__4__12, 
         que_out_25__4__11, que_out_25__4__10, que_out_25__4__9, 
         que_out_25__4__8, que_out_25__4__7, que_out_25__4__6, que_out_25__4__5, 
         que_out_25__4__4, que_out_25__4__3, que_out_25__4__2, que_out_25__4__1, 
         que_out_25__4__0, que_out_26__0__15, que_out_26__0__14, 
         que_out_26__0__13, que_out_26__0__12, que_out_26__0__11, 
         que_out_26__0__10, que_out_26__0__9, que_out_26__0__8, que_out_26__0__7, 
         que_out_26__0__6, que_out_26__0__5, que_out_26__0__4, que_out_26__0__3, 
         que_out_26__0__2, que_out_26__0__1, que_out_26__0__0, que_out_26__1__15, 
         que_out_26__1__14, que_out_26__1__13, que_out_26__1__12, 
         que_out_26__1__11, que_out_26__1__10, que_out_26__1__9, 
         que_out_26__1__8, que_out_26__1__7, que_out_26__1__6, que_out_26__1__5, 
         que_out_26__1__4, que_out_26__1__3, que_out_26__1__2, que_out_26__1__1, 
         que_out_26__1__0, que_out_26__2__15, que_out_26__2__14, 
         que_out_26__2__13, que_out_26__2__12, que_out_26__2__11, 
         que_out_26__2__10, que_out_26__2__9, que_out_26__2__8, que_out_26__2__7, 
         que_out_26__2__6, que_out_26__2__5, que_out_26__2__4, que_out_26__2__3, 
         que_out_26__2__2, que_out_26__2__1, que_out_26__2__0, que_out_26__3__15, 
         que_out_26__3__14, que_out_26__3__13, que_out_26__3__12, 
         que_out_26__3__11, que_out_26__3__10, que_out_26__3__9, 
         que_out_26__3__8, que_out_26__3__7, que_out_26__3__6, que_out_26__3__5, 
         que_out_26__3__4, que_out_26__3__3, que_out_26__3__2, que_out_26__3__1, 
         que_out_26__3__0, que_out_26__4__15, que_out_26__4__14, 
         que_out_26__4__13, que_out_26__4__12, que_out_26__4__11, 
         que_out_26__4__10, que_out_26__4__9, que_out_26__4__8, que_out_26__4__7, 
         que_out_26__4__6, que_out_26__4__5, que_out_26__4__4, que_out_26__4__3, 
         que_out_26__4__2, que_out_26__4__1, que_out_26__4__0, que_out_27__0__15, 
         que_out_27__0__14, que_out_27__0__13, que_out_27__0__12, 
         que_out_27__0__11, que_out_27__0__10, que_out_27__0__9, 
         que_out_27__0__8, que_out_27__0__7, que_out_27__0__6, que_out_27__0__5, 
         que_out_27__0__4, que_out_27__0__3, que_out_27__0__2, que_out_27__0__1, 
         que_out_27__0__0, que_out_27__1__15, que_out_27__1__14, 
         que_out_27__1__13, que_out_27__1__12, que_out_27__1__11, 
         que_out_27__1__10, que_out_27__1__9, que_out_27__1__8, que_out_27__1__7, 
         que_out_27__1__6, que_out_27__1__5, que_out_27__1__4, que_out_27__1__3, 
         que_out_27__1__2, que_out_27__1__1, que_out_27__1__0, que_out_27__2__15, 
         que_out_27__2__14, que_out_27__2__13, que_out_27__2__12, 
         que_out_27__2__11, que_out_27__2__10, que_out_27__2__9, 
         que_out_27__2__8, que_out_27__2__7, que_out_27__2__6, que_out_27__2__5, 
         que_out_27__2__4, que_out_27__2__3, que_out_27__2__2, que_out_27__2__1, 
         que_out_27__2__0, que_out_27__3__15, que_out_27__3__14, 
         que_out_27__3__13, que_out_27__3__12, que_out_27__3__11, 
         que_out_27__3__10, que_out_27__3__9, que_out_27__3__8, que_out_27__3__7, 
         que_out_27__3__6, que_out_27__3__5, que_out_27__3__4, que_out_27__3__3, 
         que_out_27__3__2, que_out_27__3__1, que_out_27__3__0, que_out_27__4__15, 
         que_out_27__4__14, que_out_27__4__13, que_out_27__4__12, 
         que_out_27__4__11, que_out_27__4__10, que_out_27__4__9, 
         que_out_27__4__8, que_out_27__4__7, que_out_27__4__6, que_out_27__4__5, 
         que_out_27__4__4, que_out_27__4__3, que_out_27__4__2, que_out_27__4__1, 
         que_out_27__4__0, sel_que_27, sel_que_26, sel_que_25, sel_que_24, 
         sel_que_23, sel_que_22, sel_que_21, sel_que_20, sel_que_19, sel_que_18, 
         sel_que_17, sel_que_16, sel_que_15, sel_que_14, sel_que_13, sel_que_12, 
         sel_que_11, sel_que_10, sel_que_9, sel_que_8, sel_que_7, sel_que_6, 
         sel_que_5, sel_que_4, sel_que_3, sel_que_2, sel_que_1, sel_que_0, nx12, 
         nx14, nx28, nx30, nx42, nx48, nx62, nx64, nx68, nx74, nx82, nx88, nx90, 
         nx94, nx100, nx104, nx114, nx118, nx122, nx130, nx136, nx144, nx150, 
         nx158, nx166, nx172, nx180, nx188, nx192, nx200, nx206, nx214, nx222, 
         nx226, nx230, nx238, nx268, nx294, nx322, nx348, nx378, nx404, nx432, 
         nx458, nx488, nx514, nx542, nx568, nx598, nx624, nx652, nx678, nx708, 
         nx734, nx762, nx788, nx818, nx844, nx872, nx898, nx928, nx954, nx982, 
         nx1008, nx1038, nx1064, nx1092, nx1118, nx1148, nx1174, nx1202, nx1228, 
         nx1258, nx1284, nx1312, nx1338, nx1368, nx1394, nx1422, nx1448, nx1478, 
         nx1504, nx1532, nx1558, nx1588, nx1614, nx1642, nx1668, nx1698, nx1724, 
         nx1752, nx1778, nx1808, nx1834, nx1862, nx1888, nx1918, nx1944, nx1972, 
         nx1998, nx2028, nx2054, nx2082, nx2108, nx2138, nx2164, nx2192, nx2218, 
         nx2248, nx2274, nx2302, nx2328, nx2358, nx2384, nx2412, nx2438, nx2468, 
         nx2494, nx2522, nx2548, nx2578, nx2604, nx2632, nx2658, nx2688, nx2714, 
         nx2742, nx2768, nx2798, nx2824, nx2852, nx2878, nx2908, nx2934, nx2962, 
         nx2988, nx3018, nx3044, nx3072, nx3098, nx3128, nx3154, nx3182, nx3208, 
         nx3238, nx3264, nx3292, nx3318, nx3348, nx3374, nx3402, nx3428, nx3458, 
         nx3484, nx3512, nx3538, nx3568, nx3594, nx3622, nx3648, nx3678, nx3704, 
         nx3732, nx3758, nx3788, nx3814, nx3842, nx3868, nx3898, nx3924, nx3952, 
         nx3978, nx4008, nx4034, nx4062, nx4088, nx4118, nx4144, nx4172, nx4198, 
         nx4228, nx4254, nx4282, nx4308, nx4338, nx4364, nx4392, nx4418, nx4448, 
         nx4474, nx4502, nx4528, nx4558, nx4584, nx4612, nx4638, nx4668, nx4694, 
         nx4722, nx4748, nx4778, nx4804, nx4832, nx4858, nx4888, nx4914, nx4942, 
         nx4968, nx4998, nx5024, nx5052, nx5078, nx5108, nx5134, nx5162, nx5188, 
         nx5218, nx5244, nx5272, nx5298, nx5328, nx5354, nx5382, nx5408, nx5438, 
         nx5464, nx5492, nx5518, nx5548, nx5574, nx5602, nx5628, nx5658, nx5684, 
         nx5712, nx5738, nx5768, nx5794, nx5822, nx5848, nx5878, nx5904, nx5932, 
         nx5958, nx5988, nx6014, nx6042, nx6068, nx6098, nx6124, nx6152, nx6178, 
         nx6208, nx6234, nx6262, nx6288, nx6318, nx6344, nx6372, nx6398, nx6428, 
         nx6454, nx6482, nx6508, nx6538, nx6564, nx6592, nx6618, nx6648, nx6674, 
         nx6702, nx6728, nx6758, nx6784, nx6812, nx6838, nx6868, nx6894, nx6922, 
         nx6948, nx6978, nx7004, nx7032, nx7058, nx7088, nx7114, nx7142, nx7168, 
         nx7198, nx7224, nx7252, nx7278, nx7308, nx7334, nx7362, nx7388, nx7418, 
         nx7444, nx7472, nx7498, nx7528, nx7554, nx7582, nx7608, nx7638, nx7664, 
         nx7692, nx7718, nx7748, nx7774, nx7802, nx7828, nx7858, nx7884, nx7912, 
         nx7938, nx7968, nx7994, nx8022, nx8048, nx8078, nx8104, nx8132, nx8158, 
         nx8188, nx8214, nx8242, nx8268, nx8298, nx8324, nx8352, nx8378, nx8408, 
         nx8434, nx8462, nx8488, nx8518, nx8544, nx8572, nx8598, nx8628, nx8654, 
         nx8682, nx8708, nx8738, nx8764, nx8792, nx8818, nx8848, nx8874, nx8902, 
         nx8928, nx8938, nx9038, nx6829, nx6833, nx6835, nx6839, nx6843, nx6847, 
         nx6875, nx6885, nx6889, nx6893, nx6897, nx6901, nx6905, nx6915, nx6927, 
         nx6931, nx6933, nx6937, nx6939, nx6943, nx6945, nx6949, nx6951, nx6955, 
         nx6957, nx6961, nx6965, nx6967, nx6971, nx6977, nx6985, nx6991, nx6999, 
         nx7007, nx7017, nx7029, nx7037, nx7043, nx7053, nx7055, nx7057, nx7061, 
         nx7063, nx7065, nx7069, nx7071, nx7073, nx7077, nx7079, nx7081, nx7087, 
         nx7089, nx7091, nx7095, nx7097, nx7099, nx7103, nx7105, nx7107, nx7111, 
         nx7113, nx7115, nx7121, nx7123, nx7125, nx7129, nx7131, nx7133, nx7137, 
         nx7139, nx7141, nx7145, nx7147, nx7149, nx7155, nx7157, nx7159, nx7163, 
         nx7165, nx7167, nx7171, nx7173, nx7175, nx7179, nx7181, nx7183, nx7189, 
         nx7191, nx7193, nx7197, nx7199, nx7201, nx7205, nx7207, nx7209, nx7213, 
         nx7215, nx7217, nx7223, nx7225, nx7227, nx7231, nx7233, nx7235, nx7239, 
         nx7241, nx7243, nx7247, nx7249, nx7251, nx7257, nx7259, nx7261, nx7265, 
         nx7267, nx7269, nx7273, nx7275, nx7277, nx7281, nx7283, nx7285, nx7291, 
         nx7293, nx7295, nx7299, nx7301, nx7303, nx7307, nx7309, nx7311, nx7315, 
         nx7317, nx7319, nx7325, nx7327, nx7329, nx7333, nx7335, nx7337, nx7341, 
         nx7343, nx7345, nx7349, nx7351, nx7353, nx7359, nx7361, nx7363, nx7367, 
         nx7369, nx7371, nx7375, nx7377, nx7379, nx7383, nx7385, nx7387, nx7393, 
         nx7395, nx7397, nx7401, nx7403, nx7405, nx7409, nx7411, nx7413, nx7417, 
         nx7419, nx7421, nx7427, nx7429, nx7431, nx7435, nx7437, nx7439, nx7443, 
         nx7445, nx7447, nx7451, nx7453, nx7455, nx7461, nx7463, nx7465, nx7469, 
         nx7471, nx7473, nx7477, nx7479, nx7481, nx7485, nx7487, nx7489, nx7495, 
         nx7497, nx7499, nx7503, nx7505, nx7507, nx7511, nx7513, nx7515, nx7519, 
         nx7521, nx7523, nx7529, nx7531, nx7533, nx7537, nx7539, nx7541, nx7545, 
         nx7547, nx7549, nx7553, nx7555, nx7557, nx7563, nx7565, nx7567, nx7571, 
         nx7573, nx7575, nx7579, nx7581, nx7583, nx7587, nx7589, nx7591, nx7597, 
         nx7599, nx7601, nx7605, nx7607, nx7609, nx7613, nx7615, nx7617, nx7621, 
         nx7623, nx7625, nx7631, nx7633, nx7635, nx7639, nx7641, nx7643, nx7647, 
         nx7649, nx7651, nx7655, nx7657, nx7659, nx7665, nx7667, nx7669, nx7673, 
         nx7675, nx7677, nx7681, nx7683, nx7685, nx7689, nx7691, nx7693, nx7699, 
         nx7701, nx7703, nx7707, nx7709, nx7711, nx7715, nx7717, nx7719, nx7723, 
         nx7725, nx7727, nx7733, nx7735, nx7737, nx7741, nx7743, nx7745, nx7749, 
         nx7751, nx7753, nx7757, nx7759, nx7761, nx7767, nx7769, nx7771, nx7775, 
         nx7777, nx7779, nx7783, nx7785, nx7787, nx7791, nx7793, nx7795, nx7801, 
         nx7803, nx7805, nx7809, nx7811, nx7813, nx7817, nx7819, nx7821, nx7825, 
         nx7827, nx7829, nx7835, nx7837, nx7839, nx7843, nx7845, nx7847, nx7851, 
         nx7853, nx7855, nx7859, nx7861, nx7863, nx7869, nx7871, nx7873, nx7877, 
         nx7879, nx7881, nx7885, nx7887, nx7889, nx7893, nx7895, nx7897, nx7903, 
         nx7905, nx7907, nx7911, nx7913, nx7915, nx7919, nx7921, nx7923, nx7927, 
         nx7929, nx7931, nx7937, nx7939, nx7941, nx7945, nx7947, nx7949, nx7953, 
         nx7955, nx7957, nx7961, nx7963, nx7965, nx7971, nx7973, nx7975, nx7979, 
         nx7981, nx7983, nx7987, nx7989, nx7991, nx7995, nx7997, nx7999, nx8005, 
         nx8007, nx8009, nx8013, nx8015, nx8017, nx8021, nx8023, nx8025, nx8029, 
         nx8031, nx8033, nx8039, nx8041, nx8043, nx8047, nx8049, nx8051, nx8055, 
         nx8057, nx8059, nx8063, nx8065, nx8067, nx8073, nx8075, nx8077, nx8081, 
         nx8083, nx8085, nx8089, nx8091, nx8093, nx8097, nx8099, nx8101, nx8107, 
         nx8109, nx8111, nx8115, nx8117, nx8119, nx8123, nx8125, nx8127, nx8131, 
         nx8133, nx8135, nx8141, nx8143, nx8145, nx8149, nx8151, nx8153, nx8157, 
         nx8159, nx8161, nx8165, nx8167, nx8169, nx8175, nx8177, nx8179, nx8183, 
         nx8185, nx8187, nx8191, nx8193, nx8195, nx8199, nx8201, nx8203, nx8209, 
         nx8211, nx8213, nx8217, nx8219, nx8221, nx8225, nx8227, nx8229, nx8233, 
         nx8235, nx8237, nx8243, nx8245, nx8247, nx8251, nx8253, nx8255, nx8259, 
         nx8261, nx8263, nx8267, nx8269, nx8271, nx8277, nx8279, nx8281, nx8285, 
         nx8287, nx8289, nx8293, nx8295, nx8297, nx8301, nx8303, nx8305, nx8311, 
         nx8313, nx8315, nx8319, nx8321, nx8323, nx8327, nx8329, nx8331, nx8335, 
         nx8337, nx8339, nx8345, nx8347, nx8349, nx8353, nx8355, nx8357, nx8361, 
         nx8363, nx8365, nx8369, nx8371, nx8373, nx8379, nx8381, nx8383, nx8387, 
         nx8389, nx8391, nx8395, nx8397, nx8399, nx8403, nx8405, nx8407, nx8413, 
         nx8415, nx8417, nx8421, nx8423, nx8425, nx8429, nx8431, nx8433, nx8437, 
         nx8439, nx8441, nx8447, nx8449, nx8451, nx8455, nx8457, nx8459, nx8463, 
         nx8465, nx8467, nx8471, nx8473, nx8475, nx8481, nx8483, nx8485, nx8489, 
         nx8491, nx8493, nx8497, nx8499, nx8501, nx8505, nx8507, nx8509, nx8515, 
         nx8517, nx8519, nx8523, nx8525, nx8527, nx8531, nx8533, nx8535, nx8539, 
         nx8541, nx8543, nx8549, nx8551, nx8553, nx8557, nx8559, nx8561, nx8565, 
         nx8567, nx8569, nx8573, nx8575, nx8577, nx8583, nx8585, nx8587, nx8591, 
         nx8593, nx8595, nx8599, nx8601, nx8603, nx8607, nx8609, nx8611, nx8617, 
         nx8619, nx8621, nx8625, nx8627, nx8629, nx8633, nx8635, nx8637, nx8641, 
         nx8643, nx8645, nx8651, nx8653, nx8655, nx8659, nx8661, nx8663, nx8667, 
         nx8669, nx8671, nx8675, nx8677, nx8679, nx8685, nx8687, nx8689, nx8693, 
         nx8695, nx8697, nx8701, nx8703, nx8705, nx8709, nx8711, nx8713, nx8719, 
         nx8721, nx8723, nx8727, nx8729, nx8731, nx8735, nx8737, nx8739, nx8743, 
         nx8745, nx8747, nx8753, nx8755, nx8757, nx8761, nx8763, nx8765, nx8769, 
         nx8771, nx8773, nx8777, nx8779, nx8781, nx8787, nx8789, nx8791, nx8795, 
         nx8797, nx8799, nx8803, nx8805, nx8807, nx8811, nx8813, nx8815, nx8821, 
         nx8823, nx8825, nx8829, nx8831, nx8833, nx8837, nx8839, nx8841, nx8845, 
         nx8847, nx8849, nx8855, nx8857, nx8859, nx8863, nx8865, nx8867, nx8871, 
         nx8873, nx8875, nx8879, nx8881, nx8883, nx8889, nx8891, nx8893, nx8897, 
         nx8899, nx8901, nx8905, nx8907, nx8909, nx8913, nx8915, nx8917, nx8923, 
         nx8925, nx8927, nx8931, nx8933, nx8935, nx8939, nx8941, nx8943, nx8947, 
         nx8949, nx8951, nx8955, nx8957, nx8959, nx8963, nx8965, nx8967, nx8970, 
         nx8973, nx8975, nx8978, nx8981, nx8983, nx8989, nx8991, nx8993, nx8997, 
         nx8999, nx9001, nx9005, nx9007, nx9009, nx9013, nx9015, nx9017, nx9023, 
         nx9025, nx9027, nx9031, nx9033, nx9035, nx9039, nx9041, nx9043, nx9047, 
         nx9049, nx9051, nx9057, nx9059, nx9061, nx9065, nx9067, nx9069, nx9073, 
         nx9075, nx9077, nx9081, nx9083, nx9085, nx9090, nx9093, nx9095, nx9098, 
         nx9101, nx9103, nx9106, nx9108, nx9110, nx9113, nx9115, nx9117, nx9121, 
         nx9123, nx9125, nx9128, nx9130, nx9132, nx9135, nx9137, nx9139, nx9142, 
         nx9144, nx9146, nx9150, nx9152, nx9154, nx9157, nx9159, nx9161, nx9164, 
         nx9166, nx9168, nx9171, nx9173, nx9175, nx9179, nx9181, nx9183, nx9186, 
         nx9188, nx9190, nx9193, nx9195, nx9197, nx9200, nx9202, nx9204, nx9208, 
         nx9210, nx9212, nx9215, nx9217, nx9219, nx9222, nx9224, nx9226, nx9229, 
         nx9231, nx9233, nx9237, nx9239, nx9241, nx9244, nx9246, nx9248, nx9251, 
         nx9253, nx9255, nx9258, nx9260, nx9262, nx9266, nx9268, nx9270, nx9273, 
         nx9275, nx9277, nx9280, nx9282, nx9284, nx9287, nx9289, nx9291, nx9295, 
         nx9297, nx9299, nx9302, nx9304, nx9306, nx9309, nx9311, nx9313, nx9316, 
         nx9318, nx9320, nx9324, nx9326, nx9328, nx9331, nx9333, nx9335, nx9338, 
         nx9340, nx9342, nx9345, nx9347, nx9349, nx9353, nx9355, nx9357, nx9360, 
         nx9362, nx9364, nx9367, nx9369, nx9371, nx9374, nx9376, nx9378, nx9382, 
         nx9384, nx9386, nx9389, nx9391, nx9393, nx9396, nx9398, nx9400, nx9403, 
         nx9405, nx9407, nx9411, nx9413, nx9415, nx9418, nx9420, nx9422, nx9425, 
         nx9427, nx9429, nx9432, nx9434, nx9436, nx9440, nx9442, nx9444, nx9447, 
         nx9449, nx9451, nx9454, nx9456, nx9458, nx9461, nx9463, nx9465, nx9469, 
         nx9471, nx9473, nx9476, nx9478, nx9480, nx9483, nx9485, nx9487, nx9490, 
         nx9492, nx9494, nx9498, nx9500, nx9502, nx9505, nx9507, nx9509, nx9512, 
         nx9514, nx9516, nx9519, nx9521, nx9523, nx9527, nx9529, nx9531, nx9534, 
         nx9536, nx9538, nx9541, nx9543, nx9545, nx9548, nx9550, nx9552, nx9556, 
         nx9558, nx9560, nx9563, nx9565, nx9567, nx9570, nx9572, nx9574, nx9577, 
         nx9579, nx9581, nx9585, nx9587, nx9589, nx9592, nx9594, nx9596, nx9599, 
         nx9601, nx9603, nx9606, nx9608, nx9610, nx9614, nx9616, nx9618, nx9621, 
         nx9623, nx9625, nx9628, nx9630, nx9632, nx9635, nx9637, nx9639, nx9648, 
         nx9650, nx9652, nx9654, nx9656, nx9658, nx9660, nx9662, nx9664, nx9666, 
         nx9668, nx9670, nx9674, nx9676, nx9678, nx9680, nx9682, nx9684, nx9686, 
         nx9688, nx9690, nx9692, nx9694, nx9696, nx9700, nx9702, nx9704, nx9706, 
         nx9708, nx9710, nx9712, nx9714, nx9716, nx9718, nx9720, nx9722, nx9726, 
         nx9728, nx9730, nx9732, nx9734, nx9736, nx9738, nx9740, nx9742, nx9744, 
         nx9746, nx9748, nx9752, nx9754, nx9756, nx9758, nx9760, nx9762, nx9764, 
         nx9766, nx9768, nx9770, nx9772, nx9774, nx9778, nx9780, nx9782, nx9784, 
         nx9786, nx9788, nx9790, nx9792, nx9794, nx9796, nx9798, nx9800, nx9804, 
         nx9806, nx9808, nx9810, nx9812, nx9814, nx9816, nx9818, nx9820, nx9822, 
         nx9824, nx9826, nx9830, nx9832, nx9834, nx9836, nx9838, nx9840, nx9842, 
         nx9844, nx9846, nx9848, nx9850, nx9852, nx9856, nx9858, nx9860, nx9862, 
         nx9864, nx9866, nx9868, nx9870, nx9872, nx9874, nx9876, nx9878, nx9882, 
         nx9884, nx9886, nx9888, nx9890, nx9892, nx9894, nx9896, nx9898, nx9900, 
         nx9902, nx9904, nx9908, nx9910, nx9912, nx9914, nx9916, nx9918, nx9920, 
         nx9922, nx9924, nx9926, nx9928, nx9930, nx9934, nx9936, nx9938, nx9940, 
         nx9942, nx9944, nx9946, nx9948, nx9950, nx9952, nx9954, nx9956, nx9960, 
         nx9962, nx9964, nx9966, nx9968, nx9970, nx9972, nx9974, nx9976, nx9978, 
         nx9980, nx9982, nx9986, nx9988, nx9990, nx9992, nx9994, nx9996, nx9998, 
         nx10000, nx10002, nx10004, nx10006, nx10008, nx10012, nx10014, nx10016, 
         nx10018, nx10020, nx10022, nx10024, nx10026, nx10028, nx10030, nx10032, 
         nx10034, nx10038, nx10040, nx10042, nx10044, nx10046, nx10048, nx10050, 
         nx10052, nx10054, nx10056, nx10058, nx10060, nx10064, nx10066, nx10068, 
         nx10070, nx10072, nx10074, nx10076, nx10078, nx10080, nx10082, nx10084, 
         nx10086, nx10090, nx10092, nx10094, nx10096, nx10098, nx10100, nx10102, 
         nx10104, nx10106, nx10108, nx10110, nx10112, nx10116, nx10118, nx10120, 
         nx10122, nx10124, nx10126, nx10128, nx10130, nx10132, nx10134, nx10136, 
         nx10138, nx10142, nx10144, nx10146, nx10148, nx10150, nx10152, nx10154, 
         nx10156, nx10158, nx10160, nx10162, nx10164, nx10168, nx10170, nx10172, 
         nx10174, nx10176, nx10178, nx10180, nx10182, nx10184, nx10186, nx10188, 
         nx10190, nx10194, nx10196, nx10198, nx10200, nx10202, nx10204, nx10206, 
         nx10208, nx10210, nx10212, nx10214, nx10216, nx10220, nx10222, nx10224, 
         nx10226, nx10228, nx10230, nx10232, nx10234, nx10236, nx10238, nx10240, 
         nx10242, nx10246, nx10248, nx10250, nx10252, nx10254, nx10256, nx10258, 
         nx10260, nx10262, nx10264, nx10266, nx10268, nx10272, nx10274, nx10276, 
         nx10278, nx10280, nx10282, nx10284, nx10286, nx10288, nx10290, nx10292, 
         nx10294, nx10298, nx10300, nx10302, nx10304, nx10306, nx10308, nx10310, 
         nx10312, nx10314, nx10316, nx10318, nx10320, nx10324, nx10326, nx10328, 
         nx10330, nx10332, nx10334, nx10336, nx10338, nx10340, nx10342, nx10344, 
         nx10346, nx10350, nx10352, nx10354, nx10356, nx10358, nx10360, nx10362, 
         nx10364, nx10366, nx10368, nx10370, nx10372, nx10374, nx10376, nx10378, 
         nx10380, nx10382, nx10384, nx10386, nx10388, nx10390, nx10392, nx10394, 
         nx10396, nx10398, nx10400, nx10402, nx10404, nx10406, nx10408, nx10410, 
         nx10412, nx10414, nx10416, nx10418, nx10420, nx10422, nx10424, nx10426, 
         nx10428, nx10430, nx10432, nx10434, nx10436, nx10438, nx10440, nx10442, 
         nx10444, nx10446, nx10448, nx10450, nx10452, nx10454, nx10456, nx10458, 
         nx10460, nx10462, nx10464, nx10466, nx10468, nx10470, nx10472, nx10474, 
         nx10476, nx10478, nx10480, nx10482, nx10484, nx10486, nx10488, nx10494, 
         nx10496, nx10498, nx10500, nx10502, nx10504, nx10506, nx10508, nx10510, 
         nx10512, nx10514, nx10516, nx10518, nx10520, nx10522, nx10524, nx10526, 
         nx10528, nx10530, nx10532, nx10534, nx10536, nx10538, nx10540, nx10542, 
         nx10544, nx10546, nx10548, nx10550, nx10552, nx10554, nx10556, nx10558, 
         nx10560, nx10562, nx10564, nx10566, nx10568, nx10570, nx10572, nx10574, 
         nx10576, nx10578, nx10580, nx10582, nx10584, nx10586, nx10588, nx10590, 
         nx10592, nx10594, nx10596, nx10598, nx10600, nx10602, nx10604, nx10606, 
         nx10608, nx10610, nx10612, nx10614, nx10616, nx10618, nx10620, nx10622, 
         nx10624, nx10626, nx10628, nx10630, nx10632, nx10634, nx10636, nx10638, 
         nx10640, nx10642, nx10644, nx10646, nx10648, nx10650, nx10652, nx10654, 
         nx10656, nx10658, nx10660, nx10662, nx10664, nx10666, nx10668, nx10690, 
         nx10692, nx10694, nx10696, nx10698, nx10700, nx10702, nx10704, nx10706, 
         nx10708, nx10710, nx10712, nx10714, nx10716, nx10718, nx10720, nx10722, 
         nx10724, nx10726, nx10728, nx10730, nx10732, nx10734, nx10736, nx10742, 
         nx10744, nx10746, nx10748;



    Queue_5 gen_queues_0_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_0__0__15), .q_0__14 (
            que_out_0__0__14), .q_0__13 (que_out_0__0__13), .q_0__12 (
            que_out_0__0__12), .q_0__11 (que_out_0__0__11), .q_0__10 (
            que_out_0__0__10), .q_0__9 (que_out_0__0__9), .q_0__8 (
            que_out_0__0__8), .q_0__7 (que_out_0__0__7), .q_0__6 (
            que_out_0__0__6), .q_0__5 (que_out_0__0__5), .q_0__4 (
            que_out_0__0__4), .q_0__3 (que_out_0__0__3), .q_0__2 (
            que_out_0__0__2), .q_0__1 (que_out_0__0__1), .q_0__0 (
            que_out_0__0__0), .q_1__15 (que_out_0__1__15), .q_1__14 (
            que_out_0__1__14), .q_1__13 (que_out_0__1__13), .q_1__12 (
            que_out_0__1__12), .q_1__11 (que_out_0__1__11), .q_1__10 (
            que_out_0__1__10), .q_1__9 (que_out_0__1__9), .q_1__8 (
            que_out_0__1__8), .q_1__7 (que_out_0__1__7), .q_1__6 (
            que_out_0__1__6), .q_1__5 (que_out_0__1__5), .q_1__4 (
            que_out_0__1__4), .q_1__3 (que_out_0__1__3), .q_1__2 (
            que_out_0__1__2), .q_1__1 (que_out_0__1__1), .q_1__0 (
            que_out_0__1__0), .q_2__15 (que_out_0__2__15), .q_2__14 (
            que_out_0__2__14), .q_2__13 (que_out_0__2__13), .q_2__12 (
            que_out_0__2__12), .q_2__11 (que_out_0__2__11), .q_2__10 (
            que_out_0__2__10), .q_2__9 (que_out_0__2__9), .q_2__8 (
            que_out_0__2__8), .q_2__7 (que_out_0__2__7), .q_2__6 (
            que_out_0__2__6), .q_2__5 (que_out_0__2__5), .q_2__4 (
            que_out_0__2__4), .q_2__3 (que_out_0__2__3), .q_2__2 (
            que_out_0__2__2), .q_2__1 (que_out_0__2__1), .q_2__0 (
            que_out_0__2__0), .q_3__15 (que_out_0__3__15), .q_3__14 (
            que_out_0__3__14), .q_3__13 (que_out_0__3__13), .q_3__12 (
            que_out_0__3__12), .q_3__11 (que_out_0__3__11), .q_3__10 (
            que_out_0__3__10), .q_3__9 (que_out_0__3__9), .q_3__8 (
            que_out_0__3__8), .q_3__7 (que_out_0__3__7), .q_3__6 (
            que_out_0__3__6), .q_3__5 (que_out_0__3__5), .q_3__4 (
            que_out_0__3__4), .q_3__3 (que_out_0__3__3), .q_3__2 (
            que_out_0__3__2), .q_3__1 (que_out_0__3__1), .q_3__0 (
            que_out_0__3__0), .q_4__15 (que_out_0__4__15), .q_4__14 (
            que_out_0__4__14), .q_4__13 (que_out_0__4__13), .q_4__12 (
            que_out_0__4__12), .q_4__11 (que_out_0__4__11), .q_4__10 (
            que_out_0__4__10), .q_4__9 (que_out_0__4__9), .q_4__8 (
            que_out_0__4__8), .q_4__7 (que_out_0__4__7), .q_4__6 (
            que_out_0__4__6), .q_4__5 (que_out_0__4__5), .q_4__4 (
            que_out_0__4__4), .q_4__3 (que_out_0__4__3), .q_4__2 (
            que_out_0__4__2), .q_4__1 (que_out_0__4__1), .q_4__0 (
            que_out_0__4__0), .clk (nx10714), .load (sel_que_0), .reset (nx10690
            )) ;
    Queue_5 gen_queues_1_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_1__0__15), .q_0__14 (
            que_out_1__0__14), .q_0__13 (que_out_1__0__13), .q_0__12 (
            que_out_1__0__12), .q_0__11 (que_out_1__0__11), .q_0__10 (
            que_out_1__0__10), .q_0__9 (que_out_1__0__9), .q_0__8 (
            que_out_1__0__8), .q_0__7 (que_out_1__0__7), .q_0__6 (
            que_out_1__0__6), .q_0__5 (que_out_1__0__5), .q_0__4 (
            que_out_1__0__4), .q_0__3 (que_out_1__0__3), .q_0__2 (
            que_out_1__0__2), .q_0__1 (que_out_1__0__1), .q_0__0 (
            que_out_1__0__0), .q_1__15 (que_out_1__1__15), .q_1__14 (
            que_out_1__1__14), .q_1__13 (que_out_1__1__13), .q_1__12 (
            que_out_1__1__12), .q_1__11 (que_out_1__1__11), .q_1__10 (
            que_out_1__1__10), .q_1__9 (que_out_1__1__9), .q_1__8 (
            que_out_1__1__8), .q_1__7 (que_out_1__1__7), .q_1__6 (
            que_out_1__1__6), .q_1__5 (que_out_1__1__5), .q_1__4 (
            que_out_1__1__4), .q_1__3 (que_out_1__1__3), .q_1__2 (
            que_out_1__1__2), .q_1__1 (que_out_1__1__1), .q_1__0 (
            que_out_1__1__0), .q_2__15 (que_out_1__2__15), .q_2__14 (
            que_out_1__2__14), .q_2__13 (que_out_1__2__13), .q_2__12 (
            que_out_1__2__12), .q_2__11 (que_out_1__2__11), .q_2__10 (
            que_out_1__2__10), .q_2__9 (que_out_1__2__9), .q_2__8 (
            que_out_1__2__8), .q_2__7 (que_out_1__2__7), .q_2__6 (
            que_out_1__2__6), .q_2__5 (que_out_1__2__5), .q_2__4 (
            que_out_1__2__4), .q_2__3 (que_out_1__2__3), .q_2__2 (
            que_out_1__2__2), .q_2__1 (que_out_1__2__1), .q_2__0 (
            que_out_1__2__0), .q_3__15 (que_out_1__3__15), .q_3__14 (
            que_out_1__3__14), .q_3__13 (que_out_1__3__13), .q_3__12 (
            que_out_1__3__12), .q_3__11 (que_out_1__3__11), .q_3__10 (
            que_out_1__3__10), .q_3__9 (que_out_1__3__9), .q_3__8 (
            que_out_1__3__8), .q_3__7 (que_out_1__3__7), .q_3__6 (
            que_out_1__3__6), .q_3__5 (que_out_1__3__5), .q_3__4 (
            que_out_1__3__4), .q_3__3 (que_out_1__3__3), .q_3__2 (
            que_out_1__3__2), .q_3__1 (que_out_1__3__1), .q_3__0 (
            que_out_1__3__0), .q_4__15 (que_out_1__4__15), .q_4__14 (
            que_out_1__4__14), .q_4__13 (que_out_1__4__13), .q_4__12 (
            que_out_1__4__12), .q_4__11 (que_out_1__4__11), .q_4__10 (
            que_out_1__4__10), .q_4__9 (que_out_1__4__9), .q_4__8 (
            que_out_1__4__8), .q_4__7 (que_out_1__4__7), .q_4__6 (
            que_out_1__4__6), .q_4__5 (que_out_1__4__5), .q_4__4 (
            que_out_1__4__4), .q_4__3 (que_out_1__4__3), .q_4__2 (
            que_out_1__4__2), .q_4__1 (que_out_1__4__1), .q_4__0 (
            que_out_1__4__0), .clk (nx10714), .load (sel_que_1), .reset (nx10690
            )) ;
    Queue_5 gen_queues_2_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_2__0__15), .q_0__14 (
            que_out_2__0__14), .q_0__13 (que_out_2__0__13), .q_0__12 (
            que_out_2__0__12), .q_0__11 (que_out_2__0__11), .q_0__10 (
            que_out_2__0__10), .q_0__9 (que_out_2__0__9), .q_0__8 (
            que_out_2__0__8), .q_0__7 (que_out_2__0__7), .q_0__6 (
            que_out_2__0__6), .q_0__5 (que_out_2__0__5), .q_0__4 (
            que_out_2__0__4), .q_0__3 (que_out_2__0__3), .q_0__2 (
            que_out_2__0__2), .q_0__1 (que_out_2__0__1), .q_0__0 (
            que_out_2__0__0), .q_1__15 (que_out_2__1__15), .q_1__14 (
            que_out_2__1__14), .q_1__13 (que_out_2__1__13), .q_1__12 (
            que_out_2__1__12), .q_1__11 (que_out_2__1__11), .q_1__10 (
            que_out_2__1__10), .q_1__9 (que_out_2__1__9), .q_1__8 (
            que_out_2__1__8), .q_1__7 (que_out_2__1__7), .q_1__6 (
            que_out_2__1__6), .q_1__5 (que_out_2__1__5), .q_1__4 (
            que_out_2__1__4), .q_1__3 (que_out_2__1__3), .q_1__2 (
            que_out_2__1__2), .q_1__1 (que_out_2__1__1), .q_1__0 (
            que_out_2__1__0), .q_2__15 (que_out_2__2__15), .q_2__14 (
            que_out_2__2__14), .q_2__13 (que_out_2__2__13), .q_2__12 (
            que_out_2__2__12), .q_2__11 (que_out_2__2__11), .q_2__10 (
            que_out_2__2__10), .q_2__9 (que_out_2__2__9), .q_2__8 (
            que_out_2__2__8), .q_2__7 (que_out_2__2__7), .q_2__6 (
            que_out_2__2__6), .q_2__5 (que_out_2__2__5), .q_2__4 (
            que_out_2__2__4), .q_2__3 (que_out_2__2__3), .q_2__2 (
            que_out_2__2__2), .q_2__1 (que_out_2__2__1), .q_2__0 (
            que_out_2__2__0), .q_3__15 (que_out_2__3__15), .q_3__14 (
            que_out_2__3__14), .q_3__13 (que_out_2__3__13), .q_3__12 (
            que_out_2__3__12), .q_3__11 (que_out_2__3__11), .q_3__10 (
            que_out_2__3__10), .q_3__9 (que_out_2__3__9), .q_3__8 (
            que_out_2__3__8), .q_3__7 (que_out_2__3__7), .q_3__6 (
            que_out_2__3__6), .q_3__5 (que_out_2__3__5), .q_3__4 (
            que_out_2__3__4), .q_3__3 (que_out_2__3__3), .q_3__2 (
            que_out_2__3__2), .q_3__1 (que_out_2__3__1), .q_3__0 (
            que_out_2__3__0), .q_4__15 (que_out_2__4__15), .q_4__14 (
            que_out_2__4__14), .q_4__13 (que_out_2__4__13), .q_4__12 (
            que_out_2__4__12), .q_4__11 (que_out_2__4__11), .q_4__10 (
            que_out_2__4__10), .q_4__9 (que_out_2__4__9), .q_4__8 (
            que_out_2__4__8), .q_4__7 (que_out_2__4__7), .q_4__6 (
            que_out_2__4__6), .q_4__5 (que_out_2__4__5), .q_4__4 (
            que_out_2__4__4), .q_4__3 (que_out_2__4__3), .q_4__2 (
            que_out_2__4__2), .q_4__1 (que_out_2__4__1), .q_4__0 (
            que_out_2__4__0), .clk (nx10714), .load (sel_que_2), .reset (nx10690
            )) ;
    Queue_5 gen_queues_3_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_3__0__15), .q_0__14 (
            que_out_3__0__14), .q_0__13 (que_out_3__0__13), .q_0__12 (
            que_out_3__0__12), .q_0__11 (que_out_3__0__11), .q_0__10 (
            que_out_3__0__10), .q_0__9 (que_out_3__0__9), .q_0__8 (
            que_out_3__0__8), .q_0__7 (que_out_3__0__7), .q_0__6 (
            que_out_3__0__6), .q_0__5 (que_out_3__0__5), .q_0__4 (
            que_out_3__0__4), .q_0__3 (que_out_3__0__3), .q_0__2 (
            que_out_3__0__2), .q_0__1 (que_out_3__0__1), .q_0__0 (
            que_out_3__0__0), .q_1__15 (que_out_3__1__15), .q_1__14 (
            que_out_3__1__14), .q_1__13 (que_out_3__1__13), .q_1__12 (
            que_out_3__1__12), .q_1__11 (que_out_3__1__11), .q_1__10 (
            que_out_3__1__10), .q_1__9 (que_out_3__1__9), .q_1__8 (
            que_out_3__1__8), .q_1__7 (que_out_3__1__7), .q_1__6 (
            que_out_3__1__6), .q_1__5 (que_out_3__1__5), .q_1__4 (
            que_out_3__1__4), .q_1__3 (que_out_3__1__3), .q_1__2 (
            que_out_3__1__2), .q_1__1 (que_out_3__1__1), .q_1__0 (
            que_out_3__1__0), .q_2__15 (que_out_3__2__15), .q_2__14 (
            que_out_3__2__14), .q_2__13 (que_out_3__2__13), .q_2__12 (
            que_out_3__2__12), .q_2__11 (que_out_3__2__11), .q_2__10 (
            que_out_3__2__10), .q_2__9 (que_out_3__2__9), .q_2__8 (
            que_out_3__2__8), .q_2__7 (que_out_3__2__7), .q_2__6 (
            que_out_3__2__6), .q_2__5 (que_out_3__2__5), .q_2__4 (
            que_out_3__2__4), .q_2__3 (que_out_3__2__3), .q_2__2 (
            que_out_3__2__2), .q_2__1 (que_out_3__2__1), .q_2__0 (
            que_out_3__2__0), .q_3__15 (que_out_3__3__15), .q_3__14 (
            que_out_3__3__14), .q_3__13 (que_out_3__3__13), .q_3__12 (
            que_out_3__3__12), .q_3__11 (que_out_3__3__11), .q_3__10 (
            que_out_3__3__10), .q_3__9 (que_out_3__3__9), .q_3__8 (
            que_out_3__3__8), .q_3__7 (que_out_3__3__7), .q_3__6 (
            que_out_3__3__6), .q_3__5 (que_out_3__3__5), .q_3__4 (
            que_out_3__3__4), .q_3__3 (que_out_3__3__3), .q_3__2 (
            que_out_3__3__2), .q_3__1 (que_out_3__3__1), .q_3__0 (
            que_out_3__3__0), .q_4__15 (que_out_3__4__15), .q_4__14 (
            que_out_3__4__14), .q_4__13 (que_out_3__4__13), .q_4__12 (
            que_out_3__4__12), .q_4__11 (que_out_3__4__11), .q_4__10 (
            que_out_3__4__10), .q_4__9 (que_out_3__4__9), .q_4__8 (
            que_out_3__4__8), .q_4__7 (que_out_3__4__7), .q_4__6 (
            que_out_3__4__6), .q_4__5 (que_out_3__4__5), .q_4__4 (
            que_out_3__4__4), .q_4__3 (que_out_3__4__3), .q_4__2 (
            que_out_3__4__2), .q_4__1 (que_out_3__4__1), .q_4__0 (
            que_out_3__4__0), .clk (nx10716), .load (sel_que_3), .reset (nx10692
            )) ;
    Queue_5 gen_queues_4_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_4__0__15), .q_0__14 (
            que_out_4__0__14), .q_0__13 (que_out_4__0__13), .q_0__12 (
            que_out_4__0__12), .q_0__11 (que_out_4__0__11), .q_0__10 (
            que_out_4__0__10), .q_0__9 (que_out_4__0__9), .q_0__8 (
            que_out_4__0__8), .q_0__7 (que_out_4__0__7), .q_0__6 (
            que_out_4__0__6), .q_0__5 (que_out_4__0__5), .q_0__4 (
            que_out_4__0__4), .q_0__3 (que_out_4__0__3), .q_0__2 (
            que_out_4__0__2), .q_0__1 (que_out_4__0__1), .q_0__0 (
            que_out_4__0__0), .q_1__15 (que_out_4__1__15), .q_1__14 (
            que_out_4__1__14), .q_1__13 (que_out_4__1__13), .q_1__12 (
            que_out_4__1__12), .q_1__11 (que_out_4__1__11), .q_1__10 (
            que_out_4__1__10), .q_1__9 (que_out_4__1__9), .q_1__8 (
            que_out_4__1__8), .q_1__7 (que_out_4__1__7), .q_1__6 (
            que_out_4__1__6), .q_1__5 (que_out_4__1__5), .q_1__4 (
            que_out_4__1__4), .q_1__3 (que_out_4__1__3), .q_1__2 (
            que_out_4__1__2), .q_1__1 (que_out_4__1__1), .q_1__0 (
            que_out_4__1__0), .q_2__15 (que_out_4__2__15), .q_2__14 (
            que_out_4__2__14), .q_2__13 (que_out_4__2__13), .q_2__12 (
            que_out_4__2__12), .q_2__11 (que_out_4__2__11), .q_2__10 (
            que_out_4__2__10), .q_2__9 (que_out_4__2__9), .q_2__8 (
            que_out_4__2__8), .q_2__7 (que_out_4__2__7), .q_2__6 (
            que_out_4__2__6), .q_2__5 (que_out_4__2__5), .q_2__4 (
            que_out_4__2__4), .q_2__3 (que_out_4__2__3), .q_2__2 (
            que_out_4__2__2), .q_2__1 (que_out_4__2__1), .q_2__0 (
            que_out_4__2__0), .q_3__15 (que_out_4__3__15), .q_3__14 (
            que_out_4__3__14), .q_3__13 (que_out_4__3__13), .q_3__12 (
            que_out_4__3__12), .q_3__11 (que_out_4__3__11), .q_3__10 (
            que_out_4__3__10), .q_3__9 (que_out_4__3__9), .q_3__8 (
            que_out_4__3__8), .q_3__7 (que_out_4__3__7), .q_3__6 (
            que_out_4__3__6), .q_3__5 (que_out_4__3__5), .q_3__4 (
            que_out_4__3__4), .q_3__3 (que_out_4__3__3), .q_3__2 (
            que_out_4__3__2), .q_3__1 (que_out_4__3__1), .q_3__0 (
            que_out_4__3__0), .q_4__15 (que_out_4__4__15), .q_4__14 (
            que_out_4__4__14), .q_4__13 (que_out_4__4__13), .q_4__12 (
            que_out_4__4__12), .q_4__11 (que_out_4__4__11), .q_4__10 (
            que_out_4__4__10), .q_4__9 (que_out_4__4__9), .q_4__8 (
            que_out_4__4__8), .q_4__7 (que_out_4__4__7), .q_4__6 (
            que_out_4__4__6), .q_4__5 (que_out_4__4__5), .q_4__4 (
            que_out_4__4__4), .q_4__3 (que_out_4__4__3), .q_4__2 (
            que_out_4__4__2), .q_4__1 (que_out_4__4__1), .q_4__0 (
            que_out_4__4__0), .clk (nx10716), .load (sel_que_4), .reset (nx10692
            )) ;
    Queue_5 gen_queues_5_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_5__0__15), .q_0__14 (
            que_out_5__0__14), .q_0__13 (que_out_5__0__13), .q_0__12 (
            que_out_5__0__12), .q_0__11 (que_out_5__0__11), .q_0__10 (
            que_out_5__0__10), .q_0__9 (que_out_5__0__9), .q_0__8 (
            que_out_5__0__8), .q_0__7 (que_out_5__0__7), .q_0__6 (
            que_out_5__0__6), .q_0__5 (que_out_5__0__5), .q_0__4 (
            que_out_5__0__4), .q_0__3 (que_out_5__0__3), .q_0__2 (
            que_out_5__0__2), .q_0__1 (que_out_5__0__1), .q_0__0 (
            que_out_5__0__0), .q_1__15 (que_out_5__1__15), .q_1__14 (
            que_out_5__1__14), .q_1__13 (que_out_5__1__13), .q_1__12 (
            que_out_5__1__12), .q_1__11 (que_out_5__1__11), .q_1__10 (
            que_out_5__1__10), .q_1__9 (que_out_5__1__9), .q_1__8 (
            que_out_5__1__8), .q_1__7 (que_out_5__1__7), .q_1__6 (
            que_out_5__1__6), .q_1__5 (que_out_5__1__5), .q_1__4 (
            que_out_5__1__4), .q_1__3 (que_out_5__1__3), .q_1__2 (
            que_out_5__1__2), .q_1__1 (que_out_5__1__1), .q_1__0 (
            que_out_5__1__0), .q_2__15 (que_out_5__2__15), .q_2__14 (
            que_out_5__2__14), .q_2__13 (que_out_5__2__13), .q_2__12 (
            que_out_5__2__12), .q_2__11 (que_out_5__2__11), .q_2__10 (
            que_out_5__2__10), .q_2__9 (que_out_5__2__9), .q_2__8 (
            que_out_5__2__8), .q_2__7 (que_out_5__2__7), .q_2__6 (
            que_out_5__2__6), .q_2__5 (que_out_5__2__5), .q_2__4 (
            que_out_5__2__4), .q_2__3 (que_out_5__2__3), .q_2__2 (
            que_out_5__2__2), .q_2__1 (que_out_5__2__1), .q_2__0 (
            que_out_5__2__0), .q_3__15 (que_out_5__3__15), .q_3__14 (
            que_out_5__3__14), .q_3__13 (que_out_5__3__13), .q_3__12 (
            que_out_5__3__12), .q_3__11 (que_out_5__3__11), .q_3__10 (
            que_out_5__3__10), .q_3__9 (que_out_5__3__9), .q_3__8 (
            que_out_5__3__8), .q_3__7 (que_out_5__3__7), .q_3__6 (
            que_out_5__3__6), .q_3__5 (que_out_5__3__5), .q_3__4 (
            que_out_5__3__4), .q_3__3 (que_out_5__3__3), .q_3__2 (
            que_out_5__3__2), .q_3__1 (que_out_5__3__1), .q_3__0 (
            que_out_5__3__0), .q_4__15 (que_out_5__4__15), .q_4__14 (
            que_out_5__4__14), .q_4__13 (que_out_5__4__13), .q_4__12 (
            que_out_5__4__12), .q_4__11 (que_out_5__4__11), .q_4__10 (
            que_out_5__4__10), .q_4__9 (que_out_5__4__9), .q_4__8 (
            que_out_5__4__8), .q_4__7 (que_out_5__4__7), .q_4__6 (
            que_out_5__4__6), .q_4__5 (que_out_5__4__5), .q_4__4 (
            que_out_5__4__4), .q_4__3 (que_out_5__4__3), .q_4__2 (
            que_out_5__4__2), .q_4__1 (que_out_5__4__1), .q_4__0 (
            que_out_5__4__0), .clk (nx10716), .load (sel_que_5), .reset (nx10692
            )) ;
    Queue_5 gen_queues_6_que (.d ({nx10512,nx10522,nx10532,nx10542,nx10552,
            nx10562,nx10572,nx10582,nx10592,nx10602,nx10612,nx10622,nx10632,
            nx10642,nx10652,nx10662}), .q_0__15 (que_out_6__0__15), .q_0__14 (
            que_out_6__0__14), .q_0__13 (que_out_6__0__13), .q_0__12 (
            que_out_6__0__12), .q_0__11 (que_out_6__0__11), .q_0__10 (
            que_out_6__0__10), .q_0__9 (que_out_6__0__9), .q_0__8 (
            que_out_6__0__8), .q_0__7 (que_out_6__0__7), .q_0__6 (
            que_out_6__0__6), .q_0__5 (que_out_6__0__5), .q_0__4 (
            que_out_6__0__4), .q_0__3 (que_out_6__0__3), .q_0__2 (
            que_out_6__0__2), .q_0__1 (que_out_6__0__1), .q_0__0 (
            que_out_6__0__0), .q_1__15 (que_out_6__1__15), .q_1__14 (
            que_out_6__1__14), .q_1__13 (que_out_6__1__13), .q_1__12 (
            que_out_6__1__12), .q_1__11 (que_out_6__1__11), .q_1__10 (
            que_out_6__1__10), .q_1__9 (que_out_6__1__9), .q_1__8 (
            que_out_6__1__8), .q_1__7 (que_out_6__1__7), .q_1__6 (
            que_out_6__1__6), .q_1__5 (que_out_6__1__5), .q_1__4 (
            que_out_6__1__4), .q_1__3 (que_out_6__1__3), .q_1__2 (
            que_out_6__1__2), .q_1__1 (que_out_6__1__1), .q_1__0 (
            que_out_6__1__0), .q_2__15 (que_out_6__2__15), .q_2__14 (
            que_out_6__2__14), .q_2__13 (que_out_6__2__13), .q_2__12 (
            que_out_6__2__12), .q_2__11 (que_out_6__2__11), .q_2__10 (
            que_out_6__2__10), .q_2__9 (que_out_6__2__9), .q_2__8 (
            que_out_6__2__8), .q_2__7 (que_out_6__2__7), .q_2__6 (
            que_out_6__2__6), .q_2__5 (que_out_6__2__5), .q_2__4 (
            que_out_6__2__4), .q_2__3 (que_out_6__2__3), .q_2__2 (
            que_out_6__2__2), .q_2__1 (que_out_6__2__1), .q_2__0 (
            que_out_6__2__0), .q_3__15 (que_out_6__3__15), .q_3__14 (
            que_out_6__3__14), .q_3__13 (que_out_6__3__13), .q_3__12 (
            que_out_6__3__12), .q_3__11 (que_out_6__3__11), .q_3__10 (
            que_out_6__3__10), .q_3__9 (que_out_6__3__9), .q_3__8 (
            que_out_6__3__8), .q_3__7 (que_out_6__3__7), .q_3__6 (
            que_out_6__3__6), .q_3__5 (que_out_6__3__5), .q_3__4 (
            que_out_6__3__4), .q_3__3 (que_out_6__3__3), .q_3__2 (
            que_out_6__3__2), .q_3__1 (que_out_6__3__1), .q_3__0 (
            que_out_6__3__0), .q_4__15 (que_out_6__4__15), .q_4__14 (
            que_out_6__4__14), .q_4__13 (que_out_6__4__13), .q_4__12 (
            que_out_6__4__12), .q_4__11 (que_out_6__4__11), .q_4__10 (
            que_out_6__4__10), .q_4__9 (que_out_6__4__9), .q_4__8 (
            que_out_6__4__8), .q_4__7 (que_out_6__4__7), .q_4__6 (
            que_out_6__4__6), .q_4__5 (que_out_6__4__5), .q_4__4 (
            que_out_6__4__4), .q_4__3 (que_out_6__4__3), .q_4__2 (
            que_out_6__4__2), .q_4__1 (que_out_6__4__1), .q_4__0 (
            que_out_6__4__0), .clk (nx10718), .load (sel_que_6), .reset (nx10694
            )) ;
    Queue_5 gen_queues_7_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_7__0__15), .q_0__14 (
            que_out_7__0__14), .q_0__13 (que_out_7__0__13), .q_0__12 (
            que_out_7__0__12), .q_0__11 (que_out_7__0__11), .q_0__10 (
            que_out_7__0__10), .q_0__9 (que_out_7__0__9), .q_0__8 (
            que_out_7__0__8), .q_0__7 (que_out_7__0__7), .q_0__6 (
            que_out_7__0__6), .q_0__5 (que_out_7__0__5), .q_0__4 (
            que_out_7__0__4), .q_0__3 (que_out_7__0__3), .q_0__2 (
            que_out_7__0__2), .q_0__1 (que_out_7__0__1), .q_0__0 (
            que_out_7__0__0), .q_1__15 (que_out_7__1__15), .q_1__14 (
            que_out_7__1__14), .q_1__13 (que_out_7__1__13), .q_1__12 (
            que_out_7__1__12), .q_1__11 (que_out_7__1__11), .q_1__10 (
            que_out_7__1__10), .q_1__9 (que_out_7__1__9), .q_1__8 (
            que_out_7__1__8), .q_1__7 (que_out_7__1__7), .q_1__6 (
            que_out_7__1__6), .q_1__5 (que_out_7__1__5), .q_1__4 (
            que_out_7__1__4), .q_1__3 (que_out_7__1__3), .q_1__2 (
            que_out_7__1__2), .q_1__1 (que_out_7__1__1), .q_1__0 (
            que_out_7__1__0), .q_2__15 (que_out_7__2__15), .q_2__14 (
            que_out_7__2__14), .q_2__13 (que_out_7__2__13), .q_2__12 (
            que_out_7__2__12), .q_2__11 (que_out_7__2__11), .q_2__10 (
            que_out_7__2__10), .q_2__9 (que_out_7__2__9), .q_2__8 (
            que_out_7__2__8), .q_2__7 (que_out_7__2__7), .q_2__6 (
            que_out_7__2__6), .q_2__5 (que_out_7__2__5), .q_2__4 (
            que_out_7__2__4), .q_2__3 (que_out_7__2__3), .q_2__2 (
            que_out_7__2__2), .q_2__1 (que_out_7__2__1), .q_2__0 (
            que_out_7__2__0), .q_3__15 (que_out_7__3__15), .q_3__14 (
            que_out_7__3__14), .q_3__13 (que_out_7__3__13), .q_3__12 (
            que_out_7__3__12), .q_3__11 (que_out_7__3__11), .q_3__10 (
            que_out_7__3__10), .q_3__9 (que_out_7__3__9), .q_3__8 (
            que_out_7__3__8), .q_3__7 (que_out_7__3__7), .q_3__6 (
            que_out_7__3__6), .q_3__5 (que_out_7__3__5), .q_3__4 (
            que_out_7__3__4), .q_3__3 (que_out_7__3__3), .q_3__2 (
            que_out_7__3__2), .q_3__1 (que_out_7__3__1), .q_3__0 (
            que_out_7__3__0), .q_4__15 (que_out_7__4__15), .q_4__14 (
            que_out_7__4__14), .q_4__13 (que_out_7__4__13), .q_4__12 (
            que_out_7__4__12), .q_4__11 (que_out_7__4__11), .q_4__10 (
            que_out_7__4__10), .q_4__9 (que_out_7__4__9), .q_4__8 (
            que_out_7__4__8), .q_4__7 (que_out_7__4__7), .q_4__6 (
            que_out_7__4__6), .q_4__5 (que_out_7__4__5), .q_4__4 (
            que_out_7__4__4), .q_4__3 (que_out_7__4__3), .q_4__2 (
            que_out_7__4__2), .q_4__1 (que_out_7__4__1), .q_4__0 (
            que_out_7__4__0), .clk (nx10720), .load (sel_que_7), .reset (nx10696
            )) ;
    Queue_5 gen_queues_8_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_8__0__15), .q_0__14 (
            que_out_8__0__14), .q_0__13 (que_out_8__0__13), .q_0__12 (
            que_out_8__0__12), .q_0__11 (que_out_8__0__11), .q_0__10 (
            que_out_8__0__10), .q_0__9 (que_out_8__0__9), .q_0__8 (
            que_out_8__0__8), .q_0__7 (que_out_8__0__7), .q_0__6 (
            que_out_8__0__6), .q_0__5 (que_out_8__0__5), .q_0__4 (
            que_out_8__0__4), .q_0__3 (que_out_8__0__3), .q_0__2 (
            que_out_8__0__2), .q_0__1 (que_out_8__0__1), .q_0__0 (
            que_out_8__0__0), .q_1__15 (que_out_8__1__15), .q_1__14 (
            que_out_8__1__14), .q_1__13 (que_out_8__1__13), .q_1__12 (
            que_out_8__1__12), .q_1__11 (que_out_8__1__11), .q_1__10 (
            que_out_8__1__10), .q_1__9 (que_out_8__1__9), .q_1__8 (
            que_out_8__1__8), .q_1__7 (que_out_8__1__7), .q_1__6 (
            que_out_8__1__6), .q_1__5 (que_out_8__1__5), .q_1__4 (
            que_out_8__1__4), .q_1__3 (que_out_8__1__3), .q_1__2 (
            que_out_8__1__2), .q_1__1 (que_out_8__1__1), .q_1__0 (
            que_out_8__1__0), .q_2__15 (que_out_8__2__15), .q_2__14 (
            que_out_8__2__14), .q_2__13 (que_out_8__2__13), .q_2__12 (
            que_out_8__2__12), .q_2__11 (que_out_8__2__11), .q_2__10 (
            que_out_8__2__10), .q_2__9 (que_out_8__2__9), .q_2__8 (
            que_out_8__2__8), .q_2__7 (que_out_8__2__7), .q_2__6 (
            que_out_8__2__6), .q_2__5 (que_out_8__2__5), .q_2__4 (
            que_out_8__2__4), .q_2__3 (que_out_8__2__3), .q_2__2 (
            que_out_8__2__2), .q_2__1 (que_out_8__2__1), .q_2__0 (
            que_out_8__2__0), .q_3__15 (que_out_8__3__15), .q_3__14 (
            que_out_8__3__14), .q_3__13 (que_out_8__3__13), .q_3__12 (
            que_out_8__3__12), .q_3__11 (que_out_8__3__11), .q_3__10 (
            que_out_8__3__10), .q_3__9 (que_out_8__3__9), .q_3__8 (
            que_out_8__3__8), .q_3__7 (que_out_8__3__7), .q_3__6 (
            que_out_8__3__6), .q_3__5 (que_out_8__3__5), .q_3__4 (
            que_out_8__3__4), .q_3__3 (que_out_8__3__3), .q_3__2 (
            que_out_8__3__2), .q_3__1 (que_out_8__3__1), .q_3__0 (
            que_out_8__3__0), .q_4__15 (que_out_8__4__15), .q_4__14 (
            que_out_8__4__14), .q_4__13 (que_out_8__4__13), .q_4__12 (
            que_out_8__4__12), .q_4__11 (que_out_8__4__11), .q_4__10 (
            que_out_8__4__10), .q_4__9 (que_out_8__4__9), .q_4__8 (
            que_out_8__4__8), .q_4__7 (que_out_8__4__7), .q_4__6 (
            que_out_8__4__6), .q_4__5 (que_out_8__4__5), .q_4__4 (
            que_out_8__4__4), .q_4__3 (que_out_8__4__3), .q_4__2 (
            que_out_8__4__2), .q_4__1 (que_out_8__4__1), .q_4__0 (
            que_out_8__4__0), .clk (nx10720), .load (sel_que_8), .reset (nx10696
            )) ;
    Queue_5 gen_queues_9_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_9__0__15), .q_0__14 (
            que_out_9__0__14), .q_0__13 (que_out_9__0__13), .q_0__12 (
            que_out_9__0__12), .q_0__11 (que_out_9__0__11), .q_0__10 (
            que_out_9__0__10), .q_0__9 (que_out_9__0__9), .q_0__8 (
            que_out_9__0__8), .q_0__7 (que_out_9__0__7), .q_0__6 (
            que_out_9__0__6), .q_0__5 (que_out_9__0__5), .q_0__4 (
            que_out_9__0__4), .q_0__3 (que_out_9__0__3), .q_0__2 (
            que_out_9__0__2), .q_0__1 (que_out_9__0__1), .q_0__0 (
            que_out_9__0__0), .q_1__15 (que_out_9__1__15), .q_1__14 (
            que_out_9__1__14), .q_1__13 (que_out_9__1__13), .q_1__12 (
            que_out_9__1__12), .q_1__11 (que_out_9__1__11), .q_1__10 (
            que_out_9__1__10), .q_1__9 (que_out_9__1__9), .q_1__8 (
            que_out_9__1__8), .q_1__7 (que_out_9__1__7), .q_1__6 (
            que_out_9__1__6), .q_1__5 (que_out_9__1__5), .q_1__4 (
            que_out_9__1__4), .q_1__3 (que_out_9__1__3), .q_1__2 (
            que_out_9__1__2), .q_1__1 (que_out_9__1__1), .q_1__0 (
            que_out_9__1__0), .q_2__15 (que_out_9__2__15), .q_2__14 (
            que_out_9__2__14), .q_2__13 (que_out_9__2__13), .q_2__12 (
            que_out_9__2__12), .q_2__11 (que_out_9__2__11), .q_2__10 (
            que_out_9__2__10), .q_2__9 (que_out_9__2__9), .q_2__8 (
            que_out_9__2__8), .q_2__7 (que_out_9__2__7), .q_2__6 (
            que_out_9__2__6), .q_2__5 (que_out_9__2__5), .q_2__4 (
            que_out_9__2__4), .q_2__3 (que_out_9__2__3), .q_2__2 (
            que_out_9__2__2), .q_2__1 (que_out_9__2__1), .q_2__0 (
            que_out_9__2__0), .q_3__15 (que_out_9__3__15), .q_3__14 (
            que_out_9__3__14), .q_3__13 (que_out_9__3__13), .q_3__12 (
            que_out_9__3__12), .q_3__11 (que_out_9__3__11), .q_3__10 (
            que_out_9__3__10), .q_3__9 (que_out_9__3__9), .q_3__8 (
            que_out_9__3__8), .q_3__7 (que_out_9__3__7), .q_3__6 (
            que_out_9__3__6), .q_3__5 (que_out_9__3__5), .q_3__4 (
            que_out_9__3__4), .q_3__3 (que_out_9__3__3), .q_3__2 (
            que_out_9__3__2), .q_3__1 (que_out_9__3__1), .q_3__0 (
            que_out_9__3__0), .q_4__15 (que_out_9__4__15), .q_4__14 (
            que_out_9__4__14), .q_4__13 (que_out_9__4__13), .q_4__12 (
            que_out_9__4__12), .q_4__11 (que_out_9__4__11), .q_4__10 (
            que_out_9__4__10), .q_4__9 (que_out_9__4__9), .q_4__8 (
            que_out_9__4__8), .q_4__7 (que_out_9__4__7), .q_4__6 (
            que_out_9__4__6), .q_4__5 (que_out_9__4__5), .q_4__4 (
            que_out_9__4__4), .q_4__3 (que_out_9__4__3), .q_4__2 (
            que_out_9__4__2), .q_4__1 (que_out_9__4__1), .q_4__0 (
            que_out_9__4__0), .clk (nx10720), .load (sel_que_9), .reset (nx10696
            )) ;
    Queue_5 gen_queues_10_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_10__0__15), .q_0__14 (
            que_out_10__0__14), .q_0__13 (que_out_10__0__13), .q_0__12 (
            que_out_10__0__12), .q_0__11 (que_out_10__0__11), .q_0__10 (
            que_out_10__0__10), .q_0__9 (que_out_10__0__9), .q_0__8 (
            que_out_10__0__8), .q_0__7 (que_out_10__0__7), .q_0__6 (
            que_out_10__0__6), .q_0__5 (que_out_10__0__5), .q_0__4 (
            que_out_10__0__4), .q_0__3 (que_out_10__0__3), .q_0__2 (
            que_out_10__0__2), .q_0__1 (que_out_10__0__1), .q_0__0 (
            que_out_10__0__0), .q_1__15 (que_out_10__1__15), .q_1__14 (
            que_out_10__1__14), .q_1__13 (que_out_10__1__13), .q_1__12 (
            que_out_10__1__12), .q_1__11 (que_out_10__1__11), .q_1__10 (
            que_out_10__1__10), .q_1__9 (que_out_10__1__9), .q_1__8 (
            que_out_10__1__8), .q_1__7 (que_out_10__1__7), .q_1__6 (
            que_out_10__1__6), .q_1__5 (que_out_10__1__5), .q_1__4 (
            que_out_10__1__4), .q_1__3 (que_out_10__1__3), .q_1__2 (
            que_out_10__1__2), .q_1__1 (que_out_10__1__1), .q_1__0 (
            que_out_10__1__0), .q_2__15 (que_out_10__2__15), .q_2__14 (
            que_out_10__2__14), .q_2__13 (que_out_10__2__13), .q_2__12 (
            que_out_10__2__12), .q_2__11 (que_out_10__2__11), .q_2__10 (
            que_out_10__2__10), .q_2__9 (que_out_10__2__9), .q_2__8 (
            que_out_10__2__8), .q_2__7 (que_out_10__2__7), .q_2__6 (
            que_out_10__2__6), .q_2__5 (que_out_10__2__5), .q_2__4 (
            que_out_10__2__4), .q_2__3 (que_out_10__2__3), .q_2__2 (
            que_out_10__2__2), .q_2__1 (que_out_10__2__1), .q_2__0 (
            que_out_10__2__0), .q_3__15 (que_out_10__3__15), .q_3__14 (
            que_out_10__3__14), .q_3__13 (que_out_10__3__13), .q_3__12 (
            que_out_10__3__12), .q_3__11 (que_out_10__3__11), .q_3__10 (
            que_out_10__3__10), .q_3__9 (que_out_10__3__9), .q_3__8 (
            que_out_10__3__8), .q_3__7 (que_out_10__3__7), .q_3__6 (
            que_out_10__3__6), .q_3__5 (que_out_10__3__5), .q_3__4 (
            que_out_10__3__4), .q_3__3 (que_out_10__3__3), .q_3__2 (
            que_out_10__3__2), .q_3__1 (que_out_10__3__1), .q_3__0 (
            que_out_10__3__0), .q_4__15 (que_out_10__4__15), .q_4__14 (
            que_out_10__4__14), .q_4__13 (que_out_10__4__13), .q_4__12 (
            que_out_10__4__12), .q_4__11 (que_out_10__4__11), .q_4__10 (
            que_out_10__4__10), .q_4__9 (que_out_10__4__9), .q_4__8 (
            que_out_10__4__8), .q_4__7 (que_out_10__4__7), .q_4__6 (
            que_out_10__4__6), .q_4__5 (que_out_10__4__5), .q_4__4 (
            que_out_10__4__4), .q_4__3 (que_out_10__4__3), .q_4__2 (
            que_out_10__4__2), .q_4__1 (que_out_10__4__1), .q_4__0 (
            que_out_10__4__0), .clk (nx10722), .load (sel_que_10), .reset (
            nx10698)) ;
    Queue_5 gen_queues_11_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_11__0__15), .q_0__14 (
            que_out_11__0__14), .q_0__13 (que_out_11__0__13), .q_0__12 (
            que_out_11__0__12), .q_0__11 (que_out_11__0__11), .q_0__10 (
            que_out_11__0__10), .q_0__9 (que_out_11__0__9), .q_0__8 (
            que_out_11__0__8), .q_0__7 (que_out_11__0__7), .q_0__6 (
            que_out_11__0__6), .q_0__5 (que_out_11__0__5), .q_0__4 (
            que_out_11__0__4), .q_0__3 (que_out_11__0__3), .q_0__2 (
            que_out_11__0__2), .q_0__1 (que_out_11__0__1), .q_0__0 (
            que_out_11__0__0), .q_1__15 (que_out_11__1__15), .q_1__14 (
            que_out_11__1__14), .q_1__13 (que_out_11__1__13), .q_1__12 (
            que_out_11__1__12), .q_1__11 (que_out_11__1__11), .q_1__10 (
            que_out_11__1__10), .q_1__9 (que_out_11__1__9), .q_1__8 (
            que_out_11__1__8), .q_1__7 (que_out_11__1__7), .q_1__6 (
            que_out_11__1__6), .q_1__5 (que_out_11__1__5), .q_1__4 (
            que_out_11__1__4), .q_1__3 (que_out_11__1__3), .q_1__2 (
            que_out_11__1__2), .q_1__1 (que_out_11__1__1), .q_1__0 (
            que_out_11__1__0), .q_2__15 (que_out_11__2__15), .q_2__14 (
            que_out_11__2__14), .q_2__13 (que_out_11__2__13), .q_2__12 (
            que_out_11__2__12), .q_2__11 (que_out_11__2__11), .q_2__10 (
            que_out_11__2__10), .q_2__9 (que_out_11__2__9), .q_2__8 (
            que_out_11__2__8), .q_2__7 (que_out_11__2__7), .q_2__6 (
            que_out_11__2__6), .q_2__5 (que_out_11__2__5), .q_2__4 (
            que_out_11__2__4), .q_2__3 (que_out_11__2__3), .q_2__2 (
            que_out_11__2__2), .q_2__1 (que_out_11__2__1), .q_2__0 (
            que_out_11__2__0), .q_3__15 (que_out_11__3__15), .q_3__14 (
            que_out_11__3__14), .q_3__13 (que_out_11__3__13), .q_3__12 (
            que_out_11__3__12), .q_3__11 (que_out_11__3__11), .q_3__10 (
            que_out_11__3__10), .q_3__9 (que_out_11__3__9), .q_3__8 (
            que_out_11__3__8), .q_3__7 (que_out_11__3__7), .q_3__6 (
            que_out_11__3__6), .q_3__5 (que_out_11__3__5), .q_3__4 (
            que_out_11__3__4), .q_3__3 (que_out_11__3__3), .q_3__2 (
            que_out_11__3__2), .q_3__1 (que_out_11__3__1), .q_3__0 (
            que_out_11__3__0), .q_4__15 (que_out_11__4__15), .q_4__14 (
            que_out_11__4__14), .q_4__13 (que_out_11__4__13), .q_4__12 (
            que_out_11__4__12), .q_4__11 (que_out_11__4__11), .q_4__10 (
            que_out_11__4__10), .q_4__9 (que_out_11__4__9), .q_4__8 (
            que_out_11__4__8), .q_4__7 (que_out_11__4__7), .q_4__6 (
            que_out_11__4__6), .q_4__5 (que_out_11__4__5), .q_4__4 (
            que_out_11__4__4), .q_4__3 (que_out_11__4__3), .q_4__2 (
            que_out_11__4__2), .q_4__1 (que_out_11__4__1), .q_4__0 (
            que_out_11__4__0), .clk (nx10722), .load (sel_que_11), .reset (
            nx10698)) ;
    Queue_5 gen_queues_12_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_12__0__15), .q_0__14 (
            que_out_12__0__14), .q_0__13 (que_out_12__0__13), .q_0__12 (
            que_out_12__0__12), .q_0__11 (que_out_12__0__11), .q_0__10 (
            que_out_12__0__10), .q_0__9 (que_out_12__0__9), .q_0__8 (
            que_out_12__0__8), .q_0__7 (que_out_12__0__7), .q_0__6 (
            que_out_12__0__6), .q_0__5 (que_out_12__0__5), .q_0__4 (
            que_out_12__0__4), .q_0__3 (que_out_12__0__3), .q_0__2 (
            que_out_12__0__2), .q_0__1 (que_out_12__0__1), .q_0__0 (
            que_out_12__0__0), .q_1__15 (que_out_12__1__15), .q_1__14 (
            que_out_12__1__14), .q_1__13 (que_out_12__1__13), .q_1__12 (
            que_out_12__1__12), .q_1__11 (que_out_12__1__11), .q_1__10 (
            que_out_12__1__10), .q_1__9 (que_out_12__1__9), .q_1__8 (
            que_out_12__1__8), .q_1__7 (que_out_12__1__7), .q_1__6 (
            que_out_12__1__6), .q_1__5 (que_out_12__1__5), .q_1__4 (
            que_out_12__1__4), .q_1__3 (que_out_12__1__3), .q_1__2 (
            que_out_12__1__2), .q_1__1 (que_out_12__1__1), .q_1__0 (
            que_out_12__1__0), .q_2__15 (que_out_12__2__15), .q_2__14 (
            que_out_12__2__14), .q_2__13 (que_out_12__2__13), .q_2__12 (
            que_out_12__2__12), .q_2__11 (que_out_12__2__11), .q_2__10 (
            que_out_12__2__10), .q_2__9 (que_out_12__2__9), .q_2__8 (
            que_out_12__2__8), .q_2__7 (que_out_12__2__7), .q_2__6 (
            que_out_12__2__6), .q_2__5 (que_out_12__2__5), .q_2__4 (
            que_out_12__2__4), .q_2__3 (que_out_12__2__3), .q_2__2 (
            que_out_12__2__2), .q_2__1 (que_out_12__2__1), .q_2__0 (
            que_out_12__2__0), .q_3__15 (que_out_12__3__15), .q_3__14 (
            que_out_12__3__14), .q_3__13 (que_out_12__3__13), .q_3__12 (
            que_out_12__3__12), .q_3__11 (que_out_12__3__11), .q_3__10 (
            que_out_12__3__10), .q_3__9 (que_out_12__3__9), .q_3__8 (
            que_out_12__3__8), .q_3__7 (que_out_12__3__7), .q_3__6 (
            que_out_12__3__6), .q_3__5 (que_out_12__3__5), .q_3__4 (
            que_out_12__3__4), .q_3__3 (que_out_12__3__3), .q_3__2 (
            que_out_12__3__2), .q_3__1 (que_out_12__3__1), .q_3__0 (
            que_out_12__3__0), .q_4__15 (que_out_12__4__15), .q_4__14 (
            que_out_12__4__14), .q_4__13 (que_out_12__4__13), .q_4__12 (
            que_out_12__4__12), .q_4__11 (que_out_12__4__11), .q_4__10 (
            que_out_12__4__10), .q_4__9 (que_out_12__4__9), .q_4__8 (
            que_out_12__4__8), .q_4__7 (que_out_12__4__7), .q_4__6 (
            que_out_12__4__6), .q_4__5 (que_out_12__4__5), .q_4__4 (
            que_out_12__4__4), .q_4__3 (que_out_12__4__3), .q_4__2 (
            que_out_12__4__2), .q_4__1 (que_out_12__4__1), .q_4__0 (
            que_out_12__4__0), .clk (nx10722), .load (sel_que_12), .reset (
            nx10698)) ;
    Queue_5 gen_queues_13_que (.d ({nx10514,nx10524,nx10534,nx10544,nx10554,
            nx10564,nx10574,nx10584,nx10594,nx10604,nx10614,nx10624,nx10634,
            nx10644,nx10654,nx10664}), .q_0__15 (que_out_13__0__15), .q_0__14 (
            que_out_13__0__14), .q_0__13 (que_out_13__0__13), .q_0__12 (
            que_out_13__0__12), .q_0__11 (que_out_13__0__11), .q_0__10 (
            que_out_13__0__10), .q_0__9 (que_out_13__0__9), .q_0__8 (
            que_out_13__0__8), .q_0__7 (que_out_13__0__7), .q_0__6 (
            que_out_13__0__6), .q_0__5 (que_out_13__0__5), .q_0__4 (
            que_out_13__0__4), .q_0__3 (que_out_13__0__3), .q_0__2 (
            que_out_13__0__2), .q_0__1 (que_out_13__0__1), .q_0__0 (
            que_out_13__0__0), .q_1__15 (que_out_13__1__15), .q_1__14 (
            que_out_13__1__14), .q_1__13 (que_out_13__1__13), .q_1__12 (
            que_out_13__1__12), .q_1__11 (que_out_13__1__11), .q_1__10 (
            que_out_13__1__10), .q_1__9 (que_out_13__1__9), .q_1__8 (
            que_out_13__1__8), .q_1__7 (que_out_13__1__7), .q_1__6 (
            que_out_13__1__6), .q_1__5 (que_out_13__1__5), .q_1__4 (
            que_out_13__1__4), .q_1__3 (que_out_13__1__3), .q_1__2 (
            que_out_13__1__2), .q_1__1 (que_out_13__1__1), .q_1__0 (
            que_out_13__1__0), .q_2__15 (que_out_13__2__15), .q_2__14 (
            que_out_13__2__14), .q_2__13 (que_out_13__2__13), .q_2__12 (
            que_out_13__2__12), .q_2__11 (que_out_13__2__11), .q_2__10 (
            que_out_13__2__10), .q_2__9 (que_out_13__2__9), .q_2__8 (
            que_out_13__2__8), .q_2__7 (que_out_13__2__7), .q_2__6 (
            que_out_13__2__6), .q_2__5 (que_out_13__2__5), .q_2__4 (
            que_out_13__2__4), .q_2__3 (que_out_13__2__3), .q_2__2 (
            que_out_13__2__2), .q_2__1 (que_out_13__2__1), .q_2__0 (
            que_out_13__2__0), .q_3__15 (que_out_13__3__15), .q_3__14 (
            que_out_13__3__14), .q_3__13 (que_out_13__3__13), .q_3__12 (
            que_out_13__3__12), .q_3__11 (que_out_13__3__11), .q_3__10 (
            que_out_13__3__10), .q_3__9 (que_out_13__3__9), .q_3__8 (
            que_out_13__3__8), .q_3__7 (que_out_13__3__7), .q_3__6 (
            que_out_13__3__6), .q_3__5 (que_out_13__3__5), .q_3__4 (
            que_out_13__3__4), .q_3__3 (que_out_13__3__3), .q_3__2 (
            que_out_13__3__2), .q_3__1 (que_out_13__3__1), .q_3__0 (
            que_out_13__3__0), .q_4__15 (que_out_13__4__15), .q_4__14 (
            que_out_13__4__14), .q_4__13 (que_out_13__4__13), .q_4__12 (
            que_out_13__4__12), .q_4__11 (que_out_13__4__11), .q_4__10 (
            que_out_13__4__10), .q_4__9 (que_out_13__4__9), .q_4__8 (
            que_out_13__4__8), .q_4__7 (que_out_13__4__7), .q_4__6 (
            que_out_13__4__6), .q_4__5 (que_out_13__4__5), .q_4__4 (
            que_out_13__4__4), .q_4__3 (que_out_13__4__3), .q_4__2 (
            que_out_13__4__2), .q_4__1 (que_out_13__4__1), .q_4__0 (
            que_out_13__4__0), .clk (nx10724), .load (sel_que_13), .reset (
            nx10700)) ;
    Queue_5 gen_queues_14_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_14__0__15), .q_0__14 (
            que_out_14__0__14), .q_0__13 (que_out_14__0__13), .q_0__12 (
            que_out_14__0__12), .q_0__11 (que_out_14__0__11), .q_0__10 (
            que_out_14__0__10), .q_0__9 (que_out_14__0__9), .q_0__8 (
            que_out_14__0__8), .q_0__7 (que_out_14__0__7), .q_0__6 (
            que_out_14__0__6), .q_0__5 (que_out_14__0__5), .q_0__4 (
            que_out_14__0__4), .q_0__3 (que_out_14__0__3), .q_0__2 (
            que_out_14__0__2), .q_0__1 (que_out_14__0__1), .q_0__0 (
            que_out_14__0__0), .q_1__15 (que_out_14__1__15), .q_1__14 (
            que_out_14__1__14), .q_1__13 (que_out_14__1__13), .q_1__12 (
            que_out_14__1__12), .q_1__11 (que_out_14__1__11), .q_1__10 (
            que_out_14__1__10), .q_1__9 (que_out_14__1__9), .q_1__8 (
            que_out_14__1__8), .q_1__7 (que_out_14__1__7), .q_1__6 (
            que_out_14__1__6), .q_1__5 (que_out_14__1__5), .q_1__4 (
            que_out_14__1__4), .q_1__3 (que_out_14__1__3), .q_1__2 (
            que_out_14__1__2), .q_1__1 (que_out_14__1__1), .q_1__0 (
            que_out_14__1__0), .q_2__15 (que_out_14__2__15), .q_2__14 (
            que_out_14__2__14), .q_2__13 (que_out_14__2__13), .q_2__12 (
            que_out_14__2__12), .q_2__11 (que_out_14__2__11), .q_2__10 (
            que_out_14__2__10), .q_2__9 (que_out_14__2__9), .q_2__8 (
            que_out_14__2__8), .q_2__7 (que_out_14__2__7), .q_2__6 (
            que_out_14__2__6), .q_2__5 (que_out_14__2__5), .q_2__4 (
            que_out_14__2__4), .q_2__3 (que_out_14__2__3), .q_2__2 (
            que_out_14__2__2), .q_2__1 (que_out_14__2__1), .q_2__0 (
            que_out_14__2__0), .q_3__15 (que_out_14__3__15), .q_3__14 (
            que_out_14__3__14), .q_3__13 (que_out_14__3__13), .q_3__12 (
            que_out_14__3__12), .q_3__11 (que_out_14__3__11), .q_3__10 (
            que_out_14__3__10), .q_3__9 (que_out_14__3__9), .q_3__8 (
            que_out_14__3__8), .q_3__7 (que_out_14__3__7), .q_3__6 (
            que_out_14__3__6), .q_3__5 (que_out_14__3__5), .q_3__4 (
            que_out_14__3__4), .q_3__3 (que_out_14__3__3), .q_3__2 (
            que_out_14__3__2), .q_3__1 (que_out_14__3__1), .q_3__0 (
            que_out_14__3__0), .q_4__15 (que_out_14__4__15), .q_4__14 (
            que_out_14__4__14), .q_4__13 (que_out_14__4__13), .q_4__12 (
            que_out_14__4__12), .q_4__11 (que_out_14__4__11), .q_4__10 (
            que_out_14__4__10), .q_4__9 (que_out_14__4__9), .q_4__8 (
            que_out_14__4__8), .q_4__7 (que_out_14__4__7), .q_4__6 (
            que_out_14__4__6), .q_4__5 (que_out_14__4__5), .q_4__4 (
            que_out_14__4__4), .q_4__3 (que_out_14__4__3), .q_4__2 (
            que_out_14__4__2), .q_4__1 (que_out_14__4__1), .q_4__0 (
            que_out_14__4__0), .clk (nx10726), .load (sel_que_14), .reset (
            nx10702)) ;
    Queue_5 gen_queues_15_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_15__0__15), .q_0__14 (
            que_out_15__0__14), .q_0__13 (que_out_15__0__13), .q_0__12 (
            que_out_15__0__12), .q_0__11 (que_out_15__0__11), .q_0__10 (
            que_out_15__0__10), .q_0__9 (que_out_15__0__9), .q_0__8 (
            que_out_15__0__8), .q_0__7 (que_out_15__0__7), .q_0__6 (
            que_out_15__0__6), .q_0__5 (que_out_15__0__5), .q_0__4 (
            que_out_15__0__4), .q_0__3 (que_out_15__0__3), .q_0__2 (
            que_out_15__0__2), .q_0__1 (que_out_15__0__1), .q_0__0 (
            que_out_15__0__0), .q_1__15 (que_out_15__1__15), .q_1__14 (
            que_out_15__1__14), .q_1__13 (que_out_15__1__13), .q_1__12 (
            que_out_15__1__12), .q_1__11 (que_out_15__1__11), .q_1__10 (
            que_out_15__1__10), .q_1__9 (que_out_15__1__9), .q_1__8 (
            que_out_15__1__8), .q_1__7 (que_out_15__1__7), .q_1__6 (
            que_out_15__1__6), .q_1__5 (que_out_15__1__5), .q_1__4 (
            que_out_15__1__4), .q_1__3 (que_out_15__1__3), .q_1__2 (
            que_out_15__1__2), .q_1__1 (que_out_15__1__1), .q_1__0 (
            que_out_15__1__0), .q_2__15 (que_out_15__2__15), .q_2__14 (
            que_out_15__2__14), .q_2__13 (que_out_15__2__13), .q_2__12 (
            que_out_15__2__12), .q_2__11 (que_out_15__2__11), .q_2__10 (
            que_out_15__2__10), .q_2__9 (que_out_15__2__9), .q_2__8 (
            que_out_15__2__8), .q_2__7 (que_out_15__2__7), .q_2__6 (
            que_out_15__2__6), .q_2__5 (que_out_15__2__5), .q_2__4 (
            que_out_15__2__4), .q_2__3 (que_out_15__2__3), .q_2__2 (
            que_out_15__2__2), .q_2__1 (que_out_15__2__1), .q_2__0 (
            que_out_15__2__0), .q_3__15 (que_out_15__3__15), .q_3__14 (
            que_out_15__3__14), .q_3__13 (que_out_15__3__13), .q_3__12 (
            que_out_15__3__12), .q_3__11 (que_out_15__3__11), .q_3__10 (
            que_out_15__3__10), .q_3__9 (que_out_15__3__9), .q_3__8 (
            que_out_15__3__8), .q_3__7 (que_out_15__3__7), .q_3__6 (
            que_out_15__3__6), .q_3__5 (que_out_15__3__5), .q_3__4 (
            que_out_15__3__4), .q_3__3 (que_out_15__3__3), .q_3__2 (
            que_out_15__3__2), .q_3__1 (que_out_15__3__1), .q_3__0 (
            que_out_15__3__0), .q_4__15 (que_out_15__4__15), .q_4__14 (
            que_out_15__4__14), .q_4__13 (que_out_15__4__13), .q_4__12 (
            que_out_15__4__12), .q_4__11 (que_out_15__4__11), .q_4__10 (
            que_out_15__4__10), .q_4__9 (que_out_15__4__9), .q_4__8 (
            que_out_15__4__8), .q_4__7 (que_out_15__4__7), .q_4__6 (
            que_out_15__4__6), .q_4__5 (que_out_15__4__5), .q_4__4 (
            que_out_15__4__4), .q_4__3 (que_out_15__4__3), .q_4__2 (
            que_out_15__4__2), .q_4__1 (que_out_15__4__1), .q_4__0 (
            que_out_15__4__0), .clk (nx10726), .load (sel_que_15), .reset (
            nx10702)) ;
    Queue_5 gen_queues_16_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_16__0__15), .q_0__14 (
            que_out_16__0__14), .q_0__13 (que_out_16__0__13), .q_0__12 (
            que_out_16__0__12), .q_0__11 (que_out_16__0__11), .q_0__10 (
            que_out_16__0__10), .q_0__9 (que_out_16__0__9), .q_0__8 (
            que_out_16__0__8), .q_0__7 (que_out_16__0__7), .q_0__6 (
            que_out_16__0__6), .q_0__5 (que_out_16__0__5), .q_0__4 (
            que_out_16__0__4), .q_0__3 (que_out_16__0__3), .q_0__2 (
            que_out_16__0__2), .q_0__1 (que_out_16__0__1), .q_0__0 (
            que_out_16__0__0), .q_1__15 (que_out_16__1__15), .q_1__14 (
            que_out_16__1__14), .q_1__13 (que_out_16__1__13), .q_1__12 (
            que_out_16__1__12), .q_1__11 (que_out_16__1__11), .q_1__10 (
            que_out_16__1__10), .q_1__9 (que_out_16__1__9), .q_1__8 (
            que_out_16__1__8), .q_1__7 (que_out_16__1__7), .q_1__6 (
            que_out_16__1__6), .q_1__5 (que_out_16__1__5), .q_1__4 (
            que_out_16__1__4), .q_1__3 (que_out_16__1__3), .q_1__2 (
            que_out_16__1__2), .q_1__1 (que_out_16__1__1), .q_1__0 (
            que_out_16__1__0), .q_2__15 (que_out_16__2__15), .q_2__14 (
            que_out_16__2__14), .q_2__13 (que_out_16__2__13), .q_2__12 (
            que_out_16__2__12), .q_2__11 (que_out_16__2__11), .q_2__10 (
            que_out_16__2__10), .q_2__9 (que_out_16__2__9), .q_2__8 (
            que_out_16__2__8), .q_2__7 (que_out_16__2__7), .q_2__6 (
            que_out_16__2__6), .q_2__5 (que_out_16__2__5), .q_2__4 (
            que_out_16__2__4), .q_2__3 (que_out_16__2__3), .q_2__2 (
            que_out_16__2__2), .q_2__1 (que_out_16__2__1), .q_2__0 (
            que_out_16__2__0), .q_3__15 (que_out_16__3__15), .q_3__14 (
            que_out_16__3__14), .q_3__13 (que_out_16__3__13), .q_3__12 (
            que_out_16__3__12), .q_3__11 (que_out_16__3__11), .q_3__10 (
            que_out_16__3__10), .q_3__9 (que_out_16__3__9), .q_3__8 (
            que_out_16__3__8), .q_3__7 (que_out_16__3__7), .q_3__6 (
            que_out_16__3__6), .q_3__5 (que_out_16__3__5), .q_3__4 (
            que_out_16__3__4), .q_3__3 (que_out_16__3__3), .q_3__2 (
            que_out_16__3__2), .q_3__1 (que_out_16__3__1), .q_3__0 (
            que_out_16__3__0), .q_4__15 (que_out_16__4__15), .q_4__14 (
            que_out_16__4__14), .q_4__13 (que_out_16__4__13), .q_4__12 (
            que_out_16__4__12), .q_4__11 (que_out_16__4__11), .q_4__10 (
            que_out_16__4__10), .q_4__9 (que_out_16__4__9), .q_4__8 (
            que_out_16__4__8), .q_4__7 (que_out_16__4__7), .q_4__6 (
            que_out_16__4__6), .q_4__5 (que_out_16__4__5), .q_4__4 (
            que_out_16__4__4), .q_4__3 (que_out_16__4__3), .q_4__2 (
            que_out_16__4__2), .q_4__1 (que_out_16__4__1), .q_4__0 (
            que_out_16__4__0), .clk (nx10726), .load (sel_que_16), .reset (
            nx10702)) ;
    Queue_5 gen_queues_17_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_17__0__15), .q_0__14 (
            que_out_17__0__14), .q_0__13 (que_out_17__0__13), .q_0__12 (
            que_out_17__0__12), .q_0__11 (que_out_17__0__11), .q_0__10 (
            que_out_17__0__10), .q_0__9 (que_out_17__0__9), .q_0__8 (
            que_out_17__0__8), .q_0__7 (que_out_17__0__7), .q_0__6 (
            que_out_17__0__6), .q_0__5 (que_out_17__0__5), .q_0__4 (
            que_out_17__0__4), .q_0__3 (que_out_17__0__3), .q_0__2 (
            que_out_17__0__2), .q_0__1 (que_out_17__0__1), .q_0__0 (
            que_out_17__0__0), .q_1__15 (que_out_17__1__15), .q_1__14 (
            que_out_17__1__14), .q_1__13 (que_out_17__1__13), .q_1__12 (
            que_out_17__1__12), .q_1__11 (que_out_17__1__11), .q_1__10 (
            que_out_17__1__10), .q_1__9 (que_out_17__1__9), .q_1__8 (
            que_out_17__1__8), .q_1__7 (que_out_17__1__7), .q_1__6 (
            que_out_17__1__6), .q_1__5 (que_out_17__1__5), .q_1__4 (
            que_out_17__1__4), .q_1__3 (que_out_17__1__3), .q_1__2 (
            que_out_17__1__2), .q_1__1 (que_out_17__1__1), .q_1__0 (
            que_out_17__1__0), .q_2__15 (que_out_17__2__15), .q_2__14 (
            que_out_17__2__14), .q_2__13 (que_out_17__2__13), .q_2__12 (
            que_out_17__2__12), .q_2__11 (que_out_17__2__11), .q_2__10 (
            que_out_17__2__10), .q_2__9 (que_out_17__2__9), .q_2__8 (
            que_out_17__2__8), .q_2__7 (que_out_17__2__7), .q_2__6 (
            que_out_17__2__6), .q_2__5 (que_out_17__2__5), .q_2__4 (
            que_out_17__2__4), .q_2__3 (que_out_17__2__3), .q_2__2 (
            que_out_17__2__2), .q_2__1 (que_out_17__2__1), .q_2__0 (
            que_out_17__2__0), .q_3__15 (que_out_17__3__15), .q_3__14 (
            que_out_17__3__14), .q_3__13 (que_out_17__3__13), .q_3__12 (
            que_out_17__3__12), .q_3__11 (que_out_17__3__11), .q_3__10 (
            que_out_17__3__10), .q_3__9 (que_out_17__3__9), .q_3__8 (
            que_out_17__3__8), .q_3__7 (que_out_17__3__7), .q_3__6 (
            que_out_17__3__6), .q_3__5 (que_out_17__3__5), .q_3__4 (
            que_out_17__3__4), .q_3__3 (que_out_17__3__3), .q_3__2 (
            que_out_17__3__2), .q_3__1 (que_out_17__3__1), .q_3__0 (
            que_out_17__3__0), .q_4__15 (que_out_17__4__15), .q_4__14 (
            que_out_17__4__14), .q_4__13 (que_out_17__4__13), .q_4__12 (
            que_out_17__4__12), .q_4__11 (que_out_17__4__11), .q_4__10 (
            que_out_17__4__10), .q_4__9 (que_out_17__4__9), .q_4__8 (
            que_out_17__4__8), .q_4__7 (que_out_17__4__7), .q_4__6 (
            que_out_17__4__6), .q_4__5 (que_out_17__4__5), .q_4__4 (
            que_out_17__4__4), .q_4__3 (que_out_17__4__3), .q_4__2 (
            que_out_17__4__2), .q_4__1 (que_out_17__4__1), .q_4__0 (
            que_out_17__4__0), .clk (nx10728), .load (sel_que_17), .reset (
            nx10704)) ;
    Queue_5 gen_queues_18_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_18__0__15), .q_0__14 (
            que_out_18__0__14), .q_0__13 (que_out_18__0__13), .q_0__12 (
            que_out_18__0__12), .q_0__11 (que_out_18__0__11), .q_0__10 (
            que_out_18__0__10), .q_0__9 (que_out_18__0__9), .q_0__8 (
            que_out_18__0__8), .q_0__7 (que_out_18__0__7), .q_0__6 (
            que_out_18__0__6), .q_0__5 (que_out_18__0__5), .q_0__4 (
            que_out_18__0__4), .q_0__3 (que_out_18__0__3), .q_0__2 (
            que_out_18__0__2), .q_0__1 (que_out_18__0__1), .q_0__0 (
            que_out_18__0__0), .q_1__15 (que_out_18__1__15), .q_1__14 (
            que_out_18__1__14), .q_1__13 (que_out_18__1__13), .q_1__12 (
            que_out_18__1__12), .q_1__11 (que_out_18__1__11), .q_1__10 (
            que_out_18__1__10), .q_1__9 (que_out_18__1__9), .q_1__8 (
            que_out_18__1__8), .q_1__7 (que_out_18__1__7), .q_1__6 (
            que_out_18__1__6), .q_1__5 (que_out_18__1__5), .q_1__4 (
            que_out_18__1__4), .q_1__3 (que_out_18__1__3), .q_1__2 (
            que_out_18__1__2), .q_1__1 (que_out_18__1__1), .q_1__0 (
            que_out_18__1__0), .q_2__15 (que_out_18__2__15), .q_2__14 (
            que_out_18__2__14), .q_2__13 (que_out_18__2__13), .q_2__12 (
            que_out_18__2__12), .q_2__11 (que_out_18__2__11), .q_2__10 (
            que_out_18__2__10), .q_2__9 (que_out_18__2__9), .q_2__8 (
            que_out_18__2__8), .q_2__7 (que_out_18__2__7), .q_2__6 (
            que_out_18__2__6), .q_2__5 (que_out_18__2__5), .q_2__4 (
            que_out_18__2__4), .q_2__3 (que_out_18__2__3), .q_2__2 (
            que_out_18__2__2), .q_2__1 (que_out_18__2__1), .q_2__0 (
            que_out_18__2__0), .q_3__15 (que_out_18__3__15), .q_3__14 (
            que_out_18__3__14), .q_3__13 (que_out_18__3__13), .q_3__12 (
            que_out_18__3__12), .q_3__11 (que_out_18__3__11), .q_3__10 (
            que_out_18__3__10), .q_3__9 (que_out_18__3__9), .q_3__8 (
            que_out_18__3__8), .q_3__7 (que_out_18__3__7), .q_3__6 (
            que_out_18__3__6), .q_3__5 (que_out_18__3__5), .q_3__4 (
            que_out_18__3__4), .q_3__3 (que_out_18__3__3), .q_3__2 (
            que_out_18__3__2), .q_3__1 (que_out_18__3__1), .q_3__0 (
            que_out_18__3__0), .q_4__15 (que_out_18__4__15), .q_4__14 (
            que_out_18__4__14), .q_4__13 (que_out_18__4__13), .q_4__12 (
            que_out_18__4__12), .q_4__11 (que_out_18__4__11), .q_4__10 (
            que_out_18__4__10), .q_4__9 (que_out_18__4__9), .q_4__8 (
            que_out_18__4__8), .q_4__7 (que_out_18__4__7), .q_4__6 (
            que_out_18__4__6), .q_4__5 (que_out_18__4__5), .q_4__4 (
            que_out_18__4__4), .q_4__3 (que_out_18__4__3), .q_4__2 (
            que_out_18__4__2), .q_4__1 (que_out_18__4__1), .q_4__0 (
            que_out_18__4__0), .clk (nx10728), .load (sel_que_18), .reset (
            nx10704)) ;
    Queue_5 gen_queues_19_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_19__0__15), .q_0__14 (
            que_out_19__0__14), .q_0__13 (que_out_19__0__13), .q_0__12 (
            que_out_19__0__12), .q_0__11 (que_out_19__0__11), .q_0__10 (
            que_out_19__0__10), .q_0__9 (que_out_19__0__9), .q_0__8 (
            que_out_19__0__8), .q_0__7 (que_out_19__0__7), .q_0__6 (
            que_out_19__0__6), .q_0__5 (que_out_19__0__5), .q_0__4 (
            que_out_19__0__4), .q_0__3 (que_out_19__0__3), .q_0__2 (
            que_out_19__0__2), .q_0__1 (que_out_19__0__1), .q_0__0 (
            que_out_19__0__0), .q_1__15 (que_out_19__1__15), .q_1__14 (
            que_out_19__1__14), .q_1__13 (que_out_19__1__13), .q_1__12 (
            que_out_19__1__12), .q_1__11 (que_out_19__1__11), .q_1__10 (
            que_out_19__1__10), .q_1__9 (que_out_19__1__9), .q_1__8 (
            que_out_19__1__8), .q_1__7 (que_out_19__1__7), .q_1__6 (
            que_out_19__1__6), .q_1__5 (que_out_19__1__5), .q_1__4 (
            que_out_19__1__4), .q_1__3 (que_out_19__1__3), .q_1__2 (
            que_out_19__1__2), .q_1__1 (que_out_19__1__1), .q_1__0 (
            que_out_19__1__0), .q_2__15 (que_out_19__2__15), .q_2__14 (
            que_out_19__2__14), .q_2__13 (que_out_19__2__13), .q_2__12 (
            que_out_19__2__12), .q_2__11 (que_out_19__2__11), .q_2__10 (
            que_out_19__2__10), .q_2__9 (que_out_19__2__9), .q_2__8 (
            que_out_19__2__8), .q_2__7 (que_out_19__2__7), .q_2__6 (
            que_out_19__2__6), .q_2__5 (que_out_19__2__5), .q_2__4 (
            que_out_19__2__4), .q_2__3 (que_out_19__2__3), .q_2__2 (
            que_out_19__2__2), .q_2__1 (que_out_19__2__1), .q_2__0 (
            que_out_19__2__0), .q_3__15 (que_out_19__3__15), .q_3__14 (
            que_out_19__3__14), .q_3__13 (que_out_19__3__13), .q_3__12 (
            que_out_19__3__12), .q_3__11 (que_out_19__3__11), .q_3__10 (
            que_out_19__3__10), .q_3__9 (que_out_19__3__9), .q_3__8 (
            que_out_19__3__8), .q_3__7 (que_out_19__3__7), .q_3__6 (
            que_out_19__3__6), .q_3__5 (que_out_19__3__5), .q_3__4 (
            que_out_19__3__4), .q_3__3 (que_out_19__3__3), .q_3__2 (
            que_out_19__3__2), .q_3__1 (que_out_19__3__1), .q_3__0 (
            que_out_19__3__0), .q_4__15 (que_out_19__4__15), .q_4__14 (
            que_out_19__4__14), .q_4__13 (que_out_19__4__13), .q_4__12 (
            que_out_19__4__12), .q_4__11 (que_out_19__4__11), .q_4__10 (
            que_out_19__4__10), .q_4__9 (que_out_19__4__9), .q_4__8 (
            que_out_19__4__8), .q_4__7 (que_out_19__4__7), .q_4__6 (
            que_out_19__4__6), .q_4__5 (que_out_19__4__5), .q_4__4 (
            que_out_19__4__4), .q_4__3 (que_out_19__4__3), .q_4__2 (
            que_out_19__4__2), .q_4__1 (que_out_19__4__1), .q_4__0 (
            que_out_19__4__0), .clk (nx10728), .load (sel_que_19), .reset (
            nx10704)) ;
    Queue_5 gen_queues_20_que (.d ({nx10516,nx10526,nx10536,nx10546,nx10556,
            nx10566,nx10576,nx10586,nx10596,nx10606,nx10616,nx10626,nx10636,
            nx10646,nx10656,nx10666}), .q_0__15 (que_out_20__0__15), .q_0__14 (
            que_out_20__0__14), .q_0__13 (que_out_20__0__13), .q_0__12 (
            que_out_20__0__12), .q_0__11 (que_out_20__0__11), .q_0__10 (
            que_out_20__0__10), .q_0__9 (que_out_20__0__9), .q_0__8 (
            que_out_20__0__8), .q_0__7 (que_out_20__0__7), .q_0__6 (
            que_out_20__0__6), .q_0__5 (que_out_20__0__5), .q_0__4 (
            que_out_20__0__4), .q_0__3 (que_out_20__0__3), .q_0__2 (
            que_out_20__0__2), .q_0__1 (que_out_20__0__1), .q_0__0 (
            que_out_20__0__0), .q_1__15 (que_out_20__1__15), .q_1__14 (
            que_out_20__1__14), .q_1__13 (que_out_20__1__13), .q_1__12 (
            que_out_20__1__12), .q_1__11 (que_out_20__1__11), .q_1__10 (
            que_out_20__1__10), .q_1__9 (que_out_20__1__9), .q_1__8 (
            que_out_20__1__8), .q_1__7 (que_out_20__1__7), .q_1__6 (
            que_out_20__1__6), .q_1__5 (que_out_20__1__5), .q_1__4 (
            que_out_20__1__4), .q_1__3 (que_out_20__1__3), .q_1__2 (
            que_out_20__1__2), .q_1__1 (que_out_20__1__1), .q_1__0 (
            que_out_20__1__0), .q_2__15 (que_out_20__2__15), .q_2__14 (
            que_out_20__2__14), .q_2__13 (que_out_20__2__13), .q_2__12 (
            que_out_20__2__12), .q_2__11 (que_out_20__2__11), .q_2__10 (
            que_out_20__2__10), .q_2__9 (que_out_20__2__9), .q_2__8 (
            que_out_20__2__8), .q_2__7 (que_out_20__2__7), .q_2__6 (
            que_out_20__2__6), .q_2__5 (que_out_20__2__5), .q_2__4 (
            que_out_20__2__4), .q_2__3 (que_out_20__2__3), .q_2__2 (
            que_out_20__2__2), .q_2__1 (que_out_20__2__1), .q_2__0 (
            que_out_20__2__0), .q_3__15 (que_out_20__3__15), .q_3__14 (
            que_out_20__3__14), .q_3__13 (que_out_20__3__13), .q_3__12 (
            que_out_20__3__12), .q_3__11 (que_out_20__3__11), .q_3__10 (
            que_out_20__3__10), .q_3__9 (que_out_20__3__9), .q_3__8 (
            que_out_20__3__8), .q_3__7 (que_out_20__3__7), .q_3__6 (
            que_out_20__3__6), .q_3__5 (que_out_20__3__5), .q_3__4 (
            que_out_20__3__4), .q_3__3 (que_out_20__3__3), .q_3__2 (
            que_out_20__3__2), .q_3__1 (que_out_20__3__1), .q_3__0 (
            que_out_20__3__0), .q_4__15 (que_out_20__4__15), .q_4__14 (
            que_out_20__4__14), .q_4__13 (que_out_20__4__13), .q_4__12 (
            que_out_20__4__12), .q_4__11 (que_out_20__4__11), .q_4__10 (
            que_out_20__4__10), .q_4__9 (que_out_20__4__9), .q_4__8 (
            que_out_20__4__8), .q_4__7 (que_out_20__4__7), .q_4__6 (
            que_out_20__4__6), .q_4__5 (que_out_20__4__5), .q_4__4 (
            que_out_20__4__4), .q_4__3 (que_out_20__4__3), .q_4__2 (
            que_out_20__4__2), .q_4__1 (que_out_20__4__1), .q_4__0 (
            que_out_20__4__0), .clk (nx10730), .load (sel_que_20), .reset (
            nx10706)) ;
    Queue_5 gen_queues_21_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_21__0__15), .q_0__14 (
            que_out_21__0__14), .q_0__13 (que_out_21__0__13), .q_0__12 (
            que_out_21__0__12), .q_0__11 (que_out_21__0__11), .q_0__10 (
            que_out_21__0__10), .q_0__9 (que_out_21__0__9), .q_0__8 (
            que_out_21__0__8), .q_0__7 (que_out_21__0__7), .q_0__6 (
            que_out_21__0__6), .q_0__5 (que_out_21__0__5), .q_0__4 (
            que_out_21__0__4), .q_0__3 (que_out_21__0__3), .q_0__2 (
            que_out_21__0__2), .q_0__1 (que_out_21__0__1), .q_0__0 (
            que_out_21__0__0), .q_1__15 (que_out_21__1__15), .q_1__14 (
            que_out_21__1__14), .q_1__13 (que_out_21__1__13), .q_1__12 (
            que_out_21__1__12), .q_1__11 (que_out_21__1__11), .q_1__10 (
            que_out_21__1__10), .q_1__9 (que_out_21__1__9), .q_1__8 (
            que_out_21__1__8), .q_1__7 (que_out_21__1__7), .q_1__6 (
            que_out_21__1__6), .q_1__5 (que_out_21__1__5), .q_1__4 (
            que_out_21__1__4), .q_1__3 (que_out_21__1__3), .q_1__2 (
            que_out_21__1__2), .q_1__1 (que_out_21__1__1), .q_1__0 (
            que_out_21__1__0), .q_2__15 (que_out_21__2__15), .q_2__14 (
            que_out_21__2__14), .q_2__13 (que_out_21__2__13), .q_2__12 (
            que_out_21__2__12), .q_2__11 (que_out_21__2__11), .q_2__10 (
            que_out_21__2__10), .q_2__9 (que_out_21__2__9), .q_2__8 (
            que_out_21__2__8), .q_2__7 (que_out_21__2__7), .q_2__6 (
            que_out_21__2__6), .q_2__5 (que_out_21__2__5), .q_2__4 (
            que_out_21__2__4), .q_2__3 (que_out_21__2__3), .q_2__2 (
            que_out_21__2__2), .q_2__1 (que_out_21__2__1), .q_2__0 (
            que_out_21__2__0), .q_3__15 (que_out_21__3__15), .q_3__14 (
            que_out_21__3__14), .q_3__13 (que_out_21__3__13), .q_3__12 (
            que_out_21__3__12), .q_3__11 (que_out_21__3__11), .q_3__10 (
            que_out_21__3__10), .q_3__9 (que_out_21__3__9), .q_3__8 (
            que_out_21__3__8), .q_3__7 (que_out_21__3__7), .q_3__6 (
            que_out_21__3__6), .q_3__5 (que_out_21__3__5), .q_3__4 (
            que_out_21__3__4), .q_3__3 (que_out_21__3__3), .q_3__2 (
            que_out_21__3__2), .q_3__1 (que_out_21__3__1), .q_3__0 (
            que_out_21__3__0), .q_4__15 (que_out_21__4__15), .q_4__14 (
            que_out_21__4__14), .q_4__13 (que_out_21__4__13), .q_4__12 (
            que_out_21__4__12), .q_4__11 (que_out_21__4__11), .q_4__10 (
            que_out_21__4__10), .q_4__9 (que_out_21__4__9), .q_4__8 (
            que_out_21__4__8), .q_4__7 (que_out_21__4__7), .q_4__6 (
            que_out_21__4__6), .q_4__5 (que_out_21__4__5), .q_4__4 (
            que_out_21__4__4), .q_4__3 (que_out_21__4__3), .q_4__2 (
            que_out_21__4__2), .q_4__1 (que_out_21__4__1), .q_4__0 (
            que_out_21__4__0), .clk (nx10732), .load (sel_que_21), .reset (
            nx10708)) ;
    Queue_5 gen_queues_22_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_22__0__15), .q_0__14 (
            que_out_22__0__14), .q_0__13 (que_out_22__0__13), .q_0__12 (
            que_out_22__0__12), .q_0__11 (que_out_22__0__11), .q_0__10 (
            que_out_22__0__10), .q_0__9 (que_out_22__0__9), .q_0__8 (
            que_out_22__0__8), .q_0__7 (que_out_22__0__7), .q_0__6 (
            que_out_22__0__6), .q_0__5 (que_out_22__0__5), .q_0__4 (
            que_out_22__0__4), .q_0__3 (que_out_22__0__3), .q_0__2 (
            que_out_22__0__2), .q_0__1 (que_out_22__0__1), .q_0__0 (
            que_out_22__0__0), .q_1__15 (que_out_22__1__15), .q_1__14 (
            que_out_22__1__14), .q_1__13 (que_out_22__1__13), .q_1__12 (
            que_out_22__1__12), .q_1__11 (que_out_22__1__11), .q_1__10 (
            que_out_22__1__10), .q_1__9 (que_out_22__1__9), .q_1__8 (
            que_out_22__1__8), .q_1__7 (que_out_22__1__7), .q_1__6 (
            que_out_22__1__6), .q_1__5 (que_out_22__1__5), .q_1__4 (
            que_out_22__1__4), .q_1__3 (que_out_22__1__3), .q_1__2 (
            que_out_22__1__2), .q_1__1 (que_out_22__1__1), .q_1__0 (
            que_out_22__1__0), .q_2__15 (que_out_22__2__15), .q_2__14 (
            que_out_22__2__14), .q_2__13 (que_out_22__2__13), .q_2__12 (
            que_out_22__2__12), .q_2__11 (que_out_22__2__11), .q_2__10 (
            que_out_22__2__10), .q_2__9 (que_out_22__2__9), .q_2__8 (
            que_out_22__2__8), .q_2__7 (que_out_22__2__7), .q_2__6 (
            que_out_22__2__6), .q_2__5 (que_out_22__2__5), .q_2__4 (
            que_out_22__2__4), .q_2__3 (que_out_22__2__3), .q_2__2 (
            que_out_22__2__2), .q_2__1 (que_out_22__2__1), .q_2__0 (
            que_out_22__2__0), .q_3__15 (que_out_22__3__15), .q_3__14 (
            que_out_22__3__14), .q_3__13 (que_out_22__3__13), .q_3__12 (
            que_out_22__3__12), .q_3__11 (que_out_22__3__11), .q_3__10 (
            que_out_22__3__10), .q_3__9 (que_out_22__3__9), .q_3__8 (
            que_out_22__3__8), .q_3__7 (que_out_22__3__7), .q_3__6 (
            que_out_22__3__6), .q_3__5 (que_out_22__3__5), .q_3__4 (
            que_out_22__3__4), .q_3__3 (que_out_22__3__3), .q_3__2 (
            que_out_22__3__2), .q_3__1 (que_out_22__3__1), .q_3__0 (
            que_out_22__3__0), .q_4__15 (que_out_22__4__15), .q_4__14 (
            que_out_22__4__14), .q_4__13 (que_out_22__4__13), .q_4__12 (
            que_out_22__4__12), .q_4__11 (que_out_22__4__11), .q_4__10 (
            que_out_22__4__10), .q_4__9 (que_out_22__4__9), .q_4__8 (
            que_out_22__4__8), .q_4__7 (que_out_22__4__7), .q_4__6 (
            que_out_22__4__6), .q_4__5 (que_out_22__4__5), .q_4__4 (
            que_out_22__4__4), .q_4__3 (que_out_22__4__3), .q_4__2 (
            que_out_22__4__2), .q_4__1 (que_out_22__4__1), .q_4__0 (
            que_out_22__4__0), .clk (nx10732), .load (sel_que_22), .reset (
            nx10708)) ;
    Queue_5 gen_queues_23_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_23__0__15), .q_0__14 (
            que_out_23__0__14), .q_0__13 (que_out_23__0__13), .q_0__12 (
            que_out_23__0__12), .q_0__11 (que_out_23__0__11), .q_0__10 (
            que_out_23__0__10), .q_0__9 (que_out_23__0__9), .q_0__8 (
            que_out_23__0__8), .q_0__7 (que_out_23__0__7), .q_0__6 (
            que_out_23__0__6), .q_0__5 (que_out_23__0__5), .q_0__4 (
            que_out_23__0__4), .q_0__3 (que_out_23__0__3), .q_0__2 (
            que_out_23__0__2), .q_0__1 (que_out_23__0__1), .q_0__0 (
            que_out_23__0__0), .q_1__15 (que_out_23__1__15), .q_1__14 (
            que_out_23__1__14), .q_1__13 (que_out_23__1__13), .q_1__12 (
            que_out_23__1__12), .q_1__11 (que_out_23__1__11), .q_1__10 (
            que_out_23__1__10), .q_1__9 (que_out_23__1__9), .q_1__8 (
            que_out_23__1__8), .q_1__7 (que_out_23__1__7), .q_1__6 (
            que_out_23__1__6), .q_1__5 (que_out_23__1__5), .q_1__4 (
            que_out_23__1__4), .q_1__3 (que_out_23__1__3), .q_1__2 (
            que_out_23__1__2), .q_1__1 (que_out_23__1__1), .q_1__0 (
            que_out_23__1__0), .q_2__15 (que_out_23__2__15), .q_2__14 (
            que_out_23__2__14), .q_2__13 (que_out_23__2__13), .q_2__12 (
            que_out_23__2__12), .q_2__11 (que_out_23__2__11), .q_2__10 (
            que_out_23__2__10), .q_2__9 (que_out_23__2__9), .q_2__8 (
            que_out_23__2__8), .q_2__7 (que_out_23__2__7), .q_2__6 (
            que_out_23__2__6), .q_2__5 (que_out_23__2__5), .q_2__4 (
            que_out_23__2__4), .q_2__3 (que_out_23__2__3), .q_2__2 (
            que_out_23__2__2), .q_2__1 (que_out_23__2__1), .q_2__0 (
            que_out_23__2__0), .q_3__15 (que_out_23__3__15), .q_3__14 (
            que_out_23__3__14), .q_3__13 (que_out_23__3__13), .q_3__12 (
            que_out_23__3__12), .q_3__11 (que_out_23__3__11), .q_3__10 (
            que_out_23__3__10), .q_3__9 (que_out_23__3__9), .q_3__8 (
            que_out_23__3__8), .q_3__7 (que_out_23__3__7), .q_3__6 (
            que_out_23__3__6), .q_3__5 (que_out_23__3__5), .q_3__4 (
            que_out_23__3__4), .q_3__3 (que_out_23__3__3), .q_3__2 (
            que_out_23__3__2), .q_3__1 (que_out_23__3__1), .q_3__0 (
            que_out_23__3__0), .q_4__15 (que_out_23__4__15), .q_4__14 (
            que_out_23__4__14), .q_4__13 (que_out_23__4__13), .q_4__12 (
            que_out_23__4__12), .q_4__11 (que_out_23__4__11), .q_4__10 (
            que_out_23__4__10), .q_4__9 (que_out_23__4__9), .q_4__8 (
            que_out_23__4__8), .q_4__7 (que_out_23__4__7), .q_4__6 (
            que_out_23__4__6), .q_4__5 (que_out_23__4__5), .q_4__4 (
            que_out_23__4__4), .q_4__3 (que_out_23__4__3), .q_4__2 (
            que_out_23__4__2), .q_4__1 (que_out_23__4__1), .q_4__0 (
            que_out_23__4__0), .clk (nx10732), .load (sel_que_23), .reset (
            nx10708)) ;
    Queue_5 gen_queues_24_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_24__0__15), .q_0__14 (
            que_out_24__0__14), .q_0__13 (que_out_24__0__13), .q_0__12 (
            que_out_24__0__12), .q_0__11 (que_out_24__0__11), .q_0__10 (
            que_out_24__0__10), .q_0__9 (que_out_24__0__9), .q_0__8 (
            que_out_24__0__8), .q_0__7 (que_out_24__0__7), .q_0__6 (
            que_out_24__0__6), .q_0__5 (que_out_24__0__5), .q_0__4 (
            que_out_24__0__4), .q_0__3 (que_out_24__0__3), .q_0__2 (
            que_out_24__0__2), .q_0__1 (que_out_24__0__1), .q_0__0 (
            que_out_24__0__0), .q_1__15 (que_out_24__1__15), .q_1__14 (
            que_out_24__1__14), .q_1__13 (que_out_24__1__13), .q_1__12 (
            que_out_24__1__12), .q_1__11 (que_out_24__1__11), .q_1__10 (
            que_out_24__1__10), .q_1__9 (que_out_24__1__9), .q_1__8 (
            que_out_24__1__8), .q_1__7 (que_out_24__1__7), .q_1__6 (
            que_out_24__1__6), .q_1__5 (que_out_24__1__5), .q_1__4 (
            que_out_24__1__4), .q_1__3 (que_out_24__1__3), .q_1__2 (
            que_out_24__1__2), .q_1__1 (que_out_24__1__1), .q_1__0 (
            que_out_24__1__0), .q_2__15 (que_out_24__2__15), .q_2__14 (
            que_out_24__2__14), .q_2__13 (que_out_24__2__13), .q_2__12 (
            que_out_24__2__12), .q_2__11 (que_out_24__2__11), .q_2__10 (
            que_out_24__2__10), .q_2__9 (que_out_24__2__9), .q_2__8 (
            que_out_24__2__8), .q_2__7 (que_out_24__2__7), .q_2__6 (
            que_out_24__2__6), .q_2__5 (que_out_24__2__5), .q_2__4 (
            que_out_24__2__4), .q_2__3 (que_out_24__2__3), .q_2__2 (
            que_out_24__2__2), .q_2__1 (que_out_24__2__1), .q_2__0 (
            que_out_24__2__0), .q_3__15 (que_out_24__3__15), .q_3__14 (
            que_out_24__3__14), .q_3__13 (que_out_24__3__13), .q_3__12 (
            que_out_24__3__12), .q_3__11 (que_out_24__3__11), .q_3__10 (
            que_out_24__3__10), .q_3__9 (que_out_24__3__9), .q_3__8 (
            que_out_24__3__8), .q_3__7 (que_out_24__3__7), .q_3__6 (
            que_out_24__3__6), .q_3__5 (que_out_24__3__5), .q_3__4 (
            que_out_24__3__4), .q_3__3 (que_out_24__3__3), .q_3__2 (
            que_out_24__3__2), .q_3__1 (que_out_24__3__1), .q_3__0 (
            que_out_24__3__0), .q_4__15 (que_out_24__4__15), .q_4__14 (
            que_out_24__4__14), .q_4__13 (que_out_24__4__13), .q_4__12 (
            que_out_24__4__12), .q_4__11 (que_out_24__4__11), .q_4__10 (
            que_out_24__4__10), .q_4__9 (que_out_24__4__9), .q_4__8 (
            que_out_24__4__8), .q_4__7 (que_out_24__4__7), .q_4__6 (
            que_out_24__4__6), .q_4__5 (que_out_24__4__5), .q_4__4 (
            que_out_24__4__4), .q_4__3 (que_out_24__4__3), .q_4__2 (
            que_out_24__4__2), .q_4__1 (que_out_24__4__1), .q_4__0 (
            que_out_24__4__0), .clk (nx10734), .load (sel_que_24), .reset (
            nx10710)) ;
    Queue_5 gen_queues_25_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_25__0__15), .q_0__14 (
            que_out_25__0__14), .q_0__13 (que_out_25__0__13), .q_0__12 (
            que_out_25__0__12), .q_0__11 (que_out_25__0__11), .q_0__10 (
            que_out_25__0__10), .q_0__9 (que_out_25__0__9), .q_0__8 (
            que_out_25__0__8), .q_0__7 (que_out_25__0__7), .q_0__6 (
            que_out_25__0__6), .q_0__5 (que_out_25__0__5), .q_0__4 (
            que_out_25__0__4), .q_0__3 (que_out_25__0__3), .q_0__2 (
            que_out_25__0__2), .q_0__1 (que_out_25__0__1), .q_0__0 (
            que_out_25__0__0), .q_1__15 (que_out_25__1__15), .q_1__14 (
            que_out_25__1__14), .q_1__13 (que_out_25__1__13), .q_1__12 (
            que_out_25__1__12), .q_1__11 (que_out_25__1__11), .q_1__10 (
            que_out_25__1__10), .q_1__9 (que_out_25__1__9), .q_1__8 (
            que_out_25__1__8), .q_1__7 (que_out_25__1__7), .q_1__6 (
            que_out_25__1__6), .q_1__5 (que_out_25__1__5), .q_1__4 (
            que_out_25__1__4), .q_1__3 (que_out_25__1__3), .q_1__2 (
            que_out_25__1__2), .q_1__1 (que_out_25__1__1), .q_1__0 (
            que_out_25__1__0), .q_2__15 (que_out_25__2__15), .q_2__14 (
            que_out_25__2__14), .q_2__13 (que_out_25__2__13), .q_2__12 (
            que_out_25__2__12), .q_2__11 (que_out_25__2__11), .q_2__10 (
            que_out_25__2__10), .q_2__9 (que_out_25__2__9), .q_2__8 (
            que_out_25__2__8), .q_2__7 (que_out_25__2__7), .q_2__6 (
            que_out_25__2__6), .q_2__5 (que_out_25__2__5), .q_2__4 (
            que_out_25__2__4), .q_2__3 (que_out_25__2__3), .q_2__2 (
            que_out_25__2__2), .q_2__1 (que_out_25__2__1), .q_2__0 (
            que_out_25__2__0), .q_3__15 (que_out_25__3__15), .q_3__14 (
            que_out_25__3__14), .q_3__13 (que_out_25__3__13), .q_3__12 (
            que_out_25__3__12), .q_3__11 (que_out_25__3__11), .q_3__10 (
            que_out_25__3__10), .q_3__9 (que_out_25__3__9), .q_3__8 (
            que_out_25__3__8), .q_3__7 (que_out_25__3__7), .q_3__6 (
            que_out_25__3__6), .q_3__5 (que_out_25__3__5), .q_3__4 (
            que_out_25__3__4), .q_3__3 (que_out_25__3__3), .q_3__2 (
            que_out_25__3__2), .q_3__1 (que_out_25__3__1), .q_3__0 (
            que_out_25__3__0), .q_4__15 (que_out_25__4__15), .q_4__14 (
            que_out_25__4__14), .q_4__13 (que_out_25__4__13), .q_4__12 (
            que_out_25__4__12), .q_4__11 (que_out_25__4__11), .q_4__10 (
            que_out_25__4__10), .q_4__9 (que_out_25__4__9), .q_4__8 (
            que_out_25__4__8), .q_4__7 (que_out_25__4__7), .q_4__6 (
            que_out_25__4__6), .q_4__5 (que_out_25__4__5), .q_4__4 (
            que_out_25__4__4), .q_4__3 (que_out_25__4__3), .q_4__2 (
            que_out_25__4__2), .q_4__1 (que_out_25__4__1), .q_4__0 (
            que_out_25__4__0), .clk (nx10734), .load (sel_que_25), .reset (
            nx10710)) ;
    Queue_5 gen_queues_26_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_26__0__15), .q_0__14 (
            que_out_26__0__14), .q_0__13 (que_out_26__0__13), .q_0__12 (
            que_out_26__0__12), .q_0__11 (que_out_26__0__11), .q_0__10 (
            que_out_26__0__10), .q_0__9 (que_out_26__0__9), .q_0__8 (
            que_out_26__0__8), .q_0__7 (que_out_26__0__7), .q_0__6 (
            que_out_26__0__6), .q_0__5 (que_out_26__0__5), .q_0__4 (
            que_out_26__0__4), .q_0__3 (que_out_26__0__3), .q_0__2 (
            que_out_26__0__2), .q_0__1 (que_out_26__0__1), .q_0__0 (
            que_out_26__0__0), .q_1__15 (que_out_26__1__15), .q_1__14 (
            que_out_26__1__14), .q_1__13 (que_out_26__1__13), .q_1__12 (
            que_out_26__1__12), .q_1__11 (que_out_26__1__11), .q_1__10 (
            que_out_26__1__10), .q_1__9 (que_out_26__1__9), .q_1__8 (
            que_out_26__1__8), .q_1__7 (que_out_26__1__7), .q_1__6 (
            que_out_26__1__6), .q_1__5 (que_out_26__1__5), .q_1__4 (
            que_out_26__1__4), .q_1__3 (que_out_26__1__3), .q_1__2 (
            que_out_26__1__2), .q_1__1 (que_out_26__1__1), .q_1__0 (
            que_out_26__1__0), .q_2__15 (que_out_26__2__15), .q_2__14 (
            que_out_26__2__14), .q_2__13 (que_out_26__2__13), .q_2__12 (
            que_out_26__2__12), .q_2__11 (que_out_26__2__11), .q_2__10 (
            que_out_26__2__10), .q_2__9 (que_out_26__2__9), .q_2__8 (
            que_out_26__2__8), .q_2__7 (que_out_26__2__7), .q_2__6 (
            que_out_26__2__6), .q_2__5 (que_out_26__2__5), .q_2__4 (
            que_out_26__2__4), .q_2__3 (que_out_26__2__3), .q_2__2 (
            que_out_26__2__2), .q_2__1 (que_out_26__2__1), .q_2__0 (
            que_out_26__2__0), .q_3__15 (que_out_26__3__15), .q_3__14 (
            que_out_26__3__14), .q_3__13 (que_out_26__3__13), .q_3__12 (
            que_out_26__3__12), .q_3__11 (que_out_26__3__11), .q_3__10 (
            que_out_26__3__10), .q_3__9 (que_out_26__3__9), .q_3__8 (
            que_out_26__3__8), .q_3__7 (que_out_26__3__7), .q_3__6 (
            que_out_26__3__6), .q_3__5 (que_out_26__3__5), .q_3__4 (
            que_out_26__3__4), .q_3__3 (que_out_26__3__3), .q_3__2 (
            que_out_26__3__2), .q_3__1 (que_out_26__3__1), .q_3__0 (
            que_out_26__3__0), .q_4__15 (que_out_26__4__15), .q_4__14 (
            que_out_26__4__14), .q_4__13 (que_out_26__4__13), .q_4__12 (
            que_out_26__4__12), .q_4__11 (que_out_26__4__11), .q_4__10 (
            que_out_26__4__10), .q_4__9 (que_out_26__4__9), .q_4__8 (
            que_out_26__4__8), .q_4__7 (que_out_26__4__7), .q_4__6 (
            que_out_26__4__6), .q_4__5 (que_out_26__4__5), .q_4__4 (
            que_out_26__4__4), .q_4__3 (que_out_26__4__3), .q_4__2 (
            que_out_26__4__2), .q_4__1 (que_out_26__4__1), .q_4__0 (
            que_out_26__4__0), .clk (nx10734), .load (sel_que_26), .reset (
            nx10710)) ;
    Queue_5 gen_queues_27_que (.d ({nx10518,nx10528,nx10538,nx10548,nx10558,
            nx10568,nx10578,nx10588,nx10598,nx10608,nx10618,nx10628,nx10638,
            nx10648,nx10658,nx10668}), .q_0__15 (que_out_27__0__15), .q_0__14 (
            que_out_27__0__14), .q_0__13 (que_out_27__0__13), .q_0__12 (
            que_out_27__0__12), .q_0__11 (que_out_27__0__11), .q_0__10 (
            que_out_27__0__10), .q_0__9 (que_out_27__0__9), .q_0__8 (
            que_out_27__0__8), .q_0__7 (que_out_27__0__7), .q_0__6 (
            que_out_27__0__6), .q_0__5 (que_out_27__0__5), .q_0__4 (
            que_out_27__0__4), .q_0__3 (que_out_27__0__3), .q_0__2 (
            que_out_27__0__2), .q_0__1 (que_out_27__0__1), .q_0__0 (
            que_out_27__0__0), .q_1__15 (que_out_27__1__15), .q_1__14 (
            que_out_27__1__14), .q_1__13 (que_out_27__1__13), .q_1__12 (
            que_out_27__1__12), .q_1__11 (que_out_27__1__11), .q_1__10 (
            que_out_27__1__10), .q_1__9 (que_out_27__1__9), .q_1__8 (
            que_out_27__1__8), .q_1__7 (que_out_27__1__7), .q_1__6 (
            que_out_27__1__6), .q_1__5 (que_out_27__1__5), .q_1__4 (
            que_out_27__1__4), .q_1__3 (que_out_27__1__3), .q_1__2 (
            que_out_27__1__2), .q_1__1 (que_out_27__1__1), .q_1__0 (
            que_out_27__1__0), .q_2__15 (que_out_27__2__15), .q_2__14 (
            que_out_27__2__14), .q_2__13 (que_out_27__2__13), .q_2__12 (
            que_out_27__2__12), .q_2__11 (que_out_27__2__11), .q_2__10 (
            que_out_27__2__10), .q_2__9 (que_out_27__2__9), .q_2__8 (
            que_out_27__2__8), .q_2__7 (que_out_27__2__7), .q_2__6 (
            que_out_27__2__6), .q_2__5 (que_out_27__2__5), .q_2__4 (
            que_out_27__2__4), .q_2__3 (que_out_27__2__3), .q_2__2 (
            que_out_27__2__2), .q_2__1 (que_out_27__2__1), .q_2__0 (
            que_out_27__2__0), .q_3__15 (que_out_27__3__15), .q_3__14 (
            que_out_27__3__14), .q_3__13 (que_out_27__3__13), .q_3__12 (
            que_out_27__3__12), .q_3__11 (que_out_27__3__11), .q_3__10 (
            que_out_27__3__10), .q_3__9 (que_out_27__3__9), .q_3__8 (
            que_out_27__3__8), .q_3__7 (que_out_27__3__7), .q_3__6 (
            que_out_27__3__6), .q_3__5 (que_out_27__3__5), .q_3__4 (
            que_out_27__3__4), .q_3__3 (que_out_27__3__3), .q_3__2 (
            que_out_27__3__2), .q_3__1 (que_out_27__3__1), .q_3__0 (
            que_out_27__3__0), .q_4__15 (que_out_27__4__15), .q_4__14 (
            que_out_27__4__14), .q_4__13 (que_out_27__4__13), .q_4__12 (
            que_out_27__4__12), .q_4__11 (que_out_27__4__11), .q_4__10 (
            que_out_27__4__10), .q_4__9 (que_out_27__4__9), .q_4__8 (
            que_out_27__4__8), .q_4__7 (que_out_27__4__7), .q_4__6 (
            que_out_27__4__6), .q_4__5 (que_out_27__4__5), .q_4__4 (
            que_out_27__4__4), .q_4__3 (que_out_27__4__3), .q_4__2 (
            que_out_27__4__2), .q_4__1 (que_out_27__4__1), .q_4__0 (
            que_out_27__4__0), .clk (nx10736), .load (sel_que_27), .reset (
            nx10712)) ;
    nand03 ix6830 (.Y (nx6829), .A0 (nx8938), .A1 (nx6833), .A2 (nx6835)) ;
    nor02ii ix8939 (.Y (nx8938), .A0 (cache_in_sel[4]), .A1 (decoder_enable)) ;
    inv01 ix6834 (.Y (nx6833), .A (cache_in_sel[1])) ;
    inv01 ix6836 (.Y (nx6835), .A (cache_in_sel[0])) ;
    nand03 ix6840 (.Y (nx6839), .A0 (nx8938), .A1 (nx6833), .A2 (nx10508)) ;
    nand03 ix6844 (.Y (nx6843), .A0 (nx8938), .A1 (nx10506), .A2 (nx6835)) ;
    nand03 ix6848 (.Y (nx6847), .A0 (nx8938), .A1 (nx10506), .A2 (nx10508)) ;
    nor02_2x ix9023 (.Y (sel_que_12), .A0 (nx6875), .A1 (nx6829)) ;
    nand02 ix6876 (.Y (nx6875), .A0 (cache_in_sel[3]), .A1 (cache_in_sel[2])) ;
    nor02_2x ix9025 (.Y (sel_que_13), .A0 (nx6875), .A1 (nx6839)) ;
    nor02_2x ix9027 (.Y (sel_que_14), .A0 (nx6843), .A1 (nx6875)) ;
    nor02_2x ix9029 (.Y (sel_que_15), .A0 (nx6875), .A1 (nx6847)) ;
    and02 ix9043 (.Y (sel_que_16), .A0 (nx6885), .A1 (nx9038)) ;
    nor02_2x ix6886 (.Y (nx6885), .A0 (cache_in_sel[2]), .A1 (cache_in_sel[3])
             ) ;
    nor03_2x ix9039 (.Y (nx9038), .A0 (nx6889), .A1 (nx10506), .A2 (nx10508)) ;
    nand02 ix6890 (.Y (nx6889), .A0 (cache_in_sel[4]), .A1 (decoder_enable)) ;
    nand04 ix6894 (.Y (nx6893), .A0 (cache_in_sel[4]), .A1 (decoder_enable), .A2 (
           nx6833), .A3 (nx10508)) ;
    nand04 ix6898 (.Y (nx6897), .A0 (cache_in_sel[4]), .A1 (decoder_enable), .A2 (
           nx10506), .A3 (nx6835)) ;
    nand04 ix6902 (.Y (nx6901), .A0 (cache_in_sel[4]), .A1 (decoder_enable), .A2 (
           nx10506), .A3 (nx10508)) ;
    and02 ix9075 (.Y (sel_que_20), .A0 (nx6905), .A1 (nx9038)) ;
    and02 ix9091 (.Y (sel_que_24), .A0 (nx6915), .A1 (nx9038)) ;
    or04 ix243 (.Y (out_column_4__0), .A0 (nx238), .A1 (nx188), .A2 (nx130), .A3 (
         nx82)) ;
    nand03 ix239 (.Y (nx238), .A0 (nx6927), .A1 (nx6951), .A2 (nx6967)) ;
    aoi222 ix6928 (.Y (nx6927), .A0 (que_out_10__4__0), .A1 (nx10298), .B0 (
           que_out_6__4__0), .B1 (nx10350), .C0 (que_out_9__4__0), .C1 (nx10324)
           ) ;
    nand02_2x ix6932 (.Y (nx6931), .A0 (cache_out_sel[3]), .A1 (nx6933)) ;
    inv01 ix6934 (.Y (nx6933), .A (cache_out_sel[0])) ;
    inv01 ix6938 (.Y (nx6937), .A (cache_out_sel[4])) ;
    inv02 ix6940 (.Y (nx6939), .A (cache_out_sel[2])) ;
    nand03 ix6946 (.Y (nx6945), .A0 (nx10502), .A1 (nx6937), .A2 (nx10498)) ;
    nor04 ix227 (.Y (nx226), .A0 (nx6949), .A1 (nx10502), .A2 (nx10494), .A3 (
          nx10498)) ;
    nand02_2x ix6950 (.Y (nx6949), .A0 (cache_out_sel[3]), .A1 (cache_out_sel[0]
              )) ;
    aoi22 ix6952 (.Y (nx6951), .A0 (que_out_5__4__0), .A1 (nx10246), .B0 (
          que_out_18__4__0), .B1 (nx10272)) ;
    nand02 ix6956 (.Y (nx6955), .A0 (nx6957), .A1 (cache_out_sel[0])) ;
    inv01 ix6958 (.Y (nx6957), .A (cache_out_sel[3])) ;
    inv01 ix6962 (.Y (nx6961), .A (cache_out_sel[1])) ;
    nor03_2x ix215 (.Y (nx214), .A0 (nx6965), .A1 (nx10498), .A2 (nx6943)) ;
    nand02_2x ix6966 (.Y (nx6965), .A0 (nx10494), .A1 (nx10504)) ;
    aoi22 ix6968 (.Y (nx6967), .A0 (que_out_17__4__0), .A1 (nx10220), .B0 (
          que_out_20__4__0), .B1 (nx10194)) ;
    nor03_2x ix201 (.Y (nx200), .A0 (nx6971), .A1 (nx10498), .A2 (nx10374)) ;
    nand02_2x ix6972 (.Y (nx6971), .A0 (nx10496), .A1 (nx6961)) ;
    nor03_2x ix193 (.Y (nx192), .A0 (nx6971), .A1 (nx6939), .A2 (nx6943)) ;
    nand03 ix189 (.Y (nx188), .A0 (nx6977), .A1 (nx6985), .A2 (nx6991)) ;
    aoi222 ix6978 (.Y (nx6977), .A0 (que_out_19__4__0), .A1 (nx10168), .B0 (
           que_out_21__4__0), .B1 (nx10142), .C0 (que_out_8__4__0), .C1 (nx10116
           )) ;
    nor03_2x ix181 (.Y (nx180), .A0 (nx6965), .A1 (nx10498), .A2 (nx10374)) ;
    nor03_2x ix173 (.Y (nx172), .A0 (nx6971), .A1 (nx6939), .A2 (nx10374)) ;
    nor04 ix167 (.Y (nx166), .A0 (nx6931), .A1 (nx10502), .A2 (nx10494), .A3 (
          nx10498)) ;
    aoi22 ix6986 (.Y (nx6985), .A0 (que_out_25__4__0), .A1 (nx10064), .B0 (
          que_out_16__4__0), .B1 (nx10090)) ;
    nor02_2x ix151 (.Y (nx150), .A0 (nx6949), .A1 (nx6971)) ;
    nor03_2x ix159 (.Y (nx158), .A0 (nx6971), .A1 (nx10498), .A2 (nx6943)) ;
    aoi22 ix6992 (.Y (nx6991), .A0 (que_out_24__4__0), .A1 (nx10038), .B0 (
          que_out_22__4__0), .B1 (nx10012)) ;
    nor02_2x ix145 (.Y (nx144), .A0 (nx6971), .A1 (nx6931)) ;
    nor03_2x ix137 (.Y (nx136), .A0 (nx6965), .A1 (nx6939), .A2 (nx6943)) ;
    nand03 ix131 (.Y (nx130), .A0 (nx6999), .A1 (nx7007), .A2 (nx7017)) ;
    aoi222 ix7000 (.Y (nx6999), .A0 (que_out_15__4__0), .A1 (nx9960), .B0 (
           que_out_3__4__0), .B1 (nx9986), .C0 (que_out_23__4__0), .C1 (nx9934)
           ) ;
    nor02_2x ix119 (.Y (nx118), .A0 (nx6949), .A1 (nx6945)) ;
    nor03_2x ix115 (.Y (nx114), .A0 (nx6965), .A1 (nx6939), .A2 (nx10374)) ;
    aoi22 ix7008 (.Y (nx7007), .A0 (que_out_27__4__0), .A1 (nx9908), .B0 (
          que_out_4__4__0), .B1 (nx9882)) ;
    nor02_2x ix105 (.Y (nx104), .A0 (nx6949), .A1 (nx6965)) ;
    and02 ix101 (.Y (nx100), .A0 (nx88), .A1 (nx28)) ;
    nor02_2x ix89 (.Y (nx88), .A0 (cache_out_sel[3]), .A1 (cache_out_sel[0])) ;
    nor03_2x ix29 (.Y (nx28), .A0 (nx10502), .A1 (nx10494), .A2 (nx6939)) ;
    aoi22 ix7018 (.Y (nx7017), .A0 (que_out_0__4__0), .A1 (nx9830), .B0 (
          que_out_2__4__0), .B1 (nx9856)) ;
    and02 ix91 (.Y (nx90), .A0 (nx88), .A1 (nx12)) ;
    nor03_2x ix13 (.Y (nx12), .A0 (nx10504), .A1 (nx10494), .A2 (nx10500)) ;
    and02 ix95 (.Y (nx94), .A0 (nx88), .A1 (nx62)) ;
    nor03_2x ix63 (.Y (nx62), .A0 (nx6961), .A1 (nx10494), .A2 (nx10500)) ;
    nand03 ix83 (.Y (nx82), .A0 (nx7029), .A1 (nx7037), .A2 (nx7043)) ;
    aoi222 ix7030 (.Y (nx7029), .A0 (que_out_26__4__0), .A1 (nx9804), .B0 (
           que_out_14__4__0), .B1 (nx9778), .C0 (que_out_11__4__0), .C1 (nx9752)
           ) ;
    nor02_2x ix75 (.Y (nx74), .A0 (nx6965), .A1 (nx6931)) ;
    nor02_2x ix69 (.Y (nx68), .A0 (nx6931), .A1 (nx6945)) ;
    aoi22 ix7038 (.Y (nx7037), .A0 (que_out_13__4__0), .A1 (nx9726), .B0 (
          que_out_7__4__0), .B1 (nx9700)) ;
    nor02_2x ix43 (.Y (nx42), .A0 (nx10374), .A1 (nx6945)) ;
    aoi22 ix7044 (.Y (nx7043), .A0 (que_out_12__4__0), .A1 (nx9674), .B0 (
          que_out_1__4__0), .B1 (nx9648)) ;
    nor04 ix15 (.Y (nx14), .A0 (nx10376), .A1 (nx10504), .A2 (nx10494), .A3 (
          nx10500)) ;
    or04 ix353 (.Y (out_column_4__1), .A0 (nx348), .A1 (nx322), .A2 (nx294), .A3 (
         nx268)) ;
    nand03 ix349 (.Y (nx348), .A0 (nx7053), .A1 (nx7055), .A2 (nx7057)) ;
    aoi222 ix7054 (.Y (nx7053), .A0 (que_out_10__4__1), .A1 (nx10298), .B0 (
           que_out_6__4__1), .B1 (nx10350), .C0 (que_out_9__4__1), .C1 (nx10324)
           ) ;
    aoi22 ix7056 (.Y (nx7055), .A0 (que_out_5__4__1), .A1 (nx10246), .B0 (
          que_out_18__4__1), .B1 (nx10272)) ;
    aoi22 ix7058 (.Y (nx7057), .A0 (que_out_17__4__1), .A1 (nx10220), .B0 (
          que_out_20__4__1), .B1 (nx10194)) ;
    nand03 ix323 (.Y (nx322), .A0 (nx7061), .A1 (nx7063), .A2 (nx7065)) ;
    aoi222 ix7062 (.Y (nx7061), .A0 (que_out_19__4__1), .A1 (nx10168), .B0 (
           que_out_21__4__1), .B1 (nx10142), .C0 (que_out_8__4__1), .C1 (nx10116
           )) ;
    aoi22 ix7064 (.Y (nx7063), .A0 (que_out_25__4__1), .A1 (nx10064), .B0 (
          que_out_16__4__1), .B1 (nx10090)) ;
    aoi22 ix7066 (.Y (nx7065), .A0 (que_out_24__4__1), .A1 (nx10038), .B0 (
          que_out_22__4__1), .B1 (nx10012)) ;
    nand03 ix295 (.Y (nx294), .A0 (nx7069), .A1 (nx7071), .A2 (nx7073)) ;
    aoi222 ix7070 (.Y (nx7069), .A0 (que_out_15__4__1), .A1 (nx9960), .B0 (
           que_out_3__4__1), .B1 (nx9986), .C0 (que_out_23__4__1), .C1 (nx9934)
           ) ;
    aoi22 ix7072 (.Y (nx7071), .A0 (que_out_27__4__1), .A1 (nx9908), .B0 (
          que_out_4__4__1), .B1 (nx9882)) ;
    aoi22 ix7074 (.Y (nx7073), .A0 (que_out_0__4__1), .A1 (nx9830), .B0 (
          que_out_2__4__1), .B1 (nx9856)) ;
    nand03 ix269 (.Y (nx268), .A0 (nx7077), .A1 (nx7079), .A2 (nx7081)) ;
    aoi222 ix7078 (.Y (nx7077), .A0 (que_out_26__4__1), .A1 (nx9804), .B0 (
           que_out_14__4__1), .B1 (nx9778), .C0 (que_out_11__4__1), .C1 (nx9752)
           ) ;
    aoi22 ix7080 (.Y (nx7079), .A0 (que_out_13__4__1), .A1 (nx9726), .B0 (
          que_out_7__4__1), .B1 (nx9700)) ;
    aoi22 ix7082 (.Y (nx7081), .A0 (que_out_12__4__1), .A1 (nx9674), .B0 (
          que_out_1__4__1), .B1 (nx9648)) ;
    or04 ix463 (.Y (out_column_4__2), .A0 (nx458), .A1 (nx432), .A2 (nx404), .A3 (
         nx378)) ;
    nand03 ix459 (.Y (nx458), .A0 (nx7087), .A1 (nx7089), .A2 (nx7091)) ;
    aoi222 ix7088 (.Y (nx7087), .A0 (que_out_10__4__2), .A1 (nx10298), .B0 (
           que_out_6__4__2), .B1 (nx10350), .C0 (que_out_9__4__2), .C1 (nx10324)
           ) ;
    aoi22 ix7090 (.Y (nx7089), .A0 (que_out_5__4__2), .A1 (nx10246), .B0 (
          que_out_18__4__2), .B1 (nx10272)) ;
    aoi22 ix7092 (.Y (nx7091), .A0 (que_out_17__4__2), .A1 (nx10220), .B0 (
          que_out_20__4__2), .B1 (nx10194)) ;
    nand03 ix433 (.Y (nx432), .A0 (nx7095), .A1 (nx7097), .A2 (nx7099)) ;
    aoi222 ix7096 (.Y (nx7095), .A0 (que_out_19__4__2), .A1 (nx10168), .B0 (
           que_out_21__4__2), .B1 (nx10142), .C0 (que_out_8__4__2), .C1 (nx10116
           )) ;
    aoi22 ix7098 (.Y (nx7097), .A0 (que_out_25__4__2), .A1 (nx10064), .B0 (
          que_out_16__4__2), .B1 (nx10090)) ;
    aoi22 ix7100 (.Y (nx7099), .A0 (que_out_24__4__2), .A1 (nx10038), .B0 (
          que_out_22__4__2), .B1 (nx10012)) ;
    nand03 ix405 (.Y (nx404), .A0 (nx7103), .A1 (nx7105), .A2 (nx7107)) ;
    aoi222 ix7104 (.Y (nx7103), .A0 (que_out_15__4__2), .A1 (nx9960), .B0 (
           que_out_3__4__2), .B1 (nx9986), .C0 (que_out_23__4__2), .C1 (nx9934)
           ) ;
    aoi22 ix7106 (.Y (nx7105), .A0 (que_out_27__4__2), .A1 (nx9908), .B0 (
          que_out_4__4__2), .B1 (nx9882)) ;
    aoi22 ix7108 (.Y (nx7107), .A0 (que_out_0__4__2), .A1 (nx9830), .B0 (
          que_out_2__4__2), .B1 (nx9856)) ;
    nand03 ix379 (.Y (nx378), .A0 (nx7111), .A1 (nx7113), .A2 (nx7115)) ;
    aoi222 ix7112 (.Y (nx7111), .A0 (que_out_26__4__2), .A1 (nx9804), .B0 (
           que_out_14__4__2), .B1 (nx9778), .C0 (que_out_11__4__2), .C1 (nx9752)
           ) ;
    aoi22 ix7114 (.Y (nx7113), .A0 (que_out_13__4__2), .A1 (nx9726), .B0 (
          que_out_7__4__2), .B1 (nx9700)) ;
    aoi22 ix7116 (.Y (nx7115), .A0 (que_out_12__4__2), .A1 (nx9674), .B0 (
          que_out_1__4__2), .B1 (nx9648)) ;
    or04 ix573 (.Y (out_column_4__3), .A0 (nx568), .A1 (nx542), .A2 (nx514), .A3 (
         nx488)) ;
    nand03 ix569 (.Y (nx568), .A0 (nx7121), .A1 (nx7123), .A2 (nx7125)) ;
    aoi222 ix7122 (.Y (nx7121), .A0 (que_out_10__4__3), .A1 (nx10298), .B0 (
           que_out_6__4__3), .B1 (nx10350), .C0 (que_out_9__4__3), .C1 (nx10324)
           ) ;
    aoi22 ix7124 (.Y (nx7123), .A0 (que_out_5__4__3), .A1 (nx10246), .B0 (
          que_out_18__4__3), .B1 (nx10272)) ;
    aoi22 ix7126 (.Y (nx7125), .A0 (que_out_17__4__3), .A1 (nx10220), .B0 (
          que_out_20__4__3), .B1 (nx10194)) ;
    nand03 ix543 (.Y (nx542), .A0 (nx7129), .A1 (nx7131), .A2 (nx7133)) ;
    aoi222 ix7130 (.Y (nx7129), .A0 (que_out_19__4__3), .A1 (nx10168), .B0 (
           que_out_21__4__3), .B1 (nx10142), .C0 (que_out_8__4__3), .C1 (nx10116
           )) ;
    aoi22 ix7132 (.Y (nx7131), .A0 (que_out_25__4__3), .A1 (nx10064), .B0 (
          que_out_16__4__3), .B1 (nx10090)) ;
    aoi22 ix7134 (.Y (nx7133), .A0 (que_out_24__4__3), .A1 (nx10038), .B0 (
          que_out_22__4__3), .B1 (nx10012)) ;
    nand03 ix515 (.Y (nx514), .A0 (nx7137), .A1 (nx7139), .A2 (nx7141)) ;
    aoi222 ix7138 (.Y (nx7137), .A0 (que_out_15__4__3), .A1 (nx9960), .B0 (
           que_out_3__4__3), .B1 (nx9986), .C0 (que_out_23__4__3), .C1 (nx9934)
           ) ;
    aoi22 ix7140 (.Y (nx7139), .A0 (que_out_27__4__3), .A1 (nx9908), .B0 (
          que_out_4__4__3), .B1 (nx9882)) ;
    aoi22 ix7142 (.Y (nx7141), .A0 (que_out_0__4__3), .A1 (nx9830), .B0 (
          que_out_2__4__3), .B1 (nx9856)) ;
    nand03 ix489 (.Y (nx488), .A0 (nx7145), .A1 (nx7147), .A2 (nx7149)) ;
    aoi222 ix7146 (.Y (nx7145), .A0 (que_out_26__4__3), .A1 (nx9804), .B0 (
           que_out_14__4__3), .B1 (nx9778), .C0 (que_out_11__4__3), .C1 (nx9752)
           ) ;
    aoi22 ix7148 (.Y (nx7147), .A0 (que_out_13__4__3), .A1 (nx9726), .B0 (
          que_out_7__4__3), .B1 (nx9700)) ;
    aoi22 ix7150 (.Y (nx7149), .A0 (que_out_12__4__3), .A1 (nx9674), .B0 (
          que_out_1__4__3), .B1 (nx9648)) ;
    or04 ix683 (.Y (out_column_4__4), .A0 (nx678), .A1 (nx652), .A2 (nx624), .A3 (
         nx598)) ;
    nand03 ix679 (.Y (nx678), .A0 (nx7155), .A1 (nx7157), .A2 (nx7159)) ;
    aoi222 ix7156 (.Y (nx7155), .A0 (que_out_10__4__4), .A1 (nx10298), .B0 (
           que_out_6__4__4), .B1 (nx10350), .C0 (que_out_9__4__4), .C1 (nx10324)
           ) ;
    aoi22 ix7158 (.Y (nx7157), .A0 (que_out_5__4__4), .A1 (nx10246), .B0 (
          que_out_18__4__4), .B1 (nx10272)) ;
    aoi22 ix7160 (.Y (nx7159), .A0 (que_out_17__4__4), .A1 (nx10220), .B0 (
          que_out_20__4__4), .B1 (nx10194)) ;
    nand03 ix653 (.Y (nx652), .A0 (nx7163), .A1 (nx7165), .A2 (nx7167)) ;
    aoi222 ix7164 (.Y (nx7163), .A0 (que_out_19__4__4), .A1 (nx10168), .B0 (
           que_out_21__4__4), .B1 (nx10142), .C0 (que_out_8__4__4), .C1 (nx10116
           )) ;
    aoi22 ix7166 (.Y (nx7165), .A0 (que_out_25__4__4), .A1 (nx10064), .B0 (
          que_out_16__4__4), .B1 (nx10090)) ;
    aoi22 ix7168 (.Y (nx7167), .A0 (que_out_24__4__4), .A1 (nx10038), .B0 (
          que_out_22__4__4), .B1 (nx10012)) ;
    nand03 ix625 (.Y (nx624), .A0 (nx7171), .A1 (nx7173), .A2 (nx7175)) ;
    aoi222 ix7172 (.Y (nx7171), .A0 (que_out_15__4__4), .A1 (nx9960), .B0 (
           que_out_3__4__4), .B1 (nx9986), .C0 (que_out_23__4__4), .C1 (nx9934)
           ) ;
    aoi22 ix7174 (.Y (nx7173), .A0 (que_out_27__4__4), .A1 (nx9908), .B0 (
          que_out_4__4__4), .B1 (nx9882)) ;
    aoi22 ix7176 (.Y (nx7175), .A0 (que_out_0__4__4), .A1 (nx9830), .B0 (
          que_out_2__4__4), .B1 (nx9856)) ;
    nand03 ix599 (.Y (nx598), .A0 (nx7179), .A1 (nx7181), .A2 (nx7183)) ;
    aoi222 ix7180 (.Y (nx7179), .A0 (que_out_26__4__4), .A1 (nx9804), .B0 (
           que_out_14__4__4), .B1 (nx9778), .C0 (que_out_11__4__4), .C1 (nx9752)
           ) ;
    aoi22 ix7182 (.Y (nx7181), .A0 (que_out_13__4__4), .A1 (nx9726), .B0 (
          que_out_7__4__4), .B1 (nx9700)) ;
    aoi22 ix7184 (.Y (nx7183), .A0 (que_out_12__4__4), .A1 (nx9674), .B0 (
          que_out_1__4__4), .B1 (nx9648)) ;
    or04 ix793 (.Y (out_column_4__5), .A0 (nx788), .A1 (nx762), .A2 (nx734), .A3 (
         nx708)) ;
    nand03 ix789 (.Y (nx788), .A0 (nx7189), .A1 (nx7191), .A2 (nx7193)) ;
    aoi222 ix7190 (.Y (nx7189), .A0 (que_out_10__4__5), .A1 (nx10298), .B0 (
           que_out_6__4__5), .B1 (nx10350), .C0 (que_out_9__4__5), .C1 (nx10324)
           ) ;
    aoi22 ix7192 (.Y (nx7191), .A0 (que_out_5__4__5), .A1 (nx10246), .B0 (
          que_out_18__4__5), .B1 (nx10272)) ;
    aoi22 ix7194 (.Y (nx7193), .A0 (que_out_17__4__5), .A1 (nx10220), .B0 (
          que_out_20__4__5), .B1 (nx10194)) ;
    nand03 ix763 (.Y (nx762), .A0 (nx7197), .A1 (nx7199), .A2 (nx7201)) ;
    aoi222 ix7198 (.Y (nx7197), .A0 (que_out_19__4__5), .A1 (nx10168), .B0 (
           que_out_21__4__5), .B1 (nx10142), .C0 (que_out_8__4__5), .C1 (nx10116
           )) ;
    aoi22 ix7200 (.Y (nx7199), .A0 (que_out_25__4__5), .A1 (nx10064), .B0 (
          que_out_16__4__5), .B1 (nx10090)) ;
    aoi22 ix7202 (.Y (nx7201), .A0 (que_out_24__4__5), .A1 (nx10038), .B0 (
          que_out_22__4__5), .B1 (nx10012)) ;
    nand03 ix735 (.Y (nx734), .A0 (nx7205), .A1 (nx7207), .A2 (nx7209)) ;
    aoi222 ix7206 (.Y (nx7205), .A0 (que_out_15__4__5), .A1 (nx9960), .B0 (
           que_out_3__4__5), .B1 (nx9986), .C0 (que_out_23__4__5), .C1 (nx9934)
           ) ;
    aoi22 ix7208 (.Y (nx7207), .A0 (que_out_27__4__5), .A1 (nx9908), .B0 (
          que_out_4__4__5), .B1 (nx9882)) ;
    aoi22 ix7210 (.Y (nx7209), .A0 (que_out_0__4__5), .A1 (nx9830), .B0 (
          que_out_2__4__5), .B1 (nx9856)) ;
    nand03 ix709 (.Y (nx708), .A0 (nx7213), .A1 (nx7215), .A2 (nx7217)) ;
    aoi222 ix7214 (.Y (nx7213), .A0 (que_out_26__4__5), .A1 (nx9804), .B0 (
           que_out_14__4__5), .B1 (nx9778), .C0 (que_out_11__4__5), .C1 (nx9752)
           ) ;
    aoi22 ix7216 (.Y (nx7215), .A0 (que_out_13__4__5), .A1 (nx9726), .B0 (
          que_out_7__4__5), .B1 (nx9700)) ;
    aoi22 ix7218 (.Y (nx7217), .A0 (que_out_12__4__5), .A1 (nx9674), .B0 (
          que_out_1__4__5), .B1 (nx9648)) ;
    or04 ix903 (.Y (out_column_4__6), .A0 (nx898), .A1 (nx872), .A2 (nx844), .A3 (
         nx818)) ;
    nand03 ix899 (.Y (nx898), .A0 (nx7223), .A1 (nx7225), .A2 (nx7227)) ;
    aoi222 ix7224 (.Y (nx7223), .A0 (que_out_10__4__6), .A1 (nx10298), .B0 (
           que_out_6__4__6), .B1 (nx10350), .C0 (que_out_9__4__6), .C1 (nx10324)
           ) ;
    aoi22 ix7226 (.Y (nx7225), .A0 (que_out_5__4__6), .A1 (nx10246), .B0 (
          que_out_18__4__6), .B1 (nx10272)) ;
    aoi22 ix7228 (.Y (nx7227), .A0 (que_out_17__4__6), .A1 (nx10220), .B0 (
          que_out_20__4__6), .B1 (nx10194)) ;
    nand03 ix873 (.Y (nx872), .A0 (nx7231), .A1 (nx7233), .A2 (nx7235)) ;
    aoi222 ix7232 (.Y (nx7231), .A0 (que_out_19__4__6), .A1 (nx10168), .B0 (
           que_out_21__4__6), .B1 (nx10142), .C0 (que_out_8__4__6), .C1 (nx10116
           )) ;
    aoi22 ix7234 (.Y (nx7233), .A0 (que_out_25__4__6), .A1 (nx10064), .B0 (
          que_out_16__4__6), .B1 (nx10090)) ;
    aoi22 ix7236 (.Y (nx7235), .A0 (que_out_24__4__6), .A1 (nx10038), .B0 (
          que_out_22__4__6), .B1 (nx10012)) ;
    nand03 ix845 (.Y (nx844), .A0 (nx7239), .A1 (nx7241), .A2 (nx7243)) ;
    aoi222 ix7240 (.Y (nx7239), .A0 (que_out_15__4__6), .A1 (nx9960), .B0 (
           que_out_3__4__6), .B1 (nx9986), .C0 (que_out_23__4__6), .C1 (nx9934)
           ) ;
    aoi22 ix7242 (.Y (nx7241), .A0 (que_out_27__4__6), .A1 (nx9908), .B0 (
          que_out_4__4__6), .B1 (nx9882)) ;
    aoi22 ix7244 (.Y (nx7243), .A0 (que_out_0__4__6), .A1 (nx9830), .B0 (
          que_out_2__4__6), .B1 (nx9856)) ;
    nand03 ix819 (.Y (nx818), .A0 (nx7247), .A1 (nx7249), .A2 (nx7251)) ;
    aoi222 ix7248 (.Y (nx7247), .A0 (que_out_26__4__6), .A1 (nx9804), .B0 (
           que_out_14__4__6), .B1 (nx9778), .C0 (que_out_11__4__6), .C1 (nx9752)
           ) ;
    aoi22 ix7250 (.Y (nx7249), .A0 (que_out_13__4__6), .A1 (nx9726), .B0 (
          que_out_7__4__6), .B1 (nx9700)) ;
    aoi22 ix7252 (.Y (nx7251), .A0 (que_out_12__4__6), .A1 (nx9674), .B0 (
          que_out_1__4__6), .B1 (nx9648)) ;
    or04 ix1013 (.Y (out_column_4__7), .A0 (nx1008), .A1 (nx982), .A2 (nx954), .A3 (
         nx928)) ;
    nand03 ix1009 (.Y (nx1008), .A0 (nx7257), .A1 (nx7259), .A2 (nx7261)) ;
    aoi222 ix7258 (.Y (nx7257), .A0 (que_out_10__4__7), .A1 (nx10300), .B0 (
           que_out_6__4__7), .B1 (nx10352), .C0 (que_out_9__4__7), .C1 (nx10326)
           ) ;
    aoi22 ix7260 (.Y (nx7259), .A0 (que_out_5__4__7), .A1 (nx10248), .B0 (
          que_out_18__4__7), .B1 (nx10274)) ;
    aoi22 ix7262 (.Y (nx7261), .A0 (que_out_17__4__7), .A1 (nx10222), .B0 (
          que_out_20__4__7), .B1 (nx10196)) ;
    nand03 ix983 (.Y (nx982), .A0 (nx7265), .A1 (nx7267), .A2 (nx7269)) ;
    aoi222 ix7266 (.Y (nx7265), .A0 (que_out_19__4__7), .A1 (nx10170), .B0 (
           que_out_21__4__7), .B1 (nx10144), .C0 (que_out_8__4__7), .C1 (nx10118
           )) ;
    aoi22 ix7268 (.Y (nx7267), .A0 (que_out_25__4__7), .A1 (nx10066), .B0 (
          que_out_16__4__7), .B1 (nx10092)) ;
    aoi22 ix7270 (.Y (nx7269), .A0 (que_out_24__4__7), .A1 (nx10040), .B0 (
          que_out_22__4__7), .B1 (nx10014)) ;
    nand03 ix955 (.Y (nx954), .A0 (nx7273), .A1 (nx7275), .A2 (nx7277)) ;
    aoi222 ix7274 (.Y (nx7273), .A0 (que_out_15__4__7), .A1 (nx9962), .B0 (
           que_out_3__4__7), .B1 (nx9988), .C0 (que_out_23__4__7), .C1 (nx9936)
           ) ;
    aoi22 ix7276 (.Y (nx7275), .A0 (que_out_27__4__7), .A1 (nx9910), .B0 (
          que_out_4__4__7), .B1 (nx9884)) ;
    aoi22 ix7278 (.Y (nx7277), .A0 (que_out_0__4__7), .A1 (nx9832), .B0 (
          que_out_2__4__7), .B1 (nx9858)) ;
    nand03 ix929 (.Y (nx928), .A0 (nx7281), .A1 (nx7283), .A2 (nx7285)) ;
    aoi222 ix7282 (.Y (nx7281), .A0 (que_out_26__4__7), .A1 (nx9806), .B0 (
           que_out_14__4__7), .B1 (nx9780), .C0 (que_out_11__4__7), .C1 (nx9754)
           ) ;
    aoi22 ix7284 (.Y (nx7283), .A0 (que_out_13__4__7), .A1 (nx9728), .B0 (
          que_out_7__4__7), .B1 (nx9702)) ;
    aoi22 ix7286 (.Y (nx7285), .A0 (que_out_12__4__7), .A1 (nx9676), .B0 (
          que_out_1__4__7), .B1 (nx9650)) ;
    or04 ix1123 (.Y (out_column_4__8), .A0 (nx1118), .A1 (nx1092), .A2 (nx1064)
         , .A3 (nx1038)) ;
    nand03 ix1119 (.Y (nx1118), .A0 (nx7291), .A1 (nx7293), .A2 (nx7295)) ;
    aoi222 ix7292 (.Y (nx7291), .A0 (que_out_10__4__8), .A1 (nx10300), .B0 (
           que_out_6__4__8), .B1 (nx10352), .C0 (que_out_9__4__8), .C1 (nx10326)
           ) ;
    aoi22 ix7294 (.Y (nx7293), .A0 (que_out_5__4__8), .A1 (nx10248), .B0 (
          que_out_18__4__8), .B1 (nx10274)) ;
    aoi22 ix7296 (.Y (nx7295), .A0 (que_out_17__4__8), .A1 (nx10222), .B0 (
          que_out_20__4__8), .B1 (nx10196)) ;
    nand03 ix1093 (.Y (nx1092), .A0 (nx7299), .A1 (nx7301), .A2 (nx7303)) ;
    aoi222 ix7300 (.Y (nx7299), .A0 (que_out_19__4__8), .A1 (nx10170), .B0 (
           que_out_21__4__8), .B1 (nx10144), .C0 (que_out_8__4__8), .C1 (nx10118
           )) ;
    aoi22 ix7302 (.Y (nx7301), .A0 (que_out_25__4__8), .A1 (nx10066), .B0 (
          que_out_16__4__8), .B1 (nx10092)) ;
    aoi22 ix7304 (.Y (nx7303), .A0 (que_out_24__4__8), .A1 (nx10040), .B0 (
          que_out_22__4__8), .B1 (nx10014)) ;
    nand03 ix1065 (.Y (nx1064), .A0 (nx7307), .A1 (nx7309), .A2 (nx7311)) ;
    aoi222 ix7308 (.Y (nx7307), .A0 (que_out_15__4__8), .A1 (nx9962), .B0 (
           que_out_3__4__8), .B1 (nx9988), .C0 (que_out_23__4__8), .C1 (nx9936)
           ) ;
    aoi22 ix7310 (.Y (nx7309), .A0 (que_out_27__4__8), .A1 (nx9910), .B0 (
          que_out_4__4__8), .B1 (nx9884)) ;
    aoi22 ix7312 (.Y (nx7311), .A0 (que_out_0__4__8), .A1 (nx9832), .B0 (
          que_out_2__4__8), .B1 (nx9858)) ;
    nand03 ix1039 (.Y (nx1038), .A0 (nx7315), .A1 (nx7317), .A2 (nx7319)) ;
    aoi222 ix7316 (.Y (nx7315), .A0 (que_out_26__4__8), .A1 (nx9806), .B0 (
           que_out_14__4__8), .B1 (nx9780), .C0 (que_out_11__4__8), .C1 (nx9754)
           ) ;
    aoi22 ix7318 (.Y (nx7317), .A0 (que_out_13__4__8), .A1 (nx9728), .B0 (
          que_out_7__4__8), .B1 (nx9702)) ;
    aoi22 ix7320 (.Y (nx7319), .A0 (que_out_12__4__8), .A1 (nx9676), .B0 (
          que_out_1__4__8), .B1 (nx9650)) ;
    or04 ix1233 (.Y (out_column_4__9), .A0 (nx1228), .A1 (nx1202), .A2 (nx1174)
         , .A3 (nx1148)) ;
    nand03 ix1229 (.Y (nx1228), .A0 (nx7325), .A1 (nx7327), .A2 (nx7329)) ;
    aoi222 ix7326 (.Y (nx7325), .A0 (que_out_10__4__9), .A1 (nx10300), .B0 (
           que_out_6__4__9), .B1 (nx10352), .C0 (que_out_9__4__9), .C1 (nx10326)
           ) ;
    aoi22 ix7328 (.Y (nx7327), .A0 (que_out_5__4__9), .A1 (nx10248), .B0 (
          que_out_18__4__9), .B1 (nx10274)) ;
    aoi22 ix7330 (.Y (nx7329), .A0 (que_out_17__4__9), .A1 (nx10222), .B0 (
          que_out_20__4__9), .B1 (nx10196)) ;
    nand03 ix1203 (.Y (nx1202), .A0 (nx7333), .A1 (nx7335), .A2 (nx7337)) ;
    aoi222 ix7334 (.Y (nx7333), .A0 (que_out_19__4__9), .A1 (nx10170), .B0 (
           que_out_21__4__9), .B1 (nx10144), .C0 (que_out_8__4__9), .C1 (nx10118
           )) ;
    aoi22 ix7336 (.Y (nx7335), .A0 (que_out_25__4__9), .A1 (nx10066), .B0 (
          que_out_16__4__9), .B1 (nx10092)) ;
    aoi22 ix7338 (.Y (nx7337), .A0 (que_out_24__4__9), .A1 (nx10040), .B0 (
          que_out_22__4__9), .B1 (nx10014)) ;
    nand03 ix1175 (.Y (nx1174), .A0 (nx7341), .A1 (nx7343), .A2 (nx7345)) ;
    aoi222 ix7342 (.Y (nx7341), .A0 (que_out_15__4__9), .A1 (nx9962), .B0 (
           que_out_3__4__9), .B1 (nx9988), .C0 (que_out_23__4__9), .C1 (nx9936)
           ) ;
    aoi22 ix7344 (.Y (nx7343), .A0 (que_out_27__4__9), .A1 (nx9910), .B0 (
          que_out_4__4__9), .B1 (nx9884)) ;
    aoi22 ix7346 (.Y (nx7345), .A0 (que_out_0__4__9), .A1 (nx9832), .B0 (
          que_out_2__4__9), .B1 (nx9858)) ;
    nand03 ix1149 (.Y (nx1148), .A0 (nx7349), .A1 (nx7351), .A2 (nx7353)) ;
    aoi222 ix7350 (.Y (nx7349), .A0 (que_out_26__4__9), .A1 (nx9806), .B0 (
           que_out_14__4__9), .B1 (nx9780), .C0 (que_out_11__4__9), .C1 (nx9754)
           ) ;
    aoi22 ix7352 (.Y (nx7351), .A0 (que_out_13__4__9), .A1 (nx9728), .B0 (
          que_out_7__4__9), .B1 (nx9702)) ;
    aoi22 ix7354 (.Y (nx7353), .A0 (que_out_12__4__9), .A1 (nx9676), .B0 (
          que_out_1__4__9), .B1 (nx9650)) ;
    or04 ix1343 (.Y (out_column_4__10), .A0 (nx1338), .A1 (nx1312), .A2 (nx1284)
         , .A3 (nx1258)) ;
    nand03 ix1339 (.Y (nx1338), .A0 (nx7359), .A1 (nx7361), .A2 (nx7363)) ;
    aoi222 ix7360 (.Y (nx7359), .A0 (que_out_10__4__10), .A1 (nx10300), .B0 (
           que_out_6__4__10), .B1 (nx10352), .C0 (que_out_9__4__10), .C1 (
           nx10326)) ;
    aoi22 ix7362 (.Y (nx7361), .A0 (que_out_5__4__10), .A1 (nx10248), .B0 (
          que_out_18__4__10), .B1 (nx10274)) ;
    aoi22 ix7364 (.Y (nx7363), .A0 (que_out_17__4__10), .A1 (nx10222), .B0 (
          que_out_20__4__10), .B1 (nx10196)) ;
    nand03 ix1313 (.Y (nx1312), .A0 (nx7367), .A1 (nx7369), .A2 (nx7371)) ;
    aoi222 ix7368 (.Y (nx7367), .A0 (que_out_19__4__10), .A1 (nx10170), .B0 (
           que_out_21__4__10), .B1 (nx10144), .C0 (que_out_8__4__10), .C1 (
           nx10118)) ;
    aoi22 ix7370 (.Y (nx7369), .A0 (que_out_25__4__10), .A1 (nx10066), .B0 (
          que_out_16__4__10), .B1 (nx10092)) ;
    aoi22 ix7372 (.Y (nx7371), .A0 (que_out_24__4__10), .A1 (nx10040), .B0 (
          que_out_22__4__10), .B1 (nx10014)) ;
    nand03 ix1285 (.Y (nx1284), .A0 (nx7375), .A1 (nx7377), .A2 (nx7379)) ;
    aoi222 ix7376 (.Y (nx7375), .A0 (que_out_15__4__10), .A1 (nx9962), .B0 (
           que_out_3__4__10), .B1 (nx9988), .C0 (que_out_23__4__10), .C1 (nx9936
           )) ;
    aoi22 ix7378 (.Y (nx7377), .A0 (que_out_27__4__10), .A1 (nx9910), .B0 (
          que_out_4__4__10), .B1 (nx9884)) ;
    aoi22 ix7380 (.Y (nx7379), .A0 (que_out_0__4__10), .A1 (nx9832), .B0 (
          que_out_2__4__10), .B1 (nx9858)) ;
    nand03 ix1259 (.Y (nx1258), .A0 (nx7383), .A1 (nx7385), .A2 (nx7387)) ;
    aoi222 ix7384 (.Y (nx7383), .A0 (que_out_26__4__10), .A1 (nx9806), .B0 (
           que_out_14__4__10), .B1 (nx9780), .C0 (que_out_11__4__10), .C1 (
           nx9754)) ;
    aoi22 ix7386 (.Y (nx7385), .A0 (que_out_13__4__10), .A1 (nx9728), .B0 (
          que_out_7__4__10), .B1 (nx9702)) ;
    aoi22 ix7388 (.Y (nx7387), .A0 (que_out_12__4__10), .A1 (nx9676), .B0 (
          que_out_1__4__10), .B1 (nx9650)) ;
    or04 ix1453 (.Y (out_column_4__11), .A0 (nx1448), .A1 (nx1422), .A2 (nx1394)
         , .A3 (nx1368)) ;
    nand03 ix1449 (.Y (nx1448), .A0 (nx7393), .A1 (nx7395), .A2 (nx7397)) ;
    aoi222 ix7394 (.Y (nx7393), .A0 (que_out_10__4__11), .A1 (nx10300), .B0 (
           que_out_6__4__11), .B1 (nx10352), .C0 (que_out_9__4__11), .C1 (
           nx10326)) ;
    aoi22 ix7396 (.Y (nx7395), .A0 (que_out_5__4__11), .A1 (nx10248), .B0 (
          que_out_18__4__11), .B1 (nx10274)) ;
    aoi22 ix7398 (.Y (nx7397), .A0 (que_out_17__4__11), .A1 (nx10222), .B0 (
          que_out_20__4__11), .B1 (nx10196)) ;
    nand03 ix1423 (.Y (nx1422), .A0 (nx7401), .A1 (nx7403), .A2 (nx7405)) ;
    aoi222 ix7402 (.Y (nx7401), .A0 (que_out_19__4__11), .A1 (nx10170), .B0 (
           que_out_21__4__11), .B1 (nx10144), .C0 (que_out_8__4__11), .C1 (
           nx10118)) ;
    aoi22 ix7404 (.Y (nx7403), .A0 (que_out_25__4__11), .A1 (nx10066), .B0 (
          que_out_16__4__11), .B1 (nx10092)) ;
    aoi22 ix7406 (.Y (nx7405), .A0 (que_out_24__4__11), .A1 (nx10040), .B0 (
          que_out_22__4__11), .B1 (nx10014)) ;
    nand03 ix1395 (.Y (nx1394), .A0 (nx7409), .A1 (nx7411), .A2 (nx7413)) ;
    aoi222 ix7410 (.Y (nx7409), .A0 (que_out_15__4__11), .A1 (nx9962), .B0 (
           que_out_3__4__11), .B1 (nx9988), .C0 (que_out_23__4__11), .C1 (nx9936
           )) ;
    aoi22 ix7412 (.Y (nx7411), .A0 (que_out_27__4__11), .A1 (nx9910), .B0 (
          que_out_4__4__11), .B1 (nx9884)) ;
    aoi22 ix7414 (.Y (nx7413), .A0 (que_out_0__4__11), .A1 (nx9832), .B0 (
          que_out_2__4__11), .B1 (nx9858)) ;
    nand03 ix1369 (.Y (nx1368), .A0 (nx7417), .A1 (nx7419), .A2 (nx7421)) ;
    aoi222 ix7418 (.Y (nx7417), .A0 (que_out_26__4__11), .A1 (nx9806), .B0 (
           que_out_14__4__11), .B1 (nx9780), .C0 (que_out_11__4__11), .C1 (
           nx9754)) ;
    aoi22 ix7420 (.Y (nx7419), .A0 (que_out_13__4__11), .A1 (nx9728), .B0 (
          que_out_7__4__11), .B1 (nx9702)) ;
    aoi22 ix7422 (.Y (nx7421), .A0 (que_out_12__4__11), .A1 (nx9676), .B0 (
          que_out_1__4__11), .B1 (nx9650)) ;
    or04 ix1563 (.Y (out_column_4__12), .A0 (nx1558), .A1 (nx1532), .A2 (nx1504)
         , .A3 (nx1478)) ;
    nand03 ix1559 (.Y (nx1558), .A0 (nx7427), .A1 (nx7429), .A2 (nx7431)) ;
    aoi222 ix7428 (.Y (nx7427), .A0 (que_out_10__4__12), .A1 (nx10300), .B0 (
           que_out_6__4__12), .B1 (nx10352), .C0 (que_out_9__4__12), .C1 (
           nx10326)) ;
    aoi22 ix7430 (.Y (nx7429), .A0 (que_out_5__4__12), .A1 (nx10248), .B0 (
          que_out_18__4__12), .B1 (nx10274)) ;
    aoi22 ix7432 (.Y (nx7431), .A0 (que_out_17__4__12), .A1 (nx10222), .B0 (
          que_out_20__4__12), .B1 (nx10196)) ;
    nand03 ix1533 (.Y (nx1532), .A0 (nx7435), .A1 (nx7437), .A2 (nx7439)) ;
    aoi222 ix7436 (.Y (nx7435), .A0 (que_out_19__4__12), .A1 (nx10170), .B0 (
           que_out_21__4__12), .B1 (nx10144), .C0 (que_out_8__4__12), .C1 (
           nx10118)) ;
    aoi22 ix7438 (.Y (nx7437), .A0 (que_out_25__4__12), .A1 (nx10066), .B0 (
          que_out_16__4__12), .B1 (nx10092)) ;
    aoi22 ix7440 (.Y (nx7439), .A0 (que_out_24__4__12), .A1 (nx10040), .B0 (
          que_out_22__4__12), .B1 (nx10014)) ;
    nand03 ix1505 (.Y (nx1504), .A0 (nx7443), .A1 (nx7445), .A2 (nx7447)) ;
    aoi222 ix7444 (.Y (nx7443), .A0 (que_out_15__4__12), .A1 (nx9962), .B0 (
           que_out_3__4__12), .B1 (nx9988), .C0 (que_out_23__4__12), .C1 (nx9936
           )) ;
    aoi22 ix7446 (.Y (nx7445), .A0 (que_out_27__4__12), .A1 (nx9910), .B0 (
          que_out_4__4__12), .B1 (nx9884)) ;
    aoi22 ix7448 (.Y (nx7447), .A0 (que_out_0__4__12), .A1 (nx9832), .B0 (
          que_out_2__4__12), .B1 (nx9858)) ;
    nand03 ix1479 (.Y (nx1478), .A0 (nx7451), .A1 (nx7453), .A2 (nx7455)) ;
    aoi222 ix7452 (.Y (nx7451), .A0 (que_out_26__4__12), .A1 (nx9806), .B0 (
           que_out_14__4__12), .B1 (nx9780), .C0 (que_out_11__4__12), .C1 (
           nx9754)) ;
    aoi22 ix7454 (.Y (nx7453), .A0 (que_out_13__4__12), .A1 (nx9728), .B0 (
          que_out_7__4__12), .B1 (nx9702)) ;
    aoi22 ix7456 (.Y (nx7455), .A0 (que_out_12__4__12), .A1 (nx9676), .B0 (
          que_out_1__4__12), .B1 (nx9650)) ;
    or04 ix1673 (.Y (out_column_4__13), .A0 (nx1668), .A1 (nx1642), .A2 (nx1614)
         , .A3 (nx1588)) ;
    nand03 ix1669 (.Y (nx1668), .A0 (nx7461), .A1 (nx7463), .A2 (nx7465)) ;
    aoi222 ix7462 (.Y (nx7461), .A0 (que_out_10__4__13), .A1 (nx10300), .B0 (
           que_out_6__4__13), .B1 (nx10352), .C0 (que_out_9__4__13), .C1 (
           nx10326)) ;
    aoi22 ix7464 (.Y (nx7463), .A0 (que_out_5__4__13), .A1 (nx10248), .B0 (
          que_out_18__4__13), .B1 (nx10274)) ;
    aoi22 ix7466 (.Y (nx7465), .A0 (que_out_17__4__13), .A1 (nx10222), .B0 (
          que_out_20__4__13), .B1 (nx10196)) ;
    nand03 ix1643 (.Y (nx1642), .A0 (nx7469), .A1 (nx7471), .A2 (nx7473)) ;
    aoi222 ix7470 (.Y (nx7469), .A0 (que_out_19__4__13), .A1 (nx10170), .B0 (
           que_out_21__4__13), .B1 (nx10144), .C0 (que_out_8__4__13), .C1 (
           nx10118)) ;
    aoi22 ix7472 (.Y (nx7471), .A0 (que_out_25__4__13), .A1 (nx10066), .B0 (
          que_out_16__4__13), .B1 (nx10092)) ;
    aoi22 ix7474 (.Y (nx7473), .A0 (que_out_24__4__13), .A1 (nx10040), .B0 (
          que_out_22__4__13), .B1 (nx10014)) ;
    nand03 ix1615 (.Y (nx1614), .A0 (nx7477), .A1 (nx7479), .A2 (nx7481)) ;
    aoi222 ix7478 (.Y (nx7477), .A0 (que_out_15__4__13), .A1 (nx9962), .B0 (
           que_out_3__4__13), .B1 (nx9988), .C0 (que_out_23__4__13), .C1 (nx9936
           )) ;
    aoi22 ix7480 (.Y (nx7479), .A0 (que_out_27__4__13), .A1 (nx9910), .B0 (
          que_out_4__4__13), .B1 (nx9884)) ;
    aoi22 ix7482 (.Y (nx7481), .A0 (que_out_0__4__13), .A1 (nx9832), .B0 (
          que_out_2__4__13), .B1 (nx9858)) ;
    nand03 ix1589 (.Y (nx1588), .A0 (nx7485), .A1 (nx7487), .A2 (nx7489)) ;
    aoi222 ix7486 (.Y (nx7485), .A0 (que_out_26__4__13), .A1 (nx9806), .B0 (
           que_out_14__4__13), .B1 (nx9780), .C0 (que_out_11__4__13), .C1 (
           nx9754)) ;
    aoi22 ix7488 (.Y (nx7487), .A0 (que_out_13__4__13), .A1 (nx9728), .B0 (
          que_out_7__4__13), .B1 (nx9702)) ;
    aoi22 ix7490 (.Y (nx7489), .A0 (que_out_12__4__13), .A1 (nx9676), .B0 (
          que_out_1__4__13), .B1 (nx9650)) ;
    or04 ix1783 (.Y (out_column_4__14), .A0 (nx1778), .A1 (nx1752), .A2 (nx1724)
         , .A3 (nx1698)) ;
    nand03 ix1779 (.Y (nx1778), .A0 (nx7495), .A1 (nx7497), .A2 (nx7499)) ;
    aoi222 ix7496 (.Y (nx7495), .A0 (que_out_10__4__14), .A1 (nx10302), .B0 (
           que_out_6__4__14), .B1 (nx10354), .C0 (que_out_9__4__14), .C1 (
           nx10328)) ;
    aoi22 ix7498 (.Y (nx7497), .A0 (que_out_5__4__14), .A1 (nx10250), .B0 (
          que_out_18__4__14), .B1 (nx10276)) ;
    aoi22 ix7500 (.Y (nx7499), .A0 (que_out_17__4__14), .A1 (nx10224), .B0 (
          que_out_20__4__14), .B1 (nx10198)) ;
    nand03 ix1753 (.Y (nx1752), .A0 (nx7503), .A1 (nx7505), .A2 (nx7507)) ;
    aoi222 ix7504 (.Y (nx7503), .A0 (que_out_19__4__14), .A1 (nx10172), .B0 (
           que_out_21__4__14), .B1 (nx10146), .C0 (que_out_8__4__14), .C1 (
           nx10120)) ;
    aoi22 ix7506 (.Y (nx7505), .A0 (que_out_25__4__14), .A1 (nx10068), .B0 (
          que_out_16__4__14), .B1 (nx10094)) ;
    aoi22 ix7508 (.Y (nx7507), .A0 (que_out_24__4__14), .A1 (nx10042), .B0 (
          que_out_22__4__14), .B1 (nx10016)) ;
    nand03 ix1725 (.Y (nx1724), .A0 (nx7511), .A1 (nx7513), .A2 (nx7515)) ;
    aoi222 ix7512 (.Y (nx7511), .A0 (que_out_15__4__14), .A1 (nx9964), .B0 (
           que_out_3__4__14), .B1 (nx9990), .C0 (que_out_23__4__14), .C1 (nx9938
           )) ;
    aoi22 ix7514 (.Y (nx7513), .A0 (que_out_27__4__14), .A1 (nx9912), .B0 (
          que_out_4__4__14), .B1 (nx9886)) ;
    aoi22 ix7516 (.Y (nx7515), .A0 (que_out_0__4__14), .A1 (nx9834), .B0 (
          que_out_2__4__14), .B1 (nx9860)) ;
    nand03 ix1699 (.Y (nx1698), .A0 (nx7519), .A1 (nx7521), .A2 (nx7523)) ;
    aoi222 ix7520 (.Y (nx7519), .A0 (que_out_26__4__14), .A1 (nx9808), .B0 (
           que_out_14__4__14), .B1 (nx9782), .C0 (que_out_11__4__14), .C1 (
           nx9756)) ;
    aoi22 ix7522 (.Y (nx7521), .A0 (que_out_13__4__14), .A1 (nx9730), .B0 (
          que_out_7__4__14), .B1 (nx9704)) ;
    aoi22 ix7524 (.Y (nx7523), .A0 (que_out_12__4__14), .A1 (nx9678), .B0 (
          que_out_1__4__14), .B1 (nx9652)) ;
    or04 ix1893 (.Y (out_column_4__15), .A0 (nx1888), .A1 (nx1862), .A2 (nx1834)
         , .A3 (nx1808)) ;
    nand03 ix1889 (.Y (nx1888), .A0 (nx7529), .A1 (nx7531), .A2 (nx7533)) ;
    aoi222 ix7530 (.Y (nx7529), .A0 (que_out_10__4__15), .A1 (nx10302), .B0 (
           que_out_6__4__15), .B1 (nx10354), .C0 (que_out_9__4__15), .C1 (
           nx10328)) ;
    aoi22 ix7532 (.Y (nx7531), .A0 (que_out_5__4__15), .A1 (nx10250), .B0 (
          que_out_18__4__15), .B1 (nx10276)) ;
    aoi22 ix7534 (.Y (nx7533), .A0 (que_out_17__4__15), .A1 (nx10224), .B0 (
          que_out_20__4__15), .B1 (nx10198)) ;
    nand03 ix1863 (.Y (nx1862), .A0 (nx7537), .A1 (nx7539), .A2 (nx7541)) ;
    aoi222 ix7538 (.Y (nx7537), .A0 (que_out_19__4__15), .A1 (nx10172), .B0 (
           que_out_21__4__15), .B1 (nx10146), .C0 (que_out_8__4__15), .C1 (
           nx10120)) ;
    aoi22 ix7540 (.Y (nx7539), .A0 (que_out_25__4__15), .A1 (nx10068), .B0 (
          que_out_16__4__15), .B1 (nx10094)) ;
    aoi22 ix7542 (.Y (nx7541), .A0 (que_out_24__4__15), .A1 (nx10042), .B0 (
          que_out_22__4__15), .B1 (nx10016)) ;
    nand03 ix1835 (.Y (nx1834), .A0 (nx7545), .A1 (nx7547), .A2 (nx7549)) ;
    aoi222 ix7546 (.Y (nx7545), .A0 (que_out_15__4__15), .A1 (nx9964), .B0 (
           que_out_3__4__15), .B1 (nx9990), .C0 (que_out_23__4__15), .C1 (nx9938
           )) ;
    aoi22 ix7548 (.Y (nx7547), .A0 (que_out_27__4__15), .A1 (nx9912), .B0 (
          que_out_4__4__15), .B1 (nx9886)) ;
    aoi22 ix7550 (.Y (nx7549), .A0 (que_out_0__4__15), .A1 (nx9834), .B0 (
          que_out_2__4__15), .B1 (nx9860)) ;
    nand03 ix1809 (.Y (nx1808), .A0 (nx7553), .A1 (nx7555), .A2 (nx7557)) ;
    aoi222 ix7554 (.Y (nx7553), .A0 (que_out_26__4__15), .A1 (nx9808), .B0 (
           que_out_14__4__15), .B1 (nx9782), .C0 (que_out_11__4__15), .C1 (
           nx9756)) ;
    aoi22 ix7556 (.Y (nx7555), .A0 (que_out_13__4__15), .A1 (nx9730), .B0 (
          que_out_7__4__15), .B1 (nx9704)) ;
    aoi22 ix7558 (.Y (nx7557), .A0 (que_out_12__4__15), .A1 (nx9678), .B0 (
          que_out_1__4__15), .B1 (nx9652)) ;
    or04 ix2003 (.Y (out_column_3__0), .A0 (nx1998), .A1 (nx1972), .A2 (nx1944)
         , .A3 (nx1918)) ;
    nand03 ix1999 (.Y (nx1998), .A0 (nx7563), .A1 (nx7565), .A2 (nx7567)) ;
    aoi222 ix7564 (.Y (nx7563), .A0 (que_out_10__3__0), .A1 (nx10302), .B0 (
           que_out_6__3__0), .B1 (nx10354), .C0 (que_out_9__3__0), .C1 (nx10328)
           ) ;
    aoi22 ix7566 (.Y (nx7565), .A0 (que_out_5__3__0), .A1 (nx10250), .B0 (
          que_out_18__3__0), .B1 (nx10276)) ;
    aoi22 ix7568 (.Y (nx7567), .A0 (que_out_17__3__0), .A1 (nx10224), .B0 (
          que_out_20__3__0), .B1 (nx10198)) ;
    nand03 ix1973 (.Y (nx1972), .A0 (nx7571), .A1 (nx7573), .A2 (nx7575)) ;
    aoi222 ix7572 (.Y (nx7571), .A0 (que_out_19__3__0), .A1 (nx10172), .B0 (
           que_out_21__3__0), .B1 (nx10146), .C0 (que_out_8__3__0), .C1 (nx10120
           )) ;
    aoi22 ix7574 (.Y (nx7573), .A0 (que_out_25__3__0), .A1 (nx10068), .B0 (
          que_out_16__3__0), .B1 (nx10094)) ;
    aoi22 ix7576 (.Y (nx7575), .A0 (que_out_24__3__0), .A1 (nx10042), .B0 (
          que_out_22__3__0), .B1 (nx10016)) ;
    nand03 ix1945 (.Y (nx1944), .A0 (nx7579), .A1 (nx7581), .A2 (nx7583)) ;
    aoi222 ix7580 (.Y (nx7579), .A0 (que_out_15__3__0), .A1 (nx9964), .B0 (
           que_out_3__3__0), .B1 (nx9990), .C0 (que_out_23__3__0), .C1 (nx9938)
           ) ;
    aoi22 ix7582 (.Y (nx7581), .A0 (que_out_27__3__0), .A1 (nx9912), .B0 (
          que_out_4__3__0), .B1 (nx9886)) ;
    aoi22 ix7584 (.Y (nx7583), .A0 (que_out_0__3__0), .A1 (nx9834), .B0 (
          que_out_2__3__0), .B1 (nx9860)) ;
    nand03 ix1919 (.Y (nx1918), .A0 (nx7587), .A1 (nx7589), .A2 (nx7591)) ;
    aoi222 ix7588 (.Y (nx7587), .A0 (que_out_26__3__0), .A1 (nx9808), .B0 (
           que_out_14__3__0), .B1 (nx9782), .C0 (que_out_11__3__0), .C1 (nx9756)
           ) ;
    aoi22 ix7590 (.Y (nx7589), .A0 (que_out_13__3__0), .A1 (nx9730), .B0 (
          que_out_7__3__0), .B1 (nx9704)) ;
    aoi22 ix7592 (.Y (nx7591), .A0 (que_out_12__3__0), .A1 (nx9678), .B0 (
          que_out_1__3__0), .B1 (nx9652)) ;
    or04 ix2113 (.Y (out_column_3__1), .A0 (nx2108), .A1 (nx2082), .A2 (nx2054)
         , .A3 (nx2028)) ;
    nand03 ix2109 (.Y (nx2108), .A0 (nx7597), .A1 (nx7599), .A2 (nx7601)) ;
    aoi222 ix7598 (.Y (nx7597), .A0 (que_out_10__3__1), .A1 (nx10302), .B0 (
           que_out_6__3__1), .B1 (nx10354), .C0 (que_out_9__3__1), .C1 (nx10328)
           ) ;
    aoi22 ix7600 (.Y (nx7599), .A0 (que_out_5__3__1), .A1 (nx10250), .B0 (
          que_out_18__3__1), .B1 (nx10276)) ;
    aoi22 ix7602 (.Y (nx7601), .A0 (que_out_17__3__1), .A1 (nx10224), .B0 (
          que_out_20__3__1), .B1 (nx10198)) ;
    nand03 ix2083 (.Y (nx2082), .A0 (nx7605), .A1 (nx7607), .A2 (nx7609)) ;
    aoi222 ix7606 (.Y (nx7605), .A0 (que_out_19__3__1), .A1 (nx10172), .B0 (
           que_out_21__3__1), .B1 (nx10146), .C0 (que_out_8__3__1), .C1 (nx10120
           )) ;
    aoi22 ix7608 (.Y (nx7607), .A0 (que_out_25__3__1), .A1 (nx10068), .B0 (
          que_out_16__3__1), .B1 (nx10094)) ;
    aoi22 ix7610 (.Y (nx7609), .A0 (que_out_24__3__1), .A1 (nx10042), .B0 (
          que_out_22__3__1), .B1 (nx10016)) ;
    nand03 ix2055 (.Y (nx2054), .A0 (nx7613), .A1 (nx7615), .A2 (nx7617)) ;
    aoi222 ix7614 (.Y (nx7613), .A0 (que_out_15__3__1), .A1 (nx9964), .B0 (
           que_out_3__3__1), .B1 (nx9990), .C0 (que_out_23__3__1), .C1 (nx9938)
           ) ;
    aoi22 ix7616 (.Y (nx7615), .A0 (que_out_27__3__1), .A1 (nx9912), .B0 (
          que_out_4__3__1), .B1 (nx9886)) ;
    aoi22 ix7618 (.Y (nx7617), .A0 (que_out_0__3__1), .A1 (nx9834), .B0 (
          que_out_2__3__1), .B1 (nx9860)) ;
    nand03 ix2029 (.Y (nx2028), .A0 (nx7621), .A1 (nx7623), .A2 (nx7625)) ;
    aoi222 ix7622 (.Y (nx7621), .A0 (que_out_26__3__1), .A1 (nx9808), .B0 (
           que_out_14__3__1), .B1 (nx9782), .C0 (que_out_11__3__1), .C1 (nx9756)
           ) ;
    aoi22 ix7624 (.Y (nx7623), .A0 (que_out_13__3__1), .A1 (nx9730), .B0 (
          que_out_7__3__1), .B1 (nx9704)) ;
    aoi22 ix7626 (.Y (nx7625), .A0 (que_out_12__3__1), .A1 (nx9678), .B0 (
          que_out_1__3__1), .B1 (nx9652)) ;
    or04 ix2223 (.Y (out_column_3__2), .A0 (nx2218), .A1 (nx2192), .A2 (nx2164)
         , .A3 (nx2138)) ;
    nand03 ix2219 (.Y (nx2218), .A0 (nx7631), .A1 (nx7633), .A2 (nx7635)) ;
    aoi222 ix7632 (.Y (nx7631), .A0 (que_out_10__3__2), .A1 (nx10302), .B0 (
           que_out_6__3__2), .B1 (nx10354), .C0 (que_out_9__3__2), .C1 (nx10328)
           ) ;
    aoi22 ix7634 (.Y (nx7633), .A0 (que_out_5__3__2), .A1 (nx10250), .B0 (
          que_out_18__3__2), .B1 (nx10276)) ;
    aoi22 ix7636 (.Y (nx7635), .A0 (que_out_17__3__2), .A1 (nx10224), .B0 (
          que_out_20__3__2), .B1 (nx10198)) ;
    nand03 ix2193 (.Y (nx2192), .A0 (nx7639), .A1 (nx7641), .A2 (nx7643)) ;
    aoi222 ix7640 (.Y (nx7639), .A0 (que_out_19__3__2), .A1 (nx10172), .B0 (
           que_out_21__3__2), .B1 (nx10146), .C0 (que_out_8__3__2), .C1 (nx10120
           )) ;
    aoi22 ix7642 (.Y (nx7641), .A0 (que_out_25__3__2), .A1 (nx10068), .B0 (
          que_out_16__3__2), .B1 (nx10094)) ;
    aoi22 ix7644 (.Y (nx7643), .A0 (que_out_24__3__2), .A1 (nx10042), .B0 (
          que_out_22__3__2), .B1 (nx10016)) ;
    nand03 ix2165 (.Y (nx2164), .A0 (nx7647), .A1 (nx7649), .A2 (nx7651)) ;
    aoi222 ix7648 (.Y (nx7647), .A0 (que_out_15__3__2), .A1 (nx9964), .B0 (
           que_out_3__3__2), .B1 (nx9990), .C0 (que_out_23__3__2), .C1 (nx9938)
           ) ;
    aoi22 ix7650 (.Y (nx7649), .A0 (que_out_27__3__2), .A1 (nx9912), .B0 (
          que_out_4__3__2), .B1 (nx9886)) ;
    aoi22 ix7652 (.Y (nx7651), .A0 (que_out_0__3__2), .A1 (nx9834), .B0 (
          que_out_2__3__2), .B1 (nx9860)) ;
    nand03 ix2139 (.Y (nx2138), .A0 (nx7655), .A1 (nx7657), .A2 (nx7659)) ;
    aoi222 ix7656 (.Y (nx7655), .A0 (que_out_26__3__2), .A1 (nx9808), .B0 (
           que_out_14__3__2), .B1 (nx9782), .C0 (que_out_11__3__2), .C1 (nx9756)
           ) ;
    aoi22 ix7658 (.Y (nx7657), .A0 (que_out_13__3__2), .A1 (nx9730), .B0 (
          que_out_7__3__2), .B1 (nx9704)) ;
    aoi22 ix7660 (.Y (nx7659), .A0 (que_out_12__3__2), .A1 (nx9678), .B0 (
          que_out_1__3__2), .B1 (nx9652)) ;
    or04 ix2333 (.Y (out_column_3__3), .A0 (nx2328), .A1 (nx2302), .A2 (nx2274)
         , .A3 (nx2248)) ;
    nand03 ix2329 (.Y (nx2328), .A0 (nx7665), .A1 (nx7667), .A2 (nx7669)) ;
    aoi222 ix7666 (.Y (nx7665), .A0 (que_out_10__3__3), .A1 (nx10302), .B0 (
           que_out_6__3__3), .B1 (nx10354), .C0 (que_out_9__3__3), .C1 (nx10328)
           ) ;
    aoi22 ix7668 (.Y (nx7667), .A0 (que_out_5__3__3), .A1 (nx10250), .B0 (
          que_out_18__3__3), .B1 (nx10276)) ;
    aoi22 ix7670 (.Y (nx7669), .A0 (que_out_17__3__3), .A1 (nx10224), .B0 (
          que_out_20__3__3), .B1 (nx10198)) ;
    nand03 ix2303 (.Y (nx2302), .A0 (nx7673), .A1 (nx7675), .A2 (nx7677)) ;
    aoi222 ix7674 (.Y (nx7673), .A0 (que_out_19__3__3), .A1 (nx10172), .B0 (
           que_out_21__3__3), .B1 (nx10146), .C0 (que_out_8__3__3), .C1 (nx10120
           )) ;
    aoi22 ix7676 (.Y (nx7675), .A0 (que_out_25__3__3), .A1 (nx10068), .B0 (
          que_out_16__3__3), .B1 (nx10094)) ;
    aoi22 ix7678 (.Y (nx7677), .A0 (que_out_24__3__3), .A1 (nx10042), .B0 (
          que_out_22__3__3), .B1 (nx10016)) ;
    nand03 ix2275 (.Y (nx2274), .A0 (nx7681), .A1 (nx7683), .A2 (nx7685)) ;
    aoi222 ix7682 (.Y (nx7681), .A0 (que_out_15__3__3), .A1 (nx9964), .B0 (
           que_out_3__3__3), .B1 (nx9990), .C0 (que_out_23__3__3), .C1 (nx9938)
           ) ;
    aoi22 ix7684 (.Y (nx7683), .A0 (que_out_27__3__3), .A1 (nx9912), .B0 (
          que_out_4__3__3), .B1 (nx9886)) ;
    aoi22 ix7686 (.Y (nx7685), .A0 (que_out_0__3__3), .A1 (nx9834), .B0 (
          que_out_2__3__3), .B1 (nx9860)) ;
    nand03 ix2249 (.Y (nx2248), .A0 (nx7689), .A1 (nx7691), .A2 (nx7693)) ;
    aoi222 ix7690 (.Y (nx7689), .A0 (que_out_26__3__3), .A1 (nx9808), .B0 (
           que_out_14__3__3), .B1 (nx9782), .C0 (que_out_11__3__3), .C1 (nx9756)
           ) ;
    aoi22 ix7692 (.Y (nx7691), .A0 (que_out_13__3__3), .A1 (nx9730), .B0 (
          que_out_7__3__3), .B1 (nx9704)) ;
    aoi22 ix7694 (.Y (nx7693), .A0 (que_out_12__3__3), .A1 (nx9678), .B0 (
          que_out_1__3__3), .B1 (nx9652)) ;
    or04 ix2443 (.Y (out_column_3__4), .A0 (nx2438), .A1 (nx2412), .A2 (nx2384)
         , .A3 (nx2358)) ;
    nand03 ix2439 (.Y (nx2438), .A0 (nx7699), .A1 (nx7701), .A2 (nx7703)) ;
    aoi222 ix7700 (.Y (nx7699), .A0 (que_out_10__3__4), .A1 (nx10302), .B0 (
           que_out_6__3__4), .B1 (nx10354), .C0 (que_out_9__3__4), .C1 (nx10328)
           ) ;
    aoi22 ix7702 (.Y (nx7701), .A0 (que_out_5__3__4), .A1 (nx10250), .B0 (
          que_out_18__3__4), .B1 (nx10276)) ;
    aoi22 ix7704 (.Y (nx7703), .A0 (que_out_17__3__4), .A1 (nx10224), .B0 (
          que_out_20__3__4), .B1 (nx10198)) ;
    nand03 ix2413 (.Y (nx2412), .A0 (nx7707), .A1 (nx7709), .A2 (nx7711)) ;
    aoi222 ix7708 (.Y (nx7707), .A0 (que_out_19__3__4), .A1 (nx10172), .B0 (
           que_out_21__3__4), .B1 (nx10146), .C0 (que_out_8__3__4), .C1 (nx10120
           )) ;
    aoi22 ix7710 (.Y (nx7709), .A0 (que_out_25__3__4), .A1 (nx10068), .B0 (
          que_out_16__3__4), .B1 (nx10094)) ;
    aoi22 ix7712 (.Y (nx7711), .A0 (que_out_24__3__4), .A1 (nx10042), .B0 (
          que_out_22__3__4), .B1 (nx10016)) ;
    nand03 ix2385 (.Y (nx2384), .A0 (nx7715), .A1 (nx7717), .A2 (nx7719)) ;
    aoi222 ix7716 (.Y (nx7715), .A0 (que_out_15__3__4), .A1 (nx9964), .B0 (
           que_out_3__3__4), .B1 (nx9990), .C0 (que_out_23__3__4), .C1 (nx9938)
           ) ;
    aoi22 ix7718 (.Y (nx7717), .A0 (que_out_27__3__4), .A1 (nx9912), .B0 (
          que_out_4__3__4), .B1 (nx9886)) ;
    aoi22 ix7720 (.Y (nx7719), .A0 (que_out_0__3__4), .A1 (nx9834), .B0 (
          que_out_2__3__4), .B1 (nx9860)) ;
    nand03 ix2359 (.Y (nx2358), .A0 (nx7723), .A1 (nx7725), .A2 (nx7727)) ;
    aoi222 ix7724 (.Y (nx7723), .A0 (que_out_26__3__4), .A1 (nx9808), .B0 (
           que_out_14__3__4), .B1 (nx9782), .C0 (que_out_11__3__4), .C1 (nx9756)
           ) ;
    aoi22 ix7726 (.Y (nx7725), .A0 (que_out_13__3__4), .A1 (nx9730), .B0 (
          que_out_7__3__4), .B1 (nx9704)) ;
    aoi22 ix7728 (.Y (nx7727), .A0 (que_out_12__3__4), .A1 (nx9678), .B0 (
          que_out_1__3__4), .B1 (nx9652)) ;
    or04 ix2553 (.Y (out_column_3__5), .A0 (nx2548), .A1 (nx2522), .A2 (nx2494)
         , .A3 (nx2468)) ;
    nand03 ix2549 (.Y (nx2548), .A0 (nx7733), .A1 (nx7735), .A2 (nx7737)) ;
    aoi222 ix7734 (.Y (nx7733), .A0 (que_out_10__3__5), .A1 (nx10304), .B0 (
           que_out_6__3__5), .B1 (nx10356), .C0 (que_out_9__3__5), .C1 (nx10330)
           ) ;
    aoi22 ix7736 (.Y (nx7735), .A0 (que_out_5__3__5), .A1 (nx10252), .B0 (
          que_out_18__3__5), .B1 (nx10278)) ;
    aoi22 ix7738 (.Y (nx7737), .A0 (que_out_17__3__5), .A1 (nx10226), .B0 (
          que_out_20__3__5), .B1 (nx10200)) ;
    nand03 ix2523 (.Y (nx2522), .A0 (nx7741), .A1 (nx7743), .A2 (nx7745)) ;
    aoi222 ix7742 (.Y (nx7741), .A0 (que_out_19__3__5), .A1 (nx10174), .B0 (
           que_out_21__3__5), .B1 (nx10148), .C0 (que_out_8__3__5), .C1 (nx10122
           )) ;
    aoi22 ix7744 (.Y (nx7743), .A0 (que_out_25__3__5), .A1 (nx10070), .B0 (
          que_out_16__3__5), .B1 (nx10096)) ;
    aoi22 ix7746 (.Y (nx7745), .A0 (que_out_24__3__5), .A1 (nx10044), .B0 (
          que_out_22__3__5), .B1 (nx10018)) ;
    nand03 ix2495 (.Y (nx2494), .A0 (nx7749), .A1 (nx7751), .A2 (nx7753)) ;
    aoi222 ix7750 (.Y (nx7749), .A0 (que_out_15__3__5), .A1 (nx9966), .B0 (
           que_out_3__3__5), .B1 (nx9992), .C0 (que_out_23__3__5), .C1 (nx9940)
           ) ;
    aoi22 ix7752 (.Y (nx7751), .A0 (que_out_27__3__5), .A1 (nx9914), .B0 (
          que_out_4__3__5), .B1 (nx9888)) ;
    aoi22 ix7754 (.Y (nx7753), .A0 (que_out_0__3__5), .A1 (nx9836), .B0 (
          que_out_2__3__5), .B1 (nx9862)) ;
    nand03 ix2469 (.Y (nx2468), .A0 (nx7757), .A1 (nx7759), .A2 (nx7761)) ;
    aoi222 ix7758 (.Y (nx7757), .A0 (que_out_26__3__5), .A1 (nx9810), .B0 (
           que_out_14__3__5), .B1 (nx9784), .C0 (que_out_11__3__5), .C1 (nx9758)
           ) ;
    aoi22 ix7760 (.Y (nx7759), .A0 (que_out_13__3__5), .A1 (nx9732), .B0 (
          que_out_7__3__5), .B1 (nx9706)) ;
    aoi22 ix7762 (.Y (nx7761), .A0 (que_out_12__3__5), .A1 (nx9680), .B0 (
          que_out_1__3__5), .B1 (nx9654)) ;
    or04 ix2663 (.Y (out_column_3__6), .A0 (nx2658), .A1 (nx2632), .A2 (nx2604)
         , .A3 (nx2578)) ;
    nand03 ix2659 (.Y (nx2658), .A0 (nx7767), .A1 (nx7769), .A2 (nx7771)) ;
    aoi222 ix7768 (.Y (nx7767), .A0 (que_out_10__3__6), .A1 (nx10304), .B0 (
           que_out_6__3__6), .B1 (nx10356), .C0 (que_out_9__3__6), .C1 (nx10330)
           ) ;
    aoi22 ix7770 (.Y (nx7769), .A0 (que_out_5__3__6), .A1 (nx10252), .B0 (
          que_out_18__3__6), .B1 (nx10278)) ;
    aoi22 ix7772 (.Y (nx7771), .A0 (que_out_17__3__6), .A1 (nx10226), .B0 (
          que_out_20__3__6), .B1 (nx10200)) ;
    nand03 ix2633 (.Y (nx2632), .A0 (nx7775), .A1 (nx7777), .A2 (nx7779)) ;
    aoi222 ix7776 (.Y (nx7775), .A0 (que_out_19__3__6), .A1 (nx10174), .B0 (
           que_out_21__3__6), .B1 (nx10148), .C0 (que_out_8__3__6), .C1 (nx10122
           )) ;
    aoi22 ix7778 (.Y (nx7777), .A0 (que_out_25__3__6), .A1 (nx10070), .B0 (
          que_out_16__3__6), .B1 (nx10096)) ;
    aoi22 ix7780 (.Y (nx7779), .A0 (que_out_24__3__6), .A1 (nx10044), .B0 (
          que_out_22__3__6), .B1 (nx10018)) ;
    nand03 ix2605 (.Y (nx2604), .A0 (nx7783), .A1 (nx7785), .A2 (nx7787)) ;
    aoi222 ix7784 (.Y (nx7783), .A0 (que_out_15__3__6), .A1 (nx9966), .B0 (
           que_out_3__3__6), .B1 (nx9992), .C0 (que_out_23__3__6), .C1 (nx9940)
           ) ;
    aoi22 ix7786 (.Y (nx7785), .A0 (que_out_27__3__6), .A1 (nx9914), .B0 (
          que_out_4__3__6), .B1 (nx9888)) ;
    aoi22 ix7788 (.Y (nx7787), .A0 (que_out_0__3__6), .A1 (nx9836), .B0 (
          que_out_2__3__6), .B1 (nx9862)) ;
    nand03 ix2579 (.Y (nx2578), .A0 (nx7791), .A1 (nx7793), .A2 (nx7795)) ;
    aoi222 ix7792 (.Y (nx7791), .A0 (que_out_26__3__6), .A1 (nx9810), .B0 (
           que_out_14__3__6), .B1 (nx9784), .C0 (que_out_11__3__6), .C1 (nx9758)
           ) ;
    aoi22 ix7794 (.Y (nx7793), .A0 (que_out_13__3__6), .A1 (nx9732), .B0 (
          que_out_7__3__6), .B1 (nx9706)) ;
    aoi22 ix7796 (.Y (nx7795), .A0 (que_out_12__3__6), .A1 (nx9680), .B0 (
          que_out_1__3__6), .B1 (nx9654)) ;
    or04 ix2773 (.Y (out_column_3__7), .A0 (nx2768), .A1 (nx2742), .A2 (nx2714)
         , .A3 (nx2688)) ;
    nand03 ix2769 (.Y (nx2768), .A0 (nx7801), .A1 (nx7803), .A2 (nx7805)) ;
    aoi222 ix7802 (.Y (nx7801), .A0 (que_out_10__3__7), .A1 (nx10304), .B0 (
           que_out_6__3__7), .B1 (nx10356), .C0 (que_out_9__3__7), .C1 (nx10330)
           ) ;
    aoi22 ix7804 (.Y (nx7803), .A0 (que_out_5__3__7), .A1 (nx10252), .B0 (
          que_out_18__3__7), .B1 (nx10278)) ;
    aoi22 ix7806 (.Y (nx7805), .A0 (que_out_17__3__7), .A1 (nx10226), .B0 (
          que_out_20__3__7), .B1 (nx10200)) ;
    nand03 ix2743 (.Y (nx2742), .A0 (nx7809), .A1 (nx7811), .A2 (nx7813)) ;
    aoi222 ix7810 (.Y (nx7809), .A0 (que_out_19__3__7), .A1 (nx10174), .B0 (
           que_out_21__3__7), .B1 (nx10148), .C0 (que_out_8__3__7), .C1 (nx10122
           )) ;
    aoi22 ix7812 (.Y (nx7811), .A0 (que_out_25__3__7), .A1 (nx10070), .B0 (
          que_out_16__3__7), .B1 (nx10096)) ;
    aoi22 ix7814 (.Y (nx7813), .A0 (que_out_24__3__7), .A1 (nx10044), .B0 (
          que_out_22__3__7), .B1 (nx10018)) ;
    nand03 ix2715 (.Y (nx2714), .A0 (nx7817), .A1 (nx7819), .A2 (nx7821)) ;
    aoi222 ix7818 (.Y (nx7817), .A0 (que_out_15__3__7), .A1 (nx9966), .B0 (
           que_out_3__3__7), .B1 (nx9992), .C0 (que_out_23__3__7), .C1 (nx9940)
           ) ;
    aoi22 ix7820 (.Y (nx7819), .A0 (que_out_27__3__7), .A1 (nx9914), .B0 (
          que_out_4__3__7), .B1 (nx9888)) ;
    aoi22 ix7822 (.Y (nx7821), .A0 (que_out_0__3__7), .A1 (nx9836), .B0 (
          que_out_2__3__7), .B1 (nx9862)) ;
    nand03 ix2689 (.Y (nx2688), .A0 (nx7825), .A1 (nx7827), .A2 (nx7829)) ;
    aoi222 ix7826 (.Y (nx7825), .A0 (que_out_26__3__7), .A1 (nx9810), .B0 (
           que_out_14__3__7), .B1 (nx9784), .C0 (que_out_11__3__7), .C1 (nx9758)
           ) ;
    aoi22 ix7828 (.Y (nx7827), .A0 (que_out_13__3__7), .A1 (nx9732), .B0 (
          que_out_7__3__7), .B1 (nx9706)) ;
    aoi22 ix7830 (.Y (nx7829), .A0 (que_out_12__3__7), .A1 (nx9680), .B0 (
          que_out_1__3__7), .B1 (nx9654)) ;
    or04 ix2883 (.Y (out_column_3__8), .A0 (nx2878), .A1 (nx2852), .A2 (nx2824)
         , .A3 (nx2798)) ;
    nand03 ix2879 (.Y (nx2878), .A0 (nx7835), .A1 (nx7837), .A2 (nx7839)) ;
    aoi222 ix7836 (.Y (nx7835), .A0 (que_out_10__3__8), .A1 (nx10304), .B0 (
           que_out_6__3__8), .B1 (nx10356), .C0 (que_out_9__3__8), .C1 (nx10330)
           ) ;
    aoi22 ix7838 (.Y (nx7837), .A0 (que_out_5__3__8), .A1 (nx10252), .B0 (
          que_out_18__3__8), .B1 (nx10278)) ;
    aoi22 ix7840 (.Y (nx7839), .A0 (que_out_17__3__8), .A1 (nx10226), .B0 (
          que_out_20__3__8), .B1 (nx10200)) ;
    nand03 ix2853 (.Y (nx2852), .A0 (nx7843), .A1 (nx7845), .A2 (nx7847)) ;
    aoi222 ix7844 (.Y (nx7843), .A0 (que_out_19__3__8), .A1 (nx10174), .B0 (
           que_out_21__3__8), .B1 (nx10148), .C0 (que_out_8__3__8), .C1 (nx10122
           )) ;
    aoi22 ix7846 (.Y (nx7845), .A0 (que_out_25__3__8), .A1 (nx10070), .B0 (
          que_out_16__3__8), .B1 (nx10096)) ;
    aoi22 ix7848 (.Y (nx7847), .A0 (que_out_24__3__8), .A1 (nx10044), .B0 (
          que_out_22__3__8), .B1 (nx10018)) ;
    nand03 ix2825 (.Y (nx2824), .A0 (nx7851), .A1 (nx7853), .A2 (nx7855)) ;
    aoi222 ix7852 (.Y (nx7851), .A0 (que_out_15__3__8), .A1 (nx9966), .B0 (
           que_out_3__3__8), .B1 (nx9992), .C0 (que_out_23__3__8), .C1 (nx9940)
           ) ;
    aoi22 ix7854 (.Y (nx7853), .A0 (que_out_27__3__8), .A1 (nx9914), .B0 (
          que_out_4__3__8), .B1 (nx9888)) ;
    aoi22 ix7856 (.Y (nx7855), .A0 (que_out_0__3__8), .A1 (nx9836), .B0 (
          que_out_2__3__8), .B1 (nx9862)) ;
    nand03 ix2799 (.Y (nx2798), .A0 (nx7859), .A1 (nx7861), .A2 (nx7863)) ;
    aoi222 ix7860 (.Y (nx7859), .A0 (que_out_26__3__8), .A1 (nx9810), .B0 (
           que_out_14__3__8), .B1 (nx9784), .C0 (que_out_11__3__8), .C1 (nx9758)
           ) ;
    aoi22 ix7862 (.Y (nx7861), .A0 (que_out_13__3__8), .A1 (nx9732), .B0 (
          que_out_7__3__8), .B1 (nx9706)) ;
    aoi22 ix7864 (.Y (nx7863), .A0 (que_out_12__3__8), .A1 (nx9680), .B0 (
          que_out_1__3__8), .B1 (nx9654)) ;
    or04 ix2993 (.Y (out_column_3__9), .A0 (nx2988), .A1 (nx2962), .A2 (nx2934)
         , .A3 (nx2908)) ;
    nand03 ix2989 (.Y (nx2988), .A0 (nx7869), .A1 (nx7871), .A2 (nx7873)) ;
    aoi222 ix7870 (.Y (nx7869), .A0 (que_out_10__3__9), .A1 (nx10304), .B0 (
           que_out_6__3__9), .B1 (nx10356), .C0 (que_out_9__3__9), .C1 (nx10330)
           ) ;
    aoi22 ix7872 (.Y (nx7871), .A0 (que_out_5__3__9), .A1 (nx10252), .B0 (
          que_out_18__3__9), .B1 (nx10278)) ;
    aoi22 ix7874 (.Y (nx7873), .A0 (que_out_17__3__9), .A1 (nx10226), .B0 (
          que_out_20__3__9), .B1 (nx10200)) ;
    nand03 ix2963 (.Y (nx2962), .A0 (nx7877), .A1 (nx7879), .A2 (nx7881)) ;
    aoi222 ix7878 (.Y (nx7877), .A0 (que_out_19__3__9), .A1 (nx10174), .B0 (
           que_out_21__3__9), .B1 (nx10148), .C0 (que_out_8__3__9), .C1 (nx10122
           )) ;
    aoi22 ix7880 (.Y (nx7879), .A0 (que_out_25__3__9), .A1 (nx10070), .B0 (
          que_out_16__3__9), .B1 (nx10096)) ;
    aoi22 ix7882 (.Y (nx7881), .A0 (que_out_24__3__9), .A1 (nx10044), .B0 (
          que_out_22__3__9), .B1 (nx10018)) ;
    nand03 ix2935 (.Y (nx2934), .A0 (nx7885), .A1 (nx7887), .A2 (nx7889)) ;
    aoi222 ix7886 (.Y (nx7885), .A0 (que_out_15__3__9), .A1 (nx9966), .B0 (
           que_out_3__3__9), .B1 (nx9992), .C0 (que_out_23__3__9), .C1 (nx9940)
           ) ;
    aoi22 ix7888 (.Y (nx7887), .A0 (que_out_27__3__9), .A1 (nx9914), .B0 (
          que_out_4__3__9), .B1 (nx9888)) ;
    aoi22 ix7890 (.Y (nx7889), .A0 (que_out_0__3__9), .A1 (nx9836), .B0 (
          que_out_2__3__9), .B1 (nx9862)) ;
    nand03 ix2909 (.Y (nx2908), .A0 (nx7893), .A1 (nx7895), .A2 (nx7897)) ;
    aoi222 ix7894 (.Y (nx7893), .A0 (que_out_26__3__9), .A1 (nx9810), .B0 (
           que_out_14__3__9), .B1 (nx9784), .C0 (que_out_11__3__9), .C1 (nx9758)
           ) ;
    aoi22 ix7896 (.Y (nx7895), .A0 (que_out_13__3__9), .A1 (nx9732), .B0 (
          que_out_7__3__9), .B1 (nx9706)) ;
    aoi22 ix7898 (.Y (nx7897), .A0 (que_out_12__3__9), .A1 (nx9680), .B0 (
          que_out_1__3__9), .B1 (nx9654)) ;
    or04 ix3103 (.Y (out_column_3__10), .A0 (nx3098), .A1 (nx3072), .A2 (nx3044)
         , .A3 (nx3018)) ;
    nand03 ix3099 (.Y (nx3098), .A0 (nx7903), .A1 (nx7905), .A2 (nx7907)) ;
    aoi222 ix7904 (.Y (nx7903), .A0 (que_out_10__3__10), .A1 (nx10304), .B0 (
           que_out_6__3__10), .B1 (nx10356), .C0 (que_out_9__3__10), .C1 (
           nx10330)) ;
    aoi22 ix7906 (.Y (nx7905), .A0 (que_out_5__3__10), .A1 (nx10252), .B0 (
          que_out_18__3__10), .B1 (nx10278)) ;
    aoi22 ix7908 (.Y (nx7907), .A0 (que_out_17__3__10), .A1 (nx10226), .B0 (
          que_out_20__3__10), .B1 (nx10200)) ;
    nand03 ix3073 (.Y (nx3072), .A0 (nx7911), .A1 (nx7913), .A2 (nx7915)) ;
    aoi222 ix7912 (.Y (nx7911), .A0 (que_out_19__3__10), .A1 (nx10174), .B0 (
           que_out_21__3__10), .B1 (nx10148), .C0 (que_out_8__3__10), .C1 (
           nx10122)) ;
    aoi22 ix7914 (.Y (nx7913), .A0 (que_out_25__3__10), .A1 (nx10070), .B0 (
          que_out_16__3__10), .B1 (nx10096)) ;
    aoi22 ix7916 (.Y (nx7915), .A0 (que_out_24__3__10), .A1 (nx10044), .B0 (
          que_out_22__3__10), .B1 (nx10018)) ;
    nand03 ix3045 (.Y (nx3044), .A0 (nx7919), .A1 (nx7921), .A2 (nx7923)) ;
    aoi222 ix7920 (.Y (nx7919), .A0 (que_out_15__3__10), .A1 (nx9966), .B0 (
           que_out_3__3__10), .B1 (nx9992), .C0 (que_out_23__3__10), .C1 (nx9940
           )) ;
    aoi22 ix7922 (.Y (nx7921), .A0 (que_out_27__3__10), .A1 (nx9914), .B0 (
          que_out_4__3__10), .B1 (nx9888)) ;
    aoi22 ix7924 (.Y (nx7923), .A0 (que_out_0__3__10), .A1 (nx9836), .B0 (
          que_out_2__3__10), .B1 (nx9862)) ;
    nand03 ix3019 (.Y (nx3018), .A0 (nx7927), .A1 (nx7929), .A2 (nx7931)) ;
    aoi222 ix7928 (.Y (nx7927), .A0 (que_out_26__3__10), .A1 (nx9810), .B0 (
           que_out_14__3__10), .B1 (nx9784), .C0 (que_out_11__3__10), .C1 (
           nx9758)) ;
    aoi22 ix7930 (.Y (nx7929), .A0 (que_out_13__3__10), .A1 (nx9732), .B0 (
          que_out_7__3__10), .B1 (nx9706)) ;
    aoi22 ix7932 (.Y (nx7931), .A0 (que_out_12__3__10), .A1 (nx9680), .B0 (
          que_out_1__3__10), .B1 (nx9654)) ;
    or04 ix3213 (.Y (out_column_3__11), .A0 (nx3208), .A1 (nx3182), .A2 (nx3154)
         , .A3 (nx3128)) ;
    nand03 ix3209 (.Y (nx3208), .A0 (nx7937), .A1 (nx7939), .A2 (nx7941)) ;
    aoi222 ix7938 (.Y (nx7937), .A0 (que_out_10__3__11), .A1 (nx10304), .B0 (
           que_out_6__3__11), .B1 (nx10356), .C0 (que_out_9__3__11), .C1 (
           nx10330)) ;
    aoi22 ix7940 (.Y (nx7939), .A0 (que_out_5__3__11), .A1 (nx10252), .B0 (
          que_out_18__3__11), .B1 (nx10278)) ;
    aoi22 ix7942 (.Y (nx7941), .A0 (que_out_17__3__11), .A1 (nx10226), .B0 (
          que_out_20__3__11), .B1 (nx10200)) ;
    nand03 ix3183 (.Y (nx3182), .A0 (nx7945), .A1 (nx7947), .A2 (nx7949)) ;
    aoi222 ix7946 (.Y (nx7945), .A0 (que_out_19__3__11), .A1 (nx10174), .B0 (
           que_out_21__3__11), .B1 (nx10148), .C0 (que_out_8__3__11), .C1 (
           nx10122)) ;
    aoi22 ix7948 (.Y (nx7947), .A0 (que_out_25__3__11), .A1 (nx10070), .B0 (
          que_out_16__3__11), .B1 (nx10096)) ;
    aoi22 ix7950 (.Y (nx7949), .A0 (que_out_24__3__11), .A1 (nx10044), .B0 (
          que_out_22__3__11), .B1 (nx10018)) ;
    nand03 ix3155 (.Y (nx3154), .A0 (nx7953), .A1 (nx7955), .A2 (nx7957)) ;
    aoi222 ix7954 (.Y (nx7953), .A0 (que_out_15__3__11), .A1 (nx9966), .B0 (
           que_out_3__3__11), .B1 (nx9992), .C0 (que_out_23__3__11), .C1 (nx9940
           )) ;
    aoi22 ix7956 (.Y (nx7955), .A0 (que_out_27__3__11), .A1 (nx9914), .B0 (
          que_out_4__3__11), .B1 (nx9888)) ;
    aoi22 ix7958 (.Y (nx7957), .A0 (que_out_0__3__11), .A1 (nx9836), .B0 (
          que_out_2__3__11), .B1 (nx9862)) ;
    nand03 ix3129 (.Y (nx3128), .A0 (nx7961), .A1 (nx7963), .A2 (nx7965)) ;
    aoi222 ix7962 (.Y (nx7961), .A0 (que_out_26__3__11), .A1 (nx9810), .B0 (
           que_out_14__3__11), .B1 (nx9784), .C0 (que_out_11__3__11), .C1 (
           nx9758)) ;
    aoi22 ix7964 (.Y (nx7963), .A0 (que_out_13__3__11), .A1 (nx9732), .B0 (
          que_out_7__3__11), .B1 (nx9706)) ;
    aoi22 ix7966 (.Y (nx7965), .A0 (que_out_12__3__11), .A1 (nx9680), .B0 (
          que_out_1__3__11), .B1 (nx9654)) ;
    or04 ix3323 (.Y (out_column_3__12), .A0 (nx3318), .A1 (nx3292), .A2 (nx3264)
         , .A3 (nx3238)) ;
    nand03 ix3319 (.Y (nx3318), .A0 (nx7971), .A1 (nx7973), .A2 (nx7975)) ;
    aoi222 ix7972 (.Y (nx7971), .A0 (que_out_10__3__12), .A1 (nx10306), .B0 (
           que_out_6__3__12), .B1 (nx10358), .C0 (que_out_9__3__12), .C1 (
           nx10332)) ;
    aoi22 ix7974 (.Y (nx7973), .A0 (que_out_5__3__12), .A1 (nx10254), .B0 (
          que_out_18__3__12), .B1 (nx10280)) ;
    aoi22 ix7976 (.Y (nx7975), .A0 (que_out_17__3__12), .A1 (nx10228), .B0 (
          que_out_20__3__12), .B1 (nx10202)) ;
    nand03 ix3293 (.Y (nx3292), .A0 (nx7979), .A1 (nx7981), .A2 (nx7983)) ;
    aoi222 ix7980 (.Y (nx7979), .A0 (que_out_19__3__12), .A1 (nx10176), .B0 (
           que_out_21__3__12), .B1 (nx10150), .C0 (que_out_8__3__12), .C1 (
           nx10124)) ;
    aoi22 ix7982 (.Y (nx7981), .A0 (que_out_25__3__12), .A1 (nx10072), .B0 (
          que_out_16__3__12), .B1 (nx10098)) ;
    aoi22 ix7984 (.Y (nx7983), .A0 (que_out_24__3__12), .A1 (nx10046), .B0 (
          que_out_22__3__12), .B1 (nx10020)) ;
    nand03 ix3265 (.Y (nx3264), .A0 (nx7987), .A1 (nx7989), .A2 (nx7991)) ;
    aoi222 ix7988 (.Y (nx7987), .A0 (que_out_15__3__12), .A1 (nx9968), .B0 (
           que_out_3__3__12), .B1 (nx9994), .C0 (que_out_23__3__12), .C1 (nx9942
           )) ;
    aoi22 ix7990 (.Y (nx7989), .A0 (que_out_27__3__12), .A1 (nx9916), .B0 (
          que_out_4__3__12), .B1 (nx9890)) ;
    aoi22 ix7992 (.Y (nx7991), .A0 (que_out_0__3__12), .A1 (nx9838), .B0 (
          que_out_2__3__12), .B1 (nx9864)) ;
    nand03 ix3239 (.Y (nx3238), .A0 (nx7995), .A1 (nx7997), .A2 (nx7999)) ;
    aoi222 ix7996 (.Y (nx7995), .A0 (que_out_26__3__12), .A1 (nx9812), .B0 (
           que_out_14__3__12), .B1 (nx9786), .C0 (que_out_11__3__12), .C1 (
           nx9760)) ;
    aoi22 ix7998 (.Y (nx7997), .A0 (que_out_13__3__12), .A1 (nx9734), .B0 (
          que_out_7__3__12), .B1 (nx9708)) ;
    aoi22 ix8000 (.Y (nx7999), .A0 (que_out_12__3__12), .A1 (nx9682), .B0 (
          que_out_1__3__12), .B1 (nx9656)) ;
    or04 ix3433 (.Y (out_column_3__13), .A0 (nx3428), .A1 (nx3402), .A2 (nx3374)
         , .A3 (nx3348)) ;
    nand03 ix3429 (.Y (nx3428), .A0 (nx8005), .A1 (nx8007), .A2 (nx8009)) ;
    aoi222 ix8006 (.Y (nx8005), .A0 (que_out_10__3__13), .A1 (nx10306), .B0 (
           que_out_6__3__13), .B1 (nx10358), .C0 (que_out_9__3__13), .C1 (
           nx10332)) ;
    aoi22 ix8008 (.Y (nx8007), .A0 (que_out_5__3__13), .A1 (nx10254), .B0 (
          que_out_18__3__13), .B1 (nx10280)) ;
    aoi22 ix8010 (.Y (nx8009), .A0 (que_out_17__3__13), .A1 (nx10228), .B0 (
          que_out_20__3__13), .B1 (nx10202)) ;
    nand03 ix3403 (.Y (nx3402), .A0 (nx8013), .A1 (nx8015), .A2 (nx8017)) ;
    aoi222 ix8014 (.Y (nx8013), .A0 (que_out_19__3__13), .A1 (nx10176), .B0 (
           que_out_21__3__13), .B1 (nx10150), .C0 (que_out_8__3__13), .C1 (
           nx10124)) ;
    aoi22 ix8016 (.Y (nx8015), .A0 (que_out_25__3__13), .A1 (nx10072), .B0 (
          que_out_16__3__13), .B1 (nx10098)) ;
    aoi22 ix8018 (.Y (nx8017), .A0 (que_out_24__3__13), .A1 (nx10046), .B0 (
          que_out_22__3__13), .B1 (nx10020)) ;
    nand03 ix3375 (.Y (nx3374), .A0 (nx8021), .A1 (nx8023), .A2 (nx8025)) ;
    aoi222 ix8022 (.Y (nx8021), .A0 (que_out_15__3__13), .A1 (nx9968), .B0 (
           que_out_3__3__13), .B1 (nx9994), .C0 (que_out_23__3__13), .C1 (nx9942
           )) ;
    aoi22 ix8024 (.Y (nx8023), .A0 (que_out_27__3__13), .A1 (nx9916), .B0 (
          que_out_4__3__13), .B1 (nx9890)) ;
    aoi22 ix8026 (.Y (nx8025), .A0 (que_out_0__3__13), .A1 (nx9838), .B0 (
          que_out_2__3__13), .B1 (nx9864)) ;
    nand03 ix3349 (.Y (nx3348), .A0 (nx8029), .A1 (nx8031), .A2 (nx8033)) ;
    aoi222 ix8030 (.Y (nx8029), .A0 (que_out_26__3__13), .A1 (nx9812), .B0 (
           que_out_14__3__13), .B1 (nx9786), .C0 (que_out_11__3__13), .C1 (
           nx9760)) ;
    aoi22 ix8032 (.Y (nx8031), .A0 (que_out_13__3__13), .A1 (nx9734), .B0 (
          que_out_7__3__13), .B1 (nx9708)) ;
    aoi22 ix8034 (.Y (nx8033), .A0 (que_out_12__3__13), .A1 (nx9682), .B0 (
          que_out_1__3__13), .B1 (nx9656)) ;
    or04 ix3543 (.Y (out_column_3__14), .A0 (nx3538), .A1 (nx3512), .A2 (nx3484)
         , .A3 (nx3458)) ;
    nand03 ix3539 (.Y (nx3538), .A0 (nx8039), .A1 (nx8041), .A2 (nx8043)) ;
    aoi222 ix8040 (.Y (nx8039), .A0 (que_out_10__3__14), .A1 (nx10306), .B0 (
           que_out_6__3__14), .B1 (nx10358), .C0 (que_out_9__3__14), .C1 (
           nx10332)) ;
    aoi22 ix8042 (.Y (nx8041), .A0 (que_out_5__3__14), .A1 (nx10254), .B0 (
          que_out_18__3__14), .B1 (nx10280)) ;
    aoi22 ix8044 (.Y (nx8043), .A0 (que_out_17__3__14), .A1 (nx10228), .B0 (
          que_out_20__3__14), .B1 (nx10202)) ;
    nand03 ix3513 (.Y (nx3512), .A0 (nx8047), .A1 (nx8049), .A2 (nx8051)) ;
    aoi222 ix8048 (.Y (nx8047), .A0 (que_out_19__3__14), .A1 (nx10176), .B0 (
           que_out_21__3__14), .B1 (nx10150), .C0 (que_out_8__3__14), .C1 (
           nx10124)) ;
    aoi22 ix8050 (.Y (nx8049), .A0 (que_out_25__3__14), .A1 (nx10072), .B0 (
          que_out_16__3__14), .B1 (nx10098)) ;
    aoi22 ix8052 (.Y (nx8051), .A0 (que_out_24__3__14), .A1 (nx10046), .B0 (
          que_out_22__3__14), .B1 (nx10020)) ;
    nand03 ix3485 (.Y (nx3484), .A0 (nx8055), .A1 (nx8057), .A2 (nx8059)) ;
    aoi222 ix8056 (.Y (nx8055), .A0 (que_out_15__3__14), .A1 (nx9968), .B0 (
           que_out_3__3__14), .B1 (nx9994), .C0 (que_out_23__3__14), .C1 (nx9942
           )) ;
    aoi22 ix8058 (.Y (nx8057), .A0 (que_out_27__3__14), .A1 (nx9916), .B0 (
          que_out_4__3__14), .B1 (nx9890)) ;
    aoi22 ix8060 (.Y (nx8059), .A0 (que_out_0__3__14), .A1 (nx9838), .B0 (
          que_out_2__3__14), .B1 (nx9864)) ;
    nand03 ix3459 (.Y (nx3458), .A0 (nx8063), .A1 (nx8065), .A2 (nx8067)) ;
    aoi222 ix8064 (.Y (nx8063), .A0 (que_out_26__3__14), .A1 (nx9812), .B0 (
           que_out_14__3__14), .B1 (nx9786), .C0 (que_out_11__3__14), .C1 (
           nx9760)) ;
    aoi22 ix8066 (.Y (nx8065), .A0 (que_out_13__3__14), .A1 (nx9734), .B0 (
          que_out_7__3__14), .B1 (nx9708)) ;
    aoi22 ix8068 (.Y (nx8067), .A0 (que_out_12__3__14), .A1 (nx9682), .B0 (
          que_out_1__3__14), .B1 (nx9656)) ;
    or04 ix3653 (.Y (out_column_3__15), .A0 (nx3648), .A1 (nx3622), .A2 (nx3594)
         , .A3 (nx3568)) ;
    nand03 ix3649 (.Y (nx3648), .A0 (nx8073), .A1 (nx8075), .A2 (nx8077)) ;
    aoi222 ix8074 (.Y (nx8073), .A0 (que_out_10__3__15), .A1 (nx10306), .B0 (
           que_out_6__3__15), .B1 (nx10358), .C0 (que_out_9__3__15), .C1 (
           nx10332)) ;
    aoi22 ix8076 (.Y (nx8075), .A0 (que_out_5__3__15), .A1 (nx10254), .B0 (
          que_out_18__3__15), .B1 (nx10280)) ;
    aoi22 ix8078 (.Y (nx8077), .A0 (que_out_17__3__15), .A1 (nx10228), .B0 (
          que_out_20__3__15), .B1 (nx10202)) ;
    nand03 ix3623 (.Y (nx3622), .A0 (nx8081), .A1 (nx8083), .A2 (nx8085)) ;
    aoi222 ix8082 (.Y (nx8081), .A0 (que_out_19__3__15), .A1 (nx10176), .B0 (
           que_out_21__3__15), .B1 (nx10150), .C0 (que_out_8__3__15), .C1 (
           nx10124)) ;
    aoi22 ix8084 (.Y (nx8083), .A0 (que_out_25__3__15), .A1 (nx10072), .B0 (
          que_out_16__3__15), .B1 (nx10098)) ;
    aoi22 ix8086 (.Y (nx8085), .A0 (que_out_24__3__15), .A1 (nx10046), .B0 (
          que_out_22__3__15), .B1 (nx10020)) ;
    nand03 ix3595 (.Y (nx3594), .A0 (nx8089), .A1 (nx8091), .A2 (nx8093)) ;
    aoi222 ix8090 (.Y (nx8089), .A0 (que_out_15__3__15), .A1 (nx9968), .B0 (
           que_out_3__3__15), .B1 (nx9994), .C0 (que_out_23__3__15), .C1 (nx9942
           )) ;
    aoi22 ix8092 (.Y (nx8091), .A0 (que_out_27__3__15), .A1 (nx9916), .B0 (
          que_out_4__3__15), .B1 (nx9890)) ;
    aoi22 ix8094 (.Y (nx8093), .A0 (que_out_0__3__15), .A1 (nx9838), .B0 (
          que_out_2__3__15), .B1 (nx9864)) ;
    nand03 ix3569 (.Y (nx3568), .A0 (nx8097), .A1 (nx8099), .A2 (nx8101)) ;
    aoi222 ix8098 (.Y (nx8097), .A0 (que_out_26__3__15), .A1 (nx9812), .B0 (
           que_out_14__3__15), .B1 (nx9786), .C0 (que_out_11__3__15), .C1 (
           nx9760)) ;
    aoi22 ix8100 (.Y (nx8099), .A0 (que_out_13__3__15), .A1 (nx9734), .B0 (
          que_out_7__3__15), .B1 (nx9708)) ;
    aoi22 ix8102 (.Y (nx8101), .A0 (que_out_12__3__15), .A1 (nx9682), .B0 (
          que_out_1__3__15), .B1 (nx9656)) ;
    or04 ix3763 (.Y (out_column_2__0), .A0 (nx3758), .A1 (nx3732), .A2 (nx3704)
         , .A3 (nx3678)) ;
    nand03 ix3759 (.Y (nx3758), .A0 (nx8107), .A1 (nx8109), .A2 (nx8111)) ;
    aoi222 ix8108 (.Y (nx8107), .A0 (que_out_10__2__0), .A1 (nx10306), .B0 (
           que_out_6__2__0), .B1 (nx10358), .C0 (que_out_9__2__0), .C1 (nx10332)
           ) ;
    aoi22 ix8110 (.Y (nx8109), .A0 (que_out_5__2__0), .A1 (nx10254), .B0 (
          que_out_18__2__0), .B1 (nx10280)) ;
    aoi22 ix8112 (.Y (nx8111), .A0 (que_out_17__2__0), .A1 (nx10228), .B0 (
          que_out_20__2__0), .B1 (nx10202)) ;
    nand03 ix3733 (.Y (nx3732), .A0 (nx8115), .A1 (nx8117), .A2 (nx8119)) ;
    aoi222 ix8116 (.Y (nx8115), .A0 (que_out_19__2__0), .A1 (nx10176), .B0 (
           que_out_21__2__0), .B1 (nx10150), .C0 (que_out_8__2__0), .C1 (nx10124
           )) ;
    aoi22 ix8118 (.Y (nx8117), .A0 (que_out_25__2__0), .A1 (nx10072), .B0 (
          que_out_16__2__0), .B1 (nx10098)) ;
    aoi22 ix8120 (.Y (nx8119), .A0 (que_out_24__2__0), .A1 (nx10046), .B0 (
          que_out_22__2__0), .B1 (nx10020)) ;
    nand03 ix3705 (.Y (nx3704), .A0 (nx8123), .A1 (nx8125), .A2 (nx8127)) ;
    aoi222 ix8124 (.Y (nx8123), .A0 (que_out_15__2__0), .A1 (nx9968), .B0 (
           que_out_3__2__0), .B1 (nx9994), .C0 (que_out_23__2__0), .C1 (nx9942)
           ) ;
    aoi22 ix8126 (.Y (nx8125), .A0 (que_out_27__2__0), .A1 (nx9916), .B0 (
          que_out_4__2__0), .B1 (nx9890)) ;
    aoi22 ix8128 (.Y (nx8127), .A0 (que_out_0__2__0), .A1 (nx9838), .B0 (
          que_out_2__2__0), .B1 (nx9864)) ;
    nand03 ix3679 (.Y (nx3678), .A0 (nx8131), .A1 (nx8133), .A2 (nx8135)) ;
    aoi222 ix8132 (.Y (nx8131), .A0 (que_out_26__2__0), .A1 (nx9812), .B0 (
           que_out_14__2__0), .B1 (nx9786), .C0 (que_out_11__2__0), .C1 (nx9760)
           ) ;
    aoi22 ix8134 (.Y (nx8133), .A0 (que_out_13__2__0), .A1 (nx9734), .B0 (
          que_out_7__2__0), .B1 (nx9708)) ;
    aoi22 ix8136 (.Y (nx8135), .A0 (que_out_12__2__0), .A1 (nx9682), .B0 (
          que_out_1__2__0), .B1 (nx9656)) ;
    or04 ix3873 (.Y (out_column_2__1), .A0 (nx3868), .A1 (nx3842), .A2 (nx3814)
         , .A3 (nx3788)) ;
    nand03 ix3869 (.Y (nx3868), .A0 (nx8141), .A1 (nx8143), .A2 (nx8145)) ;
    aoi222 ix8142 (.Y (nx8141), .A0 (que_out_10__2__1), .A1 (nx10306), .B0 (
           que_out_6__2__1), .B1 (nx10358), .C0 (que_out_9__2__1), .C1 (nx10332)
           ) ;
    aoi22 ix8144 (.Y (nx8143), .A0 (que_out_5__2__1), .A1 (nx10254), .B0 (
          que_out_18__2__1), .B1 (nx10280)) ;
    aoi22 ix8146 (.Y (nx8145), .A0 (que_out_17__2__1), .A1 (nx10228), .B0 (
          que_out_20__2__1), .B1 (nx10202)) ;
    nand03 ix3843 (.Y (nx3842), .A0 (nx8149), .A1 (nx8151), .A2 (nx8153)) ;
    aoi222 ix8150 (.Y (nx8149), .A0 (que_out_19__2__1), .A1 (nx10176), .B0 (
           que_out_21__2__1), .B1 (nx10150), .C0 (que_out_8__2__1), .C1 (nx10124
           )) ;
    aoi22 ix8152 (.Y (nx8151), .A0 (que_out_25__2__1), .A1 (nx10072), .B0 (
          que_out_16__2__1), .B1 (nx10098)) ;
    aoi22 ix8154 (.Y (nx8153), .A0 (que_out_24__2__1), .A1 (nx10046), .B0 (
          que_out_22__2__1), .B1 (nx10020)) ;
    nand03 ix3815 (.Y (nx3814), .A0 (nx8157), .A1 (nx8159), .A2 (nx8161)) ;
    aoi222 ix8158 (.Y (nx8157), .A0 (que_out_15__2__1), .A1 (nx9968), .B0 (
           que_out_3__2__1), .B1 (nx9994), .C0 (que_out_23__2__1), .C1 (nx9942)
           ) ;
    aoi22 ix8160 (.Y (nx8159), .A0 (que_out_27__2__1), .A1 (nx9916), .B0 (
          que_out_4__2__1), .B1 (nx9890)) ;
    aoi22 ix8162 (.Y (nx8161), .A0 (que_out_0__2__1), .A1 (nx9838), .B0 (
          que_out_2__2__1), .B1 (nx9864)) ;
    nand03 ix3789 (.Y (nx3788), .A0 (nx8165), .A1 (nx8167), .A2 (nx8169)) ;
    aoi222 ix8166 (.Y (nx8165), .A0 (que_out_26__2__1), .A1 (nx9812), .B0 (
           que_out_14__2__1), .B1 (nx9786), .C0 (que_out_11__2__1), .C1 (nx9760)
           ) ;
    aoi22 ix8168 (.Y (nx8167), .A0 (que_out_13__2__1), .A1 (nx9734), .B0 (
          que_out_7__2__1), .B1 (nx9708)) ;
    aoi22 ix8170 (.Y (nx8169), .A0 (que_out_12__2__1), .A1 (nx9682), .B0 (
          que_out_1__2__1), .B1 (nx9656)) ;
    or04 ix3983 (.Y (out_column_2__2), .A0 (nx3978), .A1 (nx3952), .A2 (nx3924)
         , .A3 (nx3898)) ;
    nand03 ix3979 (.Y (nx3978), .A0 (nx8175), .A1 (nx8177), .A2 (nx8179)) ;
    aoi222 ix8176 (.Y (nx8175), .A0 (que_out_10__2__2), .A1 (nx10306), .B0 (
           que_out_6__2__2), .B1 (nx10358), .C0 (que_out_9__2__2), .C1 (nx10332)
           ) ;
    aoi22 ix8178 (.Y (nx8177), .A0 (que_out_5__2__2), .A1 (nx10254), .B0 (
          que_out_18__2__2), .B1 (nx10280)) ;
    aoi22 ix8180 (.Y (nx8179), .A0 (que_out_17__2__2), .A1 (nx10228), .B0 (
          que_out_20__2__2), .B1 (nx10202)) ;
    nand03 ix3953 (.Y (nx3952), .A0 (nx8183), .A1 (nx8185), .A2 (nx8187)) ;
    aoi222 ix8184 (.Y (nx8183), .A0 (que_out_19__2__2), .A1 (nx10176), .B0 (
           que_out_21__2__2), .B1 (nx10150), .C0 (que_out_8__2__2), .C1 (nx10124
           )) ;
    aoi22 ix8186 (.Y (nx8185), .A0 (que_out_25__2__2), .A1 (nx10072), .B0 (
          que_out_16__2__2), .B1 (nx10098)) ;
    aoi22 ix8188 (.Y (nx8187), .A0 (que_out_24__2__2), .A1 (nx10046), .B0 (
          que_out_22__2__2), .B1 (nx10020)) ;
    nand03 ix3925 (.Y (nx3924), .A0 (nx8191), .A1 (nx8193), .A2 (nx8195)) ;
    aoi222 ix8192 (.Y (nx8191), .A0 (que_out_15__2__2), .A1 (nx9968), .B0 (
           que_out_3__2__2), .B1 (nx9994), .C0 (que_out_23__2__2), .C1 (nx9942)
           ) ;
    aoi22 ix8194 (.Y (nx8193), .A0 (que_out_27__2__2), .A1 (nx9916), .B0 (
          que_out_4__2__2), .B1 (nx9890)) ;
    aoi22 ix8196 (.Y (nx8195), .A0 (que_out_0__2__2), .A1 (nx9838), .B0 (
          que_out_2__2__2), .B1 (nx9864)) ;
    nand03 ix3899 (.Y (nx3898), .A0 (nx8199), .A1 (nx8201), .A2 (nx8203)) ;
    aoi222 ix8200 (.Y (nx8199), .A0 (que_out_26__2__2), .A1 (nx9812), .B0 (
           que_out_14__2__2), .B1 (nx9786), .C0 (que_out_11__2__2), .C1 (nx9760)
           ) ;
    aoi22 ix8202 (.Y (nx8201), .A0 (que_out_13__2__2), .A1 (nx9734), .B0 (
          que_out_7__2__2), .B1 (nx9708)) ;
    aoi22 ix8204 (.Y (nx8203), .A0 (que_out_12__2__2), .A1 (nx9682), .B0 (
          que_out_1__2__2), .B1 (nx9656)) ;
    or04 ix4093 (.Y (out_column_2__3), .A0 (nx4088), .A1 (nx4062), .A2 (nx4034)
         , .A3 (nx4008)) ;
    nand03 ix4089 (.Y (nx4088), .A0 (nx8209), .A1 (nx8211), .A2 (nx8213)) ;
    aoi222 ix8210 (.Y (nx8209), .A0 (que_out_10__2__3), .A1 (nx10308), .B0 (
           que_out_6__2__3), .B1 (nx10360), .C0 (que_out_9__2__3), .C1 (nx10334)
           ) ;
    aoi22 ix8212 (.Y (nx8211), .A0 (que_out_5__2__3), .A1 (nx10256), .B0 (
          que_out_18__2__3), .B1 (nx10282)) ;
    aoi22 ix8214 (.Y (nx8213), .A0 (que_out_17__2__3), .A1 (nx10230), .B0 (
          que_out_20__2__3), .B1 (nx10204)) ;
    nand03 ix4063 (.Y (nx4062), .A0 (nx8217), .A1 (nx8219), .A2 (nx8221)) ;
    aoi222 ix8218 (.Y (nx8217), .A0 (que_out_19__2__3), .A1 (nx10178), .B0 (
           que_out_21__2__3), .B1 (nx10152), .C0 (que_out_8__2__3), .C1 (nx10126
           )) ;
    aoi22 ix8220 (.Y (nx8219), .A0 (que_out_25__2__3), .A1 (nx10074), .B0 (
          que_out_16__2__3), .B1 (nx10100)) ;
    aoi22 ix8222 (.Y (nx8221), .A0 (que_out_24__2__3), .A1 (nx10048), .B0 (
          que_out_22__2__3), .B1 (nx10022)) ;
    nand03 ix4035 (.Y (nx4034), .A0 (nx8225), .A1 (nx8227), .A2 (nx8229)) ;
    aoi222 ix8226 (.Y (nx8225), .A0 (que_out_15__2__3), .A1 (nx9970), .B0 (
           que_out_3__2__3), .B1 (nx9996), .C0 (que_out_23__2__3), .C1 (nx9944)
           ) ;
    aoi22 ix8228 (.Y (nx8227), .A0 (que_out_27__2__3), .A1 (nx9918), .B0 (
          que_out_4__2__3), .B1 (nx9892)) ;
    aoi22 ix8230 (.Y (nx8229), .A0 (que_out_0__2__3), .A1 (nx9840), .B0 (
          que_out_2__2__3), .B1 (nx9866)) ;
    nand03 ix4009 (.Y (nx4008), .A0 (nx8233), .A1 (nx8235), .A2 (nx8237)) ;
    aoi222 ix8234 (.Y (nx8233), .A0 (que_out_26__2__3), .A1 (nx9814), .B0 (
           que_out_14__2__3), .B1 (nx9788), .C0 (que_out_11__2__3), .C1 (nx9762)
           ) ;
    aoi22 ix8236 (.Y (nx8235), .A0 (que_out_13__2__3), .A1 (nx9736), .B0 (
          que_out_7__2__3), .B1 (nx9710)) ;
    aoi22 ix8238 (.Y (nx8237), .A0 (que_out_12__2__3), .A1 (nx9684), .B0 (
          que_out_1__2__3), .B1 (nx9658)) ;
    or04 ix4203 (.Y (out_column_2__4), .A0 (nx4198), .A1 (nx4172), .A2 (nx4144)
         , .A3 (nx4118)) ;
    nand03 ix4199 (.Y (nx4198), .A0 (nx8243), .A1 (nx8245), .A2 (nx8247)) ;
    aoi222 ix8244 (.Y (nx8243), .A0 (que_out_10__2__4), .A1 (nx10308), .B0 (
           que_out_6__2__4), .B1 (nx10360), .C0 (que_out_9__2__4), .C1 (nx10334)
           ) ;
    aoi22 ix8246 (.Y (nx8245), .A0 (que_out_5__2__4), .A1 (nx10256), .B0 (
          que_out_18__2__4), .B1 (nx10282)) ;
    aoi22 ix8248 (.Y (nx8247), .A0 (que_out_17__2__4), .A1 (nx10230), .B0 (
          que_out_20__2__4), .B1 (nx10204)) ;
    nand03 ix4173 (.Y (nx4172), .A0 (nx8251), .A1 (nx8253), .A2 (nx8255)) ;
    aoi222 ix8252 (.Y (nx8251), .A0 (que_out_19__2__4), .A1 (nx10178), .B0 (
           que_out_21__2__4), .B1 (nx10152), .C0 (que_out_8__2__4), .C1 (nx10126
           )) ;
    aoi22 ix8254 (.Y (nx8253), .A0 (que_out_25__2__4), .A1 (nx10074), .B0 (
          que_out_16__2__4), .B1 (nx10100)) ;
    aoi22 ix8256 (.Y (nx8255), .A0 (que_out_24__2__4), .A1 (nx10048), .B0 (
          que_out_22__2__4), .B1 (nx10022)) ;
    nand03 ix4145 (.Y (nx4144), .A0 (nx8259), .A1 (nx8261), .A2 (nx8263)) ;
    aoi222 ix8260 (.Y (nx8259), .A0 (que_out_15__2__4), .A1 (nx9970), .B0 (
           que_out_3__2__4), .B1 (nx9996), .C0 (que_out_23__2__4), .C1 (nx9944)
           ) ;
    aoi22 ix8262 (.Y (nx8261), .A0 (que_out_27__2__4), .A1 (nx9918), .B0 (
          que_out_4__2__4), .B1 (nx9892)) ;
    aoi22 ix8264 (.Y (nx8263), .A0 (que_out_0__2__4), .A1 (nx9840), .B0 (
          que_out_2__2__4), .B1 (nx9866)) ;
    nand03 ix4119 (.Y (nx4118), .A0 (nx8267), .A1 (nx8269), .A2 (nx8271)) ;
    aoi222 ix8268 (.Y (nx8267), .A0 (que_out_26__2__4), .A1 (nx9814), .B0 (
           que_out_14__2__4), .B1 (nx9788), .C0 (que_out_11__2__4), .C1 (nx9762)
           ) ;
    aoi22 ix8270 (.Y (nx8269), .A0 (que_out_13__2__4), .A1 (nx9736), .B0 (
          que_out_7__2__4), .B1 (nx9710)) ;
    aoi22 ix8272 (.Y (nx8271), .A0 (que_out_12__2__4), .A1 (nx9684), .B0 (
          que_out_1__2__4), .B1 (nx9658)) ;
    or04 ix4313 (.Y (out_column_2__5), .A0 (nx4308), .A1 (nx4282), .A2 (nx4254)
         , .A3 (nx4228)) ;
    nand03 ix4309 (.Y (nx4308), .A0 (nx8277), .A1 (nx8279), .A2 (nx8281)) ;
    aoi222 ix8278 (.Y (nx8277), .A0 (que_out_10__2__5), .A1 (nx10308), .B0 (
           que_out_6__2__5), .B1 (nx10360), .C0 (que_out_9__2__5), .C1 (nx10334)
           ) ;
    aoi22 ix8280 (.Y (nx8279), .A0 (que_out_5__2__5), .A1 (nx10256), .B0 (
          que_out_18__2__5), .B1 (nx10282)) ;
    aoi22 ix8282 (.Y (nx8281), .A0 (que_out_17__2__5), .A1 (nx10230), .B0 (
          que_out_20__2__5), .B1 (nx10204)) ;
    nand03 ix4283 (.Y (nx4282), .A0 (nx8285), .A1 (nx8287), .A2 (nx8289)) ;
    aoi222 ix8286 (.Y (nx8285), .A0 (que_out_19__2__5), .A1 (nx10178), .B0 (
           que_out_21__2__5), .B1 (nx10152), .C0 (que_out_8__2__5), .C1 (nx10126
           )) ;
    aoi22 ix8288 (.Y (nx8287), .A0 (que_out_25__2__5), .A1 (nx10074), .B0 (
          que_out_16__2__5), .B1 (nx10100)) ;
    aoi22 ix8290 (.Y (nx8289), .A0 (que_out_24__2__5), .A1 (nx10048), .B0 (
          que_out_22__2__5), .B1 (nx10022)) ;
    nand03 ix4255 (.Y (nx4254), .A0 (nx8293), .A1 (nx8295), .A2 (nx8297)) ;
    aoi222 ix8294 (.Y (nx8293), .A0 (que_out_15__2__5), .A1 (nx9970), .B0 (
           que_out_3__2__5), .B1 (nx9996), .C0 (que_out_23__2__5), .C1 (nx9944)
           ) ;
    aoi22 ix8296 (.Y (nx8295), .A0 (que_out_27__2__5), .A1 (nx9918), .B0 (
          que_out_4__2__5), .B1 (nx9892)) ;
    aoi22 ix8298 (.Y (nx8297), .A0 (que_out_0__2__5), .A1 (nx9840), .B0 (
          que_out_2__2__5), .B1 (nx9866)) ;
    nand03 ix4229 (.Y (nx4228), .A0 (nx8301), .A1 (nx8303), .A2 (nx8305)) ;
    aoi222 ix8302 (.Y (nx8301), .A0 (que_out_26__2__5), .A1 (nx9814), .B0 (
           que_out_14__2__5), .B1 (nx9788), .C0 (que_out_11__2__5), .C1 (nx9762)
           ) ;
    aoi22 ix8304 (.Y (nx8303), .A0 (que_out_13__2__5), .A1 (nx9736), .B0 (
          que_out_7__2__5), .B1 (nx9710)) ;
    aoi22 ix8306 (.Y (nx8305), .A0 (que_out_12__2__5), .A1 (nx9684), .B0 (
          que_out_1__2__5), .B1 (nx9658)) ;
    or04 ix4423 (.Y (out_column_2__6), .A0 (nx4418), .A1 (nx4392), .A2 (nx4364)
         , .A3 (nx4338)) ;
    nand03 ix4419 (.Y (nx4418), .A0 (nx8311), .A1 (nx8313), .A2 (nx8315)) ;
    aoi222 ix8312 (.Y (nx8311), .A0 (que_out_10__2__6), .A1 (nx10308), .B0 (
           que_out_6__2__6), .B1 (nx10360), .C0 (que_out_9__2__6), .C1 (nx10334)
           ) ;
    aoi22 ix8314 (.Y (nx8313), .A0 (que_out_5__2__6), .A1 (nx10256), .B0 (
          que_out_18__2__6), .B1 (nx10282)) ;
    aoi22 ix8316 (.Y (nx8315), .A0 (que_out_17__2__6), .A1 (nx10230), .B0 (
          que_out_20__2__6), .B1 (nx10204)) ;
    nand03 ix4393 (.Y (nx4392), .A0 (nx8319), .A1 (nx8321), .A2 (nx8323)) ;
    aoi222 ix8320 (.Y (nx8319), .A0 (que_out_19__2__6), .A1 (nx10178), .B0 (
           que_out_21__2__6), .B1 (nx10152), .C0 (que_out_8__2__6), .C1 (nx10126
           )) ;
    aoi22 ix8322 (.Y (nx8321), .A0 (que_out_25__2__6), .A1 (nx10074), .B0 (
          que_out_16__2__6), .B1 (nx10100)) ;
    aoi22 ix8324 (.Y (nx8323), .A0 (que_out_24__2__6), .A1 (nx10048), .B0 (
          que_out_22__2__6), .B1 (nx10022)) ;
    nand03 ix4365 (.Y (nx4364), .A0 (nx8327), .A1 (nx8329), .A2 (nx8331)) ;
    aoi222 ix8328 (.Y (nx8327), .A0 (que_out_15__2__6), .A1 (nx9970), .B0 (
           que_out_3__2__6), .B1 (nx9996), .C0 (que_out_23__2__6), .C1 (nx9944)
           ) ;
    aoi22 ix8330 (.Y (nx8329), .A0 (que_out_27__2__6), .A1 (nx9918), .B0 (
          que_out_4__2__6), .B1 (nx9892)) ;
    aoi22 ix8332 (.Y (nx8331), .A0 (que_out_0__2__6), .A1 (nx9840), .B0 (
          que_out_2__2__6), .B1 (nx9866)) ;
    nand03 ix4339 (.Y (nx4338), .A0 (nx8335), .A1 (nx8337), .A2 (nx8339)) ;
    aoi222 ix8336 (.Y (nx8335), .A0 (que_out_26__2__6), .A1 (nx9814), .B0 (
           que_out_14__2__6), .B1 (nx9788), .C0 (que_out_11__2__6), .C1 (nx9762)
           ) ;
    aoi22 ix8338 (.Y (nx8337), .A0 (que_out_13__2__6), .A1 (nx9736), .B0 (
          que_out_7__2__6), .B1 (nx9710)) ;
    aoi22 ix8340 (.Y (nx8339), .A0 (que_out_12__2__6), .A1 (nx9684), .B0 (
          que_out_1__2__6), .B1 (nx9658)) ;
    or04 ix4533 (.Y (out_column_2__7), .A0 (nx4528), .A1 (nx4502), .A2 (nx4474)
         , .A3 (nx4448)) ;
    nand03 ix4529 (.Y (nx4528), .A0 (nx8345), .A1 (nx8347), .A2 (nx8349)) ;
    aoi222 ix8346 (.Y (nx8345), .A0 (que_out_10__2__7), .A1 (nx10308), .B0 (
           que_out_6__2__7), .B1 (nx10360), .C0 (que_out_9__2__7), .C1 (nx10334)
           ) ;
    aoi22 ix8348 (.Y (nx8347), .A0 (que_out_5__2__7), .A1 (nx10256), .B0 (
          que_out_18__2__7), .B1 (nx10282)) ;
    aoi22 ix8350 (.Y (nx8349), .A0 (que_out_17__2__7), .A1 (nx10230), .B0 (
          que_out_20__2__7), .B1 (nx10204)) ;
    nand03 ix4503 (.Y (nx4502), .A0 (nx8353), .A1 (nx8355), .A2 (nx8357)) ;
    aoi222 ix8354 (.Y (nx8353), .A0 (que_out_19__2__7), .A1 (nx10178), .B0 (
           que_out_21__2__7), .B1 (nx10152), .C0 (que_out_8__2__7), .C1 (nx10126
           )) ;
    aoi22 ix8356 (.Y (nx8355), .A0 (que_out_25__2__7), .A1 (nx10074), .B0 (
          que_out_16__2__7), .B1 (nx10100)) ;
    aoi22 ix8358 (.Y (nx8357), .A0 (que_out_24__2__7), .A1 (nx10048), .B0 (
          que_out_22__2__7), .B1 (nx10022)) ;
    nand03 ix4475 (.Y (nx4474), .A0 (nx8361), .A1 (nx8363), .A2 (nx8365)) ;
    aoi222 ix8362 (.Y (nx8361), .A0 (que_out_15__2__7), .A1 (nx9970), .B0 (
           que_out_3__2__7), .B1 (nx9996), .C0 (que_out_23__2__7), .C1 (nx9944)
           ) ;
    aoi22 ix8364 (.Y (nx8363), .A0 (que_out_27__2__7), .A1 (nx9918), .B0 (
          que_out_4__2__7), .B1 (nx9892)) ;
    aoi22 ix8366 (.Y (nx8365), .A0 (que_out_0__2__7), .A1 (nx9840), .B0 (
          que_out_2__2__7), .B1 (nx9866)) ;
    nand03 ix4449 (.Y (nx4448), .A0 (nx8369), .A1 (nx8371), .A2 (nx8373)) ;
    aoi222 ix8370 (.Y (nx8369), .A0 (que_out_26__2__7), .A1 (nx9814), .B0 (
           que_out_14__2__7), .B1 (nx9788), .C0 (que_out_11__2__7), .C1 (nx9762)
           ) ;
    aoi22 ix8372 (.Y (nx8371), .A0 (que_out_13__2__7), .A1 (nx9736), .B0 (
          que_out_7__2__7), .B1 (nx9710)) ;
    aoi22 ix8374 (.Y (nx8373), .A0 (que_out_12__2__7), .A1 (nx9684), .B0 (
          que_out_1__2__7), .B1 (nx9658)) ;
    or04 ix4643 (.Y (out_column_2__8), .A0 (nx4638), .A1 (nx4612), .A2 (nx4584)
         , .A3 (nx4558)) ;
    nand03 ix4639 (.Y (nx4638), .A0 (nx8379), .A1 (nx8381), .A2 (nx8383)) ;
    aoi222 ix8380 (.Y (nx8379), .A0 (que_out_10__2__8), .A1 (nx10308), .B0 (
           que_out_6__2__8), .B1 (nx10360), .C0 (que_out_9__2__8), .C1 (nx10334)
           ) ;
    aoi22 ix8382 (.Y (nx8381), .A0 (que_out_5__2__8), .A1 (nx10256), .B0 (
          que_out_18__2__8), .B1 (nx10282)) ;
    aoi22 ix8384 (.Y (nx8383), .A0 (que_out_17__2__8), .A1 (nx10230), .B0 (
          que_out_20__2__8), .B1 (nx10204)) ;
    nand03 ix4613 (.Y (nx4612), .A0 (nx8387), .A1 (nx8389), .A2 (nx8391)) ;
    aoi222 ix8388 (.Y (nx8387), .A0 (que_out_19__2__8), .A1 (nx10178), .B0 (
           que_out_21__2__8), .B1 (nx10152), .C0 (que_out_8__2__8), .C1 (nx10126
           )) ;
    aoi22 ix8390 (.Y (nx8389), .A0 (que_out_25__2__8), .A1 (nx10074), .B0 (
          que_out_16__2__8), .B1 (nx10100)) ;
    aoi22 ix8392 (.Y (nx8391), .A0 (que_out_24__2__8), .A1 (nx10048), .B0 (
          que_out_22__2__8), .B1 (nx10022)) ;
    nand03 ix4585 (.Y (nx4584), .A0 (nx8395), .A1 (nx8397), .A2 (nx8399)) ;
    aoi222 ix8396 (.Y (nx8395), .A0 (que_out_15__2__8), .A1 (nx9970), .B0 (
           que_out_3__2__8), .B1 (nx9996), .C0 (que_out_23__2__8), .C1 (nx9944)
           ) ;
    aoi22 ix8398 (.Y (nx8397), .A0 (que_out_27__2__8), .A1 (nx9918), .B0 (
          que_out_4__2__8), .B1 (nx9892)) ;
    aoi22 ix8400 (.Y (nx8399), .A0 (que_out_0__2__8), .A1 (nx9840), .B0 (
          que_out_2__2__8), .B1 (nx9866)) ;
    nand03 ix4559 (.Y (nx4558), .A0 (nx8403), .A1 (nx8405), .A2 (nx8407)) ;
    aoi222 ix8404 (.Y (nx8403), .A0 (que_out_26__2__8), .A1 (nx9814), .B0 (
           que_out_14__2__8), .B1 (nx9788), .C0 (que_out_11__2__8), .C1 (nx9762)
           ) ;
    aoi22 ix8406 (.Y (nx8405), .A0 (que_out_13__2__8), .A1 (nx9736), .B0 (
          que_out_7__2__8), .B1 (nx9710)) ;
    aoi22 ix8408 (.Y (nx8407), .A0 (que_out_12__2__8), .A1 (nx9684), .B0 (
          que_out_1__2__8), .B1 (nx9658)) ;
    or04 ix4753 (.Y (out_column_2__9), .A0 (nx4748), .A1 (nx4722), .A2 (nx4694)
         , .A3 (nx4668)) ;
    nand03 ix4749 (.Y (nx4748), .A0 (nx8413), .A1 (nx8415), .A2 (nx8417)) ;
    aoi222 ix8414 (.Y (nx8413), .A0 (que_out_10__2__9), .A1 (nx10308), .B0 (
           que_out_6__2__9), .B1 (nx10360), .C0 (que_out_9__2__9), .C1 (nx10334)
           ) ;
    aoi22 ix8416 (.Y (nx8415), .A0 (que_out_5__2__9), .A1 (nx10256), .B0 (
          que_out_18__2__9), .B1 (nx10282)) ;
    aoi22 ix8418 (.Y (nx8417), .A0 (que_out_17__2__9), .A1 (nx10230), .B0 (
          que_out_20__2__9), .B1 (nx10204)) ;
    nand03 ix4723 (.Y (nx4722), .A0 (nx8421), .A1 (nx8423), .A2 (nx8425)) ;
    aoi222 ix8422 (.Y (nx8421), .A0 (que_out_19__2__9), .A1 (nx10178), .B0 (
           que_out_21__2__9), .B1 (nx10152), .C0 (que_out_8__2__9), .C1 (nx10126
           )) ;
    aoi22 ix8424 (.Y (nx8423), .A0 (que_out_25__2__9), .A1 (nx10074), .B0 (
          que_out_16__2__9), .B1 (nx10100)) ;
    aoi22 ix8426 (.Y (nx8425), .A0 (que_out_24__2__9), .A1 (nx10048), .B0 (
          que_out_22__2__9), .B1 (nx10022)) ;
    nand03 ix4695 (.Y (nx4694), .A0 (nx8429), .A1 (nx8431), .A2 (nx8433)) ;
    aoi222 ix8430 (.Y (nx8429), .A0 (que_out_15__2__9), .A1 (nx9970), .B0 (
           que_out_3__2__9), .B1 (nx9996), .C0 (que_out_23__2__9), .C1 (nx9944)
           ) ;
    aoi22 ix8432 (.Y (nx8431), .A0 (que_out_27__2__9), .A1 (nx9918), .B0 (
          que_out_4__2__9), .B1 (nx9892)) ;
    aoi22 ix8434 (.Y (nx8433), .A0 (que_out_0__2__9), .A1 (nx9840), .B0 (
          que_out_2__2__9), .B1 (nx9866)) ;
    nand03 ix4669 (.Y (nx4668), .A0 (nx8437), .A1 (nx8439), .A2 (nx8441)) ;
    aoi222 ix8438 (.Y (nx8437), .A0 (que_out_26__2__9), .A1 (nx9814), .B0 (
           que_out_14__2__9), .B1 (nx9788), .C0 (que_out_11__2__9), .C1 (nx9762)
           ) ;
    aoi22 ix8440 (.Y (nx8439), .A0 (que_out_13__2__9), .A1 (nx9736), .B0 (
          que_out_7__2__9), .B1 (nx9710)) ;
    aoi22 ix8442 (.Y (nx8441), .A0 (que_out_12__2__9), .A1 (nx9684), .B0 (
          que_out_1__2__9), .B1 (nx9658)) ;
    or04 ix4863 (.Y (out_column_2__10), .A0 (nx4858), .A1 (nx4832), .A2 (nx4804)
         , .A3 (nx4778)) ;
    nand03 ix4859 (.Y (nx4858), .A0 (nx8447), .A1 (nx8449), .A2 (nx8451)) ;
    aoi222 ix8448 (.Y (nx8447), .A0 (que_out_10__2__10), .A1 (nx10310), .B0 (
           que_out_6__2__10), .B1 (nx10362), .C0 (que_out_9__2__10), .C1 (
           nx10336)) ;
    aoi22 ix8450 (.Y (nx8449), .A0 (que_out_5__2__10), .A1 (nx10258), .B0 (
          que_out_18__2__10), .B1 (nx10284)) ;
    aoi22 ix8452 (.Y (nx8451), .A0 (que_out_17__2__10), .A1 (nx10232), .B0 (
          que_out_20__2__10), .B1 (nx10206)) ;
    nand03 ix4833 (.Y (nx4832), .A0 (nx8455), .A1 (nx8457), .A2 (nx8459)) ;
    aoi222 ix8456 (.Y (nx8455), .A0 (que_out_19__2__10), .A1 (nx10180), .B0 (
           que_out_21__2__10), .B1 (nx10154), .C0 (que_out_8__2__10), .C1 (
           nx10128)) ;
    aoi22 ix8458 (.Y (nx8457), .A0 (que_out_25__2__10), .A1 (nx10076), .B0 (
          que_out_16__2__10), .B1 (nx10102)) ;
    aoi22 ix8460 (.Y (nx8459), .A0 (que_out_24__2__10), .A1 (nx10050), .B0 (
          que_out_22__2__10), .B1 (nx10024)) ;
    nand03 ix4805 (.Y (nx4804), .A0 (nx8463), .A1 (nx8465), .A2 (nx8467)) ;
    aoi222 ix8464 (.Y (nx8463), .A0 (que_out_15__2__10), .A1 (nx9972), .B0 (
           que_out_3__2__10), .B1 (nx9998), .C0 (que_out_23__2__10), .C1 (nx9946
           )) ;
    aoi22 ix8466 (.Y (nx8465), .A0 (que_out_27__2__10), .A1 (nx9920), .B0 (
          que_out_4__2__10), .B1 (nx9894)) ;
    aoi22 ix8468 (.Y (nx8467), .A0 (que_out_0__2__10), .A1 (nx9842), .B0 (
          que_out_2__2__10), .B1 (nx9868)) ;
    nand03 ix4779 (.Y (nx4778), .A0 (nx8471), .A1 (nx8473), .A2 (nx8475)) ;
    aoi222 ix8472 (.Y (nx8471), .A0 (que_out_26__2__10), .A1 (nx9816), .B0 (
           que_out_14__2__10), .B1 (nx9790), .C0 (que_out_11__2__10), .C1 (
           nx9764)) ;
    aoi22 ix8474 (.Y (nx8473), .A0 (que_out_13__2__10), .A1 (nx9738), .B0 (
          que_out_7__2__10), .B1 (nx9712)) ;
    aoi22 ix8476 (.Y (nx8475), .A0 (que_out_12__2__10), .A1 (nx9686), .B0 (
          que_out_1__2__10), .B1 (nx9660)) ;
    or04 ix4973 (.Y (out_column_2__11), .A0 (nx4968), .A1 (nx4942), .A2 (nx4914)
         , .A3 (nx4888)) ;
    nand03 ix4969 (.Y (nx4968), .A0 (nx8481), .A1 (nx8483), .A2 (nx8485)) ;
    aoi222 ix8482 (.Y (nx8481), .A0 (que_out_10__2__11), .A1 (nx10310), .B0 (
           que_out_6__2__11), .B1 (nx10362), .C0 (que_out_9__2__11), .C1 (
           nx10336)) ;
    aoi22 ix8484 (.Y (nx8483), .A0 (que_out_5__2__11), .A1 (nx10258), .B0 (
          que_out_18__2__11), .B1 (nx10284)) ;
    aoi22 ix8486 (.Y (nx8485), .A0 (que_out_17__2__11), .A1 (nx10232), .B0 (
          que_out_20__2__11), .B1 (nx10206)) ;
    nand03 ix4943 (.Y (nx4942), .A0 (nx8489), .A1 (nx8491), .A2 (nx8493)) ;
    aoi222 ix8490 (.Y (nx8489), .A0 (que_out_19__2__11), .A1 (nx10180), .B0 (
           que_out_21__2__11), .B1 (nx10154), .C0 (que_out_8__2__11), .C1 (
           nx10128)) ;
    aoi22 ix8492 (.Y (nx8491), .A0 (que_out_25__2__11), .A1 (nx10076), .B0 (
          que_out_16__2__11), .B1 (nx10102)) ;
    aoi22 ix8494 (.Y (nx8493), .A0 (que_out_24__2__11), .A1 (nx10050), .B0 (
          que_out_22__2__11), .B1 (nx10024)) ;
    nand03 ix4915 (.Y (nx4914), .A0 (nx8497), .A1 (nx8499), .A2 (nx8501)) ;
    aoi222 ix8498 (.Y (nx8497), .A0 (que_out_15__2__11), .A1 (nx9972), .B0 (
           que_out_3__2__11), .B1 (nx9998), .C0 (que_out_23__2__11), .C1 (nx9946
           )) ;
    aoi22 ix8500 (.Y (nx8499), .A0 (que_out_27__2__11), .A1 (nx9920), .B0 (
          que_out_4__2__11), .B1 (nx9894)) ;
    aoi22 ix8502 (.Y (nx8501), .A0 (que_out_0__2__11), .A1 (nx9842), .B0 (
          que_out_2__2__11), .B1 (nx9868)) ;
    nand03 ix4889 (.Y (nx4888), .A0 (nx8505), .A1 (nx8507), .A2 (nx8509)) ;
    aoi222 ix8506 (.Y (nx8505), .A0 (que_out_26__2__11), .A1 (nx9816), .B0 (
           que_out_14__2__11), .B1 (nx9790), .C0 (que_out_11__2__11), .C1 (
           nx9764)) ;
    aoi22 ix8508 (.Y (nx8507), .A0 (que_out_13__2__11), .A1 (nx9738), .B0 (
          que_out_7__2__11), .B1 (nx9712)) ;
    aoi22 ix8510 (.Y (nx8509), .A0 (que_out_12__2__11), .A1 (nx9686), .B0 (
          que_out_1__2__11), .B1 (nx9660)) ;
    or04 ix5083 (.Y (out_column_2__12), .A0 (nx5078), .A1 (nx5052), .A2 (nx5024)
         , .A3 (nx4998)) ;
    nand03 ix5079 (.Y (nx5078), .A0 (nx8515), .A1 (nx8517), .A2 (nx8519)) ;
    aoi222 ix8516 (.Y (nx8515), .A0 (que_out_10__2__12), .A1 (nx10310), .B0 (
           que_out_6__2__12), .B1 (nx10362), .C0 (que_out_9__2__12), .C1 (
           nx10336)) ;
    aoi22 ix8518 (.Y (nx8517), .A0 (que_out_5__2__12), .A1 (nx10258), .B0 (
          que_out_18__2__12), .B1 (nx10284)) ;
    aoi22 ix8520 (.Y (nx8519), .A0 (que_out_17__2__12), .A1 (nx10232), .B0 (
          que_out_20__2__12), .B1 (nx10206)) ;
    nand03 ix5053 (.Y (nx5052), .A0 (nx8523), .A1 (nx8525), .A2 (nx8527)) ;
    aoi222 ix8524 (.Y (nx8523), .A0 (que_out_19__2__12), .A1 (nx10180), .B0 (
           que_out_21__2__12), .B1 (nx10154), .C0 (que_out_8__2__12), .C1 (
           nx10128)) ;
    aoi22 ix8526 (.Y (nx8525), .A0 (que_out_25__2__12), .A1 (nx10076), .B0 (
          que_out_16__2__12), .B1 (nx10102)) ;
    aoi22 ix8528 (.Y (nx8527), .A0 (que_out_24__2__12), .A1 (nx10050), .B0 (
          que_out_22__2__12), .B1 (nx10024)) ;
    nand03 ix5025 (.Y (nx5024), .A0 (nx8531), .A1 (nx8533), .A2 (nx8535)) ;
    aoi222 ix8532 (.Y (nx8531), .A0 (que_out_15__2__12), .A1 (nx9972), .B0 (
           que_out_3__2__12), .B1 (nx9998), .C0 (que_out_23__2__12), .C1 (nx9946
           )) ;
    aoi22 ix8534 (.Y (nx8533), .A0 (que_out_27__2__12), .A1 (nx9920), .B0 (
          que_out_4__2__12), .B1 (nx9894)) ;
    aoi22 ix8536 (.Y (nx8535), .A0 (que_out_0__2__12), .A1 (nx9842), .B0 (
          que_out_2__2__12), .B1 (nx9868)) ;
    nand03 ix4999 (.Y (nx4998), .A0 (nx8539), .A1 (nx8541), .A2 (nx8543)) ;
    aoi222 ix8540 (.Y (nx8539), .A0 (que_out_26__2__12), .A1 (nx9816), .B0 (
           que_out_14__2__12), .B1 (nx9790), .C0 (que_out_11__2__12), .C1 (
           nx9764)) ;
    aoi22 ix8542 (.Y (nx8541), .A0 (que_out_13__2__12), .A1 (nx9738), .B0 (
          que_out_7__2__12), .B1 (nx9712)) ;
    aoi22 ix8544 (.Y (nx8543), .A0 (que_out_12__2__12), .A1 (nx9686), .B0 (
          que_out_1__2__12), .B1 (nx9660)) ;
    or04 ix5193 (.Y (out_column_2__13), .A0 (nx5188), .A1 (nx5162), .A2 (nx5134)
         , .A3 (nx5108)) ;
    nand03 ix5189 (.Y (nx5188), .A0 (nx8549), .A1 (nx8551), .A2 (nx8553)) ;
    aoi222 ix8550 (.Y (nx8549), .A0 (que_out_10__2__13), .A1 (nx10310), .B0 (
           que_out_6__2__13), .B1 (nx10362), .C0 (que_out_9__2__13), .C1 (
           nx10336)) ;
    aoi22 ix8552 (.Y (nx8551), .A0 (que_out_5__2__13), .A1 (nx10258), .B0 (
          que_out_18__2__13), .B1 (nx10284)) ;
    aoi22 ix8554 (.Y (nx8553), .A0 (que_out_17__2__13), .A1 (nx10232), .B0 (
          que_out_20__2__13), .B1 (nx10206)) ;
    nand03 ix5163 (.Y (nx5162), .A0 (nx8557), .A1 (nx8559), .A2 (nx8561)) ;
    aoi222 ix8558 (.Y (nx8557), .A0 (que_out_19__2__13), .A1 (nx10180), .B0 (
           que_out_21__2__13), .B1 (nx10154), .C0 (que_out_8__2__13), .C1 (
           nx10128)) ;
    aoi22 ix8560 (.Y (nx8559), .A0 (que_out_25__2__13), .A1 (nx10076), .B0 (
          que_out_16__2__13), .B1 (nx10102)) ;
    aoi22 ix8562 (.Y (nx8561), .A0 (que_out_24__2__13), .A1 (nx10050), .B0 (
          que_out_22__2__13), .B1 (nx10024)) ;
    nand03 ix5135 (.Y (nx5134), .A0 (nx8565), .A1 (nx8567), .A2 (nx8569)) ;
    aoi222 ix8566 (.Y (nx8565), .A0 (que_out_15__2__13), .A1 (nx9972), .B0 (
           que_out_3__2__13), .B1 (nx9998), .C0 (que_out_23__2__13), .C1 (nx9946
           )) ;
    aoi22 ix8568 (.Y (nx8567), .A0 (que_out_27__2__13), .A1 (nx9920), .B0 (
          que_out_4__2__13), .B1 (nx9894)) ;
    aoi22 ix8570 (.Y (nx8569), .A0 (que_out_0__2__13), .A1 (nx9842), .B0 (
          que_out_2__2__13), .B1 (nx9868)) ;
    nand03 ix5109 (.Y (nx5108), .A0 (nx8573), .A1 (nx8575), .A2 (nx8577)) ;
    aoi222 ix8574 (.Y (nx8573), .A0 (que_out_26__2__13), .A1 (nx9816), .B0 (
           que_out_14__2__13), .B1 (nx9790), .C0 (que_out_11__2__13), .C1 (
           nx9764)) ;
    aoi22 ix8576 (.Y (nx8575), .A0 (que_out_13__2__13), .A1 (nx9738), .B0 (
          que_out_7__2__13), .B1 (nx9712)) ;
    aoi22 ix8578 (.Y (nx8577), .A0 (que_out_12__2__13), .A1 (nx9686), .B0 (
          que_out_1__2__13), .B1 (nx9660)) ;
    or04 ix5303 (.Y (out_column_2__14), .A0 (nx5298), .A1 (nx5272), .A2 (nx5244)
         , .A3 (nx5218)) ;
    nand03 ix5299 (.Y (nx5298), .A0 (nx8583), .A1 (nx8585), .A2 (nx8587)) ;
    aoi222 ix8584 (.Y (nx8583), .A0 (que_out_10__2__14), .A1 (nx10310), .B0 (
           que_out_6__2__14), .B1 (nx10362), .C0 (que_out_9__2__14), .C1 (
           nx10336)) ;
    aoi22 ix8586 (.Y (nx8585), .A0 (que_out_5__2__14), .A1 (nx10258), .B0 (
          que_out_18__2__14), .B1 (nx10284)) ;
    aoi22 ix8588 (.Y (nx8587), .A0 (que_out_17__2__14), .A1 (nx10232), .B0 (
          que_out_20__2__14), .B1 (nx10206)) ;
    nand03 ix5273 (.Y (nx5272), .A0 (nx8591), .A1 (nx8593), .A2 (nx8595)) ;
    aoi222 ix8592 (.Y (nx8591), .A0 (que_out_19__2__14), .A1 (nx10180), .B0 (
           que_out_21__2__14), .B1 (nx10154), .C0 (que_out_8__2__14), .C1 (
           nx10128)) ;
    aoi22 ix8594 (.Y (nx8593), .A0 (que_out_25__2__14), .A1 (nx10076), .B0 (
          que_out_16__2__14), .B1 (nx10102)) ;
    aoi22 ix8596 (.Y (nx8595), .A0 (que_out_24__2__14), .A1 (nx10050), .B0 (
          que_out_22__2__14), .B1 (nx10024)) ;
    nand03 ix5245 (.Y (nx5244), .A0 (nx8599), .A1 (nx8601), .A2 (nx8603)) ;
    aoi222 ix8600 (.Y (nx8599), .A0 (que_out_15__2__14), .A1 (nx9972), .B0 (
           que_out_3__2__14), .B1 (nx9998), .C0 (que_out_23__2__14), .C1 (nx9946
           )) ;
    aoi22 ix8602 (.Y (nx8601), .A0 (que_out_27__2__14), .A1 (nx9920), .B0 (
          que_out_4__2__14), .B1 (nx9894)) ;
    aoi22 ix8604 (.Y (nx8603), .A0 (que_out_0__2__14), .A1 (nx9842), .B0 (
          que_out_2__2__14), .B1 (nx9868)) ;
    nand03 ix5219 (.Y (nx5218), .A0 (nx8607), .A1 (nx8609), .A2 (nx8611)) ;
    aoi222 ix8608 (.Y (nx8607), .A0 (que_out_26__2__14), .A1 (nx9816), .B0 (
           que_out_14__2__14), .B1 (nx9790), .C0 (que_out_11__2__14), .C1 (
           nx9764)) ;
    aoi22 ix8610 (.Y (nx8609), .A0 (que_out_13__2__14), .A1 (nx9738), .B0 (
          que_out_7__2__14), .B1 (nx9712)) ;
    aoi22 ix8612 (.Y (nx8611), .A0 (que_out_12__2__14), .A1 (nx9686), .B0 (
          que_out_1__2__14), .B1 (nx9660)) ;
    or04 ix5413 (.Y (out_column_2__15), .A0 (nx5408), .A1 (nx5382), .A2 (nx5354)
         , .A3 (nx5328)) ;
    nand03 ix5409 (.Y (nx5408), .A0 (nx8617), .A1 (nx8619), .A2 (nx8621)) ;
    aoi222 ix8618 (.Y (nx8617), .A0 (que_out_10__2__15), .A1 (nx10310), .B0 (
           que_out_6__2__15), .B1 (nx10362), .C0 (que_out_9__2__15), .C1 (
           nx10336)) ;
    aoi22 ix8620 (.Y (nx8619), .A0 (que_out_5__2__15), .A1 (nx10258), .B0 (
          que_out_18__2__15), .B1 (nx10284)) ;
    aoi22 ix8622 (.Y (nx8621), .A0 (que_out_17__2__15), .A1 (nx10232), .B0 (
          que_out_20__2__15), .B1 (nx10206)) ;
    nand03 ix5383 (.Y (nx5382), .A0 (nx8625), .A1 (nx8627), .A2 (nx8629)) ;
    aoi222 ix8626 (.Y (nx8625), .A0 (que_out_19__2__15), .A1 (nx10180), .B0 (
           que_out_21__2__15), .B1 (nx10154), .C0 (que_out_8__2__15), .C1 (
           nx10128)) ;
    aoi22 ix8628 (.Y (nx8627), .A0 (que_out_25__2__15), .A1 (nx10076), .B0 (
          que_out_16__2__15), .B1 (nx10102)) ;
    aoi22 ix8630 (.Y (nx8629), .A0 (que_out_24__2__15), .A1 (nx10050), .B0 (
          que_out_22__2__15), .B1 (nx10024)) ;
    nand03 ix5355 (.Y (nx5354), .A0 (nx8633), .A1 (nx8635), .A2 (nx8637)) ;
    aoi222 ix8634 (.Y (nx8633), .A0 (que_out_15__2__15), .A1 (nx9972), .B0 (
           que_out_3__2__15), .B1 (nx9998), .C0 (que_out_23__2__15), .C1 (nx9946
           )) ;
    aoi22 ix8636 (.Y (nx8635), .A0 (que_out_27__2__15), .A1 (nx9920), .B0 (
          que_out_4__2__15), .B1 (nx9894)) ;
    aoi22 ix8638 (.Y (nx8637), .A0 (que_out_0__2__15), .A1 (nx9842), .B0 (
          que_out_2__2__15), .B1 (nx9868)) ;
    nand03 ix5329 (.Y (nx5328), .A0 (nx8641), .A1 (nx8643), .A2 (nx8645)) ;
    aoi222 ix8642 (.Y (nx8641), .A0 (que_out_26__2__15), .A1 (nx9816), .B0 (
           que_out_14__2__15), .B1 (nx9790), .C0 (que_out_11__2__15), .C1 (
           nx9764)) ;
    aoi22 ix8644 (.Y (nx8643), .A0 (que_out_13__2__15), .A1 (nx9738), .B0 (
          que_out_7__2__15), .B1 (nx9712)) ;
    aoi22 ix8646 (.Y (nx8645), .A0 (que_out_12__2__15), .A1 (nx9686), .B0 (
          que_out_1__2__15), .B1 (nx9660)) ;
    or04 ix5523 (.Y (out_column_1__0), .A0 (nx5518), .A1 (nx5492), .A2 (nx5464)
         , .A3 (nx5438)) ;
    nand03 ix5519 (.Y (nx5518), .A0 (nx8651), .A1 (nx8653), .A2 (nx8655)) ;
    aoi222 ix8652 (.Y (nx8651), .A0 (que_out_10__1__0), .A1 (nx10310), .B0 (
           que_out_6__1__0), .B1 (nx10362), .C0 (que_out_9__1__0), .C1 (nx10336)
           ) ;
    aoi22 ix8654 (.Y (nx8653), .A0 (que_out_5__1__0), .A1 (nx10258), .B0 (
          que_out_18__1__0), .B1 (nx10284)) ;
    aoi22 ix8656 (.Y (nx8655), .A0 (que_out_17__1__0), .A1 (nx10232), .B0 (
          que_out_20__1__0), .B1 (nx10206)) ;
    nand03 ix5493 (.Y (nx5492), .A0 (nx8659), .A1 (nx8661), .A2 (nx8663)) ;
    aoi222 ix8660 (.Y (nx8659), .A0 (que_out_19__1__0), .A1 (nx10180), .B0 (
           que_out_21__1__0), .B1 (nx10154), .C0 (que_out_8__1__0), .C1 (nx10128
           )) ;
    aoi22 ix8662 (.Y (nx8661), .A0 (que_out_25__1__0), .A1 (nx10076), .B0 (
          que_out_16__1__0), .B1 (nx10102)) ;
    aoi22 ix8664 (.Y (nx8663), .A0 (que_out_24__1__0), .A1 (nx10050), .B0 (
          que_out_22__1__0), .B1 (nx10024)) ;
    nand03 ix5465 (.Y (nx5464), .A0 (nx8667), .A1 (nx8669), .A2 (nx8671)) ;
    aoi222 ix8668 (.Y (nx8667), .A0 (que_out_15__1__0), .A1 (nx9972), .B0 (
           que_out_3__1__0), .B1 (nx9998), .C0 (que_out_23__1__0), .C1 (nx9946)
           ) ;
    aoi22 ix8670 (.Y (nx8669), .A0 (que_out_27__1__0), .A1 (nx9920), .B0 (
          que_out_4__1__0), .B1 (nx9894)) ;
    aoi22 ix8672 (.Y (nx8671), .A0 (que_out_0__1__0), .A1 (nx9842), .B0 (
          que_out_2__1__0), .B1 (nx9868)) ;
    nand03 ix5439 (.Y (nx5438), .A0 (nx8675), .A1 (nx8677), .A2 (nx8679)) ;
    aoi222 ix8676 (.Y (nx8675), .A0 (que_out_26__1__0), .A1 (nx9816), .B0 (
           que_out_14__1__0), .B1 (nx9790), .C0 (que_out_11__1__0), .C1 (nx9764)
           ) ;
    aoi22 ix8678 (.Y (nx8677), .A0 (que_out_13__1__0), .A1 (nx9738), .B0 (
          que_out_7__1__0), .B1 (nx9712)) ;
    aoi22 ix8680 (.Y (nx8679), .A0 (que_out_12__1__0), .A1 (nx9686), .B0 (
          que_out_1__1__0), .B1 (nx9660)) ;
    or04 ix5633 (.Y (out_column_1__1), .A0 (nx5628), .A1 (nx5602), .A2 (nx5574)
         , .A3 (nx5548)) ;
    nand03 ix5629 (.Y (nx5628), .A0 (nx8685), .A1 (nx8687), .A2 (nx8689)) ;
    aoi222 ix8686 (.Y (nx8685), .A0 (que_out_10__1__1), .A1 (nx10312), .B0 (
           que_out_6__1__1), .B1 (nx10364), .C0 (que_out_9__1__1), .C1 (nx10338)
           ) ;
    aoi22 ix8688 (.Y (nx8687), .A0 (que_out_5__1__1), .A1 (nx10260), .B0 (
          que_out_18__1__1), .B1 (nx10286)) ;
    aoi22 ix8690 (.Y (nx8689), .A0 (que_out_17__1__1), .A1 (nx10234), .B0 (
          que_out_20__1__1), .B1 (nx10208)) ;
    nand03 ix5603 (.Y (nx5602), .A0 (nx8693), .A1 (nx8695), .A2 (nx8697)) ;
    aoi222 ix8694 (.Y (nx8693), .A0 (que_out_19__1__1), .A1 (nx10182), .B0 (
           que_out_21__1__1), .B1 (nx10156), .C0 (que_out_8__1__1), .C1 (nx10130
           )) ;
    aoi22 ix8696 (.Y (nx8695), .A0 (que_out_25__1__1), .A1 (nx10078), .B0 (
          que_out_16__1__1), .B1 (nx10104)) ;
    aoi22 ix8698 (.Y (nx8697), .A0 (que_out_24__1__1), .A1 (nx10052), .B0 (
          que_out_22__1__1), .B1 (nx10026)) ;
    nand03 ix5575 (.Y (nx5574), .A0 (nx8701), .A1 (nx8703), .A2 (nx8705)) ;
    aoi222 ix8702 (.Y (nx8701), .A0 (que_out_15__1__1), .A1 (nx9974), .B0 (
           que_out_3__1__1), .B1 (nx10000), .C0 (que_out_23__1__1), .C1 (nx9948)
           ) ;
    aoi22 ix8704 (.Y (nx8703), .A0 (que_out_27__1__1), .A1 (nx9922), .B0 (
          que_out_4__1__1), .B1 (nx9896)) ;
    aoi22 ix8706 (.Y (nx8705), .A0 (que_out_0__1__1), .A1 (nx9844), .B0 (
          que_out_2__1__1), .B1 (nx9870)) ;
    nand03 ix5549 (.Y (nx5548), .A0 (nx8709), .A1 (nx8711), .A2 (nx8713)) ;
    aoi222 ix8710 (.Y (nx8709), .A0 (que_out_26__1__1), .A1 (nx9818), .B0 (
           que_out_14__1__1), .B1 (nx9792), .C0 (que_out_11__1__1), .C1 (nx9766)
           ) ;
    aoi22 ix8712 (.Y (nx8711), .A0 (que_out_13__1__1), .A1 (nx9740), .B0 (
          que_out_7__1__1), .B1 (nx9714)) ;
    aoi22 ix8714 (.Y (nx8713), .A0 (que_out_12__1__1), .A1 (nx9688), .B0 (
          que_out_1__1__1), .B1 (nx9662)) ;
    or04 ix5743 (.Y (out_column_1__2), .A0 (nx5738), .A1 (nx5712), .A2 (nx5684)
         , .A3 (nx5658)) ;
    nand03 ix5739 (.Y (nx5738), .A0 (nx8719), .A1 (nx8721), .A2 (nx8723)) ;
    aoi222 ix8720 (.Y (nx8719), .A0 (que_out_10__1__2), .A1 (nx10312), .B0 (
           que_out_6__1__2), .B1 (nx10364), .C0 (que_out_9__1__2), .C1 (nx10338)
           ) ;
    aoi22 ix8722 (.Y (nx8721), .A0 (que_out_5__1__2), .A1 (nx10260), .B0 (
          que_out_18__1__2), .B1 (nx10286)) ;
    aoi22 ix8724 (.Y (nx8723), .A0 (que_out_17__1__2), .A1 (nx10234), .B0 (
          que_out_20__1__2), .B1 (nx10208)) ;
    nand03 ix5713 (.Y (nx5712), .A0 (nx8727), .A1 (nx8729), .A2 (nx8731)) ;
    aoi222 ix8728 (.Y (nx8727), .A0 (que_out_19__1__2), .A1 (nx10182), .B0 (
           que_out_21__1__2), .B1 (nx10156), .C0 (que_out_8__1__2), .C1 (nx10130
           )) ;
    aoi22 ix8730 (.Y (nx8729), .A0 (que_out_25__1__2), .A1 (nx10078), .B0 (
          que_out_16__1__2), .B1 (nx10104)) ;
    aoi22 ix8732 (.Y (nx8731), .A0 (que_out_24__1__2), .A1 (nx10052), .B0 (
          que_out_22__1__2), .B1 (nx10026)) ;
    nand03 ix5685 (.Y (nx5684), .A0 (nx8735), .A1 (nx8737), .A2 (nx8739)) ;
    aoi222 ix8736 (.Y (nx8735), .A0 (que_out_15__1__2), .A1 (nx9974), .B0 (
           que_out_3__1__2), .B1 (nx10000), .C0 (que_out_23__1__2), .C1 (nx9948)
           ) ;
    aoi22 ix8738 (.Y (nx8737), .A0 (que_out_27__1__2), .A1 (nx9922), .B0 (
          que_out_4__1__2), .B1 (nx9896)) ;
    aoi22 ix8740 (.Y (nx8739), .A0 (que_out_0__1__2), .A1 (nx9844), .B0 (
          que_out_2__1__2), .B1 (nx9870)) ;
    nand03 ix5659 (.Y (nx5658), .A0 (nx8743), .A1 (nx8745), .A2 (nx8747)) ;
    aoi222 ix8744 (.Y (nx8743), .A0 (que_out_26__1__2), .A1 (nx9818), .B0 (
           que_out_14__1__2), .B1 (nx9792), .C0 (que_out_11__1__2), .C1 (nx9766)
           ) ;
    aoi22 ix8746 (.Y (nx8745), .A0 (que_out_13__1__2), .A1 (nx9740), .B0 (
          que_out_7__1__2), .B1 (nx9714)) ;
    aoi22 ix8748 (.Y (nx8747), .A0 (que_out_12__1__2), .A1 (nx9688), .B0 (
          que_out_1__1__2), .B1 (nx9662)) ;
    or04 ix5853 (.Y (out_column_1__3), .A0 (nx5848), .A1 (nx5822), .A2 (nx5794)
         , .A3 (nx5768)) ;
    nand03 ix5849 (.Y (nx5848), .A0 (nx8753), .A1 (nx8755), .A2 (nx8757)) ;
    aoi222 ix8754 (.Y (nx8753), .A0 (que_out_10__1__3), .A1 (nx10312), .B0 (
           que_out_6__1__3), .B1 (nx10364), .C0 (que_out_9__1__3), .C1 (nx10338)
           ) ;
    aoi22 ix8756 (.Y (nx8755), .A0 (que_out_5__1__3), .A1 (nx10260), .B0 (
          que_out_18__1__3), .B1 (nx10286)) ;
    aoi22 ix8758 (.Y (nx8757), .A0 (que_out_17__1__3), .A1 (nx10234), .B0 (
          que_out_20__1__3), .B1 (nx10208)) ;
    nand03 ix5823 (.Y (nx5822), .A0 (nx8761), .A1 (nx8763), .A2 (nx8765)) ;
    aoi222 ix8762 (.Y (nx8761), .A0 (que_out_19__1__3), .A1 (nx10182), .B0 (
           que_out_21__1__3), .B1 (nx10156), .C0 (que_out_8__1__3), .C1 (nx10130
           )) ;
    aoi22 ix8764 (.Y (nx8763), .A0 (que_out_25__1__3), .A1 (nx10078), .B0 (
          que_out_16__1__3), .B1 (nx10104)) ;
    aoi22 ix8766 (.Y (nx8765), .A0 (que_out_24__1__3), .A1 (nx10052), .B0 (
          que_out_22__1__3), .B1 (nx10026)) ;
    nand03 ix5795 (.Y (nx5794), .A0 (nx8769), .A1 (nx8771), .A2 (nx8773)) ;
    aoi222 ix8770 (.Y (nx8769), .A0 (que_out_15__1__3), .A1 (nx9974), .B0 (
           que_out_3__1__3), .B1 (nx10000), .C0 (que_out_23__1__3), .C1 (nx9948)
           ) ;
    aoi22 ix8772 (.Y (nx8771), .A0 (que_out_27__1__3), .A1 (nx9922), .B0 (
          que_out_4__1__3), .B1 (nx9896)) ;
    aoi22 ix8774 (.Y (nx8773), .A0 (que_out_0__1__3), .A1 (nx9844), .B0 (
          que_out_2__1__3), .B1 (nx9870)) ;
    nand03 ix5769 (.Y (nx5768), .A0 (nx8777), .A1 (nx8779), .A2 (nx8781)) ;
    aoi222 ix8778 (.Y (nx8777), .A0 (que_out_26__1__3), .A1 (nx9818), .B0 (
           que_out_14__1__3), .B1 (nx9792), .C0 (que_out_11__1__3), .C1 (nx9766)
           ) ;
    aoi22 ix8780 (.Y (nx8779), .A0 (que_out_13__1__3), .A1 (nx9740), .B0 (
          que_out_7__1__3), .B1 (nx9714)) ;
    aoi22 ix8782 (.Y (nx8781), .A0 (que_out_12__1__3), .A1 (nx9688), .B0 (
          que_out_1__1__3), .B1 (nx9662)) ;
    or04 ix5963 (.Y (out_column_1__4), .A0 (nx5958), .A1 (nx5932), .A2 (nx5904)
         , .A3 (nx5878)) ;
    nand03 ix5959 (.Y (nx5958), .A0 (nx8787), .A1 (nx8789), .A2 (nx8791)) ;
    aoi222 ix8788 (.Y (nx8787), .A0 (que_out_10__1__4), .A1 (nx10312), .B0 (
           que_out_6__1__4), .B1 (nx10364), .C0 (que_out_9__1__4), .C1 (nx10338)
           ) ;
    aoi22 ix8790 (.Y (nx8789), .A0 (que_out_5__1__4), .A1 (nx10260), .B0 (
          que_out_18__1__4), .B1 (nx10286)) ;
    aoi22 ix8792 (.Y (nx8791), .A0 (que_out_17__1__4), .A1 (nx10234), .B0 (
          que_out_20__1__4), .B1 (nx10208)) ;
    nand03 ix5933 (.Y (nx5932), .A0 (nx8795), .A1 (nx8797), .A2 (nx8799)) ;
    aoi222 ix8796 (.Y (nx8795), .A0 (que_out_19__1__4), .A1 (nx10182), .B0 (
           que_out_21__1__4), .B1 (nx10156), .C0 (que_out_8__1__4), .C1 (nx10130
           )) ;
    aoi22 ix8798 (.Y (nx8797), .A0 (que_out_25__1__4), .A1 (nx10078), .B0 (
          que_out_16__1__4), .B1 (nx10104)) ;
    aoi22 ix8800 (.Y (nx8799), .A0 (que_out_24__1__4), .A1 (nx10052), .B0 (
          que_out_22__1__4), .B1 (nx10026)) ;
    nand03 ix5905 (.Y (nx5904), .A0 (nx8803), .A1 (nx8805), .A2 (nx8807)) ;
    aoi222 ix8804 (.Y (nx8803), .A0 (que_out_15__1__4), .A1 (nx9974), .B0 (
           que_out_3__1__4), .B1 (nx10000), .C0 (que_out_23__1__4), .C1 (nx9948)
           ) ;
    aoi22 ix8806 (.Y (nx8805), .A0 (que_out_27__1__4), .A1 (nx9922), .B0 (
          que_out_4__1__4), .B1 (nx9896)) ;
    aoi22 ix8808 (.Y (nx8807), .A0 (que_out_0__1__4), .A1 (nx9844), .B0 (
          que_out_2__1__4), .B1 (nx9870)) ;
    nand03 ix5879 (.Y (nx5878), .A0 (nx8811), .A1 (nx8813), .A2 (nx8815)) ;
    aoi222 ix8812 (.Y (nx8811), .A0 (que_out_26__1__4), .A1 (nx9818), .B0 (
           que_out_14__1__4), .B1 (nx9792), .C0 (que_out_11__1__4), .C1 (nx9766)
           ) ;
    aoi22 ix8814 (.Y (nx8813), .A0 (que_out_13__1__4), .A1 (nx9740), .B0 (
          que_out_7__1__4), .B1 (nx9714)) ;
    aoi22 ix8816 (.Y (nx8815), .A0 (que_out_12__1__4), .A1 (nx9688), .B0 (
          que_out_1__1__4), .B1 (nx9662)) ;
    or04 ix6073 (.Y (out_column_1__5), .A0 (nx6068), .A1 (nx6042), .A2 (nx6014)
         , .A3 (nx5988)) ;
    nand03 ix6069 (.Y (nx6068), .A0 (nx8821), .A1 (nx8823), .A2 (nx8825)) ;
    aoi222 ix8822 (.Y (nx8821), .A0 (que_out_10__1__5), .A1 (nx10312), .B0 (
           que_out_6__1__5), .B1 (nx10364), .C0 (que_out_9__1__5), .C1 (nx10338)
           ) ;
    aoi22 ix8824 (.Y (nx8823), .A0 (que_out_5__1__5), .A1 (nx10260), .B0 (
          que_out_18__1__5), .B1 (nx10286)) ;
    aoi22 ix8826 (.Y (nx8825), .A0 (que_out_17__1__5), .A1 (nx10234), .B0 (
          que_out_20__1__5), .B1 (nx10208)) ;
    nand03 ix6043 (.Y (nx6042), .A0 (nx8829), .A1 (nx8831), .A2 (nx8833)) ;
    aoi222 ix8830 (.Y (nx8829), .A0 (que_out_19__1__5), .A1 (nx10182), .B0 (
           que_out_21__1__5), .B1 (nx10156), .C0 (que_out_8__1__5), .C1 (nx10130
           )) ;
    aoi22 ix8832 (.Y (nx8831), .A0 (que_out_25__1__5), .A1 (nx10078), .B0 (
          que_out_16__1__5), .B1 (nx10104)) ;
    aoi22 ix8834 (.Y (nx8833), .A0 (que_out_24__1__5), .A1 (nx10052), .B0 (
          que_out_22__1__5), .B1 (nx10026)) ;
    nand03 ix6015 (.Y (nx6014), .A0 (nx8837), .A1 (nx8839), .A2 (nx8841)) ;
    aoi222 ix8838 (.Y (nx8837), .A0 (que_out_15__1__5), .A1 (nx9974), .B0 (
           que_out_3__1__5), .B1 (nx10000), .C0 (que_out_23__1__5), .C1 (nx9948)
           ) ;
    aoi22 ix8840 (.Y (nx8839), .A0 (que_out_27__1__5), .A1 (nx9922), .B0 (
          que_out_4__1__5), .B1 (nx9896)) ;
    aoi22 ix8842 (.Y (nx8841), .A0 (que_out_0__1__5), .A1 (nx9844), .B0 (
          que_out_2__1__5), .B1 (nx9870)) ;
    nand03 ix5989 (.Y (nx5988), .A0 (nx8845), .A1 (nx8847), .A2 (nx8849)) ;
    aoi222 ix8846 (.Y (nx8845), .A0 (que_out_26__1__5), .A1 (nx9818), .B0 (
           que_out_14__1__5), .B1 (nx9792), .C0 (que_out_11__1__5), .C1 (nx9766)
           ) ;
    aoi22 ix8848 (.Y (nx8847), .A0 (que_out_13__1__5), .A1 (nx9740), .B0 (
          que_out_7__1__5), .B1 (nx9714)) ;
    aoi22 ix8850 (.Y (nx8849), .A0 (que_out_12__1__5), .A1 (nx9688), .B0 (
          que_out_1__1__5), .B1 (nx9662)) ;
    or04 ix6183 (.Y (out_column_1__6), .A0 (nx6178), .A1 (nx6152), .A2 (nx6124)
         , .A3 (nx6098)) ;
    nand03 ix6179 (.Y (nx6178), .A0 (nx8855), .A1 (nx8857), .A2 (nx8859)) ;
    aoi222 ix8856 (.Y (nx8855), .A0 (que_out_10__1__6), .A1 (nx10312), .B0 (
           que_out_6__1__6), .B1 (nx10364), .C0 (que_out_9__1__6), .C1 (nx10338)
           ) ;
    aoi22 ix8858 (.Y (nx8857), .A0 (que_out_5__1__6), .A1 (nx10260), .B0 (
          que_out_18__1__6), .B1 (nx10286)) ;
    aoi22 ix8860 (.Y (nx8859), .A0 (que_out_17__1__6), .A1 (nx10234), .B0 (
          que_out_20__1__6), .B1 (nx10208)) ;
    nand03 ix6153 (.Y (nx6152), .A0 (nx8863), .A1 (nx8865), .A2 (nx8867)) ;
    aoi222 ix8864 (.Y (nx8863), .A0 (que_out_19__1__6), .A1 (nx10182), .B0 (
           que_out_21__1__6), .B1 (nx10156), .C0 (que_out_8__1__6), .C1 (nx10130
           )) ;
    aoi22 ix8866 (.Y (nx8865), .A0 (que_out_25__1__6), .A1 (nx10078), .B0 (
          que_out_16__1__6), .B1 (nx10104)) ;
    aoi22 ix8868 (.Y (nx8867), .A0 (que_out_24__1__6), .A1 (nx10052), .B0 (
          que_out_22__1__6), .B1 (nx10026)) ;
    nand03 ix6125 (.Y (nx6124), .A0 (nx8871), .A1 (nx8873), .A2 (nx8875)) ;
    aoi222 ix8872 (.Y (nx8871), .A0 (que_out_15__1__6), .A1 (nx9974), .B0 (
           que_out_3__1__6), .B1 (nx10000), .C0 (que_out_23__1__6), .C1 (nx9948)
           ) ;
    aoi22 ix8874 (.Y (nx8873), .A0 (que_out_27__1__6), .A1 (nx9922), .B0 (
          que_out_4__1__6), .B1 (nx9896)) ;
    aoi22 ix8876 (.Y (nx8875), .A0 (que_out_0__1__6), .A1 (nx9844), .B0 (
          que_out_2__1__6), .B1 (nx9870)) ;
    nand03 ix6099 (.Y (nx6098), .A0 (nx8879), .A1 (nx8881), .A2 (nx8883)) ;
    aoi222 ix8880 (.Y (nx8879), .A0 (que_out_26__1__6), .A1 (nx9818), .B0 (
           que_out_14__1__6), .B1 (nx9792), .C0 (que_out_11__1__6), .C1 (nx9766)
           ) ;
    aoi22 ix8882 (.Y (nx8881), .A0 (que_out_13__1__6), .A1 (nx9740), .B0 (
          que_out_7__1__6), .B1 (nx9714)) ;
    aoi22 ix8884 (.Y (nx8883), .A0 (que_out_12__1__6), .A1 (nx9688), .B0 (
          que_out_1__1__6), .B1 (nx9662)) ;
    or04 ix6293 (.Y (out_column_1__7), .A0 (nx6288), .A1 (nx6262), .A2 (nx6234)
         , .A3 (nx6208)) ;
    nand03 ix6289 (.Y (nx6288), .A0 (nx8889), .A1 (nx8891), .A2 (nx8893)) ;
    aoi222 ix8890 (.Y (nx8889), .A0 (que_out_10__1__7), .A1 (nx10312), .B0 (
           que_out_6__1__7), .B1 (nx10364), .C0 (que_out_9__1__7), .C1 (nx10338)
           ) ;
    aoi22 ix8892 (.Y (nx8891), .A0 (que_out_5__1__7), .A1 (nx10260), .B0 (
          que_out_18__1__7), .B1 (nx10286)) ;
    aoi22 ix8894 (.Y (nx8893), .A0 (que_out_17__1__7), .A1 (nx10234), .B0 (
          que_out_20__1__7), .B1 (nx10208)) ;
    nand03 ix6263 (.Y (nx6262), .A0 (nx8897), .A1 (nx8899), .A2 (nx8901)) ;
    aoi222 ix8898 (.Y (nx8897), .A0 (que_out_19__1__7), .A1 (nx10182), .B0 (
           que_out_21__1__7), .B1 (nx10156), .C0 (que_out_8__1__7), .C1 (nx10130
           )) ;
    aoi22 ix8900 (.Y (nx8899), .A0 (que_out_25__1__7), .A1 (nx10078), .B0 (
          que_out_16__1__7), .B1 (nx10104)) ;
    aoi22 ix8902 (.Y (nx8901), .A0 (que_out_24__1__7), .A1 (nx10052), .B0 (
          que_out_22__1__7), .B1 (nx10026)) ;
    nand03 ix6235 (.Y (nx6234), .A0 (nx8905), .A1 (nx8907), .A2 (nx8909)) ;
    aoi222 ix8906 (.Y (nx8905), .A0 (que_out_15__1__7), .A1 (nx9974), .B0 (
           que_out_3__1__7), .B1 (nx10000), .C0 (que_out_23__1__7), .C1 (nx9948)
           ) ;
    aoi22 ix8908 (.Y (nx8907), .A0 (que_out_27__1__7), .A1 (nx9922), .B0 (
          que_out_4__1__7), .B1 (nx9896)) ;
    aoi22 ix8910 (.Y (nx8909), .A0 (que_out_0__1__7), .A1 (nx9844), .B0 (
          que_out_2__1__7), .B1 (nx9870)) ;
    nand03 ix6209 (.Y (nx6208), .A0 (nx8913), .A1 (nx8915), .A2 (nx8917)) ;
    aoi222 ix8914 (.Y (nx8913), .A0 (que_out_26__1__7), .A1 (nx9818), .B0 (
           que_out_14__1__7), .B1 (nx9792), .C0 (que_out_11__1__7), .C1 (nx9766)
           ) ;
    aoi22 ix8916 (.Y (nx8915), .A0 (que_out_13__1__7), .A1 (nx9740), .B0 (
          que_out_7__1__7), .B1 (nx9714)) ;
    aoi22 ix8918 (.Y (nx8917), .A0 (que_out_12__1__7), .A1 (nx9688), .B0 (
          que_out_1__1__7), .B1 (nx9662)) ;
    or04 ix6403 (.Y (out_column_1__8), .A0 (nx6398), .A1 (nx6372), .A2 (nx6344)
         , .A3 (nx6318)) ;
    nand03 ix6399 (.Y (nx6398), .A0 (nx8923), .A1 (nx8925), .A2 (nx8927)) ;
    aoi222 ix8924 (.Y (nx8923), .A0 (que_out_10__1__8), .A1 (nx10314), .B0 (
           que_out_6__1__8), .B1 (nx10366), .C0 (que_out_9__1__8), .C1 (nx10340)
           ) ;
    aoi22 ix8926 (.Y (nx8925), .A0 (que_out_5__1__8), .A1 (nx10262), .B0 (
          que_out_18__1__8), .B1 (nx10288)) ;
    aoi22 ix8928 (.Y (nx8927), .A0 (que_out_17__1__8), .A1 (nx10236), .B0 (
          que_out_20__1__8), .B1 (nx10210)) ;
    nand03 ix6373 (.Y (nx6372), .A0 (nx8931), .A1 (nx8933), .A2 (nx8935)) ;
    aoi222 ix8932 (.Y (nx8931), .A0 (que_out_19__1__8), .A1 (nx10184), .B0 (
           que_out_21__1__8), .B1 (nx10158), .C0 (que_out_8__1__8), .C1 (nx10132
           )) ;
    aoi22 ix8934 (.Y (nx8933), .A0 (que_out_25__1__8), .A1 (nx10080), .B0 (
          que_out_16__1__8), .B1 (nx10106)) ;
    aoi22 ix8936 (.Y (nx8935), .A0 (que_out_24__1__8), .A1 (nx10054), .B0 (
          que_out_22__1__8), .B1 (nx10028)) ;
    nand03 ix6345 (.Y (nx6344), .A0 (nx8939), .A1 (nx8941), .A2 (nx8943)) ;
    aoi222 ix8940 (.Y (nx8939), .A0 (que_out_15__1__8), .A1 (nx9976), .B0 (
           que_out_3__1__8), .B1 (nx10002), .C0 (que_out_23__1__8), .C1 (nx9950)
           ) ;
    aoi22 ix8942 (.Y (nx8941), .A0 (que_out_27__1__8), .A1 (nx9924), .B0 (
          que_out_4__1__8), .B1 (nx9898)) ;
    aoi22 ix8944 (.Y (nx8943), .A0 (que_out_0__1__8), .A1 (nx9846), .B0 (
          que_out_2__1__8), .B1 (nx9872)) ;
    nand03 ix6319 (.Y (nx6318), .A0 (nx8947), .A1 (nx8949), .A2 (nx8951)) ;
    aoi222 ix8948 (.Y (nx8947), .A0 (que_out_26__1__8), .A1 (nx9820), .B0 (
           que_out_14__1__8), .B1 (nx9794), .C0 (que_out_11__1__8), .C1 (nx9768)
           ) ;
    aoi22 ix8950 (.Y (nx8949), .A0 (que_out_13__1__8), .A1 (nx9742), .B0 (
          que_out_7__1__8), .B1 (nx9716)) ;
    aoi22 ix8952 (.Y (nx8951), .A0 (que_out_12__1__8), .A1 (nx9690), .B0 (
          que_out_1__1__8), .B1 (nx9664)) ;
    or04 ix6513 (.Y (out_column_1__9), .A0 (nx6508), .A1 (nx6482), .A2 (nx6454)
         , .A3 (nx6428)) ;
    nand03 ix6509 (.Y (nx6508), .A0 (nx8955), .A1 (nx8957), .A2 (nx8959)) ;
    aoi222 ix8956 (.Y (nx8955), .A0 (que_out_10__1__9), .A1 (nx10314), .B0 (
           que_out_6__1__9), .B1 (nx10366), .C0 (que_out_9__1__9), .C1 (nx10340)
           ) ;
    aoi22 ix8958 (.Y (nx8957), .A0 (que_out_5__1__9), .A1 (nx10262), .B0 (
          que_out_18__1__9), .B1 (nx10288)) ;
    aoi22 ix8960 (.Y (nx8959), .A0 (que_out_17__1__9), .A1 (nx10236), .B0 (
          que_out_20__1__9), .B1 (nx10210)) ;
    nand03 ix6483 (.Y (nx6482), .A0 (nx8963), .A1 (nx8965), .A2 (nx8967)) ;
    aoi222 ix8964 (.Y (nx8963), .A0 (que_out_19__1__9), .A1 (nx10184), .B0 (
           que_out_21__1__9), .B1 (nx10158), .C0 (que_out_8__1__9), .C1 (nx10132
           )) ;
    aoi22 ix8966 (.Y (nx8965), .A0 (que_out_25__1__9), .A1 (nx10080), .B0 (
          que_out_16__1__9), .B1 (nx10106)) ;
    aoi22 ix8968 (.Y (nx8967), .A0 (que_out_24__1__9), .A1 (nx10054), .B0 (
          que_out_22__1__9), .B1 (nx10028)) ;
    nand03 ix6455 (.Y (nx6454), .A0 (nx8970), .A1 (nx8973), .A2 (nx8975)) ;
    aoi222 ix8972 (.Y (nx8970), .A0 (que_out_15__1__9), .A1 (nx9976), .B0 (
           que_out_3__1__9), .B1 (nx10002), .C0 (que_out_23__1__9), .C1 (nx9950)
           ) ;
    aoi22 ix8974 (.Y (nx8973), .A0 (que_out_27__1__9), .A1 (nx9924), .B0 (
          que_out_4__1__9), .B1 (nx9898)) ;
    aoi22 ix8976 (.Y (nx8975), .A0 (que_out_0__1__9), .A1 (nx9846), .B0 (
          que_out_2__1__9), .B1 (nx9872)) ;
    nand03 ix6429 (.Y (nx6428), .A0 (nx8978), .A1 (nx8981), .A2 (nx8983)) ;
    aoi222 ix8980 (.Y (nx8978), .A0 (que_out_26__1__9), .A1 (nx9820), .B0 (
           que_out_14__1__9), .B1 (nx9794), .C0 (que_out_11__1__9), .C1 (nx9768)
           ) ;
    aoi22 ix8982 (.Y (nx8981), .A0 (que_out_13__1__9), .A1 (nx9742), .B0 (
          que_out_7__1__9), .B1 (nx9716)) ;
    aoi22 ix8984 (.Y (nx8983), .A0 (que_out_12__1__9), .A1 (nx9690), .B0 (
          que_out_1__1__9), .B1 (nx9664)) ;
    or04 ix6623 (.Y (out_column_1__10), .A0 (nx6618), .A1 (nx6592), .A2 (nx6564)
         , .A3 (nx6538)) ;
    nand03 ix6619 (.Y (nx6618), .A0 (nx8989), .A1 (nx8991), .A2 (nx8993)) ;
    aoi222 ix8990 (.Y (nx8989), .A0 (que_out_10__1__10), .A1 (nx10314), .B0 (
           que_out_6__1__10), .B1 (nx10366), .C0 (que_out_9__1__10), .C1 (
           nx10340)) ;
    aoi22 ix8992 (.Y (nx8991), .A0 (que_out_5__1__10), .A1 (nx10262), .B0 (
          que_out_18__1__10), .B1 (nx10288)) ;
    aoi22 ix8994 (.Y (nx8993), .A0 (que_out_17__1__10), .A1 (nx10236), .B0 (
          que_out_20__1__10), .B1 (nx10210)) ;
    nand03 ix6593 (.Y (nx6592), .A0 (nx8997), .A1 (nx8999), .A2 (nx9001)) ;
    aoi222 ix8998 (.Y (nx8997), .A0 (que_out_19__1__10), .A1 (nx10184), .B0 (
           que_out_21__1__10), .B1 (nx10158), .C0 (que_out_8__1__10), .C1 (
           nx10132)) ;
    aoi22 ix9000 (.Y (nx8999), .A0 (que_out_25__1__10), .A1 (nx10080), .B0 (
          que_out_16__1__10), .B1 (nx10106)) ;
    aoi22 ix9002 (.Y (nx9001), .A0 (que_out_24__1__10), .A1 (nx10054), .B0 (
          que_out_22__1__10), .B1 (nx10028)) ;
    nand03 ix6565 (.Y (nx6564), .A0 (nx9005), .A1 (nx9007), .A2 (nx9009)) ;
    aoi222 ix9006 (.Y (nx9005), .A0 (que_out_15__1__10), .A1 (nx9976), .B0 (
           que_out_3__1__10), .B1 (nx10002), .C0 (que_out_23__1__10), .C1 (
           nx9950)) ;
    aoi22 ix9008 (.Y (nx9007), .A0 (que_out_27__1__10), .A1 (nx9924), .B0 (
          que_out_4__1__10), .B1 (nx9898)) ;
    aoi22 ix9010 (.Y (nx9009), .A0 (que_out_0__1__10), .A1 (nx9846), .B0 (
          que_out_2__1__10), .B1 (nx9872)) ;
    nand03 ix6539 (.Y (nx6538), .A0 (nx9013), .A1 (nx9015), .A2 (nx9017)) ;
    aoi222 ix9014 (.Y (nx9013), .A0 (que_out_26__1__10), .A1 (nx9820), .B0 (
           que_out_14__1__10), .B1 (nx9794), .C0 (que_out_11__1__10), .C1 (
           nx9768)) ;
    aoi22 ix9016 (.Y (nx9015), .A0 (que_out_13__1__10), .A1 (nx9742), .B0 (
          que_out_7__1__10), .B1 (nx9716)) ;
    aoi22 ix9018 (.Y (nx9017), .A0 (que_out_12__1__10), .A1 (nx9690), .B0 (
          que_out_1__1__10), .B1 (nx9664)) ;
    or04 ix6733 (.Y (out_column_1__11), .A0 (nx6728), .A1 (nx6702), .A2 (nx6674)
         , .A3 (nx6648)) ;
    nand03 ix6729 (.Y (nx6728), .A0 (nx9023), .A1 (nx9025), .A2 (nx9027)) ;
    aoi222 ix9024 (.Y (nx9023), .A0 (que_out_10__1__11), .A1 (nx10314), .B0 (
           que_out_6__1__11), .B1 (nx10366), .C0 (que_out_9__1__11), .C1 (
           nx10340)) ;
    aoi22 ix9026 (.Y (nx9025), .A0 (que_out_5__1__11), .A1 (nx10262), .B0 (
          que_out_18__1__11), .B1 (nx10288)) ;
    aoi22 ix9028 (.Y (nx9027), .A0 (que_out_17__1__11), .A1 (nx10236), .B0 (
          que_out_20__1__11), .B1 (nx10210)) ;
    nand03 ix6703 (.Y (nx6702), .A0 (nx9031), .A1 (nx9033), .A2 (nx9035)) ;
    aoi222 ix9032 (.Y (nx9031), .A0 (que_out_19__1__11), .A1 (nx10184), .B0 (
           que_out_21__1__11), .B1 (nx10158), .C0 (que_out_8__1__11), .C1 (
           nx10132)) ;
    aoi22 ix9034 (.Y (nx9033), .A0 (que_out_25__1__11), .A1 (nx10080), .B0 (
          que_out_16__1__11), .B1 (nx10106)) ;
    aoi22 ix9036 (.Y (nx9035), .A0 (que_out_24__1__11), .A1 (nx10054), .B0 (
          que_out_22__1__11), .B1 (nx10028)) ;
    nand03 ix6675 (.Y (nx6674), .A0 (nx9039), .A1 (nx9041), .A2 (nx9043)) ;
    aoi222 ix9040 (.Y (nx9039), .A0 (que_out_15__1__11), .A1 (nx9976), .B0 (
           que_out_3__1__11), .B1 (nx10002), .C0 (que_out_23__1__11), .C1 (
           nx9950)) ;
    aoi22 ix9042 (.Y (nx9041), .A0 (que_out_27__1__11), .A1 (nx9924), .B0 (
          que_out_4__1__11), .B1 (nx9898)) ;
    aoi22 ix9044 (.Y (nx9043), .A0 (que_out_0__1__11), .A1 (nx9846), .B0 (
          que_out_2__1__11), .B1 (nx9872)) ;
    nand03 ix6649 (.Y (nx6648), .A0 (nx9047), .A1 (nx9049), .A2 (nx9051)) ;
    aoi222 ix9048 (.Y (nx9047), .A0 (que_out_26__1__11), .A1 (nx9820), .B0 (
           que_out_14__1__11), .B1 (nx9794), .C0 (que_out_11__1__11), .C1 (
           nx9768)) ;
    aoi22 ix9050 (.Y (nx9049), .A0 (que_out_13__1__11), .A1 (nx9742), .B0 (
          que_out_7__1__11), .B1 (nx9716)) ;
    aoi22 ix9052 (.Y (nx9051), .A0 (que_out_12__1__11), .A1 (nx9690), .B0 (
          que_out_1__1__11), .B1 (nx9664)) ;
    or04 ix6843 (.Y (out_column_1__12), .A0 (nx6838), .A1 (nx6812), .A2 (nx6784)
         , .A3 (nx6758)) ;
    nand03 ix6839 (.Y (nx6838), .A0 (nx9057), .A1 (nx9059), .A2 (nx9061)) ;
    aoi222 ix9058 (.Y (nx9057), .A0 (que_out_10__1__12), .A1 (nx10314), .B0 (
           que_out_6__1__12), .B1 (nx10366), .C0 (que_out_9__1__12), .C1 (
           nx10340)) ;
    aoi22 ix9060 (.Y (nx9059), .A0 (que_out_5__1__12), .A1 (nx10262), .B0 (
          que_out_18__1__12), .B1 (nx10288)) ;
    aoi22 ix9062 (.Y (nx9061), .A0 (que_out_17__1__12), .A1 (nx10236), .B0 (
          que_out_20__1__12), .B1 (nx10210)) ;
    nand03 ix6813 (.Y (nx6812), .A0 (nx9065), .A1 (nx9067), .A2 (nx9069)) ;
    aoi222 ix9066 (.Y (nx9065), .A0 (que_out_19__1__12), .A1 (nx10184), .B0 (
           que_out_21__1__12), .B1 (nx10158), .C0 (que_out_8__1__12), .C1 (
           nx10132)) ;
    aoi22 ix9068 (.Y (nx9067), .A0 (que_out_25__1__12), .A1 (nx10080), .B0 (
          que_out_16__1__12), .B1 (nx10106)) ;
    aoi22 ix9070 (.Y (nx9069), .A0 (que_out_24__1__12), .A1 (nx10054), .B0 (
          que_out_22__1__12), .B1 (nx10028)) ;
    nand03 ix6785 (.Y (nx6784), .A0 (nx9073), .A1 (nx9075), .A2 (nx9077)) ;
    aoi222 ix9074 (.Y (nx9073), .A0 (que_out_15__1__12), .A1 (nx9976), .B0 (
           que_out_3__1__12), .B1 (nx10002), .C0 (que_out_23__1__12), .C1 (
           nx9950)) ;
    aoi22 ix9076 (.Y (nx9075), .A0 (que_out_27__1__12), .A1 (nx9924), .B0 (
          que_out_4__1__12), .B1 (nx9898)) ;
    aoi22 ix9078 (.Y (nx9077), .A0 (que_out_0__1__12), .A1 (nx9846), .B0 (
          que_out_2__1__12), .B1 (nx9872)) ;
    nand03 ix6759 (.Y (nx6758), .A0 (nx9081), .A1 (nx9083), .A2 (nx9085)) ;
    aoi222 ix9082 (.Y (nx9081), .A0 (que_out_26__1__12), .A1 (nx9820), .B0 (
           que_out_14__1__12), .B1 (nx9794), .C0 (que_out_11__1__12), .C1 (
           nx9768)) ;
    aoi22 ix9084 (.Y (nx9083), .A0 (que_out_13__1__12), .A1 (nx9742), .B0 (
          que_out_7__1__12), .B1 (nx9716)) ;
    aoi22 ix9086 (.Y (nx9085), .A0 (que_out_12__1__12), .A1 (nx9690), .B0 (
          que_out_1__1__12), .B1 (nx9664)) ;
    or04 ix6953 (.Y (out_column_1__13), .A0 (nx6948), .A1 (nx6922), .A2 (nx6894)
         , .A3 (nx6868)) ;
    nand03 ix6949 (.Y (nx6948), .A0 (nx9090), .A1 (nx9093), .A2 (nx9095)) ;
    aoi222 ix9092 (.Y (nx9090), .A0 (que_out_10__1__13), .A1 (nx10314), .B0 (
           que_out_6__1__13), .B1 (nx10366), .C0 (que_out_9__1__13), .C1 (
           nx10340)) ;
    aoi22 ix9094 (.Y (nx9093), .A0 (que_out_5__1__13), .A1 (nx10262), .B0 (
          que_out_18__1__13), .B1 (nx10288)) ;
    aoi22 ix9096 (.Y (nx9095), .A0 (que_out_17__1__13), .A1 (nx10236), .B0 (
          que_out_20__1__13), .B1 (nx10210)) ;
    nand03 ix6923 (.Y (nx6922), .A0 (nx9098), .A1 (nx9101), .A2 (nx9103)) ;
    aoi222 ix9100 (.Y (nx9098), .A0 (que_out_19__1__13), .A1 (nx10184), .B0 (
           que_out_21__1__13), .B1 (nx10158), .C0 (que_out_8__1__13), .C1 (
           nx10132)) ;
    aoi22 ix9102 (.Y (nx9101), .A0 (que_out_25__1__13), .A1 (nx10080), .B0 (
          que_out_16__1__13), .B1 (nx10106)) ;
    aoi22 ix9104 (.Y (nx9103), .A0 (que_out_24__1__13), .A1 (nx10054), .B0 (
          que_out_22__1__13), .B1 (nx10028)) ;
    nand03 ix6895 (.Y (nx6894), .A0 (nx9106), .A1 (nx9108), .A2 (nx9110)) ;
    aoi222 ix9107 (.Y (nx9106), .A0 (que_out_15__1__13), .A1 (nx9976), .B0 (
           que_out_3__1__13), .B1 (nx10002), .C0 (que_out_23__1__13), .C1 (
           nx9950)) ;
    aoi22 ix9109 (.Y (nx9108), .A0 (que_out_27__1__13), .A1 (nx9924), .B0 (
          que_out_4__1__13), .B1 (nx9898)) ;
    aoi22 ix9111 (.Y (nx9110), .A0 (que_out_0__1__13), .A1 (nx9846), .B0 (
          que_out_2__1__13), .B1 (nx9872)) ;
    nand03 ix6869 (.Y (nx6868), .A0 (nx9113), .A1 (nx9115), .A2 (nx9117)) ;
    aoi222 ix9114 (.Y (nx9113), .A0 (que_out_26__1__13), .A1 (nx9820), .B0 (
           que_out_14__1__13), .B1 (nx9794), .C0 (que_out_11__1__13), .C1 (
           nx9768)) ;
    aoi22 ix9116 (.Y (nx9115), .A0 (que_out_13__1__13), .A1 (nx9742), .B0 (
          que_out_7__1__13), .B1 (nx9716)) ;
    aoi22 ix9118 (.Y (nx9117), .A0 (que_out_12__1__13), .A1 (nx9690), .B0 (
          que_out_1__1__13), .B1 (nx9664)) ;
    or04 ix7063 (.Y (out_column_1__14), .A0 (nx7058), .A1 (nx7032), .A2 (nx7004)
         , .A3 (nx6978)) ;
    nand03 ix7059 (.Y (nx7058), .A0 (nx9121), .A1 (nx9123), .A2 (nx9125)) ;
    aoi222 ix9122 (.Y (nx9121), .A0 (que_out_10__1__14), .A1 (nx10314), .B0 (
           que_out_6__1__14), .B1 (nx10366), .C0 (que_out_9__1__14), .C1 (
           nx10340)) ;
    aoi22 ix9124 (.Y (nx9123), .A0 (que_out_5__1__14), .A1 (nx10262), .B0 (
          que_out_18__1__14), .B1 (nx10288)) ;
    aoi22 ix9126 (.Y (nx9125), .A0 (que_out_17__1__14), .A1 (nx10236), .B0 (
          que_out_20__1__14), .B1 (nx10210)) ;
    nand03 ix7033 (.Y (nx7032), .A0 (nx9128), .A1 (nx9130), .A2 (nx9132)) ;
    aoi222 ix9129 (.Y (nx9128), .A0 (que_out_19__1__14), .A1 (nx10184), .B0 (
           que_out_21__1__14), .B1 (nx10158), .C0 (que_out_8__1__14), .C1 (
           nx10132)) ;
    aoi22 ix9131 (.Y (nx9130), .A0 (que_out_25__1__14), .A1 (nx10080), .B0 (
          que_out_16__1__14), .B1 (nx10106)) ;
    aoi22 ix9133 (.Y (nx9132), .A0 (que_out_24__1__14), .A1 (nx10054), .B0 (
          que_out_22__1__14), .B1 (nx10028)) ;
    nand03 ix7005 (.Y (nx7004), .A0 (nx9135), .A1 (nx9137), .A2 (nx9139)) ;
    aoi222 ix9136 (.Y (nx9135), .A0 (que_out_15__1__14), .A1 (nx9976), .B0 (
           que_out_3__1__14), .B1 (nx10002), .C0 (que_out_23__1__14), .C1 (
           nx9950)) ;
    aoi22 ix9138 (.Y (nx9137), .A0 (que_out_27__1__14), .A1 (nx9924), .B0 (
          que_out_4__1__14), .B1 (nx9898)) ;
    aoi22 ix9140 (.Y (nx9139), .A0 (que_out_0__1__14), .A1 (nx9846), .B0 (
          que_out_2__1__14), .B1 (nx9872)) ;
    nand03 ix6979 (.Y (nx6978), .A0 (nx9142), .A1 (nx9144), .A2 (nx9146)) ;
    aoi222 ix9143 (.Y (nx9142), .A0 (que_out_26__1__14), .A1 (nx9820), .B0 (
           que_out_14__1__14), .B1 (nx9794), .C0 (que_out_11__1__14), .C1 (
           nx9768)) ;
    aoi22 ix9145 (.Y (nx9144), .A0 (que_out_13__1__14), .A1 (nx9742), .B0 (
          que_out_7__1__14), .B1 (nx9716)) ;
    aoi22 ix9147 (.Y (nx9146), .A0 (que_out_12__1__14), .A1 (nx9690), .B0 (
          que_out_1__1__14), .B1 (nx9664)) ;
    or04 ix7173 (.Y (out_column_1__15), .A0 (nx7168), .A1 (nx7142), .A2 (nx7114)
         , .A3 (nx7088)) ;
    nand03 ix7169 (.Y (nx7168), .A0 (nx9150), .A1 (nx9152), .A2 (nx9154)) ;
    aoi222 ix9151 (.Y (nx9150), .A0 (que_out_10__1__15), .A1 (nx10316), .B0 (
           que_out_6__1__15), .B1 (nx10368), .C0 (que_out_9__1__15), .C1 (
           nx10342)) ;
    aoi22 ix9153 (.Y (nx9152), .A0 (que_out_5__1__15), .A1 (nx10264), .B0 (
          que_out_18__1__15), .B1 (nx10290)) ;
    aoi22 ix9155 (.Y (nx9154), .A0 (que_out_17__1__15), .A1 (nx10238), .B0 (
          que_out_20__1__15), .B1 (nx10212)) ;
    nand03 ix7143 (.Y (nx7142), .A0 (nx9157), .A1 (nx9159), .A2 (nx9161)) ;
    aoi222 ix9158 (.Y (nx9157), .A0 (que_out_19__1__15), .A1 (nx10186), .B0 (
           que_out_21__1__15), .B1 (nx10160), .C0 (que_out_8__1__15), .C1 (
           nx10134)) ;
    aoi22 ix9160 (.Y (nx9159), .A0 (que_out_25__1__15), .A1 (nx10082), .B0 (
          que_out_16__1__15), .B1 (nx10108)) ;
    aoi22 ix9162 (.Y (nx9161), .A0 (que_out_24__1__15), .A1 (nx10056), .B0 (
          que_out_22__1__15), .B1 (nx10030)) ;
    nand03 ix7115 (.Y (nx7114), .A0 (nx9164), .A1 (nx9166), .A2 (nx9168)) ;
    aoi222 ix9165 (.Y (nx9164), .A0 (que_out_15__1__15), .A1 (nx9978), .B0 (
           que_out_3__1__15), .B1 (nx10004), .C0 (que_out_23__1__15), .C1 (
           nx9952)) ;
    aoi22 ix9167 (.Y (nx9166), .A0 (que_out_27__1__15), .A1 (nx9926), .B0 (
          que_out_4__1__15), .B1 (nx9900)) ;
    aoi22 ix9169 (.Y (nx9168), .A0 (que_out_0__1__15), .A1 (nx9848), .B0 (
          que_out_2__1__15), .B1 (nx9874)) ;
    nand03 ix7089 (.Y (nx7088), .A0 (nx9171), .A1 (nx9173), .A2 (nx9175)) ;
    aoi222 ix9172 (.Y (nx9171), .A0 (que_out_26__1__15), .A1 (nx9822), .B0 (
           que_out_14__1__15), .B1 (nx9796), .C0 (que_out_11__1__15), .C1 (
           nx9770)) ;
    aoi22 ix9174 (.Y (nx9173), .A0 (que_out_13__1__15), .A1 (nx9744), .B0 (
          que_out_7__1__15), .B1 (nx9718)) ;
    aoi22 ix9176 (.Y (nx9175), .A0 (que_out_12__1__15), .A1 (nx9692), .B0 (
          que_out_1__1__15), .B1 (nx9666)) ;
    or04 ix7283 (.Y (out_column_0__0), .A0 (nx7278), .A1 (nx7252), .A2 (nx7224)
         , .A3 (nx7198)) ;
    nand03 ix7279 (.Y (nx7278), .A0 (nx9179), .A1 (nx9181), .A2 (nx9183)) ;
    aoi222 ix9180 (.Y (nx9179), .A0 (que_out_10__0__0), .A1 (nx10316), .B0 (
           que_out_6__0__0), .B1 (nx10368), .C0 (que_out_9__0__0), .C1 (nx10342)
           ) ;
    aoi22 ix9182 (.Y (nx9181), .A0 (que_out_5__0__0), .A1 (nx10264), .B0 (
          que_out_18__0__0), .B1 (nx10290)) ;
    aoi22 ix9184 (.Y (nx9183), .A0 (que_out_17__0__0), .A1 (nx10238), .B0 (
          que_out_20__0__0), .B1 (nx10212)) ;
    nand03 ix7253 (.Y (nx7252), .A0 (nx9186), .A1 (nx9188), .A2 (nx9190)) ;
    aoi222 ix9187 (.Y (nx9186), .A0 (que_out_19__0__0), .A1 (nx10186), .B0 (
           que_out_21__0__0), .B1 (nx10160), .C0 (que_out_8__0__0), .C1 (nx10134
           )) ;
    aoi22 ix9189 (.Y (nx9188), .A0 (que_out_25__0__0), .A1 (nx10082), .B0 (
          que_out_16__0__0), .B1 (nx10108)) ;
    aoi22 ix9191 (.Y (nx9190), .A0 (que_out_24__0__0), .A1 (nx10056), .B0 (
          que_out_22__0__0), .B1 (nx10030)) ;
    nand03 ix7225 (.Y (nx7224), .A0 (nx9193), .A1 (nx9195), .A2 (nx9197)) ;
    aoi222 ix9194 (.Y (nx9193), .A0 (que_out_15__0__0), .A1 (nx9978), .B0 (
           que_out_3__0__0), .B1 (nx10004), .C0 (que_out_23__0__0), .C1 (nx9952)
           ) ;
    aoi22 ix9196 (.Y (nx9195), .A0 (que_out_27__0__0), .A1 (nx9926), .B0 (
          que_out_4__0__0), .B1 (nx9900)) ;
    aoi22 ix9198 (.Y (nx9197), .A0 (que_out_0__0__0), .A1 (nx9848), .B0 (
          que_out_2__0__0), .B1 (nx9874)) ;
    nand03 ix7199 (.Y (nx7198), .A0 (nx9200), .A1 (nx9202), .A2 (nx9204)) ;
    aoi222 ix9201 (.Y (nx9200), .A0 (que_out_26__0__0), .A1 (nx9822), .B0 (
           que_out_14__0__0), .B1 (nx9796), .C0 (que_out_11__0__0), .C1 (nx9770)
           ) ;
    aoi22 ix9203 (.Y (nx9202), .A0 (que_out_13__0__0), .A1 (nx9744), .B0 (
          que_out_7__0__0), .B1 (nx9718)) ;
    aoi22 ix9205 (.Y (nx9204), .A0 (que_out_12__0__0), .A1 (nx9692), .B0 (
          que_out_1__0__0), .B1 (nx9666)) ;
    or04 ix7393 (.Y (out_column_0__1), .A0 (nx7388), .A1 (nx7362), .A2 (nx7334)
         , .A3 (nx7308)) ;
    nand03 ix7389 (.Y (nx7388), .A0 (nx9208), .A1 (nx9210), .A2 (nx9212)) ;
    aoi222 ix9209 (.Y (nx9208), .A0 (que_out_10__0__1), .A1 (nx10316), .B0 (
           que_out_6__0__1), .B1 (nx10368), .C0 (que_out_9__0__1), .C1 (nx10342)
           ) ;
    aoi22 ix9211 (.Y (nx9210), .A0 (que_out_5__0__1), .A1 (nx10264), .B0 (
          que_out_18__0__1), .B1 (nx10290)) ;
    aoi22 ix9213 (.Y (nx9212), .A0 (que_out_17__0__1), .A1 (nx10238), .B0 (
          que_out_20__0__1), .B1 (nx10212)) ;
    nand03 ix7363 (.Y (nx7362), .A0 (nx9215), .A1 (nx9217), .A2 (nx9219)) ;
    aoi222 ix9216 (.Y (nx9215), .A0 (que_out_19__0__1), .A1 (nx10186), .B0 (
           que_out_21__0__1), .B1 (nx10160), .C0 (que_out_8__0__1), .C1 (nx10134
           )) ;
    aoi22 ix9218 (.Y (nx9217), .A0 (que_out_25__0__1), .A1 (nx10082), .B0 (
          que_out_16__0__1), .B1 (nx10108)) ;
    aoi22 ix9220 (.Y (nx9219), .A0 (que_out_24__0__1), .A1 (nx10056), .B0 (
          que_out_22__0__1), .B1 (nx10030)) ;
    nand03 ix7335 (.Y (nx7334), .A0 (nx9222), .A1 (nx9224), .A2 (nx9226)) ;
    aoi222 ix9223 (.Y (nx9222), .A0 (que_out_15__0__1), .A1 (nx9978), .B0 (
           que_out_3__0__1), .B1 (nx10004), .C0 (que_out_23__0__1), .C1 (nx9952)
           ) ;
    aoi22 ix9225 (.Y (nx9224), .A0 (que_out_27__0__1), .A1 (nx9926), .B0 (
          que_out_4__0__1), .B1 (nx9900)) ;
    aoi22 ix9227 (.Y (nx9226), .A0 (que_out_0__0__1), .A1 (nx9848), .B0 (
          que_out_2__0__1), .B1 (nx9874)) ;
    nand03 ix7309 (.Y (nx7308), .A0 (nx9229), .A1 (nx9231), .A2 (nx9233)) ;
    aoi222 ix9230 (.Y (nx9229), .A0 (que_out_26__0__1), .A1 (nx9822), .B0 (
           que_out_14__0__1), .B1 (nx9796), .C0 (que_out_11__0__1), .C1 (nx9770)
           ) ;
    aoi22 ix9232 (.Y (nx9231), .A0 (que_out_13__0__1), .A1 (nx9744), .B0 (
          que_out_7__0__1), .B1 (nx9718)) ;
    aoi22 ix9234 (.Y (nx9233), .A0 (que_out_12__0__1), .A1 (nx9692), .B0 (
          que_out_1__0__1), .B1 (nx9666)) ;
    or04 ix7503 (.Y (out_column_0__2), .A0 (nx7498), .A1 (nx7472), .A2 (nx7444)
         , .A3 (nx7418)) ;
    nand03 ix7499 (.Y (nx7498), .A0 (nx9237), .A1 (nx9239), .A2 (nx9241)) ;
    aoi222 ix9238 (.Y (nx9237), .A0 (que_out_10__0__2), .A1 (nx10316), .B0 (
           que_out_6__0__2), .B1 (nx10368), .C0 (que_out_9__0__2), .C1 (nx10342)
           ) ;
    aoi22 ix9240 (.Y (nx9239), .A0 (que_out_5__0__2), .A1 (nx10264), .B0 (
          que_out_18__0__2), .B1 (nx10290)) ;
    aoi22 ix9242 (.Y (nx9241), .A0 (que_out_17__0__2), .A1 (nx10238), .B0 (
          que_out_20__0__2), .B1 (nx10212)) ;
    nand03 ix7473 (.Y (nx7472), .A0 (nx9244), .A1 (nx9246), .A2 (nx9248)) ;
    aoi222 ix9245 (.Y (nx9244), .A0 (que_out_19__0__2), .A1 (nx10186), .B0 (
           que_out_21__0__2), .B1 (nx10160), .C0 (que_out_8__0__2), .C1 (nx10134
           )) ;
    aoi22 ix9247 (.Y (nx9246), .A0 (que_out_25__0__2), .A1 (nx10082), .B0 (
          que_out_16__0__2), .B1 (nx10108)) ;
    aoi22 ix9249 (.Y (nx9248), .A0 (que_out_24__0__2), .A1 (nx10056), .B0 (
          que_out_22__0__2), .B1 (nx10030)) ;
    nand03 ix7445 (.Y (nx7444), .A0 (nx9251), .A1 (nx9253), .A2 (nx9255)) ;
    aoi222 ix9252 (.Y (nx9251), .A0 (que_out_15__0__2), .A1 (nx9978), .B0 (
           que_out_3__0__2), .B1 (nx10004), .C0 (que_out_23__0__2), .C1 (nx9952)
           ) ;
    aoi22 ix9254 (.Y (nx9253), .A0 (que_out_27__0__2), .A1 (nx9926), .B0 (
          que_out_4__0__2), .B1 (nx9900)) ;
    aoi22 ix9256 (.Y (nx9255), .A0 (que_out_0__0__2), .A1 (nx9848), .B0 (
          que_out_2__0__2), .B1 (nx9874)) ;
    nand03 ix7419 (.Y (nx7418), .A0 (nx9258), .A1 (nx9260), .A2 (nx9262)) ;
    aoi222 ix9259 (.Y (nx9258), .A0 (que_out_26__0__2), .A1 (nx9822), .B0 (
           que_out_14__0__2), .B1 (nx9796), .C0 (que_out_11__0__2), .C1 (nx9770)
           ) ;
    aoi22 ix9261 (.Y (nx9260), .A0 (que_out_13__0__2), .A1 (nx9744), .B0 (
          que_out_7__0__2), .B1 (nx9718)) ;
    aoi22 ix9263 (.Y (nx9262), .A0 (que_out_12__0__2), .A1 (nx9692), .B0 (
          que_out_1__0__2), .B1 (nx9666)) ;
    or04 ix7613 (.Y (out_column_0__3), .A0 (nx7608), .A1 (nx7582), .A2 (nx7554)
         , .A3 (nx7528)) ;
    nand03 ix7609 (.Y (nx7608), .A0 (nx9266), .A1 (nx9268), .A2 (nx9270)) ;
    aoi222 ix9267 (.Y (nx9266), .A0 (que_out_10__0__3), .A1 (nx10316), .B0 (
           que_out_6__0__3), .B1 (nx10368), .C0 (que_out_9__0__3), .C1 (nx10342)
           ) ;
    aoi22 ix9269 (.Y (nx9268), .A0 (que_out_5__0__3), .A1 (nx10264), .B0 (
          que_out_18__0__3), .B1 (nx10290)) ;
    aoi22 ix9271 (.Y (nx9270), .A0 (que_out_17__0__3), .A1 (nx10238), .B0 (
          que_out_20__0__3), .B1 (nx10212)) ;
    nand03 ix7583 (.Y (nx7582), .A0 (nx9273), .A1 (nx9275), .A2 (nx9277)) ;
    aoi222 ix9274 (.Y (nx9273), .A0 (que_out_19__0__3), .A1 (nx10186), .B0 (
           que_out_21__0__3), .B1 (nx10160), .C0 (que_out_8__0__3), .C1 (nx10134
           )) ;
    aoi22 ix9276 (.Y (nx9275), .A0 (que_out_25__0__3), .A1 (nx10082), .B0 (
          que_out_16__0__3), .B1 (nx10108)) ;
    aoi22 ix9278 (.Y (nx9277), .A0 (que_out_24__0__3), .A1 (nx10056), .B0 (
          que_out_22__0__3), .B1 (nx10030)) ;
    nand03 ix7555 (.Y (nx7554), .A0 (nx9280), .A1 (nx9282), .A2 (nx9284)) ;
    aoi222 ix9281 (.Y (nx9280), .A0 (que_out_15__0__3), .A1 (nx9978), .B0 (
           que_out_3__0__3), .B1 (nx10004), .C0 (que_out_23__0__3), .C1 (nx9952)
           ) ;
    aoi22 ix9283 (.Y (nx9282), .A0 (que_out_27__0__3), .A1 (nx9926), .B0 (
          que_out_4__0__3), .B1 (nx9900)) ;
    aoi22 ix9285 (.Y (nx9284), .A0 (que_out_0__0__3), .A1 (nx9848), .B0 (
          que_out_2__0__3), .B1 (nx9874)) ;
    nand03 ix7529 (.Y (nx7528), .A0 (nx9287), .A1 (nx9289), .A2 (nx9291)) ;
    aoi222 ix9288 (.Y (nx9287), .A0 (que_out_26__0__3), .A1 (nx9822), .B0 (
           que_out_14__0__3), .B1 (nx9796), .C0 (que_out_11__0__3), .C1 (nx9770)
           ) ;
    aoi22 ix9290 (.Y (nx9289), .A0 (que_out_13__0__3), .A1 (nx9744), .B0 (
          que_out_7__0__3), .B1 (nx9718)) ;
    aoi22 ix9292 (.Y (nx9291), .A0 (que_out_12__0__3), .A1 (nx9692), .B0 (
          que_out_1__0__3), .B1 (nx9666)) ;
    or04 ix7723 (.Y (out_column_0__4), .A0 (nx7718), .A1 (nx7692), .A2 (nx7664)
         , .A3 (nx7638)) ;
    nand03 ix7719 (.Y (nx7718), .A0 (nx9295), .A1 (nx9297), .A2 (nx9299)) ;
    aoi222 ix9296 (.Y (nx9295), .A0 (que_out_10__0__4), .A1 (nx10316), .B0 (
           que_out_6__0__4), .B1 (nx10368), .C0 (que_out_9__0__4), .C1 (nx10342)
           ) ;
    aoi22 ix9298 (.Y (nx9297), .A0 (que_out_5__0__4), .A1 (nx10264), .B0 (
          que_out_18__0__4), .B1 (nx10290)) ;
    aoi22 ix9300 (.Y (nx9299), .A0 (que_out_17__0__4), .A1 (nx10238), .B0 (
          que_out_20__0__4), .B1 (nx10212)) ;
    nand03 ix7693 (.Y (nx7692), .A0 (nx9302), .A1 (nx9304), .A2 (nx9306)) ;
    aoi222 ix9303 (.Y (nx9302), .A0 (que_out_19__0__4), .A1 (nx10186), .B0 (
           que_out_21__0__4), .B1 (nx10160), .C0 (que_out_8__0__4), .C1 (nx10134
           )) ;
    aoi22 ix9305 (.Y (nx9304), .A0 (que_out_25__0__4), .A1 (nx10082), .B0 (
          que_out_16__0__4), .B1 (nx10108)) ;
    aoi22 ix9307 (.Y (nx9306), .A0 (que_out_24__0__4), .A1 (nx10056), .B0 (
          que_out_22__0__4), .B1 (nx10030)) ;
    nand03 ix7665 (.Y (nx7664), .A0 (nx9309), .A1 (nx9311), .A2 (nx9313)) ;
    aoi222 ix9310 (.Y (nx9309), .A0 (que_out_15__0__4), .A1 (nx9978), .B0 (
           que_out_3__0__4), .B1 (nx10004), .C0 (que_out_23__0__4), .C1 (nx9952)
           ) ;
    aoi22 ix9312 (.Y (nx9311), .A0 (que_out_27__0__4), .A1 (nx9926), .B0 (
          que_out_4__0__4), .B1 (nx9900)) ;
    aoi22 ix9314 (.Y (nx9313), .A0 (que_out_0__0__4), .A1 (nx9848), .B0 (
          que_out_2__0__4), .B1 (nx9874)) ;
    nand03 ix7639 (.Y (nx7638), .A0 (nx9316), .A1 (nx9318), .A2 (nx9320)) ;
    aoi222 ix9317 (.Y (nx9316), .A0 (que_out_26__0__4), .A1 (nx9822), .B0 (
           que_out_14__0__4), .B1 (nx9796), .C0 (que_out_11__0__4), .C1 (nx9770)
           ) ;
    aoi22 ix9319 (.Y (nx9318), .A0 (que_out_13__0__4), .A1 (nx9744), .B0 (
          que_out_7__0__4), .B1 (nx9718)) ;
    aoi22 ix9321 (.Y (nx9320), .A0 (que_out_12__0__4), .A1 (nx9692), .B0 (
          que_out_1__0__4), .B1 (nx9666)) ;
    or04 ix7833 (.Y (out_column_0__5), .A0 (nx7828), .A1 (nx7802), .A2 (nx7774)
         , .A3 (nx7748)) ;
    nand03 ix7829 (.Y (nx7828), .A0 (nx9324), .A1 (nx9326), .A2 (nx9328)) ;
    aoi222 ix9325 (.Y (nx9324), .A0 (que_out_10__0__5), .A1 (nx10316), .B0 (
           que_out_6__0__5), .B1 (nx10368), .C0 (que_out_9__0__5), .C1 (nx10342)
           ) ;
    aoi22 ix9327 (.Y (nx9326), .A0 (que_out_5__0__5), .A1 (nx10264), .B0 (
          que_out_18__0__5), .B1 (nx10290)) ;
    aoi22 ix9329 (.Y (nx9328), .A0 (que_out_17__0__5), .A1 (nx10238), .B0 (
          que_out_20__0__5), .B1 (nx10212)) ;
    nand03 ix7803 (.Y (nx7802), .A0 (nx9331), .A1 (nx9333), .A2 (nx9335)) ;
    aoi222 ix9332 (.Y (nx9331), .A0 (que_out_19__0__5), .A1 (nx10186), .B0 (
           que_out_21__0__5), .B1 (nx10160), .C0 (que_out_8__0__5), .C1 (nx10134
           )) ;
    aoi22 ix9334 (.Y (nx9333), .A0 (que_out_25__0__5), .A1 (nx10082), .B0 (
          que_out_16__0__5), .B1 (nx10108)) ;
    aoi22 ix9336 (.Y (nx9335), .A0 (que_out_24__0__5), .A1 (nx10056), .B0 (
          que_out_22__0__5), .B1 (nx10030)) ;
    nand03 ix7775 (.Y (nx7774), .A0 (nx9338), .A1 (nx9340), .A2 (nx9342)) ;
    aoi222 ix9339 (.Y (nx9338), .A0 (que_out_15__0__5), .A1 (nx9978), .B0 (
           que_out_3__0__5), .B1 (nx10004), .C0 (que_out_23__0__5), .C1 (nx9952)
           ) ;
    aoi22 ix9341 (.Y (nx9340), .A0 (que_out_27__0__5), .A1 (nx9926), .B0 (
          que_out_4__0__5), .B1 (nx9900)) ;
    aoi22 ix9343 (.Y (nx9342), .A0 (que_out_0__0__5), .A1 (nx9848), .B0 (
          que_out_2__0__5), .B1 (nx9874)) ;
    nand03 ix7749 (.Y (nx7748), .A0 (nx9345), .A1 (nx9347), .A2 (nx9349)) ;
    aoi222 ix9346 (.Y (nx9345), .A0 (que_out_26__0__5), .A1 (nx9822), .B0 (
           que_out_14__0__5), .B1 (nx9796), .C0 (que_out_11__0__5), .C1 (nx9770)
           ) ;
    aoi22 ix9348 (.Y (nx9347), .A0 (que_out_13__0__5), .A1 (nx9744), .B0 (
          que_out_7__0__5), .B1 (nx9718)) ;
    aoi22 ix9350 (.Y (nx9349), .A0 (que_out_12__0__5), .A1 (nx9692), .B0 (
          que_out_1__0__5), .B1 (nx9666)) ;
    or04 ix7943 (.Y (out_column_0__6), .A0 (nx7938), .A1 (nx7912), .A2 (nx7884)
         , .A3 (nx7858)) ;
    nand03 ix7939 (.Y (nx7938), .A0 (nx9353), .A1 (nx9355), .A2 (nx9357)) ;
    aoi222 ix9354 (.Y (nx9353), .A0 (que_out_10__0__6), .A1 (nx10318), .B0 (
           que_out_6__0__6), .B1 (nx10370), .C0 (que_out_9__0__6), .C1 (nx10344)
           ) ;
    aoi22 ix9356 (.Y (nx9355), .A0 (que_out_5__0__6), .A1 (nx10266), .B0 (
          que_out_18__0__6), .B1 (nx10292)) ;
    aoi22 ix9358 (.Y (nx9357), .A0 (que_out_17__0__6), .A1 (nx10240), .B0 (
          que_out_20__0__6), .B1 (nx10214)) ;
    nand03 ix7913 (.Y (nx7912), .A0 (nx9360), .A1 (nx9362), .A2 (nx9364)) ;
    aoi222 ix9361 (.Y (nx9360), .A0 (que_out_19__0__6), .A1 (nx10188), .B0 (
           que_out_21__0__6), .B1 (nx10162), .C0 (que_out_8__0__6), .C1 (nx10136
           )) ;
    aoi22 ix9363 (.Y (nx9362), .A0 (que_out_25__0__6), .A1 (nx10084), .B0 (
          que_out_16__0__6), .B1 (nx10110)) ;
    aoi22 ix9365 (.Y (nx9364), .A0 (que_out_24__0__6), .A1 (nx10058), .B0 (
          que_out_22__0__6), .B1 (nx10032)) ;
    nand03 ix7885 (.Y (nx7884), .A0 (nx9367), .A1 (nx9369), .A2 (nx9371)) ;
    aoi222 ix9368 (.Y (nx9367), .A0 (que_out_15__0__6), .A1 (nx9980), .B0 (
           que_out_3__0__6), .B1 (nx10006), .C0 (que_out_23__0__6), .C1 (nx9954)
           ) ;
    aoi22 ix9370 (.Y (nx9369), .A0 (que_out_27__0__6), .A1 (nx9928), .B0 (
          que_out_4__0__6), .B1 (nx9902)) ;
    aoi22 ix9372 (.Y (nx9371), .A0 (que_out_0__0__6), .A1 (nx9850), .B0 (
          que_out_2__0__6), .B1 (nx9876)) ;
    nand03 ix7859 (.Y (nx7858), .A0 (nx9374), .A1 (nx9376), .A2 (nx9378)) ;
    aoi222 ix9375 (.Y (nx9374), .A0 (que_out_26__0__6), .A1 (nx9824), .B0 (
           que_out_14__0__6), .B1 (nx9798), .C0 (que_out_11__0__6), .C1 (nx9772)
           ) ;
    aoi22 ix9377 (.Y (nx9376), .A0 (que_out_13__0__6), .A1 (nx9746), .B0 (
          que_out_7__0__6), .B1 (nx9720)) ;
    aoi22 ix9379 (.Y (nx9378), .A0 (que_out_12__0__6), .A1 (nx9694), .B0 (
          que_out_1__0__6), .B1 (nx9668)) ;
    or04 ix8053 (.Y (out_column_0__7), .A0 (nx8048), .A1 (nx8022), .A2 (nx7994)
         , .A3 (nx7968)) ;
    nand03 ix8049 (.Y (nx8048), .A0 (nx9382), .A1 (nx9384), .A2 (nx9386)) ;
    aoi222 ix9383 (.Y (nx9382), .A0 (que_out_10__0__7), .A1 (nx10318), .B0 (
           que_out_6__0__7), .B1 (nx10370), .C0 (que_out_9__0__7), .C1 (nx10344)
           ) ;
    aoi22 ix9385 (.Y (nx9384), .A0 (que_out_5__0__7), .A1 (nx10266), .B0 (
          que_out_18__0__7), .B1 (nx10292)) ;
    aoi22 ix9387 (.Y (nx9386), .A0 (que_out_17__0__7), .A1 (nx10240), .B0 (
          que_out_20__0__7), .B1 (nx10214)) ;
    nand03 ix8023 (.Y (nx8022), .A0 (nx9389), .A1 (nx9391), .A2 (nx9393)) ;
    aoi222 ix9390 (.Y (nx9389), .A0 (que_out_19__0__7), .A1 (nx10188), .B0 (
           que_out_21__0__7), .B1 (nx10162), .C0 (que_out_8__0__7), .C1 (nx10136
           )) ;
    aoi22 ix9392 (.Y (nx9391), .A0 (que_out_25__0__7), .A1 (nx10084), .B0 (
          que_out_16__0__7), .B1 (nx10110)) ;
    aoi22 ix9394 (.Y (nx9393), .A0 (que_out_24__0__7), .A1 (nx10058), .B0 (
          que_out_22__0__7), .B1 (nx10032)) ;
    nand03 ix7995 (.Y (nx7994), .A0 (nx9396), .A1 (nx9398), .A2 (nx9400)) ;
    aoi222 ix9397 (.Y (nx9396), .A0 (que_out_15__0__7), .A1 (nx9980), .B0 (
           que_out_3__0__7), .B1 (nx10006), .C0 (que_out_23__0__7), .C1 (nx9954)
           ) ;
    aoi22 ix9399 (.Y (nx9398), .A0 (que_out_27__0__7), .A1 (nx9928), .B0 (
          que_out_4__0__7), .B1 (nx9902)) ;
    aoi22 ix9401 (.Y (nx9400), .A0 (que_out_0__0__7), .A1 (nx9850), .B0 (
          que_out_2__0__7), .B1 (nx9876)) ;
    nand03 ix7969 (.Y (nx7968), .A0 (nx9403), .A1 (nx9405), .A2 (nx9407)) ;
    aoi222 ix9404 (.Y (nx9403), .A0 (que_out_26__0__7), .A1 (nx9824), .B0 (
           que_out_14__0__7), .B1 (nx9798), .C0 (que_out_11__0__7), .C1 (nx9772)
           ) ;
    aoi22 ix9406 (.Y (nx9405), .A0 (que_out_13__0__7), .A1 (nx9746), .B0 (
          que_out_7__0__7), .B1 (nx9720)) ;
    aoi22 ix9408 (.Y (nx9407), .A0 (que_out_12__0__7), .A1 (nx9694), .B0 (
          que_out_1__0__7), .B1 (nx9668)) ;
    or04 ix8163 (.Y (out_column_0__8), .A0 (nx8158), .A1 (nx8132), .A2 (nx8104)
         , .A3 (nx8078)) ;
    nand03 ix8159 (.Y (nx8158), .A0 (nx9411), .A1 (nx9413), .A2 (nx9415)) ;
    aoi222 ix9412 (.Y (nx9411), .A0 (que_out_10__0__8), .A1 (nx10318), .B0 (
           que_out_6__0__8), .B1 (nx10370), .C0 (que_out_9__0__8), .C1 (nx10344)
           ) ;
    aoi22 ix9414 (.Y (nx9413), .A0 (que_out_5__0__8), .A1 (nx10266), .B0 (
          que_out_18__0__8), .B1 (nx10292)) ;
    aoi22 ix9416 (.Y (nx9415), .A0 (que_out_17__0__8), .A1 (nx10240), .B0 (
          que_out_20__0__8), .B1 (nx10214)) ;
    nand03 ix8133 (.Y (nx8132), .A0 (nx9418), .A1 (nx9420), .A2 (nx9422)) ;
    aoi222 ix9419 (.Y (nx9418), .A0 (que_out_19__0__8), .A1 (nx10188), .B0 (
           que_out_21__0__8), .B1 (nx10162), .C0 (que_out_8__0__8), .C1 (nx10136
           )) ;
    aoi22 ix9421 (.Y (nx9420), .A0 (que_out_25__0__8), .A1 (nx10084), .B0 (
          que_out_16__0__8), .B1 (nx10110)) ;
    aoi22 ix9423 (.Y (nx9422), .A0 (que_out_24__0__8), .A1 (nx10058), .B0 (
          que_out_22__0__8), .B1 (nx10032)) ;
    nand03 ix8105 (.Y (nx8104), .A0 (nx9425), .A1 (nx9427), .A2 (nx9429)) ;
    aoi222 ix9426 (.Y (nx9425), .A0 (que_out_15__0__8), .A1 (nx9980), .B0 (
           que_out_3__0__8), .B1 (nx10006), .C0 (que_out_23__0__8), .C1 (nx9954)
           ) ;
    aoi22 ix9428 (.Y (nx9427), .A0 (que_out_27__0__8), .A1 (nx9928), .B0 (
          que_out_4__0__8), .B1 (nx9902)) ;
    aoi22 ix9430 (.Y (nx9429), .A0 (que_out_0__0__8), .A1 (nx9850), .B0 (
          que_out_2__0__8), .B1 (nx9876)) ;
    nand03 ix8079 (.Y (nx8078), .A0 (nx9432), .A1 (nx9434), .A2 (nx9436)) ;
    aoi222 ix9433 (.Y (nx9432), .A0 (que_out_26__0__8), .A1 (nx9824), .B0 (
           que_out_14__0__8), .B1 (nx9798), .C0 (que_out_11__0__8), .C1 (nx9772)
           ) ;
    aoi22 ix9435 (.Y (nx9434), .A0 (que_out_13__0__8), .A1 (nx9746), .B0 (
          que_out_7__0__8), .B1 (nx9720)) ;
    aoi22 ix9437 (.Y (nx9436), .A0 (que_out_12__0__8), .A1 (nx9694), .B0 (
          que_out_1__0__8), .B1 (nx9668)) ;
    or04 ix8273 (.Y (out_column_0__9), .A0 (nx8268), .A1 (nx8242), .A2 (nx8214)
         , .A3 (nx8188)) ;
    nand03 ix8269 (.Y (nx8268), .A0 (nx9440), .A1 (nx9442), .A2 (nx9444)) ;
    aoi222 ix9441 (.Y (nx9440), .A0 (que_out_10__0__9), .A1 (nx10318), .B0 (
           que_out_6__0__9), .B1 (nx10370), .C0 (que_out_9__0__9), .C1 (nx10344)
           ) ;
    aoi22 ix9443 (.Y (nx9442), .A0 (que_out_5__0__9), .A1 (nx10266), .B0 (
          que_out_18__0__9), .B1 (nx10292)) ;
    aoi22 ix9445 (.Y (nx9444), .A0 (que_out_17__0__9), .A1 (nx10240), .B0 (
          que_out_20__0__9), .B1 (nx10214)) ;
    nand03 ix8243 (.Y (nx8242), .A0 (nx9447), .A1 (nx9449), .A2 (nx9451)) ;
    aoi222 ix9448 (.Y (nx9447), .A0 (que_out_19__0__9), .A1 (nx10188), .B0 (
           que_out_21__0__9), .B1 (nx10162), .C0 (que_out_8__0__9), .C1 (nx10136
           )) ;
    aoi22 ix9450 (.Y (nx9449), .A0 (que_out_25__0__9), .A1 (nx10084), .B0 (
          que_out_16__0__9), .B1 (nx10110)) ;
    aoi22 ix9452 (.Y (nx9451), .A0 (que_out_24__0__9), .A1 (nx10058), .B0 (
          que_out_22__0__9), .B1 (nx10032)) ;
    nand03 ix8215 (.Y (nx8214), .A0 (nx9454), .A1 (nx9456), .A2 (nx9458)) ;
    aoi222 ix9455 (.Y (nx9454), .A0 (que_out_15__0__9), .A1 (nx9980), .B0 (
           que_out_3__0__9), .B1 (nx10006), .C0 (que_out_23__0__9), .C1 (nx9954)
           ) ;
    aoi22 ix9457 (.Y (nx9456), .A0 (que_out_27__0__9), .A1 (nx9928), .B0 (
          que_out_4__0__9), .B1 (nx9902)) ;
    aoi22 ix9459 (.Y (nx9458), .A0 (que_out_0__0__9), .A1 (nx9850), .B0 (
          que_out_2__0__9), .B1 (nx9876)) ;
    nand03 ix8189 (.Y (nx8188), .A0 (nx9461), .A1 (nx9463), .A2 (nx9465)) ;
    aoi222 ix9462 (.Y (nx9461), .A0 (que_out_26__0__9), .A1 (nx9824), .B0 (
           que_out_14__0__9), .B1 (nx9798), .C0 (que_out_11__0__9), .C1 (nx9772)
           ) ;
    aoi22 ix9464 (.Y (nx9463), .A0 (que_out_13__0__9), .A1 (nx9746), .B0 (
          que_out_7__0__9), .B1 (nx9720)) ;
    aoi22 ix9466 (.Y (nx9465), .A0 (que_out_12__0__9), .A1 (nx9694), .B0 (
          que_out_1__0__9), .B1 (nx9668)) ;
    or04 ix8383 (.Y (out_column_0__10), .A0 (nx8378), .A1 (nx8352), .A2 (nx8324)
         , .A3 (nx8298)) ;
    nand03 ix8379 (.Y (nx8378), .A0 (nx9469), .A1 (nx9471), .A2 (nx9473)) ;
    aoi222 ix9470 (.Y (nx9469), .A0 (que_out_10__0__10), .A1 (nx10318), .B0 (
           que_out_6__0__10), .B1 (nx10370), .C0 (que_out_9__0__10), .C1 (
           nx10344)) ;
    aoi22 ix9472 (.Y (nx9471), .A0 (que_out_5__0__10), .A1 (nx10266), .B0 (
          que_out_18__0__10), .B1 (nx10292)) ;
    aoi22 ix9474 (.Y (nx9473), .A0 (que_out_17__0__10), .A1 (nx10240), .B0 (
          que_out_20__0__10), .B1 (nx10214)) ;
    nand03 ix8353 (.Y (nx8352), .A0 (nx9476), .A1 (nx9478), .A2 (nx9480)) ;
    aoi222 ix9477 (.Y (nx9476), .A0 (que_out_19__0__10), .A1 (nx10188), .B0 (
           que_out_21__0__10), .B1 (nx10162), .C0 (que_out_8__0__10), .C1 (
           nx10136)) ;
    aoi22 ix9479 (.Y (nx9478), .A0 (que_out_25__0__10), .A1 (nx10084), .B0 (
          que_out_16__0__10), .B1 (nx10110)) ;
    aoi22 ix9481 (.Y (nx9480), .A0 (que_out_24__0__10), .A1 (nx10058), .B0 (
          que_out_22__0__10), .B1 (nx10032)) ;
    nand03 ix8325 (.Y (nx8324), .A0 (nx9483), .A1 (nx9485), .A2 (nx9487)) ;
    aoi222 ix9484 (.Y (nx9483), .A0 (que_out_15__0__10), .A1 (nx9980), .B0 (
           que_out_3__0__10), .B1 (nx10006), .C0 (que_out_23__0__10), .C1 (
           nx9954)) ;
    aoi22 ix9486 (.Y (nx9485), .A0 (que_out_27__0__10), .A1 (nx9928), .B0 (
          que_out_4__0__10), .B1 (nx9902)) ;
    aoi22 ix9488 (.Y (nx9487), .A0 (que_out_0__0__10), .A1 (nx9850), .B0 (
          que_out_2__0__10), .B1 (nx9876)) ;
    nand03 ix8299 (.Y (nx8298), .A0 (nx9490), .A1 (nx9492), .A2 (nx9494)) ;
    aoi222 ix9491 (.Y (nx9490), .A0 (que_out_26__0__10), .A1 (nx9824), .B0 (
           que_out_14__0__10), .B1 (nx9798), .C0 (que_out_11__0__10), .C1 (
           nx9772)) ;
    aoi22 ix9493 (.Y (nx9492), .A0 (que_out_13__0__10), .A1 (nx9746), .B0 (
          que_out_7__0__10), .B1 (nx9720)) ;
    aoi22 ix9495 (.Y (nx9494), .A0 (que_out_12__0__10), .A1 (nx9694), .B0 (
          que_out_1__0__10), .B1 (nx9668)) ;
    or04 ix8493 (.Y (out_column_0__11), .A0 (nx8488), .A1 (nx8462), .A2 (nx8434)
         , .A3 (nx8408)) ;
    nand03 ix8489 (.Y (nx8488), .A0 (nx9498), .A1 (nx9500), .A2 (nx9502)) ;
    aoi222 ix9499 (.Y (nx9498), .A0 (que_out_10__0__11), .A1 (nx10318), .B0 (
           que_out_6__0__11), .B1 (nx10370), .C0 (que_out_9__0__11), .C1 (
           nx10344)) ;
    aoi22 ix9501 (.Y (nx9500), .A0 (que_out_5__0__11), .A1 (nx10266), .B0 (
          que_out_18__0__11), .B1 (nx10292)) ;
    aoi22 ix9503 (.Y (nx9502), .A0 (que_out_17__0__11), .A1 (nx10240), .B0 (
          que_out_20__0__11), .B1 (nx10214)) ;
    nand03 ix8463 (.Y (nx8462), .A0 (nx9505), .A1 (nx9507), .A2 (nx9509)) ;
    aoi222 ix9506 (.Y (nx9505), .A0 (que_out_19__0__11), .A1 (nx10188), .B0 (
           que_out_21__0__11), .B1 (nx10162), .C0 (que_out_8__0__11), .C1 (
           nx10136)) ;
    aoi22 ix9508 (.Y (nx9507), .A0 (que_out_25__0__11), .A1 (nx10084), .B0 (
          que_out_16__0__11), .B1 (nx10110)) ;
    aoi22 ix9510 (.Y (nx9509), .A0 (que_out_24__0__11), .A1 (nx10058), .B0 (
          que_out_22__0__11), .B1 (nx10032)) ;
    nand03 ix8435 (.Y (nx8434), .A0 (nx9512), .A1 (nx9514), .A2 (nx9516)) ;
    aoi222 ix9513 (.Y (nx9512), .A0 (que_out_15__0__11), .A1 (nx9980), .B0 (
           que_out_3__0__11), .B1 (nx10006), .C0 (que_out_23__0__11), .C1 (
           nx9954)) ;
    aoi22 ix9515 (.Y (nx9514), .A0 (que_out_27__0__11), .A1 (nx9928), .B0 (
          que_out_4__0__11), .B1 (nx9902)) ;
    aoi22 ix9517 (.Y (nx9516), .A0 (que_out_0__0__11), .A1 (nx9850), .B0 (
          que_out_2__0__11), .B1 (nx9876)) ;
    nand03 ix8409 (.Y (nx8408), .A0 (nx9519), .A1 (nx9521), .A2 (nx9523)) ;
    aoi222 ix9520 (.Y (nx9519), .A0 (que_out_26__0__11), .A1 (nx9824), .B0 (
           que_out_14__0__11), .B1 (nx9798), .C0 (que_out_11__0__11), .C1 (
           nx9772)) ;
    aoi22 ix9522 (.Y (nx9521), .A0 (que_out_13__0__11), .A1 (nx9746), .B0 (
          que_out_7__0__11), .B1 (nx9720)) ;
    aoi22 ix9524 (.Y (nx9523), .A0 (que_out_12__0__11), .A1 (nx9694), .B0 (
          que_out_1__0__11), .B1 (nx9668)) ;
    or04 ix8603 (.Y (out_column_0__12), .A0 (nx8598), .A1 (nx8572), .A2 (nx8544)
         , .A3 (nx8518)) ;
    nand03 ix8599 (.Y (nx8598), .A0 (nx9527), .A1 (nx9529), .A2 (nx9531)) ;
    aoi222 ix9528 (.Y (nx9527), .A0 (que_out_10__0__12), .A1 (nx10318), .B0 (
           que_out_6__0__12), .B1 (nx10370), .C0 (que_out_9__0__12), .C1 (
           nx10344)) ;
    aoi22 ix9530 (.Y (nx9529), .A0 (que_out_5__0__12), .A1 (nx10266), .B0 (
          que_out_18__0__12), .B1 (nx10292)) ;
    aoi22 ix9532 (.Y (nx9531), .A0 (que_out_17__0__12), .A1 (nx10240), .B0 (
          que_out_20__0__12), .B1 (nx10214)) ;
    nand03 ix8573 (.Y (nx8572), .A0 (nx9534), .A1 (nx9536), .A2 (nx9538)) ;
    aoi222 ix9535 (.Y (nx9534), .A0 (que_out_19__0__12), .A1 (nx10188), .B0 (
           que_out_21__0__12), .B1 (nx10162), .C0 (que_out_8__0__12), .C1 (
           nx10136)) ;
    aoi22 ix9537 (.Y (nx9536), .A0 (que_out_25__0__12), .A1 (nx10084), .B0 (
          que_out_16__0__12), .B1 (nx10110)) ;
    aoi22 ix9539 (.Y (nx9538), .A0 (que_out_24__0__12), .A1 (nx10058), .B0 (
          que_out_22__0__12), .B1 (nx10032)) ;
    nand03 ix8545 (.Y (nx8544), .A0 (nx9541), .A1 (nx9543), .A2 (nx9545)) ;
    aoi222 ix9542 (.Y (nx9541), .A0 (que_out_15__0__12), .A1 (nx9980), .B0 (
           que_out_3__0__12), .B1 (nx10006), .C0 (que_out_23__0__12), .C1 (
           nx9954)) ;
    aoi22 ix9544 (.Y (nx9543), .A0 (que_out_27__0__12), .A1 (nx9928), .B0 (
          que_out_4__0__12), .B1 (nx9902)) ;
    aoi22 ix9546 (.Y (nx9545), .A0 (que_out_0__0__12), .A1 (nx9850), .B0 (
          que_out_2__0__12), .B1 (nx9876)) ;
    nand03 ix8519 (.Y (nx8518), .A0 (nx9548), .A1 (nx9550), .A2 (nx9552)) ;
    aoi222 ix9549 (.Y (nx9548), .A0 (que_out_26__0__12), .A1 (nx9824), .B0 (
           que_out_14__0__12), .B1 (nx9798), .C0 (que_out_11__0__12), .C1 (
           nx9772)) ;
    aoi22 ix9551 (.Y (nx9550), .A0 (que_out_13__0__12), .A1 (nx9746), .B0 (
          que_out_7__0__12), .B1 (nx9720)) ;
    aoi22 ix9553 (.Y (nx9552), .A0 (que_out_12__0__12), .A1 (nx9694), .B0 (
          que_out_1__0__12), .B1 (nx9668)) ;
    or04 ix8713 (.Y (out_column_0__13), .A0 (nx8708), .A1 (nx8682), .A2 (nx8654)
         , .A3 (nx8628)) ;
    nand03 ix8709 (.Y (nx8708), .A0 (nx9556), .A1 (nx9558), .A2 (nx9560)) ;
    aoi222 ix9557 (.Y (nx9556), .A0 (que_out_10__0__13), .A1 (nx10320), .B0 (
           que_out_6__0__13), .B1 (nx10372), .C0 (que_out_9__0__13), .C1 (
           nx10346)) ;
    aoi22 ix9559 (.Y (nx9558), .A0 (que_out_5__0__13), .A1 (nx10268), .B0 (
          que_out_18__0__13), .B1 (nx10294)) ;
    aoi22 ix9561 (.Y (nx9560), .A0 (que_out_17__0__13), .A1 (nx10242), .B0 (
          que_out_20__0__13), .B1 (nx10216)) ;
    nand03 ix8683 (.Y (nx8682), .A0 (nx9563), .A1 (nx9565), .A2 (nx9567)) ;
    aoi222 ix9564 (.Y (nx9563), .A0 (que_out_19__0__13), .A1 (nx10190), .B0 (
           que_out_21__0__13), .B1 (nx10164), .C0 (que_out_8__0__13), .C1 (
           nx10138)) ;
    aoi22 ix9566 (.Y (nx9565), .A0 (que_out_25__0__13), .A1 (nx10086), .B0 (
          que_out_16__0__13), .B1 (nx10112)) ;
    aoi22 ix9568 (.Y (nx9567), .A0 (que_out_24__0__13), .A1 (nx10060), .B0 (
          que_out_22__0__13), .B1 (nx10034)) ;
    nand03 ix8655 (.Y (nx8654), .A0 (nx9570), .A1 (nx9572), .A2 (nx9574)) ;
    aoi222 ix9571 (.Y (nx9570), .A0 (que_out_15__0__13), .A1 (nx9982), .B0 (
           que_out_3__0__13), .B1 (nx10008), .C0 (que_out_23__0__13), .C1 (
           nx9956)) ;
    aoi22 ix9573 (.Y (nx9572), .A0 (que_out_27__0__13), .A1 (nx9930), .B0 (
          que_out_4__0__13), .B1 (nx9904)) ;
    aoi22 ix9575 (.Y (nx9574), .A0 (que_out_0__0__13), .A1 (nx9852), .B0 (
          que_out_2__0__13), .B1 (nx9878)) ;
    nand03 ix8629 (.Y (nx8628), .A0 (nx9577), .A1 (nx9579), .A2 (nx9581)) ;
    aoi222 ix9578 (.Y (nx9577), .A0 (que_out_26__0__13), .A1 (nx9826), .B0 (
           que_out_14__0__13), .B1 (nx9800), .C0 (que_out_11__0__13), .C1 (
           nx9774)) ;
    aoi22 ix9580 (.Y (nx9579), .A0 (que_out_13__0__13), .A1 (nx9748), .B0 (
          que_out_7__0__13), .B1 (nx9722)) ;
    aoi22 ix9582 (.Y (nx9581), .A0 (que_out_12__0__13), .A1 (nx9696), .B0 (
          que_out_1__0__13), .B1 (nx9670)) ;
    or04 ix8823 (.Y (out_column_0__14), .A0 (nx8818), .A1 (nx8792), .A2 (nx8764)
         , .A3 (nx8738)) ;
    nand03 ix8819 (.Y (nx8818), .A0 (nx9585), .A1 (nx9587), .A2 (nx9589)) ;
    aoi222 ix9586 (.Y (nx9585), .A0 (que_out_10__0__14), .A1 (nx10320), .B0 (
           que_out_6__0__14), .B1 (nx10372), .C0 (que_out_9__0__14), .C1 (
           nx10346)) ;
    aoi22 ix9588 (.Y (nx9587), .A0 (que_out_5__0__14), .A1 (nx10268), .B0 (
          que_out_18__0__14), .B1 (nx10294)) ;
    aoi22 ix9590 (.Y (nx9589), .A0 (que_out_17__0__14), .A1 (nx10242), .B0 (
          que_out_20__0__14), .B1 (nx10216)) ;
    nand03 ix8793 (.Y (nx8792), .A0 (nx9592), .A1 (nx9594), .A2 (nx9596)) ;
    aoi222 ix9593 (.Y (nx9592), .A0 (que_out_19__0__14), .A1 (nx10190), .B0 (
           que_out_21__0__14), .B1 (nx10164), .C0 (que_out_8__0__14), .C1 (
           nx10138)) ;
    aoi22 ix9595 (.Y (nx9594), .A0 (que_out_25__0__14), .A1 (nx10086), .B0 (
          que_out_16__0__14), .B1 (nx10112)) ;
    aoi22 ix9597 (.Y (nx9596), .A0 (que_out_24__0__14), .A1 (nx10060), .B0 (
          que_out_22__0__14), .B1 (nx10034)) ;
    nand03 ix8765 (.Y (nx8764), .A0 (nx9599), .A1 (nx9601), .A2 (nx9603)) ;
    aoi222 ix9600 (.Y (nx9599), .A0 (que_out_15__0__14), .A1 (nx9982), .B0 (
           que_out_3__0__14), .B1 (nx10008), .C0 (que_out_23__0__14), .C1 (
           nx9956)) ;
    aoi22 ix9602 (.Y (nx9601), .A0 (que_out_27__0__14), .A1 (nx9930), .B0 (
          que_out_4__0__14), .B1 (nx9904)) ;
    aoi22 ix9604 (.Y (nx9603), .A0 (que_out_0__0__14), .A1 (nx9852), .B0 (
          que_out_2__0__14), .B1 (nx9878)) ;
    nand03 ix8739 (.Y (nx8738), .A0 (nx9606), .A1 (nx9608), .A2 (nx9610)) ;
    aoi222 ix9607 (.Y (nx9606), .A0 (que_out_26__0__14), .A1 (nx9826), .B0 (
           que_out_14__0__14), .B1 (nx9800), .C0 (que_out_11__0__14), .C1 (
           nx9774)) ;
    aoi22 ix9609 (.Y (nx9608), .A0 (que_out_13__0__14), .A1 (nx9748), .B0 (
          que_out_7__0__14), .B1 (nx9722)) ;
    aoi22 ix9611 (.Y (nx9610), .A0 (que_out_12__0__14), .A1 (nx9696), .B0 (
          que_out_1__0__14), .B1 (nx9670)) ;
    or04 ix8933 (.Y (out_column_0__15), .A0 (nx8928), .A1 (nx8902), .A2 (nx8874)
         , .A3 (nx8848)) ;
    nand03 ix8929 (.Y (nx8928), .A0 (nx9614), .A1 (nx9616), .A2 (nx9618)) ;
    aoi222 ix9615 (.Y (nx9614), .A0 (que_out_10__0__15), .A1 (nx10320), .B0 (
           que_out_6__0__15), .B1 (nx10372), .C0 (que_out_9__0__15), .C1 (
           nx10346)) ;
    aoi22 ix9617 (.Y (nx9616), .A0 (que_out_5__0__15), .A1 (nx10268), .B0 (
          que_out_18__0__15), .B1 (nx10294)) ;
    aoi22 ix9619 (.Y (nx9618), .A0 (que_out_17__0__15), .A1 (nx10242), .B0 (
          que_out_20__0__15), .B1 (nx10216)) ;
    nand03 ix8903 (.Y (nx8902), .A0 (nx9621), .A1 (nx9623), .A2 (nx9625)) ;
    aoi222 ix9622 (.Y (nx9621), .A0 (que_out_19__0__15), .A1 (nx10190), .B0 (
           que_out_21__0__15), .B1 (nx10164), .C0 (que_out_8__0__15), .C1 (
           nx10138)) ;
    aoi22 ix9624 (.Y (nx9623), .A0 (que_out_25__0__15), .A1 (nx10086), .B0 (
          que_out_16__0__15), .B1 (nx10112)) ;
    aoi22 ix9626 (.Y (nx9625), .A0 (que_out_24__0__15), .A1 (nx10060), .B0 (
          que_out_22__0__15), .B1 (nx10034)) ;
    nand03 ix8875 (.Y (nx8874), .A0 (nx9628), .A1 (nx9630), .A2 (nx9632)) ;
    aoi222 ix9629 (.Y (nx9628), .A0 (que_out_15__0__15), .A1 (nx9982), .B0 (
           que_out_3__0__15), .B1 (nx10008), .C0 (que_out_23__0__15), .C1 (
           nx9956)) ;
    aoi22 ix9631 (.Y (nx9630), .A0 (que_out_27__0__15), .A1 (nx9930), .B0 (
          que_out_4__0__15), .B1 (nx9904)) ;
    aoi22 ix9633 (.Y (nx9632), .A0 (que_out_0__0__15), .A1 (nx9852), .B0 (
          que_out_2__0__15), .B1 (nx9878)) ;
    nand03 ix8849 (.Y (nx8848), .A0 (nx9635), .A1 (nx9637), .A2 (nx9639)) ;
    aoi222 ix9636 (.Y (nx9635), .A0 (que_out_26__0__15), .A1 (nx9826), .B0 (
           que_out_14__0__15), .B1 (nx9800), .C0 (que_out_11__0__15), .C1 (
           nx9774)) ;
    aoi22 ix9638 (.Y (nx9637), .A0 (que_out_13__0__15), .A1 (nx9748), .B0 (
          que_out_7__0__15), .B1 (nx9722)) ;
    aoi22 ix9640 (.Y (nx9639), .A0 (que_out_12__0__15), .A1 (nx9696), .B0 (
          que_out_1__0__15), .B1 (nx9670)) ;
    inv02 ix6944 (.Y (nx6943), .A (nx88)) ;
    inv02 ix9647 (.Y (nx9648), .A (nx10378)) ;
    inv02 ix9649 (.Y (nx9650), .A (nx10378)) ;
    inv02 ix9651 (.Y (nx9652), .A (nx10378)) ;
    inv02 ix9653 (.Y (nx9654), .A (nx10378)) ;
    inv02 ix9655 (.Y (nx9656), .A (nx10378)) ;
    inv02 ix9657 (.Y (nx9658), .A (nx10378)) ;
    inv02 ix9659 (.Y (nx9660), .A (nx10378)) ;
    inv02 ix9661 (.Y (nx9662), .A (nx10380)) ;
    inv02 ix9663 (.Y (nx9664), .A (nx10380)) ;
    inv02 ix9665 (.Y (nx9666), .A (nx10380)) ;
    inv02 ix9667 (.Y (nx9668), .A (nx10380)) ;
    inv02 ix9669 (.Y (nx9670), .A (nx10380)) ;
    inv02 ix9673 (.Y (nx9674), .A (nx10382)) ;
    inv02 ix9675 (.Y (nx9676), .A (nx10382)) ;
    inv02 ix9677 (.Y (nx9678), .A (nx10382)) ;
    inv02 ix9679 (.Y (nx9680), .A (nx10382)) ;
    inv02 ix9681 (.Y (nx9682), .A (nx10382)) ;
    inv02 ix9683 (.Y (nx9684), .A (nx10382)) ;
    inv02 ix9685 (.Y (nx9686), .A (nx10382)) ;
    inv02 ix9687 (.Y (nx9688), .A (nx10384)) ;
    inv02 ix9689 (.Y (nx9690), .A (nx10384)) ;
    inv02 ix9691 (.Y (nx9692), .A (nx10384)) ;
    inv02 ix9693 (.Y (nx9694), .A (nx10384)) ;
    inv02 ix9695 (.Y (nx9696), .A (nx10384)) ;
    inv02 ix9699 (.Y (nx9700), .A (nx10386)) ;
    inv02 ix9701 (.Y (nx9702), .A (nx10386)) ;
    inv02 ix9703 (.Y (nx9704), .A (nx10386)) ;
    inv02 ix9705 (.Y (nx9706), .A (nx10386)) ;
    inv02 ix9707 (.Y (nx9708), .A (nx10386)) ;
    inv02 ix9709 (.Y (nx9710), .A (nx10386)) ;
    inv02 ix9711 (.Y (nx9712), .A (nx10386)) ;
    inv02 ix9713 (.Y (nx9714), .A (nx10388)) ;
    inv02 ix9715 (.Y (nx9716), .A (nx10388)) ;
    inv02 ix9717 (.Y (nx9718), .A (nx10388)) ;
    inv02 ix9719 (.Y (nx9720), .A (nx10388)) ;
    inv02 ix9721 (.Y (nx9722), .A (nx10388)) ;
    inv02 ix9725 (.Y (nx9726), .A (nx10390)) ;
    inv02 ix9727 (.Y (nx9728), .A (nx10390)) ;
    inv02 ix9729 (.Y (nx9730), .A (nx10390)) ;
    inv02 ix9731 (.Y (nx9732), .A (nx10390)) ;
    inv02 ix9733 (.Y (nx9734), .A (nx10390)) ;
    inv02 ix9735 (.Y (nx9736), .A (nx10390)) ;
    inv02 ix9737 (.Y (nx9738), .A (nx10390)) ;
    inv02 ix9739 (.Y (nx9740), .A (nx10392)) ;
    inv02 ix9741 (.Y (nx9742), .A (nx10392)) ;
    inv02 ix9743 (.Y (nx9744), .A (nx10392)) ;
    inv02 ix9745 (.Y (nx9746), .A (nx10392)) ;
    inv02 ix9747 (.Y (nx9748), .A (nx10392)) ;
    inv02 ix9751 (.Y (nx9752), .A (nx10394)) ;
    inv02 ix9753 (.Y (nx9754), .A (nx10394)) ;
    inv02 ix9755 (.Y (nx9756), .A (nx10394)) ;
    inv02 ix9757 (.Y (nx9758), .A (nx10394)) ;
    inv02 ix9759 (.Y (nx9760), .A (nx10394)) ;
    inv02 ix9761 (.Y (nx9762), .A (nx10394)) ;
    inv02 ix9763 (.Y (nx9764), .A (nx10394)) ;
    inv02 ix9765 (.Y (nx9766), .A (nx10396)) ;
    inv02 ix9767 (.Y (nx9768), .A (nx10396)) ;
    inv02 ix9769 (.Y (nx9770), .A (nx10396)) ;
    inv02 ix9771 (.Y (nx9772), .A (nx10396)) ;
    inv02 ix9773 (.Y (nx9774), .A (nx10396)) ;
    inv02 ix9777 (.Y (nx9778), .A (nx10398)) ;
    inv02 ix9779 (.Y (nx9780), .A (nx10398)) ;
    inv02 ix9781 (.Y (nx9782), .A (nx10398)) ;
    inv02 ix9783 (.Y (nx9784), .A (nx10398)) ;
    inv02 ix9785 (.Y (nx9786), .A (nx10398)) ;
    inv02 ix9787 (.Y (nx9788), .A (nx10398)) ;
    inv02 ix9789 (.Y (nx9790), .A (nx10398)) ;
    inv02 ix9791 (.Y (nx9792), .A (nx10400)) ;
    inv02 ix9793 (.Y (nx9794), .A (nx10400)) ;
    inv02 ix9795 (.Y (nx9796), .A (nx10400)) ;
    inv02 ix9797 (.Y (nx9798), .A (nx10400)) ;
    inv02 ix9799 (.Y (nx9800), .A (nx10400)) ;
    inv02 ix9803 (.Y (nx9804), .A (nx10402)) ;
    inv02 ix9805 (.Y (nx9806), .A (nx10402)) ;
    inv02 ix9807 (.Y (nx9808), .A (nx10402)) ;
    inv02 ix9809 (.Y (nx9810), .A (nx10402)) ;
    inv02 ix9811 (.Y (nx9812), .A (nx10402)) ;
    inv02 ix9813 (.Y (nx9814), .A (nx10402)) ;
    inv02 ix9815 (.Y (nx9816), .A (nx10402)) ;
    inv02 ix9817 (.Y (nx9818), .A (nx10404)) ;
    inv02 ix9819 (.Y (nx9820), .A (nx10404)) ;
    inv02 ix9821 (.Y (nx9822), .A (nx10404)) ;
    inv02 ix9823 (.Y (nx9824), .A (nx10404)) ;
    inv02 ix9825 (.Y (nx9826), .A (nx10404)) ;
    inv02 ix9829 (.Y (nx9830), .A (nx10406)) ;
    inv02 ix9831 (.Y (nx9832), .A (nx10406)) ;
    inv02 ix9833 (.Y (nx9834), .A (nx10406)) ;
    inv02 ix9835 (.Y (nx9836), .A (nx10406)) ;
    inv02 ix9837 (.Y (nx9838), .A (nx10406)) ;
    inv02 ix9839 (.Y (nx9840), .A (nx10406)) ;
    inv02 ix9841 (.Y (nx9842), .A (nx10406)) ;
    inv02 ix9843 (.Y (nx9844), .A (nx10408)) ;
    inv02 ix9845 (.Y (nx9846), .A (nx10408)) ;
    inv02 ix9847 (.Y (nx9848), .A (nx10408)) ;
    inv02 ix9849 (.Y (nx9850), .A (nx10408)) ;
    inv02 ix9851 (.Y (nx9852), .A (nx10408)) ;
    inv02 ix9855 (.Y (nx9856), .A (nx10410)) ;
    inv02 ix9857 (.Y (nx9858), .A (nx10410)) ;
    inv02 ix9859 (.Y (nx9860), .A (nx10410)) ;
    inv02 ix9861 (.Y (nx9862), .A (nx10410)) ;
    inv02 ix9863 (.Y (nx9864), .A (nx10410)) ;
    inv02 ix9865 (.Y (nx9866), .A (nx10410)) ;
    inv02 ix9867 (.Y (nx9868), .A (nx10410)) ;
    inv02 ix9869 (.Y (nx9870), .A (nx10412)) ;
    inv02 ix9871 (.Y (nx9872), .A (nx10412)) ;
    inv02 ix9873 (.Y (nx9874), .A (nx10412)) ;
    inv02 ix9875 (.Y (nx9876), .A (nx10412)) ;
    inv02 ix9877 (.Y (nx9878), .A (nx10412)) ;
    inv02 ix9881 (.Y (nx9882), .A (nx10414)) ;
    inv02 ix9883 (.Y (nx9884), .A (nx10414)) ;
    inv02 ix9885 (.Y (nx9886), .A (nx10414)) ;
    inv02 ix9887 (.Y (nx9888), .A (nx10414)) ;
    inv02 ix9889 (.Y (nx9890), .A (nx10414)) ;
    inv02 ix9891 (.Y (nx9892), .A (nx10414)) ;
    inv02 ix9893 (.Y (nx9894), .A (nx10414)) ;
    inv02 ix9895 (.Y (nx9896), .A (nx10416)) ;
    inv02 ix9897 (.Y (nx9898), .A (nx10416)) ;
    inv02 ix9899 (.Y (nx9900), .A (nx10416)) ;
    inv02 ix9901 (.Y (nx9902), .A (nx10416)) ;
    inv02 ix9903 (.Y (nx9904), .A (nx10416)) ;
    inv02 ix9907 (.Y (nx9908), .A (nx10418)) ;
    inv02 ix9909 (.Y (nx9910), .A (nx10418)) ;
    inv02 ix9911 (.Y (nx9912), .A (nx10418)) ;
    inv02 ix9913 (.Y (nx9914), .A (nx10418)) ;
    inv02 ix9915 (.Y (nx9916), .A (nx10418)) ;
    inv02 ix9917 (.Y (nx9918), .A (nx10418)) ;
    inv02 ix9919 (.Y (nx9920), .A (nx10418)) ;
    inv02 ix9921 (.Y (nx9922), .A (nx10420)) ;
    inv02 ix9923 (.Y (nx9924), .A (nx10420)) ;
    inv02 ix9925 (.Y (nx9926), .A (nx10420)) ;
    inv02 ix9927 (.Y (nx9928), .A (nx10420)) ;
    inv02 ix9929 (.Y (nx9930), .A (nx10420)) ;
    inv02 ix9933 (.Y (nx9934), .A (nx10422)) ;
    inv02 ix9935 (.Y (nx9936), .A (nx10422)) ;
    inv02 ix9937 (.Y (nx9938), .A (nx10422)) ;
    inv02 ix9939 (.Y (nx9940), .A (nx10422)) ;
    inv02 ix9941 (.Y (nx9942), .A (nx10422)) ;
    inv02 ix9943 (.Y (nx9944), .A (nx10422)) ;
    inv02 ix9945 (.Y (nx9946), .A (nx10422)) ;
    inv02 ix9947 (.Y (nx9948), .A (nx10424)) ;
    inv02 ix9949 (.Y (nx9950), .A (nx10424)) ;
    inv02 ix9951 (.Y (nx9952), .A (nx10424)) ;
    inv02 ix9953 (.Y (nx9954), .A (nx10424)) ;
    inv02 ix9955 (.Y (nx9956), .A (nx10424)) ;
    inv02 ix9959 (.Y (nx9960), .A (nx10426)) ;
    inv02 ix9961 (.Y (nx9962), .A (nx10426)) ;
    inv02 ix9963 (.Y (nx9964), .A (nx10426)) ;
    inv02 ix9965 (.Y (nx9966), .A (nx10426)) ;
    inv02 ix9967 (.Y (nx9968), .A (nx10426)) ;
    inv02 ix9969 (.Y (nx9970), .A (nx10426)) ;
    inv02 ix9971 (.Y (nx9972), .A (nx10426)) ;
    inv02 ix9973 (.Y (nx9974), .A (nx10428)) ;
    inv02 ix9975 (.Y (nx9976), .A (nx10428)) ;
    inv02 ix9977 (.Y (nx9978), .A (nx10428)) ;
    inv02 ix9979 (.Y (nx9980), .A (nx10428)) ;
    inv02 ix9981 (.Y (nx9982), .A (nx10428)) ;
    inv02 ix9985 (.Y (nx9986), .A (nx10430)) ;
    inv02 ix9987 (.Y (nx9988), .A (nx10430)) ;
    inv02 ix9989 (.Y (nx9990), .A (nx10430)) ;
    inv02 ix9991 (.Y (nx9992), .A (nx10430)) ;
    inv02 ix9993 (.Y (nx9994), .A (nx10430)) ;
    inv02 ix9995 (.Y (nx9996), .A (nx10430)) ;
    inv02 ix9997 (.Y (nx9998), .A (nx10430)) ;
    inv02 ix9999 (.Y (nx10000), .A (nx10432)) ;
    inv02 ix10001 (.Y (nx10002), .A (nx10432)) ;
    inv02 ix10003 (.Y (nx10004), .A (nx10432)) ;
    inv02 ix10005 (.Y (nx10006), .A (nx10432)) ;
    inv02 ix10007 (.Y (nx10008), .A (nx10432)) ;
    inv02 ix10011 (.Y (nx10012), .A (nx10434)) ;
    inv02 ix10013 (.Y (nx10014), .A (nx10434)) ;
    inv02 ix10015 (.Y (nx10016), .A (nx10434)) ;
    inv02 ix10017 (.Y (nx10018), .A (nx10434)) ;
    inv02 ix10019 (.Y (nx10020), .A (nx10434)) ;
    inv02 ix10021 (.Y (nx10022), .A (nx10434)) ;
    inv02 ix10023 (.Y (nx10024), .A (nx10434)) ;
    inv02 ix10025 (.Y (nx10026), .A (nx10436)) ;
    inv02 ix10027 (.Y (nx10028), .A (nx10436)) ;
    inv02 ix10029 (.Y (nx10030), .A (nx10436)) ;
    inv02 ix10031 (.Y (nx10032), .A (nx10436)) ;
    inv02 ix10033 (.Y (nx10034), .A (nx10436)) ;
    inv02 ix10037 (.Y (nx10038), .A (nx10438)) ;
    inv02 ix10039 (.Y (nx10040), .A (nx10438)) ;
    inv02 ix10041 (.Y (nx10042), .A (nx10438)) ;
    inv02 ix10043 (.Y (nx10044), .A (nx10438)) ;
    inv02 ix10045 (.Y (nx10046), .A (nx10438)) ;
    inv02 ix10047 (.Y (nx10048), .A (nx10438)) ;
    inv02 ix10049 (.Y (nx10050), .A (nx10438)) ;
    inv02 ix10051 (.Y (nx10052), .A (nx10440)) ;
    inv02 ix10053 (.Y (nx10054), .A (nx10440)) ;
    inv02 ix10055 (.Y (nx10056), .A (nx10440)) ;
    inv02 ix10057 (.Y (nx10058), .A (nx10440)) ;
    inv02 ix10059 (.Y (nx10060), .A (nx10440)) ;
    inv02 ix10063 (.Y (nx10064), .A (nx10442)) ;
    inv02 ix10065 (.Y (nx10066), .A (nx10442)) ;
    inv02 ix10067 (.Y (nx10068), .A (nx10442)) ;
    inv02 ix10069 (.Y (nx10070), .A (nx10442)) ;
    inv02 ix10071 (.Y (nx10072), .A (nx10442)) ;
    inv02 ix10073 (.Y (nx10074), .A (nx10442)) ;
    inv02 ix10075 (.Y (nx10076), .A (nx10442)) ;
    inv02 ix10077 (.Y (nx10078), .A (nx10444)) ;
    inv02 ix10079 (.Y (nx10080), .A (nx10444)) ;
    inv02 ix10081 (.Y (nx10082), .A (nx10444)) ;
    inv02 ix10083 (.Y (nx10084), .A (nx10444)) ;
    inv02 ix10085 (.Y (nx10086), .A (nx10444)) ;
    inv02 ix10089 (.Y (nx10090), .A (nx10446)) ;
    inv02 ix10091 (.Y (nx10092), .A (nx10446)) ;
    inv02 ix10093 (.Y (nx10094), .A (nx10446)) ;
    inv02 ix10095 (.Y (nx10096), .A (nx10446)) ;
    inv02 ix10097 (.Y (nx10098), .A (nx10446)) ;
    inv02 ix10099 (.Y (nx10100), .A (nx10446)) ;
    inv02 ix10101 (.Y (nx10102), .A (nx10446)) ;
    inv02 ix10103 (.Y (nx10104), .A (nx10448)) ;
    inv02 ix10105 (.Y (nx10106), .A (nx10448)) ;
    inv02 ix10107 (.Y (nx10108), .A (nx10448)) ;
    inv02 ix10109 (.Y (nx10110), .A (nx10448)) ;
    inv02 ix10111 (.Y (nx10112), .A (nx10448)) ;
    inv02 ix10115 (.Y (nx10116), .A (nx10450)) ;
    inv02 ix10117 (.Y (nx10118), .A (nx10450)) ;
    inv02 ix10119 (.Y (nx10120), .A (nx10450)) ;
    inv02 ix10121 (.Y (nx10122), .A (nx10450)) ;
    inv02 ix10123 (.Y (nx10124), .A (nx10450)) ;
    inv02 ix10125 (.Y (nx10126), .A (nx10450)) ;
    inv02 ix10127 (.Y (nx10128), .A (nx10450)) ;
    inv02 ix10129 (.Y (nx10130), .A (nx10452)) ;
    inv02 ix10131 (.Y (nx10132), .A (nx10452)) ;
    inv02 ix10133 (.Y (nx10134), .A (nx10452)) ;
    inv02 ix10135 (.Y (nx10136), .A (nx10452)) ;
    inv02 ix10137 (.Y (nx10138), .A (nx10452)) ;
    inv02 ix10141 (.Y (nx10142), .A (nx10454)) ;
    inv02 ix10143 (.Y (nx10144), .A (nx10454)) ;
    inv02 ix10145 (.Y (nx10146), .A (nx10454)) ;
    inv02 ix10147 (.Y (nx10148), .A (nx10454)) ;
    inv02 ix10149 (.Y (nx10150), .A (nx10454)) ;
    inv02 ix10151 (.Y (nx10152), .A (nx10454)) ;
    inv02 ix10153 (.Y (nx10154), .A (nx10454)) ;
    inv02 ix10155 (.Y (nx10156), .A (nx10456)) ;
    inv02 ix10157 (.Y (nx10158), .A (nx10456)) ;
    inv02 ix10159 (.Y (nx10160), .A (nx10456)) ;
    inv02 ix10161 (.Y (nx10162), .A (nx10456)) ;
    inv02 ix10163 (.Y (nx10164), .A (nx10456)) ;
    inv02 ix10167 (.Y (nx10168), .A (nx10458)) ;
    inv02 ix10169 (.Y (nx10170), .A (nx10458)) ;
    inv02 ix10171 (.Y (nx10172), .A (nx10458)) ;
    inv02 ix10173 (.Y (nx10174), .A (nx10458)) ;
    inv02 ix10175 (.Y (nx10176), .A (nx10458)) ;
    inv02 ix10177 (.Y (nx10178), .A (nx10458)) ;
    inv02 ix10179 (.Y (nx10180), .A (nx10458)) ;
    inv02 ix10181 (.Y (nx10182), .A (nx10460)) ;
    inv02 ix10183 (.Y (nx10184), .A (nx10460)) ;
    inv02 ix10185 (.Y (nx10186), .A (nx10460)) ;
    inv02 ix10187 (.Y (nx10188), .A (nx10460)) ;
    inv02 ix10189 (.Y (nx10190), .A (nx10460)) ;
    inv02 ix10193 (.Y (nx10194), .A (nx10462)) ;
    inv02 ix10195 (.Y (nx10196), .A (nx10462)) ;
    inv02 ix10197 (.Y (nx10198), .A (nx10462)) ;
    inv02 ix10199 (.Y (nx10200), .A (nx10462)) ;
    inv02 ix10201 (.Y (nx10202), .A (nx10462)) ;
    inv02 ix10203 (.Y (nx10204), .A (nx10462)) ;
    inv02 ix10205 (.Y (nx10206), .A (nx10462)) ;
    inv02 ix10207 (.Y (nx10208), .A (nx10464)) ;
    inv02 ix10209 (.Y (nx10210), .A (nx10464)) ;
    inv02 ix10211 (.Y (nx10212), .A (nx10464)) ;
    inv02 ix10213 (.Y (nx10214), .A (nx10464)) ;
    inv02 ix10215 (.Y (nx10216), .A (nx10464)) ;
    inv02 ix10219 (.Y (nx10220), .A (nx10466)) ;
    inv02 ix10221 (.Y (nx10222), .A (nx10466)) ;
    inv02 ix10223 (.Y (nx10224), .A (nx10466)) ;
    inv02 ix10225 (.Y (nx10226), .A (nx10466)) ;
    inv02 ix10227 (.Y (nx10228), .A (nx10466)) ;
    inv02 ix10229 (.Y (nx10230), .A (nx10466)) ;
    inv02 ix10231 (.Y (nx10232), .A (nx10466)) ;
    inv02 ix10233 (.Y (nx10234), .A (nx10468)) ;
    inv02 ix10235 (.Y (nx10236), .A (nx10468)) ;
    inv02 ix10237 (.Y (nx10238), .A (nx10468)) ;
    inv02 ix10239 (.Y (nx10240), .A (nx10468)) ;
    inv02 ix10241 (.Y (nx10242), .A (nx10468)) ;
    inv02 ix10245 (.Y (nx10246), .A (nx10470)) ;
    inv02 ix10247 (.Y (nx10248), .A (nx10470)) ;
    inv02 ix10249 (.Y (nx10250), .A (nx10470)) ;
    inv02 ix10251 (.Y (nx10252), .A (nx10470)) ;
    inv02 ix10253 (.Y (nx10254), .A (nx10470)) ;
    inv02 ix10255 (.Y (nx10256), .A (nx10470)) ;
    inv02 ix10257 (.Y (nx10258), .A (nx10470)) ;
    inv02 ix10259 (.Y (nx10260), .A (nx10472)) ;
    inv02 ix10261 (.Y (nx10262), .A (nx10472)) ;
    inv02 ix10263 (.Y (nx10264), .A (nx10472)) ;
    inv02 ix10265 (.Y (nx10266), .A (nx10472)) ;
    inv02 ix10267 (.Y (nx10268), .A (nx10472)) ;
    inv02 ix10271 (.Y (nx10272), .A (nx10474)) ;
    inv02 ix10273 (.Y (nx10274), .A (nx10474)) ;
    inv02 ix10275 (.Y (nx10276), .A (nx10474)) ;
    inv02 ix10277 (.Y (nx10278), .A (nx10474)) ;
    inv02 ix10279 (.Y (nx10280), .A (nx10474)) ;
    inv02 ix10281 (.Y (nx10282), .A (nx10474)) ;
    inv02 ix10283 (.Y (nx10284), .A (nx10474)) ;
    inv02 ix10285 (.Y (nx10286), .A (nx10476)) ;
    inv02 ix10287 (.Y (nx10288), .A (nx10476)) ;
    inv02 ix10289 (.Y (nx10290), .A (nx10476)) ;
    inv02 ix10291 (.Y (nx10292), .A (nx10476)) ;
    inv02 ix10293 (.Y (nx10294), .A (nx10476)) ;
    inv02 ix10297 (.Y (nx10298), .A (nx10478)) ;
    inv02 ix10299 (.Y (nx10300), .A (nx10478)) ;
    inv02 ix10301 (.Y (nx10302), .A (nx10478)) ;
    inv02 ix10303 (.Y (nx10304), .A (nx10478)) ;
    inv02 ix10305 (.Y (nx10306), .A (nx10478)) ;
    inv02 ix10307 (.Y (nx10308), .A (nx10478)) ;
    inv02 ix10309 (.Y (nx10310), .A (nx10478)) ;
    inv02 ix10311 (.Y (nx10312), .A (nx10480)) ;
    inv02 ix10313 (.Y (nx10314), .A (nx10480)) ;
    inv02 ix10315 (.Y (nx10316), .A (nx10480)) ;
    inv02 ix10317 (.Y (nx10318), .A (nx10480)) ;
    inv02 ix10319 (.Y (nx10320), .A (nx10480)) ;
    inv02 ix10323 (.Y (nx10324), .A (nx10482)) ;
    inv02 ix10325 (.Y (nx10326), .A (nx10482)) ;
    inv02 ix10327 (.Y (nx10328), .A (nx10482)) ;
    inv02 ix10329 (.Y (nx10330), .A (nx10482)) ;
    inv02 ix10331 (.Y (nx10332), .A (nx10482)) ;
    inv02 ix10333 (.Y (nx10334), .A (nx10482)) ;
    inv02 ix10335 (.Y (nx10336), .A (nx10482)) ;
    inv02 ix10337 (.Y (nx10338), .A (nx10484)) ;
    inv02 ix10339 (.Y (nx10340), .A (nx10484)) ;
    inv02 ix10341 (.Y (nx10342), .A (nx10484)) ;
    inv02 ix10343 (.Y (nx10344), .A (nx10484)) ;
    inv02 ix10345 (.Y (nx10346), .A (nx10484)) ;
    inv02 ix10349 (.Y (nx10350), .A (nx10486)) ;
    inv02 ix10351 (.Y (nx10352), .A (nx10486)) ;
    inv02 ix10353 (.Y (nx10354), .A (nx10486)) ;
    inv02 ix10355 (.Y (nx10356), .A (nx10486)) ;
    inv02 ix10357 (.Y (nx10358), .A (nx10486)) ;
    inv02 ix10359 (.Y (nx10360), .A (nx10486)) ;
    inv02 ix10361 (.Y (nx10362), .A (nx10486)) ;
    inv02 ix10363 (.Y (nx10364), .A (nx10488)) ;
    inv02 ix10365 (.Y (nx10366), .A (nx10488)) ;
    inv02 ix10367 (.Y (nx10368), .A (nx10488)) ;
    inv02 ix10369 (.Y (nx10370), .A (nx10488)) ;
    inv02 ix10371 (.Y (nx10372), .A (nx10488)) ;
    buf02 ix10373 (.Y (nx10374), .A (nx6955)) ;
    buf02 ix10375 (.Y (nx10376), .A (nx6955)) ;
    inv02 ix10377 (.Y (nx10378), .A (nx14)) ;
    inv02 ix10379 (.Y (nx10380), .A (nx14)) ;
    inv02 ix10381 (.Y (nx10382), .A (nx30)) ;
    inv02 ix10383 (.Y (nx10384), .A (nx30)) ;
    inv02 ix10385 (.Y (nx10386), .A (nx42)) ;
    inv02 ix10387 (.Y (nx10388), .A (nx42)) ;
    inv02 ix10389 (.Y (nx10390), .A (nx48)) ;
    inv02 ix10391 (.Y (nx10392), .A (nx48)) ;
    inv02 ix10393 (.Y (nx10394), .A (nx64)) ;
    inv02 ix10395 (.Y (nx10396), .A (nx64)) ;
    inv02 ix10397 (.Y (nx10398), .A (nx68)) ;
    inv02 ix10399 (.Y (nx10400), .A (nx68)) ;
    inv02 ix10401 (.Y (nx10402), .A (nx74)) ;
    inv02 ix10403 (.Y (nx10404), .A (nx74)) ;
    inv02 ix10405 (.Y (nx10406), .A (nx90)) ;
    inv02 ix10407 (.Y (nx10408), .A (nx90)) ;
    inv02 ix10409 (.Y (nx10410), .A (nx94)) ;
    inv02 ix10411 (.Y (nx10412), .A (nx94)) ;
    inv02 ix10413 (.Y (nx10414), .A (nx100)) ;
    inv02 ix10415 (.Y (nx10416), .A (nx100)) ;
    inv02 ix10417 (.Y (nx10418), .A (nx104)) ;
    inv02 ix10419 (.Y (nx10420), .A (nx104)) ;
    inv02 ix10421 (.Y (nx10422), .A (nx114)) ;
    inv02 ix10423 (.Y (nx10424), .A (nx114)) ;
    inv02 ix10425 (.Y (nx10426), .A (nx118)) ;
    inv02 ix10427 (.Y (nx10428), .A (nx118)) ;
    inv02 ix10429 (.Y (nx10430), .A (nx122)) ;
    inv02 ix10431 (.Y (nx10432), .A (nx122)) ;
    inv02 ix10433 (.Y (nx10434), .A (nx136)) ;
    inv02 ix10435 (.Y (nx10436), .A (nx136)) ;
    inv02 ix10437 (.Y (nx10438), .A (nx144)) ;
    inv02 ix10439 (.Y (nx10440), .A (nx144)) ;
    inv02 ix10441 (.Y (nx10442), .A (nx150)) ;
    inv02 ix10443 (.Y (nx10444), .A (nx150)) ;
    inv02 ix10445 (.Y (nx10446), .A (nx158)) ;
    inv02 ix10447 (.Y (nx10448), .A (nx158)) ;
    inv02 ix10449 (.Y (nx10450), .A (nx166)) ;
    inv02 ix10451 (.Y (nx10452), .A (nx166)) ;
    inv02 ix10453 (.Y (nx10454), .A (nx172)) ;
    inv02 ix10455 (.Y (nx10456), .A (nx172)) ;
    inv02 ix10457 (.Y (nx10458), .A (nx180)) ;
    inv02 ix10459 (.Y (nx10460), .A (nx180)) ;
    inv02 ix10461 (.Y (nx10462), .A (nx192)) ;
    inv02 ix10463 (.Y (nx10464), .A (nx192)) ;
    inv02 ix10465 (.Y (nx10466), .A (nx200)) ;
    inv02 ix10467 (.Y (nx10468), .A (nx200)) ;
    inv02 ix10469 (.Y (nx10470), .A (nx206)) ;
    inv02 ix10471 (.Y (nx10472), .A (nx206)) ;
    inv02 ix10473 (.Y (nx10474), .A (nx214)) ;
    inv02 ix10475 (.Y (nx10476), .A (nx214)) ;
    inv02 ix10477 (.Y (nx10478), .A (nx222)) ;
    inv02 ix10479 (.Y (nx10480), .A (nx222)) ;
    inv02 ix10481 (.Y (nx10482), .A (nx226)) ;
    inv02 ix10483 (.Y (nx10484), .A (nx226)) ;
    inv02 ix10485 (.Y (nx10486), .A (nx230)) ;
    inv02 ix10487 (.Y (nx10488), .A (nx230)) ;
    nor02ii ix8951 (.Y (sel_que_0), .A0 (nx6829), .A1 (nx6885)) ;
    nor02ii ix8961 (.Y (sel_que_1), .A0 (nx6839), .A1 (nx6885)) ;
    nor02ii ix8971 (.Y (sel_que_2), .A0 (nx6843), .A1 (nx6885)) ;
    nor02ii ix8979 (.Y (sel_que_3), .A0 (nx6847), .A1 (nx6885)) ;
    nor02ii ix8987 (.Y (sel_que_4), .A0 (nx6829), .A1 (nx6905)) ;
    nor02ii ix8991 (.Y (sel_que_5), .A0 (nx6839), .A1 (nx6905)) ;
    nor02ii ix8995 (.Y (sel_que_6), .A0 (nx6843), .A1 (nx6905)) ;
    nor02ii ix8999 (.Y (sel_que_7), .A0 (nx6847), .A1 (nx6905)) ;
    nor02ii ix9007 (.Y (sel_que_8), .A0 (nx6829), .A1 (nx6915)) ;
    nor02ii ix9011 (.Y (sel_que_9), .A0 (nx6839), .A1 (nx6915)) ;
    nor02ii ix9015 (.Y (sel_que_10), .A0 (nx6843), .A1 (nx6915)) ;
    nor02ii ix9019 (.Y (sel_que_11), .A0 (nx6847), .A1 (nx6915)) ;
    nor02ii ix9053 (.Y (sel_que_17), .A0 (nx6893), .A1 (nx6885)) ;
    nor02ii ix9063 (.Y (sel_que_18), .A0 (nx6897), .A1 (nx6885)) ;
    nor02ii ix9071 (.Y (sel_que_19), .A0 (nx6901), .A1 (nx6885)) ;
    nor02ii ix6906 (.Y (nx6905), .A0 (cache_in_sel[3]), .A1 (cache_in_sel[2])) ;
    nor02ii ix9079 (.Y (sel_que_21), .A0 (nx6893), .A1 (nx6905)) ;
    nor02ii ix9083 (.Y (sel_que_22), .A0 (nx6897), .A1 (nx6905)) ;
    nor02ii ix9087 (.Y (sel_que_23), .A0 (nx6901), .A1 (nx6905)) ;
    nor02ii ix6916 (.Y (nx6915), .A0 (cache_in_sel[2]), .A1 (cache_in_sel[3])) ;
    nor02ii ix9095 (.Y (sel_que_25), .A0 (nx6893), .A1 (nx6915)) ;
    nor02ii ix9099 (.Y (sel_que_26), .A0 (nx6897), .A1 (nx6915)) ;
    nor02ii ix9103 (.Y (sel_que_27), .A0 (nx6901), .A1 (nx6915)) ;
    nor02ii ix223 (.Y (nx222), .A0 (nx6931), .A1 (nx62)) ;
    nor02ii ix231 (.Y (nx230), .A0 (nx6945), .A1 (nx88)) ;
    nor02ii ix207 (.Y (nx206), .A0 (nx10374), .A1 (nx28)) ;
    nor02ii ix123 (.Y (nx122), .A0 (nx10374), .A1 (nx62)) ;
    nor02ii ix65 (.Y (nx64), .A0 (nx6949), .A1 (nx62)) ;
    nor02ii ix49 (.Y (nx48), .A0 (nx6949), .A1 (nx28)) ;
    nor02ii ix31 (.Y (nx30), .A0 (nx6931), .A1 (nx28)) ;
    inv02 ix10493 (.Y (nx10494), .A (nx6937)) ;
    inv02 ix10495 (.Y (nx10496), .A (nx6937)) ;
    inv02 ix10497 (.Y (nx10498), .A (nx6939)) ;
    inv02 ix10499 (.Y (nx10500), .A (nx6939)) ;
    inv01 ix10501 (.Y (nx10502), .A (nx6961)) ;
    inv01 ix10503 (.Y (nx10504), .A (nx6961)) ;
    inv02 ix10505 (.Y (nx10506), .A (nx6833)) ;
    inv02 ix10507 (.Y (nx10508), .A (nx6835)) ;
    inv01 ix10509 (.Y (nx10510), .A (in_word[15])) ;
    inv01 ix10511 (.Y (nx10512), .A (nx10510)) ;
    inv01 ix10513 (.Y (nx10514), .A (nx10510)) ;
    inv01 ix10515 (.Y (nx10516), .A (nx10510)) ;
    inv01 ix10517 (.Y (nx10518), .A (nx10510)) ;
    inv01 ix10519 (.Y (nx10520), .A (in_word[14])) ;
    inv01 ix10521 (.Y (nx10522), .A (nx10520)) ;
    inv01 ix10523 (.Y (nx10524), .A (nx10520)) ;
    inv01 ix10525 (.Y (nx10526), .A (nx10520)) ;
    inv01 ix10527 (.Y (nx10528), .A (nx10520)) ;
    inv01 ix10529 (.Y (nx10530), .A (in_word[13])) ;
    inv01 ix10531 (.Y (nx10532), .A (nx10530)) ;
    inv01 ix10533 (.Y (nx10534), .A (nx10530)) ;
    inv01 ix10535 (.Y (nx10536), .A (nx10530)) ;
    inv01 ix10537 (.Y (nx10538), .A (nx10530)) ;
    inv01 ix10539 (.Y (nx10540), .A (in_word[12])) ;
    inv01 ix10541 (.Y (nx10542), .A (nx10540)) ;
    inv01 ix10543 (.Y (nx10544), .A (nx10540)) ;
    inv01 ix10545 (.Y (nx10546), .A (nx10540)) ;
    inv01 ix10547 (.Y (nx10548), .A (nx10540)) ;
    inv01 ix10549 (.Y (nx10550), .A (in_word[11])) ;
    inv01 ix10551 (.Y (nx10552), .A (nx10550)) ;
    inv01 ix10553 (.Y (nx10554), .A (nx10550)) ;
    inv01 ix10555 (.Y (nx10556), .A (nx10550)) ;
    inv01 ix10557 (.Y (nx10558), .A (nx10550)) ;
    inv01 ix10559 (.Y (nx10560), .A (in_word[10])) ;
    inv01 ix10561 (.Y (nx10562), .A (nx10560)) ;
    inv01 ix10563 (.Y (nx10564), .A (nx10560)) ;
    inv01 ix10565 (.Y (nx10566), .A (nx10560)) ;
    inv01 ix10567 (.Y (nx10568), .A (nx10560)) ;
    inv01 ix10569 (.Y (nx10570), .A (in_word[9])) ;
    inv01 ix10571 (.Y (nx10572), .A (nx10570)) ;
    inv01 ix10573 (.Y (nx10574), .A (nx10570)) ;
    inv01 ix10575 (.Y (nx10576), .A (nx10570)) ;
    inv01 ix10577 (.Y (nx10578), .A (nx10570)) ;
    inv01 ix10579 (.Y (nx10580), .A (in_word[8])) ;
    inv01 ix10581 (.Y (nx10582), .A (nx10580)) ;
    inv01 ix10583 (.Y (nx10584), .A (nx10580)) ;
    inv01 ix10585 (.Y (nx10586), .A (nx10580)) ;
    inv01 ix10587 (.Y (nx10588), .A (nx10580)) ;
    inv01 ix10589 (.Y (nx10590), .A (in_word[7])) ;
    inv01 ix10591 (.Y (nx10592), .A (nx10590)) ;
    inv01 ix10593 (.Y (nx10594), .A (nx10590)) ;
    inv01 ix10595 (.Y (nx10596), .A (nx10590)) ;
    inv01 ix10597 (.Y (nx10598), .A (nx10590)) ;
    inv01 ix10599 (.Y (nx10600), .A (in_word[6])) ;
    inv01 ix10601 (.Y (nx10602), .A (nx10600)) ;
    inv01 ix10603 (.Y (nx10604), .A (nx10600)) ;
    inv01 ix10605 (.Y (nx10606), .A (nx10600)) ;
    inv01 ix10607 (.Y (nx10608), .A (nx10600)) ;
    inv01 ix10609 (.Y (nx10610), .A (in_word[5])) ;
    inv01 ix10611 (.Y (nx10612), .A (nx10610)) ;
    inv01 ix10613 (.Y (nx10614), .A (nx10610)) ;
    inv01 ix10615 (.Y (nx10616), .A (nx10610)) ;
    inv01 ix10617 (.Y (nx10618), .A (nx10610)) ;
    inv01 ix10619 (.Y (nx10620), .A (in_word[4])) ;
    inv01 ix10621 (.Y (nx10622), .A (nx10620)) ;
    inv01 ix10623 (.Y (nx10624), .A (nx10620)) ;
    inv01 ix10625 (.Y (nx10626), .A (nx10620)) ;
    inv01 ix10627 (.Y (nx10628), .A (nx10620)) ;
    inv01 ix10629 (.Y (nx10630), .A (in_word[3])) ;
    inv01 ix10631 (.Y (nx10632), .A (nx10630)) ;
    inv01 ix10633 (.Y (nx10634), .A (nx10630)) ;
    inv01 ix10635 (.Y (nx10636), .A (nx10630)) ;
    inv01 ix10637 (.Y (nx10638), .A (nx10630)) ;
    inv01 ix10639 (.Y (nx10640), .A (in_word[2])) ;
    inv01 ix10641 (.Y (nx10642), .A (nx10640)) ;
    inv01 ix10643 (.Y (nx10644), .A (nx10640)) ;
    inv01 ix10645 (.Y (nx10646), .A (nx10640)) ;
    inv01 ix10647 (.Y (nx10648), .A (nx10640)) ;
    inv01 ix10649 (.Y (nx10650), .A (in_word[1])) ;
    inv01 ix10651 (.Y (nx10652), .A (nx10650)) ;
    inv01 ix10653 (.Y (nx10654), .A (nx10650)) ;
    inv01 ix10655 (.Y (nx10656), .A (nx10650)) ;
    inv01 ix10657 (.Y (nx10658), .A (nx10650)) ;
    inv01 ix10659 (.Y (nx10660), .A (in_word[0])) ;
    inv01 ix10661 (.Y (nx10662), .A (nx10660)) ;
    inv01 ix10663 (.Y (nx10664), .A (nx10660)) ;
    inv01 ix10665 (.Y (nx10666), .A (nx10660)) ;
    inv01 ix10667 (.Y (nx10668), .A (nx10660)) ;
    inv02 ix10689 (.Y (nx10690), .A (nx10742)) ;
    inv02 ix10691 (.Y (nx10692), .A (nx10742)) ;
    inv02 ix10693 (.Y (nx10694), .A (nx10742)) ;
    inv02 ix10695 (.Y (nx10696), .A (nx10742)) ;
    inv02 ix10697 (.Y (nx10698), .A (nx10742)) ;
    inv02 ix10699 (.Y (nx10700), .A (nx10742)) ;
    inv02 ix10701 (.Y (nx10702), .A (nx10742)) ;
    inv02 ix10703 (.Y (nx10704), .A (nx10744)) ;
    inv02 ix10705 (.Y (nx10706), .A (nx10744)) ;
    inv02 ix10707 (.Y (nx10708), .A (nx10744)) ;
    inv02 ix10709 (.Y (nx10710), .A (nx10744)) ;
    inv02 ix10711 (.Y (nx10712), .A (nx10744)) ;
    inv02 ix10713 (.Y (nx10714), .A (nx10746)) ;
    inv02 ix10715 (.Y (nx10716), .A (nx10746)) ;
    inv02 ix10717 (.Y (nx10718), .A (nx10746)) ;
    inv02 ix10719 (.Y (nx10720), .A (nx10746)) ;
    inv02 ix10721 (.Y (nx10722), .A (nx10746)) ;
    inv02 ix10723 (.Y (nx10724), .A (nx10746)) ;
    inv02 ix10725 (.Y (nx10726), .A (nx10746)) ;
    inv02 ix10727 (.Y (nx10728), .A (nx10748)) ;
    inv02 ix10729 (.Y (nx10730), .A (nx10748)) ;
    inv02 ix10731 (.Y (nx10732), .A (nx10748)) ;
    inv02 ix10733 (.Y (nx10734), .A (nx10748)) ;
    inv02 ix10735 (.Y (nx10736), .A (nx10748)) ;
    inv02 ix10741 (.Y (nx10742), .A (reset)) ;
    inv02 ix10743 (.Y (nx10744), .A (reset)) ;
    inv02 ix10745 (.Y (nx10746), .A (clk)) ;
    inv02 ix10747 (.Y (nx10748), .A (clk)) ;
endmodule


module Queue_5 ( d, q_0__15, q_0__14, q_0__13, q_0__12, q_0__11, q_0__10, q_0__9, 
                 q_0__8, q_0__7, q_0__6, q_0__5, q_0__4, q_0__3, q_0__2, q_0__1, 
                 q_0__0, q_1__15, q_1__14, q_1__13, q_1__12, q_1__11, q_1__10, 
                 q_1__9, q_1__8, q_1__7, q_1__6, q_1__5, q_1__4, q_1__3, q_1__2, 
                 q_1__1, q_1__0, q_2__15, q_2__14, q_2__13, q_2__12, q_2__11, 
                 q_2__10, q_2__9, q_2__8, q_2__7, q_2__6, q_2__5, q_2__4, q_2__3, 
                 q_2__2, q_2__1, q_2__0, q_3__15, q_3__14, q_3__13, q_3__12, 
                 q_3__11, q_3__10, q_3__9, q_3__8, q_3__7, q_3__6, q_3__5, 
                 q_3__4, q_3__3, q_3__2, q_3__1, q_3__0, q_4__15, q_4__14, 
                 q_4__13, q_4__12, q_4__11, q_4__10, q_4__9, q_4__8, q_4__7, 
                 q_4__6, q_4__5, q_4__4, q_4__3, q_4__2, q_4__1, q_4__0, clk, 
                 load, reset ) ;

    input [15:0]d ;
    output q_0__15 ;
    output q_0__14 ;
    output q_0__13 ;
    output q_0__12 ;
    output q_0__11 ;
    output q_0__10 ;
    output q_0__9 ;
    output q_0__8 ;
    output q_0__7 ;
    output q_0__6 ;
    output q_0__5 ;
    output q_0__4 ;
    output q_0__3 ;
    output q_0__2 ;
    output q_0__1 ;
    output q_0__0 ;
    output q_1__15 ;
    output q_1__14 ;
    output q_1__13 ;
    output q_1__12 ;
    output q_1__11 ;
    output q_1__10 ;
    output q_1__9 ;
    output q_1__8 ;
    output q_1__7 ;
    output q_1__6 ;
    output q_1__5 ;
    output q_1__4 ;
    output q_1__3 ;
    output q_1__2 ;
    output q_1__1 ;
    output q_1__0 ;
    output q_2__15 ;
    output q_2__14 ;
    output q_2__13 ;
    output q_2__12 ;
    output q_2__11 ;
    output q_2__10 ;
    output q_2__9 ;
    output q_2__8 ;
    output q_2__7 ;
    output q_2__6 ;
    output q_2__5 ;
    output q_2__4 ;
    output q_2__3 ;
    output q_2__2 ;
    output q_2__1 ;
    output q_2__0 ;
    output q_3__15 ;
    output q_3__14 ;
    output q_3__13 ;
    output q_3__12 ;
    output q_3__11 ;
    output q_3__10 ;
    output q_3__9 ;
    output q_3__8 ;
    output q_3__7 ;
    output q_3__6 ;
    output q_3__5 ;
    output q_3__4 ;
    output q_3__3 ;
    output q_3__2 ;
    output q_3__1 ;
    output q_3__0 ;
    output q_4__15 ;
    output q_4__14 ;
    output q_4__13 ;
    output q_4__12 ;
    output q_4__11 ;
    output q_4__10 ;
    output q_4__9 ;
    output q_4__8 ;
    output q_4__7 ;
    output q_4__6 ;
    output q_4__5 ;
    output q_4__4 ;
    output q_4__3 ;
    output q_4__2 ;
    output q_4__1 ;
    output q_4__0 ;
    input clk ;
    input load ;
    input reset ;

    wire nx393, nx403, nx413, nx423, nx433, nx443, nx453, nx463, nx473, nx483, 
         nx493, nx503, nx513, nx523, nx533, nx543, nx553, nx563, nx573, nx583, 
         nx593, nx603, nx613, nx623, nx633, nx643, nx653, nx663, nx673, nx683, 
         nx693, nx703, nx713, nx723, nx733, nx743, nx753, nx763, nx773, nx783, 
         nx793, nx803, nx813, nx823, nx833, nx843, nx853, nx863, nx873, nx883, 
         nx893, nx903, nx913, nx923, nx933, nx943, nx953, nx963, nx973, nx983, 
         nx993, nx1003, nx1013, nx1023, nx1033, nx1043, nx1053, nx1063, nx1073, 
         nx1083, nx1093, nx1103, nx1113, nx1123, nx1133, nx1143, nx1153, nx1163, 
         nx1173, nx1183, nx1440, nx1442, nx1444, nx1446, nx1448, nx1450, nx1452, 
         nx1454, nx1456, nx1458, nx1460, nx1462, nx1466, nx1468, nx1470, nx1472, 
         nx1474, nx1476, nx1478, nx1480, nx1482, nx1484, nx1486, nx1488, nx1492, 
         nx1494, nx1496, nx1498, nx1500, nx1502, nx1504, nx1506, nx1508, nx1510, 
         nx1512, nx1514, nx1516, nx1518, nx1520, nx1522, nx1524, nx1526;
    wire [79:0] \$dummy ;




    dffr gen_regs_4_regi_reg_q_0 (.Q (q_4__0), .QB (\$dummy [0]), .D (nx433), .CLK (
         nx1492), .R (nx1466)) ;
    mux21_ni ix434 (.Y (nx433), .A0 (q_4__0), .A1 (q_3__0), .S0 (nx1440)) ;
    dffr gen_regs_3_regi_reg_q_0 (.Q (q_3__0), .QB (\$dummy [1]), .D (nx423), .CLK (
         nx1492), .R (nx1466)) ;
    mux21_ni ix424 (.Y (nx423), .A0 (q_3__0), .A1 (q_2__0), .S0 (nx1440)) ;
    dffr gen_regs_2_regi_reg_q_0 (.Q (q_2__0), .QB (\$dummy [2]), .D (nx413), .CLK (
         nx1492), .R (nx1466)) ;
    mux21_ni ix414 (.Y (nx413), .A0 (q_2__0), .A1 (q_1__0), .S0 (nx1440)) ;
    dffr gen_regs_1_regi_reg_q_0 (.Q (q_1__0), .QB (\$dummy [3]), .D (nx403), .CLK (
         nx1492), .R (nx1466)) ;
    mux21_ni ix404 (.Y (nx403), .A0 (q_1__0), .A1 (q_0__0), .S0 (nx1440)) ;
    dffr reg0_reg_q_0 (.Q (q_0__0), .QB (\$dummy [4]), .D (nx393), .CLK (nx1492)
         , .R (nx1466)) ;
    mux21_ni ix394 (.Y (nx393), .A0 (q_0__0), .A1 (d[0]), .S0 (nx1440)) ;
    dffr gen_regs_4_regi_reg_q_1 (.Q (q_4__1), .QB (\$dummy [5]), .D (nx483), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix484 (.Y (nx483), .A0 (q_4__1), .A1 (q_3__1), .S0 (nx1442)) ;
    dffr gen_regs_3_regi_reg_q_1 (.Q (q_3__1), .QB (\$dummy [6]), .D (nx473), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix474 (.Y (nx473), .A0 (q_3__1), .A1 (q_2__1), .S0 (nx1442)) ;
    dffr gen_regs_2_regi_reg_q_1 (.Q (q_2__1), .QB (\$dummy [7]), .D (nx463), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix464 (.Y (nx463), .A0 (q_2__1), .A1 (q_1__1), .S0 (nx1442)) ;
    dffr gen_regs_1_regi_reg_q_1 (.Q (q_1__1), .QB (\$dummy [8]), .D (nx453), .CLK (
         nx1492), .R (nx1466)) ;
    mux21_ni ix454 (.Y (nx453), .A0 (q_1__1), .A1 (q_0__1), .S0 (nx1440)) ;
    dffr reg0_reg_q_1 (.Q (q_0__1), .QB (\$dummy [9]), .D (nx443), .CLK (nx1492)
         , .R (nx1466)) ;
    mux21_ni ix444 (.Y (nx443), .A0 (q_0__1), .A1 (d[1]), .S0 (nx1440)) ;
    dffr gen_regs_4_regi_reg_q_2 (.Q (q_4__2), .QB (\$dummy [10]), .D (nx533), .CLK (
         nx1496), .R (nx1470)) ;
    mux21_ni ix534 (.Y (nx533), .A0 (q_4__2), .A1 (q_3__2), .S0 (nx1444)) ;
    dffr gen_regs_3_regi_reg_q_2 (.Q (q_3__2), .QB (\$dummy [11]), .D (nx523), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix524 (.Y (nx523), .A0 (q_3__2), .A1 (q_2__2), .S0 (nx1442)) ;
    dffr gen_regs_2_regi_reg_q_2 (.Q (q_2__2), .QB (\$dummy [12]), .D (nx513), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix514 (.Y (nx513), .A0 (q_2__2), .A1 (q_1__2), .S0 (nx1442)) ;
    dffr gen_regs_1_regi_reg_q_2 (.Q (q_1__2), .QB (\$dummy [13]), .D (nx503), .CLK (
         nx1494), .R (nx1468)) ;
    mux21_ni ix504 (.Y (nx503), .A0 (q_1__2), .A1 (q_0__2), .S0 (nx1442)) ;
    dffr reg0_reg_q_2 (.Q (q_0__2), .QB (\$dummy [14]), .D (nx493), .CLK (nx1494
         ), .R (nx1468)) ;
    mux21_ni ix494 (.Y (nx493), .A0 (q_0__2), .A1 (d[2]), .S0 (nx1442)) ;
    dffr gen_regs_4_regi_reg_q_3 (.Q (q_4__3), .QB (\$dummy [15]), .D (nx583), .CLK (
         nx1496), .R (nx1470)) ;
    mux21_ni ix584 (.Y (nx583), .A0 (q_4__3), .A1 (q_3__3), .S0 (nx1444)) ;
    dffr gen_regs_3_regi_reg_q_3 (.Q (q_3__3), .QB (\$dummy [16]), .D (nx573), .CLK (
         nx1496), .R (nx1470)) ;
    mux21_ni ix574 (.Y (nx573), .A0 (q_3__3), .A1 (q_2__3), .S0 (nx1444)) ;
    dffr gen_regs_2_regi_reg_q_3 (.Q (q_2__3), .QB (\$dummy [17]), .D (nx563), .CLK (
         nx1496), .R (nx1470)) ;
    mux21_ni ix564 (.Y (nx563), .A0 (q_2__3), .A1 (q_1__3), .S0 (nx1444)) ;
    dffr gen_regs_1_regi_reg_q_3 (.Q (q_1__3), .QB (\$dummy [18]), .D (nx553), .CLK (
         nx1496), .R (nx1470)) ;
    mux21_ni ix554 (.Y (nx553), .A0 (q_1__3), .A1 (q_0__3), .S0 (nx1444)) ;
    dffr reg0_reg_q_3 (.Q (q_0__3), .QB (\$dummy [19]), .D (nx543), .CLK (nx1496
         ), .R (nx1470)) ;
    mux21_ni ix544 (.Y (nx543), .A0 (q_0__3), .A1 (d[3]), .S0 (nx1444)) ;
    dffr gen_regs_4_regi_reg_q_4 (.Q (q_4__4), .QB (\$dummy [20]), .D (nx633), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix634 (.Y (nx633), .A0 (q_4__4), .A1 (q_3__4), .S0 (nx1446)) ;
    dffr gen_regs_3_regi_reg_q_4 (.Q (q_3__4), .QB (\$dummy [21]), .D (nx623), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix624 (.Y (nx623), .A0 (q_3__4), .A1 (q_2__4), .S0 (nx1446)) ;
    dffr gen_regs_2_regi_reg_q_4 (.Q (q_2__4), .QB (\$dummy [22]), .D (nx613), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix614 (.Y (nx613), .A0 (q_2__4), .A1 (q_1__4), .S0 (nx1446)) ;
    dffr gen_regs_1_regi_reg_q_4 (.Q (q_1__4), .QB (\$dummy [23]), .D (nx603), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix604 (.Y (nx603), .A0 (q_1__4), .A1 (q_0__4), .S0 (nx1446)) ;
    dffr reg0_reg_q_4 (.Q (q_0__4), .QB (\$dummy [24]), .D (nx593), .CLK (nx1496
         ), .R (nx1470)) ;
    mux21_ni ix594 (.Y (nx593), .A0 (q_0__4), .A1 (d[4]), .S0 (nx1444)) ;
    dffr gen_regs_4_regi_reg_q_5 (.Q (q_4__5), .QB (\$dummy [25]), .D (nx683), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix684 (.Y (nx683), .A0 (q_4__5), .A1 (q_3__5), .S0 (nx1448)) ;
    dffr gen_regs_3_regi_reg_q_5 (.Q (q_3__5), .QB (\$dummy [26]), .D (nx673), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix674 (.Y (nx673), .A0 (q_3__5), .A1 (q_2__5), .S0 (nx1448)) ;
    dffr gen_regs_2_regi_reg_q_5 (.Q (q_2__5), .QB (\$dummy [27]), .D (nx663), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix664 (.Y (nx663), .A0 (q_2__5), .A1 (q_1__5), .S0 (nx1446)) ;
    dffr gen_regs_1_regi_reg_q_5 (.Q (q_1__5), .QB (\$dummy [28]), .D (nx653), .CLK (
         nx1498), .R (nx1472)) ;
    mux21_ni ix654 (.Y (nx653), .A0 (q_1__5), .A1 (q_0__5), .S0 (nx1446)) ;
    dffr reg0_reg_q_5 (.Q (q_0__5), .QB (\$dummy [29]), .D (nx643), .CLK (nx1498
         ), .R (nx1472)) ;
    mux21_ni ix644 (.Y (nx643), .A0 (q_0__5), .A1 (d[5]), .S0 (nx1446)) ;
    dffr gen_regs_4_regi_reg_q_6 (.Q (q_4__6), .QB (\$dummy [30]), .D (nx733), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix734 (.Y (nx733), .A0 (q_4__6), .A1 (q_3__6), .S0 (nx1448)) ;
    dffr gen_regs_3_regi_reg_q_6 (.Q (q_3__6), .QB (\$dummy [31]), .D (nx723), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix724 (.Y (nx723), .A0 (q_3__6), .A1 (q_2__6), .S0 (nx1448)) ;
    dffr gen_regs_2_regi_reg_q_6 (.Q (q_2__6), .QB (\$dummy [32]), .D (nx713), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix714 (.Y (nx713), .A0 (q_2__6), .A1 (q_1__6), .S0 (nx1448)) ;
    dffr gen_regs_1_regi_reg_q_6 (.Q (q_1__6), .QB (\$dummy [33]), .D (nx703), .CLK (
         nx1500), .R (nx1474)) ;
    mux21_ni ix704 (.Y (nx703), .A0 (q_1__6), .A1 (q_0__6), .S0 (nx1448)) ;
    dffr reg0_reg_q_6 (.Q (q_0__6), .QB (\$dummy [34]), .D (nx693), .CLK (nx1500
         ), .R (nx1474)) ;
    mux21_ni ix694 (.Y (nx693), .A0 (q_0__6), .A1 (d[6]), .S0 (nx1448)) ;
    dffr gen_regs_4_regi_reg_q_7 (.Q (q_4__7), .QB (\$dummy [35]), .D (nx783), .CLK (
         nx1502), .R (nx1476)) ;
    mux21_ni ix784 (.Y (nx783), .A0 (q_4__7), .A1 (q_3__7), .S0 (nx1450)) ;
    dffr gen_regs_3_regi_reg_q_7 (.Q (q_3__7), .QB (\$dummy [36]), .D (nx773), .CLK (
         nx1502), .R (nx1476)) ;
    mux21_ni ix774 (.Y (nx773), .A0 (q_3__7), .A1 (q_2__7), .S0 (nx1450)) ;
    dffr gen_regs_2_regi_reg_q_7 (.Q (q_2__7), .QB (\$dummy [37]), .D (nx763), .CLK (
         nx1502), .R (nx1476)) ;
    mux21_ni ix764 (.Y (nx763), .A0 (q_2__7), .A1 (q_1__7), .S0 (nx1450)) ;
    dffr gen_regs_1_regi_reg_q_7 (.Q (q_1__7), .QB (\$dummy [38]), .D (nx753), .CLK (
         nx1502), .R (nx1476)) ;
    mux21_ni ix754 (.Y (nx753), .A0 (q_1__7), .A1 (q_0__7), .S0 (nx1450)) ;
    dffr reg0_reg_q_7 (.Q (q_0__7), .QB (\$dummy [39]), .D (nx743), .CLK (nx1502
         ), .R (nx1476)) ;
    mux21_ni ix744 (.Y (nx743), .A0 (q_0__7), .A1 (d[7]), .S0 (nx1450)) ;
    dffr gen_regs_4_regi_reg_q_8 (.Q (q_4__8), .QB (\$dummy [40]), .D (nx833), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix834 (.Y (nx833), .A0 (q_4__8), .A1 (q_3__8), .S0 (nx1452)) ;
    dffr gen_regs_3_regi_reg_q_8 (.Q (q_3__8), .QB (\$dummy [41]), .D (nx823), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix824 (.Y (nx823), .A0 (q_3__8), .A1 (q_2__8), .S0 (nx1452)) ;
    dffr gen_regs_2_regi_reg_q_8 (.Q (q_2__8), .QB (\$dummy [42]), .D (nx813), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix814 (.Y (nx813), .A0 (q_2__8), .A1 (q_1__8), .S0 (nx1452)) ;
    dffr gen_regs_1_regi_reg_q_8 (.Q (q_1__8), .QB (\$dummy [43]), .D (nx803), .CLK (
         nx1502), .R (nx1476)) ;
    mux21_ni ix804 (.Y (nx803), .A0 (q_1__8), .A1 (q_0__8), .S0 (nx1450)) ;
    dffr reg0_reg_q_8 (.Q (q_0__8), .QB (\$dummy [44]), .D (nx793), .CLK (nx1502
         ), .R (nx1476)) ;
    mux21_ni ix794 (.Y (nx793), .A0 (q_0__8), .A1 (d[8]), .S0 (nx1450)) ;
    dffr gen_regs_4_regi_reg_q_9 (.Q (q_4__9), .QB (\$dummy [45]), .D (nx883), .CLK (
         nx1506), .R (nx1480)) ;
    mux21_ni ix884 (.Y (nx883), .A0 (q_4__9), .A1 (q_3__9), .S0 (nx1454)) ;
    dffr gen_regs_3_regi_reg_q_9 (.Q (q_3__9), .QB (\$dummy [46]), .D (nx873), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix874 (.Y (nx873), .A0 (q_3__9), .A1 (q_2__9), .S0 (nx1452)) ;
    dffr gen_regs_2_regi_reg_q_9 (.Q (q_2__9), .QB (\$dummy [47]), .D (nx863), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix864 (.Y (nx863), .A0 (q_2__9), .A1 (q_1__9), .S0 (nx1452)) ;
    dffr gen_regs_1_regi_reg_q_9 (.Q (q_1__9), .QB (\$dummy [48]), .D (nx853), .CLK (
         nx1504), .R (nx1478)) ;
    mux21_ni ix854 (.Y (nx853), .A0 (q_1__9), .A1 (q_0__9), .S0 (nx1452)) ;
    dffr reg0_reg_q_9 (.Q (q_0__9), .QB (\$dummy [49]), .D (nx843), .CLK (nx1504
         ), .R (nx1478)) ;
    mux21_ni ix844 (.Y (nx843), .A0 (q_0__9), .A1 (d[9]), .S0 (nx1452)) ;
    dffr gen_regs_4_regi_reg_q_10 (.Q (q_4__10), .QB (\$dummy [50]), .D (nx933)
         , .CLK (nx1506), .R (nx1480)) ;
    mux21_ni ix934 (.Y (nx933), .A0 (q_4__10), .A1 (q_3__10), .S0 (nx1454)) ;
    dffr gen_regs_3_regi_reg_q_10 (.Q (q_3__10), .QB (\$dummy [51]), .D (nx923)
         , .CLK (nx1506), .R (nx1480)) ;
    mux21_ni ix924 (.Y (nx923), .A0 (q_3__10), .A1 (q_2__10), .S0 (nx1454)) ;
    dffr gen_regs_2_regi_reg_q_10 (.Q (q_2__10), .QB (\$dummy [52]), .D (nx913)
         , .CLK (nx1506), .R (nx1480)) ;
    mux21_ni ix914 (.Y (nx913), .A0 (q_2__10), .A1 (q_1__10), .S0 (nx1454)) ;
    dffr gen_regs_1_regi_reg_q_10 (.Q (q_1__10), .QB (\$dummy [53]), .D (nx903)
         , .CLK (nx1506), .R (nx1480)) ;
    mux21_ni ix904 (.Y (nx903), .A0 (q_1__10), .A1 (q_0__10), .S0 (nx1454)) ;
    dffr reg0_reg_q_10 (.Q (q_0__10), .QB (\$dummy [54]), .D (nx893), .CLK (
         nx1506), .R (nx1480)) ;
    mux21_ni ix894 (.Y (nx893), .A0 (q_0__10), .A1 (d[10]), .S0 (nx1454)) ;
    dffr gen_regs_4_regi_reg_q_11 (.Q (q_4__11), .QB (\$dummy [55]), .D (nx983)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix984 (.Y (nx983), .A0 (q_4__11), .A1 (q_3__11), .S0 (nx1456)) ;
    dffr gen_regs_3_regi_reg_q_11 (.Q (q_3__11), .QB (\$dummy [56]), .D (nx973)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix974 (.Y (nx973), .A0 (q_3__11), .A1 (q_2__11), .S0 (nx1456)) ;
    dffr gen_regs_2_regi_reg_q_11 (.Q (q_2__11), .QB (\$dummy [57]), .D (nx963)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix964 (.Y (nx963), .A0 (q_2__11), .A1 (q_1__11), .S0 (nx1456)) ;
    dffr gen_regs_1_regi_reg_q_11 (.Q (q_1__11), .QB (\$dummy [58]), .D (nx953)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix954 (.Y (nx953), .A0 (q_1__11), .A1 (q_0__11), .S0 (nx1456)) ;
    dffr reg0_reg_q_11 (.Q (q_0__11), .QB (\$dummy [59]), .D (nx943), .CLK (
         nx1506), .R (nx1480)) ;
    mux21_ni ix944 (.Y (nx943), .A0 (q_0__11), .A1 (d[11]), .S0 (nx1454)) ;
    dffr gen_regs_4_regi_reg_q_12 (.Q (q_4__12), .QB (\$dummy [60]), .D (nx1033)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1034 (.Y (nx1033), .A0 (q_4__12), .A1 (q_3__12), .S0 (nx1458)) ;
    dffr gen_regs_3_regi_reg_q_12 (.Q (q_3__12), .QB (\$dummy [61]), .D (nx1023)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1024 (.Y (nx1023), .A0 (q_3__12), .A1 (q_2__12), .S0 (nx1458)) ;
    dffr gen_regs_2_regi_reg_q_12 (.Q (q_2__12), .QB (\$dummy [62]), .D (nx1013)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix1014 (.Y (nx1013), .A0 (q_2__12), .A1 (q_1__12), .S0 (nx1456)) ;
    dffr gen_regs_1_regi_reg_q_12 (.Q (q_1__12), .QB (\$dummy [63]), .D (nx1003)
         , .CLK (nx1508), .R (nx1482)) ;
    mux21_ni ix1004 (.Y (nx1003), .A0 (q_1__12), .A1 (q_0__12), .S0 (nx1456)) ;
    dffr reg0_reg_q_12 (.Q (q_0__12), .QB (\$dummy [64]), .D (nx993), .CLK (
         nx1508), .R (nx1482)) ;
    mux21_ni ix994 (.Y (nx993), .A0 (q_0__12), .A1 (d[12]), .S0 (nx1456)) ;
    dffr gen_regs_4_regi_reg_q_13 (.Q (q_4__13), .QB (\$dummy [65]), .D (nx1083)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1084 (.Y (nx1083), .A0 (q_4__13), .A1 (q_3__13), .S0 (nx1458)) ;
    dffr gen_regs_3_regi_reg_q_13 (.Q (q_3__13), .QB (\$dummy [66]), .D (nx1073)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1074 (.Y (nx1073), .A0 (q_3__13), .A1 (q_2__13), .S0 (nx1458)) ;
    dffr gen_regs_2_regi_reg_q_13 (.Q (q_2__13), .QB (\$dummy [67]), .D (nx1063)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1064 (.Y (nx1063), .A0 (q_2__13), .A1 (q_1__13), .S0 (nx1458)) ;
    dffr gen_regs_1_regi_reg_q_13 (.Q (q_1__13), .QB (\$dummy [68]), .D (nx1053)
         , .CLK (nx1510), .R (nx1484)) ;
    mux21_ni ix1054 (.Y (nx1053), .A0 (q_1__13), .A1 (q_0__13), .S0 (nx1458)) ;
    dffr reg0_reg_q_13 (.Q (q_0__13), .QB (\$dummy [69]), .D (nx1043), .CLK (
         nx1510), .R (nx1484)) ;
    mux21_ni ix1044 (.Y (nx1043), .A0 (q_0__13), .A1 (d[13]), .S0 (nx1458)) ;
    dffr gen_regs_4_regi_reg_q_14 (.Q (q_4__14), .QB (\$dummy [70]), .D (nx1133)
         , .CLK (nx1512), .R (nx1486)) ;
    mux21_ni ix1134 (.Y (nx1133), .A0 (q_4__14), .A1 (q_3__14), .S0 (nx1460)) ;
    dffr gen_regs_3_regi_reg_q_14 (.Q (q_3__14), .QB (\$dummy [71]), .D (nx1123)
         , .CLK (nx1512), .R (nx1486)) ;
    mux21_ni ix1124 (.Y (nx1123), .A0 (q_3__14), .A1 (q_2__14), .S0 (nx1460)) ;
    dffr gen_regs_2_regi_reg_q_14 (.Q (q_2__14), .QB (\$dummy [72]), .D (nx1113)
         , .CLK (nx1512), .R (nx1486)) ;
    mux21_ni ix1114 (.Y (nx1113), .A0 (q_2__14), .A1 (q_1__14), .S0 (nx1460)) ;
    dffr gen_regs_1_regi_reg_q_14 (.Q (q_1__14), .QB (\$dummy [73]), .D (nx1103)
         , .CLK (nx1512), .R (nx1486)) ;
    mux21_ni ix1104 (.Y (nx1103), .A0 (q_1__14), .A1 (q_0__14), .S0 (nx1460)) ;
    dffr reg0_reg_q_14 (.Q (q_0__14), .QB (\$dummy [74]), .D (nx1093), .CLK (
         nx1512), .R (nx1486)) ;
    mux21_ni ix1094 (.Y (nx1093), .A0 (q_0__14), .A1 (d[14]), .S0 (nx1460)) ;
    dffr gen_regs_4_regi_reg_q_15 (.Q (q_4__15), .QB (\$dummy [75]), .D (nx1183)
         , .CLK (nx1514), .R (nx1488)) ;
    mux21_ni ix1184 (.Y (nx1183), .A0 (q_4__15), .A1 (q_3__15), .S0 (nx1462)) ;
    dffr gen_regs_3_regi_reg_q_15 (.Q (q_3__15), .QB (\$dummy [76]), .D (nx1173)
         , .CLK (nx1514), .R (nx1488)) ;
    mux21_ni ix1174 (.Y (nx1173), .A0 (q_3__15), .A1 (q_2__15), .S0 (nx1462)) ;
    dffr gen_regs_2_regi_reg_q_15 (.Q (q_2__15), .QB (\$dummy [77]), .D (nx1163)
         , .CLK (nx1514), .R (nx1488)) ;
    mux21_ni ix1164 (.Y (nx1163), .A0 (q_2__15), .A1 (q_1__15), .S0 (nx1462)) ;
    dffr gen_regs_1_regi_reg_q_15 (.Q (q_1__15), .QB (\$dummy [78]), .D (nx1153)
         , .CLK (nx1512), .R (nx1486)) ;
    mux21_ni ix1154 (.Y (nx1153), .A0 (q_1__15), .A1 (q_0__15), .S0 (nx1460)) ;
    dffr reg0_reg_q_15 (.Q (q_0__15), .QB (\$dummy [79]), .D (nx1143), .CLK (
         nx1512), .R (nx1486)) ;
    mux21_ni ix1144 (.Y (nx1143), .A0 (q_0__15), .A1 (d[15]), .S0 (nx1460)) ;
    inv02 ix1439 (.Y (nx1440), .A (nx1516)) ;
    inv02 ix1441 (.Y (nx1442), .A (nx1516)) ;
    inv02 ix1443 (.Y (nx1444), .A (nx1516)) ;
    inv02 ix1445 (.Y (nx1446), .A (nx1516)) ;
    inv02 ix1447 (.Y (nx1448), .A (nx1516)) ;
    inv02 ix1449 (.Y (nx1450), .A (nx1516)) ;
    inv02 ix1451 (.Y (nx1452), .A (nx1516)) ;
    inv02 ix1453 (.Y (nx1454), .A (nx1518)) ;
    inv02 ix1455 (.Y (nx1456), .A (nx1518)) ;
    inv02 ix1457 (.Y (nx1458), .A (nx1518)) ;
    inv02 ix1459 (.Y (nx1460), .A (nx1518)) ;
    inv02 ix1461 (.Y (nx1462), .A (nx1518)) ;
    inv02 ix1465 (.Y (nx1466), .A (nx1520)) ;
    inv02 ix1467 (.Y (nx1468), .A (nx1520)) ;
    inv02 ix1469 (.Y (nx1470), .A (nx1520)) ;
    inv02 ix1471 (.Y (nx1472), .A (nx1520)) ;
    inv02 ix1473 (.Y (nx1474), .A (nx1520)) ;
    inv02 ix1475 (.Y (nx1476), .A (nx1520)) ;
    inv02 ix1477 (.Y (nx1478), .A (nx1520)) ;
    inv02 ix1479 (.Y (nx1480), .A (nx1522)) ;
    inv02 ix1481 (.Y (nx1482), .A (nx1522)) ;
    inv02 ix1483 (.Y (nx1484), .A (nx1522)) ;
    inv02 ix1485 (.Y (nx1486), .A (nx1522)) ;
    inv02 ix1487 (.Y (nx1488), .A (nx1522)) ;
    inv02 ix1491 (.Y (nx1492), .A (nx1524)) ;
    inv02 ix1493 (.Y (nx1494), .A (nx1524)) ;
    inv02 ix1495 (.Y (nx1496), .A (nx1524)) ;
    inv02 ix1497 (.Y (nx1498), .A (nx1524)) ;
    inv02 ix1499 (.Y (nx1500), .A (nx1524)) ;
    inv02 ix1501 (.Y (nx1502), .A (nx1524)) ;
    inv02 ix1503 (.Y (nx1504), .A (nx1524)) ;
    inv02 ix1505 (.Y (nx1506), .A (nx1526)) ;
    inv02 ix1507 (.Y (nx1508), .A (nx1526)) ;
    inv02 ix1509 (.Y (nx1510), .A (nx1526)) ;
    inv02 ix1511 (.Y (nx1512), .A (nx1526)) ;
    inv02 ix1513 (.Y (nx1514), .A (nx1526)) ;
    inv02 ix1515 (.Y (nx1516), .A (load)) ;
    inv02 ix1517 (.Y (nx1518), .A (load)) ;
    inv02 ix1519 (.Y (nx1520), .A (reset)) ;
    inv02 ix1521 (.Y (nx1522), .A (reset)) ;
    inv02 ix1523 (.Y (nx1524), .A (clk)) ;
    inv02 ix1525 (.Y (nx1526), .A (clk)) ;
endmodule

