library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;

entity control_unit_test is
end control_unit_test;

architecture mixed of control_unit_test is
begin
end mixed;